module frisc (
	tin_pdata_8_8_, tin_pdata_0_0_, tin_pdata_7_7_, preset_0_0_, tin_pdata_2_2_, tin_pdata_9_9_, tin_pdata_1_1_, tin_pdata_4_4_, 
	pclk, pirq_0_0_, tin_pdata_10_10_, tin_pdata_3_3_, tin_pdata_6_6_, tin_pdata_15_15_, tin_pdata_11_11_, tin_pdata_14_14_, tin_pdata_12_12_, tin_pdata_5_5_, 
	preset, tin_pdata_13_13_, ppeakb_7_7_, ppeakp_12_12_, ppeakp_0_0_, ppeaka_7_7_, ppeaki_15_15_, ppeaki_11_11_, ppeaki_3_3_, paddress_3_3_, 
	pdata_8_8_, pdata_0_0_, ppeakb_14_14_, ppeakb_10_10_, ppeakb_8_8_, ppeakp_1_1_, ppeaka_14_14_, ppeaka_10_10_, ppeaka_8_8_, ppeaki_4_4_, 
	paddress_15_15_, paddress_11_11_, paddress_2_2_, ppeakb_9_9_, ppeakp_2_2_, ppeaka_9_9_, ppeaks_12_12_, ppeaks_0_0_, ppeaki_5_5_, paddress_5_5_, 
	pdata_7_7_, ppeakb_15_15_, ppeakp_3_3_, pwr_0_0_, ppeaks_1_1_, ppeaki_6_6_, paddress_4_4_, piack_0_0_, ppeakp_13_13_, ppeakp_4_4_, 
	ppeaka_15_15_, ppeaka_11_11_, ppeaks_2_2_, ppeaki_7_7_, paddress_10_10_, paddress_7_7_, pdata_2_2_, ppeakp_5_5_, ppeaks_13_13_, ppeaks_3_3_, 
	ppeaki_14_14_, ppeaki_10_10_, ppeaki_8_8_, paddress_6_6_, ppeakp_6_6_, ppeaks_4_4_, ppeaki_9_9_, paddress_9_9_, pdata_9_9_, pdata_1_1_, 
	ppeakb_11_11_, ppeakp_7_7_, ppeaks_5_5_, paddress_13_13_, paddress_8_8_, ppeakp_14_14_, ppeakp_10_10_, ppeakp_8_8_, ppeaks_6_6_, ppeaki_13_13_, 
	pdata_4_4_, ppeakb_0_0_, ppeakp_9_9_, ppeaka_0_0_, ppeaks_7_7_, ppeakb_1_1_, ppeaka_1_1_, ppeaks_10_10_, ppeaks_8_8_, pdata_10_10_, 
	pdata_3_3_, ppeakb_12_12_, ppeakb_2_2_, ppeaka_12_12_, ppeaka_2_2_, ppeaks_15_15_, ppeaks_9_9_, ppeakb_3_3_, ppeakp_15_15_, ppeakp_11_11_, 
	ppeaka_13_13_, ppeaka_3_3_, paddress_14_14_, paddress_12_12_, pdata_6_6_, ppeakb_13_13_, ppeakb_4_4_, pdn, ppeaka_4_4_, ppeaki_0_0_, 
	prd_0_0_, pdata_15_15_, pdata_11_11_, ppeakb_5_5_, ppeaka_5_5_, ppeaks_14_14_, ppeaki_1_1_, paddress_1_1_, pdata_14_14_, pdata_12_12_, 
	pdata_5_5_, ppeakb_6_6_, ppeaka_6_6_, ppeaks_11_11_, ppeaki_12_12_, ppeaki_2_2_, paddress_0_0_, pdata_13_13_);

input tin_pdata_8_8_;
input tin_pdata_0_0_;
input tin_pdata_7_7_;
input preset_0_0_;
input tin_pdata_2_2_;
input tin_pdata_9_9_;
input tin_pdata_1_1_;
input tin_pdata_4_4_;
input pclk;
input pirq_0_0_;
input tin_pdata_10_10_;
input tin_pdata_3_3_;
input tin_pdata_6_6_;
input tin_pdata_15_15_;
input tin_pdata_11_11_;
input tin_pdata_14_14_;
input tin_pdata_12_12_;
input tin_pdata_5_5_;
input preset;
input tin_pdata_13_13_;
output ppeakb_7_7_;
output ppeakp_12_12_;
output ppeakp_0_0_;
output ppeaka_7_7_;
output ppeaki_15_15_;
output ppeaki_11_11_;
output ppeaki_3_3_;
output paddress_3_3_;
output pdata_8_8_;
output pdata_0_0_;
output ppeakb_14_14_;
output ppeakb_10_10_;
output ppeakb_8_8_;
output ppeakp_1_1_;
output ppeaka_14_14_;
output ppeaka_10_10_;
output ppeaka_8_8_;
output ppeaki_4_4_;
output paddress_15_15_;
output paddress_11_11_;
output paddress_2_2_;
output ppeakb_9_9_;
output ppeakp_2_2_;
output ppeaka_9_9_;
output ppeaks_12_12_;
output ppeaks_0_0_;
output ppeaki_5_5_;
output paddress_5_5_;
output pdata_7_7_;
output ppeakb_15_15_;
output ppeakp_3_3_;
output pwr_0_0_;
output ppeaks_1_1_;
output ppeaki_6_6_;
output paddress_4_4_;
output piack_0_0_;
output ppeakp_13_13_;
output ppeakp_4_4_;
output ppeaka_15_15_;
output ppeaka_11_11_;
output ppeaks_2_2_;
output ppeaki_7_7_;
output paddress_10_10_;
output paddress_7_7_;
output pdata_2_2_;
output ppeakp_5_5_;
output ppeaks_13_13_;
output ppeaks_3_3_;
output ppeaki_14_14_;
output ppeaki_10_10_;
output ppeaki_8_8_;
output paddress_6_6_;
output ppeakp_6_6_;
output ppeaks_4_4_;
output ppeaki_9_9_;
output paddress_9_9_;
output pdata_9_9_;
output pdata_1_1_;
output ppeakb_11_11_;
output ppeakp_7_7_;
output ppeaks_5_5_;
output paddress_13_13_;
output paddress_8_8_;
output ppeakp_14_14_;
output ppeakp_10_10_;
output ppeakp_8_8_;
output ppeaks_6_6_;
output ppeaki_13_13_;
output pdata_4_4_;
output ppeakb_0_0_;
output ppeakp_9_9_;
output ppeaka_0_0_;
output ppeaks_7_7_;
output ppeakb_1_1_;
output ppeaka_1_1_;
output ppeaks_10_10_;
output ppeaks_8_8_;
output pdata_10_10_;
output pdata_3_3_;
output ppeakb_12_12_;
output ppeakb_2_2_;
output ppeaka_12_12_;
output ppeaka_2_2_;
output ppeaks_15_15_;
output ppeaks_9_9_;
output ppeakb_3_3_;
output ppeakp_15_15_;
output ppeakp_11_11_;
output ppeaka_13_13_;
output ppeaka_3_3_;
output paddress_14_14_;
output paddress_12_12_;
output pdata_6_6_;
output ppeakb_13_13_;
output ppeakb_4_4_;
output pdn;
output ppeaka_4_4_;
output ppeaki_0_0_;
output prd_0_0_;
output pdata_15_15_;
output pdata_11_11_;
output ppeakb_5_5_;
output ppeaka_5_5_;
output ppeaks_14_14_;
output ppeaki_1_1_;
output paddress_1_1_;
output pdata_14_14_;
output pdata_12_12_;
output pdata_5_5_;
output ppeakb_6_6_;
output ppeaka_6_6_;
output ppeaks_11_11_;
output ppeaki_12_12_;
output ppeaki_2_2_;
output paddress_0_0_;
output pdata_13_13_;
wire wire4244;
wire wire4259;
wire wire4274;
wire wire4289;
wire wire4304;
wire wire4319;
wire wire4334;
wire wire4349;
wire wire4364;
wire wire4379;
wire wire4394;
wire wire4409;
wire wire4424;
wire wire4439;
wire wire4454;
wire wire4469;
wire wire4484;
wire wire4499;
wire wire4514;
wire wire4529;
wire wire4544;
wire wire4559;
wire wire4574;
wire wire4589;
wire wire4604;
wire wire4619;
wire wire4634;
wire wire4649;
wire wire4664;
wire wire4679;
wire wire4709;
wire wire4724;
wire wire4739;
wire wire4754;
wire wire4769;
wire wire4784;
wire wire4799;
wire wire4814;
wire wire4829;
wire wire4844;
wire wire4859;
wire wire4874;
wire wire4889;
wire wire4904;
wire wire4919;
wire wire4934;
wire wire4949;
wire wire4964;
wire wire4979;
wire wire4994;
wire wire5009;
wire wire5024;
wire wire5039;
wire wire5054;
wire wire5069;
wire wire5084;
wire wire5099;
wire wire5114;
wire wire5129;
wire wire5144;
wire wire5159;
wire wire5174;
wire wire5189;
wire wire5204;
wire wire5219;
wire wire5234;
wire wire5249;
wire wire5264;
wire wire5279;
wire wire5294;
wire wire5309;
wire wire5324;
wire wire5339;
wire wire5354;
wire wire5369;
wire wire5384;
wire wire5399;
wire wire5414;
wire wire5429;
wire wire5444;
wire wire5459;
wire wire5474;
wire wire5489;
wire wire5504;
wire wire5519;
wire wire5534;
wire wire5549;
wire wire5564;
wire wire5579;
wire wire5609;
wire wire5624;
wire wire5639;
wire wire5654;
wire wire5669;
wire wire5684;
wire wire5699;
wire wire5714;
wire wire5729;
wire wire5744;
wire wire5759;
wire wire5774;
wire wire5789;
wire wire5804;
wire wire5819;
wire wire5834;
wire wire5849;
wire wire5864;
wire wire5879;
wire wire5894;
wire wire5909;
wire wire5924;
wire wire5939;
wire wire5954;
wire wire5969;
wire wire5984;
wire wire5999;
wire wire6014;
wire wire6029;
wire wire6044;
wire wire6059;
wire wire6074;
wire wire6089;
wire wire6104;
wire wire6119;
wire wire6134;
wire wire6149;
wire wire6164;
wire wire6179;
wire wire6194;
wire wire6209;
wire wire6224;
wire wire6239;
wire wire6254;
wire wire6269;
wire wire6284;
wire wire6299;
wire wire6314;
wire wire6329;
wire wire6344;
wire wire6359;
wire wire6374;
wire wire6389;
wire wire6404;
wire wire6419;
wire wire6434;
wire wire6449;
wire wire6464;
wire wire6479;
wire wire6494;
wire wire6509;
wire wire6524;
wire wire6539;
wire wire6554;
wire wire6569;
wire wire6584;
wire wire6599;
wire wire6614;
wire wire6629;
wire wire6644;
wire wire6659;
wire wire6674;
wire wire6689;
wire wire6704;
wire wire6719;
wire wire6734;
wire wire6749;
wire wire6764;
wire wire6779;
wire wire6794;
wire wire6824;
wire wire6839;
wire wire6854;
wire wire6869;
wire wire6884;
wire wire6899;
wire wire6914;
wire wire6929;
wire wire6944;
wire wire6959;
wire wire6974;
wire wire6989;
wire wire7004;
wire wire7019;
wire wire7034;
wire wire7064;
wire wire7079;
wire wire7094;
wire wire7109;
wire wire7124;
wire wire7139;
wire wire7154;
wire wire7169;
wire wire7184;
wire wire7199;
wire wire7214;
wire wire7229;
wire wire7244;
wire wire7259;
wire wire7274;
wire wire7289;
wire wire7304;
wire wire7319;
wire wire7334;
wire wire7349;
wire wire7364;
wire wire7379;
wire wire7394;
wire wire7409;
wire wire7424;
wire wire7439;
wire wire7454;
wire wire7469;
wire wire7484;
wire wire7499;
wire wire7514;
wire wire7529;
wire wire7544;
wire wire7559;
wire wire7574;
wire wire7589;
wire wire7604;
wire wire7634;
wire wire7649;
wire wire7664;
wire wire7679;
wire wire7694;
wire wire7709;
wire wire7724;
wire wire7739;
wire wire7754;
wire wire7769;
wire wire7784;
wire wire7799;
wire wire7814;
wire wire7829;
wire wire7844;
wire wire7859;
wire wire7874;
wire wire7889;
wire wire7904;
wire wire7919;
wire wire7934;
wire wire7949;
wire wire7964;
wire wire7979;
wire wire8009;
wire wire8024;
wire wire8039;
wire wire8054;
wire wire8069;
wire wire8084;
wire wire8099;
wire wire8114;
wire wire8129;
wire wire8144;
wire wire8159;
wire wire8174;
wire wire8189;
wire wire8204;
wire wire8219;
wire wire8234;
wire wire8249;
wire wire8264;
wire wire8294;
wire wire8309;
wire wire8324;
wire wire8339;
wire wire8354;
wire wire8369;
wire wire8384;
wire wire8399;
wire wire8414;
wire wire8429;
wire wire8444;
wire wire8459;
wire wire8474;
wire wire8489;
wire wire8504;
wire wire8519;
wire wire8534;
wire wire8549;
wire wire8564;
wire wire8579;
wire wire8594;
wire wire8609;
wire wire8624;
wire wire8639;
wire wire8654;
wire wire8669;
wire wire8684;
wire wire8699;
wire wire8714;
wire wire8729;
wire wire8744;
wire wire8759;
wire wire8774;
wire wire8789;
wire wire8819;
wire wire8834;
wire wire8849;
wire wire8864;
wire wire8879;
wire wire8894;
wire wire8909;
wire wire8924;
wire wire8939;
wire wire8954;
wire wire8969;
wire wire8984;
wire wire8999;
wire wire9014;
wire wire9029;
wire wire9044;
wire wire9059;
wire wire9074;
wire wire9089;
wire wire9104;
wire wire9119;
wire wire9134;
wire wire9149;
wire wire9164;
wire wire9179;
wire wire9194;
wire wire9209;
wire wire9224;
wire wire9239;
wire wire9254;
wire wire9269;
wire wire9284;
wire wire9299;
wire wire9314;
wire wire9329;
wire wire9344;
wire wire9359;
wire wire9374;
wire wire9389;
wire wire9404;
wire wire9419;
wire wire9449;
wire wire9464;
wire wire9479;
wire wire9494;
wire wire9509;
wire wire9524;
wire wire9539;
wire wire9554;
wire wire9569;
wire wire9584;
wire wire9599;
wire wire9614;
wire wire9629;
wire wire9644;
wire wire9659;
wire wire9674;
wire wire9689;
wire wire9704;
wire wire9719;
wire wire9734;
wire wire9749;
wire wire9779;
wire wire9794;
wire wire9809;
wire wire9824;
wire wire9839;
wire wire9854;
wire wire9869;
wire wire9884;
wire wire9899;
wire wire9914;
wire wire9929;
wire wire9944;
wire wire9959;
wire wire9989;
wire wire10004;
wire wire10019;
wire wire10034;
wire wire10049;
wire wire10064;
wire wire10079;
wire wire10094;
wire wire10109;
wire wire10124;
wire wire10139;
wire wire10154;
wire wire10184;
wire wire10199;
wire wire10214;
wire wire10229;
wire wire10244;
wire wire10259;
wire wire10274;
wire wire10289;
wire wire10319;
wire wire10334;
wire wire10349;
wire wire10364;
wire wire10379;
wire wire10409;
wire wire10424;
wire wire10439;
wire wire10454;
wire wire10469;
wire wire10484;
wire wire10499;
wire wire10514;
wire wire10529;
wire wire10544;
wire wire10559;
wire wire10574;
wire wire10589;
wire wire10604;
wire wire10619;
wire wire10634;
wire wire10664;
wire wire10679;
wire wire10694;
wire wire10709;
wire wire10724;
wire wire10739;
wire wire10754;
wire wire10769;
wire wire10784;
wire wire10799;
wire wire10814;
wire wire10829;
wire wire10859;
wire wire10874;
wire wire10889;
wire wire10904;
wire wire10934;
wire wire10949;
wire wire10964;
wire wire10979;
wire wire10994;
wire wire11024;
wire wire11039;
wire wire11054;
wire wire11069;
wire wire11084;
wire wire11099;
wire wire11129;
wire wire11144;
wire wire11159;
wire wire11174;
wire wire11189;
wire wire11204;
wire wire11219;
wire wire11234;
wire wire11249;
wire wire11264;
wire wire11279;
wire wire11294;
wire wire11309;
wire wire11324;
wire wire11339;
wire wire11354;
wire wire11384;
wire wire11399;
wire wire11414;
wire wire11429;
wire wire11444;
wire wire11459;
wire wire11474;
wire wire11489;
wire wire11504;
wire wire11519;
wire wire11534;
wire wire11549;
wire wire11564;
wire wire11579;
wire wire11594;
wire wire11609;
wire wire11624;
wire wire11639;
wire wire11654;
wire wire11669;
wire wire11684;
wire wire11699;
wire wire11714;
wire wire11729;
wire wire11744;
wire wire11759;
wire wire11774;
wire wire11789;
wire wire11804;
wire wire11819;
wire wire11864;
wire wire11879;
wire wire11894;
wire wire11909;
wire wire11924;
wire wire11939;
wire wire11984;
wire wire11999;
wire wire12014;
wire wire12029;
wire wire12044;
wire wire12059;
wire wire12074;
wire wire12089;
wire wire12119;
wire wire12134;
wire wire12149;
wire wire12164;
wire wire12179;
wire wire12194;
wire wire12209;
wire wire12239;
wire wire12254;
wire wire12269;
wire wire12284;
wire wire12314;
wire wire12329;
wire wire12344;
wire wire12359;
wire wire12374;
wire wire12389;
wire wire12404;
wire wire12419;
wire wire12434;
wire wire12449;
wire wire12464;
wire wire12479;
wire wire12494;
wire wire12524;
wire wire12539;
wire wire12554;
wire wire12569;
wire wire12584;
wire wire12599;
wire wire12614;
wire wire12629;
wire wire12644;
wire wire12659;
wire wire12674;
wire wire12689;
wire wire12704;
wire wire12749;
wire wire12764;
wire wire12779;
wire wire12809;
wire wire12824;
wire wire12839;
wire wire12854;
wire wire12869;
wire wire12884;
wire wire12899;
wire wire12914;
wire wire12929;
wire wire12944;
wire wire12989;
wire wire13004;
wire wire13019;
wire wire13034;
wire wire13049;
wire wire13064;
wire wire13079;
wire wire13094;
wire wire13109;
wire wire13124;
wire wire13139;
wire wire13169;
wire wire13184;
wire wire13199;
wire wire13214;
wire wire13229;
wire wire13244;
wire wire13259;
wire wire13274;
wire wire13289;
wire wire13304;
wire wire13319;
wire wire13334;
wire wire13349;
wire wire13364;
wire wire13379;
wire wire13394;
wire wire13409;
wire wire13424;
wire wire13439;
wire wire13454;
wire wire13469;
wire wire13484;
wire wire13499;
wire wire13514;
wire wire13544;
wire wire13559;
wire wire13574;
wire wire13589;
wire wire13604;
wire wire13619;
wire wire13634;
wire wire13649;
wire wire13664;
wire wire13679;
wire wire13694;
wire wire13709;
wire wire13724;
wire wire13739;
wire wire13754;
wire wire13784;
wire wire13799;
wire wire13814;
wire wire13829;
wire wire13844;
wire wire13859;
wire wire13874;
wire wire13889;
wire wire13904;
wire wire13919;
wire wire13934;
wire wire13949;
wire wire13964;
wire wire13979;
wire wire13994;
wire wire14009;
wire wire14024;
wire wire14039;
wire wire14054;
wire wire14069;
wire wire14084;
wire wire14099;
wire wire14114;
wire wire14129;
wire wire14144;
wire wire14159;
wire wire14174;
wire wire14189;
wire wire14219;
wire wire14234;
wire wire14249;
wire wire14264;
wire wire14279;
wire wire14294;
wire wire14309;
wire wire14324;
wire wire14339;
wire wire14354;
wire wire14369;
wire wire14384;
wire wire14399;
wire wire14414;
wire wire14429;
wire wire14444;
wire wire14459;
wire wire14474;
wire wire14489;
wire wire14504;
wire wire14519;
wire wire14534;
wire wire14549;
wire wire14564;
wire wire14579;
wire wire14594;
wire wire14609;
wire wire14624;
wire wire14639;
wire wire14669;
wire wire14684;
wire wire14699;
wire wire14714;
wire wire14729;
wire wire14744;
wire wire14759;
wire wire14774;
wire wire14789;
wire wire14804;
wire wire14819;
wire wire14834;
wire wire14849;
wire wire14864;
wire wire14879;
wire wire14894;
wire wire14909;
wire wire14924;
wire wire14939;
wire wire14969;
wire wire14984;
wire wire14999;
wire wire15014;
wire wire15029;
wire wire15044;
wire wire15059;
wire wire15074;
wire wire15089;
wire wire15104;
wire wire15119;
wire wire15134;
wire wire15149;
wire wire15164;
wire wire15179;
wire wire15194;
wire wire15209;
wire wire15224;
wire wire15239;
wire wire15254;
wire wire15269;
wire wire15284;
wire wire15299;
wire wire15314;
wire wire15329;
wire wire15344;
wire wire15359;
wire wire15374;
wire wire15389;
wire wire15404;
wire wire15419;
wire wire15434;
wire wire15449;
wire wire15464;
wire wire15479;
wire wire15494;
wire wire15509;
wire wire15524;
wire wire15539;
wire wire15554;
wire wire15569;
wire wire15584;
wire wire15599;
wire wire15614;
wire wire15629;
wire wire15644;
wire wire15659;
wire wire15674;
wire wire15689;
wire wire15704;
wire wire15719;
wire wire15734;
wire wire15764;
wire wire15779;
wire wire15794;
wire wire15809;
wire wire15824;
wire wire15839;
wire wire15854;
wire wire15869;
wire wire15884;
wire wire15899;
wire wire15914;
wire wire15929;
wire wire15944;
wire wire15959;
wire wire15974;
wire wire15989;
wire wire16004;
wire wire16019;
wire wire16034;
wire wire16049;
wire wire16064;
wire wire16079;
wire wire16094;
wire wire16109;
wire wire16904;
wire wire16917;
wire wire16928;
wire wire16941;
wire wire16956;
wire wire16969;
wire wire16980;
wire wire16993;
wire wire17008;
wire wire17021;
wire wire17032;
wire wire17045;
wire wire17058;
wire wire17073;
wire wire17086;
wire wire17097;
wire wire17110;
wire wire17123;
wire wire17138;
wire wire17151;
wire wire17162;
wire wire17175;
wire wire17188;
wire wire17203;
wire wire17214;
wire wire17227;
wire wire17240;
wire wire17253;
wire wire17268;
wire wire17279;
wire wire17292;
wire wire17305;
wire wire17318;
wire wire17333;
wire wire17346;
wire wire17357;
wire wire17370;
wire wire17383;
wire wire17396;
wire wire17411;
wire wire17422;
wire wire17435;
wire wire17461;
wire wire17476;
wire wire17489;
wire wire17502;
wire wire17513;
wire wire17526;
wire wire17539;
wire wire17554;
wire wire17567;
wire wire17578;
wire wire17591;
wire wire17604;
wire wire17619;
wire wire17632;
wire wire17643;
wire wire17656;
wire wire17669;
wire wire17684;
wire wire17697;
wire wire17708;
wire wire17723;
wire wire17736;
wire wire17747;
wire wire17760;
wire wire17775;
wire wire17788;
wire wire17799;
wire wire17812;
wire wire17825;
wire wire17840;
wire wire17851;
wire wire17866;
wire wire17879;
wire wire17892;
wire wire17905;
wire wire17918;
wire wire17931;
wire wire17944;
wire wire17957;
wire wire17970;
wire wire17983;
wire wire17994;
wire wire18007;
wire wire18022;
wire wire18033;
wire wire18048;
wire wire18059;
wire wire18072;
wire wire18085;
wire wire18100;
wire wire18111;
wire wire18126;
wire wire18139;
wire wire18150;
wire wire18165;
wire wire18176;
wire wire18191;
wire wire18204;
wire wire18215;
wire wire18228;
wire wire18243;
wire wire18254;
wire wire18269;
wire wire18282;
wire wire18293;
wire wire18306;
wire wire18319;
wire wire18334;
wire wire18347;
wire wire18360;
wire wire18371;
wire wire18384;
wire wire18397;
wire wire18412;
wire wire18423;
wire wire18436;
wire wire18449;
wire wire18464;
wire wire18475;
wire wire18488;
wire wire18501;
wire wire18514;
wire wire18529;
wire wire18542;
wire wire18555;
wire wire18568;
wire wire18581;
wire wire18594;
wire wire18605;
wire wire18618;
wire wire18633;
wire wire18644;
wire wire4305;
wire wire4260;
wire wire4269;
wire wire4298;
wire wire4392;
wire wire4397;
wire wire4226;
wire wire4352;
wire wire4280;
wire wire4353;
wire wire4243;
wire wire4253;
wire wire4354;
wire wire4245;
wire wire4252;
wire wire4375;
wire wire19360;
wire wire4340;
wire wire19390;
wire wire4308;
wire wire4306;
wire wire4317;
wire wire4381;
wire wire19368;
wire wire19359;
wire wire4377;
wire wire4277;
wire wire4278;
wire wire19088;
wire wire4350;
wire wire19092;
wire wire4345;
wire wire19103;
wire wire4330;
wire wire4374;
wire wire19060;
wire wire4360;
wire wire19097;
wire wire4331;
wire wire4332;
wire wire19061;
wire wire19091;
wire wire4336;
wire wire4365;
wire wire19367;
wire wire19387;
wire wire19070;
wire wire19096;
wire wire19072;
wire wire19087;
wire wire19082;
wire wire19396;
wire wire4383;
wire wire19073;
wire wire4307;
wire wire4325;
wire wire19068;
wire wire19065;
wire wire4357;
wire wire1427;
wire wire4199;
wire wire4358;
wire wire1342;
wire wire1353;
wire wire4359;
wire wire1412;
wire wire1397;
wire wire4316;
wire wire4327;
wire wire1439;
wire wire1368;
wire wire4368;
wire wire1386;
wire wire1411;
wire wire1398;
wire wire1434;
wire wire1413;
wire wire4341;
wire wire4351;
wire wire4369;
wire wire4378;
wire wire4382;
wire wire4467;
wire wire4458;
wire nrq21_7;
wire nrq13_4;
wire wire4300;
wire ndn7_2;
wire wire4466;
wire nen3_5;
wire nrq3_11;
wire nrq8_2;
wire nen2_3;
wire wire4235;
wire wire4513;
wire wire4241;
wire nrq10_4;
wire nrq4_14;
wire nrq14_8;
wire nen3_2;
wire n_n2344;
wire nsl8_2;
wire nrq7_2;
wire nrq1_4;
wire wire3723;
wire wire3744;
wire wire3738;
wire wire3718;
wire n_n3925;
wire ndn_latch3_9;
wire wire3740;
wire ndn_latch12_11;
wire wire3715;
wire ndn_latch13_2;
wire ndn_latch24_2;
wire wire3746;
wire wire3747;
wire nrq23_3;
wire wire3770;
wire wire3775;
wire nrq3_5;
wire nrq14_3;
wire nrq4_9;
wire wire3727;
wire nrq17_3;
wire wire3711;
wire nrq15_5;
wire nrq21_5;
wire nrq4_5;
wire nrq4_2;
wire wire3750;
wire wire3754;
wire n_n2333;
wire n_n3712;
wire n_n2326;
wire n_n2314;
wire n_n2325;
wire n_n2316;
wire n_n2318;
wire n_n2323;
wire n_n2317;
wire n_n2315;
wire n_n2321;
wire n_n2324;
wire n_n2320;
wire n_n2322;
wire n_n2319;
wire wire3784;
wire wire4468;
wire wire4470;
wire wire4391;
wire wire4483;
wire wire4273;
wire n_n2453;
wire n_n2452;
wire wire4465;
wire wire4471;
wire wire4459;
wire wire4480;
wire wire4472;
wire wire4205;
wire n_n2772;
wire wire4234;
wire wire4242;
wire n_n2443;
wire n_n2449;
wire n_n3711;
wire n_n2442;
wire n_n2446;
wire n_n2447;
wire n_n2445;
wire n_n2441;
wire n_n2440;
wire n_n2444;
wire n_n2454;
wire n_n2450;
wire n_n2451;
wire n_n2448;
wire n_n3081;
wire n_n3714;
wire wire3720;
wire nlbr8_2_e;
wire wire4265;
wire wire4488;
wire n_n2475;
wire n_n3713;
wire n_n2472;
wire wire4292;
wire n_n2484;
wire n_n2474;
wire n_n2479;
wire n_n2483;
wire n_n2485;
wire n_n2482;
wire n_n2480;
wire n_n2486;
wire n_n2473;
wire n_n2471;
wire n_n2487;
wire n_n2476;
wire n_n2478;
wire n_n2477;
wire n_n2481;
wire wire4024;
wire wire19749;
wire wire19466;
wire wire19739;
wire wire19514;
wire wire19741;
wire wire19531;
wire wire4438;
wire wire19727;
wire wire19456;
wire wire4440;
wire wire19735;
wire wire19504;
wire wire19725;
wire wire19479;
wire wire19731;
wire wire19474;
wire wire4301;
wire wire19747;
wire wire19721;
wire wire19452;
wire wire19733;
wire wire19737;
wire wire19520;
wire wire19495;
wire wire19171;
wire wire19221;
wire wire19205;
wire wire19232;
wire wire19157;
wire wire19180;
wire wire4388;
wire wire4511;
wire wire19227;
wire wire19153;
wire wire4496;
wire wire19191;
wire wire19215;
wire wire4410;
wire wire19729;
wire wire19196;
wire wire19175;
wire wire19743;
wire wire4450;
wire wire19167;
wire wire4451;
wire wire4457;
wire wire4507;
wire wire4452;
wire wire4508;
wire wire19989;
wire wire4453;
wire wire18861;
wire wire4455;
wire wire4456;
wire wire4509;
wire wire4202;
wire wire4204;
wire wire4207;
wire wire4208;
wire wire4209;
wire wire4211;
wire wire4212;
wire wire4215;
wire wire4266;
wire wire4219;
wire wire4303;
wire wire4224;
wire wire4225;
wire wire4515;
wire wire1914;
wire wire1915;
wire wire1918;
wire wire1920;
wire wire1921;
wire wire1922;
wire wire1923;
wire wire1926;
wire wire1927;
wire wire1928;
wire wire1929;
wire wire1930;
wire wire1935;
wire wire1936;
wire wire1944;
wire wire1946;
wire wire1947;
wire wire1948;
wire wire1949;
wire wire1952;
wire wire1953;
wire wire1954;
wire wire1955;
wire wire1956;
wire wire1961;
wire wire1963;
wire wire1964;
wire wire1965;
wire wire1966;
wire wire1969;
wire wire1970;
wire wire1971;
wire wire1972;
wire wire1973;
wire wire1976;
wire wire1978;
wire wire1979;
wire wire1980;
wire wire1981;
wire wire1984;
wire wire1985;
wire wire1986;
wire wire1987;
wire wire1988;
wire wire1991;
wire wire1992;
wire wire1995;
wire wire1997;
wire wire1998;
wire wire1999;
wire wire2000;
wire wire2003;
wire wire2004;
wire wire2005;
wire wire2006;
wire wire2007;
wire wire2010;
wire wire2012;
wire wire2013;
wire wire2014;
wire wire2015;
wire wire2018;
wire wire2019;
wire wire2020;
wire wire2021;
wire wire2022;
wire wire2028;
wire wire2029;
wire wire2032;
wire wire2034;
wire wire2035;
wire wire2036;
wire wire2037;
wire wire2040;
wire wire2041;
wire wire2042;
wire wire2043;
wire wire2044;
wire wire2045;
wire wire2049;
wire wire2050;
wire wire2051;
wire wire2055;
wire wire2057;
wire wire2058;
wire wire2059;
wire wire2060;
wire wire2063;
wire wire2064;
wire wire2065;
wire wire2066;
wire wire2067;
wire wire2068;
wire wire2069;
wire wire2070;
wire wire2076;
wire wire2077;
wire wire2080;
wire wire2081;
wire wire2084;
wire wire2085;
wire wire2088;
wire wire2089;
wire wire2092;
wire wire2100;
wire wire2101;
wire wire2107;
wire wire2108;
wire wire2116;
wire wire2117;
wire wire2179;
wire wire2184;
wire wire2185;
wire wire2187;
wire wire2188;
wire wire2193;
wire wire2195;
wire wire2196;
wire wire2197;
wire wire2198;
wire wire2201;
wire wire2202;
wire wire2203;
wire wire2204;
wire wire2205;
wire wire2210;
wire wire2212;
wire wire2213;
wire wire2214;
wire wire2215;
wire wire2218;
wire wire2219;
wire wire2220;
wire wire2221;
wire wire2222;
wire wire2231;
wire wire2233;
wire wire2234;
wire wire2235;
wire wire2236;
wire wire2239;
wire wire2240;
wire wire2241;
wire wire2242;
wire wire2243;
wire wire2246;
wire wire2255;
wire wire2260;
wire wire2262;
wire wire2263;
wire wire2264;
wire wire2265;
wire wire2268;
wire wire2269;
wire wire2270;
wire wire2271;
wire wire2272;
wire wire2276;
wire wire2280;
wire wire2281;
wire wire2286;
wire wire2288;
wire wire2289;
wire wire2290;
wire wire2291;
wire wire2294;
wire wire2295;
wire wire2296;
wire wire2297;
wire wire2298;
wire wire2303;
wire wire2305;
wire wire2306;
wire wire2307;
wire wire2308;
wire wire2311;
wire wire2312;
wire wire2313;
wire wire2314;
wire wire2315;
wire wire2319;
wire wire2320;
wire wire2324;
wire wire2325;
wire wire2329;
wire wire2330;
wire wire2336;
wire wire2337;
wire wire2341;
wire wire2342;
wire wire2344;
wire wire2345;
wire wire2351;
wire wire2352;
wire wire2354;
wire wire2355;
wire wire2358;
wire wire2360;
wire wire2361;
wire wire2362;
wire wire2363;
wire wire2366;
wire wire2367;
wire wire2368;
wire wire2369;
wire wire2370;
wire wire2374;
wire wire2375;
wire wire2378;
wire wire2380;
wire wire2381;
wire wire2382;
wire wire2383;
wire wire2386;
wire wire2387;
wire wire2388;
wire wire2389;
wire wire2390;
wire wire2391;
wire wire2392;
wire wire2394;
wire wire2400;
wire wire2402;
wire wire2404;
wire wire2408;
wire wire2410;
wire wire2411;
wire wire2412;
wire wire2413;
wire wire2414;
wire wire2415;
wire wire2416;
wire wire2417;
wire wire2423;
wire wire2425;
wire wire2428;
wire wire2429;
wire wire2430;
wire wire2431;
wire wire2432;
wire wire2433;
wire wire2434;
wire wire2435;
wire wire2436;
wire wire2437;
wire wire2438;
wire wire2440;
wire wire2441;
wire wire2443;
wire wire2445;
wire wire2446;
wire wire2447;
wire wire2449;
wire wire2450;
wire wire2451;
wire wire2452;
wire wire2453;
wire wire2454;
wire wire2455;
wire wire2456;
wire wire2457;
wire wire2458;
wire wire2459;
wire wire2460;
wire wire2461;
wire wire2462;
wire wire2463;
wire wire2464;
wire wire2465;
wire wire2466;
wire wire2468;
wire wire2469;
wire wire2472;
wire wire2473;
wire wire2474;
wire wire2476;
wire wire2479;
wire wire2480;
wire wire2481;
wire wire2482;
wire wire2483;
wire wire2484;
wire wire2485;
wire wire2486;
wire wire2488;
wire wire2489;
wire wire2491;
wire wire2492;
wire wire2498;
wire wire2500;
wire wire2501;
wire wire2503;
wire wire2508;
wire wire2509;
wire wire2510;
wire wire2511;
wire wire2512;
wire wire2513;
wire wire2519;
wire wire2521;
wire wire2524;
wire wire2525;
wire wire2526;
wire wire2527;
wire wire2528;
wire wire2529;
wire wire2530;
wire wire2531;
wire wire2532;
wire wire2533;
wire wire2534;
wire wire2536;
wire wire2537;
wire wire2539;
wire wire2541;
wire wire2542;
wire wire2543;
wire wire2545;
wire wire2546;
wire wire2547;
wire wire2548;
wire wire2549;
wire wire2550;
wire wire2551;
wire wire2552;
wire wire2553;
wire wire2554;
wire wire2555;
wire wire2556;
wire wire2557;
wire wire2558;
wire wire2559;
wire wire2560;
wire wire2561;
wire wire2562;
wire wire2563;
wire wire2564;
wire wire2565;
wire wire2566;
wire wire2567;
wire wire2568;
wire wire2569;
wire wire2570;
wire wire2571;
wire wire2572;
wire wire2573;
wire wire2574;
wire wire2576;
wire wire2577;
wire wire2578;
wire wire2579;
wire wire2580;
wire wire2581;
wire wire2582;
wire wire2583;
wire wire2584;
wire wire2585;
wire wire2586;
wire wire2587;
wire wire2592;
wire wire2594;
wire wire2595;
wire wire2597;
wire wire2598;
wire wire2599;
wire wire2602;
wire wire2607;
wire wire2608;
wire wire2609;
wire wire2610;
wire wire2611;
wire wire2612;
wire wire2614;
wire wire2618;
wire wire2620;
wire wire2623;
wire wire2625;
wire wire2626;
wire wire2627;
wire wire2629;
wire wire2630;
wire wire2631;
wire wire2632;
wire wire2633;
wire wire2634;
wire wire2635;
wire wire2636;
wire wire2637;
wire wire2638;
wire wire2639;
wire wire2641;
wire wire2642;
wire wire2644;
wire wire2646;
wire wire2647;
wire wire2648;
wire wire2649;
wire wire2650;
wire wire2651;
wire wire2652;
wire wire2653;
wire wire2654;
wire wire2655;
wire wire2656;
wire wire2657;
wire wire2658;
wire wire2659;
wire wire2660;
wire wire2661;
wire wire2662;
wire wire2663;
wire wire2665;
wire wire2666;
wire wire2669;
wire wire2670;
wire wire2671;
wire wire2673;
wire wire2676;
wire wire2678;
wire wire2679;
wire wire2680;
wire wire2681;
wire wire2682;
wire wire2683;
wire wire2684;
wire wire2685;
wire wire2686;
wire wire2687;
wire wire2688;
wire wire2689;
wire wire2694;
wire wire2696;
wire wire2697;
wire wire2699;
wire wire2700;
wire wire2701;
wire wire2702;
wire wire2703;
wire wire2704;
wire wire2706;
wire wire2709;
wire wire2710;
wire wire2711;
wire wire2712;
wire wire2713;
wire wire2714;
wire wire2716;
wire wire2722;
wire wire2725;
wire wire2727;
wire wire2728;
wire wire2729;
wire wire2731;
wire wire2732;
wire wire2733;
wire wire2734;
wire wire2735;
wire wire2736;
wire wire2737;
wire wire2738;
wire wire2739;
wire wire2740;
wire wire2741;
wire wire2743;
wire wire2744;
wire wire2746;
wire wire2748;
wire wire2749;
wire wire2750;
wire wire2751;
wire wire2752;
wire wire2753;
wire wire2754;
wire wire2755;
wire wire2756;
wire wire2757;
wire wire2758;
wire wire2759;
wire wire2760;
wire wire2761;
wire wire2762;
wire wire2763;
wire wire2764;
wire wire2765;
wire wire2766;
wire wire2767;
wire wire2768;
wire wire2771;
wire wire2772;
wire wire2773;
wire wire2775;
wire wire2778;
wire wire2780;
wire wire2781;
wire wire2782;
wire wire2783;
wire wire2784;
wire wire2785;
wire wire2786;
wire wire2787;
wire wire2788;
wire wire2789;
wire wire2790;
wire wire2791;
wire wire2800;
wire wire2802;
wire wire2803;
wire wire2804;
wire wire2805;
wire wire2806;
wire wire2807;
wire wire2809;
wire wire2810;
wire wire2812;
wire wire2814;
wire wire2816;
wire wire2817;
wire wire2818;
wire wire2819;
wire wire2820;
wire wire2821;
wire wire2822;
wire wire2823;
wire wire2826;
wire wire2830;
wire wire2834;
wire wire2836;
wire wire2837;
wire wire2839;
wire wire2840;
wire wire2841;
wire wire2843;
wire wire2844;
wire wire2845;
wire wire2846;
wire wire2847;
wire wire2848;
wire wire2849;
wire wire2850;
wire wire2851;
wire wire2852;
wire wire2853;
wire wire2854;
wire wire2855;
wire wire2856;
wire wire2857;
wire wire2858;
wire wire2859;
wire wire2860;
wire wire2861;
wire wire2862;
wire wire2863;
wire wire2864;
wire wire2865;
wire wire2866;
wire wire2867;
wire wire2868;
wire wire2869;
wire wire2870;
wire wire2872;
wire wire2873;
wire wire2874;
wire wire2875;
wire wire2876;
wire wire2877;
wire wire2878;
wire wire2879;
wire wire2880;
wire wire2881;
wire wire2882;
wire wire2883;
wire wire2892;
wire wire2894;
wire wire2895;
wire wire2897;
wire wire2899;
wire wire2900;
wire wire2901;
wire wire2906;
wire wire2908;
wire wire2909;
wire wire2910;
wire wire2911;
wire wire2912;
wire wire2913;
wire wire2914;
wire wire2915;
wire wire2918;
wire wire2922;
wire wire2924;
wire wire2926;
wire wire2927;
wire wire2929;
wire wire2930;
wire wire2931;
wire wire2933;
wire wire2934;
wire wire2935;
wire wire2936;
wire wire2937;
wire wire2938;
wire wire2939;
wire wire2940;
wire wire2941;
wire wire2942;
wire wire2943;
wire wire2944;
wire wire2945;
wire wire2946;
wire wire2949;
wire wire2950;
wire wire2951;
wire wire2952;
wire wire2955;
wire wire2956;
wire wire2957;
wire wire2959;
wire wire2962;
wire wire2963;
wire wire2966;
wire wire2972;
wire wire2974;
wire wire2977;
wire wire2978;
wire wire2979;
wire wire2981;
wire wire2982;
wire wire2986;
wire wire2988;
wire wire2989;
wire wire2990;
wire wire2991;
wire wire2992;
wire wire2993;
wire wire2994;
wire wire2995;
wire wire2996;
wire wire3000;
wire wire3004;
wire wire3005;
wire wire3007;
wire wire3008;
wire wire3009;
wire wire3012;
wire wire3013;
wire wire3014;
wire wire3015;
wire wire3016;
wire wire3017;
wire wire3018;
wire wire3019;
wire wire3020;
wire wire3021;
wire wire3023;
wire wire3024;
wire wire3026;
wire wire3032;
wire wire3034;
wire wire3037;
wire wire3038;
wire wire3039;
wire wire3040;
wire wire3041;
wire wire3043;
wire wire3044;
wire wire3049;
wire wire3050;
wire wire3051;
wire wire3052;
wire wire3053;
wire wire3054;
wire wire3055;
wire wire3056;
wire wire3060;
wire wire3064;
wire wire3066;
wire wire3067;
wire wire3069;
wire wire3070;
wire wire3073;
wire wire3074;
wire wire3075;
wire wire3077;
wire wire3080;
wire wire3081;
wire wire3082;
wire wire3083;
wire wire3084;
wire wire3085;
wire wire3086;
wire wire3087;
wire wire3089;
wire wire3090;
wire wire3092;
wire wire3098;
wire wire3100;
wire wire3102;
wire wire3103;
wire wire3105;
wire wire3107;
wire wire3108;
wire wire3109;
wire wire3111;
wire wire3113;
wire wire3114;
wire wire3115;
wire wire3116;
wire wire3120;
wire wire3121;
wire wire3124;
wire wire3132;
wire wire3134;
wire wire3136;
wire wire3137;
wire wire3138;
wire wire3139;
wire wire3140;
wire wire3141;
wire wire3142;
wire wire3143;
wire wire3144;
wire wire3145;
wire wire3146;
wire wire3150;
wire wire3151;
wire wire3154;
wire wire3162;
wire wire3164;
wire wire3166;
wire wire3167;
wire wire3168;
wire wire3169;
wire wire3173;
wire wire3174;
wire wire3175;
wire wire3176;
wire wire3180;
wire wire3183;
wire wire3185;
wire wire3191;
wire wire3193;
wire wire3195;
wire wire3197;
wire wire3198;
wire wire3200;
wire wire3201;
wire wire3203;
wire wire3204;
wire wire3205;
wire wire3209;
wire wire3212;
wire wire3214;
wire wire3218;
wire wire3219;
wire wire3220;
wire wire3221;
wire wire3222;
wire wire3223;
wire wire3224;
wire wire3225;
wire wire3226;
wire wire3227;
wire wire3228;
wire wire3230;
wire wire3232;
wire wire3234;
wire wire3236;
wire wire3237;
wire wire3241;
wire wire3242;
wire wire3247;
wire wire3249;
wire wire3251;
wire wire3253;
wire wire3254;
wire wire3259;
wire wire3260;
wire wire3261;
wire wire3262;
wire wire3263;
wire wire3264;
wire wire3265;
wire wire3266;
wire wire3267;
wire wire3268;
wire wire3269;
wire wire3270;
wire wire3271;
wire wire3274;
wire wire3276;
wire wire3278;
wire wire3280;
wire wire3281;
wire wire3282;
wire wire3283;
wire wire3284;
wire wire3285;
wire wire3286;
wire wire3287;
wire wire3289;
wire wire3290;
wire wire3292;
wire wire3293;
wire wire3294;
wire wire3297;
wire wire3299;
wire wire3301;
wire wire3303;
wire wire3304;
wire wire3315;
wire wire3317;
wire wire3322;
wire wire3325;
wire wire3327;
wire wire3329;
wire wire3331;
wire wire3333;
wire wire3334;
wire wire3345;
wire wire3347;
wire wire3350;
wire wire3352;
wire wire3353;
wire wire3357;
wire wire3359;
wire wire3361;
wire wire3363;
wire wire3364;
wire wire3370;
wire wire3375;
wire wire3377;
wire wire3382;
wire wire3387;
wire wire3389;
wire wire3391;
wire wire3393;
wire wire3395;
wire wire3396;
wire wire3405;
wire wire3407;
wire wire3410;
wire wire3412;
wire wire3413;
wire wire3414;
wire wire3417;
wire wire3419;
wire wire3421;
wire wire3423;
wire wire3425;
wire wire3426;
wire wire3430;
wire wire3432;
wire wire3441;
wire wire3443;
wire wire3445;
wire wire3447;
wire wire3448;
wire wire3450;
wire wire3453;
wire wire3454;
wire wire3455;
wire wire3459;
wire wire3462;
wire wire3464;
wire wire3466;
wire wire3469;
wire wire3471;
wire wire3478;
wire wire3480;
wire wire3481;
wire wire3482;
wire wire3483;
wire wire3484;
wire wire3487;
wire wire3488;
wire wire3491;
wire wire3492;
wire wire3496;
wire wire3499;
wire wire3501;
wire wire3506;
wire wire3515;
wire wire3517;
wire wire3519;
wire wire3522;
wire wire3531;
wire wire3533;
wire wire3538;
wire wire3540;
wire wire3549;
wire wire3551;
wire wire3552;
wire wire3553;
wire wire3555;
wire wire3557;
wire wire3559;
wire wire3562;
wire wire3563;
wire wire3568;
wire wire3570;
wire wire3575;
wire wire3577;
wire wire3582;
wire wire3588;
wire wire3590;
wire wire3592;
wire wire3598;
wire wire3599;
wire wire3600;
wire wire3602;
wire wire3603;
wire wire3605;
wire wire3606;
wire wire3611;
wire wire3612;
wire wire3613;
wire wire3614;
wire wire3616;
wire wire3620;
wire wire3622;
wire wire3624;
wire wire3633;
wire wire3634;
wire wire3635;
wire wire3637;
wire wire3640;
wire wire3642;
wire wire3650;
wire wire3651;
wire wire3653;
wire wire3654;
wire wire3655;
wire wire3657;
wire wire3659;
wire wire3660;
wire wire3661;
wire wire3663;
wire wire3664;
wire wire3665;
wire wire3666;
wire wire3667;
wire wire3668;
wire wire3669;
wire wire3670;
wire wire3671;
wire wire3672;
wire wire3673;
wire wire3675;
wire wire3676;
wire wire3678;
wire wire3679;
wire wire3680;
wire wire3681;
wire wire3682;
wire wire3683;
wire wire3684;
wire wire3685;
wire wire3686;
wire wire3687;
wire wire3688;
wire wire3689;
wire wire3691;
wire wire3692;
wire wire3694;
wire wire3699;
wire wire3701;
wire wire3706;
wire wire3713;
wire wire3716;
wire wire3719;
wire wire3721;
wire wire3725;
wire wire3730;
wire wire3731;
wire wire3733;
wire wire3735;
wire wire3737;
wire wire3741;
wire wire3743;
wire wire3749;
wire wire3751;
wire wire3757;
wire wire3759;
wire wire3768;
wire wire3769;
wire wire3771;
wire wire3773;
wire wire3777;
wire wire3788;
wire wire3789;
wire wire3791;
wire wire3792;
wire wire3793;
wire wire3795;
wire wire3797;
wire wire3798;
wire wire3799;
wire wire3801;
wire wire3802;
wire wire3803;
wire wire3804;
wire wire3805;
wire wire3806;
wire wire3807;
wire wire3808;
wire wire3809;
wire wire3810;
wire wire3811;
wire wire3813;
wire wire3814;
wire wire3816;
wire wire3818;
wire wire3819;
wire wire3820;
wire wire3825;
wire wire3834;
wire wire3836;
wire wire3838;
wire wire3842;
wire wire3843;
wire wire3844;
wire wire3846;
wire wire3848;
wire wire3849;
wire wire3850;
wire wire3851;
wire wire3853;
wire wire3857;
wire wire3858;
wire wire3859;
wire wire3860;
wire wire3862;
wire wire3866;
wire wire3868;
wire wire3875;
wire wire3876;
wire wire3877;
wire wire3878;
wire wire3879;
wire wire3881;
wire wire3884;
wire wire3886;
wire wire3894;
wire wire3895;
wire wire3897;
wire wire3898;
wire wire3899;
wire wire3901;
wire wire3903;
wire wire3904;
wire wire3905;
wire wire3907;
wire wire3908;
wire wire3909;
wire wire3910;
wire wire3911;
wire wire3912;
wire wire3913;
wire wire3914;
wire wire3915;
wire wire3916;
wire wire3917;
wire wire3919;
wire wire3920;
wire wire3922;
wire wire3924;
wire wire3925;
wire wire3926;
wire wire3929;
wire wire3931;
wire wire3938;
wire wire3940;
wire wire3942;
wire wire3945;
wire wire3947;
wire wire3948;
wire wire3950;
wire wire3953;
wire wire3955;
wire wire3956;
wire wire3957;
wire wire3960;
wire wire3961;
wire wire3963;
wire wire3967;
wire wire3970;
wire wire3972;
wire wire3974;
wire wire3981;
wire wire3982;
wire wire3983;
wire wire3984;
wire wire3985;
wire wire3988;
wire wire3990;
wire wire3992;
wire wire4000;
wire wire4001;
wire wire4003;
wire wire4004;
wire wire4005;
wire wire4007;
wire wire4008;
wire wire4009;
wire wire4010;
wire wire4011;
wire wire4012;
wire wire4013;
wire wire4014;
wire wire4015;
wire wire4016;
wire wire4017;
wire wire4019;
wire wire4020;
wire wire4022;
wire wire4023;
wire wire4025;
wire wire4026;
wire wire4027;
wire wire4028;
wire wire4029;
wire wire4030;
wire wire4031;
wire wire4032;
wire wire4033;
wire wire4034;
wire wire4036;
wire wire4037;
wire wire4039;
wire wire4041;
wire wire4042;
wire wire4043;
wire wire4047;
wire wire4056;
wire wire4058;
wire wire4060;
wire wire4062;
wire wire4065;
wire wire4067;
wire wire4073;
wire wire4074;
wire wire4075;
wire wire4076;
wire wire4077;
wire wire4079;
wire wire4080;
wire wire4085;
wire wire4088;
wire wire4090;
wire wire4092;
wire wire4099;
wire wire4100;
wire wire4101;
wire wire4102;
wire wire4103;
wire wire4105;
wire wire4108;
wire wire4120;
wire wire4121;
wire wire4123;
wire wire4124;
wire wire4125;
wire wire4127;
wire wire4128;
wire wire4129;
wire wire4130;
wire wire4131;
wire wire4132;
wire wire4133;
wire wire4134;
wire wire4135;
wire wire4136;
wire wire4137;
wire wire4139;
wire wire4140;
wire wire4142;
wire wire4143;
wire wire4144;
wire wire4145;
wire wire4146;
wire wire4147;
wire wire4148;
wire wire4149;
wire wire4150;
wire wire4151;
wire wire4152;
wire wire4153;
wire wire4155;
wire wire4156;
wire wire4158;
wire wire4160;
wire wire4161;
wire wire4162;
wire wire4163;
wire wire4164;
wire wire4165;
wire wire4166;
wire wire4167;
wire wire4168;
wire wire4169;
wire wire4171;
wire wire4172;
wire wire4174;
wire wire4175;
wire wire4176;
wire wire4177;
wire wire4178;
wire wire4179;
wire wire4180;
wire wire4181;
wire wire4183;
wire wire4184;
wire wire4186;
wire wire4188;
wire wire4196;
wire wire4213;
wire wire4218;
wire wire4227;
wire wire4230;
wire wire4246;
wire wire4247;
wire wire4249;
wire wire4250;
wire wire4251;
wire wire4257;
wire wire4262;
wire wire4263;
wire wire4291;
wire wire4406;
wire wire4492;
wire wire4493;
wire wire4494;
wire wire4497;
wire wire4506;
wire wire4523;
wire wire4524;
wire wire4525;
wire wire4526;
wire wire4527;
wire wire4528;
wire wire4530;
wire wire4531;
wire wire4532;
wire wire4536;
wire wire4549;
wire wire4551;
wire wire4553;
wire wire4554;
wire wire4555;
wire wire4557;
wire wire4558;
wire wire4560;
wire wire4561;
wire wire4562;
wire wire4563;
wire wire4564;
wire wire4566;
wire wire4567;
wire wire4568;
wire wire4569;
wire wire4571;
wire wire4572;
wire wire4575;
wire wire4576;
wire wire4577;
wire wire4578;
wire wire4579;
wire wire4581;
wire wire4582;
wire wire4583;
wire wire4584;
wire wire4585;
wire wire4586;
wire wire4587;
wire wire4590;
wire wire4591;
wire wire4593;
wire wire4596;
wire wire4597;
wire wire4598;
wire wire4599;
wire wire4601;
wire wire4602;
wire wire4606;
wire wire4607;
wire wire4608;
wire wire4611;
wire wire4614;
wire wire4615;
wire wire4616;
wire wire4617;
wire wire4618;
wire wire4620;
wire wire4621;
wire wire4622;
wire wire4624;
wire wire4626;
wire wire4628;
wire wire4629;
wire wire4643;
wire wire4648;
wire wire4657;
wire wire4667;
wire wire4669;
wire wire4673;
wire wire4680;
wire wire4682;
wire wire4683;
wire wire4686;
wire wire4688;
wire wire4690;
wire wire4693;
wire wire4694;
wire wire4697;
wire wire4698;
wire wire4702;
wire wire4710;
wire wire4711;
wire wire4712;
wire wire4713;
wire wire4714;
wire wire4716;
wire wire4717;
wire wire4719;
wire wire4725;
wire wire4734;
wire wire4736;
wire wire4738;
wire wire4741;
wire wire4742;
wire wire4744;
wire wire4746;
wire wire4747;
wire wire4749;
wire wire4750;
wire wire4751;
wire wire4752;
wire wire4753;
wire wire4755;
wire wire4756;
wire wire4757;
wire wire4758;
wire wire4759;
wire wire4761;
wire wire4763;
wire wire4764;
wire wire4766;
wire wire4768;
wire wire4770;
wire wire4771;
wire wire4773;
wire wire4774;
wire wire4776;
wire wire4777;
wire wire4779;
wire wire4780;
wire wire4783;
wire wire4785;
wire wire4786;
wire wire4788;
wire wire4792;
wire wire4793;
wire wire4794;
wire wire4795;
wire wire4796;
wire wire4797;
wire wire4798;
wire wire4800;
wire wire4802;
wire wire4803;
wire wire4806;
wire wire4807;
wire wire4828;
wire wire4834;
wire wire4849;
wire wire4852;
wire wire4853;
wire wire4854;
wire wire4855;
wire wire4856;
wire wire4857;
wire wire4858;
wire wire4861;
wire wire4862;
wire wire4863;
wire wire4864;
wire wire4866;
wire wire4867;
wire wire4868;
wire wire4870;
wire wire4871;
wire wire4872;
wire wire4873;
wire wire4875;
wire wire4876;
wire wire4877;
wire wire4879;
wire wire4881;
wire wire4882;
wire wire4883;
wire wire4884;
wire wire4885;
wire wire4886;
wire wire4888;
wire wire4890;
wire wire4891;
wire wire4892;
wire wire4893;
wire wire4894;
wire wire4902;
wire wire4916;
wire wire4918;
wire wire4920;
wire wire4921;
wire wire4922;
wire wire4923;
wire wire4924;
wire wire4926;
wire wire4928;
wire wire4929;
wire wire4930;
wire wire4931;
wire wire4932;
wire wire4933;
wire wire4935;
wire wire4937;
wire wire4938;
wire wire4939;
wire wire4941;
wire wire4942;
wire wire4943;
wire wire4944;
wire wire4946;
wire wire4947;
wire wire4948;
wire wire4950;
wire wire4951;
wire wire4952;
wire wire4978;
wire wire4986;
wire wire4988;
wire wire4989;
wire wire4990;
wire wire4991;
wire wire4992;
wire wire4993;
wire wire4995;
wire wire4997;
wire wire4998;
wire wire4999;
wire wire5000;
wire wire5001;
wire wire5002;
wire wire5003;
wire wire5005;
wire wire5006;
wire wire5007;
wire wire5008;
wire wire5010;
wire wire5011;
wire wire5012;
wire wire5014;
wire wire5016;
wire wire5017;
wire wire5018;
wire wire5019;
wire wire5020;
wire wire5021;
wire wire5023;
wire wire5025;
wire wire5026;
wire wire5027;
wire wire5028;
wire wire5029;
wire wire5031;
wire wire5033;
wire wire5034;
wire wire5035;
wire wire5036;
wire wire5037;
wire wire5038;
wire wire5040;
wire wire5042;
wire wire5043;
wire wire5044;
wire wire5045;
wire wire5046;
wire wire5047;
wire wire5057;
wire wire5058;
wire wire5063;
wire wire5068;
wire wire5073;
wire wire5088;
wire wire5091;
wire wire5094;
wire wire5096;
wire wire5097;
wire wire5098;
wire wire5106;
wire wire5113;
wire wire5116;
wire wire5117;
wire wire5118;
wire wire5121;
wire wire5123;
wire wire5124;
wire wire5125;
wire wire5126;
wire wire5132;
wire wire5133;
wire wire5139;
wire wire5143;
wire wire5145;
wire wire5157;
wire wire5158;
wire wire5164;
wire wire5166;
wire wire5171;
wire wire5172;
wire wire5182;
wire wire5184;
wire wire5185;
wire wire5186;
wire wire5190;
wire wire5192;
wire wire5194;
wire wire5196;
wire wire5197;
wire wire5201;
wire wire5203;
wire wire5205;
wire wire5206;
wire wire5208;
wire wire5211;
wire wire5212;
wire wire5213;
wire wire5218;
wire wire5221;
wire wire5222;
wire wire5223;
wire wire5228;
wire wire5230;
wire wire5231;
wire wire5232;
wire wire5235;
wire wire5237;
wire wire5238;
wire wire5239;
wire wire5241;
wire wire5243;
wire wire5245;
wire wire5247;
wire wire5248;
wire wire5250;
wire wire5254;
wire wire5257;
wire wire5258;
wire wire5259;
wire wire5261;
wire wire5263;
wire wire5265;
wire wire5266;
wire wire5271;
wire wire5272;
wire wire5273;
wire wire5274;
wire wire5275;
wire wire5277;
wire wire5283;
wire wire5286;
wire wire5287;
wire wire5288;
wire wire5289;
wire wire5290;
wire wire5291;
wire wire5292;
wire wire5295;
wire wire5297;
wire wire5298;
wire wire5299;
wire wire5313;
wire wire5320;
wire wire5322;
wire wire5323;
wire wire5325;
wire wire5327;
wire wire5329;
wire wire5331;
wire wire5332;
wire wire5334;
wire wire5344;
wire wire5346;
wire wire5349;
wire wire5350;
wire wire5353;
wire wire5355;
wire wire5358;
wire wire5363;
wire wire5368;
wire wire5385;
wire wire5389;
wire wire5398;
wire wire5403;
wire wire5407;
wire wire5409;
wire wire5410;
wire wire5411;
wire wire5413;
wire wire5418;
wire wire5426;
wire wire5427;
wire wire5428;
wire wire5430;
wire wire5431;
wire wire5432;
wire wire5433;
wire wire5434;
wire wire5436;
wire wire5437;
wire wire5438;
wire wire5440;
wire wire5441;
wire wire5443;
wire wire5451;
wire wire5452;
wire wire5453;
wire wire5455;
wire wire5456;
wire wire5457;
wire wire5464;
wire wire5467;
wire wire5468;
wire wire5471;
wire wire5472;
wire wire5473;
wire wire5476;
wire wire5479;
wire wire5483;
wire wire5484;
wire wire5485;
wire wire5486;
wire wire5487;
wire wire5488;
wire wire5490;
wire wire5492;
wire wire5493;
wire wire5496;
wire wire5497;
wire wire5498;
wire wire5499;
wire wire5500;
wire wire5501;
wire wire5502;
wire wire5503;
wire wire5506;
wire wire5507;
wire wire5509;
wire wire5513;
wire wire5514;
wire wire5520;
wire wire5522;
wire wire5528;
wire wire5582;
wire wire17517;
wire wire17519;
wire wire17520;
wire wire17521;
wire wire17522;
wire wire17523;
wire wire17524;
wire wire17525;
wire wire17527;
wire wire17528;
wire wire17529;
wire wire17530;
wire wire17532;
wire wire17533;
wire wire17534;
wire wire17535;
wire wire17536;
wire wire17537;
wire wire17538;
wire wire17540;
wire wire17541;
wire wire17542;
wire wire17543;
wire wire17545;
wire wire17546;
wire wire17547;
wire wire17555;
wire wire17556;
wire wire17557;
wire wire17558;
wire wire17562;
wire wire17564;
wire wire17566;
wire wire17568;
wire wire17572;
wire wire17574;
wire wire17576;
wire wire17577;
wire wire17580;
wire wire17582;
wire wire17593;
wire wire17594;
wire wire17595;
wire wire17597;
wire wire17599;
wire wire17600;
wire wire17601;
wire wire17602;
wire wire17603;
wire wire17605;
wire wire17606;
wire wire17607;
wire wire17608;
wire wire17610;
wire wire17615;
wire wire17616;
wire wire17617;
wire wire17621;
wire wire17626;
wire wire17627;
wire wire17628;
wire wire17631;
wire wire17638;
wire wire17639;
wire wire17640;
wire wire17641;
wire wire17642;
wire wire17647;
wire wire17649;
wire wire17650;
wire wire17652;
wire wire17654;
wire wire17657;
wire wire17658;
wire wire17659;
wire wire17660;
wire wire17662;
wire wire17668;
wire wire17670;
wire wire17671;
wire wire17672;
wire wire17673;
wire wire17678;
wire wire17688;
wire wire17689;
wire wire17690;
wire wire17691;
wire wire17694;
wire wire17695;
wire wire17696;
wire wire17698;
wire wire17699;
wire wire17703;
wire wire17704;
wire wire17705;
wire wire17709;
wire wire17710;
wire wire17711;
wire wire17712;
wire wire17714;
wire wire17715;
wire wire17716;
wire wire17717;
wire wire17718;
wire wire17719;
wire wire17720;
wire wire17722;
wire wire17724;
wire wire17727;
wire wire17728;
wire wire17731;
wire wire17738;
wire wire17742;
wire wire17743;
wire wire17745;
wire wire17746;
wire wire17748;
wire wire17749;
wire wire17753;
wire wire17754;
wire wire17756;
wire wire17757;
wire wire17758;
wire wire17759;
wire wire17763;
wire wire17764;
wire wire17768;
wire wire17769;
wire wire17770;
wire wire17771;
wire wire17774;
wire wire17776;
wire wire17780;
wire wire17781;
wire wire17784;
wire wire17785;
wire wire17787;
wire wire17792;
wire wire17793;
wire wire17796;
wire wire17797;
wire wire17801;
wire wire17805;
wire wire17808;
wire wire17809;
wire wire17813;
wire wire17826;
wire wire17829;
wire wire17830;
wire wire17833;
wire wire17834;
wire wire17836;
wire wire17837;
wire wire17841;
wire wire17842;
wire wire17844;
wire wire17845;
wire wire17846;
wire wire17865;
wire wire17868;
wire wire17871;
wire wire17873;
wire wire17875;
wire wire17877;
wire wire17880;
wire wire17883;
wire wire17885;
wire wire17887;
wire wire17889;
wire wire17891;
wire wire17894;
wire wire17896;
wire wire17898;
wire wire17900;
wire wire17901;
wire wire17902;
wire wire17903;
wire wire17904;
wire wire17906;
wire wire17909;
wire wire17911;
wire wire17913;
wire wire17915;
wire wire17917;
wire wire17920;
wire wire17924;
wire wire17925;
wire wire17926;
wire wire17927;
wire wire17928;
wire wire17932;
wire wire17937;
wire wire17939;
wire wire17941;
wire wire17943;
wire wire17946;
wire wire17949;
wire wire17951;
wire wire17953;
wire wire17955;
wire wire17958;
wire wire17961;
wire wire17963;
wire wire17964;
wire wire17965;
wire wire17966;
wire wire17969;
wire wire17979;
wire wire17981;
wire wire17984;
wire wire17987;
wire wire17989;
wire wire17991;
wire wire17993;
wire wire17996;
wire wire17998;
wire wire18001;
wire wire18003;
wire wire18005;
wire wire18008;
wire wire18010;
wire wire18013;
wire wire18014;
wire wire18015;
wire wire18016;
wire wire18017;
wire wire18037;
wire wire18039;
wire wire18040;
wire wire18043;
wire wire18047;
wire wire18049;
wire wire18050;
wire wire18051;
wire wire18052;
wire wire18056;
wire wire18057;
wire wire18060;
wire wire18068;
wire wire18069;
wire wire18070;
wire wire18071;
wire wire18073;
wire wire18078;
wire wire18079;
wire wire18080;
wire wire18114;
wire wire18115;
wire wire18117;
wire wire18120;
wire wire18124;
wire wire18125;
wire wire18127;
wire wire18128;
wire wire18130;
wire wire18134;
wire wire18135;
wire wire18144;
wire wire18145;
wire wire18146;
wire wire18147;
wire wire18148;
wire wire18153;
wire wire18160;
wire wire18161;
wire wire18162;
wire wire18163;
wire wire18164;
wire wire18170;
wire wire18171;
wire wire18172;
wire wire18189;
wire wire18190;
wire wire18192;
wire wire18196;
wire wire18201;
wire wire18202;
wire wire18203;
wire wire18208;
wire wire18209;
wire wire18217;
wire wire18218;
wire wire18219;
wire wire18221;
wire wire18222;
wire wire18226;
wire wire18234;
wire wire18235;
wire wire18236;
wire wire18237;
wire wire18238;
wire wire18242;
wire wire18244;
wire wire18245;
wire wire18253;
wire wire18261;
wire wire18262;
wire wire18263;
wire wire18264;
wire wire18265;
wire wire18270;
wire wire18276;
wire wire18277;
wire wire18278;
wire wire18279;
wire wire18280;
wire wire18286;
wire wire18287;
wire wire18288;
wire wire18291;
wire wire18300;
wire wire18301;
wire wire18302;
wire wire18303;
wire wire18304;
wire wire18309;
wire wire18310;
wire wire18312;
wire wire18315;
wire wire18316;
wire wire18320;
wire wire18327;
wire wire18328;
wire wire18329;
wire wire18330;
wire wire18331;
wire wire18336;
wire wire18338;
wire wire18339;
wire wire18342;
wire wire18343;
wire wire18353;
wire wire18354;
wire wire18355;
wire wire18356;
wire wire18357;
wire wire18362;
wire wire18369;
wire wire18370;
wire wire18372;
wire wire18373;
wire wire18374;
wire wire18379;
wire wire18380;
wire wire18381;
wire wire18385;
wire wire18386;
wire wire18401;
wire wire18402;
wire wire18403;
wire wire18406;
wire wire18408;
wire wire18414;
wire wire18416;
wire wire18417;
wire wire18421;
wire wire18427;
wire wire18429;
wire wire18430;
wire wire18445;
wire wire18446;
wire wire18447;
wire wire18451;
wire wire18455;
wire wire18456;
wire wire18457;
wire wire18458;
wire wire18459;
wire wire18463;
wire wire18470;
wire wire18471;
wire wire18472;
wire wire18476;
wire wire18477;
wire wire18479;
wire wire18481;
wire wire18487;
wire wire18489;
wire wire18490;
wire wire18491;
wire wire18492;
wire wire18497;
wire wire18505;
wire wire18507;
wire wire18508;
wire wire18511;
wire wire18512;
wire wire18513;
wire wire18517;
wire wire18522;
wire wire18523;
wire wire18524;
wire wire18534;
wire wire18535;
wire wire18536;
wire wire18539;
wire wire18548;
wire wire18549;
wire wire18550;
wire wire18553;
wire wire18554;
wire wire18556;
wire wire18559;
wire wire18564;
wire wire18565;
wire wire18566;
wire wire18574;
wire wire18575;
wire wire18576;
wire wire18577;
wire wire18578;
wire wire18583;
wire wire18591;
wire wire18592;
wire wire18593;
wire wire18598;
wire wire18599;
wire wire18607;
wire wire18608;
wire wire18609;
wire wire18611;
wire wire18612;
wire wire18616;
wire wire18617;
wire wire18619;
wire wire18622;
wire wire18627;
wire wire18628;
wire wire18629;
wire wire18637;
wire wire18638;
wire wire18639;
wire wire18640;
wire wire18641;
wire wire18646;
wire wire18653;
wire wire18654;
wire wire18655;
wire wire18658;
wire wire18659;
wire wire18666;
wire wire18667;
wire wire18668;
wire wire18669;
wire wire18670;
wire wire18674;
wire wire18675;
wire wire18676;
wire wire18679;
wire wire18684;
wire wire18685;
wire wire18686;
wire wire18695;
wire wire18696;
wire wire18697;
wire wire18706;
wire wire18707;
wire wire18708;
wire wire18711;
wire wire18712;
wire wire18714;
wire wire18721;
wire wire18722;
wire wire18723;
wire wire18724;
wire wire18725;
wire wire18729;
wire wire18734;
wire wire18735;
wire wire18736;
wire wire18739;
wire wire18743;
wire wire18744;
wire wire18745;
wire wire18746;
wire wire18747;
wire wire18751;
wire wire18758;
wire wire18759;
wire wire18760;
wire wire18763;
wire wire18764;
wire wire18766;
wire wire18773;
wire wire18774;
wire wire18775;
wire wire18776;
wire wire18777;
wire wire18781;
wire wire18783;
wire wire18784;
wire wire18785;
wire wire18786;
wire wire18789;
wire wire18790;
wire wire18792;
wire wire18793;
wire wire18795;
wire wire18796;
wire wire18797;
wire wire18798;
wire wire18799;
wire wire18804;
wire wire18805;
wire wire18806;
wire wire18807;
wire wire18808;
wire wire18813;
wire wire18814;
wire wire18815;
wire wire18816;
wire wire18819;
wire wire18820;
wire wire18821;
wire wire18822;
wire wire18823;
wire wire18828;
wire wire18829;
wire wire18830;
wire wire18832;
wire wire18833;
wire wire18834;
wire wire18835;
wire wire18836;
wire wire18837;
wire wire18838;
wire wire18839;
wire wire18842;
wire wire18843;
wire wire18845;
wire wire18851;
wire wire18852;
wire wire18853;
wire wire18854;
wire wire18855;
wire wire18860;
wire wire18862;
wire wire18865;
wire wire18866;
wire wire18867;
wire wire18868;
wire wire18869;
wire wire18874;
wire wire18875;
wire wire18876;
wire wire18880;
wire wire18881;
wire wire18882;
wire wire18883;
wire wire18884;
wire wire18889;
wire wire18890;
wire wire18891;
wire wire18892;
wire wire18897;
wire wire18898;
wire wire18899;
wire wire18900;
wire wire18901;
wire wire18902;
wire wire18904;
wire wire18905;
wire wire18906;
wire wire18909;
wire wire18910;
wire wire18911;
wire wire18912;
wire wire18914;
wire wire18919;
wire wire18920;
wire wire18923;
wire wire18924;
wire wire18925;
wire wire18926;
wire wire18927;
wire wire18932;
wire wire18933;
wire wire18936;
wire wire18937;
wire wire18938;
wire wire18939;
wire wire18940;
wire wire18945;
wire wire18946;
wire wire18947;
wire wire18948;
wire wire18951;
wire wire18952;
wire wire18953;
wire wire18954;
wire wire18958;
wire wire18959;
wire wire18960;
wire wire18961;
wire wire18962;
wire wire18963;
wire wire18964;
wire wire18966;
wire wire18967;
wire wire18968;
wire wire18969;
wire wire18970;
wire wire18971;
wire wire18972;
wire wire18973;
wire wire18974;
wire wire18975;
wire wire18981;
wire wire18982;
wire wire18983;
wire wire18985;
wire wire18986;
wire wire18987;
wire wire18989;
wire wire18990;
wire wire18991;
wire wire18992;
wire wire18993;
wire wire18994;
wire wire18995;
wire wire18996;
wire wire18999;
wire wire19000;
wire wire19001;
wire wire19003;
wire wire19004;
wire wire19009;
wire wire19010;
wire wire19011;
wire wire19012;
wire wire19013;
wire wire19018;
wire wire19019;
wire wire19022;
wire wire19028;
wire wire19029;
wire wire19030;
wire wire19031;
wire wire19032;
wire wire19037;
wire wire19038;
wire wire19039;
wire wire19042;
wire wire19043;
wire wire19044;
wire wire19045;
wire wire19046;
wire wire19051;
wire wire19052;
wire wire19057;
wire wire19058;
wire wire19059;
wire wire19062;
wire wire19063;
wire wire19074;
wire wire19075;
wire wire19076;
wire wire19080;
wire wire19081;
wire wire19083;
wire wire19084;
wire wire19085;
wire wire19094;
wire wire19095;
wire wire19100;
wire wire19101;
wire wire19102;
wire wire19104;
wire wire19105;
wire wire19110;
wire wire19111;
wire wire19115;
wire wire19116;
wire wire19117;
wire wire19118;
wire wire19119;
wire wire19124;
wire wire19125;
wire wire19126;
wire wire19127;
wire wire19130;
wire wire19132;
wire wire19134;
wire wire19135;
wire wire19136;
wire wire19140;
wire wire19141;
wire wire19142;
wire wire19144;
wire wire19145;
wire wire19150;
wire wire19151;
wire wire19152;
wire wire19154;
wire wire19155;
wire wire19156;
wire wire19158;
wire wire19159;
wire wire19163;
wire wire19164;
reg ndout;

reg ppeakb_12_12_;

reg ppeakb_1_1_;

reg ppeaka_6_6_;

reg wire4295;

reg wire4310;

reg ppeaks_5_5_;

reg ppeakp_10_10_;

reg wire4355;

reg wire4370;

reg wire4385;

reg wire4400;

reg wire4415;

reg wire4430;

reg wire4445;

reg wire4460;

reg wire4475;

reg wire4490;

reg wire4505;

reg wire4520;

reg wire4535;

reg wire4550;

reg wire4565;

reg wire4580;

reg wire4595;

reg wire4610;

reg wire4625;

reg wire4640;

reg wire4655;

reg wire4670;

reg wire4700;

reg wire4715;

reg wire4730;

reg wire4745;

reg wire4760;

reg wire4775;

reg wire4790;

reg wire4805;

reg wire4820;

reg wire4835;

reg wire4850;

reg wire4865;

reg wire4880;

reg wire4895;

reg wire4910;

reg wire4925;

reg wire4940;

reg wire4955;

reg wire4970;

reg ppeakb_0_0_;

reg ppeaka_7_7_;

reg wire5015;

reg wire5030;

reg ppeaks_4_4_;

reg ppeakp_11_11_;

reg wire5075;

reg wire5090;

reg wire5105;

reg wire5120;

reg wire5135;

reg wire5150;

reg wire5165;

reg wire5180;

reg wire5195;

reg wire5210;

reg wire5225;

reg wire5240;

reg wire5255;

reg wire5270;

reg wire5285;

reg wire5300;

reg wire5315;

reg wire5330;

reg wire5345;

reg wire5360;

reg wire5375;

reg wire5390;

reg wire5405;

reg wire5420;

reg wire5435;

reg wire5450;

reg wire5465;

reg wire5480;

reg wire5495;

reg wire5510;

reg wire5525;

reg wire5540;

reg wire5555;

reg wire5570;

reg wire5600;

reg wire5615;

reg wire5630;

reg wire5645;

reg wire5660;

reg wire5675;

reg ppeakb_10_10_;

reg ppeaka_8_8_;

reg wire5720;

reg ppeaks_14_14_;

reg ppeaks_7_7_;

reg ppeakp_12_12_;

reg wire5780;

reg wire5795;

reg wire5810;

reg wire5825;

reg wire5840;

reg wire5855;

reg wire5870;

reg wire5885;

reg wire5900;

reg wire5915;

reg wire5930;

reg wire5945;

reg wire5960;

reg wire5975;

reg wire5990;

reg wire6005;

reg wire6020;

reg wire6035;

reg wire6050;

reg wire6065;

reg wire6080;

reg wire6095;

reg wire6110;

reg wire6125;

reg wire6140;

reg wire6155;

reg wire6170;

reg wire6185;

reg wire6200;

reg wire6215;

reg wire6230;

reg wire6245;

reg wire6260;

reg wire6275;

reg wire6290;

reg wire6305;

reg wire6320;

reg wire6335;

reg wire6350;

reg wire6365;

reg ppeakb_11_11_;

reg ppeakb_2_2_;

reg wire6410;

reg ppeaks_15_15_;

reg ppeaks_6_6_;

reg ppeakp_13_13_;

reg wire6470;

reg wire6485;

reg wire6500;

reg wire6515;

reg wire6530;

reg wire6545;

reg wire6560;

reg wire6575;

reg wire6590;

reg wire6605;

reg wire6620;

reg wire6635;

reg wire6650;

reg wire6665;

reg wire6680;

reg wire6695;

reg wire6710;

reg wire6725;

reg wire6740;

reg wire6755;

reg wire6770;

reg wire6785;

reg wire6815;

reg wire6830;

reg wire6845;

reg wire6860;

reg wire6875;

reg wire6890;

reg wire6905;

reg wire6920;

reg wire6935;

reg wire6950;

reg wire6965;

reg wire6980;

reg wire6995;

reg wire7010;

reg wire7025;

reg wire7055;

reg ppeaks_12_12_;

reg ppeaks_1_1_;

reg ppeakp_3_3_;

reg wire7115;

reg wire7130;

reg wire7145;

reg wire7160;

reg wire7175;

reg wire7190;

reg wire7205;

reg wire7220;

reg wire7235;

reg wire7250;

reg wire7265;

reg wire7280;

reg wire7295;

reg wire7310;

reg wire7325;

reg wire7340;

reg wire7355;

reg wire7370;

reg wire7385;

reg wire7400;

reg wire7415;

reg wire7430;

reg wire7445;

reg wire7460;

reg wire7475;

reg wire7490;

reg wire7505;

reg wire7520;

reg wire7535;

reg wire7550;

reg wire7565;

reg wire7580;

reg wire7595;

reg wire7625;

reg wire7640;

reg wire7655;

reg wire7670;

reg wire7685;

reg ppeaks_13_13_;

reg ppeakp_7_7_;

reg ppeakp_2_2_;

reg wire7745;

reg wire7760;

reg wire7775;

reg wire7790;

reg wire7805;

reg wire7820;

reg wire7835;

reg wire7850;

reg wire7865;

reg wire7880;

reg wire7895;

reg wire7910;

reg wire7925;

reg wire7940;

reg wire7955;

reg wire7970;

reg wire8000;

reg wire8015;

reg wire8030;

reg wire8045;

reg wire8060;

reg wire8075;

reg wire8090;

reg wire8105;

reg wire8120;

reg wire8135;

reg wire8150;

reg wire8165;

reg wire8180;

reg wire8195;

reg wire8210;

reg wire8225;

reg wire8240;

reg wire8255;

reg wire8285;

reg wire8300;

reg wire8315;

reg wire8330;

reg ppeaks_3_3_;

reg ppeakp_8_8_;

reg ppeakp_1_1_;

reg wire8390;

reg wire8405;

reg wire8420;

reg wire8435;

reg wire8450;

reg wire8465;

reg wire8480;

reg wire8495;

reg wire8510;

reg wire8525;

reg wire8540;

reg wire8555;

reg wire8570;

reg wire8585;

reg wire8600;

reg wire8615;

reg wire8630;

reg wire8645;

reg wire8660;

reg wire8675;

reg wire8690;

reg wire8705;

reg wire8720;

reg wire8735;

reg wire8750;

reg wire8765;

reg wire8780;

reg wire8810;

reg wire8825;

reg wire8840;

reg wire8855;

reg wire8870;

reg wire8885;

reg wire8900;

reg wire8915;

reg wire8930;

reg wire8945;

reg wire8960;

reg wire8975;

reg ppeaks_11_11_;

reg ppeaks_2_2_;

reg ppeakp_9_9_;

reg ppeakp_0_0_;

reg wire9050;

reg wire9065;

reg wire9080;

reg wire9095;

reg wire9110;

reg wire9125;

reg wire9140;

reg wire9155;

reg wire9170;

reg wire9185;

reg wire9200;

reg wire9215;

reg wire9230;

reg wire9245;

reg wire9260;

reg wire9275;

reg wire9290;

reg wire9305;

reg wire9320;

reg wire9335;

reg wire9350;

reg wire9365;

reg wire9380;

reg wire9395;

reg wire9410;

reg wire9440;

reg wire9455;

reg wire9470;

reg wire9485;

reg wire9500;

reg wire9515;

reg wire9530;

reg wire9545;

reg wire9560;

reg wire9575;

reg wire9590;

reg wire9605;

reg wire9620;

reg wire9635;

reg wire9650;

reg wire9665;

reg wire9680;

reg ppeaki_6_6_;

reg wire9710;

reg wire9725;

reg wire9740;

reg wire9770;

reg wire9785;

reg wire9800;

reg wire9815;

reg wire9830;

reg wire9845;

reg wire9860;

reg wire9875;

reg wire9890;

reg wire9905;

reg wire9920;

reg wire9935;

reg wire9950;

reg wire9980;

reg wire9995;

reg wire10010;

reg wire10025;

reg wire10040;

reg wire10055;

reg wire10070;

reg wire10085;

reg wire10100;

reg wire10115;

reg wire10130;

reg wire10145;

reg wire10175;

reg wire10190;

reg wire10205;

reg wire10220;

reg ppeaki_15_15_;

reg ppeaki_4_4_;

reg wire10265;

reg wire10280;

reg wire10310;

reg wire10325;

reg wire10340;

reg wire10355;

reg wire10370;

reg wire10400;

reg wire10415;

reg wire10430;

reg wire10445;

reg wire10460;

reg wire10475;

reg wire10490;

reg wire10505;

reg ppeaki_14_14_;

reg ppeaki_5_5_;

reg wire10550;

reg wire10565;

reg wire10580;

reg wire10595;

reg wire10610;

reg wire10625;

reg wire10655;

reg wire10670;

reg wire10685;

reg wire10700;

reg wire10715;

reg wire10730;

reg wire10745;

reg wire10760;

reg wire10775;

reg wire10790;

reg wire10805;

reg wire10820;

reg wire10850;

reg wire10865;

reg wire10880;

reg wire10895;

reg wire10925;

reg wire10940;

reg wire10955;

reg wire10970;

reg wire10985;

reg wire11015;

reg wire11030;

reg wire11045;

reg wire11060;

reg wire11075;

reg wire11090;

reg wire11120;

reg wire11135;

reg wire11150;

reg wire11165;

reg wire11180;

reg wire11195;

reg wire11210;

reg wire11225;

reg wire11240;

reg wire11255;

reg wire11270;

reg wire11285;

reg wire11300;

reg wire11315;

reg wire11330;

reg wire11345;

reg wire11375;

reg wire11390;

reg wire11405;

reg wire11420;

reg wire11435;

reg wire11450;

reg wire11465;

reg wire11480;

reg wire11495;

reg wire11510;

reg wire11525;

reg wire11540;

reg wire11555;

reg wire11570;

reg wire11585;

reg wire11600;

reg wire11615;

reg wire11630;

reg wire11645;

reg wire11660;

reg wire11675;

reg wire11690;

reg wire11705;

reg wire11720;

reg wire11735;

reg wire11750;

reg wire11765;

reg wire11780;

reg wire11795;

reg wire11810;

reg ppeaki_9_9_;

reg ppeakb_14_14_;

reg wire11885;

reg wire11900;

reg wire11915;

reg wire11930;

reg ppeaki_8_8_;

reg ppeakb_15_15_;

reg wire12005;

reg wire12020;

reg wire12035;

reg wire12050;

reg wire12065;

reg wire12080;

reg ppeaki_7_7_;

reg wire12125;

reg wire12140;

reg wire12155;

reg wire12170;

reg wire12185;

reg wire12200;

reg ppeakb_13_13_;

reg wire12245;

reg wire12260;

reg wire12275;

reg ppeaki_13_13_;

reg ppeaki_2_2_;

reg wire12335;

reg wire12350;

reg wire12365;

reg wire12380;

reg wire12395;

reg wire12410;

reg wire12425;

reg wire12440;

reg wire12455;

reg wire12470;

reg wire12485;

reg ppeaki_12_12_;

reg ppeaki_3_3_;

reg wire12545;

reg wire12560;

reg wire12575;

reg wire12590;

reg wire12605;

reg wire12620;

reg wire12635;

reg wire12650;

reg wire12665;

reg wire12680;

reg wire12695;

reg ppeaki_11_11_;

reg ppeaki_0_0_;

reg wire12770;

reg wire12800;

reg wire12815;

reg wire12830;

reg wire12845;

reg wire12860;

reg wire12875;

reg wire12890;

reg wire12905;

reg wire12920;

reg wire12935;

reg ppeaki_10_10_;

reg ppeaki_1_1_;

reg wire13010;

reg wire13025;

reg wire13040;

reg wire13055;

reg wire13070;

reg wire13085;

reg wire13100;

reg wire13115;

reg wire13130;

reg wire13160;

reg wire13175;

reg ppeakb_4_4_;

reg ppeaka_9_9_;

reg wire13220;

reg wire13235;

reg wire13250;

reg wire13265;

reg wire13280;

reg wire13295;

reg wire13310;

reg wire13325;

reg wire13340;

reg wire13355;

reg wire13370;

reg wire13385;

reg wire13400;

reg wire13415;

reg wire13430;

reg wire13445;

reg wire13460;

reg wire13475;

reg wire13490;

reg wire13505;

reg ppeakb_5_5_;

reg wire13550;

reg ppeakp_6_6_;

reg wire13580;

reg wire13595;

reg wire13610;

reg wire13625;

reg wire13640;

reg wire13655;

reg wire13670;

reg wire13685;

reg wire13700;

reg wire13715;

reg wire13730;

reg wire13745;

reg wire13775;

reg wire13790;

reg wire13805;

reg wire13820;

reg wire13835;

reg wire13850;

reg wire13865;

reg wire13880;

reg wire13895;

reg ppeaka_11_11_;

reg ppeaka_0_0_;

reg ppeakp_5_5_;

reg wire13955;

reg wire13970;

reg wire13985;

reg wire14000;

reg wire14015;

reg wire14030;

reg wire14045;

reg wire14060;

reg wire14075;

reg wire14090;

reg wire14105;

reg wire14120;

reg wire14135;

reg wire14150;

reg wire14165;

reg wire14180;

reg wire14210;

reg wire14225;

reg wire14240;

reg wire14255;

reg wire14270;

reg wire14285;

reg ppeakb_3_3_;

reg ppeaka_10_10_;

reg ppeaka_1_1_;

reg ppeakp_4_4_;

reg wire14360;

reg wire14375;

reg wire14390;

reg wire14405;

reg wire14420;

reg wire14435;

reg wire14450;

reg wire14465;

reg wire14480;

reg wire14495;

reg wire14510;

reg wire14525;

reg wire14540;

reg wire14555;

reg wire14570;

reg wire14585;

reg wire14600;

reg wire14615;

reg wire14630;

reg wire14660;

reg wire14675;

reg wire14690;

reg wire14705;

reg ppeakb_8_8_;

reg ppeaka_13_13_;

reg ppeaka_2_2_;

reg wire14765;

reg ppeaks_9_9_;

reg ppeakp_14_14_;

reg wire14810;

reg wire14825;

reg wire14840;

reg wire14855;

reg wire14870;

reg wire14885;

reg wire14900;

reg wire14915;

reg wire14930;

reg wire14960;

reg wire14975;

reg wire14990;

reg wire15005;

reg wire15020;

reg wire15035;

reg wire15050;

reg wire15065;

reg wire15080;

reg ppeakb_9_9_;

reg ppeaka_12_12_;

reg ppeaka_3_3_;

reg wire15140;

reg ppeaks_8_8_;

reg ppeakp_15_15_;

reg wire15185;

reg wire15200;

reg wire15215;

reg wire15230;

reg wire15245;

reg wire15260;

reg wire15275;

reg wire15290;

reg wire15305;

reg wire15320;

reg wire15335;

reg wire15350;

reg wire15365;

reg wire15380;

reg wire15395;

reg wire15410;

reg wire15425;

reg wire15440;

reg ppeakb_6_6_;

reg ppeaka_15_15_;

reg ppeaka_4_4_;

reg wire15500;

reg wire15515;

reg ppeaks_0_0_;

reg wire15545;

reg wire15560;

reg wire15575;

reg wire15590;

reg wire15605;

reg wire15620;

reg wire15635;

reg wire15650;

reg wire15665;

reg wire15680;

reg wire15695;

reg wire15710;

reg wire15725;

reg wire15755;

reg wire15770;

reg wire15785;

reg ppeakb_7_7_;

reg ppeaka_14_14_;

reg ppeaka_5_5_;

reg wire15845;

reg wire15860;

reg ppeaks_10_10_;

reg wire15890;

reg wire15905;

reg wire15920;

reg wire15935;

reg wire15950;

reg wire15965;

reg wire15980;

reg wire15995;

reg wire16010;

reg wire16025;

reg wire16040;

reg wire16055;

reg wire16070;

reg wire16085;

reg wire16100;

reg paddress_8_8_;

reg wire16907;

reg wire16920;

reg wire16933;

reg paddress_9_9_;

reg wire16959;

reg wire16972;

reg wire16985;

reg wire16998;

reg wire17011;

reg wire17024;

reg wire17037;

reg wire17050;

reg wire17063;

reg wire17076;

reg wire17089;

reg wire17102;

reg wire17115;

reg wire17128;

reg wire17141;

reg wire17154;

reg wire17167;

reg wire17180;

reg wire17193;

reg wire17206;

reg wire17219;

reg wire17232;

reg wire17245;

reg wire17258;

reg wire17271;

reg wire17284;

reg wire17297;

reg wire17310;

reg wire17323;

reg wire17336;

reg wire17349;

reg wire17362;

reg wire17375;

reg wire17388;

reg paddress_11_11_;

reg wire17414;

reg wire17427;

reg wire17453;

reg paddress_10_10_;

reg wire17479;

reg wire17492;

reg wire17505;

reg wire17518;

reg wire17531;

reg wire17544;

reg paddress_13_13_;

reg wire17570;

reg wire17583;

reg wire17596;

reg wire17609;

reg paddress_12_12_;

reg wire17635;

reg wire17648;

reg wire17661;

reg wire17674;

reg paddress_15_15_;

reg wire17700;

reg wire17713;

reg paddress_14_14_;

reg wire17739;

reg wire17752;

reg wire17765;

reg wire17778;

reg wire17791;

reg wire17804;

reg wire17817;

reg pwr_0_0_;

reg wire17843;

reg wire17856;

reg wire17869;

reg wire17882;

reg prd_0_0_;

reg wire17908;

reg wire17921;

reg wire17934;

reg wire17947;

reg wire17960;

reg wire17973;

reg wire17986;

reg wire17999;

reg wire18012;

reg wire18025;

reg wire18038;

reg pdn;

reg wire18064;

reg wire18077;

reg wire18090;

reg wire18103;

reg wire18116;

reg wire18129;

reg wire18142;

reg wire18155;

reg wire18168;

reg wire18181;

reg wire18194;

reg wire18207;

reg wire18220;

reg wire18233;

reg wire18246;

reg paddress_0_0_;

reg piack_0_0_;

reg wire18285;

reg wire18298;

reg wire18311;

reg paddress_1_1_;

reg wire18337;

reg wire18350;

reg wire18363;

reg wire18376;

reg wire18389;

reg paddress_2_2_;

reg wire18415;

reg wire18428;

reg wire18441;

reg paddress_3_3_;

reg wire18467;

reg wire18480;

reg wire18493;

reg wire18506;

reg paddress_4_4_;

reg paddress_5_5_;

reg wire18545;

reg paddress_6_6_;

reg wire18571;

reg wire18584;

reg wire18597;

reg wire18610;

reg paddress_7_7_;

reg wire18636;

always  @(posedge pclk)
	ndout<=wire4244;

 always  @(posedge pclk)
	ppeakb_12_12_<=wire4259;

 always  @(posedge pclk)
	ppeakb_1_1_<=wire4274;

 always  @(posedge pclk)
	ppeaka_6_6_<=wire4289;

 always  @(posedge pclk)
	wire4295<=wire4304;

 always  @(posedge pclk)
	wire4310<=wire4319;

 always  @(posedge pclk)
	ppeaks_5_5_<=wire4334;

 always  @(posedge pclk)
	ppeakp_10_10_<=wire4349;

 always  @(posedge pclk)
	wire4355<=wire4364;

 always  @(posedge pclk)
	wire4370<=wire4379;

 always  @(posedge pclk)
	wire4385<=wire4394;

 always  @(posedge pclk)
	wire4400<=wire4409;

 always  @(posedge pclk)
	wire4415<=wire4424;

 always  @(posedge pclk)
	wire4430<=wire4439;

 always  @(posedge pclk)
	wire4445<=wire4454;

 always  @(posedge pclk)
	wire4460<=wire4469;

 always  @(posedge pclk)
	wire4475<=wire4484;

 always  @(posedge pclk)
	wire4490<=wire4499;

 always  @(posedge pclk)
	wire4505<=wire4514;

 always  @(posedge pclk)
	wire4520<=wire4529;

 always  @(posedge pclk)
	wire4535<=wire4544;

 always  @(posedge pclk)
	wire4550<=wire4559;

 always  @(posedge pclk)
	wire4565<=wire4574;

 always  @(posedge pclk)
	wire4580<=wire4589;

 always  @(posedge pclk)
	wire4595<=wire4604;

 always  @(posedge pclk)
	wire4610<=wire4619;

 always  @(posedge pclk)
	wire4625<=wire4634;

 always  @(posedge pclk)
	wire4640<=wire4649;

 always  @(posedge pclk)
	wire4655<=wire4664;

 always  @(posedge pclk)
	wire4670<=wire4679;

 always  @(posedge pclk)
	wire4700<=wire4709;

 always  @(posedge pclk)
	wire4715<=wire4724;

 always  @(posedge pclk)
	wire4730<=wire4739;

 always  @(posedge pclk)
	wire4745<=wire4754;

 always  @(posedge pclk)
	wire4760<=wire4769;

 always  @(posedge pclk)
	wire4775<=wire4784;

 always  @(posedge pclk)
	wire4790<=wire4799;

 always  @(posedge pclk)
	wire4805<=wire4814;

 always  @(posedge pclk)
	wire4820<=wire4829;

 always  @(posedge pclk)
	wire4835<=wire4844;

 always  @(posedge pclk)
	wire4850<=wire4859;

 always  @(posedge pclk)
	wire4865<=wire4874;

 always  @(posedge pclk)
	wire4880<=wire4889;

 always  @(posedge pclk)
	wire4895<=wire4904;

 always  @(posedge pclk)
	wire4910<=wire4919;

 always  @(posedge pclk)
	wire4925<=wire4934;

 always  @(posedge pclk)
	wire4940<=wire4949;

 always  @(posedge pclk)
	wire4955<=wire4964;

 always  @(posedge pclk)
	wire4970<=wire4979;

 always  @(posedge pclk)
	ppeakb_0_0_<=wire4994;

 always  @(posedge pclk)
	ppeaka_7_7_<=wire5009;

 always  @(posedge pclk)
	wire5015<=wire5024;

 always  @(posedge pclk)
	wire5030<=wire5039;

 always  @(posedge pclk)
	ppeaks_4_4_<=wire5054;

 always  @(posedge pclk)
	ppeakp_11_11_<=wire5069;

 always  @(posedge pclk)
	wire5075<=wire5084;

 always  @(posedge pclk)
	wire5090<=wire5099;

 always  @(posedge pclk)
	wire5105<=wire5114;

 always  @(posedge pclk)
	wire5120<=wire5129;

 always  @(posedge pclk)
	wire5135<=wire5144;

 always  @(posedge pclk)
	wire5150<=wire5159;

 always  @(posedge pclk)
	wire5165<=wire5174;

 always  @(posedge pclk)
	wire5180<=wire5189;

 always  @(posedge pclk)
	wire5195<=wire5204;

 always  @(posedge pclk)
	wire5210<=wire5219;

 always  @(posedge pclk)
	wire5225<=wire5234;

 always  @(posedge pclk)
	wire5240<=wire5249;

 always  @(posedge pclk)
	wire5255<=wire5264;

 always  @(posedge pclk)
	wire5270<=wire5279;

 always  @(posedge pclk)
	wire5285<=wire5294;

 always  @(posedge pclk)
	wire5300<=wire5309;

 always  @(posedge pclk)
	wire5315<=wire5324;

 always  @(posedge pclk)
	wire5330<=wire5339;

 always  @(posedge pclk)
	wire5345<=wire5354;

 always  @(posedge pclk)
	wire5360<=wire5369;

 always  @(posedge pclk)
	wire5375<=wire5384;

 always  @(posedge pclk)
	wire5390<=wire5399;

 always  @(posedge pclk)
	wire5405<=wire5414;

 always  @(posedge pclk)
	wire5420<=wire5429;

 always  @(posedge pclk)
	wire5435<=wire5444;

 always  @(posedge pclk)
	wire5450<=wire5459;

 always  @(posedge pclk)
	wire5465<=wire5474;

 always  @(posedge pclk)
	wire5480<=wire5489;

 always  @(posedge pclk)
	wire5495<=wire5504;

 always  @(posedge pclk)
	wire5510<=wire5519;

 always  @(posedge pclk)
	wire5525<=wire5534;

 always  @(posedge pclk)
	wire5540<=wire5549;

 always  @(posedge pclk)
	wire5555<=wire5564;

 always  @(posedge pclk)
	wire5570<=wire5579;

 always  @(posedge pclk)
	wire5600<=wire5609;

 always  @(posedge pclk)
	wire5615<=wire5624;

 always  @(posedge pclk)
	wire5630<=wire5639;

 always  @(posedge pclk)
	wire5645<=wire5654;

 always  @(posedge pclk)
	wire5660<=wire5669;

 always  @(posedge pclk)
	wire5675<=wire5684;

 always  @(posedge pclk)
	ppeakb_10_10_<=wire5699;

 always  @(posedge pclk)
	ppeaka_8_8_<=wire5714;

 always  @(posedge pclk)
	wire5720<=wire5729;

 always  @(posedge pclk)
	ppeaks_14_14_<=wire5744;

 always  @(posedge pclk)
	ppeaks_7_7_<=wire5759;

 always  @(posedge pclk)
	ppeakp_12_12_<=wire5774;

 always  @(posedge pclk)
	wire5780<=wire5789;

 always  @(posedge pclk)
	wire5795<=wire5804;

 always  @(posedge pclk)
	wire5810<=wire5819;

 always  @(posedge pclk)
	wire5825<=wire5834;

 always  @(posedge pclk)
	wire5840<=wire5849;

 always  @(posedge pclk)
	wire5855<=wire5864;

 always  @(posedge pclk)
	wire5870<=wire5879;

 always  @(posedge pclk)
	wire5885<=wire5894;

 always  @(posedge pclk)
	wire5900<=wire5909;

 always  @(posedge pclk)
	wire5915<=wire5924;

 always  @(posedge pclk)
	wire5930<=wire5939;

 always  @(posedge pclk)
	wire5945<=wire5954;

 always  @(posedge pclk)
	wire5960<=wire5969;

 always  @(posedge pclk)
	wire5975<=wire5984;

 always  @(posedge pclk)
	wire5990<=wire5999;

 always  @(posedge pclk)
	wire6005<=wire6014;

 always  @(posedge pclk)
	wire6020<=wire6029;

 always  @(posedge pclk)
	wire6035<=wire6044;

 always  @(posedge pclk)
	wire6050<=wire6059;

 always  @(posedge pclk)
	wire6065<=wire6074;

 always  @(posedge pclk)
	wire6080<=wire6089;

 always  @(posedge pclk)
	wire6095<=wire6104;

 always  @(posedge pclk)
	wire6110<=wire6119;

 always  @(posedge pclk)
	wire6125<=wire6134;

 always  @(posedge pclk)
	wire6140<=wire6149;

 always  @(posedge pclk)
	wire6155<=wire6164;

 always  @(posedge pclk)
	wire6170<=wire6179;

 always  @(posedge pclk)
	wire6185<=wire6194;

 always  @(posedge pclk)
	wire6200<=wire6209;

 always  @(posedge pclk)
	wire6215<=wire6224;

 always  @(posedge pclk)
	wire6230<=wire6239;

 always  @(posedge pclk)
	wire6245<=wire6254;

 always  @(posedge pclk)
	wire6260<=wire6269;

 always  @(posedge pclk)
	wire6275<=wire6284;

 always  @(posedge pclk)
	wire6290<=wire6299;

 always  @(posedge pclk)
	wire6305<=wire6314;

 always  @(posedge pclk)
	wire6320<=wire6329;

 always  @(posedge pclk)
	wire6335<=wire6344;

 always  @(posedge pclk)
	wire6350<=wire6359;

 always  @(posedge pclk)
	wire6365<=wire6374;

 always  @(posedge pclk)
	ppeakb_11_11_<=wire6389;

 always  @(posedge pclk)
	ppeakb_2_2_<=wire6404;

 always  @(posedge pclk)
	wire6410<=wire6419;

 always  @(posedge pclk)
	ppeaks_15_15_<=wire6434;

 always  @(posedge pclk)
	ppeaks_6_6_<=wire6449;

 always  @(posedge pclk)
	ppeakp_13_13_<=wire6464;

 always  @(posedge pclk)
	wire6470<=wire6479;

 always  @(posedge pclk)
	wire6485<=wire6494;

 always  @(posedge pclk)
	wire6500<=wire6509;

 always  @(posedge pclk)
	wire6515<=wire6524;

 always  @(posedge pclk)
	wire6530<=wire6539;

 always  @(posedge pclk)
	wire6545<=wire6554;

 always  @(posedge pclk)
	wire6560<=wire6569;

 always  @(posedge pclk)
	wire6575<=wire6584;

 always  @(posedge pclk)
	wire6590<=wire6599;

 always  @(posedge pclk)
	wire6605<=wire6614;

 always  @(posedge pclk)
	wire6620<=wire6629;

 always  @(posedge pclk)
	wire6635<=wire6644;

 always  @(posedge pclk)
	wire6650<=wire6659;

 always  @(posedge pclk)
	wire6665<=wire6674;

 always  @(posedge pclk)
	wire6680<=wire6689;

 always  @(posedge pclk)
	wire6695<=wire6704;

 always  @(posedge pclk)
	wire6710<=wire6719;

 always  @(posedge pclk)
	wire6725<=wire6734;

 always  @(posedge pclk)
	wire6740<=wire6749;

 always  @(posedge pclk)
	wire6755<=wire6764;

 always  @(posedge pclk)
	wire6770<=wire6779;

 always  @(posedge pclk)
	wire6785<=wire6794;

 always  @(posedge pclk)
	wire6815<=wire6824;

 always  @(posedge pclk)
	wire6830<=wire6839;

 always  @(posedge pclk)
	wire6845<=wire6854;

 always  @(posedge pclk)
	wire6860<=wire6869;

 always  @(posedge pclk)
	wire6875<=wire6884;

 always  @(posedge pclk)
	wire6890<=wire6899;

 always  @(posedge pclk)
	wire6905<=wire6914;

 always  @(posedge pclk)
	wire6920<=wire6929;

 always  @(posedge pclk)
	wire6935<=wire6944;

 always  @(posedge pclk)
	wire6950<=wire6959;

 always  @(posedge pclk)
	wire6965<=wire6974;

 always  @(posedge pclk)
	wire6980<=wire6989;

 always  @(posedge pclk)
	wire6995<=wire7004;

 always  @(posedge pclk)
	wire7010<=wire7019;

 always  @(posedge pclk)
	wire7025<=wire7034;

 always  @(posedge pclk)
	wire7055<=wire7064;

 always  @(posedge pclk)
	ppeaks_12_12_<=wire7079;

 always  @(posedge pclk)
	ppeaks_1_1_<=wire7094;

 always  @(posedge pclk)
	ppeakp_3_3_<=wire7109;

 always  @(posedge pclk)
	wire7115<=wire7124;

 always  @(posedge pclk)
	wire7130<=wire7139;

 always  @(posedge pclk)
	wire7145<=wire7154;

 always  @(posedge pclk)
	wire7160<=wire7169;

 always  @(posedge pclk)
	wire7175<=wire7184;

 always  @(posedge pclk)
	wire7190<=wire7199;

 always  @(posedge pclk)
	wire7205<=wire7214;

 always  @(posedge pclk)
	wire7220<=wire7229;

 always  @(posedge pclk)
	wire7235<=wire7244;

 always  @(posedge pclk)
	wire7250<=wire7259;

 always  @(posedge pclk)
	wire7265<=wire7274;

 always  @(posedge pclk)
	wire7280<=wire7289;

 always  @(posedge pclk)
	wire7295<=wire7304;

 always  @(posedge pclk)
	wire7310<=wire7319;

 always  @(posedge pclk)
	wire7325<=wire7334;

 always  @(posedge pclk)
	wire7340<=wire7349;

 always  @(posedge pclk)
	wire7355<=wire7364;

 always  @(posedge pclk)
	wire7370<=wire7379;

 always  @(posedge pclk)
	wire7385<=wire7394;

 always  @(posedge pclk)
	wire7400<=wire7409;

 always  @(posedge pclk)
	wire7415<=wire7424;

 always  @(posedge pclk)
	wire7430<=wire7439;

 always  @(posedge pclk)
	wire7445<=wire7454;

 always  @(posedge pclk)
	wire7460<=wire7469;

 always  @(posedge pclk)
	wire7475<=wire7484;

 always  @(posedge pclk)
	wire7490<=wire7499;

 always  @(posedge pclk)
	wire7505<=wire7514;

 always  @(posedge pclk)
	wire7520<=wire7529;

 always  @(posedge pclk)
	wire7535<=wire7544;

 always  @(posedge pclk)
	wire7550<=wire7559;

 always  @(posedge pclk)
	wire7565<=wire7574;

 always  @(posedge pclk)
	wire7580<=wire7589;

 always  @(posedge pclk)
	wire7595<=wire7604;

 always  @(posedge pclk)
	wire7625<=wire7634;

 always  @(posedge pclk)
	wire7640<=wire7649;

 always  @(posedge pclk)
	wire7655<=wire7664;

 always  @(posedge pclk)
	wire7670<=wire7679;

 always  @(posedge pclk)
	wire7685<=wire7694;

 always  @(posedge pclk)
	ppeaks_13_13_<=wire7709;

 always  @(posedge pclk)
	ppeakp_7_7_<=wire7724;

 always  @(posedge pclk)
	ppeakp_2_2_<=wire7739;

 always  @(posedge pclk)
	wire7745<=wire7754;

 always  @(posedge pclk)
	wire7760<=wire7769;

 always  @(posedge pclk)
	wire7775<=wire7784;

 always  @(posedge pclk)
	wire7790<=wire7799;

 always  @(posedge pclk)
	wire7805<=wire7814;

 always  @(posedge pclk)
	wire7820<=wire7829;

 always  @(posedge pclk)
	wire7835<=wire7844;

 always  @(posedge pclk)
	wire7850<=wire7859;

 always  @(posedge pclk)
	wire7865<=wire7874;

 always  @(posedge pclk)
	wire7880<=wire7889;

 always  @(posedge pclk)
	wire7895<=wire7904;

 always  @(posedge pclk)
	wire7910<=wire7919;

 always  @(posedge pclk)
	wire7925<=wire7934;

 always  @(posedge pclk)
	wire7940<=wire7949;

 always  @(posedge pclk)
	wire7955<=wire7964;

 always  @(posedge pclk)
	wire7970<=wire7979;

 always  @(posedge pclk)
	wire8000<=wire8009;

 always  @(posedge pclk)
	wire8015<=wire8024;

 always  @(posedge pclk)
	wire8030<=wire8039;

 always  @(posedge pclk)
	wire8045<=wire8054;

 always  @(posedge pclk)
	wire8060<=wire8069;

 always  @(posedge pclk)
	wire8075<=wire8084;

 always  @(posedge pclk)
	wire8090<=wire8099;

 always  @(posedge pclk)
	wire8105<=wire8114;

 always  @(posedge pclk)
	wire8120<=wire8129;

 always  @(posedge pclk)
	wire8135<=wire8144;

 always  @(posedge pclk)
	wire8150<=wire8159;

 always  @(posedge pclk)
	wire8165<=wire8174;

 always  @(posedge pclk)
	wire8180<=wire8189;

 always  @(posedge pclk)
	wire8195<=wire8204;

 always  @(posedge pclk)
	wire8210<=wire8219;

 always  @(posedge pclk)
	wire8225<=wire8234;

 always  @(posedge pclk)
	wire8240<=wire8249;

 always  @(posedge pclk)
	wire8255<=wire8264;

 always  @(posedge pclk)
	wire8285<=wire8294;

 always  @(posedge pclk)
	wire8300<=wire8309;

 always  @(posedge pclk)
	wire8315<=wire8324;

 always  @(posedge pclk)
	wire8330<=wire8339;

 always  @(posedge pclk)
	ppeaks_3_3_<=wire8354;

 always  @(posedge pclk)
	ppeakp_8_8_<=wire8369;

 always  @(posedge pclk)
	ppeakp_1_1_<=wire8384;

 always  @(posedge pclk)
	wire8390<=wire8399;

 always  @(posedge pclk)
	wire8405<=wire8414;

 always  @(posedge pclk)
	wire8420<=wire8429;

 always  @(posedge pclk)
	wire8435<=wire8444;

 always  @(posedge pclk)
	wire8450<=wire8459;

 always  @(posedge pclk)
	wire8465<=wire8474;

 always  @(posedge pclk)
	wire8480<=wire8489;

 always  @(posedge pclk)
	wire8495<=wire8504;

 always  @(posedge pclk)
	wire8510<=wire8519;

 always  @(posedge pclk)
	wire8525<=wire8534;

 always  @(posedge pclk)
	wire8540<=wire8549;

 always  @(posedge pclk)
	wire8555<=wire8564;

 always  @(posedge pclk)
	wire8570<=wire8579;

 always  @(posedge pclk)
	wire8585<=wire8594;

 always  @(posedge pclk)
	wire8600<=wire8609;

 always  @(posedge pclk)
	wire8615<=wire8624;

 always  @(posedge pclk)
	wire8630<=wire8639;

 always  @(posedge pclk)
	wire8645<=wire8654;

 always  @(posedge pclk)
	wire8660<=wire8669;

 always  @(posedge pclk)
	wire8675<=wire8684;

 always  @(posedge pclk)
	wire8690<=wire8699;

 always  @(posedge pclk)
	wire8705<=wire8714;

 always  @(posedge pclk)
	wire8720<=wire8729;

 always  @(posedge pclk)
	wire8735<=wire8744;

 always  @(posedge pclk)
	wire8750<=wire8759;

 always  @(posedge pclk)
	wire8765<=wire8774;

 always  @(posedge pclk)
	wire8780<=wire8789;

 always  @(posedge pclk)
	wire8810<=wire8819;

 always  @(posedge pclk)
	wire8825<=wire8834;

 always  @(posedge pclk)
	wire8840<=wire8849;

 always  @(posedge pclk)
	wire8855<=wire8864;

 always  @(posedge pclk)
	wire8870<=wire8879;

 always  @(posedge pclk)
	wire8885<=wire8894;

 always  @(posedge pclk)
	wire8900<=wire8909;

 always  @(posedge pclk)
	wire8915<=wire8924;

 always  @(posedge pclk)
	wire8930<=wire8939;

 always  @(posedge pclk)
	wire8945<=wire8954;

 always  @(posedge pclk)
	wire8960<=wire8969;

 always  @(posedge pclk)
	wire8975<=wire8984;

 always  @(posedge pclk)
	ppeaks_11_11_<=wire8999;

 always  @(posedge pclk)
	ppeaks_2_2_<=wire9014;

 always  @(posedge pclk)
	ppeakp_9_9_<=wire9029;

 always  @(posedge pclk)
	ppeakp_0_0_<=wire9044;

 always  @(posedge pclk)
	wire9050<=wire9059;

 always  @(posedge pclk)
	wire9065<=wire9074;

 always  @(posedge pclk)
	wire9080<=wire9089;

 always  @(posedge pclk)
	wire9095<=wire9104;

 always  @(posedge pclk)
	wire9110<=wire9119;

 always  @(posedge pclk)
	wire9125<=wire9134;

 always  @(posedge pclk)
	wire9140<=wire9149;

 always  @(posedge pclk)
	wire9155<=wire9164;

 always  @(posedge pclk)
	wire9170<=wire9179;

 always  @(posedge pclk)
	wire9185<=wire9194;

 always  @(posedge pclk)
	wire9200<=wire9209;

 always  @(posedge pclk)
	wire9215<=wire9224;

 always  @(posedge pclk)
	wire9230<=wire9239;

 always  @(posedge pclk)
	wire9245<=wire9254;

 always  @(posedge pclk)
	wire9260<=wire9269;

 always  @(posedge pclk)
	wire9275<=wire9284;

 always  @(posedge pclk)
	wire9290<=wire9299;

 always  @(posedge pclk)
	wire9305<=wire9314;

 always  @(posedge pclk)
	wire9320<=wire9329;

 always  @(posedge pclk)
	wire9335<=wire9344;

 always  @(posedge pclk)
	wire9350<=wire9359;

 always  @(posedge pclk)
	wire9365<=wire9374;

 always  @(posedge pclk)
	wire9380<=wire9389;

 always  @(posedge pclk)
	wire9395<=wire9404;

 always  @(posedge pclk)
	wire9410<=wire9419;

 always  @(posedge pclk)
	wire9440<=wire9449;

 always  @(posedge pclk)
	wire9455<=wire9464;

 always  @(posedge pclk)
	wire9470<=wire9479;

 always  @(posedge pclk)
	wire9485<=wire9494;

 always  @(posedge pclk)
	wire9500<=wire9509;

 always  @(posedge pclk)
	wire9515<=wire9524;

 always  @(posedge pclk)
	wire9530<=wire9539;

 always  @(posedge pclk)
	wire9545<=wire9554;

 always  @(posedge pclk)
	wire9560<=wire9569;

 always  @(posedge pclk)
	wire9575<=wire9584;

 always  @(posedge pclk)
	wire9590<=wire9599;

 always  @(posedge pclk)
	wire9605<=wire9614;

 always  @(posedge pclk)
	wire9620<=wire9629;

 always  @(posedge pclk)
	wire9635<=wire9644;

 always  @(posedge pclk)
	wire9650<=wire9659;

 always  @(posedge pclk)
	wire9665<=wire9674;

 always  @(posedge pclk)
	wire9680<=wire9689;

 always  @(posedge pclk)
	ppeaki_6_6_<=wire9704;

 always  @(posedge pclk)
	wire9710<=wire9719;

 always  @(posedge pclk)
	wire9725<=wire9734;

 always  @(posedge pclk)
	wire9740<=wire9749;

 always  @(posedge pclk)
	wire9770<=wire9779;

 always  @(posedge pclk)
	wire9785<=wire9794;

 always  @(posedge pclk)
	wire9800<=wire9809;

 always  @(posedge pclk)
	wire9815<=wire9824;

 always  @(posedge pclk)
	wire9830<=wire9839;

 always  @(posedge pclk)
	wire9845<=wire9854;

 always  @(posedge pclk)
	wire9860<=wire9869;

 always  @(posedge pclk)
	wire9875<=wire9884;

 always  @(posedge pclk)
	wire9890<=wire9899;

 always  @(posedge pclk)
	wire9905<=wire9914;

 always  @(posedge pclk)
	wire9920<=wire9929;

 always  @(posedge pclk)
	wire9935<=wire9944;

 always  @(posedge pclk)
	wire9950<=wire9959;

 always  @(posedge pclk)
	wire9980<=wire9989;

 always  @(posedge pclk)
	wire9995<=wire10004;

 always  @(posedge pclk)
	wire10010<=wire10019;

 always  @(posedge pclk)
	wire10025<=wire10034;

 always  @(posedge pclk)
	wire10040<=wire10049;

 always  @(posedge pclk)
	wire10055<=wire10064;

 always  @(posedge pclk)
	wire10070<=wire10079;

 always  @(posedge pclk)
	wire10085<=wire10094;

 always  @(posedge pclk)
	wire10100<=wire10109;

 always  @(posedge pclk)
	wire10115<=wire10124;

 always  @(posedge pclk)
	wire10130<=wire10139;

 always  @(posedge pclk)
	wire10145<=wire10154;

 always  @(posedge pclk)
	wire10175<=wire10184;

 always  @(posedge pclk)
	wire10190<=wire10199;

 always  @(posedge pclk)
	wire10205<=wire10214;

 always  @(posedge pclk)
	wire10220<=wire10229;

 always  @(posedge pclk)
	ppeaki_15_15_<=wire10244;

 always  @(posedge pclk)
	ppeaki_4_4_<=wire10259;

 always  @(posedge pclk)
	wire10265<=wire10274;

 always  @(posedge pclk)
	wire10280<=wire10289;

 always  @(posedge pclk)
	wire10310<=wire10319;

 always  @(posedge pclk)
	wire10325<=wire10334;

 always  @(posedge pclk)
	wire10340<=wire10349;

 always  @(posedge pclk)
	wire10355<=wire10364;

 always  @(posedge pclk)
	wire10370<=wire10379;

 always  @(posedge pclk)
	wire10400<=wire10409;

 always  @(posedge pclk)
	wire10415<=wire10424;

 always  @(posedge pclk)
	wire10430<=wire10439;

 always  @(posedge pclk)
	wire10445<=wire10454;

 always  @(posedge pclk)
	wire10460<=wire10469;

 always  @(posedge pclk)
	wire10475<=wire10484;

 always  @(posedge pclk)
	wire10490<=wire10499;

 always  @(posedge pclk)
	wire10505<=wire10514;

 always  @(posedge pclk)
	ppeaki_14_14_<=wire10529;

 always  @(posedge pclk)
	ppeaki_5_5_<=wire10544;

 always  @(posedge pclk)
	wire10550<=wire10559;

 always  @(posedge pclk)
	wire10565<=wire10574;

 always  @(posedge pclk)
	wire10580<=wire10589;

 always  @(posedge pclk)
	wire10595<=wire10604;

 always  @(posedge pclk)
	wire10610<=wire10619;

 always  @(posedge pclk)
	wire10625<=wire10634;

 always  @(posedge pclk)
	wire10655<=wire10664;

 always  @(posedge pclk)
	wire10670<=wire10679;

 always  @(posedge pclk)
	wire10685<=wire10694;

 always  @(posedge pclk)
	wire10700<=wire10709;

 always  @(posedge pclk)
	wire10715<=wire10724;

 always  @(posedge pclk)
	wire10730<=wire10739;

 always  @(posedge pclk)
	wire10745<=wire10754;

 always  @(posedge pclk)
	wire10760<=wire10769;

 always  @(posedge pclk)
	wire10775<=wire10784;

 always  @(posedge pclk)
	wire10790<=wire10799;

 always  @(posedge pclk)
	wire10805<=wire10814;

 always  @(posedge pclk)
	wire10820<=wire10829;

 always  @(posedge pclk)
	wire10850<=wire10859;

 always  @(posedge pclk)
	wire10865<=wire10874;

 always  @(posedge pclk)
	wire10880<=wire10889;

 always  @(posedge pclk)
	wire10895<=wire10904;

 always  @(posedge pclk)
	wire10925<=wire10934;

 always  @(posedge pclk)
	wire10940<=wire10949;

 always  @(posedge pclk)
	wire10955<=wire10964;

 always  @(posedge pclk)
	wire10970<=wire10979;

 always  @(posedge pclk)
	wire10985<=wire10994;

 always  @(posedge pclk)
	wire11015<=wire11024;

 always  @(posedge pclk)
	wire11030<=wire11039;

 always  @(posedge pclk)
	wire11045<=wire11054;

 always  @(posedge pclk)
	wire11060<=wire11069;

 always  @(posedge pclk)
	wire11075<=wire11084;

 always  @(posedge pclk)
	wire11090<=wire11099;

 always  @(posedge pclk)
	wire11120<=wire11129;

 always  @(posedge pclk)
	wire11135<=wire11144;

 always  @(posedge pclk)
	wire11150<=wire11159;

 always  @(posedge pclk)
	wire11165<=wire11174;

 always  @(posedge pclk)
	wire11180<=wire11189;

 always  @(posedge pclk)
	wire11195<=wire11204;

 always  @(posedge pclk)
	wire11210<=wire11219;

 always  @(posedge pclk)
	wire11225<=wire11234;

 always  @(posedge pclk)
	wire11240<=wire11249;

 always  @(posedge pclk)
	wire11255<=wire11264;

 always  @(posedge pclk)
	wire11270<=wire11279;

 always  @(posedge pclk)
	wire11285<=wire11294;

 always  @(posedge pclk)
	wire11300<=wire11309;

 always  @(posedge pclk)
	wire11315<=wire11324;

 always  @(posedge pclk)
	wire11330<=wire11339;

 always  @(posedge pclk)
	wire11345<=wire11354;

 always  @(posedge pclk)
	wire11375<=wire11384;

 always  @(posedge pclk)
	wire11390<=wire11399;

 always  @(posedge pclk)
	wire11405<=wire11414;

 always  @(posedge pclk)
	wire11420<=wire11429;

 always  @(posedge pclk)
	wire11435<=wire11444;

 always  @(posedge pclk)
	wire11450<=wire11459;

 always  @(posedge pclk)
	wire11465<=wire11474;

 always  @(posedge pclk)
	wire11480<=wire11489;

 always  @(posedge pclk)
	wire11495<=wire11504;

 always  @(posedge pclk)
	wire11510<=wire11519;

 always  @(posedge pclk)
	wire11525<=wire11534;

 always  @(posedge pclk)
	wire11540<=wire11549;

 always  @(posedge pclk)
	wire11555<=wire11564;

 always  @(posedge pclk)
	wire11570<=wire11579;

 always  @(posedge pclk)
	wire11585<=wire11594;

 always  @(posedge pclk)
	wire11600<=wire11609;

 always  @(posedge pclk)
	wire11615<=wire11624;

 always  @(posedge pclk)
	wire11630<=wire11639;

 always  @(posedge pclk)
	wire11645<=wire11654;

 always  @(posedge pclk)
	wire11660<=wire11669;

 always  @(posedge pclk)
	wire11675<=wire11684;

 always  @(posedge pclk)
	wire11690<=wire11699;

 always  @(posedge pclk)
	wire11705<=wire11714;

 always  @(posedge pclk)
	wire11720<=wire11729;

 always  @(posedge pclk)
	wire11735<=wire11744;

 always  @(posedge pclk)
	wire11750<=wire11759;

 always  @(posedge pclk)
	wire11765<=wire11774;

 always  @(posedge pclk)
	wire11780<=wire11789;

 always  @(posedge pclk)
	wire11795<=wire11804;

 always  @(posedge pclk)
	wire11810<=wire11819;

 always  @(posedge pclk)
	ppeaki_9_9_<=wire11864;

 always  @(posedge pclk)
	ppeakb_14_14_<=wire11879;

 always  @(posedge pclk)
	wire11885<=wire11894;

 always  @(posedge pclk)
	wire11900<=wire11909;

 always  @(posedge pclk)
	wire11915<=wire11924;

 always  @(posedge pclk)
	wire11930<=wire11939;

 always  @(posedge pclk)
	ppeaki_8_8_<=wire11984;

 always  @(posedge pclk)
	ppeakb_15_15_<=wire11999;

 always  @(posedge pclk)
	wire12005<=wire12014;

 always  @(posedge pclk)
	wire12020<=wire12029;

 always  @(posedge pclk)
	wire12035<=wire12044;

 always  @(posedge pclk)
	wire12050<=wire12059;

 always  @(posedge pclk)
	wire12065<=wire12074;

 always  @(posedge pclk)
	wire12080<=wire12089;

 always  @(posedge pclk)
	ppeaki_7_7_<=wire12119;

 always  @(posedge pclk)
	wire12125<=wire12134;

 always  @(posedge pclk)
	wire12140<=wire12149;

 always  @(posedge pclk)
	wire12155<=wire12164;

 always  @(posedge pclk)
	wire12170<=wire12179;

 always  @(posedge pclk)
	wire12185<=wire12194;

 always  @(posedge pclk)
	wire12200<=wire12209;

 always  @(posedge pclk)
	ppeakb_13_13_<=wire12239;

 always  @(posedge pclk)
	wire12245<=wire12254;

 always  @(posedge pclk)
	wire12260<=wire12269;

 always  @(posedge pclk)
	wire12275<=wire12284;

 always  @(posedge pclk)
	ppeaki_13_13_<=wire12314;

 always  @(posedge pclk)
	ppeaki_2_2_<=wire12329;

 always  @(posedge pclk)
	wire12335<=wire12344;

 always  @(posedge pclk)
	wire12350<=wire12359;

 always  @(posedge pclk)
	wire12365<=wire12374;

 always  @(posedge pclk)
	wire12380<=wire12389;

 always  @(posedge pclk)
	wire12395<=wire12404;

 always  @(posedge pclk)
	wire12410<=wire12419;

 always  @(posedge pclk)
	wire12425<=wire12434;

 always  @(posedge pclk)
	wire12440<=wire12449;

 always  @(posedge pclk)
	wire12455<=wire12464;

 always  @(posedge pclk)
	wire12470<=wire12479;

 always  @(posedge pclk)
	wire12485<=wire12494;

 always  @(posedge pclk)
	ppeaki_12_12_<=wire12524;

 always  @(posedge pclk)
	ppeaki_3_3_<=wire12539;

 always  @(posedge pclk)
	wire12545<=wire12554;

 always  @(posedge pclk)
	wire12560<=wire12569;

 always  @(posedge pclk)
	wire12575<=wire12584;

 always  @(posedge pclk)
	wire12590<=wire12599;

 always  @(posedge pclk)
	wire12605<=wire12614;

 always  @(posedge pclk)
	wire12620<=wire12629;

 always  @(posedge pclk)
	wire12635<=wire12644;

 always  @(posedge pclk)
	wire12650<=wire12659;

 always  @(posedge pclk)
	wire12665<=wire12674;

 always  @(posedge pclk)
	wire12680<=wire12689;

 always  @(posedge pclk)
	wire12695<=wire12704;

 always  @(posedge pclk)
	ppeaki_11_11_<=wire12749;

 always  @(posedge pclk)
	ppeaki_0_0_<=wire12764;

 always  @(posedge pclk)
	wire12770<=wire12779;

 always  @(posedge pclk)
	wire12800<=wire12809;

 always  @(posedge pclk)
	wire12815<=wire12824;

 always  @(posedge pclk)
	wire12830<=wire12839;

 always  @(posedge pclk)
	wire12845<=wire12854;

 always  @(posedge pclk)
	wire12860<=wire12869;

 always  @(posedge pclk)
	wire12875<=wire12884;

 always  @(posedge pclk)
	wire12890<=wire12899;

 always  @(posedge pclk)
	wire12905<=wire12914;

 always  @(posedge pclk)
	wire12920<=wire12929;

 always  @(posedge pclk)
	wire12935<=wire12944;

 always  @(posedge pclk)
	ppeaki_10_10_<=wire12989;

 always  @(posedge pclk)
	ppeaki_1_1_<=wire13004;

 always  @(posedge pclk)
	wire13010<=wire13019;

 always  @(posedge pclk)
	wire13025<=wire13034;

 always  @(posedge pclk)
	wire13040<=wire13049;

 always  @(posedge pclk)
	wire13055<=wire13064;

 always  @(posedge pclk)
	wire13070<=wire13079;

 always  @(posedge pclk)
	wire13085<=wire13094;

 always  @(posedge pclk)
	wire13100<=wire13109;

 always  @(posedge pclk)
	wire13115<=wire13124;

 always  @(posedge pclk)
	wire13130<=wire13139;

 always  @(posedge pclk)
	wire13160<=wire13169;

 always  @(posedge pclk)
	wire13175<=wire13184;

 always  @(posedge pclk)
	ppeakb_4_4_<=wire13199;

 always  @(posedge pclk)
	ppeaka_9_9_<=wire13214;

 always  @(posedge pclk)
	wire13220<=wire13229;

 always  @(posedge pclk)
	wire13235<=wire13244;

 always  @(posedge pclk)
	wire13250<=wire13259;

 always  @(posedge pclk)
	wire13265<=wire13274;

 always  @(posedge pclk)
	wire13280<=wire13289;

 always  @(posedge pclk)
	wire13295<=wire13304;

 always  @(posedge pclk)
	wire13310<=wire13319;

 always  @(posedge pclk)
	wire13325<=wire13334;

 always  @(posedge pclk)
	wire13340<=wire13349;

 always  @(posedge pclk)
	wire13355<=wire13364;

 always  @(posedge pclk)
	wire13370<=wire13379;

 always  @(posedge pclk)
	wire13385<=wire13394;

 always  @(posedge pclk)
	wire13400<=wire13409;

 always  @(posedge pclk)
	wire13415<=wire13424;

 always  @(posedge pclk)
	wire13430<=wire13439;

 always  @(posedge pclk)
	wire13445<=wire13454;

 always  @(posedge pclk)
	wire13460<=wire13469;

 always  @(posedge pclk)
	wire13475<=wire13484;

 always  @(posedge pclk)
	wire13490<=wire13499;

 always  @(posedge pclk)
	wire13505<=wire13514;

 always  @(posedge pclk)
	ppeakb_5_5_<=wire13544;

 always  @(posedge pclk)
	wire13550<=wire13559;

 always  @(posedge pclk)
	ppeakp_6_6_<=wire13574;

 always  @(posedge pclk)
	wire13580<=wire13589;

 always  @(posedge pclk)
	wire13595<=wire13604;

 always  @(posedge pclk)
	wire13610<=wire13619;

 always  @(posedge pclk)
	wire13625<=wire13634;

 always  @(posedge pclk)
	wire13640<=wire13649;

 always  @(posedge pclk)
	wire13655<=wire13664;

 always  @(posedge pclk)
	wire13670<=wire13679;

 always  @(posedge pclk)
	wire13685<=wire13694;

 always  @(posedge pclk)
	wire13700<=wire13709;

 always  @(posedge pclk)
	wire13715<=wire13724;

 always  @(posedge pclk)
	wire13730<=wire13739;

 always  @(posedge pclk)
	wire13745<=wire13754;

 always  @(posedge pclk)
	wire13775<=wire13784;

 always  @(posedge pclk)
	wire13790<=wire13799;

 always  @(posedge pclk)
	wire13805<=wire13814;

 always  @(posedge pclk)
	wire13820<=wire13829;

 always  @(posedge pclk)
	wire13835<=wire13844;

 always  @(posedge pclk)
	wire13850<=wire13859;

 always  @(posedge pclk)
	wire13865<=wire13874;

 always  @(posedge pclk)
	wire13880<=wire13889;

 always  @(posedge pclk)
	wire13895<=wire13904;

 always  @(posedge pclk)
	ppeaka_11_11_<=wire13919;

 always  @(posedge pclk)
	ppeaka_0_0_<=wire13934;

 always  @(posedge pclk)
	ppeakp_5_5_<=wire13949;

 always  @(posedge pclk)
	wire13955<=wire13964;

 always  @(posedge pclk)
	wire13970<=wire13979;

 always  @(posedge pclk)
	wire13985<=wire13994;

 always  @(posedge pclk)
	wire14000<=wire14009;

 always  @(posedge pclk)
	wire14015<=wire14024;

 always  @(posedge pclk)
	wire14030<=wire14039;

 always  @(posedge pclk)
	wire14045<=wire14054;

 always  @(posedge pclk)
	wire14060<=wire14069;

 always  @(posedge pclk)
	wire14075<=wire14084;

 always  @(posedge pclk)
	wire14090<=wire14099;

 always  @(posedge pclk)
	wire14105<=wire14114;

 always  @(posedge pclk)
	wire14120<=wire14129;

 always  @(posedge pclk)
	wire14135<=wire14144;

 always  @(posedge pclk)
	wire14150<=wire14159;

 always  @(posedge pclk)
	wire14165<=wire14174;

 always  @(posedge pclk)
	wire14180<=wire14189;

 always  @(posedge pclk)
	wire14210<=wire14219;

 always  @(posedge pclk)
	wire14225<=wire14234;

 always  @(posedge pclk)
	wire14240<=wire14249;

 always  @(posedge pclk)
	wire14255<=wire14264;

 always  @(posedge pclk)
	wire14270<=wire14279;

 always  @(posedge pclk)
	wire14285<=wire14294;

 always  @(posedge pclk)
	ppeakb_3_3_<=wire14309;

 always  @(posedge pclk)
	ppeaka_10_10_<=wire14324;

 always  @(posedge pclk)
	ppeaka_1_1_<=wire14339;

 always  @(posedge pclk)
	ppeakp_4_4_<=wire14354;

 always  @(posedge pclk)
	wire14360<=wire14369;

 always  @(posedge pclk)
	wire14375<=wire14384;

 always  @(posedge pclk)
	wire14390<=wire14399;

 always  @(posedge pclk)
	wire14405<=wire14414;

 always  @(posedge pclk)
	wire14420<=wire14429;

 always  @(posedge pclk)
	wire14435<=wire14444;

 always  @(posedge pclk)
	wire14450<=wire14459;

 always  @(posedge pclk)
	wire14465<=wire14474;

 always  @(posedge pclk)
	wire14480<=wire14489;

 always  @(posedge pclk)
	wire14495<=wire14504;

 always  @(posedge pclk)
	wire14510<=wire14519;

 always  @(posedge pclk)
	wire14525<=wire14534;

 always  @(posedge pclk)
	wire14540<=wire14549;

 always  @(posedge pclk)
	wire14555<=wire14564;

 always  @(posedge pclk)
	wire14570<=wire14579;

 always  @(posedge pclk)
	wire14585<=wire14594;

 always  @(posedge pclk)
	wire14600<=wire14609;

 always  @(posedge pclk)
	wire14615<=wire14624;

 always  @(posedge pclk)
	wire14630<=wire14639;

 always  @(posedge pclk)
	wire14660<=wire14669;

 always  @(posedge pclk)
	wire14675<=wire14684;

 always  @(posedge pclk)
	wire14690<=wire14699;

 always  @(posedge pclk)
	wire14705<=wire14714;

 always  @(posedge pclk)
	ppeakb_8_8_<=wire14729;

 always  @(posedge pclk)
	ppeaka_13_13_<=wire14744;

 always  @(posedge pclk)
	ppeaka_2_2_<=wire14759;

 always  @(posedge pclk)
	wire14765<=wire14774;

 always  @(posedge pclk)
	ppeaks_9_9_<=wire14789;

 always  @(posedge pclk)
	ppeakp_14_14_<=wire14804;

 always  @(posedge pclk)
	wire14810<=wire14819;

 always  @(posedge pclk)
	wire14825<=wire14834;

 always  @(posedge pclk)
	wire14840<=wire14849;

 always  @(posedge pclk)
	wire14855<=wire14864;

 always  @(posedge pclk)
	wire14870<=wire14879;

 always  @(posedge pclk)
	wire14885<=wire14894;

 always  @(posedge pclk)
	wire14900<=wire14909;

 always  @(posedge pclk)
	wire14915<=wire14924;

 always  @(posedge pclk)
	wire14930<=wire14939;

 always  @(posedge pclk)
	wire14960<=wire14969;

 always  @(posedge pclk)
	wire14975<=wire14984;

 always  @(posedge pclk)
	wire14990<=wire14999;

 always  @(posedge pclk)
	wire15005<=wire15014;

 always  @(posedge pclk)
	wire15020<=wire15029;

 always  @(posedge pclk)
	wire15035<=wire15044;

 always  @(posedge pclk)
	wire15050<=wire15059;

 always  @(posedge pclk)
	wire15065<=wire15074;

 always  @(posedge pclk)
	wire15080<=wire15089;

 always  @(posedge pclk)
	ppeakb_9_9_<=wire15104;

 always  @(posedge pclk)
	ppeaka_12_12_<=wire15119;

 always  @(posedge pclk)
	ppeaka_3_3_<=wire15134;

 always  @(posedge pclk)
	wire15140<=wire15149;

 always  @(posedge pclk)
	ppeaks_8_8_<=wire15164;

 always  @(posedge pclk)
	ppeakp_15_15_<=wire15179;

 always  @(posedge pclk)
	wire15185<=wire15194;

 always  @(posedge pclk)
	wire15200<=wire15209;

 always  @(posedge pclk)
	wire15215<=wire15224;

 always  @(posedge pclk)
	wire15230<=wire15239;

 always  @(posedge pclk)
	wire15245<=wire15254;

 always  @(posedge pclk)
	wire15260<=wire15269;

 always  @(posedge pclk)
	wire15275<=wire15284;

 always  @(posedge pclk)
	wire15290<=wire15299;

 always  @(posedge pclk)
	wire15305<=wire15314;

 always  @(posedge pclk)
	wire15320<=wire15329;

 always  @(posedge pclk)
	wire15335<=wire15344;

 always  @(posedge pclk)
	wire15350<=wire15359;

 always  @(posedge pclk)
	wire15365<=wire15374;

 always  @(posedge pclk)
	wire15380<=wire15389;

 always  @(posedge pclk)
	wire15395<=wire15404;

 always  @(posedge pclk)
	wire15410<=wire15419;

 always  @(posedge pclk)
	wire15425<=wire15434;

 always  @(posedge pclk)
	wire15440<=wire15449;

 always  @(posedge pclk)
	ppeakb_6_6_<=wire15464;

 always  @(posedge pclk)
	ppeaka_15_15_<=wire15479;

 always  @(posedge pclk)
	ppeaka_4_4_<=wire15494;

 always  @(posedge pclk)
	wire15500<=wire15509;

 always  @(posedge pclk)
	wire15515<=wire15524;

 always  @(posedge pclk)
	ppeaks_0_0_<=wire15539;

 always  @(posedge pclk)
	wire15545<=wire15554;

 always  @(posedge pclk)
	wire15560<=wire15569;

 always  @(posedge pclk)
	wire15575<=wire15584;

 always  @(posedge pclk)
	wire15590<=wire15599;

 always  @(posedge pclk)
	wire15605<=wire15614;

 always  @(posedge pclk)
	wire15620<=wire15629;

 always  @(posedge pclk)
	wire15635<=wire15644;

 always  @(posedge pclk)
	wire15650<=wire15659;

 always  @(posedge pclk)
	wire15665<=wire15674;

 always  @(posedge pclk)
	wire15680<=wire15689;

 always  @(posedge pclk)
	wire15695<=wire15704;

 always  @(posedge pclk)
	wire15710<=wire15719;

 always  @(posedge pclk)
	wire15725<=wire15734;

 always  @(posedge pclk)
	wire15755<=wire15764;

 always  @(posedge pclk)
	wire15770<=wire15779;

 always  @(posedge pclk)
	wire15785<=wire15794;

 always  @(posedge pclk)
	ppeakb_7_7_<=wire15809;

 always  @(posedge pclk)
	ppeaka_14_14_<=wire15824;

 always  @(posedge pclk)
	ppeaka_5_5_<=wire15839;

 always  @(posedge pclk)
	wire15845<=wire15854;

 always  @(posedge pclk)
	wire15860<=wire15869;

 always  @(posedge pclk)
	ppeaks_10_10_<=wire15884;

 always  @(posedge pclk)
	wire15890<=wire15899;

 always  @(posedge pclk)
	wire15905<=wire15914;

 always  @(posedge pclk)
	wire15920<=wire15929;

 always  @(posedge pclk)
	wire15935<=wire15944;

 always  @(posedge pclk)
	wire15950<=wire15959;

 always  @(posedge pclk)
	wire15965<=wire15974;

 always  @(posedge pclk)
	wire15980<=wire15989;

 always  @(posedge pclk)
	wire15995<=wire16004;

 always  @(posedge pclk)
	wire16010<=wire16019;

 always  @(posedge pclk)
	wire16025<=wire16034;

 always  @(posedge pclk)
	wire16040<=wire16049;

 always  @(posedge pclk)
	wire16055<=wire16064;

 always  @(posedge pclk)
	wire16070<=wire16079;

 always  @(posedge pclk)
	wire16085<=wire16094;

 always  @(posedge pclk)
	wire16100<=wire16109;

 always  @(posedge pclk)
	paddress_8_8_<=wire16904;

 always  @(posedge pclk)
	wire16907<=wire16917;

 always  @(posedge pclk)
	wire16920<=wire16928;

 always  @(posedge pclk)
	wire16933<=wire16941;

 always  @(posedge pclk)
	paddress_9_9_<=wire16956;

 always  @(posedge pclk)
	wire16959<=wire16969;

 always  @(posedge pclk)
	wire16972<=wire16980;

 always  @(posedge pclk)
	wire16985<=wire16993;

 always  @(posedge pclk)
	wire16998<=wire17008;

 always  @(posedge pclk)
	wire17011<=wire17021;

 always  @(posedge pclk)
	wire17024<=wire17032;

 always  @(posedge pclk)
	wire17037<=wire17045;

 always  @(posedge pclk)
	wire17050<=wire17058;

 always  @(posedge pclk)
	wire17063<=wire17073;

 always  @(posedge pclk)
	wire17076<=wire17086;

 always  @(posedge pclk)
	wire17089<=wire17097;

 always  @(posedge pclk)
	wire17102<=wire17110;

 always  @(posedge pclk)
	wire17115<=wire17123;

 always  @(posedge pclk)
	wire17128<=wire17138;

 always  @(posedge pclk)
	wire17141<=wire17151;

 always  @(posedge pclk)
	wire17154<=wire17162;

 always  @(posedge pclk)
	wire17167<=wire17175;

 always  @(posedge pclk)
	wire17180<=wire17188;

 always  @(posedge pclk)
	wire17193<=wire17203;

 always  @(posedge pclk)
	wire17206<=wire17214;

 always  @(posedge pclk)
	wire17219<=wire17227;

 always  @(posedge pclk)
	wire17232<=wire17240;

 always  @(posedge pclk)
	wire17245<=wire17253;

 always  @(posedge pclk)
	wire17258<=wire17268;

 always  @(posedge pclk)
	wire17271<=wire17279;

 always  @(posedge pclk)
	wire17284<=wire17292;

 always  @(posedge pclk)
	wire17297<=wire17305;

 always  @(posedge pclk)
	wire17310<=wire17318;

 always  @(posedge pclk)
	wire17323<=wire17333;

 always  @(posedge pclk)
	wire17336<=wire17346;

 always  @(posedge pclk)
	wire17349<=wire17357;

 always  @(posedge pclk)
	wire17362<=wire17370;

 always  @(posedge pclk)
	wire17375<=wire17383;

 always  @(posedge pclk)
	wire17388<=wire17396;

 always  @(posedge pclk)
	paddress_11_11_<=wire17411;

 always  @(posedge pclk)
	wire17414<=wire17422;

 always  @(posedge pclk)
	wire17427<=wire17435;

 always  @(posedge pclk)
	wire17453<=wire17461;

 always  @(posedge pclk)
	paddress_10_10_<=wire17476;

 always  @(posedge pclk)
	wire17479<=wire17489;

 always  @(posedge pclk)
	wire17492<=wire17502;

 always  @(posedge pclk)
	wire17505<=wire17513;

 always  @(posedge pclk)
	wire17518<=wire17526;

 always  @(posedge pclk)
	wire17531<=wire17539;

 always  @(posedge pclk)
	wire17544<=wire17554;

 always  @(posedge pclk)
	paddress_13_13_<=wire17567;

 always  @(posedge pclk)
	wire17570<=wire17578;

 always  @(posedge pclk)
	wire17583<=wire17591;

 always  @(posedge pclk)
	wire17596<=wire17604;

 always  @(posedge pclk)
	wire17609<=wire17619;

 always  @(posedge pclk)
	paddress_12_12_<=wire17632;

 always  @(posedge pclk)
	wire17635<=wire17643;

 always  @(posedge pclk)
	wire17648<=wire17656;

 always  @(posedge pclk)
	wire17661<=wire17669;

 always  @(posedge pclk)
	wire17674<=wire17684;

 always  @(posedge pclk)
	paddress_15_15_<=wire17697;

 always  @(posedge pclk)
	wire17700<=wire17708;

 always  @(posedge pclk)
	wire17713<=wire17723;

 always  @(posedge pclk)
	paddress_14_14_<=wire17736;

 always  @(posedge pclk)
	wire17739<=wire17747;

 always  @(posedge pclk)
	wire17752<=wire17760;

 always  @(posedge pclk)
	wire17765<=wire17775;

 always  @(posedge pclk)
	wire17778<=wire17788;

 always  @(posedge pclk)
	wire17791<=wire17799;

 always  @(posedge pclk)
	wire17804<=wire17812;

 always  @(posedge pclk)
	wire17817<=wire17825;

 always  @(posedge pclk)
	pwr_0_0_<=wire17840;

 always  @(posedge pclk)
	wire17843<=wire17851;

 always  @(posedge pclk)
	wire17856<=wire17866;

 always  @(posedge pclk)
	wire17869<=wire17879;

 always  @(posedge pclk)
	wire17882<=wire17892;

 always  @(posedge pclk)
	prd_0_0_<=wire17905;

 always  @(posedge pclk)
	wire17908<=wire17918;

 always  @(posedge pclk)
	wire17921<=wire17931;

 always  @(posedge pclk)
	wire17934<=wire17944;

 always  @(posedge pclk)
	wire17947<=wire17957;

 always  @(posedge pclk)
	wire17960<=wire17970;

 always  @(posedge pclk)
	wire17973<=wire17983;

 always  @(posedge pclk)
	wire17986<=wire17994;

 always  @(posedge pclk)
	wire17999<=wire18007;

 always  @(posedge pclk)
	wire18012<=wire18022;

 always  @(posedge pclk)
	wire18025<=wire18033;

 always  @(posedge pclk)
	wire18038<=wire18048;

 always  @(posedge pclk)
	pdn<=wire18059;

 always  @(posedge pclk)
	wire18064<=wire18072;

 always  @(posedge pclk)
	wire18077<=wire18085;

 always  @(posedge pclk)
	wire18090<=wire18100;

 always  @(posedge pclk)
	wire18103<=wire18111;

 always  @(posedge pclk)
	wire18116<=wire18126;

 always  @(posedge pclk)
	wire18129<=wire18139;

 always  @(posedge pclk)
	wire18142<=wire18150;

 always  @(posedge pclk)
	wire18155<=wire18165;

 always  @(posedge pclk)
	wire18168<=wire18176;

 always  @(posedge pclk)
	wire18181<=wire18191;

 always  @(posedge pclk)
	wire18194<=wire18204;

 always  @(posedge pclk)
	wire18207<=wire18215;

 always  @(posedge pclk)
	wire18220<=wire18228;

 always  @(posedge pclk)
	wire18233<=wire18243;

 always  @(posedge pclk)
	wire18246<=wire18254;

 always  @(posedge pclk)
	paddress_0_0_<=wire18269;

 always  @(posedge pclk)
	piack_0_0_<=wire18282;

 always  @(posedge pclk)
	wire18285<=wire18293;

 always  @(posedge pclk)
	wire18298<=wire18306;

 always  @(posedge pclk)
	wire18311<=wire18319;

 always  @(posedge pclk)
	paddress_1_1_<=wire18334;

 always  @(posedge pclk)
	wire18337<=wire18347;

 always  @(posedge pclk)
	wire18350<=wire18360;

 always  @(posedge pclk)
	wire18363<=wire18371;

 always  @(posedge pclk)
	wire18376<=wire18384;

 always  @(posedge pclk)
	wire18389<=wire18397;

 always  @(posedge pclk)
	paddress_2_2_<=wire18412;

 always  @(posedge pclk)
	wire18415<=wire18423;

 always  @(posedge pclk)
	wire18428<=wire18436;

 always  @(posedge pclk)
	wire18441<=wire18449;

 always  @(posedge pclk)
	paddress_3_3_<=wire18464;

 always  @(posedge pclk)
	wire18467<=wire18475;

 always  @(posedge pclk)
	wire18480<=wire18488;

 always  @(posedge pclk)
	wire18493<=wire18501;

 always  @(posedge pclk)
	wire18506<=wire18514;

 always  @(posedge pclk)
	paddress_4_4_<=wire18529;

 always  @(posedge pclk)
	paddress_5_5_<=wire18542;

 always  @(posedge pclk)
	wire18545<=wire18555;

 always  @(posedge pclk)
	paddress_6_6_<=wire18568;

 always  @(posedge pclk)
	wire18571<=wire18581;

 always  @(posedge pclk)
	wire18584<=wire18594;

 always  @(posedge pclk)
	wire18597<=wire18605;

 always  @(posedge pclk)
	wire18610<=wire18618;

 always  @(posedge pclk)
	paddress_7_7_<=wire18633;

 always  @(posedge pclk)
	wire18636<=wire18644;

 assign pdata_8_8_ = ( wire16959  &  wire17882 ) | ( tin_pdata_8_8_  &  (~ wire17882) ) ;
 assign pdata_0_0_ = ( tin_pdata_0_0_  &  (~ wire17479) ) | ( wire17479  &  wire18337 ) ;
 assign pdata_7_7_ = ( wire16907  &  wire17869 ) | ( tin_pdata_7_7_  &  (~ wire17869) ) ;
 assign pdata_2_2_ = ( wire17323  &  wire18181 ) | ( tin_pdata_2_2_  &  (~ wire18181) ) ;
 assign pdata_9_9_ = ( wire17765  &  wire18571 ) | ( tin_pdata_9_9_  &  (~ wire18571) ) ;
 assign pdata_1_1_ = ( wire17258  &  wire18116 ) | ( tin_pdata_1_1_  &  (~ wire18116) ) ;
 assign pdata_4_4_ = ( wire17193  &  wire18038 ) | ( tin_pdata_4_4_  &  (~ wire18038) ) ;
 assign pdata_10_10_ = ( tin_pdata_10_10_  &  (~ wire17011) ) | ( wire17011  &  wire17921 ) ;
 assign pdata_3_3_ = ( wire17128  &  wire17960 ) | ( tin_pdata_3_3_  &  (~ wire17960) ) ;
 assign pdata_6_6_ = ( wire17063  &  wire17934 ) | ( tin_pdata_6_6_  &  (~ wire17934) ) ;
 assign pdata_15_15_ = ( wire17076  &  wire17947 ) | ( tin_pdata_15_15_  &  (~ wire17947) ) ;
 assign pdata_11_11_ = ( tin_pdata_11_11_  &  (~ wire17336) ) | ( wire17336  &  wire18194 ) ;
 assign pdata_14_14_ = ( wire17778  &  wire18584 ) | ( tin_pdata_14_14_  &  (~ wire18584) ) ;
 assign pdata_12_12_ = ( tin_pdata_12_12_  &  (~ wire17141) ) | ( wire17141  &  wire17973 ) ;
 assign pdata_5_5_ = ( wire16998  &  wire17908 ) | ( tin_pdata_5_5_  &  (~ wire17908) ) ;
 assign pdata_13_13_ = ( wire17492  &  wire18350 ) | ( tin_pdata_13_13_  &  (~ wire18350) ) ;
 assign wire4244 = ( wire5582 ) | ( pdata_2_2_  &  wire4305 ) ;
 assign wire4259 = ( wire17615 ) | ( wire17616 ) | ( wire17621 ) ;
 assign wire4274 = ( wire17626 ) | ( wire17627 ) | ( wire17631 ) ;
 assign wire4289 = ( wire17641 ) | ( wire17642 ) | ( wire17647 ) ;
 assign wire4304 = ( wire5455 ) | ( wire5456 ) | ( wire17652 ) ;
 assign wire4319 = ( wire5451 ) | ( wire5452 ) | ( wire17654 ) ;
 assign wire4334 = ( wire17672 ) | ( wire17673 ) | ( wire17678 ) ;
 assign wire4349 = ( wire5407 ) | ( wire5410 ) | ( wire5411 ) | ( wire17705 ) ;
 assign wire4364 = ( wire5403 ) | ( pdata_0_0_  &  wire4352 ) ;
 assign wire4379 = ( wire5398 ) | ( pdata_11_11_  &  wire4352 ) ;
 assign wire4394 = ( (~ preset)  &  pdata_6_6_  &  nrq10_4 ) | ( (~ preset)  &  wire4385  &  (~ nrq10_4) ) ;
 assign wire4409 = ( wire5389 ) | ( pdata_1_1_  &  wire4353 ) ;
 assign wire4424 = ( wire5385 ) | ( pdata_12_12_  &  wire4353 ) ;
 assign wire4439 = ( (~ preset)  &  pdata_7_7_  &  nrq14_3 ) | ( (~ preset)  &  wire4430  &  (~ nrq14_3) ) ;
 assign wire4454 = ( (~ preset)  &  pdata_2_2_  &  nrq14_3 ) | ( (~ preset)  &  wire4445  &  (~ nrq14_3) ) ;
 assign wire4469 = ( (~ preset)  &  pdata_13_13_  &  nrq14_3 ) | ( (~ preset)  &  wire4460  &  (~ nrq14_3) ) ;
 assign wire4484 = ( wire5368 ) | ( pdata_8_8_  &  wire4354 ) ;
 assign wire4499 = ( wire5363 ) | ( pdata_3_3_  &  wire18384 ) ;
 assign wire4514 = ( wire5358 ) | ( pdata_14_14_  &  wire18384 ) ;
 assign wire4529 = ( wire5353 ) | ( wire5355 ) ;
 assign wire4544 = ( wire5349 ) | ( wire5350 ) ;
 assign wire4559 = ( wire5344 ) | ( wire5346 ) ;
 assign wire4574 = ( (~ preset)  &  pdata_5_5_  &  nrq23_3 ) | ( (~ preset)  &  wire4565  &  (~ nrq23_3) ) ;
 assign wire4589 = ( (~ preset)  &  pdata_0_0_  &  nrq23_3 ) | ( (~ preset)  &  wire4580  &  (~ nrq23_3) ) ;
 assign wire4604 = ( (~ preset)  &  pdata_11_11_  &  nrq23_3 ) | ( (~ preset)  &  wire4595  &  (~ nrq23_3) ) ;
 assign wire4619 = ( wire5334 ) | ( pdata_6_6_  &  wire4375 ) ;
 assign wire4634 = ( wire17461  &  wire19360 ) | ( wire4625  &  wire4340 ) ;
 assign wire4649 = ( wire4640  &  wire4340 ) | ( wire17461  &  wire19390 ) ;
 assign wire4664 = ( wire5143 ) | ( wire5145 ) ;
 assign wire4679 = ( wire5139 ) | ( wire4670  &  wire4253 ) ;
 assign wire4709 = ( wire5132 ) | ( wire5133 ) ;
 assign wire4724 = ( wire5126 ) | ( wire4715  &  wire4317 ) ;
 assign wire4739 = ( wire4730  &  wire4317 ) | ( wire4381  &  wire19368 ) ;
 assign wire4754 = ( wire5073 ) | ( wire18501  &  wire19359 ) ;
 assign wire4769 = ( wire5068 ) | ( wire4760  &  wire4252 ) ;
 assign wire4784 = ( wire5063 ) | ( wire4775  &  wire4252 ) ;
 assign wire4799 = ( wire5057 ) | ( wire5058 ) ;
 assign wire4814 = ( wire4805  &  wire4277 ) | ( wire19360  &  wire4278 ) ;
 assign wire4829 = ( wire4820  &  wire4277 ) | ( wire19390  &  wire4278 ) ;
 assign wire4844 = ( (~ preset)  &  wire19088  &  nrq4_2 ) | ( (~ preset)  &  wire4835  &  (~ nrq4_2) ) ;
 assign wire4859 = ( wire4902 ) | ( wire19092  &  wire4345 ) ;
 assign wire4874 = ( wire4865  &  wire4330 ) | ( wire19103  &  wire4374 ) ;
 assign wire4889 = ( wire4834 ) | ( wire4374  &  wire4388  &  wire4511 ) | ( wire4374  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire4904 = ( wire4828 ) | ( wire19060  &  wire4360 ) ;
 assign wire4919 = ( wire4910  &  wire4331 ) | ( wire19097  &  wire4332 ) ;
 assign wire4934 = ( wire4925  &  wire4277 ) | ( wire4278  &  wire19061 ) ;
 assign wire4949 = ( wire4940  &  wire4277 ) | ( wire4278  &  wire19091 ) ;
 assign wire4964 = ( wire4955  &  wire4336 ) | ( wire19088  &  wire4365 ) ;
 assign wire4979 = ( wire4807 ) | ( pdata_1_1_  &  wire4305 ) ;
 assign wire4994 = ( wire18037 ) | ( wire18039 ) | ( wire18043 ) ;
 assign wire5009 = ( wire18051 ) | ( wire18052 ) | ( wire18056 ) ;
 assign wire5024 = ( wire4773 ) | ( wire4774 ) | ( wire18057 ) ;
 assign wire5039 = ( wire4768 ) | ( wire4770 ) | ( wire18060 ) ;
 assign wire5054 = ( wire18071 ) | ( wire18073 ) | ( wire18078 ) ;
 assign wire5069 = ( wire4742 ) | ( wire4746 ) | ( wire4747 ) | ( wire18080 ) ;
 assign wire5084 = ( wire4741 ) | ( pdata_1_1_  &  wire4352 ) ;
 assign wire5099 = ( wire4738 ) | ( pdata_10_10_  &  wire4352 ) ;
 assign wire5114 = ( wire4736 ) | ( pdata_2_2_  &  wire4353 ) ;
 assign wire5129 = ( wire4734 ) | ( pdata_11_11_  &  wire4353 ) ;
 assign wire5144 = ( (~ preset)  &  pdata_8_8_  &  nrq14_3 ) | ( (~ preset)  &  wire5135  &  (~ nrq14_3) ) ;
 assign wire5159 = ( (~ preset)  &  pdata_1_1_  &  nrq14_3 ) | ( (~ preset)  &  wire5150  &  (~ nrq14_3) ) ;
 assign wire5174 = ( (~ preset)  &  pdata_14_14_  &  nrq14_3 ) | ( (~ preset)  &  wire5165  &  (~ nrq14_3) ) ;
 assign wire5189 = ( wire4725 ) | ( pdata_7_7_  &  wire4354 ) ;
 assign wire5204 = ( wire4719 ) | ( pdata_4_4_  &  wire18384 ) ;
 assign wire5219 = ( wire4717 ) | ( pdata_13_13_  &  wire18384 ) ;
 assign wire5234 = ( wire4714 ) | ( wire4716 ) ;
 assign wire5249 = ( wire4712 ) | ( wire4713 ) ;
 assign wire5264 = ( wire4710 ) | ( wire4711 ) ;
 assign wire5279 = ( (~ preset)  &  pdata_4_4_  &  nrq23_3 ) | ( (~ preset)  &  wire5270  &  (~ nrq23_3) ) ;
 assign wire5294 = ( (~ preset)  &  pdata_1_1_  &  nrq23_3 ) | ( (~ preset)  &  wire5285  &  (~ nrq23_3) ) ;
 assign wire5309 = ( (~ preset)  &  pdata_10_10_  &  nrq23_3 ) | ( (~ preset)  &  wire5300  &  (~ nrq23_3) ) ;
 assign wire5324 = ( wire4702 ) | ( pdata_7_7_  &  wire4375 ) ;
 assign wire5339 = ( wire4698 ) | ( wire17461  &  (~ n_n2471)  &  n_n2487 ) | ( wire17461  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire5354 = ( wire4697 ) | ( wire5345  &  wire4340 ) ;
 assign wire5369 = ( wire4694 ) | ( wire19390  &  wire4308 ) ;
 assign wire5384 = ( wire4693 ) | ( wire5375  &  wire4253 ) ;
 assign wire5399 = ( wire4690 ) | ( wire4306  &  (~ n_n2471)  &  n_n2487 ) | ( wire4306  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire5414 = ( wire4688 ) | ( wire4306  &  wire19359 ) ;
 assign wire5429 = ( wire4686 ) | ( wire5420  &  wire4317 ) ;
 assign wire5444 = ( wire5435  &  wire4317 ) | ( wire4381  &  wire19367 ) ;
 assign wire5459 = ( wire4682 ) | ( wire4683 ) ;
 assign wire5474 = ( wire4680 ) | ( wire17305  &  wire19359 ) ;
 assign wire5489 = ( wire5480  &  wire4252 ) | ( wire4245  &  wire19367 ) ;
 assign wire5504 = ( wire4673 ) | ( wire4377  &  wire19387 ) ;
 assign wire5519 = ( wire4669 ) | ( wire5510  &  wire4277 ) ;
 assign wire5534 = ( wire4667 ) | ( wire5525  &  wire4277 ) ;
 assign wire5549 = ( (~ preset)  &  wire19070  &  nrq4_2 ) | ( (~ preset)  &  wire5540  &  (~ nrq4_2) ) ;
 assign wire5564 = ( wire4657 ) | ( wire4345  &  wire19096 ) ;
 assign wire5579 = ( wire5570  &  wire4330 ) | ( wire4374  &  wire19097 ) ;
 assign wire5609 = ( wire4648 ) | ( wire4360  &  wire19072 ) ;
 assign wire5624 = ( wire5615  &  wire4331 ) | ( wire19103  &  wire4332 ) ;
 assign wire5639 = ( wire4643 ) | ( wire17240  &  wire19072 ) ;
 assign wire5654 = ( wire5645  &  wire4277 ) | ( wire4278  &  wire19087 ) ;
 assign wire5669 = ( wire5660  &  wire4336 ) | ( wire4365  &  wire19082 ) ;
 assign wire5684 = ( wire4629 ) | ( pdata_0_0_  &  wire4305 ) ;
 assign wire5699 = ( wire18114 ) | ( wire18115 ) | ( wire18120 ) ;
 assign wire5714 = ( wire18128 ) | ( wire18130 ) | ( wire18134 ) ;
 assign wire5729 = ( wire4596 ) | ( wire4597 ) | ( wire18135 ) ;
 assign wire5744 = ( wire18147 ) | ( wire18148 ) | ( wire18153 ) ;
 assign wire5759 = ( wire18163 ) | ( wire18164 ) | ( wire18170 ) ;
 assign wire5774 = ( wire4551 ) | ( wire4554 ) | ( wire4555 ) | ( wire18172 ) ;
 assign wire5789 = ( wire4549 ) | ( pdata_2_2_  &  wire4352 ) ;
 assign wire5804 = ( (~ preset)  &  pdata_4_4_  &  nrq10_4 ) | ( (~ preset)  &  wire5795  &  (~ nrq10_4) ) ;
 assign wire5819 = ( (~ preset)  &  pdata_8_8_  &  nrq10_4 ) | ( (~ preset)  &  wire5810  &  (~ nrq10_4) ) ;
 assign wire5834 = ( (~ preset)  &  pdata_9_9_  &  nrq14_3 ) | ( (~ preset)  &  wire5825  &  (~ nrq14_3) ) ;
 assign wire5849 = ( (~ preset)  &  pdata_4_4_  &  nrq14_3 ) | ( (~ preset)  &  wire5840  &  (~ nrq14_3) ) ;
 assign wire5864 = ( (~ preset)  &  pdata_11_11_  &  nrq14_3 ) | ( (~ preset)  &  wire5855  &  (~ nrq14_3) ) ;
 assign wire5879 = ( wire4536 ) | ( pdata_6_6_  &  wire4354 ) ;
 assign wire5894 = ( wire4532 ) | ( pdata_5_5_  &  wire18384 ) ;
 assign wire5909 = ( wire4530 ) | ( wire4531 ) ;
 assign wire5924 = ( wire4527 ) | ( wire4528 ) ;
 assign wire5939 = ( wire4525 ) | ( wire4526 ) ;
 assign wire5954 = ( wire4523 ) | ( wire4524 ) ;
 assign wire5969 = ( (~ preset)  &  pdata_7_7_  &  nrq23_3 ) | ( (~ preset)  &  wire5960  &  (~ nrq23_3) ) ;
 assign wire5984 = ( (~ preset)  &  pdata_14_14_  &  nrq23_3 ) | ( (~ preset)  &  wire5975  &  (~ nrq23_3) ) ;
 assign wire5999 = ( (~ preset)  &  pdata_9_9_  &  nrq23_3 ) | ( (~ preset)  &  wire5990  &  (~ nrq23_3) ) ;
 assign wire6014 = ( wire4506 ) | ( pdata_8_8_  &  wire4375 ) ;
 assign wire6029 = ( wire6020  &  wire4340 ) | ( wire17461  &  wire19396 ) ;
 assign wire6044 = ( wire4497 ) | ( wire6035  &  wire4340 ) ;
 assign wire6059 = ( wire4493 ) | ( wire4494 ) ;
 assign wire6074 = ( wire4492 ) | ( wire6065  &  wire4253 ) ;
 assign wire6089 = ( wire6080  &  wire4253 ) | ( wire4243  &  wire19367 ) ;
 assign wire6104 = ( wire4291 ) | ( wire4406 ) ;
 assign wire6119 = ( wire6110  &  wire4317 ) | ( wire4381  &  wire19387 ) ;
 assign wire6134 = ( wire4263 ) | ( wire18501  &  (~ n_n2471)  &  n_n2487 ) | ( wire18501  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire6149 = ( wire4257 ) | ( wire4262 ) ;
 assign wire6164 = ( wire4250 ) | ( wire4251 ) ;
 assign wire6179 = ( wire4249 ) | ( wire6170  &  wire4252 ) ;
 assign wire6194 = ( wire4246 ) | ( wire4247 ) ;
 assign wire6209 = ( wire6200  &  wire4277 ) | ( wire4278  &  wire19396 ) ;
 assign wire6224 = ( wire6215  &  wire4277 ) | ( wire4278  &  wire19367 ) ;
 assign wire6239 = ( (~ preset)  &  wire19103  &  nrq4_2 ) | ( (~ preset)  &  wire6230  &  (~ nrq4_2) ) ;
 assign wire6254 = ( wire4230 ) | ( wire19070  &  wire4383 ) ;
 assign wire6269 = ( wire4227 ) | ( wire4345  &  wire19061 ) ;
 assign wire6284 = ( wire4218 ) | ( wire4360  &  wire19073 ) ;
 assign wire6299 = ( wire4213 ) | ( wire4360  &  wire19096 ) ;
 assign wire6314 = ( wire6305  &  wire4331 ) | ( wire4332  &  wire19061 ) ;
 assign wire6329 = ( wire4196 ) | ( wire4307  &  wire4388  &  wire4511 ) | ( wire4307  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire6344 = ( wire6335  &  wire4277 ) | ( wire4278  &  wire19068 ) ;
 assign wire6359 = ( wire6350  &  wire4336 ) | ( wire4365  &  wire19072 ) ;
 assign wire6374 = ( wire4188 ) | ( wire4365  &  wire4388  &  wire4511 ) | ( wire4365  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire6389 = ( wire18189 ) | ( wire18190 ) | ( wire18196 ) ;
 assign wire6404 = ( wire18201 ) | ( wire18202 ) | ( wire18208 ) ;
 assign wire6419 = ( wire4160 ) | ( wire4161 ) | ( wire18209 ) ;
 assign wire6434 = ( wire18221 ) | ( wire18222 ) | ( wire18226 ) ;
 assign wire6449 = ( wire18237 ) | ( wire18238 ) | ( wire18242 ) ;
 assign wire6464 = ( wire4121 ) | ( wire4124 ) | ( wire4125 ) | ( wire18245 ) ;
 assign wire6479 = ( wire4120 ) | ( pdata_12_12_  &  wire4352 ) ;
 assign wire6494 = ( (~ preset)  &  pdata_5_5_  &  nrq10_4 ) | ( (~ preset)  &  wire6485  &  (~ nrq10_4) ) ;
 assign wire6509 = ( (~ preset)  &  pdata_7_7_  &  nrq10_4 ) | ( (~ preset)  &  wire6500  &  (~ nrq10_4) ) ;
 assign wire6524 = ( (~ preset)  &  pdata_10_10_  &  nrq14_3 ) | ( (~ preset)  &  wire6515  &  (~ nrq14_3) ) ;
 assign wire6539 = ( (~ preset)  &  pdata_3_3_  &  nrq14_3 ) | ( (~ preset)  &  wire6530  &  (~ nrq14_3) ) ;
 assign wire6554 = ( (~ preset)  &  pdata_12_12_  &  nrq14_3 ) | ( (~ preset)  &  wire6545  &  (~ nrq14_3) ) ;
 assign wire6569 = ( wire4108 ) | ( pdata_5_5_  &  wire4354 ) ;
 assign wire6584 = ( wire4105 ) | ( pdata_6_6_  &  wire18384 ) ;
 assign wire6599 = ( wire4103 ) | ( pdata_15_15_  &  wire18384 ) ;
 assign wire6614 = ( wire4101 ) | ( wire4102 ) ;
 assign wire6629 = ( wire4099 ) | ( wire4100 ) ;
 assign wire6644 = ( (~ preset)  &  pdata_6_6_  &  nrq23_3 ) | ( (~ preset)  &  wire6635  &  (~ nrq23_3) ) ;
 assign wire6659 = ( (~ preset)  &  pdata_15_15_  &  nrq23_3 ) | ( (~ preset)  &  wire6650  &  (~ nrq23_3) ) ;
 assign wire6674 = ( (~ preset)  &  pdata_8_8_  &  nrq23_3 ) | ( (~ preset)  &  wire6665  &  (~ nrq23_3) ) ;
 assign wire6689 = ( wire4092 ) | ( pdata_9_9_  &  wire4375 ) ;
 assign wire6704 = ( wire4090 ) | ( wire6695  &  wire4340 ) ;
 assign wire6719 = ( wire4088 ) | ( wire6710  &  wire4340 ) ;
 assign wire6734 = ( wire4085 ) | ( wire4308  &  wire19367 ) ;
 assign wire6749 = ( wire6740  &  wire4253 ) | ( wire4243  &  wire19387 ) ;
 assign wire6764 = ( wire6755  &  wire4253 ) | ( wire4243  &  wire19368 ) ;
 assign wire6779 = ( wire4079 ) | ( wire4080 ) ;
 assign wire6794 = ( wire4077 ) | ( wire6785  &  wire4317 ) ;
 assign wire6824 = ( wire4075 ) | ( wire4076 ) ;
 assign wire6839 = ( wire4073 ) | ( wire4074 ) ;
 assign wire6854 = ( wire6845  &  wire4252 ) | ( wire4245  &  wire19396 ) ;
 assign wire6869 = ( wire6860  &  wire4252 ) | ( wire4245  &  wire19390 ) ;
 assign wire6884 = ( wire4067 ) | ( wire6875  &  wire4277 ) ;
 assign wire6899 = ( wire4065 ) | ( wire6890  &  wire4277 ) ;
 assign wire6914 = ( (~ preset)  &  wire19082  &  nrq4_2 ) | ( (~ preset)  &  wire6905  &  (~ nrq4_2) ) ;
 assign wire6929 = ( wire4062 ) | ( wire19072  &  wire4383 ) ;
 assign wire6944 = ( wire4060 ) | ( wire4345  &  wire19073 ) ;
 assign wire6959 = ( wire4058 ) | ( wire4360  &  wire19061 ) ;
 assign wire6974 = ( wire4056 ) | ( wire19092  &  wire4360 ) ;
 assign wire6989 = ( wire6980  &  wire4331 ) | ( wire4332  &  wire19065 ) ;
 assign wire7004 = ( wire19082  &  wire4307 ) | ( wire6995  &  wire4325 ) ;
 assign wire7019 = ( wire4047 ) | ( wire4278  &  wire4388  &  wire4511 ) | ( wire4278  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire7034 = ( wire7025  &  wire4336 ) | ( wire4365  &  wire19070 ) ;
 assign wire7064 = ( wire4041 ) | ( wire4042 ) | ( wire18253 ) ;
 assign wire7079 = ( wire18264 ) | ( wire18265 ) | ( wire18270 ) ;
 assign wire7094 = ( wire18279 ) | ( wire18280 ) | ( wire18286 ) ;
 assign wire7109 = ( wire4001 ) | ( wire4004 ) | ( wire4005 ) | ( wire18288 ) ;
 assign wire7124 = ( wire4000 ) | ( pdata_7_7_  &  wire4352 ) ;
 assign wire7139 = ( (~ preset)  &  pdata_2_2_  &  nrq10_4 ) | ( (~ preset)  &  wire7130  &  (~ nrq10_4) ) ;
 assign wire7154 = ( (~ preset)  &  pdata_11_11_  &  nrq14_3 ) | ( (~ preset)  &  wire7145  &  (~ nrq14_3) ) ;
 assign wire7169 = ( (~ preset)  &  pdata_6_6_  &  nrq14_3 ) | ( (~ preset)  &  wire7160  &  (~ nrq14_3) ) ;
 assign wire7184 = ( wire3992 ) | ( pdata_1_1_  &  wire4354 ) ;
 assign wire7199 = ( wire3990 ) | ( pdata_12_12_  &  wire4354 ) ;
 assign wire7214 = ( wire3988 ) | ( pdata_15_15_  &  wire4354 ) ;
 assign wire7229 = ( wire3985 ) | ( pdata_10_10_  &  wire18384 ) ;
 assign wire7244 = ( wire3983 ) | ( wire3984 ) ;
 assign wire7259 = ( wire3981 ) | ( wire3982 ) ;
 assign wire7274 = ( (~ preset)  &  pdata_9_9_  &  nrq23_3 ) | ( (~ preset)  &  wire7265  &  (~ nrq23_3) ) ;
 assign wire7289 = ( (~ preset)  &  pdata_4_4_  &  nrq23_3 ) | ( (~ preset)  &  wire7280  &  (~ nrq23_3) ) ;
 assign wire7304 = ( (~ preset)  &  pdata_15_15_  &  nrq23_3 ) | ( (~ preset)  &  wire7295  &  (~ nrq23_3) ) ;
 assign wire7319 = ( wire3974 ) | ( pdata_2_2_  &  wire4375 ) ;
 assign wire7334 = ( wire3972 ) | ( pdata_13_13_  &  wire4375 ) ;
 assign wire7349 = ( wire3970 ) | ( wire7340  &  wire4340 ) ;
 assign wire7364 = ( wire3967 ) | ( wire4308  &  wire19368 ) ;
 assign wire7379 = ( wire7370  &  wire4253 ) | ( wire4243  &  wire19359 ) ;
 assign wire7394 = ( wire3963 ) | ( wire4306  &  wire19396 ) ;
 assign wire7409 = ( wire3961 ) | ( wire4306  &  wire19367 ) ;
 assign wire7424 = ( wire3960 ) | ( wire4381  &  (~ n_n2471)  &  n_n2487 ) | ( wire4381  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire7439 = ( wire3957 ) | ( wire7430  &  wire4317 ) ;
 assign wire7454 = ( wire3955 ) | ( wire3956 ) ;
 assign wire7469 = ( wire3953 ) | ( wire17305  &  wire19390 ) ;
 assign wire7484 = ( wire7475  &  wire4252 ) | ( wire4245  &  wire19387 ) ;
 assign wire7499 = ( wire3950 ) | ( wire4377  &  (~ n_n2471)  &  n_n2487 ) | ( wire4377  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire7514 = ( wire3947 ) | ( wire3948 ) ;
 assign wire7529 = ( wire3945 ) | ( wire7520  &  wire4277 ) ;
 assign wire7544 = ( (~ preset)  &  wire19065  &  nrq4_2 ) | ( (~ preset)  &  wire7535  &  (~ nrq4_2) ) ;
 assign wire7559 = ( wire3942 ) | ( wire19060  &  wire4383 ) ;
 assign wire7574 = ( wire3940 ) | ( wire4345  &  wire19097 ) ;
 assign wire7589 = ( wire3938 ) | ( wire4345  &  wire19068 ) ;
 assign wire7604 = ( wire7595  &  wire4330 ) | ( wire4374  &  wire19072 ) ;
 assign wire7634 = ( wire19088  &  wire4307 ) | ( wire7625  &  wire4325 ) ;
 assign wire7649 = ( wire3931 ) | ( wire17240  &  wire19073 ) ;
 assign wire7664 = ( wire3929 ) | ( wire17240  &  wire19096 ) ;
 assign wire7679 = ( wire7670  &  wire4277 ) | ( wire4278  &  wire19082 ) ;
 assign wire7694 = ( wire3924 ) | ( wire3925 ) | ( wire18291 ) ;
 assign wire7709 = ( wire18303 ) | ( wire18304 ) | ( wire18309 ) ;
 assign wire7724 = ( wire3901 ) | ( wire3904 ) | ( wire3905 ) | ( wire18312 ) ;
 assign wire7739 = ( wire3895 ) | ( wire3898 ) | ( wire3899 ) | ( wire18316 ) ;
 assign wire7754 = ( wire3894 ) | ( pdata_6_6_  &  wire4352 ) ;
 assign wire7769 = ( (~ preset)  &  pdata_3_3_  &  nrq10_4 ) | ( (~ preset)  &  wire7760  &  (~ nrq10_4) ) ;
 assign wire7784 = ( (~ preset)  &  pdata_12_12_  &  nrq14_3 ) | ( (~ preset)  &  wire7775  &  (~ nrq14_3) ) ;
 assign wire7799 = ( (~ preset)  &  pdata_5_5_  &  nrq14_3 ) | ( (~ preset)  &  wire7790  &  (~ nrq14_3) ) ;
 assign wire7814 = ( wire3886 ) | ( pdata_2_2_  &  wire4354 ) ;
 assign wire7829 = ( wire3884 ) | ( pdata_11_11_  &  wire4354 ) ;
 assign wire7844 = ( wire3881 ) | ( pdata_0_0_  &  wire18384 ) ;
 assign wire7859 = ( wire3879 ) | ( pdata_9_9_  &  wire18384 ) ;
 assign wire7874 = ( wire3877 ) | ( wire3878 ) ;
 assign wire7889 = ( wire3875 ) | ( wire3876 ) ;
 assign wire7904 = ( (~ preset)  &  pdata_8_8_  &  nrq23_3 ) | ( (~ preset)  &  wire7895  &  (~ nrq23_3) ) ;
 assign wire7919 = ( (~ preset)  &  pdata_5_5_  &  nrq23_3 ) | ( (~ preset)  &  wire7910  &  (~ nrq23_3) ) ;
 assign wire7934 = ( (~ preset)  &  pdata_14_14_  &  nrq23_3 ) | ( (~ preset)  &  wire7925  &  (~ nrq23_3) ) ;
 assign wire7949 = ( wire3868 ) | ( pdata_3_3_  &  wire4375 ) ;
 assign wire7964 = ( wire3866 ) | ( pdata_12_12_  &  wire4375 ) ;
 assign wire7979 = ( wire7970  &  wire4340 ) | ( wire17461  &  wire19359 ) ;
 assign wire8009 = ( wire3862 ) | ( wire8000  &  wire4253 ) ;
 assign wire8024 = ( wire3859 ) | ( wire3860 ) ;
 assign wire8039 = ( wire3857 ) | ( wire3858 ) ;
 assign wire8054 = ( wire8045  &  wire4317 ) | ( wire19360  &  wire4381 ) ;
 assign wire8069 = ( wire3853 ) | ( wire8060  &  wire4317 ) ;
 assign wire8084 = ( wire3851 ) | ( wire18501  &  wire19387 ) ;
 assign wire8099 = ( wire3849 ) | ( wire3850 ) ;
 assign wire8114 = ( wire3848 ) | ( wire8105  &  wire4252 ) ;
 assign wire8129 = ( wire3846 ) | ( wire19360  &  wire4377 ) ;
 assign wire8144 = ( wire3843 ) | ( wire3844 ) ;
 assign wire8159 = ( wire3842 ) | ( wire19368  &  wire4377 ) ;
 assign wire8174 = ( (~ preset)  &  wire19097  &  nrq4_2 ) | ( (~ preset)  &  wire8165  &  (~ nrq4_2) ) ;
 assign wire8189 = ( wire3838 ) | ( wire19092  &  wire4383 ) ;
 assign wire8204 = ( wire3836 ) | ( wire4345  &  wire19065 ) ;
 assign wire8219 = ( wire3834 ) | ( wire4345  &  wire4388  &  wire4511 ) | ( wire4345  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire8234 = ( wire8225  &  wire4330 ) | ( wire4374  &  wire19070 ) ;
 assign wire8249 = ( wire8240  &  wire4331 ) | ( wire4332  &  wire19073 ) ;
 assign wire8264 = ( wire19070  &  wire4307 ) | ( wire8255  &  wire4325 ) ;
 assign wire8294 = ( wire3825 ) | ( wire17240  &  wire19091 ) ;
 assign wire8309 = ( wire8300  &  wire4277 ) | ( wire4278  &  wire19103 ) ;
 assign wire8324 = ( wire8315  &  wire4336 ) | ( wire4365  &  wire19068 ) ;
 assign wire8339 = ( wire3818 ) | ( wire3819 ) | ( wire18320 ) ;
 assign wire8354 = ( wire18330 ) | ( wire18331 ) | ( wire18336 ) ;
 assign wire8369 = ( wire3795 ) | ( wire3798 ) | ( wire3799 ) | ( wire18339 ) ;
 assign wire8384 = ( wire3789 ) | ( wire3792 ) | ( wire3793 ) | ( wire18343 ) ;
 assign wire8399 = ( wire3788 ) | ( pdata_9_9_  &  wire4352 ) ;
 assign wire8414 = ( (~ preset)  &  pdata_0_0_  &  nrq10_4 ) | ( (~ preset)  &  wire8405  &  (~ nrq10_4) ) ;
 assign wire8429 = ( (~ preset)  &  pdata_13_13_  &  nrq14_3 ) | ( (~ preset)  &  wire8420  &  (~ nrq14_3) ) ;
 assign wire8444 = ( (~ preset)  &  pdata_8_8_  &  nrq14_3 ) | ( (~ preset)  &  wire8435  &  (~ nrq14_3) ) ;
 assign wire8459 = ( (~ preset)  &  pdata_15_15_  &  nrq14_3 ) | ( (~ preset)  &  wire8450  &  (~ nrq14_3) ) ;
 assign wire8474 = ( wire3777 ) | ( pdata_10_10_  &  wire4354 ) ;
 assign wire8489 = ( wire3773 ) | ( pdata_1_1_  &  wire18384 ) ;
 assign wire8504 = ( wire3771 ) | ( pdata_12_12_  &  wire18384 ) ;
 assign wire8519 = ( wire3768 ) | ( wire3769 ) ;
 assign wire8534 = ( (~ preset)  &  pdata_0_0_  &  nrq23_3 ) | ( (~ preset)  &  wire8525  &  (~ nrq23_3) ) ;
 assign wire8549 = ( (~ preset)  &  pdata_11_11_  &  nrq23_3 ) | ( (~ preset)  &  wire8540  &  (~ nrq23_3) ) ;
 assign wire8564 = ( (~ preset)  &  pdata_2_2_  &  nrq23_3 ) | ( (~ preset)  &  wire8555  &  (~ nrq23_3) ) ;
 assign wire8579 = ( (~ preset)  &  pdata_13_13_  &  nrq23_3 ) | ( (~ preset)  &  wire8570  &  (~ nrq23_3) ) ;
 assign wire8594 = ( wire3759 ) | ( pdata_4_4_  &  wire4375 ) ;
 assign wire8609 = ( wire3757 ) | ( pdata_15_15_  &  wire4375 ) ;
 assign wire8624 = ( wire8615  &  wire4340 ) | ( wire17461  &  wire19387 ) ;
 assign wire8639 = ( wire3751 ) | ( wire4243  &  (~ n_n2471)  &  n_n2487 ) | ( wire4243  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire8654 = ( wire3749 ) | ( wire8645  &  wire4253 ) ;
 assign wire8669 = ( wire3743 ) | ( wire19360  &  wire4306 ) ;
 assign wire8684 = ( wire3741 ) | ( wire19390  &  wire4306 ) ;
 assign wire8699 = ( wire3737 ) | ( wire8690  &  wire4317 ) ;
 assign wire8714 = ( wire3735 ) | ( wire8705  &  wire4317 ) ;
 assign wire8729 = ( wire3733 ) | ( wire18501  &  wire19396 ) ;
 assign wire8744 = ( wire3731 ) | ( wire17305  &  wire19367 ) ;
 assign wire8759 = ( wire3730 ) | ( wire8750  &  wire4252 ) ;
 assign wire8774 = ( wire8765  &  wire4252 ) | ( wire4245  &  wire19368 ) ;
 assign wire8789 = ( wire3725 ) | ( wire19359  &  wire4377 ) ;
 assign wire8819 = ( wire3721 ) | ( wire8810  &  wire4277 ) ;
 assign wire8834 = ( wire3719 ) | ( wire19096  &  wire4383 ) ;
 assign wire8849 = ( wire3716 ) | ( wire4345  &  wire19082 ) ;
 assign wire8864 = ( wire3713 ) | ( wire4345  &  wire19091 ) ;
 assign wire8879 = ( wire8870  &  wire4330 ) | ( wire19088  &  wire4374 ) ;
 assign wire8894 = ( wire8885  &  wire4330 ) | ( wire4374  &  wire19087 ) ;
 assign wire8909 = ( wire3706 ) | ( wire4360  &  wire19070 ) ;
 assign wire8924 = ( wire19072  &  wire4307 ) | ( wire8915  &  wire4325 ) ;
 assign wire8939 = ( wire3701 ) | ( wire17240  &  wire19065 ) ;
 assign wire8954 = ( wire3699 ) | ( wire17240  &  wire19060 ) ;
 assign wire8969 = ( wire8960  &  wire4277 ) | ( wire4278  &  wire19097 ) ;
 assign wire8984 = ( wire8975  &  wire4336 ) | ( wire19103  &  wire4365 ) ;
 assign wire8999 = ( wire18356 ) | ( wire18357 ) | ( wire18362 ) ;
 assign wire9014 = ( wire18373 ) | ( wire18374 ) | ( wire18379 ) ;
 assign wire9029 = ( wire3657 ) | ( wire3660 ) | ( wire3661 ) | ( wire18381 ) ;
 assign wire9044 = ( wire3651 ) | ( wire3654 ) | ( wire3655 ) | ( wire18386 ) ;
 assign wire9059 = ( wire3650 ) | ( pdata_8_8_  &  wire4352 ) ;
 assign wire9074 = ( (~ preset)  &  pdata_1_1_  &  nrq10_4 ) | ( (~ preset)  &  wire9065  &  (~ nrq10_4) ) ;
 assign wire9089 = ( (~ preset)  &  pdata_14_14_  &  nrq14_3 ) | ( (~ preset)  &  wire9080  &  (~ nrq14_3) ) ;
 assign wire9104 = ( (~ preset)  &  pdata_7_7_  &  nrq14_3 ) | ( (~ preset)  &  wire9095  &  (~ nrq14_3) ) ;
 assign wire9119 = ( wire3642 ) | ( pdata_0_0_  &  wire4354 ) ;
 assign wire9134 = ( wire3640 ) | ( pdata_9_9_  &  wire4354 ) ;
 assign wire9149 = ( wire3637 ) | ( pdata_2_2_  &  wire18384 ) ;
 assign wire9164 = ( wire3635 ) | ( pdata_11_11_  &  wire18384 ) ;
 assign wire9179 = ( wire3633 ) | ( wire3634 ) ;
 assign wire9194 = ( (~ preset)  &  pdata_1_1_  &  nrq23_3 ) | ( (~ preset)  &  wire9185  &  (~ nrq23_3) ) ;
 assign wire9209 = ( (~ preset)  &  pdata_10_10_  &  nrq23_3 ) | ( (~ preset)  &  wire9200  &  (~ nrq23_3) ) ;
 assign wire9224 = ( (~ preset)  &  pdata_3_3_  &  nrq23_3 ) | ( (~ preset)  &  wire9215  &  (~ nrq23_3) ) ;
 assign wire9239 = ( (~ preset)  &  pdata_12_12_  &  nrq23_3 ) | ( (~ preset)  &  wire9230  &  (~ nrq23_3) ) ;
 assign wire9254 = ( wire3624 ) | ( pdata_5_5_  &  wire4375 ) ;
 assign wire9269 = ( wire3622 ) | ( pdata_14_14_  &  wire4375 ) ;
 assign wire9284 = ( wire3620 ) | ( wire9275  &  wire4340 ) ;
 assign wire9299 = ( wire9290  &  wire4253 ) | ( wire4243  &  wire19360 ) ;
 assign wire9314 = ( wire3616 ) | ( wire9305  &  wire4253 ) ;
 assign wire9329 = ( wire3613 ) | ( wire3614 ) ;
 assign wire9344 = ( wire3611 ) | ( wire3612 ) ;
 assign wire9359 = ( wire9350  &  wire4317 ) | ( wire4381  &  wire19396 ) ;
 assign wire9374 = ( wire9365  &  wire4317 ) | ( wire19390  &  wire4381 ) ;
 assign wire9389 = ( wire3605 ) | ( wire3606 ) ;
 assign wire9404 = ( wire3603 ) | ( wire17305  &  wire19368 ) ;
 assign wire9419 = ( wire3602 ) | ( wire9410  &  wire4252 ) ;
 assign wire9449 = ( wire3599 ) | ( wire3600 ) ;
 assign wire9464 = ( wire3598 ) | ( wire4278  &  (~ n_n2471)  &  n_n2487 ) | ( wire4278  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire9479 = ( wire9470  &  wire4277 ) | ( wire19359  &  wire4278 ) ;
 assign wire9494 = ( (~ preset)  &  wire19061  &  nrq4_2 ) | ( (~ preset)  &  wire9485  &  (~ nrq4_2) ) ;
 assign wire9509 = ( wire3592 ) | ( wire19091  &  wire4383 ) ;
 assign wire9524 = ( wire3590 ) | ( wire4345  &  wire19103 ) ;
 assign wire9539 = ( wire3588 ) | ( wire4345  &  wire19087 ) ;
 assign wire9554 = ( wire9545  &  wire4330 ) | ( wire4374  &  wire19082 ) ;
 assign wire9569 = ( wire9560  &  wire4330 ) | ( wire4374  &  wire19068 ) ;
 assign wire9584 = ( wire3582 ) | ( wire19088  &  wire4360 ) ;
 assign wire9599 = ( wire19060  &  wire4307 ) | ( wire9590  &  wire4325 ) ;
 assign wire9614 = ( wire3577 ) | ( wire17240  &  wire19061 ) ;
 assign wire9629 = ( wire3575 ) | ( wire17240  &  wire19092 ) ;
 assign wire9644 = ( wire9635  &  wire4277 ) | ( wire4278  &  wire19065 ) ;
 assign wire9659 = ( wire9650  &  wire4277 ) | ( wire4278  &  wire19096 ) ;
 assign wire9674 = ( wire3570 ) | ( pdata_1_1_  &  wire4357 ) ;
 assign wire9689 = ( wire3568 ) | ( pdata_12_12_  &  wire4357 ) ;
 assign wire9704 = ( wire3562 ) | ( wire3563 ) | ( wire1427  &  wire4199 ) ;
 assign wire9719 = ( (~ preset)  &  pdata_2_2_  &  nrq23_3 ) | ( (~ preset)  &  wire9710  &  (~ nrq23_3) ) ;
 assign wire9734 = ( wire3559 ) | ( wire9725  &  wire4253 ) ;
 assign wire9749 = ( wire3557 ) | ( wire9740  &  wire4253 ) ;
 assign wire9779 = ( wire3555 ) | ( wire9770  &  wire4252 ) ;
 assign wire9794 = ( wire3552 ) | ( wire3553 ) ;
 assign wire9809 = ( wire3551 ) | ( wire19087  &  wire4383 ) ;
 assign wire9824 = ( wire3549 ) | ( wire4345  &  wire19070 ) ;
 assign wire9839 = ( wire9830  &  wire4330 ) | ( wire4374  &  wire19061 ) ;
 assign wire9854 = ( wire9845  &  wire4330 ) | ( wire4374  &  wire19091 ) ;
 assign wire9869 = ( wire19092  &  wire4307 ) | ( wire9860  &  wire4325 ) ;
 assign wire9884 = ( wire3540 ) | ( wire17240  &  wire19103 ) ;
 assign wire9899 = ( wire3538 ) | ( wire17240  &  wire4388  &  wire4511 ) | ( wire17240  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire9914 = ( wire9905  &  wire4277 ) | ( wire4278  &  wire19060 ) ;
 assign wire9929 = ( wire9920  &  wire4336 ) | ( wire19097  &  wire4365 ) ;
 assign wire9944 = ( wire3533 ) | ( pdata_0_0_  &  wire4357 ) ;
 assign wire9959 = ( wire3531 ) | ( pdata_6_6_  &  wire4358 ) ;
 assign wire9989 = ( (~ preset)  &  pdata_12_12_  &  nrq23_3 ) | ( (~ preset)  &  wire9980  &  (~ nrq23_3) ) ;
 assign wire10004 = ( wire9995  &  wire4253 ) | ( wire4243  &  wire19396 ) ;
 assign wire10019 = ( wire10010  &  wire4253 ) | ( wire4243  &  wire19390 ) ;
 assign wire10034 = ( wire3522 ) | ( wire4245  &  (~ n_n2471)  &  n_n2487 ) | ( wire4245  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire10049 = ( wire10040  &  wire4252 ) | ( wire4245  &  wire19359 ) ;
 assign wire10064 = ( wire3519 ) | ( wire4377  &  wire19367 ) ;
 assign wire10079 = ( wire3517 ) | ( wire4383  &  wire19068 ) ;
 assign wire10094 = ( wire3515 ) | ( wire19088  &  wire4345 ) ;
 assign wire10109 = ( wire10100  &  wire4330 ) | ( wire4374  &  wire19065 ) ;
 assign wire10124 = ( wire10115  &  wire4330 ) | ( wire4374  &  wire19096 ) ;
 assign wire10139 = ( wire19096  &  wire4307 ) | ( wire10130  &  wire4325 ) ;
 assign wire10154 = ( wire3506 ) | ( wire17240  &  wire19097 ) ;
 assign wire10184 = ( wire10175  &  wire4277 ) | ( wire4278  &  wire19072 ) ;
 assign wire10199 = ( wire10190  &  wire4336 ) | ( wire4365  &  wire19087 ) ;
 assign wire10214 = ( wire3501 ) | ( pdata_10_10_  &  wire4357 ) ;
 assign wire10229 = ( wire3499 ) | ( pdata_5_5_  &  wire4358 ) ;
 assign wire10244 = ( wire3496 ) | ( wire12200  &  wire5513 ) | ( wire12200  &  wire5514 ) ;
 assign wire10259 = ( wire3491 ) | ( wire3492 ) | ( wire4199  &  wire1342 ) ;
 assign wire10274 = ( (~ preset)  &  pdata_6_6_  &  nrq23_3 ) | ( (~ preset)  &  wire10265  &  (~ nrq23_3) ) ;
 assign wire10289 = ( wire3487 ) | ( wire3488 ) ;
 assign wire10319 = ( wire10310  &  wire4252 ) | ( wire4245  &  wire19360 ) ;
 assign wire10334 = ( wire3483 ) | ( wire3484 ) ;
 assign wire10349 = ( wire3481 ) | ( wire3482 ) ;
 assign wire10364 = ( wire3480 ) | ( wire4383  &  wire4388  &  wire4511 ) | ( wire4383  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire10379 = ( wire3478 ) | ( wire4345  &  wire19060 ) ;
 assign wire10409 = ( wire10400  &  wire4330 ) | ( wire19092  &  wire4374 ) ;
 assign wire10424 = ( wire19091  &  wire4307 ) | ( wire10415  &  wire4325 ) ;
 assign wire10439 = ( wire3471 ) | ( wire17240  &  wire19088 ) ;
 assign wire10454 = ( wire3469 ) | ( wire17240  &  wire19087 ) ;
 assign wire10469 = ( wire10460  &  wire4277 ) | ( wire4278  &  wire19070 ) ;
 assign wire10484 = ( wire3466 ) | ( pdata_2_2_  &  wire4357 ) ;
 assign wire10499 = ( wire3464 ) | ( pdata_11_11_  &  wire4357 ) ;
 assign wire10514 = ( wire3462 ) | ( pdata_4_4_  &  wire4358 ) ;
 assign wire10529 = ( wire3459 ) | ( wire12080  &  wire5513 ) | ( wire12080  &  wire5514 ) ;
 assign wire10544 = ( wire3454 ) | ( wire3455 ) | ( wire4199  &  wire1353 ) ;
 assign wire10559 = ( wire3453 ) | ( pdata_0_0_  &  wire4375 ) ;
 assign wire10574 = ( wire3450 ) | ( wire4306  &  wire19387 ) ;
 assign wire10589 = ( wire3448 ) | ( wire4306  &  wire19368 ) ;
 assign wire10604 = ( wire3447 ) | ( wire10595  &  wire4252 ) ;
 assign wire10619 = ( wire3445 ) | ( wire4377  &  wire19396 ) ;
 assign wire10634 = ( wire3443 ) | ( wire19390  &  wire4377 ) ;
 assign wire10664 = ( wire3441 ) | ( wire4345  &  wire19072 ) ;
 assign wire10679 = ( wire10670  &  wire4330 ) | ( wire4374  &  wire19073 ) ;
 assign wire10694 = ( wire10685  &  wire4330 ) | ( wire4374  &  wire19060 ) ;
 assign wire10709 = ( wire19087  &  wire4307 ) | ( wire10700  &  wire4325 ) ;
 assign wire10724 = ( wire3432 ) | ( wire17240  &  wire19082 ) ;
 assign wire10739 = ( wire3430 ) | ( wire17240  &  wire19068 ) ;
 assign wire10754 = ( wire10745  &  wire4277 ) | ( wire4278  &  wire19088 ) ;
 assign wire10769 = ( wire3426 ) | ( pdata_13_13_  &  wire4305 ) ;
 assign wire10784 = ( wire3425 ) | ( pdata_8_8_  &  wire4357 ) ;
 assign wire10799 = ( wire3423 ) | ( pdata_3_3_  &  wire4358 ) ;
 assign wire10814 = ( wire3421 ) | ( pdata_1_1_  &  wire4359 ) ;
 assign wire10829 = ( wire3419 ) | ( pdata_12_12_  &  wire4359 ) ;
 assign wire10859 = ( wire3417 ) | ( pdata_10_10_  &  wire4375 ) ;
 assign wire10874 = ( wire3414 ) | ( wire10865  &  wire4317 ) ;
 assign wire10889 = ( wire3412 ) | ( wire3413 ) ;
 assign wire10904 = ( wire3410 ) | ( wire10895  &  wire4277 ) ;
 assign wire10934 = ( (~ preset)  &  wire19092  &  nrq4_2 ) | ( (~ preset)  &  wire10925  &  (~ nrq4_2) ) ;
 assign wire10949 = ( wire3407 ) | ( wire4360  &  wire19065 ) ;
 assign wire10964 = ( wire3405 ) | ( wire4360  &  wire19087 ) ;
 assign wire10979 = ( wire10970  &  wire4331 ) | ( wire4332  &  wire19070 ) ;
 assign wire10994 = ( wire10985  &  wire4325 ) | ( wire4307  &  wire19068 ) ;
 assign wire11024 = ( wire11015  &  wire4336 ) | ( wire19092  &  wire4365 ) ;
 assign wire11039 = ( wire3396 ) | ( pdata_12_12_  &  wire4305 ) ;
 assign wire11054 = ( wire3395 ) | ( pdata_9_9_  &  wire4357 ) ;
 assign wire11069 = ( wire3393 ) | ( pdata_2_2_  &  wire4358 ) ;
 assign wire11084 = ( wire3391 ) | ( pdata_7_7_  &  wire4358 ) ;
 assign wire11099 = ( wire3389 ) | ( pdata_13_13_  &  wire4359 ) ;
 assign wire11129 = ( wire3387 ) | ( wire11120  &  wire4340 ) ;
 assign wire11144 = ( wire11135  &  wire4317 ) | ( wire4381  &  wire19359 ) ;
 assign wire11159 = ( wire3382 ) | ( wire18501  &  wire19360 ) ;
 assign wire11174 = ( wire11165  &  wire4277 ) | ( wire4278  &  wire19387 ) ;
 assign wire11189 = ( wire11180  &  wire4277 ) | ( wire19368  &  wire4278 ) ;
 assign wire11204 = ( wire3377 ) | ( wire4360  &  wire19097 ) ;
 assign wire11219 = ( wire3375 ) | ( wire4360  &  wire19091 ) ;
 assign wire11234 = ( wire11225  &  wire4331 ) | ( wire4332  &  wire19072 ) ;
 assign wire11249 = ( wire3370 ) | ( wire17240  &  wire19070 ) ;
 assign wire11264 = ( wire11255  &  wire4336 ) | ( wire4365  &  wire19073 ) ;
 assign wire11279 = ( wire11270  &  wire4336 ) | ( wire19060  &  wire4365 ) ;
 assign wire11294 = ( wire3364 ) | ( pdata_15_15_  &  wire4305 ) ;
 assign wire11309 = ( wire3363 ) | ( pdata_6_6_  &  wire4357 ) ;
 assign wire11324 = ( wire3361 ) | ( pdata_1_1_  &  wire4358 ) ;
 assign wire11339 = ( wire3359 ) | ( pdata_8_8_  &  wire4358 ) ;
 assign wire11354 = ( wire3357 ) | ( pdata_3_3_  &  wire4359 ) ;
 assign wire11384 = ( wire11375  &  wire4340 ) | ( wire17461  &  wire19367 ) ;
 assign wire11399 = ( wire3352 ) | ( wire3353 ) ;
 assign wire11414 = ( wire3350 ) | ( wire11405  &  wire4277 ) ;
 assign wire11429 = ( (~ preset)  &  wire19072  &  nrq4_2 ) | ( (~ preset)  &  wire11420  &  (~ nrq4_2) ) ;
 assign wire11444 = ( wire3347 ) | ( wire19103  &  wire4360 ) ;
 assign wire11459 = ( wire3345 ) | ( wire4360  &  wire4388  &  wire4511 ) | ( wire4360  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire11474 = ( wire11465  &  wire4331 ) | ( wire4332  &  wire19082 ) ;
 assign wire11489 = ( wire11480  &  wire4277 ) | ( wire4278  &  wire19073 ) ;
 assign wire11504 = ( wire11495  &  wire4336 ) | ( wire19061  &  wire4365 ) ;
 assign wire11519 = ( wire11510  &  wire4336 ) | ( wire19091  &  wire4365 ) ;
 assign wire11534 = ( wire3334 ) | ( pdata_14_14_  &  wire4305 ) ;
 assign wire11549 = ( wire3333 ) | ( pdata_7_7_  &  wire4357 ) ;
 assign wire11564 = ( wire3331 ) | ( pdata_0_0_  &  wire4358 ) ;
 assign wire11579 = ( wire3329 ) | ( pdata_9_9_  &  wire4358 ) ;
 assign wire11594 = ( wire3327 ) | ( pdata_2_2_  &  wire4359 ) ;
 assign wire11609 = ( wire3325 ) | ( pdata_11_11_  &  wire4359 ) ;
 assign wire11624 = ( wire3322 ) | ( wire18501  &  wire19390 ) ;
 assign wire11639 = ( (~ preset)  &  wire19073  &  nrq4_2 ) | ( (~ preset)  &  wire11630  &  (~ nrq4_2) ) ;
 assign wire11654 = ( (~ preset)  &  wire19060  &  nrq4_2 ) | ( (~ preset)  &  wire11645  &  (~ nrq4_2) ) ;
 assign wire11669 = ( wire3317 ) | ( wire4360  &  wire19082 ) ;
 assign wire11684 = ( wire3315 ) | ( wire4360  &  wire19068 ) ;
 assign wire11699 = ( wire11690  &  wire4331 ) | ( wire19088  &  wire4332 ) ;
 assign wire11714 = ( wire11705  &  wire4277 ) | ( wire4278  &  wire19092 ) ;
 assign wire11729 = ( wire11720  &  wire4336 ) | ( wire4365  &  wire19065 ) ;
 assign wire11744 = ( wire11735  &  wire4336 ) | ( wire4365  &  wire19096 ) ;
 assign wire11759 = ( wire3304 ) | ( pdata_9_9_  &  wire4305 ) ;
 assign wire11774 = ( wire3303 ) | ( pdata_4_4_  &  wire4357 ) ;
 assign wire11789 = ( wire3301 ) | ( pdata_15_15_  &  wire4357 ) ;
 assign wire11804 = ( wire3299 ) | ( pdata_10_10_  &  wire4358 ) ;
 assign wire11819 = ( wire3297 ) | ( pdata_5_5_  &  wire4359 ) ;
 assign wire11864 = ( wire3293 ) | ( wire3294 ) | ( wire4199  &  wire1412 ) ;
 assign wire11879 = ( wire18401 ) | ( wire18402 ) | ( wire18406 ) ;
 assign wire11894 = ( wire3280 ) | ( pdata_5_5_  &  wire4357 ) ;
 assign wire11909 = ( wire3278 ) | ( pdata_14_14_  &  wire4357 ) ;
 assign wire11924 = ( wire3276 ) | ( pdata_11_11_  &  wire4358 ) ;
 assign wire11939 = ( wire3274 ) | ( pdata_4_4_  &  wire4359 ) ;
 assign wire11984 = ( wire3270 ) | ( wire3271 ) | ( wire4199  &  wire1397 ) ;
 assign wire11999 = ( wire3268 ) | ( wire18414 ) | ( wire18416 ) | ( wire18417 ) ;
 assign wire12014 = ( wire12005  &  wire4316 ) | ( wire19061  &  wire4327 ) ;
 assign wire12029 = ( wire3254 ) | ( pdata_11_11_  &  wire4305 ) ;
 assign wire12044 = ( wire3253 ) | ( pdata_13_13_  &  wire4357 ) ;
 assign wire12059 = ( wire3251 ) | ( pdata_12_12_  &  wire4358 ) ;
 assign wire12074 = ( wire3249 ) | ( pdata_7_7_  &  wire4359 ) ;
 assign wire12089 = ( wire3247 ) | ( pdata_14_14_  &  wire4359 ) ;
 assign wire12119 = ( wire3241 ) | ( wire3242 ) | ( wire4199  &  wire1439 ) ;
 assign wire12134 = ( wire12125  &  wire4316 ) | ( wire19096  &  wire4327 ) ;
 assign wire12149 = ( wire3237 ) | ( pdata_10_10_  &  wire4305 ) ;
 assign wire12164 = ( wire3236 ) | ( pdata_3_3_  &  wire4357 ) ;
 assign wire12179 = ( wire3234 ) | ( pdata_13_13_  &  wire4358 ) ;
 assign wire12194 = ( wire3232 ) | ( pdata_6_6_  &  wire4359 ) ;
 assign wire12209 = ( wire3230 ) | ( pdata_15_15_  &  wire4359 ) ;
 assign wire12239 = ( wire3227 ) | ( wire18427 ) | ( wire18429 ) | ( wire18430 ) ;
 assign wire12254 = ( wire19103  &  wire4307 ) | ( wire12245  &  wire4325 ) ;
 assign wire12269 = ( wire3214 ) | ( pdata_14_14_  &  wire4358 ) ;
 assign wire12284 = ( wire3212 ) | ( pdata_9_9_  &  wire4359 ) ;
 assign wire12314 = ( wire3209 ) | ( wire11090  &  wire5513 ) | ( wire11090  &  wire5514 ) ;
 assign wire12329 = ( wire3204 ) | ( wire3205 ) | ( wire4199  &  wire1368 ) ;
 assign wire12344 = ( wire3203 ) | ( wire12335  &  wire4280 ) ;
 assign wire12359 = ( wire3200 ) | ( wire3201 ) ;
 assign wire12374 = ( wire3198 ) | ( wire16928  &  wire19368 ) ;
 assign wire12389 = ( wire3197 ) | ( wire19061  &  wire4368 ) ;
 assign wire12404 = ( wire3195 ) | ( wire19091  &  wire4368 ) ;
 assign wire12419 = ( wire3193 ) | ( wire19088  &  wire4383 ) ;
 assign wire12434 = ( wire3191 ) | ( wire4332  &  wire4388  &  wire4511 ) | ( wire4332  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire12449 = ( wire12440  &  wire4316 ) | ( wire19060  &  wire4327 ) ;
 assign wire12464 = ( wire19097  &  wire4307 ) | ( wire12455  &  wire4325 ) ;
 assign wire12479 = ( wire3185 ) | ( pdata_15_15_  &  wire4358 ) ;
 assign wire12494 = ( wire3183 ) | ( pdata_8_8_  &  wire4359 ) ;
 assign wire12524 = ( wire3180 ) | ( wire10820  &  wire5513 ) | ( wire10820  &  wire5514 ) ;
 assign wire12539 = ( wire3175 ) | ( wire3176 ) | ( wire4199  &  wire1386 ) ;
 assign wire12554 = ( wire3173 ) | ( wire3174 ) ;
 assign wire12569 = ( wire12560  &  wire4280 ) | ( wire18176  &  wire19387 ) ;
 assign wire12584 = ( wire3169 ) | ( wire16928  &  wire19396 ) ;
 assign wire12599 = ( wire3167 ) | ( wire3168 ) ;
 assign wire12614 = ( wire3166 ) | ( wire19073  &  wire4368 ) ;
 assign wire12629 = ( wire3164 ) | ( wire19087  &  wire4368 ) ;
 assign wire12644 = ( wire3162 ) | ( wire19082  &  wire4383 ) ;
 assign wire12659 = ( wire12650  &  wire4331 ) | ( wire4332  &  wire19068 ) ;
 assign wire12674 = ( wire12665  &  wire4316 ) | ( wire19092  &  wire4327 ) ;
 assign wire12689 = ( wire12680  &  wire4325 ) | ( wire4307  &  wire19065 ) ;
 assign wire12704 = ( wire3154 ) | ( pdata_0_0_  &  wire4359 ) ;
 assign wire12749 = ( wire3150 ) | ( wire3151 ) | ( wire4199  &  wire1411 ) ;
 assign wire12764 = ( wire3145 ) | ( wire3146 ) | ( wire4199  &  wire1398 ) ;
 assign wire12779 = ( wire3143 ) | ( wire3144 ) ;
 assign wire12809 = ( wire3141 ) | ( wire3142 ) ;
 assign wire12824 = ( wire3139 ) | ( wire3140 ) ;
 assign wire12839 = ( wire3137 ) | ( wire3138 ) ;
 assign wire12854 = ( wire3136 ) | ( wire19097  &  wire4368 ) ;
 assign wire12869 = ( wire3134 ) | ( wire19092  &  wire4368 ) ;
 assign wire12884 = ( wire3132 ) | ( wire19103  &  wire4383 ) ;
 assign wire12899 = ( wire12890  &  wire4316 ) | ( wire19073  &  wire4327 ) ;
 assign wire12914 = ( wire12905  &  wire4316 ) | ( wire19070  &  wire4327 ) ;
 assign wire12929 = ( wire19061  &  wire4307 ) | ( wire12920  &  wire4325 ) ;
 assign wire12944 = ( wire3124 ) | ( pdata_10_10_  &  wire4359 ) ;
 assign wire12989 = ( wire3120 ) | ( wire3121 ) | ( wire4199  &  wire1434 ) ;
 assign wire13004 = ( wire3115 ) | ( wire3116 ) | ( wire4199  &  wire1413 ) ;
 assign wire13019 = ( wire3113 ) | ( wire3114 ) ;
 assign wire13034 = ( wire3111 ) | ( wire4308  &  (~ n_n2471)  &  n_n2487 ) | ( wire4308  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire13049 = ( wire3109 ) | ( wire4308  &  wire19359 ) ;
 assign wire13064 = ( wire3107 ) | ( wire3108 ) ;
 assign wire13079 = ( wire3105 ) | ( wire16928  &  wire19367 ) ;
 assign wire13094 = ( wire3103 ) | ( wire17305  &  wire19387 ) ;
 assign wire13109 = ( wire3102 ) | ( wire19065  &  wire4368 ) ;
 assign wire13124 = ( wire3100 ) | ( wire19096  &  wire4368 ) ;
 assign wire13139 = ( wire3098 ) | ( wire19097  &  wire4383 ) ;
 assign wire13169 = ( wire13160  &  wire4316 ) | ( wire19072  &  wire4327 ) ;
 assign wire13184 = ( wire19073  &  wire4307 ) | ( wire13175  &  wire4325 ) ;
 assign wire13199 = ( wire18445 ) | ( wire18446 ) | ( wire18451 ) ;
 assign wire13214 = ( wire18458 ) | ( wire18459 ) | ( wire18463 ) ;
 assign wire13229 = ( wire3066 ) | ( pdata_3_3_  &  wire4352 ) ;
 assign wire13244 = ( wire3064 ) | ( pdata_14_14_  &  wire4352 ) ;
 assign wire13259 = ( (~ preset)  &  pdata_14_14_  &  nrq10_4 ) | ( (~ preset)  &  wire13250  &  (~ nrq10_4) ) ;
 assign wire13274 = ( wire3060 ) | ( pdata_9_9_  &  wire4353 ) ;
 assign wire13289 = ( (~ preset)  &  pdata_4_4_  &  nrq14_3 ) | ( (~ preset)  &  wire13280  &  (~ nrq14_3) ) ;
 assign wire13304 = ( wire3055 ) | ( wire3056 ) ;
 assign wire13319 = ( wire3053 ) | ( wire3054 ) ;
 assign wire13334 = ( wire3051 ) | ( wire3052 ) ;
 assign wire13349 = ( wire3049 ) | ( wire3050 ) ;
 assign wire13364 = ( wire13355  &  wire4280 ) | ( wire18176  &  wire19396 ) ;
 assign wire13379 = ( wire13370  &  wire4280 ) | ( wire18176  &  wire19367 ) ;
 assign wire13394 = ( wire3043 ) | ( wire3044 ) ;
 assign wire13409 = ( wire3041 ) | ( wire16928  &  (~ n_n2471)  &  n_n2487 ) | ( wire16928  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire13424 = ( wire3039 ) | ( wire3040 ) ;
 assign wire13439 = ( wire3037 ) | ( wire3038 ) ;
 assign wire13454 = ( (~ preset)  &  wire19068  &  nrq4_2 ) | ( (~ preset)  &  wire13445  &  (~ nrq4_2) ) ;
 assign wire13469 = ( wire3034 ) | ( wire19072  &  wire4368 ) ;
 assign wire13484 = ( wire3032 ) | ( wire4383  &  wire19065 ) ;
 assign wire13499 = ( wire13490  &  wire4331 ) | ( wire4332  &  wire19096 ) ;
 assign wire13514 = ( wire13505  &  wire4316 ) | ( wire19082  &  wire4327 ) ;
 assign wire13544 = ( wire18470 ) | ( wire18471 ) | ( wire18476 ) ;
 assign wire13559 = ( wire3012 ) | ( wire3013 ) | ( wire18477 ) ;
 assign wire13574 = ( wire3005 ) | ( wire3008 ) | ( wire3009 ) | ( wire18481 ) ;
 assign wire13589 = ( wire3004 ) | ( pdata_15_15_  &  wire4352 ) ;
 assign wire13604 = ( (~ preset)  &  pdata_13_13_  &  nrq10_4 ) | ( (~ preset)  &  wire13595  &  (~ nrq10_4) ) ;
 assign wire13619 = ( wire3000 ) | ( pdata_10_10_  &  wire4353 ) ;
 assign wire13634 = ( (~ preset)  &  pdata_3_3_  &  nrq14_3 ) | ( (~ preset)  &  wire13625  &  (~ nrq14_3) ) ;
 assign wire13649 = ( wire2995 ) | ( wire2996 ) ;
 assign wire13664 = ( wire2993 ) | ( wire2994 ) ;
 assign wire13679 = ( wire2991 ) | ( wire2992 ) ;
 assign wire13694 = ( wire2989 ) | ( wire2990 ) ;
 assign wire13709 = ( wire2988 ) | ( wire13700  &  wire4340 ) ;
 assign wire13724 = ( wire2986 ) | ( wire13715  &  wire4280 ) ;
 assign wire13739 = ( wire13730  &  wire4280 ) | ( wire18176  &  wire19368 ) ;
 assign wire13754 = ( wire2981 ) | ( wire2982 ) ;
 assign wire13784 = ( wire2979 ) | ( wire16928  &  wire19390 ) ;
 assign wire13799 = ( wire2977 ) | ( wire2978 ) ;
 assign wire13814 = ( (~ preset)  &  wire19087  &  nrq4_2 ) | ( (~ preset)  &  wire13805  &  (~ nrq4_2) ) ;
 assign wire13829 = ( wire2974 ) | ( wire19060  &  wire4368 ) ;
 assign wire13844 = ( wire2972 ) | ( wire19061  &  wire4383 ) ;
 assign wire13859 = ( wire13850  &  wire4331 ) | ( wire19092  &  wire4332 ) ;
 assign wire13874 = ( wire13865  &  wire4316 ) | ( wire19088  &  wire4327 ) ;
 assign wire13889 = ( wire2966 ) | ( wire4327  &  wire4388  &  wire4511 ) | ( wire4327  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire13904 = ( wire2963 ) | ( pdata_8_8_  &  wire4305 ) ;
 assign wire13919 = ( wire18491 ) | ( wire18492 ) | ( wire18497 ) ;
 assign wire13934 = ( wire2946 ) | ( wire18507 ) | ( wire18511 ) ;
 assign wire13949 = ( wire2927 ) | ( wire2930 ) | ( wire2931 ) | ( wire18513 ) ;
 assign wire13964 = ( wire2926 ) | ( pdata_5_5_  &  wire4352 ) ;
 assign wire13979 = ( wire2924 ) | ( pdata_0_0_  &  wire4353 ) ;
 assign wire13994 = ( wire2922 ) | ( pdata_7_7_  &  wire4353 ) ;
 assign wire14009 = ( (~ preset)  &  pdata_2_2_  &  nrq14_3 ) | ( (~ preset)  &  wire14000  &  (~ nrq14_3) ) ;
 assign wire14024 = ( wire2918 ) | ( pdata_13_13_  &  wire4354 ) ;
 assign wire14039 = ( wire2915 ) | ( pdata_8_8_  &  wire18384 ) ;
 assign wire14054 = ( wire2913 ) | ( wire2914 ) ;
 assign wire14069 = ( wire2911 ) | ( wire2912 ) ;
 assign wire14084 = ( wire2909 ) | ( wire2910 ) ;
 assign wire14099 = ( wire2908 ) | ( pdata_11_11_  &  wire4375 ) ;
 assign wire14114 = ( wire2906 ) | ( wire14105  &  wire4280 ) ;
 assign wire14129 = ( wire14120  &  wire4280 ) | ( wire18176  &  wire19390 ) ;
 assign wire14144 = ( wire2901 ) | ( wire4308  &  wire19387 ) ;
 assign wire14159 = ( wire2899 ) | ( wire2900 ) ;
 assign wire14174 = ( wire2897 ) | ( wire16928  &  wire19359 ) ;
 assign wire14189 = ( wire2895 ) | ( wire17305  &  wire19396 ) ;
 assign wire14219 = ( wire2894 ) | ( wire19088  &  wire4368 ) ;
 assign wire14234 = ( wire2892 ) | ( wire4383  &  wire19073 ) ;
 assign wire14249 = ( wire14240  &  wire4331 ) | ( wire4332  &  wire19087 ) ;
 assign wire14264 = ( wire14255  &  wire4316 ) | ( wire19097  &  wire4327 ) ;
 assign wire14279 = ( wire14270  &  wire4316 ) | ( wire19068  &  wire4327 ) ;
 assign wire14294 = ( wire2883 ) | ( pdata_7_7_  &  wire4305 ) ;
 assign wire14309 = ( wire2881 ) | ( wire18522 ) | ( wire18523 ) | ( wire18524 ) ;
 assign wire14324 = ( wire2870 ) | ( wire18535 ) | ( wire18539 ) ;
 assign wire14339 = ( wire2856 ) | ( wire18549 ) | ( wire18553 ) ;
 assign wire14354 = ( wire2837 ) | ( wire2840 ) | ( wire2841 ) | ( wire18556 ) ;
 assign wire14369 = ( wire2836 ) | ( pdata_4_4_  &  wire4352 ) ;
 assign wire14384 = ( wire2834 ) | ( pdata_13_13_  &  wire4352 ) ;
 assign wire14399 = ( (~ preset)  &  pdata_15_15_  &  nrq10_4 ) | ( (~ preset)  &  wire14390  &  (~ nrq10_4) ) ;
 assign wire14414 = ( wire2830 ) | ( pdata_8_8_  &  wire4353 ) ;
 assign wire14429 = ( (~ preset)  &  pdata_1_1_  &  nrq14_3 ) | ( (~ preset)  &  wire14420  &  (~ nrq14_3) ) ;
 assign wire14444 = ( wire2826 ) | ( pdata_14_14_  &  wire4354 ) ;
 assign wire14459 = ( wire2823 ) | ( pdata_7_7_  &  wire18384 ) ;
 assign wire14474 = ( wire2821 ) | ( wire2822 ) ;
 assign wire14489 = ( wire2819 ) | ( wire2820 ) ;
 assign wire14504 = ( wire2817 ) | ( wire2818 ) ;
 assign wire14519 = ( wire2816 ) | ( pdata_1_1_  &  wire4375 ) ;
 assign wire14534 = ( wire2814 ) | ( wire14525  &  wire4280 ) ;
 assign wire14549 = ( wire2812 ) | ( wire14540  &  wire4280 ) ;
 assign wire14564 = ( wire2809 ) | ( wire2810 ) ;
 assign wire14579 = ( wire2807 ) | ( wire16928  &  wire19360 ) ;
 assign wire14594 = ( wire2805 ) | ( wire2806 ) ;
 assign wire14609 = ( wire2803 ) | ( wire2804 ) ;
 assign wire14624 = ( wire2802 ) | ( wire4350  &  wire4388  &  wire4511 ) | ( wire4350  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire14639 = ( wire2800 ) | ( wire19070  &  wire4368 ) ;
 assign wire14669 = ( wire14660  &  wire4331 ) | ( wire4332  &  wire19091 ) ;
 assign wire14684 = ( wire14675  &  wire4316 ) | ( wire19103  &  wire4327 ) ;
 assign wire14699 = ( wire14690  &  wire4316 ) | ( wire19087  &  wire4327 ) ;
 assign wire14714 = ( wire2791 ) | ( pdata_6_6_  &  wire4305 ) ;
 assign wire14729 = ( wire2789 ) | ( wire18564 ) | ( wire18565 ) | ( wire18566 ) ;
 assign wire14744 = ( wire18577 ) | ( wire18578 ) | ( wire18583 ) ;
 assign wire14759 = ( wire2764 ) | ( wire18592 ) | ( wire18598 ) ;
 assign wire14774 = ( wire2748 ) | ( wire2749 ) | ( wire18599 ) ;
 assign wire14789 = ( wire18611 ) | ( wire18612 ) | ( wire18616 ) ;
 assign wire14804 = ( wire2725 ) | ( wire2728 ) | ( wire2729 ) | ( wire18619 ) ;
 assign wire14819 = ( (~ preset)  &  pdata_10_10_  &  nrq10_4 ) | ( (~ preset)  &  wire14810  &  (~ nrq10_4) ) ;
 assign wire14834 = ( wire2722 ) | ( pdata_5_5_  &  wire4353 ) ;
 assign wire14849 = ( (~ preset)  &  pdata_0_0_  &  nrq14_3 ) | ( (~ preset)  &  wire14840  &  (~ nrq14_3) ) ;
 assign wire14864 = ( (~ preset)  &  pdata_9_9_  &  nrq14_3 ) | ( (~ preset)  &  wire14855  &  (~ nrq14_3) ) ;
 assign wire14879 = ( wire2716 ) | ( pdata_4_4_  &  wire4354 ) ;
 assign wire14894 = ( wire2713 ) | ( wire2714 ) ;
 assign wire14909 = ( wire2711 ) | ( wire2712 ) ;
 assign wire14924 = ( wire2709 ) | ( wire2710 ) ;
 assign wire14939 = ( (~ preset)  &  pdata_7_7_  &  nrq23_3 ) | ( (~ preset)  &  wire14930  &  (~ nrq23_3) ) ;
 assign wire14969 = ( wire2706 ) | ( wire14960  &  wire4280 ) ;
 assign wire14984 = ( wire2703 ) | ( wire2704 ) ;
 assign wire14999 = ( wire2701 ) | ( wire2702 ) ;
 assign wire15014 = ( wire2699 ) | ( wire2700 ) ;
 assign wire15029 = ( wire2697 ) | ( wire17305  &  wire19360 ) ;
 assign wire15044 = ( wire2696 ) | ( wire19103  &  wire4368 ) ;
 assign wire15059 = ( wire2694 ) | ( wire4368  &  wire4388  &  wire4511 ) | ( wire4368  &  (~ wire4388)  &  (~ wire4511) ) ;
 assign wire15074 = ( wire15065  &  wire4316 ) | ( wire19091  &  wire4327 ) ;
 assign wire15089 = ( wire2689 ) | ( pdata_5_5_  &  wire4305 ) ;
 assign wire15104 = ( wire2687 ) | ( wire18627 ) | ( wire18628 ) | ( wire18629 ) ;
 assign wire15119 = ( wire18640 ) | ( wire18641 ) | ( wire18646 ) ;
 assign wire15134 = ( wire2662 ) | ( wire18654 ) | ( wire18658 ) ;
 assign wire15149 = ( wire2646 ) | ( wire2647 ) | ( wire18659 ) ;
 assign wire15164 = ( wire18669 ) | ( wire18670 ) | ( wire18674 ) ;
 assign wire15179 = ( wire2623 ) | ( wire2626 ) | ( wire2627 ) | ( wire18676 ) ;
 assign wire15194 = ( (~ preset)  &  pdata_9_9_  &  nrq10_4 ) | ( (~ preset)  &  wire15185  &  (~ nrq10_4) ) ;
 assign wire15209 = ( wire2620 ) | ( pdata_6_6_  &  wire4353 ) ;
 assign wire15224 = ( wire2618 ) | ( pdata_15_15_  &  wire4353 ) ;
 assign wire15239 = ( (~ preset)  &  pdata_10_10_  &  nrq14_3 ) | ( (~ preset)  &  wire15230  &  (~ nrq14_3) ) ;
 assign wire15254 = ( wire2614 ) | ( pdata_3_3_  &  wire4354 ) ;
 assign wire15269 = ( wire2611 ) | ( wire2612 ) ;
 assign wire15284 = ( wire2609 ) | ( wire2610 ) ;
 assign wire15299 = ( wire2607 ) | ( wire2608 ) ;
 assign wire15314 = ( (~ preset)  &  pdata_13_13_  &  nrq23_3 ) | ( (~ preset)  &  wire15305  &  (~ nrq23_3) ) ;
 assign wire15329 = ( wire15320  &  wire4340 ) | ( wire17461  &  wire19368 ) ;
 assign wire15344 = ( wire2602 ) | ( wire15335  &  wire4280 ) ;
 assign wire15359 = ( wire2599 ) | ( wire4308  &  wire19396 ) ;
 assign wire15374 = ( wire2597 ) | ( wire2598 ) ;
 assign wire15389 = ( wire2595 ) | ( wire17305  &  (~ n_n2471)  &  n_n2487 ) | ( wire17305  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire15404 = ( wire2594 ) | ( wire19082  &  wire4368 ) ;
 assign wire15419 = ( wire2592 ) | ( wire19068  &  wire4368 ) ;
 assign wire15434 = ( wire15425  &  wire4316 ) | ( wire19065  &  wire4327 ) ;
 assign wire15449 = ( wire2587 ) | ( pdata_4_4_  &  wire4305 ) ;
 assign wire15464 = ( wire2585 ) | ( wire18684 ) | ( wire18685 ) | ( wire18686 ) ;
 assign wire15479 = ( wire2574 ) | ( wire18695 ) | ( wire18696 ) | ( wire18697 ) ;
 assign wire15494 = ( wire2561 ) | ( wire18707 ) | ( wire18711 ) ;
 assign wire15509 = ( wire2545 ) | ( wire2546 ) | ( wire18712 ) ;
 assign wire15524 = ( wire2541 ) | ( wire2542 ) | ( wire18714 ) ;
 assign wire15539 = ( wire18724 ) | ( wire18725 ) | ( wire18729 ) ;
 assign wire15554 = ( (~ preset)  &  pdata_12_12_  &  nrq10_4 ) | ( (~ preset)  &  wire15545  &  (~ nrq10_4) ) ;
 assign wire15569 = ( wire2521 ) | ( pdata_3_3_  &  wire4353 ) ;
 assign wire15584 = ( wire2519 ) | ( pdata_14_14_  &  wire4353 ) ;
 assign wire15599 = ( (~ preset)  &  pdata_5_5_  &  nrq14_3 ) | ( (~ preset)  &  wire15590  &  (~ nrq14_3) ) ;
 assign wire15614 = ( (~ preset)  &  pdata_0_0_  &  nrq14_3 ) | ( (~ preset)  &  wire15605  &  (~ nrq14_3) ) ;
 assign wire15629 = ( wire2512 ) | ( wire2513 ) ;
 assign wire15644 = ( wire2510 ) | ( wire2511 ) ;
 assign wire15659 = ( wire2508 ) | ( wire2509 ) ;
 assign wire15674 = ( (~ preset)  &  pdata_3_3_  &  nrq23_3 ) | ( (~ preset)  &  wire15665  &  (~ nrq23_3) ) ;
 assign wire15689 = ( wire15680  &  wire4280 ) | ( wire18176  &  wire19360 ) ;
 assign wire15704 = ( wire2503 ) | ( wire15695  &  wire4280 ) ;
 assign wire15719 = ( wire2500 ) | ( wire2501 ) ;
 assign wire15734 = ( wire2498 ) | ( wire18501  &  wire19368 ) ;
 assign wire15764 = ( (~ preset)  &  wire19091  &  nrq4_2 ) | ( (~ preset)  &  wire15755  &  (~ nrq4_2) ) ;
 assign wire15779 = ( wire15770  &  wire4331 ) | ( wire19060  &  wire4332 ) ;
 assign wire15794 = ( wire2492 ) | ( pdata_3_3_  &  wire4305 ) ;
 assign wire15809 = ( wire18734 ) | ( wire18735 ) | ( wire18739 ) ;
 assign wire15824 = ( wire18746 ) | ( wire18747 ) | ( wire18751 ) ;
 assign wire15839 = ( wire2465 ) | ( wire18759 ) | ( wire18763 ) ;
 assign wire15854 = ( wire2449 ) | ( wire2450 ) | ( wire18764 ) ;
 assign wire15869 = ( wire2445 ) | ( wire2446 ) | ( wire18766 ) ;
 assign wire15884 = ( wire18776 ) | ( wire18777 ) | ( wire18781 ) ;
 assign wire15899 = ( (~ preset)  &  pdata_11_11_  &  nrq10_4 ) | ( (~ preset)  &  wire15890  &  (~ nrq10_4) ) ;
 assign wire15914 = ( wire2425 ) | ( pdata_4_4_  &  wire4353 ) ;
 assign wire15929 = ( wire2423 ) | ( pdata_13_13_  &  wire4353 ) ;
 assign wire15944 = ( (~ preset)  &  pdata_6_6_  &  nrq14_3 ) | ( (~ preset)  &  wire15935  &  (~ nrq14_3) ) ;
 assign wire15959 = ( (~ preset)  &  pdata_15_15_  &  nrq14_3 ) | ( (~ preset)  &  wire15950  &  (~ nrq14_3) ) ;
 assign wire15974 = ( wire2416 ) | ( wire2417 ) ;
 assign wire15989 = ( wire2414 ) | ( wire2415 ) ;
 assign wire16004 = ( wire2412 ) | ( wire2413 ) ;
 assign wire16019 = ( wire2410 ) | ( wire2411 ) ;
 assign wire16034 = ( wire2408 ) | ( wire18176  &  (~ n_n2471)  &  n_n2487 ) | ( wire18176  &  n_n2471  &  (~ n_n2487) ) ;
 assign wire16049 = ( wire16040  &  wire4280 ) | ( wire18176  &  wire19359 ) ;
 assign wire16064 = ( wire2404 ) | ( wire19360  &  wire4308 ) ;
 assign wire16079 = ( wire2402 ) | ( wire18501  &  wire19367 ) ;
 assign wire16094 = ( wire2400 ) | ( wire16928  &  wire19387 ) ;
 assign wire16109 = ( (~ preset)  &  wire19096  &  nrq4_2 ) | ( (~ preset)  &  wire16100  &  (~ nrq4_2) ) ;
 assign wire16904 = ( wire18813 ) | ( wire18814 ) ;
 assign wire16917 = ( wire2374 ) | ( wire18815 ) ;
 assign wire16928 = ( (~ preset)  &  (~ wire16920)  &  nrq7_2  &  wire3720 ) ;
 assign wire16941 = ( wire17396 ) | ( nrq7_2  &  wire3718  &  wire18816 ) ;
 assign wire16956 = ( wire18828 ) | ( wire18829 ) ;
 assign wire16969 = ( wire2354 ) | ( wire18830 ) ;
 assign wire16980 = ( (~ preset)  &  (~ wire16920)  &  wire16972 ) ;
 assign wire16993 = ( (~ preset)  &  wire16985  &  (~ wire18389) ) ;
 assign wire17008 = ( wire2351 ) | ( wire18832 ) ;
 assign wire17021 = ( (~ preset)  &  wire17011 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17032 = ( (~ preset)  &  (~ pdn) ) ;
 assign wire17045 = ( (~ preset)  &  wire17037  &  (~ wire17102) ) | ( (~ preset)  &  (~ wire17102)  &  wire18025 ) ;
 assign wire17058 = ( (~ preset)  &  (~ wire17050)  &  wire17115 ) ;
 assign wire17073 = ( wire2344 ) | ( wire18833 ) ;
 assign wire17086 = ( wire2341 ) | ( wire18834 ) ;
 assign wire17097 = ( (~ preset)  &  (~ pdn)  &  wire17089 ) ;
 assign wire17110 = ( (~ preset)  &  wire17037  &  (~ wire17102) ) ;
 assign wire17123 = ( wire17058 ) | ( nrq7_2  &  wire3750  &  wire18835 ) ;
 assign wire17138 = ( wire2336 ) | ( wire18836 ) ;
 assign wire17151 = ( (~ preset)  &  wire17141 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17162 = ( (~ preset)  &  (~ wire17102)  &  wire17154 ) ;
 assign wire17175 = ( (~ preset)  &  (~ wire17167)  &  nrq7_2  &  wire3727 ) ;
 assign wire17188 = ( wire17240 ) | ( nrq7_2  &  wire3754  &  wire18837 ) ;
 assign wire17203 = ( wire2329 ) | ( wire18838 ) ;
 assign wire17214 = ( wire17279 ) | ( nrq7_2  &  wire3715  &  wire18839 ) ;
 assign wire17227 = ( (~ preset)  &  (~ wire17050)  &  wire17219 ) ;
 assign wire17240 = ( (~ preset)  &  wire17180  &  (~ wire17232) ) ;
 assign wire17253 = ( (~ preset)  &  wire17245  &  (~ nrq7_2) ) | ( (~ preset)  &  wire17245  &  (~ wire3746) ) ;
 assign wire17268 = ( wire2324 ) | ( wire18842 ) ;
 assign wire17279 = ( (~ preset)  &  wire17206  &  (~ wire17271) ) ;
 assign wire17292 = ( wire18384 ) | ( nrq7_2  &  wire3738  &  wire18843 ) ;
 assign wire17305 = ( (~ preset)  &  (~ wire17297)  &  nrq7_2  &  wire3747 ) ;
 assign wire17318 = ( (~ preset)  &  wire17310  &  (~ wire17388) ) ;
 assign wire17333 = ( wire2319 ) | ( wire18845 ) ;
 assign wire17346 = ( (~ preset)  &  wire17336 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17357 = ( (~ preset)  &  (~ wire17271)  &  wire17349 ) ;
 assign wire17370 = ( (~ preset)  &  (~ wire17167)  &  wire17362 ) ;
 assign wire17383 = ( (~ preset)  &  (~ wire17297)  &  wire17375 ) ;
 assign wire17396 = ( (~ preset)  &  wire16933  &  (~ wire17388) ) ;
 assign wire17411 = ( wire18860 ) | ( wire18862 ) ;
 assign wire17422 = ( (~ preset)  &  (~ wire17414)  &  wire17843 ) ;
 assign wire17435 = ( (~ preset)  &  wire17427  &  (~ wire17700) ) | ( (~ preset)  &  wire17518  &  (~ wire17700) ) ;
 assign wire17461 = ( (~ preset)  &  nrq7_2  &  wire17710  &  wire17716 ) ;
 assign wire17476 = ( wire18874 ) | ( wire18875 ) ;
 assign wire17489 = ( (~ preset)  &  wire17479 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17502 = ( wire2280 ) | ( wire18876 ) ;
 assign wire17513 = ( (~ preset)  &  (~ wire17414)  &  wire17505 ) ;
 assign wire17526 = ( (~ preset)  &  wire17518  &  (~ wire17700) ) | ( (~ preset)  &  (~ wire17700)  &  wire17817 ) ;
 assign wire17539 = ( wire2276 ) | ( wire17531  &  wire4466 ) ;
 assign wire17554 = ( (~ preset)  &  ppeaki_7_7_  &  nlbr8_2_e ) | ( (~ preset)  &  wire17544  &  (~ nlbr8_2_e) ) ;
 assign wire17567 = ( wire18889 ) | ( wire18890 ) ;
 assign wire17578 = ( (~ preset)  &  wire17570  &  (~ nrq3_11) ) | ( (~ preset)  &  nen3_5  &  (~ nrq3_11) ) ;
 assign wire17591 = ( (~ preset)  &  wire17583  &  (~ wire17700) ) | ( (~ preset)  &  wire17648  &  (~ wire17700) ) ;
 assign wire17604 = ( wire2246 ) | ( (~ nrq3_11)  &  wire18906 ) ;
 assign wire17619 = ( (~ preset)  &  ppeaki_6_6_  &  nlbr8_2_e ) | ( (~ preset)  &  wire17609  &  (~ nlbr8_2_e) ) ;
 assign wire17632 = ( wire18919 ) | ( wire18920 ) ;
 assign wire17643 = ( (~ preset)  &  wire17570  &  (~ nrq3_11) ) | ( (~ preset)  &  wire17635  &  (~ nrq3_11) ) ;
 assign wire17656 = ( (~ preset)  &  wire17427  &  (~ wire17700) ) | ( (~ preset)  &  wire17648  &  (~ wire17700) ) ;
 assign wire17669 = ( (~ preset)  &  wire18897  &  wire18898  &  wire18901 ) ;
 assign wire17684 = ( (~ preset)  &  ppeaki_5_5_  &  nlbr8_2_e ) | ( (~ preset)  &  wire17674  &  (~ nlbr8_2_e) ) ;
 assign wire17697 = ( wire18932 ) | ( wire18933 ) ;
 assign wire17708 = ( (~ preset)  &  (~ wire17700)  &  wire18142 ) ;
 assign wire17723 = ( (~ preset)  &  ppeaki_4_4_  &  nlbr8_2_e ) | ( (~ preset)  &  wire17713  &  (~ nlbr8_2_e) ) ;
 assign wire17736 = ( wire18945 ) | ( wire18946 ) ;
 assign wire17747 = ( (~ preset)  &  (~ wire17700)  &  wire17739 ) ;
 assign wire17760 = ( wire17752  &  wire4466 ) | ( wire4466  &  nrq7_2  &  wire17710 ) ;
 assign wire17775 = ( wire2187 ) | ( wire18947 ) ;
 assign wire17788 = ( wire2184 ) | ( wire18948 ) ;
 assign wire17799 = ( (~ preset)  &  (~ wire17414)  &  wire17791 ) | ( (~ preset)  &  (~ wire17414)  &  nen2_3 ) ;
 assign wire17812 = ( (~ preset)  &  (~ pdn)  &  nrq3_11 ) ;
 assign wire17825 = ( wire2179 ) | ( (~ preset)  &  (~ wire17700)  &  wire17817 ) ;
 assign wire17840 = ( wire18962 ) | ( wire18963 ) | ( wire18964 ) ;
 assign wire17851 = ( (~ preset)  &  (~ wire17414)  &  wire17843 ) | ( (~ preset)  &  (~ wire17414)  &  wire17791  &  (~ wire17843) ) ;
 assign wire17866 = ( (~ preset)  &  wire17856 ) | ( (~ preset)  &  wire4513 ) ;
 assign wire17879 = ( (~ preset)  &  wire17869 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17892 = ( (~ preset)  &  wire17882 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17905 = ( wire18994 ) | ( wire18995 ) | ( wire18999 ) ;
 assign wire17918 = ( (~ preset)  &  wire17908 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17931 = ( wire2116 ) | ( wire19000 ) ;
 assign wire17944 = ( (~ preset)  &  wire17934 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17957 = ( (~ preset)  &  wire17947 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17970 = ( (~ preset)  &  wire17960 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire17983 = ( wire2107 ) | ( wire19001 ) ;
 assign wire17994 = ( (~ preset)  &  wire17635  &  (~ nrq3_11) ) | ( (~ preset)  &  wire17986  &  (~ nrq3_11) ) ;
 assign wire18007 = ( (~ preset)  &  (~ wire17700)  &  wire17999 ) | ( (~ preset)  &  (~ wire17700)  &  wire18077 ) ;
 assign wire18022 = ( wire2100 ) | ( wire2101 ) ;
 assign wire18033 = ( wire18025  &  wire4458 ) | ( wire4458  &  nrq7_2  &  wire3740 ) ;
 assign wire18048 = ( (~ preset)  &  wire18038 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18059 = ( (~ preset)  &  (~ pdn)  &  wire17414 ) | ( (~ preset)  &  (~ pdn)  &  nrq3_11 ) ;
 assign wire18072 = ( wire2092 ) | ( (~ preset)  &  (~ pdn)  &  wire18064 ) ;
 assign wire18085 = ( (~ preset)  &  wire17583  &  (~ wire17700) ) | ( (~ preset)  &  (~ wire17700)  &  wire18077 ) ;
 assign wire18100 = ( wire2088 ) | ( wire2089 ) ;
 assign wire18111 = ( (~ preset)  &  wire18103  &  (~ wire18168) ) ;
 assign wire18126 = ( (~ preset)  &  wire18116 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18139 = ( wire2084 ) | ( wire2085 ) ;
 assign wire18150 = ( (~ preset)  &  (~ wire17700)  &  wire18142 ) | ( (~ preset)  &  (~ wire17700)  &  wire18220 ) ;
 assign wire18165 = ( wire2080 ) | ( wire2081 ) ;
 assign wire18176 = ( (~ preset)  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire18191 = ( (~ preset)  &  wire18181 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18204 = ( wire2076 ) | ( wire19004 ) ;
 assign wire18215 = ( (~ preset)  &  (~ pdn)  &  wire18207 ) | ( (~ preset)  &  (~ pdn)  &  wire4513 ) ;
 assign wire18228 = ( (~ preset)  &  (~ wire17700)  &  wire17999 ) | ( (~ preset)  &  (~ wire17700)  &  wire18220 ) ;
 assign wire18243 = ( wire2069 ) | ( wire2070 ) ;
 assign wire18254 = ( (~ preset)  &  (~ wire17453)  &  wire18246 ) ;
 assign wire18269 = ( wire19018 ) | ( wire19019 ) ;
 assign wire18282 = ( wire17708 ) | ( wire2050 ) | ( wire2051 ) ;
 assign wire18293 = ( wire2049 ) | ( nrq7_2  &  wire3723  &  wire19022 ) ;
 assign wire18306 = ( (~ preset)  &  wire18298  &  (~ wire18376) ) ;
 assign wire18319 = ( (~ preset)  &  wire18311  &  (~ wire18389) ) | ( (~ preset)  &  (~ wire18389)  &  wire18506 ) ;
 assign wire18334 = ( wire19037 ) | ( wire19038 ) ;
 assign wire18347 = ( wire2028 ) | ( wire19039 ) ;
 assign wire18360 = ( (~ preset)  &  wire18350 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18371 = ( (~ preset)  &  wire18363  &  (~ wire18415) ) | ( (~ preset)  &  wire18285  &  (~ wire18363)  &  (~ wire18415) ) ;
 assign wire18384 = ( (~ preset)  &  wire17284  &  (~ wire18376) ) ;
 assign wire18397 = ( (~ preset)  &  wire18311  &  (~ wire18389) ) ;
 assign wire18412 = ( wire19051 ) | ( wire19052 ) ;
 assign wire18423 = ( (~ preset)  &  wire18363  &  (~ wire18415) ) ;
 assign wire18436 = ( (~ preset)  &  wire18428  &  (~ wire18493) ) ;
 assign wire18449 = ( (~ preset)  &  (~ wire17232)  &  wire18441 ) ;
 assign wire18464 = ( wire19074 ) | ( wire19075 ) ;
 assign wire18475 = ( wire1991 ) | ( wire1992 ) ;
 assign wire18488 = ( (~ preset)  &  (~ wire18415)  &  wire18480 ) ;
 assign wire18501 = ( (~ preset)  &  (~ wire18493)  &  nrq7_2  &  wire3711 ) ;
 assign wire18514 = ( wire18506  &  wire4467 ) | ( wire4467  &  nrq7_2  &  wire3744 ) ;
 assign wire18529 = ( wire19094 ) | ( wire19095 ) ;
 assign wire18542 = ( wire19110 ) | ( wire19111 ) ;
 assign wire18555 = ( (~ preset)  &  pdn  &  wire18545 ) | ( (~ preset)  &  (~ pdn)  &  n_n3081 ) | ( (~ preset)  &  wire18545  &  n_n3081 ) ;
 assign wire18568 = ( wire19124 ) | ( wire19125 ) ;
 assign wire18581 = ( (~ preset)  &  wire18571 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18594 = ( (~ preset)  &  wire18584 ) | ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  wire4242 ) ;
 assign wire18605 = ( wire1936 ) | ( (~ preset)  &  (~ pdn)  &  wire18597 ) ;
 assign wire18618 = ( wire19135 ) | ( wire19136 ) | ( wire18610  &  wire4466 ) ;
 assign wire18633 = ( wire19150 ) | ( wire19151 ) ;
 assign wire18644 = ( wire1915 ) | ( wire19163 ) | ( wire19164 ) ;
 assign wire4305 = ( (~ preset)  &  wire17791  &  (~ wire17843) ) ;
 assign wire4260 = ( wire4199  &  n_n2344  &  wire3775  &  n_n2772 ) ;
 assign wire4269 = ( wire4199  &  n_n2344  &  wire3770  &  n_n2772 ) ;
 assign wire4298 = ( wire4226  &  n_n2772 ) | ( wire4199  &  n_n2333  &  n_n2772 ) ;
 assign wire4392 = ( wire4199  &  n_n2344  &  wire3784  &  n_n2772 ) ;
 assign wire4397 = ( wire4199  &  n_n2772  &  wire4215 ) ;
 assign wire4226 = ( n_n3925  &  wire5514 ) | ( n_n3925  &  (~ wire4202)  &  wire4266 ) ;
 assign wire4352 = ( (~ preset)  &  wire17453  &  (~ wire18246) ) ;
 assign wire4280 = ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire17710) ) | ( (~ preset)  &  (~ wire17711) ) ;
 assign wire4353 = ( (~ preset)  &  wire17102  &  (~ wire17154) ) ;
 assign wire4243 = ( (~ preset)  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire4253 = ( (~ preset)  &  wire18285 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3723) ) ;
 assign wire4354 = ( (~ preset)  &  wire17167  &  (~ wire17362) ) ;
 assign wire4245 = ( (~ preset)  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire4252 = ( (~ preset)  &  wire18506 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3744) ) ;
 assign wire4375 = ( (~ preset)  &  (~ wire17310)  &  wire17388 ) ;
 assign wire19360 = ( n_n2486  &  (~ n_n2471)  &  wire4457 ) | ( (~ n_n2486)  &  (~ n_n2471)  &  (~ wire4457) ) | ( n_n2486  &  n_n2471  &  n_n2487  &  wire4457 ) | ( (~ n_n2486)  &  n_n2471  &  (~ n_n2487)  &  wire4457 ) | ( (~ n_n2486)  &  n_n2471  &  n_n2487  &  (~ wire4457) ) | ( n_n2486  &  n_n2471  &  (~ n_n2487)  &  (~ wire4457) ) ;
 assign wire4340 = ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire17710) ) | ( (~ preset)  &  (~ wire17716) ) ;
 assign wire19390 = ( n_n2475  &  wire19739  &  wire5157 ) | ( (~ n_n2475)  &  (~ wire19739)  &  wire5157 ) | ( n_n2475  &  wire19739  &  wire5158 ) | ( (~ n_n2475)  &  (~ wire19739)  &  wire5158 ) | ( (~ n_n2475)  &  wire19739  &  (~ wire5157)  &  (~ wire5158) ) | ( n_n2475  &  (~ wire19739)  &  (~ wire5157)  &  (~ wire5158) ) ;
 assign wire4308 = ( (~ preset)  &  (~ wire18103)  &  wire18168 ) ;
 assign wire4306 = ( (~ preset)  &  wire18285  &  (~ wire18363) ) ;
 assign wire4317 = ( (~ preset)  &  wire17284 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3738) ) ;
 assign wire4381 = ( (~ preset)  &  (~ wire17284)  &  nrq7_2  &  wire3738 ) ;
 assign wire19368 = ( wire19731  &  wire19474  &  wire4301 ) | ( (~ n_n2473)  &  (~ wire19731)  &  (~ wire4301) ) | ( n_n2473  &  (~ wire19731)  &  wire19474  &  wire4301 ) | ( n_n2473  &  wire19731  &  (~ wire19474)  &  wire4301 ) | ( (~ n_n2473)  &  wire19731  &  (~ wire19474)  &  (~ wire4301) ) | ( n_n2473  &  (~ wire19731)  &  (~ wire19474)  &  (~ wire4301) ) ;
 assign wire19359 = ( n_n2478  &  wire19747  &  wire5164 ) | ( (~ n_n2478)  &  (~ wire19747)  &  wire5164 ) | ( n_n2478  &  wire19747  &  wire5166 ) | ( (~ n_n2478)  &  (~ wire19747)  &  wire5166 ) | ( (~ n_n2478)  &  wire19747  &  (~ wire5164)  &  (~ wire5166) ) | ( n_n2478  &  (~ wire19747)  &  (~ wire5164)  &  (~ wire5166) ) ;
 assign wire4377 = ( (~ preset)  &  (~ wire18311)  &  wire18506 ) ;
 assign wire4277 = ( (~ preset)  &  wire16933 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3718) ) ;
 assign wire4278 = ( (~ preset)  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire19088 = ( (~ ppeaka_6_6_)  &  (~ n_n2449)  &  wire19171 ) | ( (~ ndn_latch24_2)  &  (~ n_n2449)  &  wire19171 ) | ( (~ ppeaka_6_6_)  &  n_n2449  &  (~ wire19171) ) | ( (~ ndn_latch24_2)  &  n_n2449  &  (~ wire19171) ) | ( ppeaka_6_6_  &  ndn_latch24_2  &  n_n2449  &  wire19171 ) | ( ppeaka_6_6_  &  ndn_latch24_2  &  (~ n_n2449)  &  (~ wire19171) ) ;
 assign wire4350 = ( (~ preset)  &  nrq4_2 ) ;
 assign wire19092 = ( (~ ppeaka_10_10_)  &  (~ n_n2445)  &  wire19205 ) | ( (~ ndn_latch24_2)  &  (~ n_n2445)  &  wire19205 ) | ( (~ ppeaka_10_10_)  &  n_n2445  &  (~ wire19205) ) | ( (~ ndn_latch24_2)  &  n_n2445  &  (~ wire19205) ) | ( ppeaka_10_10_  &  ndn_latch24_2  &  n_n2445  &  wire19205 ) | ( ppeaka_10_10_  &  ndn_latch24_2  &  (~ n_n2445)  &  (~ wire19205) ) ;
 assign wire4345 = ( (~ preset)  &  wire17635  &  (~ wire17986) ) ;
 assign wire19103 = ( (~ ppeaka_4_4_)  &  (~ n_n2451)  &  wire19180 ) | ( (~ ndn_latch24_2)  &  (~ n_n2451)  &  wire19180 ) | ( (~ ppeaka_4_4_)  &  n_n2451  &  (~ wire19180) ) | ( (~ ndn_latch24_2)  &  n_n2451  &  (~ wire19180) ) | ( ppeaka_4_4_  &  ndn_latch24_2  &  n_n2451  &  wire19180 ) | ( ppeaka_4_4_  &  ndn_latch24_2  &  (~ n_n2451)  &  (~ wire19180) ) ;
 assign wire4330 = ( (~ preset)  &  wire18025 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3740) ) ;
 assign wire4374 = ( (~ preset)  &  (~ wire18025)  &  nrq7_2  &  wire3740 ) ;
 assign wire19060 = ( (~ ppeaka_9_9_)  &  (~ n_n2446)  &  wire19227 ) | ( (~ ndn_latch24_2)  &  (~ n_n2446)  &  wire19227 ) | ( (~ ppeaka_9_9_)  &  n_n2446  &  (~ wire19227) ) | ( (~ ndn_latch24_2)  &  n_n2446  &  (~ wire19227) ) | ( ppeaka_9_9_  &  ndn_latch24_2  &  n_n2446  &  wire19227 ) | ( ppeaka_9_9_  &  ndn_latch24_2  &  (~ n_n2446)  &  (~ wire19227) ) ;
 assign wire4360 = ( (~ preset)  &  (~ wire17037)  &  wire18025 ) ;
 assign wire19097 = ( (~ ppeaka_3_3_)  &  (~ n_n2452)  &  wire19153 ) | ( (~ ndn_latch24_2)  &  (~ n_n2452)  &  wire19153 ) | ( (~ ppeaka_3_3_)  &  n_n2452  &  (~ wire19153) ) | ( (~ ndn_latch24_2)  &  n_n2452  &  (~ wire19153) ) | ( ppeaka_3_3_  &  ndn_latch24_2  &  n_n2452  &  wire19153 ) | ( ppeaka_3_3_  &  ndn_latch24_2  &  (~ n_n2452)  &  (~ wire19153) ) ;
 assign wire4331 = ( (~ preset)  &  wire17206 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3715) ) ;
 assign wire4332 = ( (~ preset)  &  (~ wire17206)  &  nrq7_2  &  wire3715 ) ;
 assign wire19061 = ( nrq21_7  &  (~ n_n2454)  &  wire4496 ) | ( nrq21_7  &  n_n2454  &  (~ wire4496) ) | ( (~ n_n2454)  &  wire4496  &  (~ wire4451) ) | ( n_n2454  &  (~ wire4496)  &  (~ wire4451) ) | ( (~ nrq21_7)  &  n_n2454  &  wire4496  &  wire4451 ) | ( (~ nrq21_7)  &  (~ n_n2454)  &  (~ wire4496)  &  wire4451 ) ;
 assign wire19091 = ( (~ ppeaka_12_12_)  &  (~ n_n2443)  &  wire19191 ) | ( (~ ndn_latch24_2)  &  (~ n_n2443)  &  wire19191 ) | ( (~ ppeaka_12_12_)  &  n_n2443  &  (~ wire19191) ) | ( (~ ndn_latch24_2)  &  n_n2443  &  (~ wire19191) ) | ( ppeaka_12_12_  &  ndn_latch24_2  &  n_n2443  &  wire19191 ) | ( ppeaka_12_12_  &  ndn_latch24_2  &  (~ n_n2443)  &  (~ wire19191) ) ;
 assign wire4336 = ( (~ preset)  &  wire17245 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3746) ) ;
 assign wire4365 = ( (~ preset)  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire19367 = ( n_n2474  &  wire19514  &  wire4410 ) | ( n_n2474  &  wire19733  &  wire4410 ) | ( wire19514  &  wire19733  &  wire4410 ) | ( (~ n_n2474)  &  (~ wire19514)  &  (~ wire4410) ) | ( (~ n_n2474)  &  (~ wire19733)  &  (~ wire4410) ) | ( (~ wire19514)  &  (~ wire19733)  &  (~ wire4410) ) ;
 assign wire19387 = ( n_n2481  &  wire19729  &  wire5171 ) | ( (~ n_n2481)  &  (~ wire19729)  &  wire5171 ) | ( n_n2481  &  wire19729  &  wire5172 ) | ( (~ n_n2481)  &  (~ wire19729)  &  wire5172 ) | ( (~ n_n2481)  &  wire19729  &  (~ wire5171)  &  (~ wire5172) ) | ( n_n2481  &  (~ wire19729)  &  (~ wire5171)  &  (~ wire5172) ) ;
 assign wire19070 = ( (~ ppeaka_7_7_)  &  (~ n_n2448)  &  wire19221 ) | ( (~ ndn_latch24_2)  &  (~ n_n2448)  &  wire19221 ) | ( (~ ppeaka_7_7_)  &  n_n2448  &  (~ wire19221) ) | ( (~ ndn_latch24_2)  &  n_n2448  &  (~ wire19221) ) | ( ppeaka_7_7_  &  ndn_latch24_2  &  n_n2448  &  wire19221 ) | ( ppeaka_7_7_  &  ndn_latch24_2  &  (~ n_n2448)  &  (~ wire19221) ) ;
 assign wire19096 = ( (~ ppeaka_11_11_)  &  (~ n_n2444)  &  wire19232 ) | ( (~ ndn_latch24_2)  &  (~ n_n2444)  &  wire19232 ) | ( (~ ppeaka_11_11_)  &  n_n2444  &  (~ wire19232) ) | ( (~ ndn_latch24_2)  &  n_n2444  &  (~ wire19232) ) | ( ppeaka_11_11_  &  ndn_latch24_2  &  n_n2444  &  wire19232 ) | ( ppeaka_11_11_  &  ndn_latch24_2  &  (~ n_n2444)  &  (~ wire19232) ) ;
 assign wire19072 = ( (~ ppeaka_8_8_)  &  (~ n_n2447)  &  wire19196 ) | ( (~ ndn_latch24_2)  &  (~ n_n2447)  &  wire19196 ) | ( (~ ppeaka_8_8_)  &  n_n2447  &  (~ wire19196) ) | ( (~ ndn_latch24_2)  &  n_n2447  &  (~ wire19196) ) | ( ppeaka_8_8_  &  ndn_latch24_2  &  n_n2447  &  wire19196 ) | ( ppeaka_8_8_  &  ndn_latch24_2  &  (~ n_n2447)  &  (~ wire19196) ) ;
 assign wire19087 = ( (~ ppeaka_13_13_)  &  (~ n_n2442)  &  wire19215 ) | ( (~ ndn_latch24_2)  &  (~ n_n2442)  &  wire19215 ) | ( (~ ppeaka_13_13_)  &  n_n2442  &  (~ wire19215) ) | ( (~ ndn_latch24_2)  &  n_n2442  &  (~ wire19215) ) | ( ppeaka_13_13_  &  ndn_latch24_2  &  n_n2442  &  wire19215 ) | ( ppeaka_13_13_  &  ndn_latch24_2  &  (~ n_n2442)  &  (~ wire19215) ) ;
 assign wire19082 = ( (~ ppeaka_5_5_)  &  (~ n_n2450)  &  wire19157 ) | ( (~ ndn_latch24_2)  &  (~ n_n2450)  &  wire19157 ) | ( (~ ppeaka_5_5_)  &  n_n2450  &  (~ wire19157) ) | ( (~ ndn_latch24_2)  &  n_n2450  &  (~ wire19157) ) | ( ppeaka_5_5_  &  ndn_latch24_2  &  n_n2450  &  wire19157 ) | ( ppeaka_5_5_  &  ndn_latch24_2  &  (~ n_n2450)  &  (~ wire19157) ) ;
 assign wire19396 = ( n_n2484  &  wire19452  &  wire5190 ) | ( (~ n_n2484)  &  (~ wire19452)  &  wire5190 ) | ( n_n2484  &  wire19452  &  wire17770 ) | ( (~ n_n2484)  &  (~ wire19452)  &  wire17770 ) | ( (~ n_n2484)  &  wire19452  &  (~ wire5190)  &  (~ wire17770) ) | ( n_n2484  &  (~ wire19452)  &  (~ wire5190)  &  (~ wire17770) ) ;
 assign wire4383 = ( (~ preset)  &  (~ wire17999)  &  wire18077 ) ;
 assign wire19073 = ( (~ wire4273)  &  (~ wire17906)  &  wire17913 ) | ( (~ ppeaks_0_0_)  &  wire4273  &  (~ wire17913) ) | ( (~ ppeaks_0_0_)  &  wire17906  &  (~ wire17913) ) | ( (~ wire4273)  &  wire17906  &  (~ wire17913) ) ;
 assign wire4307 = ( (~ preset)  &  (~ wire17180)  &  nrq7_2  &  wire3754 ) ;
 assign wire4325 = ( (~ preset)  &  wire17180 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3754) ) ;
 assign wire19068 = ( (~ ppeaka_14_14_)  &  (~ n_n2441)  &  wire19175 ) | ( (~ ndn_latch24_2)  &  (~ n_n2441)  &  wire19175 ) | ( (~ ppeaka_14_14_)  &  n_n2441  &  (~ wire19175) ) | ( (~ ndn_latch24_2)  &  n_n2441  &  (~ wire19175) ) | ( ppeaka_14_14_  &  ndn_latch24_2  &  n_n2441  &  wire19175 ) | ( ppeaka_14_14_  &  ndn_latch24_2  &  (~ n_n2441)  &  (~ wire19175) ) ;
 assign wire19065 = ( (~ ppeaka_2_2_)  &  (~ n_n2453)  &  wire19167 ) | ( (~ ndn_latch24_2)  &  (~ n_n2453)  &  wire19167 ) | ( (~ ppeaka_2_2_)  &  n_n2453  &  (~ wire19167) ) | ( (~ ndn_latch24_2)  &  n_n2453  &  (~ wire19167) ) | ( ppeaka_2_2_  &  ndn_latch24_2  &  n_n2453  &  wire19167 ) | ( ppeaka_2_2_  &  ndn_latch24_2  &  (~ n_n2453)  &  (~ wire19167) ) ;
 assign wire4357 = ( (~ preset)  &  wire17414  &  (~ wire17505) ) ;
 assign wire1427 = ( ppeaki_14_14_  &  n_n2344 ) | ( ppeaki_10_10_  &  wire4292 ) ;
 assign wire4199 = ( (~ preset)  &  wire18636 ) | ( (~ preset)  &  (~ nrq7_2)  &  wire17582 ) ;
 assign wire4358 = ( (~ preset)  &  (~ wire18142)  &  wire18220 ) ;
 assign wire1342 = ( ppeaki_12_12_  &  n_n2344 ) | ( ppeaki_8_8_  &  wire4292 ) ;
 assign wire1353 = ( ppeaki_13_13_  &  n_n2344 ) | ( ppeaki_9_9_  &  wire4292 ) ;
 assign wire4359 = ( (~ preset)  &  wire17570  &  (~ wire17635) ) ;
 assign wire1412 = ( ppeaki_13_13_  &  wire4292 ) ;
 assign wire1397 = ( ppeaki_12_12_  &  wire4292 ) ;
 assign wire4316 = ( (~ preset)  &  wire17115 ) | ( (~ preset)  &  (~ nrq7_2) ) | ( (~ preset)  &  (~ wire3750) ) ;
 assign wire4327 = ( (~ preset)  &  (~ wire17115)  &  nrq7_2  &  wire3750 ) ;
 assign wire1439 = ( ppeaki_15_15_  &  n_n2344 ) | ( ppeaki_11_11_  &  wire4292 ) ;
 assign wire1368 = ( ppeaki_10_10_  &  n_n2344 ) | ( ppeaki_6_6_  &  wire4292 ) ;
 assign wire4368 = ( (~ preset)  &  wire17427  &  (~ wire17648) ) ;
 assign wire1386 = ( ppeaki_11_11_  &  n_n2344 ) | ( ppeaki_7_7_  &  wire4292 ) ;
 assign wire1411 = ( ppeaki_15_15_  &  wire4292 ) ;
 assign wire1398 = ( ppeaki_8_8_  &  n_n2344 ) | ( ppeaki_4_4_  &  wire4292 ) ;
 assign wire1434 = ( ppeaki_14_14_  &  wire4292 ) ;
 assign wire1413 = ( ppeaki_9_9_  &  n_n2344 ) | ( ppeaki_5_5_  &  wire4292 ) ;
 assign wire4341 = ( (~ preset)  &  nrq4_5  &  wire18795 ) | ( (~ preset)  &  nrq4_5  &  wire18796 ) ;
 assign wire4351 = ( (~ preset)  &  nrq23_3  &  wire18795 ) | ( (~ preset)  &  nrq23_3  &  wire18796 ) ;
 assign wire4369 = ( (~ preset)  &  nrq4_9  &  wire18795 ) | ( (~ preset)  &  nrq4_9  &  wire18796 ) ;
 assign wire4378 = ( (~ preset)  &  ndn_latch12_11  &  wire18795 ) | ( (~ preset)  &  ndn_latch12_11  &  wire18796 ) ;
 assign wire4382 = ( (~ preset)  &  nrq17_3  &  wire18795 ) | ( (~ preset)  &  nrq17_3  &  wire18796 ) ;
 assign wire4467 = ( (~ preset)  &  (~ wire18389) ) ;
 assign wire4458 = ( (~ preset)  &  (~ wire17102) ) ;
 assign nrq21_7 = ( wire17180  &  (~ wire17232) ) ;
 assign nrq13_4 = ( wire17206  &  (~ wire17271) ) ;
 assign wire4300 = ( (~ preset)  &  (~ wire17700) ) ;
 assign ndn7_2 = ( wire18636 ) | ( (~ nrq7_2)  &  wire17582 ) ;
 assign wire4466 = ( (~ preset)  &  (~ wire18636)  &  nrq7_2 ) | ( (~ preset)  &  (~ wire18636)  &  (~ wire17582) ) ;
 assign nen3_5 = ( wire18467 ) | ( nen3_2  &  (~ n_n3925) ) ;
 assign nrq3_11 = ( wire18904 ) | ( wire18900  &  wire18901  &  wire18902 ) ;
 assign nrq8_2 = ( (~ wire18610)  &  n_n2344  &  (~ nsl8_2)  &  nrq7_2 ) ;
 assign nen2_3 = ( preset_0_0_  &  (~ pdn)  &  (~ wire17024) ) | ( (~ pdn)  &  wire17024  &  wire18545 ) ;
 assign wire4235 = ( (~ wire17518)  &  wire17817 ) | ( (~ wire17037)  &  wire18025 ) ;
 assign wire4513 = ( (~ wire5528)  &  (~ wire17599)  &  wire17601 ) | ( (~ wire5528)  &  (~ wire17600)  &  wire17601 ) ;
 assign wire4241 = ( wire17461 ) | ( wire18176 ) | ( wire18798 ) | ( wire18799 ) ;
 assign nrq10_4 = ( (~ wire18168)  &  nrq7_2  &  wire3770  &  wire17710 ) ;
 assign nrq4_14 = ( wire17999  &  (~ wire18220) ) ;
 assign nrq14_8 = ( wire18363  &  (~ wire18415) ) ;
 assign nen3_2 = ( (~ preset_0_0_)  &  (~ pdn)  &  (~ wire17024) ) | ( (~ preset_0_0_)  &  (~ pdn)  &  (~ wire18545) ) | ( (~ pdn)  &  wire17024  &  (~ wire18545) ) ;
 assign n_n2344 = ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) ;
 assign nsl8_2 = ( wire17555 ) | ( wire17556 ) | ( wire17557 ) | ( wire17558 ) ;
 assign nrq7_2 = ( wire17580 ) | ( (~ nsl8_2)  &  wire17564 ) | ( (~ nsl8_2)  &  wire17574 ) ;
 assign nrq1_4 = ( pdn  &  (~ wire17089) ) ;
 assign wire3723 = ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign wire3744 = ( n_n3712  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) ;
 assign wire3738 = ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) ;
 assign wire3718 = ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) ;
 assign n_n3925 = ( pirq_0_0_  &  (~ wire18064) ) | ( wire18064  &  wire18129 ) ;
 assign ndn_latch3_9 = ( wire17635  &  (~ wire17986) ) ;
 assign wire3740 = ( (~ n_n3712)  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) ;
 assign ndn_latch12_11 = ( (~ wire17037)  &  wire18025 ) ;
 assign wire3715 = ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) ;
 assign ndn_latch13_2 = ( (~ wire17206)  &  nrq7_2  &  wire3715 ) ;
 assign ndn_latch24_2 = ( (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire3746 = ( n_n3712  &  n_n3711  &  n_n3714  &  n_n3713 ) ;
 assign wire3747 = ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) ;
 assign nrq23_3 = ( (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire3770 = ( wire17602  &  wire17603 ) | ( wire4471  &  wire17605 ) ;
 assign wire3775 = ( wire17606  &  wire17607 ) | ( wire4471  &  wire17608 ) ;
 assign nrq3_5 = ( (~ wire17570)  &  wire18467 ) | ( (~ wire17570)  &  nen3_2  &  (~ n_n3925) ) ;
 assign nrq14_3 = ( (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign nrq4_9 = ( (~ wire17583)  &  wire17648 ) ;
 assign wire3727 = ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) ;
 assign nrq17_3 = ( (~ wire17284)  &  nrq7_2  &  wire3738 ) ;
 assign wire3711 = ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign nrq15_5 = ( (~ wire17115)  &  nrq7_2  &  wire3750 ) ;
 assign nrq21_5 = ( (~ wire17180)  &  nrq7_2  &  wire3754 ) ;
 assign nrq4_5 = ( (~ wire17518)  &  wire17817 ) ;
 assign nrq4_2 = ( (~ wire17817)  &  (~ wire18467)  &  nen3_2  &  n_n3925 ) ;
 assign wire3750 = ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) ;
 assign wire3754 = ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  n_n3713 ) ;
 assign n_n2333 = ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign n_n3712 = ( ppeaki_2_2_  &  (~ wire17531) ) | ( wire17531  &  wire18012 ) ;
 assign n_n2326 = ( wire4470  &  wire17517 ) | ( wire4468  &  wire17519 ) ;
 assign n_n2314 = ( wire4470  &  wire4483 ) | ( wire17520  &  wire17521 ) ;
 assign n_n2325 = ( wire4471  &  wire17522 ) | ( wire4465  &  wire17523 ) ;
 assign n_n2316 = ( wire4483  &  wire17524 ) | ( wire4459  &  wire17525 ) ;
 assign n_n2318 = ( wire4470  &  wire4480 ) | ( wire4391  &  wire17527 ) ;
 assign n_n2323 = ( wire4472  &  wire17528 ) | ( wire4465  &  wire17529 ) ;
 assign n_n2317 = ( wire4483  &  wire17530 ) | ( wire4459  &  wire17532 ) ;
 assign n_n2315 = ( wire4483  &  wire4472 ) | ( wire17533  &  wire17534 ) ;
 assign n_n2321 = ( wire4480  &  wire17535 ) | ( wire4459  &  wire17536 ) ;
 assign n_n2324 = ( wire4471  &  wire17537 ) | ( wire4465  &  wire17538 ) ;
 assign n_n2320 = ( wire4480  &  wire17540 ) | ( wire4459  &  wire17541 ) ;
 assign n_n2322 = ( wire4470  &  wire17542 ) | ( wire4465  &  wire17543 ) ;
 assign n_n2319 = ( wire4480  &  wire4472 ) | ( wire4391  &  wire17545 ) ;
 assign wire3784 = ( wire4472  &  wire17546 ) | ( wire4468  &  wire17547 ) ;
 assign wire4468 = ( (~ wire17609)  &  wire17674 ) ;
 assign wire4470 = ( ppeaki_4_4_  &  ppeaki_5_5_ ) ;
 assign wire4391 = ( wire17544  &  wire17752 ) ;
 assign wire4483 = ( ppeaki_6_6_  &  ppeaki_7_7_  &  (~ wire17752) ) ;
 assign wire4273 = ( ndn_latch13_2 ) | ( nrq15_5 ) | ( nrq21_5 ) | ( wire17865 ) ;
 assign n_n2453 = ( wire17900 ) | ( ppeaks_2_2_  &  wire4273 ) ;
 assign n_n2452 = ( wire17894 ) | ( ppeaks_3_3_  &  wire4273 ) ;
 assign wire4465 = ( (~ wire17544)  &  wire17609  &  wire17752 ) ;
 assign wire4471 = ( (~ ppeaki_5_5_)  &  (~ ppeaki_7_7_)  &  (~ wire17752) ) ;
 assign wire4459 = ( wire17544  &  (~ wire17674)  &  wire17752 ) ;
 assign wire4480 = ( (~ ppeaki_6_6_)  &  ppeaki_7_7_  &  (~ wire17752) ) ;
 assign wire4472 = ( (~ ppeaki_4_4_)  &  ppeaki_5_5_ ) ;
 assign wire4205 = ( pdn  &  (~ wire17089) ) | ( (~ wire17596)  &  wire4513 ) ;
 assign n_n2772 = ( wire18636 ) | ( wire4205 ) | ( (~ nrq7_2)  &  wire17582 ) ;
 assign wire4234 = ( nrq4_9 ) | ( (~ wire17284)  &  nrq7_2  &  wire3738 ) ;
 assign wire4242 = ( wire4235 ) | ( ndn_latch13_2 ) | ( nrq15_5 ) | ( nrq21_5 ) ;
 assign n_n2443 = ( wire18005 ) | ( ppeaks_12_12_  &  wire4273 ) ;
 assign n_n2449 = ( wire17873 ) | ( ppeaks_6_6_  &  wire4273 ) ;
 assign n_n3711 = ( ppeaki_3_3_  &  (~ wire17531) ) | ( wire17531  &  wire18090 ) ;
 assign n_n2442 = ( wire17998 ) | ( ppeaks_13_13_  &  wire4273 ) ;
 assign n_n2446 = ( wire17949 ) | ( ppeaks_9_9_  &  wire4273 ) ;
 assign n_n2447 = ( wire17955 ) | ( ppeaks_8_8_  &  wire4273 ) ;
 assign n_n2445 = ( wire17941 ) | ( ppeaks_10_10_  &  wire4273 ) ;
 assign n_n2441 = ( wire17991 ) | ( ppeaks_14_14_  &  wire4273 ) ;
 assign n_n2440 = ( wire17984 ) | ( ppeaks_15_15_  &  wire4273 ) ;
 assign n_n2444 = ( wire18013 ) | ( ppeaks_11_11_  &  wire4273 ) ;
 assign n_n2454 = ( wire17920 ) | ( ppeaks_1_1_  &  wire4273 ) ;
 assign n_n2450 = ( wire17880 ) | ( ppeaks_5_5_  &  wire4273 ) ;
 assign n_n2451 = ( wire17887 ) | ( ppeaks_4_4_  &  wire4273 ) ;
 assign n_n2448 = ( wire17963 ) | ( ppeaks_7_7_  &  wire4273 ) ;
 assign n_n3081 = ( preset_0_0_  &  (~ wire17024) ) | ( wire17024  &  wire18545 ) ;
 assign n_n3714 = ( ppeaki_0_0_  &  (~ wire17531) ) | ( wire17531  &  wire18155 ) ;
 assign wire3720 = ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) ;
 assign nlbr8_2_e = ( (~ wire17752)  &  (~ nsl8_2)  &  nrq7_2  &  wire17709 ) ;
 assign wire4265 = ( wire17717 ) | ( wire17718 ) | ( (~ wire18103)  &  wire18168 ) ;
 assign wire4488 = ( wire17037  &  (~ wire17102) ) | ( wire17284  &  (~ wire18376) ) ;
 assign n_n2475 = ( wire17742 ) | ( ppeaks_12_12_  &  wire4265 ) | ( ppeaks_12_12_  &  wire17719 ) ;
 assign n_n3713 = ( ppeaki_1_1_  &  (~ wire17531) ) | ( wire17531  &  wire18233 ) ;
 assign n_n2472 = ( wire17841 ) | ( ppeaks_15_15_  &  wire4265 ) | ( ppeaks_15_15_  &  wire17719 ) ;
 assign wire4292 = ( n_n3712  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) | ( n_n3712  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) | ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) | ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) | ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign n_n2484 = ( wire17768 ) | ( ppeaks_3_3_  &  wire4265 ) | ( ppeaks_3_3_  &  wire17719 ) ;
 assign n_n2474 = ( wire17829 ) | ( ppeaks_13_13_  &  wire4265 ) | ( ppeaks_13_13_  &  wire17719 ) ;
 assign n_n2479 = ( wire17796 ) | ( ppeaks_8_8_  &  wire4265 ) | ( ppeaks_8_8_  &  wire17719 ) ;
 assign n_n2483 = ( wire17774 ) | ( ppeaks_4_4_  &  wire4265 ) | ( ppeaks_4_4_  &  wire17719 ) ;
 assign n_n2485 = ( wire17763 ) | ( ppeaks_2_2_  &  wire4265 ) | ( ppeaks_2_2_  &  wire17719 ) ;
 assign n_n2482 = ( wire17780 ) | ( ppeaks_5_5_  &  wire4265 ) | ( ppeaks_5_5_  &  wire17719 ) ;
 assign n_n2480 = ( wire17792 ) | ( ppeaks_7_7_  &  wire4265 ) | ( ppeaks_7_7_  &  wire17719 ) ;
 assign n_n2486 = ( wire17731 ) | ( ppeaks_1_1_  &  wire4265 ) | ( ppeaks_1_1_  &  wire17719 ) ;
 assign n_n2473 = ( wire17833 ) | ( ppeaks_14_14_  &  wire4265 ) | ( ppeaks_14_14_  &  wire17719 ) ;
 assign n_n2471 = ( ndn_latch24_2 ) | ( nrq17_3 ) | ( wire4265 ) | ( wire17722 ) ;
 assign n_n2487 = ( wire17727 ) | ( ppeaks_0_0_  &  wire4265 ) | ( ppeaks_0_0_  &  wire17719 ) ;
 assign n_n2476 = ( wire17813 ) | ( ppeaks_11_11_  &  wire4265 ) | ( ppeaks_11_11_  &  wire17719 ) ;
 assign n_n2478 = ( wire17801 ) | ( ppeaks_9_9_  &  wire4265 ) | ( ppeaks_9_9_  &  wire17719 ) ;
 assign n_n2477 = ( wire17808 ) | ( ppeaks_10_10_  &  wire4265 ) | ( ppeaks_10_10_  &  wire17719 ) ;
 assign n_n2481 = ( wire17784 ) | ( ppeaks_6_6_  &  wire4265 ) | ( ppeaks_6_6_  &  wire17719 ) ;
 assign wire4024 = ( wire17688 ) | ( wire17689 ) | ( wire17690 ) | ( wire17691 ) ;
 assign wire19749 = ( wire4265  &  wire4457 ) | ( wire4457  &  wire17719 ) | ( wire4457  &  wire17722 ) | ( (~ wire4265)  &  (~ wire4457)  &  (~ wire17719)  &  (~ wire17722) ) ;
 assign wire19466 = ( n_n2486  &  n_n2471  &  n_n2487 ) | ( n_n2486  &  n_n2471  &  wire4457 ) | ( n_n2471  &  n_n2487  &  wire4457 ) | ( n_n2486  &  (~ n_n2471)  &  (~ wire4457) ) ;
 assign wire19739 = ( wire17758 ) | ( (~ ppeaka_12_12_)  &  (~ wire5271)  &  (~ wire5272) ) ;
 assign wire19514 = ( n_n2475  &  wire19739 ) | ( n_n2475  &  wire5157 ) | ( wire19739  &  wire5157 ) | ( n_n2475  &  wire5158 ) | ( wire19739  &  wire5158 ) ;
 assign wire19741 = ( wire5273 ) | ( wire5274 ) | ( (~ ppeaka_11_11_)  &  (~ wire4455) ) ;
 assign wire19531 = ( n_n2477  &  wire19735 ) | ( n_n2477  &  wire19504 ) | ( wire19735  &  wire19504 ) ;
 assign wire4438 = ( n_n2476 ) | ( wire5273 ) | ( wire5274 ) | ( wire5275 ) ;
 assign wire19727 = ( wire17748 ) | ( wire4508  &  (~ wire5288)  &  (~ wire5289) ) ;
 assign wire19456 = ( n_n2483  &  wire19725 ) | ( n_n2483  &  wire19479 ) | ( wire19725  &  wire19479 ) ;
 assign wire4440 = ( n_n2482 ) | ( wire5286 ) | ( wire17748 ) ;
 assign wire19735 = ( (~ wire4455)  &  wire5277 ) | ( wire19743  &  wire4455  &  (~ wire5277) ) | ( (~ wire19743)  &  (~ wire4455)  &  wire17753 ) | ( wire4455  &  (~ wire5277)  &  (~ wire17753) ) ;
 assign wire19504 = ( n_n2478  &  wire19747 ) | ( n_n2478  &  wire5164 ) | ( wire19747  &  wire5164 ) | ( n_n2478  &  wire5166 ) | ( wire19747  &  wire5166 ) ;
 assign wire19725 = ( (~ wire4452)  &  wire5288 ) | ( (~ nrq10_4)  &  (~ wire19749)  &  (~ wire4452) ) | ( nrq10_4  &  wire4452  &  (~ wire5288) ) | ( wire19749  &  wire4452  &  (~ wire5288) ) ;
 assign wire19479 = ( n_n2484  &  wire19452 ) | ( n_n2484  &  wire5190 ) | ( wire19452  &  wire5190 ) | ( n_n2484  &  wire17770 ) | ( wire19452  &  wire17770 ) ;
 assign wire19731 = ( wire5106 ) | ( wire17836 ) ;
 assign wire19474 = ( n_n2474  &  wire19514 ) | ( n_n2474  &  wire19733 ) | ( wire19514  &  wire19733 ) ;
 assign wire4301 = ( n_n2472  &  wire5088 ) | ( n_n2472  &  wire5091 ) | ( n_n2472  &  wire17846 ) | ( (~ n_n2472)  &  (~ wire5088)  &  (~ wire5091)  &  (~ wire17846) ) ;
 assign wire19747 = ( wire5241 ) | ( wire5243 ) | ( (~ nrq10_4)  &  (~ wire19989) ) ;
 assign wire19721 = ( wire5290 ) | ( wire5291 ) | ( (~ ppeaka_2_2_)  &  (~ wire4457) ) ;
 assign wire19452 = ( n_n2485  &  wire19466 ) | ( n_n2485  &  wire19721 ) | ( wire19466  &  wire19721 ) ;
 assign wire19733 = ( (~ wire4453)  &  wire5271 ) | ( (~ wire4453)  &  wire5272 ) | ( wire4453  &  (~ wire5271)  &  (~ wire5272) ) ;
 assign wire19737 = ( (~ wire19989)  &  wire4456 ) | ( wire19989  &  (~ wire4456) ) ;
 assign wire19520 = ( n_n2481  &  wire19729 ) | ( n_n2481  &  wire5171 ) | ( wire19729  &  wire5171 ) | ( n_n2481  &  wire5172 ) | ( wire19729  &  wire5172 ) ;
 assign wire19495 = ( n_n2480  &  wire19520 ) | ( n_n2480  &  (~ wire19989)  &  wire4456 ) | ( wire19520  &  (~ wire19989)  &  wire4456 ) | ( n_n2480  &  wire19989  &  (~ wire4456) ) | ( wire19520  &  wire19989  &  (~ wire4456) ) ;
 assign wire19171 = ( n_n2450  &  wire19157 ) | ( n_n2450  &  wire17928 ) | ( wire19157  &  wire17928 ) ;
 assign wire19221 = ( n_n2449  &  wire19171 ) | ( n_n2449  &  wire17932 ) | ( wire19171  &  wire17932 ) ;
 assign wire19205 = ( n_n2446  &  wire19227 ) | ( n_n2446  &  wire17966 ) | ( wire19227  &  wire17966 ) ;
 assign wire19232 = ( n_n2445  &  wire19205 ) | ( n_n2445  &  wire17969 ) | ( wire19205  &  wire17969 ) ;
 assign wire19157 = ( n_n2451  &  wire19180 ) | ( n_n2451  &  wire17927 ) | ( wire19180  &  wire17927 ) ;
 assign wire19180 = ( n_n2452  &  wire19153 ) | ( n_n2452  &  wire17926 ) | ( wire19153  &  wire17926 ) ;
 assign wire4388 = ( n_n2441  &  (~ n_n2440)  &  wire19175 ) | ( (~ n_n2441)  &  n_n2440  &  (~ wire19175) ) | ( n_n2441  &  (~ n_n2440)  &  wire18017 ) | ( (~ n_n2440)  &  wire19175  &  wire18017 ) | ( (~ n_n2441)  &  n_n2440  &  (~ wire18017) ) | ( n_n2440  &  (~ wire19175)  &  (~ wire18017) ) ;
 assign wire4511 = ( (~ ppeaka_15_15_) ) | ( wire16933 ) | ( (~ nrq7_2) ) | ( (~ wire3718) ) ;
 assign wire19227 = ( n_n2447  &  wire19196 ) | ( n_n2447  &  wire17965 ) | ( wire19196  &  wire17965 ) ;
 assign wire19153 = ( n_n2453  &  wire19167 ) | ( n_n2453  &  wire17925 ) | ( wire19167  &  wire17925 ) ;
 assign wire4496 = ( (~ wire4273)  &  (~ wire17906) ) | ( (~ ppeaks_0_0_)  &  (~ wire17913) ) | ( (~ wire4273)  &  (~ wire17913) ) ;
 assign wire19191 = ( n_n2444  &  wire19232 ) | ( n_n2444  &  wire18014 ) | ( wire19232  &  wire18014 ) ;
 assign wire19215 = ( n_n2443  &  wire19191 ) | ( n_n2443  &  wire18015 ) | ( wire19191  &  wire18015 ) ;
 assign wire4410 = ( n_n2473  &  wire5106 ) | ( n_n2473  &  wire17836 ) | ( (~ n_n2473)  &  (~ wire5106)  &  (~ wire17836) ) ;
 assign wire19729 = ( (~ ppeaka_6_6_)  &  (~ wire19989) ) | ( (~ nrq10_4)  &  (~ wire19989) ) | ( (~ wire19989)  &  wire17785 ) ;
 assign wire19196 = ( n_n2448  &  wire19221 ) | ( n_n2448  &  wire17964 ) | ( wire19221  &  wire17964 ) ;
 assign wire19175 = ( n_n2442  &  wire19215 ) | ( n_n2442  &  wire18016 ) | ( wire19215  &  wire18016 ) ;
 assign wire19743 = ( (~ ppeaka_8_8_)  &  (~ wire19989) ) | ( (~ nrq10_4)  &  (~ wire19989) ) | ( ppeaka_7_7_  &  (~ ppeaka_8_8_)  &  nrq10_4 ) | ( (~ ppeaka_7_7_)  &  ppeaka_8_8_  &  nrq10_4  &  wire19989 ) ;
 assign wire4450 = ( n_n2479 ) | ( wire19743 ) ;
 assign wire19167 = ( nrq21_7  &  n_n2454 ) | ( n_n2454  &  (~ wire4451) ) | ( nrq21_7  &  (~ n_n2454)  &  wire17924 ) | ( (~ n_n2454)  &  (~ wire4451)  &  wire17924 ) | ( (~ nrq21_7)  &  n_n2454  &  wire4451  &  wire17924 ) ;
 assign wire4451 = ( (~ ppeaka_1_1_) ) | ( wire16933 ) | ( (~ nrq7_2) ) | ( (~ wire3718) ) ;
 assign wire4457 = ( (~ ppeaka_1_1_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4507 = ( (~ ppeaka_2_2_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4452 = ( (~ ppeaka_4_4_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4508 = ( (~ ppeaka_5_5_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire19989 = ( wire5283 ) | ( (~ wire5286)  &  (~ wire17748)  &  wire17749 ) ;
 assign wire4453 = ( (~ ppeaka_13_13_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire18861 = ( wire5277 ) | ( (~ ppeaka_8_8_)  &  (~ ppeaka_9_9_)  &  (~ wire19743) ) ;
 assign wire4455 = ( (~ ppeaka_10_10_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4456 = ( (~ ppeaka_7_7_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4509 = ( (~ ppeaka_11_11_) ) | ( (~ nrq7_2) ) | ( (~ wire17710) ) | ( (~ wire17711) ) ;
 assign wire4202 = ( n_n3081 ) | ( (~ wire5528)  &  (~ wire17599) ) | ( (~ wire5528)  &  (~ wire17600) ) ;
 assign wire4204 = ( n_n3712  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) ;
 assign wire4207 = ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) ;
 assign wire4208 = ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) ;
 assign wire4209 = ( n_n3712  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) | ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign wire4211 = ( wire4209 ) | ( n_n2344  &  wire3784 ) ;
 assign wire4212 = ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) ;
 assign wire4215 = ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign wire4266 = ( (~ preset)  &  pdn  &  (~ wire17089) ) ;
 assign wire4219 = ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign wire4303 = ( (~ preset)  &  nrq3_5  &  wire18795 ) | ( (~ preset)  &  nrq3_5  &  wire18796 ) ;
 assign wire4224 = ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  (~ n_n3713) ) ;
 assign wire4225 = ( n_n3712  &  n_n3711  &  n_n3714  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  n_n3714  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  n_n3713 ) | ( n_n3712  &  (~ n_n3711)  &  (~ n_n3714)  &  n_n3713 ) | ( (~ n_n3712)  &  n_n3711  &  n_n3714  &  (~ n_n3713) ) | ( n_n3712  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) | ( (~ n_n3712)  &  n_n3711  &  (~ n_n3714)  &  (~ n_n3713) ) ;
 assign wire4515 = ( wire5520 ) | ( (~ preset)  &  (~ n_n2772) ) | ( (~ preset)  &  wire5522 ) ;
 assign wire1914 = ( (~ preset)  &  wire16920  &  nrq7_2 ) ;
 assign wire1915 = ( nrq7_2  &  wire1935 ) | ( nrq7_2  &  wire19135 ) | ( nrq7_2  &  wire19136 ) ;
 assign wire1918 = ( wire8255  &  wire17240  &  wire18795 ) | ( wire8255  &  wire17240  &  wire18796 ) ;
 assign wire1920 = ( wire6065  &  wire18423  &  wire18795 ) | ( wire6065  &  wire18423  &  wire18796 ) ;
 assign wire1921 = ( wire9410  &  wire18397  &  wire18795 ) | ( wire9410  &  wire18397  &  wire18796 ) ;
 assign wire1922 = ( wire10970  &  wire17279  &  wire18795 ) | ( wire10970  &  wire17279  &  wire18796 ) ;
 assign wire1923 = ( ppeaks_7_7_  &  wire4241  &  wire18795 ) | ( ppeaks_7_7_  &  wire4241  &  wire18796 ) ;
 assign wire1926 = ( (~ preset)  &  paddress_7_7_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire1927 = ( wire12905  &  wire17058  &  wire18795 ) | ( wire12905  &  wire17058  &  wire18796 ) ;
 assign wire1928 = ( wire11075  &  n_n3925  &  wire4303 ) ;
 assign wire1929 = ( ppeaka_7_7_  &  wire2391 ) | ( ppeaka_7_7_  &  wire2392 ) ;
 assign wire1930 = ( ppeakp_7_7_  &  wire2394 ) | ( ppeakp_7_7_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire1935 = ( wire18610  &  wire4466 ) ;
 assign wire1936 = ( (~ preset)  &  wire18900  &  wire18901  &  wire19126 ) ;
 assign wire1944 = ( wire7625  &  wire17240  &  wire18795 ) | ( wire7625  &  wire17240  &  wire18796 ) ;
 assign wire1946 = ( wire6740  &  wire18423  &  wire18795 ) | ( wire6740  &  wire18423  &  wire18796 ) ;
 assign wire1947 = ( wire7475  &  wire18397  &  wire18795 ) | ( wire7475  &  wire18397  &  wire18796 ) ;
 assign wire1948 = ( wire11690  &  wire17279  &  wire18795 ) | ( wire11690  &  wire17279  &  wire18796 ) ;
 assign wire1949 = ( ppeaks_6_6_  &  wire4241  &  wire18795 ) | ( ppeaks_6_6_  &  wire4241  &  wire18796 ) ;
 assign wire1952 = ( (~ preset)  &  paddress_6_6_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire1953 = ( wire13865  &  wire17058  &  wire18795 ) | ( wire13865  &  wire17058  &  wire18796 ) ;
 assign wire1954 = ( wire9950  &  n_n3925  &  wire4303 ) ;
 assign wire1955 = ( ppeaka_6_6_  &  wire2391 ) | ( ppeaka_6_6_  &  wire2392 ) ;
 assign wire1956 = ( ppeakp_6_6_  &  wire2394 ) | ( ppeakp_6_6_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire1961 = ( wire6995  &  wire17240  &  wire18795 ) | ( wire6995  &  wire17240  &  wire18796 ) ;
 assign wire1963 = ( wire4670  &  wire18423  &  wire18795 ) | ( wire4670  &  wire18423  &  wire18796 ) ;
 assign wire1964 = ( wire8105  &  wire18397  &  wire18795 ) | ( wire8105  &  wire18397  &  wire18796 ) ;
 assign wire1965 = ( wire11465  &  wire17279  &  wire18795 ) | ( wire11465  &  wire17279  &  wire18796 ) ;
 assign wire1966 = ( ppeaks_5_5_  &  wire4241  &  wire18795 ) | ( ppeaks_5_5_  &  wire4241  &  wire18796 ) ;
 assign wire1969 = ( (~ preset)  &  paddress_5_5_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire1970 = ( wire13505  &  wire17058  &  wire18795 ) | ( wire13505  &  wire17058  &  wire18796 ) ;
 assign wire1971 = ( wire10220  &  n_n3925  &  wire4303 ) ;
 assign wire1972 = ( ppeaka_5_5_  &  wire2391 ) | ( ppeaka_5_5_  &  wire2392 ) ;
 assign wire1973 = ( ppeakp_5_5_  &  wire2394 ) | ( ppeakp_5_5_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire1976 = ( wire12245  &  wire17240  &  wire18795 ) | ( wire12245  &  wire17240  &  wire18796 ) ;
 assign wire1978 = ( wire5375  &  wire18423  &  wire18795 ) | ( wire5375  &  wire18423  &  wire18796 ) ;
 assign wire1979 = ( wire6170  &  wire18397  &  wire18795 ) | ( wire6170  &  wire18397  &  wire18796 ) ;
 assign wire1980 = ( wire5615  &  wire17279  &  wire18795 ) | ( wire5615  &  wire17279  &  wire18796 ) ;
 assign wire1981 = ( ppeaks_4_4_  &  wire4241  &  wire18795 ) | ( ppeaks_4_4_  &  wire4241  &  wire18796 ) ;
 assign wire1984 = ( (~ preset)  &  paddress_4_4_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire1985 = ( wire14675  &  wire17058  &  wire18795 ) | ( wire14675  &  wire17058  &  wire18796 ) ;
 assign wire1986 = ( wire10505  &  n_n3925  &  wire4303 ) ;
 assign wire1987 = ( ppeaka_4_4_  &  wire2391 ) | ( ppeaka_4_4_  &  wire2392 ) ;
 assign wire1988 = ( ppeakp_4_4_  &  wire2394 ) | ( ppeakp_4_4_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire1991 = ( (~ wire18467)  &  nen3_2  &  n_n3925  &  wire19076 ) ;
 assign wire1992 = ( wire17032  &  wire18467 ) | ( wire17032  &  nen3_2  &  (~ n_n3925) ) ;
 assign wire1995 = ( wire12455  &  wire17240  &  wire18795 ) | ( wire12455  &  wire17240  &  wire18796 ) ;
 assign wire1997 = ( wire9995  &  wire18423  &  wire18795 ) | ( wire9995  &  wire18423  &  wire18796 ) ;
 assign wire1998 = ( wire6845  &  wire18397  &  wire18795 ) | ( wire6845  &  wire18397  &  wire18796 ) ;
 assign wire1999 = ( wire4910  &  wire17279  &  wire18795 ) | ( wire4910  &  wire17279  &  wire18796 ) ;
 assign wire2000 = ( ppeaks_3_3_  &  wire4241  &  wire18795 ) | ( ppeaks_3_3_  &  wire4241  &  wire18796 ) ;
 assign wire2003 = ( (~ preset)  &  paddress_3_3_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2004 = ( wire14255  &  wire17058  &  wire18795 ) | ( wire14255  &  wire17058  &  wire18796 ) ;
 assign wire2005 = ( wire10790  &  n_n3925  &  wire4303 ) ;
 assign wire2006 = ( ppeaka_3_3_  &  wire2391 ) | ( ppeaka_3_3_  &  wire2392 ) ;
 assign wire2007 = ( ppeakp_3_3_  &  wire2394 ) | ( ppeakp_3_3_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2010 = ( wire12680  &  wire17240  &  wire18795 ) | ( wire12680  &  wire17240  &  wire18796 ) ;
 assign wire2012 = ( wire9725  &  wire18423  &  wire18795 ) | ( wire9725  &  wire18423  &  wire18796 ) ;
 assign wire2013 = ( wire4760  &  wire18397  &  wire18795 ) | ( wire4760  &  wire18397  &  wire18796 ) ;
 assign wire2014 = ( wire6980  &  wire17279  &  wire18795 ) | ( wire6980  &  wire17279  &  wire18796 ) ;
 assign wire2015 = ( ppeaks_2_2_  &  wire4241  &  wire18795 ) | ( ppeaks_2_2_  &  wire4241  &  wire18796 ) ;
 assign wire2018 = ( (~ preset)  &  paddress_2_2_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2019 = ( wire15425  &  wire17058  &  wire18795 ) | ( wire15425  &  wire17058  &  wire18796 ) ;
 assign wire2020 = ( wire11060  &  n_n3925  &  wire4303 ) ;
 assign wire2021 = ( ppeaka_2_2_  &  wire2391 ) | ( ppeaka_2_2_  &  wire2392 ) ;
 assign wire2022 = ( ppeakp_2_2_  &  wire2394 ) | ( ppeakp_2_2_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2028 = ( (~ preset)  &  wire18337  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2029 = ( (~ preset)  &  ppeaka_0_0_  &  wire4234 ) ;
 assign wire2032 = ( wire12920  &  wire17240  &  wire18795 ) | ( wire12920  &  wire17240  &  wire18796 ) ;
 assign wire2034 = ( wire9290  &  wire18423  &  wire18795 ) | ( wire9290  &  wire18423  &  wire18796 ) ;
 assign wire2035 = ( wire10310  &  wire18397  &  wire18795 ) | ( wire10310  &  wire18397  &  wire18796 ) ;
 assign wire2036 = ( wire6305  &  wire17279  &  wire18795 ) | ( wire6305  &  wire17279  &  wire18796 ) ;
 assign wire2037 = ( ppeaks_1_1_  &  wire4241  &  wire18795 ) | ( ppeaks_1_1_  &  wire4241  &  wire18796 ) ;
 assign wire2040 = ( (~ preset)  &  paddress_1_1_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2041 = ( wire12005  &  wire17058  &  wire18795 ) | ( wire12005  &  wire17058  &  wire18796 ) ;
 assign wire2042 = ( wire11315  &  n_n3925  &  wire4303 ) ;
 assign wire2043 = ( ppeaka_1_1_  &  wire2391 ) | ( ppeaka_1_1_  &  wire2392 ) ;
 assign wire2044 = ( ppeakp_1_1_  &  wire2394 ) | ( ppeakp_1_1_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2045 = ( (~ preset)  &  nrq4_14  &  wire18795 ) | ( (~ preset)  &  nrq4_14  &  wire18796 ) ;
 assign wire2049 = ( (~ preset)  &  wire18285  &  (~ wire18415) ) ;
 assign wire2050 = ( (~ preset)  &  piack_0_0_  &  wire17739 ) ;
 assign wire2051 = ( (~ preset)  &  piack_0_0_  &  (~ wire17700) ) ;
 assign wire2055 = ( wire13175  &  wire17240  &  wire18795 ) | ( wire13175  &  wire17240  &  wire18796 ) ;
 assign wire2057 = ( wire8630  &  wire18423  &  wire18795 ) | ( wire8630  &  wire18423  &  wire18796 ) ;
 assign wire2058 = ( wire10025  &  wire18397  &  wire18795 ) | ( wire10025  &  wire18397  &  wire18796 ) ;
 assign wire2059 = ( wire8240  &  wire17279  &  wire18795 ) | ( wire8240  &  wire17279  &  wire18796 ) ;
 assign wire2060 = ( ppeaks_0_0_  &  wire4241  &  wire18795 ) | ( ppeaks_0_0_  &  wire4241  &  wire18796 ) ;
 assign wire2063 = ( (~ preset)  &  paddress_0_0_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2064 = ( wire12890  &  wire17058  &  wire18795 ) | ( wire12890  &  wire17058  &  wire18796 ) ;
 assign wire2065 = ( wire11555  &  n_n3925  &  wire4303 ) ;
 assign wire2066 = ( ppeaka_0_0_  &  wire2391 ) | ( ppeaka_0_0_  &  wire2392 ) ;
 assign wire2067 = ( ppeakp_0_0_  &  wire2394 ) | ( ppeakp_0_0_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2068 = ( wire17422  &  wire18795 ) | ( wire17422  &  wire18796 ) ;
 assign wire2069 = ( (~ preset)  &  wire17531  &  wire18233 ) | ( (~ preset)  &  wire18233  &  (~ nrq7_2) ) ;
 assign wire2070 = ( (~ preset)  &  ppeaki_1_1_  &  (~ wire17531)  &  nrq7_2 ) ;
 assign wire2076 = ( (~ preset)  &  wire18194  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2077 = ( (~ preset)  &  ppeaka_11_11_  &  wire4234 ) ;
 assign wire2080 = ( (~ preset)  &  wire17531  &  wire18155 ) | ( (~ preset)  &  wire18155  &  (~ nrq7_2) ) ;
 assign wire2081 = ( (~ preset)  &  ppeaki_0_0_  &  (~ wire17531)  &  nrq7_2 ) ;
 assign wire2084 = ( wire18467  &  wire19003 ) | ( (~ nen3_2)  &  wire19003 ) | ( nen3_2  &  (~ n_n3925)  &  wire19003 ) ;
 assign wire2085 = ( (~ preset)  &  (~ wire18467)  &  nen3_2  &  n_n3925 ) ;
 assign wire2088 = ( (~ preset)  &  wire17531  &  wire18090 ) | ( (~ preset)  &  wire18090  &  (~ nrq7_2) ) ;
 assign wire2089 = ( (~ preset)  &  ppeaki_3_3_  &  (~ wire17531)  &  nrq7_2 ) ;
 assign wire2092 = ( wire17032  &  (~ wire18467)  &  nen3_2  &  n_n3925 ) ;
 assign wire2100 = ( (~ preset)  &  wire17531  &  wire18012 ) | ( (~ preset)  &  wire18012  &  (~ nrq7_2) ) ;
 assign wire2101 = ( (~ preset)  &  ppeaki_2_2_  &  (~ wire17531)  &  nrq7_2 ) ;
 assign wire2107 = ( (~ preset)  &  wire17973  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2108 = ( (~ preset)  &  ppeaka_12_12_  &  wire4234 ) ;
 assign wire2116 = ( (~ preset)  &  wire17921  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2117 = ( (~ preset)  &  ppeaka_10_10_  &  wire4234 ) ;
 assign wire2179 = ( (~ wire18467)  &  wire4300  &  nen3_2  &  n_n3925 ) ;
 assign wire2184 = ( (~ preset)  &  wire17778  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2185 = ( (~ preset)  &  ppeaka_14_14_  &  wire4234 ) ;
 assign wire2187 = ( (~ preset)  &  wire17765  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2188 = ( (~ preset)  &  ppeaka_9_9_  &  wire4234 ) ;
 assign wire2193 = ( wire10985  &  wire17240  &  wire18795 ) | ( wire10985  &  wire17240  &  wire18796 ) ;
 assign wire2195 = ( wire6080  &  wire18423  &  wire18795 ) | ( wire6080  &  wire18423  &  wire18796 ) ;
 assign wire2196 = ( wire5480  &  wire18397  &  wire18795 ) | ( wire5480  &  wire18397  &  wire18796 ) ;
 assign wire2197 = ( wire12650  &  wire17279  &  wire18795 ) | ( wire12650  &  wire17279  &  wire18796 ) ;
 assign wire2198 = ( ppeaks_14_14_  &  wire4241  &  wire18795 ) | ( ppeaks_14_14_  &  wire4241  &  wire18796 ) ;
 assign wire2201 = ( (~ preset)  &  paddress_14_14_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2202 = ( wire14270  &  wire17058  &  wire18795 ) | ( wire14270  &  wire17058  &  wire18796 ) ;
 assign wire2203 = ( wire12260  &  n_n3925  &  wire4303 ) ;
 assign wire2204 = ( ppeaka_14_14_  &  wire2391 ) | ( ppeaka_14_14_  &  wire2392 ) ;
 assign wire2205 = ( ppeakp_14_14_  &  wire2394 ) | ( ppeakp_14_14_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2210 = ( wire6320  &  wire17240  &  wire18795 ) | ( wire6320  &  wire17240  &  wire18796 ) ;
 assign wire2212 = ( wire6755  &  wire18423  &  wire18795 ) | ( wire6755  &  wire18423  &  wire18796 ) ;
 assign wire2213 = ( wire8765  &  wire18397  &  wire18795 ) | ( wire8765  &  wire18397  &  wire18796 ) ;
 assign wire2214 = ( wire12425  &  wire17279  &  wire18795 ) | ( wire12425  &  wire17279  &  wire18796 ) ;
 assign wire2215 = ( ppeaks_15_15_  &  wire4241  &  wire18795 ) | ( ppeaks_15_15_  &  wire4241  &  wire18796 ) ;
 assign wire2218 = ( (~ preset)  &  paddress_15_15_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2219 = ( wire13880  &  wire17058  &  wire18795 ) | ( wire13880  &  wire17058  &  wire18796 ) ;
 assign wire2220 = ( wire12470  &  n_n3925  &  wire4303 ) ;
 assign wire2221 = ( ppeaka_15_15_  &  wire2391 ) | ( ppeaka_15_15_  &  wire2392 ) ;
 assign wire2222 = ( ppeakp_15_15_  &  wire2394 ) | ( ppeakp_15_15_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2231 = ( wire10415  &  wire17240  &  wire18795 ) | ( wire10415  &  wire17240  &  wire18796 ) ;
 assign wire2233 = ( wire10010  &  wire18423  &  wire18795 ) | ( wire10010  &  wire18423  &  wire18796 ) ;
 assign wire2234 = ( wire6860  &  wire18397  &  wire18795 ) | ( wire6860  &  wire18397  &  wire18796 ) ;
 assign wire2235 = ( wire14660  &  wire17279  &  wire18795 ) | ( wire14660  &  wire17279  &  wire18796 ) ;
 assign wire2236 = ( ppeaks_12_12_  &  wire4241  &  wire18795 ) | ( ppeaks_12_12_  &  wire4241  &  wire18796 ) ;
 assign wire2239 = ( (~ preset)  &  paddress_12_12_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2240 = ( wire15065  &  wire17058  &  wire18795 ) | ( wire15065  &  wire17058  &  wire18796 ) ;
 assign wire2241 = ( wire12050  &  n_n3925  &  wire4303 ) ;
 assign wire2242 = ( ppeaka_12_12_  &  wire2391 ) | ( ppeaka_12_12_  &  wire2392 ) ;
 assign wire2243 = ( ppeakp_12_12_  &  wire2394 ) | ( ppeakp_12_12_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2246 = ( (~ wire18897)  &  wire18905 ) | ( (~ wire18898)  &  wire18905 ) | ( (~ wire18901)  &  wire18905 ) ;
 assign wire2255 = ( wire17986  &  wire5528 ) | ( wire17986  &  wire17599  &  wire17600 ) ;
 assign wire2260 = ( wire10700  &  wire17240  &  wire18795 ) | ( wire10700  &  wire17240  &  wire18796 ) ;
 assign wire2262 = ( wire9740  &  wire18423  &  wire18795 ) | ( wire9740  &  wire18423  &  wire18796 ) ;
 assign wire2263 = ( wire4775  &  wire18397  &  wire18795 ) | ( wire4775  &  wire18397  &  wire18796 ) ;
 assign wire2264 = ( wire14240  &  wire17279  &  wire18795 ) | ( wire14240  &  wire17279  &  wire18796 ) ;
 assign wire2265 = ( ppeaks_13_13_  &  wire4241  &  wire18795 ) | ( ppeaks_13_13_  &  wire4241  &  wire18796 ) ;
 assign wire2268 = ( (~ preset)  &  paddress_13_13_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2269 = ( wire14690  &  wire17058  &  wire18795 ) | ( wire14690  &  wire17058  &  wire18796 ) ;
 assign wire2270 = ( wire12170  &  n_n3925  &  wire4303 ) ;
 assign wire2271 = ( ppeaka_13_13_  &  wire2391 ) | ( ppeaka_13_13_  &  wire2392 ) ;
 assign wire2272 = ( ppeakp_13_13_  &  wire2394 ) | ( ppeakp_13_13_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2276 = ( (~ preset)  &  (~ wire18636)  &  nrq7_2 ) ;
 assign wire2280 = ( (~ preset)  &  wire17492  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2281 = ( (~ preset)  &  ppeaka_13_13_  &  wire4234 ) ;
 assign wire2286 = ( wire9860  &  wire17240  &  wire18795 ) | ( wire9860  &  wire17240  &  wire18796 ) ;
 assign wire2288 = ( wire9305  &  wire18423  &  wire18795 ) | ( wire9305  &  wire18423  &  wire18796 ) ;
 assign wire2289 = ( wire9770  &  wire18397  &  wire18795 ) | ( wire9770  &  wire18397  &  wire18796 ) ;
 assign wire2290 = ( wire13850  &  wire17279  &  wire18795 ) | ( wire13850  &  wire17279  &  wire18796 ) ;
 assign wire2291 = ( ppeaks_10_10_  &  wire4241  &  wire18795 ) | ( ppeaks_10_10_  &  wire4241  &  wire18796 ) ;
 assign wire2294 = ( (~ preset)  &  paddress_10_10_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2295 = ( wire12665  &  wire17058  &  wire18795 ) | ( wire12665  &  wire17058  &  wire18796 ) ;
 assign wire2296 = ( wire11795  &  n_n3925  &  wire4303 ) ;
 assign wire2297 = ( ppeaka_10_10_  &  wire2391 ) | ( ppeaka_10_10_  &  wire2392 ) ;
 assign wire2298 = ( ppeakp_10_10_  &  wire2394 ) | ( ppeakp_10_10_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2303 = ( wire10130  &  wire17240  &  wire18795 ) | ( wire10130  &  wire17240  &  wire18796 ) ;
 assign wire2305 = ( wire8645  &  wire18423  &  wire18795 ) | ( wire8645  &  wire18423  &  wire18796 ) ;
 assign wire2306 = ( wire10595  &  wire18397  &  wire18795 ) | ( wire10595  &  wire18397  &  wire18796 ) ;
 assign wire2307 = ( wire13490  &  wire17279  &  wire18795 ) | ( wire13490  &  wire17279  &  wire18796 ) ;
 assign wire2308 = ( ppeaks_11_11_  &  wire4241  &  wire18795 ) | ( ppeaks_11_11_  &  wire4241  &  wire18796 ) ;
 assign wire2311 = ( (~ preset)  &  paddress_11_11_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2312 = ( wire12125  &  wire17058  &  wire18795 ) | ( wire12125  &  wire17058  &  wire18796 ) ;
 assign wire2313 = ( wire11915  &  n_n3925  &  wire4303 ) ;
 assign wire2314 = ( ppeaka_11_11_  &  wire2391 ) | ( ppeaka_11_11_  &  wire2392 ) ;
 assign wire2315 = ( ppeakp_11_11_  &  wire2394 ) | ( ppeakp_11_11_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2319 = ( (~ preset)  &  wire17323  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2320 = ( (~ preset)  &  ppeaka_2_2_  &  wire4234 ) ;
 assign wire2324 = ( (~ preset)  &  wire17258  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2325 = ( (~ preset)  &  ppeaka_1_1_  &  wire4234 ) ;
 assign wire2329 = ( (~ preset)  &  wire17193  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2330 = ( (~ preset)  &  ppeaka_4_4_  &  wire4234 ) ;
 assign wire2336 = ( (~ preset)  &  wire17128  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2337 = ( (~ preset)  &  ppeaka_3_3_  &  wire4234 ) ;
 assign wire2341 = ( (~ preset)  &  wire17076  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2342 = ( (~ preset)  &  ppeaka_15_15_  &  wire4234 ) ;
 assign wire2344 = ( (~ preset)  &  wire17063  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2345 = ( (~ preset)  &  ppeaka_6_6_  &  wire4234 ) ;
 assign wire2351 = ( (~ preset)  &  wire16998  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2352 = ( (~ preset)  &  ppeaka_5_5_  &  wire4234 ) ;
 assign wire2354 = ( (~ preset)  &  wire16959  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2355 = ( (~ preset)  &  ppeaka_8_8_  &  wire4234 ) ;
 assign wire2358 = ( wire9590  &  wire17240  &  wire18795 ) | ( wire9590  &  wire17240  &  wire18796 ) ;
 assign wire2360 = ( wire7370  &  wire18423  &  wire18795 ) | ( wire7370  &  wire18423  &  wire18796 ) ;
 assign wire2361 = ( wire10040  &  wire18397  &  wire18795 ) | ( wire10040  &  wire18397  &  wire18796 ) ;
 assign wire2362 = ( wire15770  &  wire17279  &  wire18795 ) | ( wire15770  &  wire17279  &  wire18796 ) ;
 assign wire2363 = ( ppeaks_9_9_  &  wire4241  &  wire18795 ) | ( ppeaks_9_9_  &  wire4241  &  wire18796 ) ;
 assign wire2366 = ( (~ preset)  &  paddress_9_9_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2367 = ( wire12440  &  wire17058  &  wire18795 ) | ( wire12440  &  wire17058  &  wire18796 ) ;
 assign wire2368 = ( wire11570  &  n_n3925  &  wire4303 ) ;
 assign wire2369 = ( ppeaka_9_9_  &  wire2391 ) | ( ppeaka_9_9_  &  wire2392 ) ;
 assign wire2370 = ( ppeakp_9_9_  &  wire2394 ) | ( ppeakp_9_9_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2374 = ( (~ preset)  &  wire16907  &  (~ wire4234)  &  (~ wire4242) ) ;
 assign wire2375 = ( (~ preset)  &  ppeaka_7_7_  &  wire4234 ) ;
 assign wire2378 = ( wire8915  &  wire17240  &  wire18795 ) | ( wire8915  &  wire17240  &  wire18796 ) ;
 assign wire2380 = ( wire8000  &  wire18423  &  wire18795 ) | ( wire8000  &  wire18423  &  wire18796 ) ;
 assign wire2381 = ( wire8750  &  wire18397  &  wire18795 ) | ( wire8750  &  wire18397  &  wire18796 ) ;
 assign wire2382 = ( wire11225  &  wire17279  &  wire18795 ) | ( wire11225  &  wire17279  &  wire18796 ) ;
 assign wire2383 = ( ppeaks_8_8_  &  wire4241  &  wire18795 ) | ( ppeaks_8_8_  &  wire4241  &  wire18796 ) ;
 assign wire2386 = ( (~ preset)  &  paddress_8_8_  &  (~ wire18795)  &  (~ wire18796) ) ;
 assign wire2387 = ( wire13160  &  wire17058  &  wire18795 ) | ( wire13160  &  wire17058  &  wire18796 ) ;
 assign wire2388 = ( wire11330  &  n_n3925  &  wire4303 ) ;
 assign wire2389 = ( ppeaka_8_8_  &  wire2391 ) | ( ppeaka_8_8_  &  wire2392 ) ;
 assign wire2390 = ( ppeakp_8_8_  &  wire2394 ) | ( ppeakp_8_8_  &  (~ n_n3925)  &  wire4303 ) ;
 assign wire2391 = ( (~ preset)  &  nrq14_3  &  wire18795 ) | ( (~ preset)  &  nrq14_3  &  wire18796 ) ;
 assign wire2392 = ( wire17175  &  wire18795 ) | ( wire17175  &  wire18796 ) ;
 assign wire2394 = ( wire17110  &  wire18795 ) | ( wire17110  &  wire18796 ) ;
 assign wire2400 = ( (~ preset)  &  wire16085  &  (~ nrq7_2) ) | ( (~ preset)  &  wire16085  &  (~ wire17714) ) ;
 assign wire2402 = ( (~ preset)  &  wire16070  &  (~ nrq7_2) ) | ( (~ preset)  &  wire16070  &  (~ wire17712) ) ;
 assign wire2404 = ( (~ preset)  &  wire16055  &  wire18103 ) | ( (~ preset)  &  wire16055  &  (~ wire18168) ) ;
 assign wire2408 = ( wire16025  &  wire4280 ) ;
 assign wire2410 = ( (~ preset)  &  wire16010  &  (~ nrq7_2) ) | ( (~ preset)  &  wire16010  &  (~ wire17715) ) ;
 assign wire2411 = ( (~ preset)  &  pdata_9_9_  &  nrq7_2  &  wire17715 ) ;
 assign wire2412 = ( (~ preset)  &  wire15995  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15995  &  (~ wire17715) ) ;
 assign wire2413 = ( (~ preset)  &  pdata_0_0_  &  nrq7_2  &  wire17715 ) ;
 assign wire2414 = ( (~ preset)  &  wire15980  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15980  &  (~ wire17714) ) ;
 assign wire2415 = ( (~ preset)  &  pdata_7_7_  &  nrq7_2  &  wire17714 ) ;
 assign wire2416 = ( (~ preset)  &  wire15965  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15965  &  (~ wire17712) ) ;
 assign wire2417 = ( (~ preset)  &  pdata_14_14_  &  nrq7_2  &  wire17712 ) ;
 assign wire2423 = ( (~ preset)  &  wire15920  &  (~ wire17102) ) | ( (~ preset)  &  wire15920  &  wire17154 ) ;
 assign wire2425 = ( (~ preset)  &  wire15905  &  (~ wire17102) ) | ( (~ preset)  &  wire15905  &  wire17154 ) ;
 assign wire2428 = ( wire9860  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire2429 = ( wire10205  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire2430 = ( wire12665  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire2431 = ( wire13850  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2432 = ( wire10400  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2433 = ( wire6155  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire2434 = ( wire8135  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire2435 = ( wire14585  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire2436 = ( wire5450  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire2437 = ( wire8060  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire2438 = ( wire8810  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2440 = ( wire12860  &  wire4226  &  n_n2772 ) ;
 assign wire2441 = ( wire4700  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2443 = ( ppeaks_10_10_  &  wire17660 ) | ( ppeaks_10_10_  &  wire17662 ) ;
 assign wire2445 = ( wire15665  &  wire4199  &  wire3744 ) ;
 assign wire2446 = ( wire15860  &  wire4515 ) | ( wire15860  &  wire17649 ) | ( wire15860  &  wire17650 ) ;
 assign wire2447 = ( wire13130  &  n_n3925  &  wire5513 ) | ( wire13130  &  n_n3925  &  wire5514 ) ;
 assign wire2449 = ( wire9980  &  wire4199  &  wire3744 ) ;
 assign wire2450 = ( wire15845  &  wire4515 ) | ( wire15845  &  wire17649 ) | ( wire15845  &  wire17650 ) ;
 assign wire2451 = ( wire9500  &  n_n3925  &  wire5513 ) | ( wire9500  &  n_n3925  &  wire5514 ) ;
 assign wire2452 = ( ppeaka_6_6_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2453 = ( wire8330  &  wire4199  &  wire4207 ) ;
 assign wire2454 = ( wire5660  &  wire4199  &  wire3746 ) ;
 assign wire2455 = ( ppeakb_5_5_  &  wire4199  &  wire4215 ) ;
 assign wire2456 = ( wire6560  &  wire4199  &  wire3727 ) ;
 assign wire2457 = ( wire11465  &  wire4199  &  wire3715 ) ;
 assign wire2458 = ( wire15590  &  wire4199  &  wire3723 ) ;
 assign wire2459 = ( wire14105  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2460 = ( wire7670  &  wire4199  &  wire3718 ) ;
 assign wire2461 = ( (~ ppeaka_5_5_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2462 = ( (~ ppeakb_5_5_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2463 = ( ppeakp_5_5_  &  wire4226 ) | ( ppeakp_5_5_  &  wire4199  &  n_n2333 ) ;
 assign wire2464 = ( wire14825  &  wire4199  &  wire3740 ) ;
 assign wire2465 = ( ppeaka_5_5_  &  wire4515 ) | ( ppeaka_5_5_  &  wire4199  &  wire3744 ) ;
 assign wire2466 = ( wire8315  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire2468 = ( wire14435  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire2469 = ( wire15140  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire2472 = ( wire12650  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2473 = ( wire15575  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2474 = ( wire6335  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2476 = ( wire9080  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2479 = ( ppeaka_14_14_  &  wire4515 ) | ( ppeaka_14_14_  &  wire4199  &  wire3744 ) ;
 assign wire2480 = ( ppeaka_7_7_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire2481 = ( wire13340  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire2482 = ( wire14930  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire2483 = ( wire15980  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire2484 = ( wire5915  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire2485 = ( wire14450  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire2486 = ( wire5315  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2488 = ( wire7055  &  wire4226  &  n_n2772 ) ;
 assign wire2489 = ( wire9095  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2491 = ( ppeakb_7_7_  &  wire4515 ) | ( ppeakb_7_7_  &  wire4199  &  wire4211 ) ;
 assign wire2492 = ( (~ preset)  &  wire15785  &  (~ wire17791) ) | ( (~ preset)  &  wire15785  &  wire17843 ) ;
 assign wire2498 = ( (~ preset)  &  wire15725  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15725  &  (~ wire17712) ) ;
 assign wire2500 = ( (~ preset)  &  wire15710  &  wire18103 ) | ( (~ preset)  &  wire15710  &  (~ wire18168) ) ;
 assign wire2501 = ( wire4308  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4308  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4308  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4308  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire2503 = ( wire18176  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire18176  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire18176  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire18176  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire2508 = ( (~ preset)  &  wire15650  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15650  &  (~ wire17715) ) ;
 assign wire2509 = ( (~ preset)  &  pdata_1_1_  &  nrq7_2  &  wire17715 ) ;
 assign wire2510 = ( (~ preset)  &  wire15635  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15635  &  (~ wire17714) ) ;
 assign wire2511 = ( (~ preset)  &  pdata_6_6_  &  nrq7_2  &  wire17714 ) ;
 assign wire2512 = ( (~ preset)  &  wire15620  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15620  &  (~ wire17712) ) ;
 assign wire2513 = ( (~ preset)  &  pdata_15_15_  &  nrq7_2  &  wire17712 ) ;
 assign wire2519 = ( (~ preset)  &  wire15575  &  (~ wire17102) ) | ( (~ preset)  &  wire15575  &  wire17154 ) ;
 assign wire2521 = ( (~ preset)  &  wire15560  &  (~ wire17102) ) | ( (~ preset)  &  wire15560  &  wire17154 ) ;
 assign wire2524 = ( wire13175  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire2525 = ( wire9935  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire2526 = ( wire12890  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire2527 = ( wire8240  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2528 = ( wire10670  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2529 = ( wire15380  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire2530 = ( wire7490  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire2531 = ( wire13400  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire2532 = ( wire6125  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire2533 = ( wire7415  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire2534 = ( wire9455  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2536 = ( wire12605  &  wire4226  &  n_n2772 ) ;
 assign wire2537 = ( wire5390  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2539 = ( ppeaks_0_0_  &  wire17660 ) | ( ppeaks_0_0_  &  wire17662 ) ;
 assign wire2541 = ( wire9710  &  wire4199  &  wire3744 ) ;
 assign wire2542 = ( wire15515  &  wire4515 ) | ( wire15515  &  wire17649 ) | ( wire15515  &  wire17650 ) ;
 assign wire2543 = ( wire13475  &  n_n3925  &  wire5513 ) | ( wire13475  &  n_n3925  &  wire5514 ) ;
 assign wire2545 = ( wire15305  &  wire4199  &  wire3744 ) ;
 assign wire2546 = ( wire15500  &  wire4515 ) | ( wire15500  &  wire17649 ) | ( wire15500  &  wire17650 ) ;
 assign wire2547 = ( wire9800  &  n_n3925  &  wire5513 ) | ( wire9800  &  n_n3925  &  wire5514 ) ;
 assign wire2548 = ( ppeaka_5_5_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2549 = ( wire14765  &  wire4199  &  wire4207 ) ;
 assign wire2550 = ( wire8975  &  wire4199  &  wire3746 ) ;
 assign wire2551 = ( ppeakb_4_4_  &  wire4199  &  wire4215 ) ;
 assign wire2552 = ( wire14870  &  wire4199  &  wire3727 ) ;
 assign wire2553 = ( wire5615  &  wire4199  &  wire3715 ) ;
 assign wire2554 = ( wire13280  &  wire4199  &  wire3723 ) ;
 assign wire2555 = ( wire14525  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2556 = ( wire8300  &  wire4199  &  wire3718 ) ;
 assign wire2557 = ( (~ ppeaka_4_4_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2558 = ( (~ ppeakb_4_4_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2559 = ( ppeakp_4_4_  &  wire4226 ) | ( ppeakp_4_4_  &  wire4199  &  n_n2333 ) ;
 assign wire2560 = ( wire15905  &  wire4199  &  wire3740 ) ;
 assign wire2561 = ( ppeaka_4_4_  &  wire4515 ) | ( ppeaka_4_4_  &  wire4199  &  wire3744 ) ;
 assign wire2562 = ( wire13550  &  wire4199  &  wire4207 ) ;
 assign wire2563 = ( wire6365  &  wire4199  &  wire3746 ) ;
 assign wire2564 = ( ppeakb_15_15_  &  wire4199  &  wire4215 ) ;
 assign wire2565 = ( wire7205  &  wire4199  &  wire3727 ) ;
 assign wire2566 = ( wire12425  &  wire4199  &  wire3715 ) ;
 assign wire2567 = ( wire15950  &  wire4199  &  wire3723 ) ;
 assign wire2568 = ( wire13730  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2569 = ( wire7010  &  wire4199  &  wire3718 ) ;
 assign wire2570 = ( (~ ppeaka_15_15_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2571 = ( (~ ppeakb_15_15_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2572 = ( ppeakp_15_15_  &  wire4226 ) | ( ppeakp_15_15_  &  wire4199  &  n_n2333 ) ;
 assign wire2573 = ( wire15215  &  wire4199  &  wire3740 ) ;
 assign wire2574 = ( ppeaka_15_15_  &  wire4515 ) | ( ppeaka_15_15_  &  wire4199  &  wire3744 ) ;
 assign wire2576 = ( ppeaka_6_6_  &  wire4199  &  wire4224 ) ;
 assign wire2577 = ( wire7865  &  wire4199  &  wire3711 ) ;
 assign wire2578 = ( wire6575  &  wire4199  &  wire3738 ) ;
 assign wire2579 = ( wire15635  &  wire4199  &  wire3720 ) ;
 assign wire2580 = ( wire7160  &  wire4199  &  wire3723 ) ;
 assign wire2581 = ( wire4385  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2582 = ( wire4610  &  wire4199  &  wire3718 ) ;
 assign wire2583 = ( wire7745  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2584 = ( wire10265  &  wire4199  &  wire3744 ) ;
 assign wire2585 = ( ppeakb_6_6_  &  wire4515 ) | ( ppeakb_6_6_  &  wire4199  &  wire4211 ) ;
 assign wire2586 = ( wire7685  &  n_n3925  &  wire5513 ) | ( wire7685  &  n_n3925  &  wire5514 ) ;
 assign wire2587 = ( (~ preset)  &  wire15440  &  (~ wire17791) ) | ( (~ preset)  &  wire15440  &  wire17843 ) ;
 assign wire2592 = ( (~ preset)  &  wire15410  &  (~ wire17427) ) | ( (~ preset)  &  wire15410  &  wire17648 ) ;
 assign wire2594 = ( (~ preset)  &  wire15395  &  (~ wire17427) ) | ( (~ preset)  &  wire15395  &  wire17648 ) ;
 assign wire2595 = ( (~ preset)  &  wire15380  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15380  &  (~ wire17715) ) ;
 assign wire2597 = ( (~ preset)  &  wire15365  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15365  &  (~ wire17714) ) ;
 assign wire2598 = ( wire16928  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire16928  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire16928  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire16928  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire2599 = ( (~ preset)  &  wire15350  &  wire18103 ) | ( (~ preset)  &  wire15350  &  (~ wire18168) ) ;
 assign wire2602 = ( wire18176  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire18176  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire18176  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire18176  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire2607 = ( (~ preset)  &  wire15290  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15290  &  (~ wire17715) ) ;
 assign wire2608 = ( (~ preset)  &  pdata_2_2_  &  nrq7_2  &  wire17715 ) ;
 assign wire2609 = ( (~ preset)  &  wire15275  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15275  &  (~ wire17714) ) ;
 assign wire2610 = ( (~ preset)  &  pdata_9_9_  &  nrq7_2  &  wire17714 ) ;
 assign wire2611 = ( (~ preset)  &  wire15260  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15260  &  (~ wire17712) ) ;
 assign wire2612 = ( (~ preset)  &  pdata_12_12_  &  nrq7_2  &  wire17712 ) ;
 assign wire2614 = ( (~ preset)  &  wire15245  &  (~ wire17167) ) | ( (~ preset)  &  wire15245  &  wire17362 ) ;
 assign wire2618 = ( (~ preset)  &  wire15215  &  (~ wire17102) ) | ( (~ preset)  &  wire15215  &  wire17154 ) ;
 assign wire2620 = ( (~ preset)  &  wire15200  &  (~ wire17102) ) | ( (~ preset)  &  wire15200  &  wire17154 ) ;
 assign wire2623 = ( ppeaka_15_15_  &  wire5413 ) | ( ppeaka_15_15_  &  wire17694 ) ;
 assign wire2625 = ( wire11285  &  n_n3081  &  wire4266 ) ;
 assign wire2626 = ( ppeakp_15_15_  &  wire17696 ) | ( ppeakp_15_15_  &  wire17698 ) | ( ppeakp_15_15_  &  wire17703 ) ;
 assign wire2627 = ( ppeakb_15_15_  &  wire4199  &  wire3744 ) ;
 assign wire2629 = ( wire8915  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire2630 = ( wire10775  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire2631 = ( wire13160  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire2632 = ( wire11225  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2633 = ( wire7595  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2634 = ( wire12590  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire2635 = ( wire9440  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire2636 = ( wire15365  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire2637 = ( wire6815  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire2638 = ( wire10865  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire2639 = ( wire7520  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2641 = ( wire13460  &  wire4226  &  n_n2772 ) ;
 assign wire2642 = ( wire6095  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2644 = ( ppeaks_8_8_  &  wire17660 ) | ( ppeaks_8_8_  &  wire17662 ) ;
 assign wire2646 = ( wire5975  &  wire4199  &  wire3744 ) ;
 assign wire2647 = ( wire15140  &  wire4515 ) | ( wire15140  &  wire17649 ) | ( wire15140  &  wire17650 ) ;
 assign wire2648 = ( wire10070  &  n_n3925  &  wire5513 ) | ( wire10070  &  n_n3925  &  wire5514 ) ;
 assign wire2649 = ( ppeaka_4_4_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2650 = ( wire15860  &  wire4199  &  wire4207 ) ;
 assign wire2651 = ( wire9920  &  wire4199  &  wire3746 ) ;
 assign wire2652 = ( ppeakb_3_3_  &  wire4199  &  wire4215 ) ;
 assign wire2653 = ( wire15245  &  wire4199  &  wire3727 ) ;
 assign wire2654 = ( wire4910  &  wire4199  &  wire3715 ) ;
 assign wire2655 = ( wire13625  &  wire4199  &  wire3723 ) ;
 assign wire2656 = ( wire13355  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2657 = ( wire8960  &  wire4199  &  wire3718 ) ;
 assign wire2658 = ( (~ ppeaka_3_3_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2659 = ( (~ ppeakb_3_3_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2660 = ( ppeakp_3_3_  &  wire4226 ) | ( ppeakp_3_3_  &  wire4199  &  n_n2333 ) ;
 assign wire2661 = ( wire15560  &  wire4199  &  wire3740 ) ;
 assign wire2662 = ( ppeaka_3_3_  &  wire4515 ) | ( ppeaka_3_3_  &  wire4199  &  wire3744 ) ;
 assign wire2663 = ( wire11510  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire2665 = ( wire7190  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire2666 = ( wire15845  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire2669 = ( wire14660  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2670 = ( wire4415  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2671 = ( wire4940  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2673 = ( wire7775  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2676 = ( ppeaka_12_12_  &  wire4515 ) | ( ppeaka_12_12_  &  wire4199  &  wire3744 ) ;
 assign wire2678 = ( ppeaka_9_9_  &  wire4199  &  wire4224 ) ;
 assign wire2679 = ( wire4520  &  wire4199  &  wire3711 ) ;
 assign wire2680 = ( wire7850  &  wire4199  &  wire3738 ) ;
 assign wire2681 = ( wire15275  &  wire4199  &  wire3720 ) ;
 assign wire2682 = ( wire14855  &  wire4199  &  wire3723 ) ;
 assign wire2683 = ( wire15185  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2684 = ( wire6680  &  wire4199  &  wire3718 ) ;
 assign wire2685 = ( wire8390  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2686 = ( wire5990  &  wire4199  &  wire3744 ) ;
 assign wire2687 = ( ppeakb_9_9_  &  wire4515 ) | ( ppeakb_9_9_  &  wire4199  &  wire4211 ) ;
 assign wire2688 = ( wire5720  &  n_n3925  &  wire5513 ) | ( wire5720  &  n_n3925  &  wire5514 ) ;
 assign wire2689 = ( (~ preset)  &  wire15080  &  (~ wire17791) ) | ( (~ preset)  &  wire15080  &  wire17843 ) ;
 assign wire2694 = ( (~ preset)  &  wire15050  &  (~ wire17427) ) | ( (~ preset)  &  wire15050  &  wire17648 ) ;
 assign wire2696 = ( (~ preset)  &  wire15035  &  (~ wire17427) ) | ( (~ preset)  &  wire15035  &  wire17648 ) ;
 assign wire2697 = ( (~ preset)  &  wire15020  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15020  &  (~ wire17715) ) ;
 assign wire2699 = ( (~ preset)  &  wire15005  &  (~ nrq7_2) ) | ( (~ preset)  &  wire15005  &  (~ wire17714) ) ;
 assign wire2700 = ( wire16928  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire16928  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire16928  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire16928  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire2701 = ( (~ preset)  &  wire14990  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14990  &  (~ wire17712) ) ;
 assign wire2702 = ( wire18501  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire18501  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire18501  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire18501  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire2703 = ( (~ preset)  &  wire14975  &  wire18103 ) | ( (~ preset)  &  wire14975  &  (~ wire18168) ) ;
 assign wire2704 = ( wire4308  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4308  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4308  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4308  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire2706 = ( wire18176  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire18176  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire18176  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire18176  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire2709 = ( (~ preset)  &  wire14915  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14915  &  (~ wire17715) ) ;
 assign wire2710 = ( (~ preset)  &  pdata_3_3_  &  nrq7_2  &  wire17715 ) ;
 assign wire2711 = ( (~ preset)  &  wire14900  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14900  &  (~ wire17714) ) ;
 assign wire2712 = ( (~ preset)  &  pdata_8_8_  &  nrq7_2  &  wire17714 ) ;
 assign wire2713 = ( (~ preset)  &  wire14885  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14885  &  (~ wire17712) ) ;
 assign wire2714 = ( (~ preset)  &  pdata_13_13_  &  nrq7_2  &  wire17712 ) ;
 assign wire2716 = ( (~ preset)  &  wire14870  &  (~ wire17167) ) | ( (~ preset)  &  wire14870  &  wire17362 ) ;
 assign wire2722 = ( (~ preset)  &  wire14825  &  (~ wire17102) ) | ( (~ preset)  &  wire14825  &  wire17154 ) ;
 assign wire2725 = ( ppeaka_14_14_  &  wire5413 ) | ( ppeaka_14_14_  &  wire17694 ) ;
 assign wire2727 = ( wire11525  &  n_n3081  &  wire4266 ) ;
 assign wire2728 = ( ppeakp_14_14_  &  wire17696 ) | ( ppeakp_14_14_  &  wire17698 ) | ( ppeakp_14_14_  &  wire17703 ) ;
 assign wire2729 = ( ppeakb_14_14_  &  wire4199  &  wire3744 ) ;
 assign wire2731 = ( wire9590  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire2732 = ( wire11045  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire2733 = ( wire12440  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire2734 = ( wire15770  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2735 = ( wire10685  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2736 = ( wire5465  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire2737 = ( wire8780  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire2738 = ( wire14165  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire2739 = ( wire4745  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire2740 = ( wire11135  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire2741 = ( wire9470  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2743 = ( wire13820  &  wire4226  &  n_n2772 ) ;
 assign wire2744 = ( wire5405  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2746 = ( ppeaks_9_9_  &  wire17660 ) | ( ppeaks_9_9_  &  wire17662 ) ;
 assign wire2748 = ( wire5270  &  wire4199  &  wire3744 ) ;
 assign wire2749 = ( wire14765  &  wire4515 ) | ( wire14765  &  wire17649 ) | ( wire14765  &  wire17650 ) ;
 assign wire2750 = ( wire12875  &  n_n3925  &  wire5513 ) | ( wire12875  &  n_n3925  &  wire5514 ) ;
 assign wire2751 = ( ppeaka_3_3_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2752 = ( wire15515  &  wire4199  &  wire4207 ) ;
 assign wire2753 = ( wire11720  &  wire4199  &  wire3746 ) ;
 assign wire2754 = ( ppeakb_2_2_  &  wire4199  &  wire4215 ) ;
 assign wire2755 = ( wire7805  &  wire4199  &  wire3727 ) ;
 assign wire2756 = ( wire6980  &  wire4199  &  wire3715 ) ;
 assign wire2757 = ( wire14000  &  wire4199  &  wire3723 ) ;
 assign wire2758 = ( wire13715  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2759 = ( wire9635  &  wire4199  &  wire3718 ) ;
 assign wire2760 = ( (~ ppeaka_2_2_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2761 = ( (~ ppeakb_2_2_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2762 = ( ppeakp_2_2_  &  wire4226 ) | ( ppeakp_2_2_  &  wire4199  &  n_n2333 ) ;
 assign wire2763 = ( wire5105  &  wire4199  &  wire3740 ) ;
 assign wire2764 = ( ppeaka_2_2_  &  wire4515 ) | ( ppeaka_2_2_  &  wire4199  &  wire3744 ) ;
 assign wire2765 = ( wire10190  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire2766 = ( ppeakb_13_13_  &  wire4199  &  n_n2772  &  wire4215 ) ;
 assign wire2767 = ( wire14015  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire2768 = ( wire15500  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire2771 = ( wire14240  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2772 = ( wire15920  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2773 = ( wire5645  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2775 = ( wire8420  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2778 = ( ppeaka_13_13_  &  wire4515 ) | ( ppeaka_13_13_  &  wire4199  &  wire3744 ) ;
 assign wire2780 = ( ppeaka_8_8_  &  wire4199  &  wire4224 ) ;
 assign wire2781 = ( wire6605  &  wire4199  &  wire3711 ) ;
 assign wire2782 = ( wire14030  &  wire4199  &  wire3738 ) ;
 assign wire2783 = ( wire14900  &  wire4199  &  wire3720 ) ;
 assign wire2784 = ( wire8435  &  wire4199  &  wire3723 ) ;
 assign wire2785 = ( wire5810  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2786 = ( wire6005  &  wire4199  &  wire3718 ) ;
 assign wire2787 = ( wire9050  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2788 = ( wire6665  &  wire4199  &  wire3744 ) ;
 assign wire2789 = ( ppeakb_8_8_  &  wire4515 ) | ( ppeakb_8_8_  &  wire4199  &  wire4211 ) ;
 assign wire2790 = ( wire6410  &  n_n3925  &  wire5513 ) | ( wire6410  &  n_n3925  &  wire5514 ) ;
 assign wire2791 = ( (~ preset)  &  wire14705  &  (~ wire17791) ) | ( (~ preset)  &  wire14705  &  wire17843 ) ;
 assign wire2800 = ( (~ preset)  &  wire14630  &  (~ wire17427) ) | ( (~ preset)  &  wire14630  &  wire17648 ) ;
 assign wire2802 = ( (~ preset)  &  wire14615  &  (~ nrq4_2) ) ;
 assign wire2803 = ( (~ preset)  &  wire14600  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14600  &  (~ wire17715) ) ;
 assign wire2804 = ( wire17305  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire17305  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire17305  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire17305  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire2805 = ( (~ preset)  &  wire14585  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14585  &  (~ wire17714) ) ;
 assign wire2806 = ( wire16928  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire16928  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire16928  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire16928  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire2807 = ( (~ preset)  &  wire14570  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14570  &  (~ wire17714) ) ;
 assign wire2809 = ( (~ preset)  &  wire14555  &  wire18103 ) | ( (~ preset)  &  wire14555  &  (~ wire18168) ) ;
 assign wire2810 = ( wire4308  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4308  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4308  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4308  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire2812 = ( wire18176  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire18176  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire18176  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire18176  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire2814 = ( wire18176  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire18176  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire18176  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire18176  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire2816 = ( (~ preset)  &  wire14510  &  wire17310 ) | ( (~ preset)  &  wire14510  &  (~ wire17388) ) ;
 assign wire2817 = ( (~ preset)  &  wire14495  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14495  &  (~ wire17715) ) ;
 assign wire2818 = ( (~ preset)  &  pdata_4_4_  &  nrq7_2  &  wire17715 ) ;
 assign wire2819 = ( (~ preset)  &  wire14480  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14480  &  (~ wire17714) ) ;
 assign wire2820 = ( (~ preset)  &  pdata_11_11_  &  nrq7_2  &  wire17714 ) ;
 assign wire2821 = ( (~ preset)  &  wire14465  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14465  &  (~ wire17714) ) ;
 assign wire2822 = ( (~ preset)  &  pdata_2_2_  &  nrq7_2  &  wire17714 ) ;
 assign wire2823 = ( (~ preset)  &  wire14450  &  (~ wire17284) ) | ( (~ preset)  &  wire14450  &  wire18376 ) ;
 assign wire2826 = ( (~ preset)  &  wire14435  &  (~ wire17167) ) | ( (~ preset)  &  wire14435  &  wire17362 ) ;
 assign wire2830 = ( (~ preset)  &  wire14405  &  (~ wire17102) ) | ( (~ preset)  &  wire14405  &  wire17154 ) ;
 assign wire2834 = ( (~ preset)  &  wire14375  &  (~ wire17453) ) | ( (~ preset)  &  wire14375  &  wire18246 ) ;
 assign wire2836 = ( (~ preset)  &  wire14360  &  (~ wire17453) ) | ( (~ preset)  &  wire14360  &  wire18246 ) ;
 assign wire2837 = ( ppeaka_4_4_  &  wire5413 ) | ( ppeaka_4_4_  &  wire17694 ) ;
 assign wire2839 = ( wire15440  &  n_n3081  &  wire4266 ) ;
 assign wire2840 = ( ppeakp_4_4_  &  wire17696 ) | ( ppeakp_4_4_  &  wire17698 ) | ( ppeakp_4_4_  &  wire17703 ) ;
 assign wire2841 = ( ppeakb_4_4_  &  wire4199  &  wire3744 ) ;
 assign wire2843 = ( ppeaka_2_2_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2844 = ( wire5030  &  wire4199  &  wire4207 ) ;
 assign wire2845 = ( wire11495  &  wire4199  &  wire3746 ) ;
 assign wire2846 = ( ppeakb_1_1_  &  wire4199  &  wire4215 ) ;
 assign wire2847 = ( wire7175  &  wire4199  &  wire3727 ) ;
 assign wire2848 = ( wire6305  &  wire4199  &  wire3715 ) ;
 assign wire2849 = ( wire14420  &  wire4199  &  wire3723 ) ;
 assign wire2850 = ( wire15680  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2851 = ( wire4925  &  wire4199  &  wire3718 ) ;
 assign wire2852 = ( (~ ppeaka_1_1_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2853 = ( (~ ppeakb_1_1_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2854 = ( ppeakp_1_1_  &  wire4226 ) | ( ppeakp_1_1_  &  wire4199  &  n_n2333 ) ;
 assign wire2855 = ( wire4400  &  wire4199  &  wire3740 ) ;
 assign wire2856 = ( ppeaka_1_1_  &  wire4515 ) | ( ppeaka_1_1_  &  wire4199  &  wire3744 ) ;
 assign wire2857 = ( ppeaka_11_11_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2858 = ( wire5015  &  wire4199  &  wire4207 ) ;
 assign wire2859 = ( wire11015  &  wire4199  &  wire3746 ) ;
 assign wire2860 = ( ppeakb_10_10_  &  wire4199  &  wire4215 ) ;
 assign wire2861 = ( wire8465  &  wire4199  &  wire3727 ) ;
 assign wire2862 = ( wire13850  &  wire4199  &  wire3715 ) ;
 assign wire2863 = ( wire6515  &  wire4199  &  wire3723 ) ;
 assign wire2864 = ( wire14960  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2865 = ( wire11705  &  wire4199  &  wire3718 ) ;
 assign wire2866 = ( (~ ppeaka_10_10_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2867 = ( (~ ppeakb_10_10_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2868 = ( ppeakp_10_10_  &  wire4226 ) | ( ppeakp_10_10_  &  wire4199  &  n_n2333 ) ;
 assign wire2869 = ( wire13610  &  wire4199  &  wire3740 ) ;
 assign wire2870 = ( ppeaka_10_10_  &  wire4515 ) | ( ppeaka_10_10_  &  wire4199  &  wire3744 ) ;
 assign wire2872 = ( ppeaka_3_3_  &  wire4199  &  wire4224 ) ;
 assign wire2873 = ( wire8510  &  wire4199  &  wire3711 ) ;
 assign wire2874 = ( wire4490  &  wire4199  &  wire3738 ) ;
 assign wire2875 = ( wire14045  &  wire4199  &  wire3720 ) ;
 assign wire2876 = ( wire6530  &  wire4199  &  wire3723 ) ;
 assign wire2877 = ( wire7760  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2878 = ( wire7940  &  wire4199  &  wire3718 ) ;
 assign wire2879 = ( wire13220  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2880 = ( wire9215  &  wire4199  &  wire3744 ) ;
 assign wire2881 = ( ppeakb_3_3_  &  wire4515 ) | ( ppeakb_3_3_  &  wire4199  &  wire4211 ) ;
 assign wire2882 = ( wire15860  &  n_n3925  &  wire5513 ) | ( wire15860  &  n_n3925  &  wire5514 ) ;
 assign wire2883 = ( (~ preset)  &  wire14285  &  (~ wire17791) ) | ( (~ preset)  &  wire14285  &  wire17843 ) ;
 assign wire2892 = ( (~ preset)  &  wire14225  &  wire17999 ) | ( (~ preset)  &  wire14225  &  (~ wire18077) ) ;
 assign wire2894 = ( (~ preset)  &  wire14210  &  (~ wire17427) ) | ( (~ preset)  &  wire14210  &  wire17648 ) ;
 assign wire2895 = ( (~ preset)  &  wire14180  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14180  &  (~ wire17715) ) ;
 assign wire2897 = ( (~ preset)  &  wire14165  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14165  &  (~ wire17714) ) ;
 assign wire2899 = ( (~ preset)  &  wire14150  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14150  &  (~ wire17714) ) ;
 assign wire2900 = ( wire16928  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire16928  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire16928  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire16928  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire2901 = ( (~ preset)  &  wire14135  &  wire18103 ) | ( (~ preset)  &  wire14135  &  (~ wire18168) ) ;
 assign wire2906 = ( wire18176  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire18176  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire18176  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire18176  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire2908 = ( (~ preset)  &  wire14090  &  wire17310 ) | ( (~ preset)  &  wire14090  &  (~ wire17388) ) ;
 assign wire2909 = ( (~ preset)  &  wire14075  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14075  &  (~ wire17715) ) ;
 assign wire2910 = ( (~ preset)  &  pdata_5_5_  &  nrq7_2  &  wire17715 ) ;
 assign wire2911 = ( (~ preset)  &  wire14060  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14060  &  (~ wire17714) ) ;
 assign wire2912 = ( (~ preset)  &  pdata_10_10_  &  nrq7_2  &  wire17714 ) ;
 assign wire2913 = ( (~ preset)  &  wire14045  &  (~ nrq7_2) ) | ( (~ preset)  &  wire14045  &  (~ wire17714) ) ;
 assign wire2914 = ( (~ preset)  &  pdata_3_3_  &  nrq7_2  &  wire17714 ) ;
 assign wire2915 = ( (~ preset)  &  wire14030  &  (~ wire17284) ) | ( (~ preset)  &  wire14030  &  wire18376 ) ;
 assign wire2918 = ( (~ preset)  &  wire14015  &  (~ wire17167) ) | ( (~ preset)  &  wire14015  &  wire17362 ) ;
 assign wire2922 = ( (~ preset)  &  wire13985  &  (~ wire17102) ) | ( (~ preset)  &  wire13985  &  wire17154 ) ;
 assign wire2924 = ( (~ preset)  &  wire13970  &  (~ wire17102) ) | ( (~ preset)  &  wire13970  &  wire17154 ) ;
 assign wire2926 = ( (~ preset)  &  wire13955  &  (~ wire17453) ) | ( (~ preset)  &  wire13955  &  wire18246 ) ;
 assign wire2927 = ( ppeaka_5_5_  &  wire5413 ) | ( ppeaka_5_5_  &  wire17694 ) ;
 assign wire2929 = ( wire15080  &  n_n3081  &  wire4266 ) ;
 assign wire2930 = ( ppeakp_5_5_  &  wire17696 ) | ( ppeakp_5_5_  &  wire17698 ) | ( ppeakp_5_5_  &  wire17703 ) ;
 assign wire2931 = ( ppeakb_5_5_  &  wire4199  &  wire3744 ) ;
 assign wire2933 = ( ppeaka_1_1_  &  wire4199  &  n_n2344  &  wire3784 ) ;
 assign wire2934 = ( wire4310  &  wire4199  &  wire4207 ) ;
 assign wire2935 = ( wire11255  &  wire4199  &  wire3746 ) ;
 assign wire2936 = ( ppeakb_0_0_  &  wire4199  &  wire4215 ) ;
 assign wire2937 = ( wire9110  &  wire4199  &  wire3727 ) ;
 assign wire2938 = ( wire8240  &  wire4199  &  wire3715 ) ;
 assign wire2939 = ( wire14840  &  wire4199  &  wire3723 ) ;
 assign wire2940 = ( wire16025  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire2941 = ( wire11480  &  wire4199  &  wire3718 ) ;
 assign wire2942 = ( (~ ppeaka_0_0_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2943 = ( (~ ppeakb_0_0_)  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire2944 = ( ppeakp_0_0_  &  wire4226 ) | ( ppeakp_0_0_  &  wire4199  &  n_n2333 ) ;
 assign wire2945 = ( wire13970  &  wire4199  &  wire3740 ) ;
 assign wire2946 = ( ppeaka_0_0_  &  wire4515 ) | ( ppeaka_0_0_  &  wire4199  &  wire3744 ) ;
 assign wire2949 = ( wire11735  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire2950 = ( ppeakb_11_11_  &  wire4199  &  n_n2772  &  wire4215 ) ;
 assign wire2951 = ( wire7820  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire2952 = ( wire4295  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire2955 = ( wire13490  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire2956 = ( wire5120  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire2957 = ( wire9650  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire2959 = ( wire7145  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire2962 = ( ppeaka_11_11_  &  wire4515 ) | ( ppeaka_11_11_  &  wire4199  &  wire3744 ) ;
 assign wire2963 = ( (~ preset)  &  wire13895  &  (~ wire17791) ) | ( (~ preset)  &  wire13895  &  wire17843 ) ;
 assign wire2966 = ( wire13880  &  wire4316 ) ;
 assign wire2972 = ( (~ preset)  &  wire13835  &  wire17999 ) | ( (~ preset)  &  wire13835  &  (~ wire18077) ) ;
 assign wire2974 = ( (~ preset)  &  wire13820  &  (~ wire17427) ) | ( (~ preset)  &  wire13820  &  wire17648 ) ;
 assign wire2977 = ( (~ preset)  &  wire13790  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13790  &  (~ wire17715) ) ;
 assign wire2978 = ( wire17305  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire17305  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire17305  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire17305  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire2979 = ( (~ preset)  &  wire13775  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13775  &  (~ wire17714) ) ;
 assign wire2981 = ( (~ preset)  &  wire13745  &  wire18103 ) | ( (~ preset)  &  wire13745  &  (~ wire18168) ) ;
 assign wire2982 = ( wire4308  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4308  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4308  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4308  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire2986 = ( wire18176  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire18176  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire18176  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire18176  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire2988 = ( wire17461  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire17461  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire17461  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire17461  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire2989 = ( (~ preset)  &  wire13685  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13685  &  (~ wire17715) ) ;
 assign wire2990 = ( (~ preset)  &  pdata_6_6_  &  nrq7_2  &  wire17715 ) ;
 assign wire2991 = ( (~ preset)  &  wire13670  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13670  &  (~ wire17714) ) ;
 assign wire2992 = ( (~ preset)  &  pdata_13_13_  &  nrq7_2  &  wire17714 ) ;
 assign wire2993 = ( (~ preset)  &  wire13655  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13655  &  (~ wire17714) ) ;
 assign wire2994 = ( (~ preset)  &  pdata_0_0_  &  nrq7_2  &  wire17714 ) ;
 assign wire2995 = ( (~ preset)  &  wire13640  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13640  &  (~ wire17712) ) ;
 assign wire2996 = ( (~ preset)  &  pdata_2_2_  &  nrq7_2  &  wire17712 ) ;
 assign wire3000 = ( (~ preset)  &  wire13610  &  (~ wire17102) ) | ( (~ preset)  &  wire13610  &  wire17154 ) ;
 assign wire3004 = ( (~ preset)  &  wire13580  &  (~ wire17453) ) | ( (~ preset)  &  wire13580  &  wire18246 ) ;
 assign wire3005 = ( ppeaka_6_6_  &  wire5413 ) | ( ppeaka_6_6_  &  wire17694 ) ;
 assign wire3007 = ( wire14705  &  n_n3081  &  wire4266 ) ;
 assign wire3008 = ( ppeakp_6_6_  &  wire17696 ) | ( ppeakp_6_6_  &  wire17698 ) | ( ppeakp_6_6_  &  wire17703 ) ;
 assign wire3009 = ( ppeakb_6_6_  &  wire4199  &  wire3744 ) ;
 assign wire3012 = ( wire6650  &  wire4199  &  wire3744 ) ;
 assign wire3013 = ( wire13550  &  wire4515 ) | ( wire13550  &  wire17649 ) | ( wire13550  &  wire17650 ) ;
 assign wire3014 = ( wire10355  &  n_n3925  &  wire5513 ) | ( wire10355  &  n_n3925  &  wire5514 ) ;
 assign wire3015 = ( ppeaka_5_5_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire3016 = ( wire14075  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3017 = ( wire7910  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3018 = ( wire5240  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3019 = ( wire7235  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3020 = ( wire5885  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3021 = ( wire9245  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3023 = ( wire8330  &  wire4226  &  n_n2772 ) ;
 assign wire3024 = ( wire7790  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3026 = ( ppeakb_5_5_  &  wire4515 ) | ( ppeakb_5_5_  &  wire4199  &  wire4211 ) ;
 assign wire3032 = ( (~ preset)  &  wire13475  &  wire17999 ) | ( (~ preset)  &  wire13475  &  (~ wire18077) ) ;
 assign wire3034 = ( (~ preset)  &  wire13460  &  (~ wire17427) ) | ( (~ preset)  &  wire13460  &  wire17648 ) ;
 assign wire3037 = ( (~ preset)  &  wire13430  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13430  &  (~ wire17715) ) ;
 assign wire3038 = ( wire17305  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire17305  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire17305  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire17305  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3039 = ( (~ preset)  &  wire13415  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13415  &  (~ wire17714) ) ;
 assign wire3040 = ( wire16928  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire16928  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire16928  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire16928  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3041 = ( (~ preset)  &  wire13400  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13400  &  (~ wire17714) ) ;
 assign wire3043 = ( (~ preset)  &  wire13385  &  wire18103 ) | ( (~ preset)  &  wire13385  &  (~ wire18168) ) ;
 assign wire3044 = ( wire4308  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4308  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4308  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4308  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3049 = ( (~ preset)  &  wire13340  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13340  &  (~ wire17715) ) ;
 assign wire3050 = ( (~ preset)  &  pdata_7_7_  &  nrq7_2  &  wire17715 ) ;
 assign wire3051 = ( (~ preset)  &  wire13325  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13325  &  (~ wire17714) ) ;
 assign wire3052 = ( (~ preset)  &  pdata_12_12_  &  nrq7_2  &  wire17714 ) ;
 assign wire3053 = ( (~ preset)  &  wire13310  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13310  &  (~ wire17714) ) ;
 assign wire3054 = ( (~ preset)  &  pdata_1_1_  &  nrq7_2  &  wire17714 ) ;
 assign wire3055 = ( (~ preset)  &  wire13295  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13295  &  (~ wire17712) ) ;
 assign wire3056 = ( (~ preset)  &  pdata_1_1_  &  nrq7_2  &  wire17712 ) ;
 assign wire3060 = ( (~ preset)  &  wire13265  &  (~ wire17102) ) | ( (~ preset)  &  wire13265  &  wire17154 ) ;
 assign wire3064 = ( (~ preset)  &  wire13235  &  (~ wire17453) ) | ( (~ preset)  &  wire13235  &  wire18246 ) ;
 assign wire3066 = ( (~ preset)  &  wire13220  &  (~ wire17453) ) | ( (~ preset)  &  wire13220  &  wire18246 ) ;
 assign wire3067 = ( wire11270  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire3069 = ( wire9125  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire3070 = ( wire5720  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire3073 = ( wire15770  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire3074 = ( wire13265  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire3075 = ( wire9905  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3077 = ( wire5825  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3080 = ( ppeaka_9_9_  &  wire4515 ) | ( ppeaka_9_9_  &  wire4199  &  wire3744 ) ;
 assign wire3081 = ( ppeaka_4_4_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire3082 = ( wire14495  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3083 = ( wire7280  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3084 = ( wire12545  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3085 = ( wire9170  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3086 = ( wire5195  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3087 = ( wire8585  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3089 = ( wire14765  &  wire4226  &  n_n2772 ) ;
 assign wire3090 = ( wire5840  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3092 = ( ppeakb_4_4_  &  wire4515 ) | ( ppeakb_4_4_  &  wire4199  &  wire4211 ) ;
 assign wire3098 = ( (~ preset)  &  wire13130  &  wire17999 ) | ( (~ preset)  &  wire13130  &  (~ wire18077) ) ;
 assign wire3100 = ( (~ preset)  &  wire13115  &  (~ wire17427) ) | ( (~ preset)  &  wire13115  &  wire17648 ) ;
 assign wire3102 = ( (~ preset)  &  wire13100  &  (~ wire17427) ) | ( (~ preset)  &  wire13100  &  wire17648 ) ;
 assign wire3103 = ( (~ preset)  &  wire13085  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13085  &  (~ wire17715) ) ;
 assign wire3105 = ( (~ preset)  &  wire13070  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13070  &  (~ wire17714) ) ;
 assign wire3107 = ( (~ preset)  &  wire13055  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13055  &  (~ wire17714) ) ;
 assign wire3108 = ( wire16928  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire16928  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire16928  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire16928  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3109 = ( (~ preset)  &  wire13040  &  wire18103 ) | ( (~ preset)  &  wire13040  &  (~ wire18168) ) ;
 assign wire3111 = ( (~ preset)  &  wire13025  &  wire18103 ) | ( (~ preset)  &  wire13025  &  (~ wire18168) ) ;
 assign wire3113 = ( (~ preset)  &  wire13010  &  (~ nrq7_2) ) | ( (~ preset)  &  wire13010  &  (~ wire17715) ) ;
 assign wire3114 = ( (~ preset)  &  pdata_8_8_  &  nrq7_2  &  wire17715 ) ;
 assign wire3115 = ( (~ preset)  &  ppeaki_1_1_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_1_1_  &  wire5522 ) ;
 assign wire3116 = ( wire10805  &  wire5514 ) | ( wire10805  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3120 = ( (~ preset)  &  ppeaki_10_10_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_10_10_  &  wire5522 ) ;
 assign wire3121 = ( wire12935  &  wire5514 ) | ( wire12935  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3124 = ( (~ preset)  &  wire12935  &  (~ wire17570) ) | ( (~ preset)  &  wire12935  &  wire17635 ) ;
 assign wire3132 = ( (~ preset)  &  wire12875  &  wire17999 ) | ( (~ preset)  &  wire12875  &  (~ wire18077) ) ;
 assign wire3134 = ( (~ preset)  &  wire12860  &  (~ wire17427) ) | ( (~ preset)  &  wire12860  &  wire17648 ) ;
 assign wire3136 = ( (~ preset)  &  wire12845  &  (~ wire17427) ) | ( (~ preset)  &  wire12845  &  wire17648 ) ;
 assign wire3137 = ( (~ preset)  &  wire12830  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12830  &  (~ wire17715) ) ;
 assign wire3138 = ( wire17305  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire17305  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire17305  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire17305  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire3139 = ( (~ preset)  &  wire12815  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12815  &  (~ wire17714) ) ;
 assign wire3140 = ( wire16928  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire16928  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire16928  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire16928  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3141 = ( (~ preset)  &  wire12800  &  wire18103 ) | ( (~ preset)  &  wire12800  &  (~ wire18168) ) ;
 assign wire3142 = ( wire4308  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4308  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4308  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4308  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3143 = ( (~ preset)  &  wire12770  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12770  &  (~ wire17714) ) ;
 assign wire3144 = ( (~ preset)  &  pdata_14_14_  &  nrq7_2  &  wire17714 ) ;
 assign wire3145 = ( (~ preset)  &  ppeaki_0_0_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_0_0_  &  wire5522 ) ;
 assign wire3146 = ( wire12695  &  wire5514 ) | ( wire12695  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3150 = ( (~ preset)  &  ppeaki_11_11_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_11_11_  &  wire5522 ) ;
 assign wire3151 = ( wire11600  &  wire5514 ) | ( wire11600  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3154 = ( (~ preset)  &  wire12695  &  (~ wire17570) ) | ( (~ preset)  &  wire12695  &  wire17635 ) ;
 assign wire3162 = ( (~ preset)  &  wire12635  &  wire17999 ) | ( (~ preset)  &  wire12635  &  (~ wire18077) ) ;
 assign wire3164 = ( (~ preset)  &  wire12620  &  (~ wire17427) ) | ( (~ preset)  &  wire12620  &  wire17648 ) ;
 assign wire3166 = ( (~ preset)  &  wire12605  &  (~ wire17427) ) | ( (~ preset)  &  wire12605  &  wire17648 ) ;
 assign wire3167 = ( (~ preset)  &  wire12590  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12590  &  (~ wire17715) ) ;
 assign wire3168 = ( wire17305  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire17305  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire17305  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire17305  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3169 = ( (~ preset)  &  wire12575  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12575  &  (~ wire17714) ) ;
 assign wire3173 = ( (~ preset)  &  wire12545  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12545  &  (~ wire17714) ) ;
 assign wire3174 = ( (~ preset)  &  pdata_4_4_  &  nrq7_2  &  wire17714 ) ;
 assign wire3175 = ( (~ preset)  &  ppeaki_3_3_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_3_3_  &  wire5522 ) ;
 assign wire3176 = ( wire11345  &  wire5514 ) | ( wire11345  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3180 = ( (~ preset)  &  ppeaki_12_12_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_12_12_  &  wire5522 ) ;
 assign wire3183 = ( (~ preset)  &  wire12485  &  (~ wire17570) ) | ( (~ preset)  &  wire12485  &  wire17635 ) ;
 assign wire3185 = ( (~ preset)  &  wire12470  &  wire18142 ) | ( (~ preset)  &  wire12470  &  (~ wire18220) ) ;
 assign wire3191 = ( wire12425  &  wire4331 ) ;
 assign wire3193 = ( (~ preset)  &  wire12410  &  wire17999 ) | ( (~ preset)  &  wire12410  &  (~ wire18077) ) ;
 assign wire3195 = ( (~ preset)  &  wire12395  &  (~ wire17427) ) | ( (~ preset)  &  wire12395  &  wire17648 ) ;
 assign wire3197 = ( (~ preset)  &  wire12380  &  (~ wire17427) ) | ( (~ preset)  &  wire12380  &  wire17648 ) ;
 assign wire3198 = ( (~ preset)  &  wire12365  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12365  &  (~ wire17714) ) ;
 assign wire3200 = ( (~ preset)  &  wire12350  &  (~ nrq7_2) ) | ( (~ preset)  &  wire12350  &  (~ wire17714) ) ;
 assign wire3201 = ( wire16928  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire16928  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire16928  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire16928  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire3203 = ( wire18176  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire18176  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire18176  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire18176  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire3204 = ( (~ preset)  &  ppeaki_2_2_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_2_2_  &  wire5522 ) ;
 assign wire3205 = ( wire11585  &  wire5514 ) | ( wire11585  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3209 = ( (~ preset)  &  ppeaki_13_13_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_13_13_  &  wire5522 ) ;
 assign wire3212 = ( (~ preset)  &  wire12275  &  (~ wire17570) ) | ( (~ preset)  &  wire12275  &  wire17635 ) ;
 assign wire3214 = ( (~ preset)  &  wire12260  &  wire18142 ) | ( (~ preset)  &  wire12260  &  (~ wire18220) ) ;
 assign wire3218 = ( ppeaka_13_13_  &  wire4199  &  wire4224 ) ;
 assign wire3219 = ( wire14885  &  wire4199  &  wire3711 ) ;
 assign wire3220 = ( wire5210  &  wire4199  &  wire3738 ) ;
 assign wire3221 = ( wire13670  &  wire4199  &  wire3720 ) ;
 assign wire3222 = ( wire4460  &  wire4199  &  wire3723 ) ;
 assign wire3223 = ( wire13595  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire3224 = ( wire7325  &  wire4199  &  wire3718 ) ;
 assign wire3225 = ( wire14375  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire3226 = ( wire8570  &  wire4199  &  wire3744 ) ;
 assign wire3227 = ( ppeakb_13_13_  &  wire4515 ) | ( ppeakb_13_13_  &  wire4199  &  wire4211 ) ;
 assign wire3228 = ( wire15500  &  n_n3925  &  wire5513 ) | ( wire15500  &  n_n3925  &  wire5514 ) ;
 assign wire3230 = ( (~ preset)  &  wire12200  &  (~ wire17570) ) | ( (~ preset)  &  wire12200  &  wire17635 ) ;
 assign wire3232 = ( (~ preset)  &  wire12185  &  (~ wire17570) ) | ( (~ preset)  &  wire12185  &  wire17635 ) ;
 assign wire3234 = ( (~ preset)  &  wire12170  &  wire18142 ) | ( (~ preset)  &  wire12170  &  (~ wire18220) ) ;
 assign wire3236 = ( (~ preset)  &  wire12155  &  (~ wire17414) ) | ( (~ preset)  &  wire12155  &  wire17505 ) ;
 assign wire3237 = ( (~ preset)  &  wire12140  &  (~ wire17791) ) | ( (~ preset)  &  wire12140  &  wire17843 ) ;
 assign wire3241 = ( (~ preset)  &  ppeaki_7_7_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_7_7_  &  wire5522 ) ;
 assign wire3242 = ( wire12065  &  wire5514 ) | ( wire12065  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3247 = ( (~ preset)  &  wire12080  &  (~ wire17570) ) | ( (~ preset)  &  wire12080  &  wire17635 ) ;
 assign wire3249 = ( (~ preset)  &  wire12065  &  (~ wire17570) ) | ( (~ preset)  &  wire12065  &  wire17635 ) ;
 assign wire3251 = ( (~ preset)  &  wire12050  &  wire18142 ) | ( (~ preset)  &  wire12050  &  (~ wire18220) ) ;
 assign wire3253 = ( (~ preset)  &  wire12035  &  (~ wire17414) ) | ( (~ preset)  &  wire12035  &  wire17505 ) ;
 assign wire3254 = ( (~ preset)  &  wire12020  &  (~ wire17791) ) | ( (~ preset)  &  wire12020  &  wire17843 ) ;
 assign wire3259 = ( ppeaka_15_15_  &  wire4199  &  wire4224 ) ;
 assign wire3260 = ( wire15620  &  wire4199  &  wire3711 ) ;
 assign wire3261 = ( wire6590  &  wire4199  &  wire3738 ) ;
 assign wire3262 = ( wire4535  &  wire4199  &  wire3720 ) ;
 assign wire3263 = ( wire8450  &  wire4199  &  wire3723 ) ;
 assign wire3264 = ( wire14390  &  wire4199  &  n_n2344  &  wire3770 ) ;
 assign wire3265 = ( wire8600  &  wire4199  &  wire3718 ) ;
 assign wire3266 = ( wire13580  &  wire4199  &  n_n2344  &  wire3775 ) ;
 assign wire3267 = ( wire7295  &  wire4199  &  wire3744 ) ;
 assign wire3268 = ( ppeakb_15_15_  &  wire4515 ) | ( ppeakb_15_15_  &  wire4199  &  wire4211 ) ;
 assign wire3269 = ( wire13550  &  n_n3925  &  wire5513 ) | ( wire13550  &  n_n3925  &  wire5514 ) ;
 assign wire3270 = ( (~ preset)  &  ppeaki_8_8_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_8_8_  &  wire5522 ) ;
 assign wire3271 = ( wire12485  &  wire5514 ) | ( wire12485  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3274 = ( (~ preset)  &  wire11930  &  (~ wire17570) ) | ( (~ preset)  &  wire11930  &  wire17635 ) ;
 assign wire3276 = ( (~ preset)  &  wire11915  &  wire18142 ) | ( (~ preset)  &  wire11915  &  (~ wire18220) ) ;
 assign wire3278 = ( (~ preset)  &  wire11900  &  (~ wire17414) ) | ( (~ preset)  &  wire11900  &  wire17505 ) ;
 assign wire3280 = ( (~ preset)  &  wire11885  &  (~ wire17414) ) | ( (~ preset)  &  wire11885  &  wire17505 ) ;
 assign wire3281 = ( ppeaka_14_14_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire3282 = ( wire7250  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3283 = ( wire7925  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3284 = ( wire12770  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3285 = ( wire15965  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3286 = ( wire4505  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3287 = ( wire9260  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3289 = ( wire15140  &  wire4226  &  n_n2772 ) ;
 assign wire3290 = ( wire5165  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3292 = ( ppeakb_14_14_  &  wire4515 ) | ( ppeakb_14_14_  &  wire4199  &  wire4211 ) ;
 assign wire3293 = ( (~ preset)  &  ppeaki_9_9_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_9_9_  &  wire5522 ) ;
 assign wire3294 = ( wire12275  &  wire5514 ) | ( wire12275  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3297 = ( (~ preset)  &  wire11810  &  (~ wire17570) ) | ( (~ preset)  &  wire11810  &  wire17635 ) ;
 assign wire3299 = ( (~ preset)  &  wire11795  &  wire18142 ) | ( (~ preset)  &  wire11795  &  (~ wire18220) ) ;
 assign wire3301 = ( (~ preset)  &  wire11780  &  (~ wire17414) ) | ( (~ preset)  &  wire11780  &  wire17505 ) ;
 assign wire3303 = ( (~ preset)  &  wire11765  &  (~ wire17414) ) | ( (~ preset)  &  wire11765  &  wire17505 ) ;
 assign wire3304 = ( (~ preset)  &  wire11750  &  (~ wire17791) ) | ( (~ preset)  &  wire11750  &  wire17843 ) ;
 assign wire3315 = ( (~ preset)  &  wire11675  &  wire17037 ) | ( (~ preset)  &  wire11675  &  (~ wire18025) ) ;
 assign wire3317 = ( (~ preset)  &  wire11660  &  wire17037 ) | ( (~ preset)  &  wire11660  &  (~ wire18025) ) ;
 assign wire3322 = ( (~ preset)  &  wire11615  &  (~ nrq7_2) ) | ( (~ preset)  &  wire11615  &  (~ wire17712) ) ;
 assign wire3325 = ( (~ preset)  &  wire11600  &  (~ wire17570) ) | ( (~ preset)  &  wire11600  &  wire17635 ) ;
 assign wire3327 = ( (~ preset)  &  wire11585  &  (~ wire17570) ) | ( (~ preset)  &  wire11585  &  wire17635 ) ;
 assign wire3329 = ( (~ preset)  &  wire11570  &  wire18142 ) | ( (~ preset)  &  wire11570  &  (~ wire18220) ) ;
 assign wire3331 = ( (~ preset)  &  wire11555  &  wire18142 ) | ( (~ preset)  &  wire11555  &  (~ wire18220) ) ;
 assign wire3333 = ( (~ preset)  &  wire11540  &  (~ wire17414) ) | ( (~ preset)  &  wire11540  &  wire17505 ) ;
 assign wire3334 = ( (~ preset)  &  wire11525  &  (~ wire17791) ) | ( (~ preset)  &  wire11525  &  wire17843 ) ;
 assign wire3345 = ( (~ preset)  &  wire11450  &  wire17037 ) | ( (~ preset)  &  wire11450  &  (~ wire18025) ) ;
 assign wire3347 = ( (~ preset)  &  wire11435  &  wire17037 ) | ( (~ preset)  &  wire11435  &  (~ wire18025) ) ;
 assign wire3350 = ( wire4278  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4278  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4278  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4278  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire3352 = ( (~ preset)  &  wire11390  &  (~ nrq7_2) ) | ( (~ preset)  &  wire11390  &  (~ wire17712) ) ;
 assign wire3353 = ( wire18501  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire18501  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire18501  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire18501  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3357 = ( (~ preset)  &  wire11345  &  (~ wire17570) ) | ( (~ preset)  &  wire11345  &  wire17635 ) ;
 assign wire3359 = ( (~ preset)  &  wire11330  &  wire18142 ) | ( (~ preset)  &  wire11330  &  (~ wire18220) ) ;
 assign wire3361 = ( (~ preset)  &  wire11315  &  wire18142 ) | ( (~ preset)  &  wire11315  &  (~ wire18220) ) ;
 assign wire3363 = ( (~ preset)  &  wire11300  &  (~ wire17414) ) | ( (~ preset)  &  wire11300  &  wire17505 ) ;
 assign wire3364 = ( (~ preset)  &  wire11285  &  (~ wire17791) ) | ( (~ preset)  &  wire11285  &  wire17843 ) ;
 assign wire3370 = ( (~ preset)  &  wire11240  &  (~ wire17180) ) | ( (~ preset)  &  wire11240  &  wire17232 ) ;
 assign wire3375 = ( (~ preset)  &  wire11210  &  wire17037 ) | ( (~ preset)  &  wire11210  &  (~ wire18025) ) ;
 assign wire3377 = ( (~ preset)  &  wire11195  &  wire17037 ) | ( (~ preset)  &  wire11195  &  (~ wire18025) ) ;
 assign wire3382 = ( (~ preset)  &  wire11150  &  (~ nrq7_2) ) | ( (~ preset)  &  wire11150  &  (~ wire17712) ) ;
 assign wire3387 = ( wire17461  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire17461  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire17461  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire17461  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire3389 = ( (~ preset)  &  wire11090  &  (~ wire17570) ) | ( (~ preset)  &  wire11090  &  wire17635 ) ;
 assign wire3391 = ( (~ preset)  &  wire11075  &  wire18142 ) | ( (~ preset)  &  wire11075  &  (~ wire18220) ) ;
 assign wire3393 = ( (~ preset)  &  wire11060  &  wire18142 ) | ( (~ preset)  &  wire11060  &  (~ wire18220) ) ;
 assign wire3395 = ( (~ preset)  &  wire11045  &  (~ wire17414) ) | ( (~ preset)  &  wire11045  &  wire17505 ) ;
 assign wire3396 = ( (~ preset)  &  wire11030  &  (~ wire17791) ) | ( (~ preset)  &  wire11030  &  wire17843 ) ;
 assign wire3405 = ( (~ preset)  &  wire10955  &  wire17037 ) | ( (~ preset)  &  wire10955  &  (~ wire18025) ) ;
 assign wire3407 = ( (~ preset)  &  wire10940  &  wire17037 ) | ( (~ preset)  &  wire10940  &  (~ wire18025) ) ;
 assign wire3410 = ( wire4278  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4278  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4278  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4278  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3412 = ( (~ preset)  &  wire10880  &  (~ nrq7_2) ) | ( (~ preset)  &  wire10880  &  (~ wire17712) ) ;
 assign wire3413 = ( wire18501  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire18501  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire18501  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire18501  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire3414 = ( wire4381  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4381  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4381  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4381  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3417 = ( (~ preset)  &  wire10850  &  wire17310 ) | ( (~ preset)  &  wire10850  &  (~ wire17388) ) ;
 assign wire3419 = ( (~ preset)  &  wire10820  &  (~ wire17570) ) | ( (~ preset)  &  wire10820  &  wire17635 ) ;
 assign wire3421 = ( (~ preset)  &  wire10805  &  (~ wire17570) ) | ( (~ preset)  &  wire10805  &  wire17635 ) ;
 assign wire3423 = ( (~ preset)  &  wire10790  &  wire18142 ) | ( (~ preset)  &  wire10790  &  (~ wire18220) ) ;
 assign wire3425 = ( (~ preset)  &  wire10775  &  (~ wire17414) ) | ( (~ preset)  &  wire10775  &  wire17505 ) ;
 assign wire3426 = ( (~ preset)  &  wire10760  &  (~ wire17791) ) | ( (~ preset)  &  wire10760  &  wire17843 ) ;
 assign wire3430 = ( (~ preset)  &  wire10730  &  (~ wire17180) ) | ( (~ preset)  &  wire10730  &  wire17232 ) ;
 assign wire3432 = ( (~ preset)  &  wire10715  &  (~ wire17180) ) | ( (~ preset)  &  wire10715  &  wire17232 ) ;
 assign wire3441 = ( (~ preset)  &  wire10655  &  (~ wire17635) ) | ( (~ preset)  &  wire10655  &  wire17986 ) ;
 assign wire3443 = ( (~ preset)  &  wire10625  &  wire18311 ) | ( (~ preset)  &  wire10625  &  (~ wire18506) ) ;
 assign wire3445 = ( (~ preset)  &  wire10610  &  wire18311 ) | ( (~ preset)  &  wire10610  &  (~ wire18506) ) ;
 assign wire3447 = ( wire4245  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4245  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4245  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4245  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3448 = ( (~ preset)  &  wire10580  &  (~ wire18285) ) | ( (~ preset)  &  wire10580  &  wire18363 ) ;
 assign wire3450 = ( (~ preset)  &  wire10565  &  (~ wire18285) ) | ( (~ preset)  &  wire10565  &  wire18363 ) ;
 assign wire3453 = ( (~ preset)  &  wire10550  &  wire17310 ) | ( (~ preset)  &  wire10550  &  (~ wire17388) ) ;
 assign wire3454 = ( (~ preset)  &  ppeaki_5_5_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_5_5_  &  wire5522 ) ;
 assign wire3455 = ( wire11810  &  wire5514 ) | ( wire11810  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3459 = ( (~ preset)  &  ppeaki_14_14_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_14_14_  &  wire5522 ) ;
 assign wire3462 = ( (~ preset)  &  wire10505  &  wire18142 ) | ( (~ preset)  &  wire10505  &  (~ wire18220) ) ;
 assign wire3464 = ( (~ preset)  &  wire10490  &  (~ wire17414) ) | ( (~ preset)  &  wire10490  &  wire17505 ) ;
 assign wire3466 = ( (~ preset)  &  wire10475  &  (~ wire17414) ) | ( (~ preset)  &  wire10475  &  wire17505 ) ;
 assign wire3469 = ( (~ preset)  &  wire10445  &  (~ wire17180) ) | ( (~ preset)  &  wire10445  &  wire17232 ) ;
 assign wire3471 = ( (~ preset)  &  wire10430  &  (~ wire17180) ) | ( (~ preset)  &  wire10430  &  wire17232 ) ;
 assign wire3478 = ( (~ preset)  &  wire10370  &  (~ wire17635) ) | ( (~ preset)  &  wire10370  &  wire17986 ) ;
 assign wire3480 = ( (~ preset)  &  wire10355  &  wire17999 ) | ( (~ preset)  &  wire10355  &  (~ wire18077) ) ;
 assign wire3481 = ( wire4377  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4377  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4377  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4377  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3482 = ( (~ preset)  &  wire10340  &  wire18311 ) | ( (~ preset)  &  wire10340  &  (~ wire18506) ) ;
 assign wire3483 = ( wire4377  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4377  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4377  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4377  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire3484 = ( (~ preset)  &  wire10325  &  wire18311 ) | ( (~ preset)  &  wire10325  &  (~ wire18506) ) ;
 assign wire3487 = ( (~ preset)  &  wire10280  &  (~ wire18285) ) | ( (~ preset)  &  wire10280  &  wire18363 ) ;
 assign wire3488 = ( wire4306  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4306  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4306  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4306  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3491 = ( (~ preset)  &  ppeaki_4_4_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_4_4_  &  wire5522 ) ;
 assign wire3492 = ( wire11930  &  wire5514 ) | ( wire11930  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3496 = ( (~ preset)  &  ppeaki_15_15_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_15_15_  &  wire5522 ) ;
 assign wire3499 = ( (~ preset)  &  wire10220  &  wire18142 ) | ( (~ preset)  &  wire10220  &  (~ wire18220) ) ;
 assign wire3501 = ( (~ preset)  &  wire10205  &  (~ wire17414) ) | ( (~ preset)  &  wire10205  &  wire17505 ) ;
 assign wire3506 = ( (~ preset)  &  wire10145  &  (~ wire17180) ) | ( (~ preset)  &  wire10145  &  wire17232 ) ;
 assign wire3515 = ( (~ preset)  &  wire10085  &  (~ wire17635) ) | ( (~ preset)  &  wire10085  &  wire17986 ) ;
 assign wire3517 = ( (~ preset)  &  wire10070  &  wire17999 ) | ( (~ preset)  &  wire10070  &  (~ wire18077) ) ;
 assign wire3519 = ( (~ preset)  &  wire10055  &  wire18311 ) | ( (~ preset)  &  wire10055  &  (~ wire18506) ) ;
 assign wire3522 = ( wire10025  &  wire4252 ) ;
 assign wire3531 = ( (~ preset)  &  wire9950  &  wire18142 ) | ( (~ preset)  &  wire9950  &  (~ wire18220) ) ;
 assign wire3533 = ( (~ preset)  &  wire9935  &  (~ wire17414) ) | ( (~ preset)  &  wire9935  &  wire17505 ) ;
 assign wire3538 = ( (~ preset)  &  wire9890  &  (~ wire17180) ) | ( (~ preset)  &  wire9890  &  wire17232 ) ;
 assign wire3540 = ( (~ preset)  &  wire9875  &  (~ wire17180) ) | ( (~ preset)  &  wire9875  &  wire17232 ) ;
 assign wire3549 = ( (~ preset)  &  wire9815  &  (~ wire17635) ) | ( (~ preset)  &  wire9815  &  wire17986 ) ;
 assign wire3551 = ( (~ preset)  &  wire9800  &  wire17999 ) | ( (~ preset)  &  wire9800  &  (~ wire18077) ) ;
 assign wire3552 = ( wire4377  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4377  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4377  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4377  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire3553 = ( (~ preset)  &  wire9785  &  wire18311 ) | ( (~ preset)  &  wire9785  &  (~ wire18506) ) ;
 assign wire3555 = ( wire4245  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4245  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4245  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4245  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3557 = ( wire4243  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4243  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4243  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4243  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3559 = ( wire4243  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4243  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4243  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4243  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire3562 = ( (~ preset)  &  ppeaki_6_6_  &  (~ n_n2772) ) | ( (~ preset)  &  ppeaki_6_6_  &  wire5522 ) ;
 assign wire3563 = ( wire12185  &  wire5514 ) | ( wire12185  &  (~ wire4202)  &  wire4266 ) ;
 assign wire3568 = ( (~ preset)  &  wire9680  &  (~ wire17414) ) | ( (~ preset)  &  wire9680  &  wire17505 ) ;
 assign wire3570 = ( (~ preset)  &  wire9665  &  (~ wire17414) ) | ( (~ preset)  &  wire9665  &  wire17505 ) ;
 assign wire3575 = ( (~ preset)  &  wire9620  &  (~ wire17180) ) | ( (~ preset)  &  wire9620  &  wire17232 ) ;
 assign wire3577 = ( (~ preset)  &  wire9605  &  (~ wire17180) ) | ( (~ preset)  &  wire9605  &  wire17232 ) ;
 assign wire3582 = ( (~ preset)  &  wire9575  &  wire17037 ) | ( (~ preset)  &  wire9575  &  (~ wire18025) ) ;
 assign wire3588 = ( (~ preset)  &  wire9530  &  (~ wire17635) ) | ( (~ preset)  &  wire9530  &  wire17986 ) ;
 assign wire3590 = ( (~ preset)  &  wire9515  &  (~ wire17635) ) | ( (~ preset)  &  wire9515  &  wire17986 ) ;
 assign wire3592 = ( (~ preset)  &  wire9500  &  wire17999 ) | ( (~ preset)  &  wire9500  &  (~ wire18077) ) ;
 assign wire3598 = ( wire9455  &  wire4277 ) ;
 assign wire3599 = ( wire4377  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4377  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4377  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4377  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3600 = ( (~ preset)  &  wire9440  &  wire18311 ) | ( (~ preset)  &  wire9440  &  (~ wire18506) ) ;
 assign wire3602 = ( wire4245  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4245  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4245  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4245  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire3603 = ( (~ preset)  &  wire9395  &  (~ nrq7_2) ) | ( (~ preset)  &  wire9395  &  (~ wire17715) ) ;
 assign wire3605 = ( (~ preset)  &  wire9380  &  (~ nrq7_2) ) | ( (~ preset)  &  wire9380  &  (~ wire17712) ) ;
 assign wire3606 = ( wire18501  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire18501  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire18501  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire18501  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire3611 = ( (~ preset)  &  wire9335  &  (~ wire18285) ) | ( (~ preset)  &  wire9335  &  wire18363 ) ;
 assign wire3612 = ( wire4306  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4306  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4306  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4306  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3613 = ( (~ preset)  &  wire9320  &  (~ wire18285) ) | ( (~ preset)  &  wire9320  &  wire18363 ) ;
 assign wire3614 = ( wire4306  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4306  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4306  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4306  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire3616 = ( wire4243  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4243  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4243  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4243  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3620 = ( wire17461  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire17461  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire17461  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire17461  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire3622 = ( (~ preset)  &  wire9260  &  wire17310 ) | ( (~ preset)  &  wire9260  &  (~ wire17388) ) ;
 assign wire3624 = ( (~ preset)  &  wire9245  &  wire17310 ) | ( (~ preset)  &  wire9245  &  (~ wire17388) ) ;
 assign wire3633 = ( (~ preset)  &  wire9170  &  (~ nrq7_2) ) | ( (~ preset)  &  wire9170  &  (~ wire17712) ) ;
 assign wire3634 = ( (~ preset)  &  pdata_4_4_  &  nrq7_2  &  wire17712 ) ;
 assign wire3635 = ( (~ preset)  &  wire9155  &  (~ wire17284) ) | ( (~ preset)  &  wire9155  &  wire18376 ) ;
 assign wire3637 = ( (~ preset)  &  wire9140  &  (~ wire17284) ) | ( (~ preset)  &  wire9140  &  wire18376 ) ;
 assign wire3640 = ( (~ preset)  &  wire9125  &  (~ wire17167) ) | ( (~ preset)  &  wire9125  &  wire17362 ) ;
 assign wire3642 = ( (~ preset)  &  wire9110  &  (~ wire17167) ) | ( (~ preset)  &  wire9110  &  wire17362 ) ;
 assign wire3650 = ( (~ preset)  &  wire9050  &  (~ wire17453) ) | ( (~ preset)  &  wire9050  &  wire18246 ) ;
 assign wire3651 = ( ppeaka_0_0_  &  wire5413 ) | ( ppeaka_0_0_  &  wire17694 ) ;
 assign wire3653 = ( wire5675  &  n_n3081  &  wire4266 ) ;
 assign wire3654 = ( ppeakp_0_0_  &  wire17696 ) | ( ppeakp_0_0_  &  wire17698 ) | ( ppeakp_0_0_  &  wire17703 ) ;
 assign wire3655 = ( ppeakb_0_0_  &  wire4199  &  wire3744 ) ;
 assign wire3657 = ( ppeaka_9_9_  &  wire5413 ) | ( ppeaka_9_9_  &  wire17694 ) ;
 assign wire3659 = ( wire11750  &  n_n3081  &  wire4266 ) ;
 assign wire3660 = ( ppeakp_9_9_  &  wire17696 ) | ( ppeakp_9_9_  &  wire17698 ) | ( ppeakp_9_9_  &  wire17703 ) ;
 assign wire3661 = ( ppeakb_9_9_  &  wire4199  &  wire3744 ) ;
 assign wire3663 = ( wire12680  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire3664 = ( wire10475  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire3665 = ( wire15425  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire3666 = ( wire6980  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire3667 = ( wire10100  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire3668 = ( wire14600  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3669 = ( wire10325  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3670 = ( wire14150  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3671 = ( wire10880  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3672 = ( wire8690  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3673 = ( wire5510  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3675 = ( wire13100  &  wire4226  &  n_n2772 ) ;
 assign wire3676 = ( wire9320  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3678 = ( ppeaks_2_2_  &  wire17660 ) | ( ppeaks_2_2_  &  wire17662 ) ;
 assign wire3679 = ( wire10130  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire3680 = ( wire10490  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire3681 = ( wire12125  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire3682 = ( wire13490  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire3683 = ( wire10115  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire3684 = ( wire6830  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3685 = ( wire7505  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3686 = ( wire13415  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3687 = ( wire11390  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3688 = ( wire7430  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3689 = ( wire5525  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3691 = ( wire13115  &  wire4226  &  n_n2772 ) ;
 assign wire3692 = ( wire9335  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3694 = ( ppeaks_11_11_  &  wire17660 ) | ( ppeaks_11_11_  &  wire17662 ) ;
 assign wire3699 = ( (~ preset)  &  wire8945  &  (~ wire17180) ) | ( (~ preset)  &  wire8945  &  wire17232 ) ;
 assign wire3701 = ( (~ preset)  &  wire8930  &  (~ wire17180) ) | ( (~ preset)  &  wire8930  &  wire17232 ) ;
 assign wire3706 = ( (~ preset)  &  wire8900  &  wire17037 ) | ( (~ preset)  &  wire8900  &  (~ wire18025) ) ;
 assign wire3713 = ( (~ preset)  &  wire8855  &  (~ wire17635) ) | ( (~ preset)  &  wire8855  &  wire17986 ) ;
 assign wire3716 = ( (~ preset)  &  wire8840  &  (~ wire17635) ) | ( (~ preset)  &  wire8840  &  wire17986 ) ;
 assign wire3719 = ( (~ preset)  &  wire8825  &  wire17999 ) | ( (~ preset)  &  wire8825  &  (~ wire18077) ) ;
 assign wire3721 = ( wire4278  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4278  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4278  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4278  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3725 = ( (~ preset)  &  wire8780  &  wire18311 ) | ( (~ preset)  &  wire8780  &  (~ wire18506) ) ;
 assign wire3730 = ( wire4245  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4245  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4245  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4245  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3731 = ( (~ preset)  &  wire8735  &  (~ nrq7_2) ) | ( (~ preset)  &  wire8735  &  (~ wire17715) ) ;
 assign wire3733 = ( (~ preset)  &  wire8720  &  (~ nrq7_2) ) | ( (~ preset)  &  wire8720  &  (~ wire17712) ) ;
 assign wire3735 = ( wire4381  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4381  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4381  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4381  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3737 = ( wire4381  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4381  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4381  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4381  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire3741 = ( (~ preset)  &  wire8675  &  (~ wire18285) ) | ( (~ preset)  &  wire8675  &  wire18363 ) ;
 assign wire3743 = ( (~ preset)  &  wire8660  &  (~ wire18285) ) | ( (~ preset)  &  wire8660  &  wire18363 ) ;
 assign wire3749 = ( wire4243  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4243  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4243  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4243  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3751 = ( wire8630  &  wire4253 ) ;
 assign wire3757 = ( (~ preset)  &  wire8600  &  wire17310 ) | ( (~ preset)  &  wire8600  &  (~ wire17388) ) ;
 assign wire3759 = ( (~ preset)  &  wire8585  &  wire17310 ) | ( (~ preset)  &  wire8585  &  (~ wire17388) ) ;
 assign wire3768 = ( (~ preset)  &  wire8510  &  (~ nrq7_2) ) | ( (~ preset)  &  wire8510  &  (~ wire17712) ) ;
 assign wire3769 = ( (~ preset)  &  pdata_3_3_  &  nrq7_2  &  wire17712 ) ;
 assign wire3771 = ( (~ preset)  &  wire8495  &  (~ wire17284) ) | ( (~ preset)  &  wire8495  &  wire18376 ) ;
 assign wire3773 = ( (~ preset)  &  wire8480  &  (~ wire17284) ) | ( (~ preset)  &  wire8480  &  wire18376 ) ;
 assign wire3777 = ( (~ preset)  &  wire8465  &  (~ wire17167) ) | ( (~ preset)  &  wire8465  &  wire17362 ) ;
 assign wire3788 = ( (~ preset)  &  wire8390  &  (~ wire17453) ) | ( (~ preset)  &  wire8390  &  wire18246 ) ;
 assign wire3789 = ( ppeaka_1_1_  &  wire5413 ) | ( ppeaka_1_1_  &  wire17694 ) ;
 assign wire3791 = ( wire4970  &  n_n3081  &  wire4266 ) ;
 assign wire3792 = ( ppeakp_1_1_  &  wire17696 ) | ( ppeakp_1_1_  &  wire17698 ) | ( ppeakp_1_1_  &  wire17703 ) ;
 assign wire3793 = ( ppeakb_1_1_  &  wire4199  &  wire3744 ) ;
 assign wire3795 = ( ppeaka_8_8_  &  wire5413 ) | ( ppeaka_8_8_  &  wire17694 ) ;
 assign wire3797 = ( wire13895  &  n_n3081  &  wire4266 ) ;
 assign wire3798 = ( ppeakp_8_8_  &  wire17696 ) | ( ppeakp_8_8_  &  wire17698 ) | ( ppeakp_8_8_  &  wire17703 ) ;
 assign wire3799 = ( ppeakb_8_8_  &  wire4199  &  wire3744 ) ;
 assign wire3801 = ( wire12455  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire3802 = ( wire12155  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire3803 = ( wire14255  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire3804 = ( wire4910  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire3805 = ( wire5570  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire3806 = ( wire14180  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3807 = ( wire10610  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3808 = ( wire12575  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3809 = ( wire8720  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3810 = ( wire9350  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3811 = ( wire6200  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3813 = ( wire12845  &  wire4226  &  n_n2772 ) ;
 assign wire3814 = ( wire7385  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3816 = ( ppeaks_3_3_  &  wire17660 ) | ( ppeaks_3_3_  &  wire17662 ) ;
 assign wire3818 = ( wire4565  &  wire4199  &  wire3744 ) ;
 assign wire3819 = ( wire8330  &  wire4515 ) | ( wire8330  &  wire17649 ) | ( wire8330  &  wire17650 ) ;
 assign wire3820 = ( wire12635  &  n_n3925  &  wire5513 ) | ( wire12635  &  n_n3925  &  wire5514 ) ;
 assign wire3825 = ( (~ preset)  &  wire8285  &  (~ wire17180) ) | ( (~ preset)  &  wire8285  &  wire17232 ) ;
 assign wire3834 = ( (~ preset)  &  wire8210  &  (~ wire17635) ) | ( (~ preset)  &  wire8210  &  wire17986 ) ;
 assign wire3836 = ( (~ preset)  &  wire8195  &  (~ wire17635) ) | ( (~ preset)  &  wire8195  &  wire17986 ) ;
 assign wire3838 = ( (~ preset)  &  wire8180  &  wire17999 ) | ( (~ preset)  &  wire8180  &  (~ wire18077) ) ;
 assign wire3842 = ( (~ preset)  &  wire8150  &  wire18311 ) | ( (~ preset)  &  wire8150  &  (~ wire18506) ) ;
 assign wire3843 = ( wire4377  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4377  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4377  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4377  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3844 = ( (~ preset)  &  wire8135  &  wire18311 ) | ( (~ preset)  &  wire8135  &  (~ wire18506) ) ;
 assign wire3846 = ( (~ preset)  &  wire8120  &  wire18311 ) | ( (~ preset)  &  wire8120  &  (~ wire18506) ) ;
 assign wire3848 = ( wire4245  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4245  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4245  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4245  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3849 = ( (~ preset)  &  wire8090  &  (~ nrq7_2) ) | ( (~ preset)  &  wire8090  &  (~ wire17715) ) ;
 assign wire3850 = ( wire17305  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire17305  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire17305  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire17305  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3851 = ( (~ preset)  &  wire8075  &  (~ nrq7_2) ) | ( (~ preset)  &  wire8075  &  (~ wire17712) ) ;
 assign wire3853 = ( wire4381  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4381  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4381  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4381  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire3857 = ( (~ preset)  &  wire8030  &  (~ wire18285) ) | ( (~ preset)  &  wire8030  &  wire18363 ) ;
 assign wire3858 = ( wire4306  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4306  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4306  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4306  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire3859 = ( (~ preset)  &  wire8015  &  (~ wire18285) ) | ( (~ preset)  &  wire8015  &  wire18363 ) ;
 assign wire3860 = ( wire4306  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4306  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4306  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4306  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire3862 = ( wire4243  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4243  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4243  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4243  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3866 = ( (~ preset)  &  wire7955  &  wire17310 ) | ( (~ preset)  &  wire7955  &  (~ wire17388) ) ;
 assign wire3868 = ( (~ preset)  &  wire7940  &  wire17310 ) | ( (~ preset)  &  wire7940  &  (~ wire17388) ) ;
 assign wire3875 = ( (~ preset)  &  wire7880  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7880  &  (~ wire17715) ) ;
 assign wire3876 = ( (~ preset)  &  pdata_15_15_  &  nrq7_2  &  wire17715 ) ;
 assign wire3877 = ( (~ preset)  &  wire7865  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7865  &  (~ wire17712) ) ;
 assign wire3878 = ( (~ preset)  &  pdata_6_6_  &  nrq7_2  &  wire17712 ) ;
 assign wire3879 = ( (~ preset)  &  wire7850  &  (~ wire17284) ) | ( (~ preset)  &  wire7850  &  wire18376 ) ;
 assign wire3881 = ( (~ preset)  &  wire7835  &  (~ wire17284) ) | ( (~ preset)  &  wire7835  &  wire18376 ) ;
 assign wire3884 = ( (~ preset)  &  wire7820  &  (~ wire17167) ) | ( (~ preset)  &  wire7820  &  wire17362 ) ;
 assign wire3886 = ( (~ preset)  &  wire7805  &  (~ wire17167) ) | ( (~ preset)  &  wire7805  &  wire17362 ) ;
 assign wire3894 = ( (~ preset)  &  wire7745  &  (~ wire17453) ) | ( (~ preset)  &  wire7745  &  wire18246 ) ;
 assign wire3895 = ( ppeaka_2_2_  &  wire5413 ) | ( ppeaka_2_2_  &  wire17694 ) ;
 assign wire3897 = ( ndout  &  n_n3081  &  wire4266 ) ;
 assign wire3898 = ( ppeakp_2_2_  &  wire17696 ) | ( ppeakp_2_2_  &  wire17698 ) | ( ppeakp_2_2_  &  wire17703 ) ;
 assign wire3899 = ( ppeakb_2_2_  &  wire4199  &  wire3744 ) ;
 assign wire3901 = ( ppeaka_7_7_  &  wire5413 ) | ( ppeaka_7_7_  &  wire17694 ) ;
 assign wire3903 = ( wire14285  &  n_n3081  &  wire4266 ) ;
 assign wire3904 = ( ppeakp_7_7_  &  wire17696 ) | ( ppeakp_7_7_  &  wire17698 ) | ( ppeakp_7_7_  &  wire17703 ) ;
 assign wire3905 = ( ppeakb_7_7_  &  wire4199  &  wire3744 ) ;
 assign wire3907 = ( wire10700  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire3908 = ( wire12035  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire3909 = ( wire14690  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire3910 = ( wire14240  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire3911 = ( wire8885  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire3912 = ( wire8090  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire3913 = ( wire10340  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire3914 = ( wire12815  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire3915 = ( wire14990  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire3916 = ( wire8705  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire3917 = ( wire6890  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire3919 = ( wire12620  &  wire4226  &  n_n2772 ) ;
 assign wire3920 = ( wire8030  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire3922 = ( ppeaks_13_13_  &  wire17660 ) | ( ppeaks_13_13_  &  wire17662 ) ;
 assign wire3924 = ( wire6635  &  wire4199  &  wire3744 ) ;
 assign wire3925 = ( wire7685  &  wire4515 ) | ( wire7685  &  wire17649 ) | ( wire7685  &  wire17650 ) ;
 assign wire3926 = ( wire12410  &  n_n3925  &  wire5513 ) | ( wire12410  &  n_n3925  &  wire5514 ) ;
 assign wire3929 = ( (~ preset)  &  wire7655  &  (~ wire17180) ) | ( (~ preset)  &  wire7655  &  wire17232 ) ;
 assign wire3931 = ( (~ preset)  &  wire7640  &  (~ wire17180) ) | ( (~ preset)  &  wire7640  &  wire17232 ) ;
 assign wire3938 = ( (~ preset)  &  wire7580  &  (~ wire17635) ) | ( (~ preset)  &  wire7580  &  wire17986 ) ;
 assign wire3940 = ( (~ preset)  &  wire7565  &  (~ wire17635) ) | ( (~ preset)  &  wire7565  &  wire17986 ) ;
 assign wire3942 = ( (~ preset)  &  wire7550  &  wire17999 ) | ( (~ preset)  &  wire7550  &  (~ wire18077) ) ;
 assign wire3945 = ( wire4278  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4278  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4278  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4278  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3947 = ( wire4377  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4377  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4377  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4377  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3948 = ( (~ preset)  &  wire7505  &  wire18311 ) | ( (~ preset)  &  wire7505  &  (~ wire18506) ) ;
 assign wire3950 = ( (~ preset)  &  wire7490  &  wire18311 ) | ( (~ preset)  &  wire7490  &  (~ wire18506) ) ;
 assign wire3953 = ( (~ preset)  &  wire7460  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7460  &  (~ wire17715) ) ;
 assign wire3955 = ( (~ preset)  &  wire7445  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7445  &  (~ wire17712) ) ;
 assign wire3956 = ( wire18501  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire18501  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire18501  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire18501  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire3957 = ( wire4381  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4381  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4381  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4381  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire3960 = ( wire7415  &  wire4317 ) ;
 assign wire3961 = ( (~ preset)  &  wire7400  &  (~ wire18285) ) | ( (~ preset)  &  wire7400  &  wire18363 ) ;
 assign wire3963 = ( (~ preset)  &  wire7385  &  (~ wire18285) ) | ( (~ preset)  &  wire7385  &  wire18363 ) ;
 assign wire3967 = ( (~ preset)  &  wire7355  &  wire18103 ) | ( (~ preset)  &  wire7355  &  (~ wire18168) ) ;
 assign wire3970 = ( wire17461  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire17461  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire17461  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire17461  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire3972 = ( (~ preset)  &  wire7325  &  wire17310 ) | ( (~ preset)  &  wire7325  &  (~ wire17388) ) ;
 assign wire3974 = ( (~ preset)  &  wire7310  &  wire17310 ) | ( (~ preset)  &  wire7310  &  (~ wire17388) ) ;
 assign wire3981 = ( (~ preset)  &  wire7250  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7250  &  (~ wire17715) ) ;
 assign wire3982 = ( (~ preset)  &  pdata_14_14_  &  nrq7_2  &  wire17715 ) ;
 assign wire3983 = ( (~ preset)  &  wire7235  &  (~ nrq7_2) ) | ( (~ preset)  &  wire7235  &  (~ wire17712) ) ;
 assign wire3984 = ( (~ preset)  &  pdata_5_5_  &  nrq7_2  &  wire17712 ) ;
 assign wire3985 = ( (~ preset)  &  wire7220  &  (~ wire17284) ) | ( (~ preset)  &  wire7220  &  wire18376 ) ;
 assign wire3988 = ( (~ preset)  &  wire7205  &  (~ wire17167) ) | ( (~ preset)  &  wire7205  &  wire17362 ) ;
 assign wire3990 = ( (~ preset)  &  wire7190  &  (~ wire17167) ) | ( (~ preset)  &  wire7190  &  wire17362 ) ;
 assign wire3992 = ( (~ preset)  &  wire7175  &  (~ wire17167) ) | ( (~ preset)  &  wire7175  &  wire17362 ) ;
 assign wire4000 = ( (~ preset)  &  wire7115  &  (~ wire17453) ) | ( (~ preset)  &  wire7115  &  wire18246 ) ;
 assign wire4001 = ( ppeaka_3_3_  &  wire5413 ) | ( ppeaka_3_3_  &  wire17694 ) ;
 assign wire4003 = ( wire15785  &  n_n3081  &  wire4266 ) ;
 assign wire4004 = ( ppeakp_3_3_  &  wire17696 ) | ( ppeakp_3_3_  &  wire17698 ) | ( ppeakp_3_3_  &  wire17703 ) ;
 assign wire4005 = ( ppeakb_3_3_  &  wire4199  &  wire3744 ) ;
 assign wire4007 = ( wire12920  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4008 = ( wire9665  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4009 = ( wire12005  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4010 = ( wire6305  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4011 = ( wire9830  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4012 = ( wire15020  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4013 = ( wire8120  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4014 = ( wire14570  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4015 = ( wire11150  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4016 = ( wire8045  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4017 = ( wire4805  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4019 = ( wire12380  &  wire4226  &  n_n2772 ) ;
 assign wire4020 = ( wire8660  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4022 = ( ppeaks_1_1_  &  wire17660 ) | ( ppeaks_1_1_  &  wire17662 ) ;
 assign wire4023 = ( wire10415  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4025 = ( wire9680  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4026 = ( wire15065  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4027 = ( wire14660  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4028 = ( wire9845  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4029 = ( wire7460  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4030 = ( wire10625  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4031 = ( wire13775  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4032 = ( wire11615  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4033 = ( wire9365  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4034 = ( wire4820  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4036 = ( wire12395  &  wire4226  &  n_n2772 ) ;
 assign wire4037 = ( wire8675  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4039 = ( ppeaks_12_12_  &  wire17660 ) | ( ppeaks_12_12_  &  wire17662 ) ;
 assign wire4041 = ( wire5960  &  wire4199  &  wire3744 ) ;
 assign wire4042 = ( wire7055  &  wire4515 ) | ( wire7055  &  wire17649 ) | ( wire7055  &  wire17650 ) ;
 assign wire4043 = ( wire6245  &  n_n3925  &  wire5513 ) | ( wire6245  &  n_n3925  &  wire5514 ) ;
 assign wire4047 = ( wire7010  &  wire4277 ) ;
 assign wire4056 = ( (~ preset)  &  wire6965  &  wire17037 ) | ( (~ preset)  &  wire6965  &  (~ wire18025) ) ;
 assign wire4058 = ( (~ preset)  &  wire6950  &  wire17037 ) | ( (~ preset)  &  wire6950  &  (~ wire18025) ) ;
 assign wire4060 = ( (~ preset)  &  wire6935  &  (~ wire17635) ) | ( (~ preset)  &  wire6935  &  wire17986 ) ;
 assign wire4062 = ( (~ preset)  &  wire6920  &  wire17999 ) | ( (~ preset)  &  wire6920  &  (~ wire18077) ) ;
 assign wire4065 = ( wire4278  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4278  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4278  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4278  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire4067 = ( wire4278  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4278  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4278  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4278  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire4073 = ( (~ preset)  &  wire6830  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6830  &  (~ wire17715) ) ;
 assign wire4074 = ( wire17305  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire17305  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire17305  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire17305  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire4075 = ( (~ preset)  &  wire6815  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6815  &  (~ wire17712) ) ;
 assign wire4076 = ( wire18501  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire18501  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire18501  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire18501  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire4077 = ( wire4381  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4381  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4381  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4381  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire4079 = ( (~ preset)  &  wire6770  &  (~ wire18285) ) | ( (~ preset)  &  wire6770  &  wire18363 ) ;
 assign wire4080 = ( wire4306  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4306  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4306  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4306  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire4085 = ( (~ preset)  &  wire6725  &  wire18103 ) | ( (~ preset)  &  wire6725  &  (~ wire18168) ) ;
 assign wire4088 = ( wire17461  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire17461  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire17461  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire17461  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire4090 = ( wire17461  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire17461  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire17461  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire17461  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire4092 = ( (~ preset)  &  wire6680  &  wire17310 ) | ( (~ preset)  &  wire6680  &  (~ wire17388) ) ;
 assign wire4099 = ( (~ preset)  &  wire6620  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6620  &  (~ wire17715) ) ;
 assign wire4100 = ( (~ preset)  &  pdata_13_13_  &  nrq7_2  &  wire17715 ) ;
 assign wire4101 = ( (~ preset)  &  wire6605  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6605  &  (~ wire17712) ) ;
 assign wire4102 = ( (~ preset)  &  pdata_8_8_  &  nrq7_2  &  wire17712 ) ;
 assign wire4103 = ( (~ preset)  &  wire6590  &  (~ wire17284) ) | ( (~ preset)  &  wire6590  &  wire18376 ) ;
 assign wire4105 = ( (~ preset)  &  wire6575  &  (~ wire17284) ) | ( (~ preset)  &  wire6575  &  wire18376 ) ;
 assign wire4108 = ( (~ preset)  &  wire6560  &  (~ wire17167) ) | ( (~ preset)  &  wire6560  &  wire17362 ) ;
 assign wire4120 = ( (~ preset)  &  wire6470  &  (~ wire17453) ) | ( (~ preset)  &  wire6470  &  wire18246 ) ;
 assign wire4121 = ( ppeaka_13_13_  &  wire5413 ) | ( ppeaka_13_13_  &  wire17694 ) ;
 assign wire4123 = ( wire10760  &  n_n3081  &  wire4266 ) ;
 assign wire4124 = ( ppeakp_13_13_  &  wire17696 ) | ( ppeakp_13_13_  &  wire17698 ) | ( ppeakp_13_13_  &  wire17703 ) ;
 assign wire4125 = ( ppeakb_13_13_  &  wire4199  &  wire3744 ) ;
 assign wire4127 = ( wire7625  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4128 = ( wire11300  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4129 = ( wire13865  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4130 = ( wire11690  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4131 = ( wire8870  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4132 = ( wire13085  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4133 = ( wire5495  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4134 = ( wire16085  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4135 = ( wire8075  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4136 = ( wire6110  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4137 = ( wire11165  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4139 = ( wire14210  &  wire4226  &  n_n2772 ) ;
 assign wire4140 = ( wire10565  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4142 = ( ppeaks_6_6_  &  wire17660 ) | ( ppeaks_6_6_  &  wire17662 ) ;
 assign wire4143 = ( wire6320  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4144 = ( wire11780  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4145 = ( wire13880  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4146 = ( wire12425  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4147 = ( wire4880  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4148 = ( wire9395  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4149 = ( wire8150  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4150 = ( wire12365  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4151 = ( wire15725  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4152 = ( wire4730  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4153 = ( wire11180  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4155 = ( wire15050  &  wire4226  &  n_n2772 ) ;
 assign wire4156 = ( wire10580  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4158 = ( ppeaks_15_15_  &  wire17660 ) | ( ppeaks_15_15_  &  wire17662 ) ;
 assign wire4160 = ( wire7895  &  wire4199  &  wire3744 ) ;
 assign wire4161 = ( wire6410  &  wire4515 ) | ( wire6410  &  wire17649 ) | ( wire6410  &  wire17650 ) ;
 assign wire4162 = ( wire6920  &  n_n3925  &  wire5513 ) | ( wire6920  &  n_n3925  &  wire5514 ) ;
 assign wire4163 = ( ppeaka_2_2_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire4164 = ( wire15290  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4165 = ( wire8555  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4166 = ( wire14465  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4167 = ( wire13640  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4168 = ( wire9140  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4169 = ( wire7310  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4171 = ( wire15515  &  wire4226  &  n_n2772 ) ;
 assign wire4172 = ( wire4445  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4174 = ( ppeakb_2_2_  &  wire4515 ) | ( ppeakb_2_2_  &  wire4199  &  wire4211 ) ;
 assign wire4175 = ( ppeaka_11_11_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire4176 = ( wire5255  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4177 = ( wire4595  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4178 = ( wire14480  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4179 = ( wire5930  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4180 = ( wire9155  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4181 = ( wire14090  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4183 = ( wire4295  &  wire4226  &  n_n2772 ) ;
 assign wire4184 = ( wire5855  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4186 = ( ppeakb_11_11_  &  wire4515 ) | ( ppeakb_11_11_  &  wire4199  &  wire4211 ) ;
 assign wire4188 = ( wire6365  &  wire4336 ) ;
 assign wire4196 = ( wire6320  &  wire4325 ) ;
 assign wire4213 = ( (~ preset)  &  wire6290  &  wire17037 ) | ( (~ preset)  &  wire6290  &  (~ wire18025) ) ;
 assign wire4218 = ( (~ preset)  &  wire6275  &  wire17037 ) | ( (~ preset)  &  wire6275  &  (~ wire18025) ) ;
 assign wire4227 = ( (~ preset)  &  wire6260  &  (~ wire17635) ) | ( (~ preset)  &  wire6260  &  wire17986 ) ;
 assign wire4230 = ( (~ preset)  &  wire6245  &  wire17999 ) | ( (~ preset)  &  wire6245  &  (~ wire18077) ) ;
 assign wire4246 = ( wire4377  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4377  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4377  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4377  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire4247 = ( (~ preset)  &  wire6185  &  wire18311 ) | ( (~ preset)  &  wire6185  &  (~ wire18506) ) ;
 assign wire4249 = ( wire4245  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4245  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4245  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4245  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire4250 = ( (~ preset)  &  wire6155  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6155  &  (~ wire17715) ) ;
 assign wire4251 = ( wire17305  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire17305  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire17305  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire17305  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire4257 = ( (~ preset)  &  wire6140  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6140  &  (~ wire17712) ) ;
 assign wire4262 = ( wire18501  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire18501  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire18501  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire18501  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire4263 = ( (~ preset)  &  wire6125  &  (~ nrq7_2) ) | ( (~ preset)  &  wire6125  &  (~ wire17712) ) ;
 assign wire4291 = ( (~ preset)  &  wire6095  &  (~ wire18285) ) | ( (~ preset)  &  wire6095  &  wire18363 ) ;
 assign wire4406 = ( wire4306  &  n_n2479  &  wire19495  &  wire19743 ) | ( wire4306  &  (~ n_n2479)  &  (~ wire19495)  &  wire19743 ) | ( wire4306  &  (~ n_n2479)  &  wire19495  &  (~ wire19743) ) | ( wire4306  &  n_n2479  &  (~ wire19495)  &  (~ wire19743) ) ;
 assign wire4492 = ( wire4243  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4243  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4243  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4243  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire4493 = ( (~ preset)  &  wire6050  &  wire18103 ) | ( (~ preset)  &  wire6050  &  (~ wire18168) ) ;
 assign wire4494 = ( wire4308  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4308  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4308  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4308  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire4497 = ( wire17461  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire17461  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire17461  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire17461  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire4506 = ( (~ preset)  &  wire6005  &  wire17310 ) | ( (~ preset)  &  wire6005  &  (~ wire17388) ) ;
 assign wire4523 = ( (~ preset)  &  wire5945  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5945  &  (~ wire17715) ) ;
 assign wire4524 = ( (~ preset)  &  pdata_12_12_  &  nrq7_2  &  wire17715 ) ;
 assign wire4525 = ( (~ preset)  &  wire5930  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5930  &  (~ wire17712) ) ;
 assign wire4526 = ( (~ preset)  &  pdata_11_11_  &  nrq7_2  &  wire17712 ) ;
 assign wire4527 = ( (~ preset)  &  wire5915  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5915  &  (~ wire17712) ) ;
 assign wire4528 = ( (~ preset)  &  pdata_7_7_  &  nrq7_2  &  wire17712 ) ;
 assign wire4530 = ( (~ preset)  &  wire5900  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5900  &  (~ wire17712) ) ;
 assign wire4531 = ( (~ preset)  &  pdata_0_0_  &  nrq7_2  &  wire17712 ) ;
 assign wire4532 = ( (~ preset)  &  wire5885  &  (~ wire17284) ) | ( (~ preset)  &  wire5885  &  wire18376 ) ;
 assign wire4536 = ( (~ preset)  &  wire5870  &  (~ wire17167) ) | ( (~ preset)  &  wire5870  &  wire17362 ) ;
 assign wire4549 = ( (~ preset)  &  wire5780  &  (~ wire17453) ) | ( (~ preset)  &  wire5780  &  wire18246 ) ;
 assign wire4551 = ( ppeaka_12_12_  &  wire5413 ) | ( ppeaka_12_12_  &  wire17694 ) ;
 assign wire4553 = ( wire11030  &  n_n3081  &  wire4266 ) ;
 assign wire4554 = ( ppeakp_12_12_  &  wire17696 ) | ( ppeakp_12_12_  &  wire17698 ) | ( ppeakp_12_12_  &  wire17703 ) ;
 assign wire4555 = ( ppeakb_12_12_  &  wire4199  &  wire3744 ) ;
 assign wire4557 = ( wire8255  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4558 = ( wire11540  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4560 = ( wire12905  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4561 = ( wire10970  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4562 = ( wire8225  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4563 = ( wire12830  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4564 = ( wire4790  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4566 = ( wire15005  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4567 = ( wire6140  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4568 = ( wire6785  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4569 = ( wire11405  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4571 = ( wire14630  &  wire4226  &  n_n2772 ) ;
 assign wire4572 = ( wire6770  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4575 = ( ppeaks_7_7_  &  wire17660 ) | ( ppeaks_7_7_  &  wire17662 ) ;
 assign wire4576 = ( wire10985  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4577 = ( wire11900  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4578 = ( wire14270  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4579 = ( wire12650  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4581 = ( wire9560  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4582 = ( wire8735  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4583 = ( wire10055  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4584 = ( wire13070  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4585 = ( wire16070  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4586 = ( wire5435  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4587 = ( wire6215  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4590 = ( wire15410  &  wire4226  &  n_n2772 ) ;
 assign wire4591 = ( wire7400  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4593 = ( ppeaks_14_14_  &  wire17660 ) | ( ppeaks_14_14_  &  wire17662 ) ;
 assign wire4596 = ( wire7265  &  wire4199  &  wire3744 ) ;
 assign wire4597 = ( wire5720  &  wire4515 ) | ( wire5720  &  wire17649 ) | ( wire5720  &  wire17650 ) ;
 assign wire4598 = ( wire7550  &  n_n3925  &  wire5513 ) | ( wire7550  &  n_n3925  &  wire5514 ) ;
 assign wire4599 = ( wire6350  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire4601 = ( wire4475  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire4602 = ( wire6410  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire4606 = ( wire11225  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4607 = ( wire14405  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4608 = ( wire10175  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4611 = ( wire5135  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4614 = ( ppeaka_8_8_  &  wire4515 ) | ( ppeaka_8_8_  &  wire4199  &  wire3744 ) ;
 assign wire4615 = ( ppeaka_10_10_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire4616 = ( wire4550  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4617 = ( wire5300  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4618 = ( wire14060  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4620 = ( wire5225  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4621 = ( wire7220  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4622 = ( wire10850  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4624 = ( wire5015  &  wire4226  &  n_n2772 ) ;
 assign wire4626 = ( wire15230  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4628 = ( ppeakb_10_10_  &  wire4515 ) | ( ppeakb_10_10_  &  wire4199  &  wire4211 ) ;
 assign wire4629 = ( (~ preset)  &  wire5675  &  (~ wire17791) ) | ( (~ preset)  &  wire5675  &  wire17843 ) ;
 assign wire4643 = ( (~ preset)  &  wire5630  &  (~ wire17180) ) | ( (~ preset)  &  wire5630  &  wire17232 ) ;
 assign wire4648 = ( (~ preset)  &  wire5600  &  wire17037 ) | ( (~ preset)  &  wire5600  &  (~ wire18025) ) ;
 assign wire4657 = ( (~ preset)  &  wire5555  &  (~ wire17635) ) | ( (~ preset)  &  wire5555  &  wire17986 ) ;
 assign wire4667 = ( wire4278  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4278  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4278  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4278  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire4669 = ( wire4278  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4278  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4278  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4278  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire4673 = ( (~ preset)  &  wire5495  &  wire18311 ) | ( (~ preset)  &  wire5495  &  (~ wire18506) ) ;
 assign wire4680 = ( (~ preset)  &  wire5465  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5465  &  (~ wire17715) ) ;
 assign wire4682 = ( (~ preset)  &  wire5450  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5450  &  (~ wire17712) ) ;
 assign wire4683 = ( wire18501  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire18501  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire18501  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire18501  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire4686 = ( wire4381  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4381  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4381  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4381  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire4688 = ( (~ preset)  &  wire5405  &  (~ wire18285) ) | ( (~ preset)  &  wire5405  &  wire18363 ) ;
 assign wire4690 = ( (~ preset)  &  wire5390  &  (~ wire18285) ) | ( (~ preset)  &  wire5390  &  wire18363 ) ;
 assign wire4693 = ( wire4243  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4243  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4243  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4243  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire4694 = ( (~ preset)  &  wire5360  &  wire18103 ) | ( (~ preset)  &  wire5360  &  (~ wire18168) ) ;
 assign wire4697 = ( wire17461  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire17461  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire17461  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire17461  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire4698 = ( wire5330  &  wire4340 ) ;
 assign wire4702 = ( (~ preset)  &  wire5315  &  wire17310 ) | ( (~ preset)  &  wire5315  &  (~ wire17388) ) ;
 assign wire4710 = ( (~ preset)  &  wire5255  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5255  &  (~ wire17715) ) ;
 assign wire4711 = ( (~ preset)  &  pdata_11_11_  &  nrq7_2  &  wire17715 ) ;
 assign wire4712 = ( (~ preset)  &  wire5240  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5240  &  (~ wire17714) ) ;
 assign wire4713 = ( (~ preset)  &  pdata_5_5_  &  nrq7_2  &  wire17714 ) ;
 assign wire4714 = ( (~ preset)  &  wire5225  &  (~ nrq7_2) ) | ( (~ preset)  &  wire5225  &  (~ wire17712) ) ;
 assign wire4716 = ( (~ preset)  &  pdata_10_10_  &  nrq7_2  &  wire17712 ) ;
 assign wire4717 = ( (~ preset)  &  wire5210  &  (~ wire17284) ) | ( (~ preset)  &  wire5210  &  wire18376 ) ;
 assign wire4719 = ( (~ preset)  &  wire5195  &  (~ wire17284) ) | ( (~ preset)  &  wire5195  &  wire18376 ) ;
 assign wire4725 = ( (~ preset)  &  wire5180  &  (~ wire17167) ) | ( (~ preset)  &  wire5180  &  wire17362 ) ;
 assign wire4734 = ( (~ preset)  &  wire5120  &  (~ wire17102) ) | ( (~ preset)  &  wire5120  &  wire17154 ) ;
 assign wire4736 = ( (~ preset)  &  wire5105  &  (~ wire17102) ) | ( (~ preset)  &  wire5105  &  wire17154 ) ;
 assign wire4738 = ( (~ preset)  &  wire5090  &  (~ wire17453) ) | ( (~ preset)  &  wire5090  &  wire18246 ) ;
 assign wire4741 = ( (~ preset)  &  wire5075  &  (~ wire17453) ) | ( (~ preset)  &  wire5075  &  wire18246 ) ;
 assign wire4742 = ( ppeaka_11_11_  &  wire5413 ) | ( ppeaka_11_11_  &  wire17694 ) ;
 assign wire4744 = ( wire12020  &  n_n3081  &  wire4266 ) ;
 assign wire4746 = ( ppeakp_11_11_  &  wire17696 ) | ( ppeakp_11_11_  &  wire17698 ) | ( ppeakp_11_11_  &  wire17703 ) ;
 assign wire4747 = ( ppeakb_11_11_  &  wire4199  &  wire3744 ) ;
 assign wire4749 = ( wire12245  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire4750 = ( wire11765  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire4751 = ( wire14675  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire4752 = ( wire5615  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4753 = ( wire4865  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4755 = ( wire13790  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4756 = ( wire9785  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4757 = ( wire12350  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4758 = ( wire9380  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4759 = ( wire4715  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4761 = ( wire6875  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4763 = ( wire15035  &  wire4226  &  n_n2772 ) ;
 assign wire4764 = ( wire8015  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4766 = ( ppeaks_4_4_  &  wire17660 ) | ( ppeaks_4_4_  &  wire17662 ) ;
 assign wire4768 = ( wire9185  &  wire4199  &  wire3744 ) ;
 assign wire4770 = ( wire5030  &  wire4515 ) | ( wire5030  &  wire17649 ) | ( wire5030  &  wire17650 ) ;
 assign wire4771 = ( wire13835  &  n_n3925  &  wire5513 ) | ( wire13835  &  n_n3925  &  wire5514 ) ;
 assign wire4773 = ( wire9200  &  wire4199  &  wire3744 ) ;
 assign wire4774 = ( wire5015  &  wire4515 ) | ( wire5015  &  wire17649 ) | ( wire5015  &  wire17650 ) ;
 assign wire4776 = ( wire8180  &  n_n3925  &  wire5513 ) | ( wire8180  &  n_n3925  &  wire5514 ) ;
 assign wire4777 = ( wire7025  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire4779 = ( wire5180  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire4780 = ( wire7055  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire4783 = ( wire10970  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire4785 = ( wire13985  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire4786 = ( wire10460  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4788 = ( wire4430  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4792 = ( ppeaka_7_7_  &  wire4515 ) | ( ppeaka_7_7_  &  wire4199  &  wire3744 ) ;
 assign wire4793 = ( ppeaka_0_0_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire4794 = ( wire15995  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire4795 = ( wire4580  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire4796 = ( wire13655  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire4797 = ( wire5900  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire4798 = ( wire7835  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire4800 = ( wire10550  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire4802 = ( wire4310  &  wire4226  &  n_n2772 ) ;
 assign wire4803 = ( wire15605  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire4806 = ( ppeakb_0_0_  &  wire4515 ) | ( ppeakb_0_0_  &  wire4199  &  wire4211 ) ;
 assign wire4807 = ( (~ preset)  &  wire4970  &  (~ wire17791) ) | ( (~ preset)  &  wire4970  &  wire17843 ) ;
 assign wire4828 = ( (~ preset)  &  wire4895  &  wire17037 ) | ( (~ preset)  &  wire4895  &  (~ wire18025) ) ;
 assign wire4834 = ( wire4880  &  wire4330 ) ;
 assign wire4849 = ( wire11915  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4852 = ( ppeakp_11_11_  &  ndn_latch12_11 ) | ( ppeakp_11_11_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4853 = ( wire16100  &  wire17427  &  (~ wire17648) ) ;
 assign wire4854 = ( wire10130  &  wire17180  &  (~ wire17232) ) ;
 assign wire4855 = ( ppeaka_11_11_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4856 = ( wire13115  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4857 = ( ppeakb_11_11_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4858 = ( wire12050  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4861 = ( ppeakp_12_12_  &  ndn_latch12_11 ) | ( ppeakp_12_12_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4862 = ( wire15755  &  wire17427  &  (~ wire17648) ) ;
 assign wire4863 = ( wire10415  &  wire17180  &  (~ wire17232) ) ;
 assign wire4864 = ( ppeaka_12_12_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4866 = ( wire12395  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4867 = ( ppeakb_12_12_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4868 = ( wire12170  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4870 = ( ppeakp_13_13_  &  ndn_latch12_11 ) | ( ppeakp_13_13_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4871 = ( wire13805  &  wire17427  &  (~ wire17648) ) ;
 assign wire4872 = ( wire10700  &  wire17180  &  (~ wire17232) ) ;
 assign wire4873 = ( ppeaka_13_13_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4875 = ( wire12620  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4876 = ( ppeakb_13_13_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4877 = ( wire12260  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4879 = ( ppeakp_14_14_  &  ndn_latch12_11 ) | ( ppeakp_14_14_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4881 = ( wire13445  &  wire17427  &  (~ wire17648) ) ;
 assign wire4882 = ( wire10985  &  wire17180  &  (~ wire17232) ) ;
 assign wire4883 = ( ppeaka_14_14_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4884 = ( wire15410  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4885 = ( ppeakb_14_14_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4886 = ( wire12470  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4888 = ( ppeakp_15_15_  &  ndn_latch12_11 ) | ( ppeakp_15_15_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4890 = ( wire14615  &  wire17427  &  (~ wire17648) ) ;
 assign wire4891 = ( wire6320  &  wire17180  &  (~ wire17232) ) ;
 assign wire4892 = ( ppeaka_15_15_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4893 = ( wire15050  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4894 = ( ppeakb_15_15_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4902 = ( (~ preset)  &  wire4850  &  (~ wire17635) ) | ( (~ preset)  &  wire4850  &  wire17986 ) ;
 assign wire4916 = ( wire11075  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4918 = ( ppeakp_7_7_  &  ndn_latch12_11 ) | ( ppeakp_7_7_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4920 = ( wire5540  &  wire17427  &  (~ wire17648) ) ;
 assign wire4921 = ( wire8255  &  wire17180  &  (~ wire17232) ) ;
 assign wire4922 = ( ppeaka_7_7_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4923 = ( wire14630  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4924 = ( ppeakb_7_7_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4926 = ( wire11330  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4928 = ( ppeakp_8_8_  &  ndn_latch12_11 ) | ( ppeakp_8_8_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4929 = ( wire11420  &  wire17427  &  (~ wire17648) ) ;
 assign wire4930 = ( wire8915  &  wire17180  &  (~ wire17232) ) ;
 assign wire4931 = ( ppeaka_8_8_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4932 = ( wire13460  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4933 = ( ppeakb_8_8_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4935 = ( wire11570  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4937 = ( ppeakp_9_9_  &  ndn_latch12_11 ) | ( ppeakp_9_9_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4938 = ( wire11645  &  wire17427  &  (~ wire17648) ) ;
 assign wire4939 = ( wire9590  &  wire17180  &  (~ wire17232) ) ;
 assign wire4941 = ( ppeaka_9_9_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4942 = ( wire13820  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4943 = ( ppeakb_9_9_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4944 = ( wire11795  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4946 = ( ppeakp_10_10_  &  ndn_latch12_11 ) | ( ppeakp_10_10_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4947 = ( wire10925  &  wire17427  &  (~ wire17648) ) ;
 assign wire4948 = ( wire9860  &  wire17180  &  (~ wire17232) ) ;
 assign wire4950 = ( ppeaka_10_10_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4951 = ( wire12860  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4952 = ( ppeakb_10_10_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4978 = ( ppeaka_0_0_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4986 = ( wire11555  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4988 = ( ppeakp_0_0_  &  ndn_latch12_11 ) | ( ppeakp_0_0_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4989 = ( wire11630  &  wire17427  &  (~ wire17648) ) ;
 assign wire4990 = ( wire13175  &  wire17180  &  (~ wire17232) ) ;
 assign wire4991 = ( ppeaka_0_0_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire4992 = ( wire12605  &  (~ wire17999)  &  wire18077 ) ;
 assign wire4993 = ( ppeakb_0_0_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire4995 = ( wire11315  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire4997 = ( ppeakp_1_1_  &  ndn_latch12_11 ) | ( ppeakp_1_1_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire4998 = ( wire9485  &  wire17427  &  (~ wire17648) ) ;
 assign wire4999 = ( wire12920  &  wire17180  &  (~ wire17232) ) ;
 assign wire5000 = ( ppeaka_1_1_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5001 = ( wire12380  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5002 = ( ppeakb_1_1_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5003 = ( wire11060  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire5005 = ( ppeakp_2_2_  &  ndn_latch12_11 ) | ( ppeakp_2_2_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire5006 = ( wire7535  &  wire17427  &  (~ wire17648) ) ;
 assign wire5007 = ( wire12680  &  wire17180  &  (~ wire17232) ) ;
 assign wire5008 = ( ppeaka_2_2_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5010 = ( wire13100  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5011 = ( ppeakb_2_2_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5012 = ( wire10790  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire5014 = ( ppeakp_3_3_  &  ndn_latch12_11 ) | ( ppeakp_3_3_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire5016 = ( wire8165  &  wire17427  &  (~ wire17648) ) ;
 assign wire5017 = ( wire12455  &  wire17180  &  (~ wire17232) ) ;
 assign wire5018 = ( ppeaka_3_3_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5019 = ( wire12845  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5020 = ( ppeakb_3_3_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5021 = ( wire10505  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire5023 = ( ppeakp_4_4_  &  ndn_latch12_11 ) | ( ppeakp_4_4_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire5025 = ( wire6230  &  wire17427  &  (~ wire17648) ) ;
 assign wire5026 = ( wire12245  &  wire17180  &  (~ wire17232) ) ;
 assign wire5027 = ( ppeaka_4_4_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5028 = ( wire15035  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5029 = ( ppeakb_4_4_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5031 = ( wire10220  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire5033 = ( ppeakp_5_5_  &  ndn_latch12_11 ) | ( ppeakp_5_5_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire5034 = ( wire6905  &  wire17427  &  (~ wire17648) ) ;
 assign wire5035 = ( wire6995  &  wire17180  &  (~ wire17232) ) ;
 assign wire5036 = ( ppeaka_5_5_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5037 = ( wire15395  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5038 = ( ppeakb_5_5_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5040 = ( wire9950  &  wire17635  &  (~ wire17986)  &  n_n3925 ) ;
 assign wire5042 = ( ppeakp_6_6_  &  ndn_latch12_11 ) | ( ppeakp_6_6_  &  (~ n_n3925)  &  ndn_latch3_9 ) ;
 assign wire5043 = ( wire4835  &  wire17427  &  (~ wire17648) ) ;
 assign wire5044 = ( wire7625  &  wire17180  &  (~ wire17232) ) ;
 assign wire5045 = ( ppeaka_6_6_  &  (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire5046 = ( wire14210  &  (~ wire17999)  &  wire18077 ) ;
 assign wire5047 = ( ppeakb_6_6_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire5057 = ( wire4377  &  n_n2480  &  wire19737  &  wire19520 ) | ( wire4377  &  (~ n_n2480)  &  (~ wire19737)  &  wire19520 ) | ( wire4377  &  (~ n_n2480)  &  wire19737  &  (~ wire19520) ) | ( wire4377  &  n_n2480  &  (~ wire19737)  &  (~ wire19520) ) ;
 assign wire5058 = ( (~ preset)  &  wire4790  &  wire18311 ) | ( (~ preset)  &  wire4790  &  (~ wire18506) ) ;
 assign wire5063 = ( wire4245  &  n_n2474  &  wire19514  &  wire19733 ) | ( wire4245  &  (~ n_n2474)  &  (~ wire19514)  &  wire19733 ) | ( wire4245  &  (~ n_n2474)  &  wire19514  &  (~ wire19733) ) | ( wire4245  &  n_n2474  &  (~ wire19514)  &  (~ wire19733) ) ;
 assign wire5068 = ( wire4245  &  n_n2485  &  wire19466  &  wire19721 ) | ( wire4245  &  (~ n_n2485)  &  (~ wire19466)  &  wire19721 ) | ( wire4245  &  (~ n_n2485)  &  wire19466  &  (~ wire19721) ) | ( wire4245  &  n_n2485  &  (~ wire19466)  &  (~ wire19721) ) ;
 assign wire5073 = ( (~ preset)  &  wire4745  &  (~ nrq7_2) ) | ( (~ preset)  &  wire4745  &  (~ wire17712) ) ;
 assign wire5088 = ( (~ wire5106)  &  (~ wire17836)  &  wire17844 ) ;
 assign wire5091 = ( (~ ppeaka_15_15_)  &  (~ wire4453) ) | ( (~ ppeaka_15_15_)  &  (~ wire5271)  &  (~ wire5272) ) ;
 assign wire5094 = ( wire6755  &  wire18285  &  (~ wire18363) ) ;
 assign wire5096 = ( ppeaka_15_15_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5097 = ( ppeakb_15_15_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5098 = ( wire13550  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5106 = ( (~ ppeaka_14_14_)  &  (~ wire4453) ) | ( (~ ppeaka_14_14_)  &  (~ wire5271)  &  (~ wire5272) ) ;
 assign wire5113 = ( wire9740  &  wire18285  &  (~ wire18363) ) ;
 assign wire5116 = ( ppeaka_13_13_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5117 = ( ppeakb_13_13_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5118 = ( wire15500  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5121 = ( wire6080  &  wire18285  &  (~ wire18363) ) ;
 assign wire5123 = ( ppeaka_14_14_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5124 = ( ppeakb_14_14_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5125 = ( wire15140  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5126 = ( wire4381  &  n_n2483  &  wire19725  &  wire19479 ) | ( wire4381  &  (~ n_n2483)  &  (~ wire19725)  &  wire19479 ) | ( wire4381  &  (~ n_n2483)  &  wire19725  &  (~ wire19479) ) | ( wire4381  &  n_n2483  &  (~ wire19725)  &  (~ wire19479) ) ;
 assign wire5132 = ( (~ preset)  &  wire4700  &  (~ wire18285) ) | ( (~ preset)  &  wire4700  &  wire18363 ) ;
 assign wire5133 = ( wire4306  &  n_n2477  &  wire19735  &  wire19504 ) | ( wire4306  &  (~ n_n2477)  &  (~ wire19735)  &  wire19504 ) | ( wire4306  &  (~ n_n2477)  &  wire19735  &  (~ wire19504) ) | ( wire4306  &  n_n2477  &  (~ wire19735)  &  (~ wire19504) ) ;
 assign wire5139 = ( wire4243  &  n_n2482  &  wire19727  &  wire19456 ) | ( wire4243  &  (~ n_n2482)  &  (~ wire19727)  &  wire19456 ) | ( wire4243  &  (~ n_n2482)  &  wire19727  &  (~ wire19456) ) | ( wire4243  &  n_n2482  &  (~ wire19727)  &  (~ wire19456) ) ;
 assign wire5143 = ( (~ preset)  &  wire4655  &  wire18103 ) | ( (~ preset)  &  wire4655  &  (~ wire18168) ) ;
 assign wire5145 = ( wire4308  &  n_n2476  &  wire19741  &  wire19531 ) | ( wire4308  &  (~ n_n2476)  &  (~ wire19741)  &  wire19531 ) | ( wire4308  &  (~ n_n2476)  &  wire19741  &  (~ wire19531) ) | ( wire4308  &  n_n2476  &  (~ wire19741)  &  (~ wire19531) ) ;
 assign wire5157 = ( n_n2477  &  wire4438  &  wire19735 ) | ( n_n2477  &  wire4438  &  wire19504 ) | ( wire4438  &  wire19735  &  wire19504 ) ;
 assign wire5158 = ( n_n2476  &  wire5273 ) | ( n_n2476  &  wire5274 ) | ( n_n2476  &  wire5275 ) ;
 assign wire5164 = ( n_n2480  &  wire19737  &  wire4450 ) | ( n_n2480  &  wire19520  &  wire4450 ) | ( wire19737  &  wire19520  &  wire4450 ) ;
 assign wire5166 = ( n_n2479  &  wire19743 ) ;
 assign wire5171 = ( n_n2483  &  wire4440  &  wire19725 ) | ( n_n2483  &  wire4440  &  wire19479 ) | ( wire4440  &  wire19725  &  wire19479 ) ;
 assign wire5172 = ( n_n2482  &  wire5286 ) | ( n_n2482  &  wire17748 ) ;
 assign wire5182 = ( wire9725  &  wire18285  &  (~ wire18363) ) ;
 assign wire5184 = ( ppeaka_2_2_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5185 = ( ppeakb_2_2_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5186 = ( wire15515  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5190 = ( (~ ppeaka_3_3_)  &  nrq10_4  &  (~ wire5288) ) | ( (~ ppeaka_3_3_)  &  wire19749  &  (~ wire5288) ) ;
 assign wire5192 = ( wire9995  &  wire18285  &  (~ wire18363) ) ;
 assign wire5194 = ( ppeaka_3_3_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5196 = ( ppeakb_3_3_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5197 = ( wire15860  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5201 = ( wire5375  &  wire18285  &  (~ wire18363) ) ;
 assign wire5203 = ( ppeaka_4_4_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5205 = ( ppeakb_4_4_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5206 = ( wire14765  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5208 = ( wire4670  &  wire18285  &  (~ wire18363) ) ;
 assign wire5211 = ( ppeaka_5_5_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5212 = ( ppeakb_5_5_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5213 = ( wire8330  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5218 = ( wire6740  &  wire18285  &  (~ wire18363) ) ;
 assign wire5221 = ( ppeaka_6_6_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5222 = ( ppeakb_6_6_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5223 = ( wire7685  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5228 = ( wire6065  &  wire18285  &  (~ wire18363) ) ;
 assign wire5230 = ( ppeaka_7_7_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5231 = ( ppeakb_7_7_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5232 = ( wire7055  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5235 = ( wire8000  &  wire18285  &  (~ wire18363) ) ;
 assign wire5237 = ( ppeaka_8_8_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5238 = ( ppeakb_8_8_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5239 = ( wire6410  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5241 = ( (~ ppeaka_8_8_)  &  ppeaka_9_9_  &  (~ wire19743)  &  (~ wire5277) ) ;
 assign wire5243 = ( ppeaka_8_8_  &  (~ ppeaka_9_9_)  &  (~ wire5277) ) | ( (~ ppeaka_9_9_)  &  wire19743  &  (~ wire5277) ) ;
 assign wire5245 = ( wire7370  &  wire18285  &  (~ wire18363) ) ;
 assign wire5247 = ( ppeaka_9_9_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5248 = ( ppeakb_9_9_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5250 = ( wire5720  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5254 = ( wire9305  &  wire18285  &  (~ wire18363) ) ;
 assign wire5257 = ( ppeaka_10_10_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5258 = ( ppeakb_10_10_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5259 = ( wire5015  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5261 = ( wire8645  &  wire18285  &  (~ wire18363) ) ;
 assign wire5263 = ( ppeaka_11_11_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5265 = ( ppeakb_11_11_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5266 = ( wire4295  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5271 = ( (~ wire5273)  &  (~ wire5274)  &  (~ wire5275)  &  wire17756 ) ;
 assign wire5272 = ( (~ nrq10_4)  &  wire19989 ) | ( (~ nrq10_4)  &  (~ wire19743)  &  wire17753 ) ;
 assign wire5273 = ( wire5277  &  wire17754 ) | ( (~ wire19743)  &  wire17753  &  wire17754 ) ;
 assign wire5274 = ( wire19743  &  wire4509  &  (~ wire5277) ) | ( wire4509  &  (~ wire5277)  &  (~ wire17753) ) ;
 assign wire5275 = ( (~ ppeaka_11_11_)  &  (~ wire4455) ) ;
 assign wire5277 = ( (~ nrq7_2)  &  wire19989 ) | ( wire19989  &  (~ wire17710) ) | ( wire19989  &  (~ wire17711) ) ;
 assign wire5283 = ( (~ nrq10_4)  &  (~ wire19749) ) | ( (~ nrq10_4)  &  wire5288 ) ;
 assign wire5286 = ( nrq10_4  &  wire4508  &  (~ wire5288) ) | ( wire19749  &  wire4508  &  (~ wire5288) ) ;
 assign wire5287 = ( (~ ppeaka_5_5_)  &  (~ wire4452) ) ;
 assign wire5288 = ( (~ wire5290)  &  (~ wire5291)  &  (~ wire5292)  &  wire17745 ) ;
 assign wire5289 = ( (~ nrq7_2)  &  (~ wire19749) ) | ( (~ wire19749)  &  (~ wire17710) ) | ( (~ wire19749)  &  (~ wire17711) ) ;
 assign wire5290 = ( (~ wire4265)  &  (~ wire17719)  &  (~ wire17722)  &  wire17743 ) ;
 assign wire5291 = ( wire4265  &  wire4507 ) | ( wire4507  &  wire17719 ) | ( wire4507  &  wire17722 ) ;
 assign wire5292 = ( (~ ppeaka_2_2_)  &  (~ wire4457) ) ;
 assign wire5295 = ( wire10010  &  wire18285  &  (~ wire18363) ) ;
 assign wire5297 = ( ppeaka_12_12_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5298 = ( ppeakb_12_12_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5299 = ( wire15845  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5313 = ( ppeaka_0_0_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5320 = ( wire8630  &  wire18285  &  (~ wire18363) ) ;
 assign wire5322 = ( ppeaka_0_0_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5323 = ( ppeakb_0_0_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5325 = ( wire4310  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5327 = ( wire9290  &  wire18285  &  (~ wire18363) ) ;
 assign wire5329 = ( ppeaka_1_1_  &  (~ wire18285)  &  nrq7_2  &  wire3723 ) ;
 assign wire5331 = ( ppeakb_1_1_  &  nrq7_2  &  wire17710  &  wire17711 ) ;
 assign wire5332 = ( wire5030  &  (~ wire18506)  &  nrq7_2  &  wire3744 ) ;
 assign wire5334 = ( (~ preset)  &  wire4610  &  wire17310 ) | ( (~ preset)  &  wire4610  &  (~ wire17388) ) ;
 assign wire5344 = ( (~ preset)  &  wire4550  &  (~ nrq7_2) ) | ( (~ preset)  &  wire4550  &  (~ wire17715) ) ;
 assign wire5346 = ( (~ preset)  &  pdata_10_10_  &  nrq7_2  &  wire17715 ) ;
 assign wire5349 = ( (~ preset)  &  wire4535  &  (~ nrq7_2) ) | ( (~ preset)  &  wire4535  &  (~ wire17714) ) ;
 assign wire5350 = ( (~ preset)  &  pdata_15_15_  &  nrq7_2  &  wire17714 ) ;
 assign wire5353 = ( (~ preset)  &  wire4520  &  (~ nrq7_2) ) | ( (~ preset)  &  wire4520  &  (~ wire17712) ) ;
 assign wire5355 = ( (~ preset)  &  pdata_9_9_  &  nrq7_2  &  wire17712 ) ;
 assign wire5358 = ( (~ preset)  &  wire4505  &  (~ wire17284) ) | ( (~ preset)  &  wire4505  &  wire18376 ) ;
 assign wire5363 = ( (~ preset)  &  wire4490  &  (~ wire17284) ) | ( (~ preset)  &  wire4490  &  wire18376 ) ;
 assign wire5368 = ( (~ preset)  &  wire4475  &  (~ wire17167) ) | ( (~ preset)  &  wire4475  &  wire17362 ) ;
 assign wire5385 = ( (~ preset)  &  wire4415  &  (~ wire17102) ) | ( (~ preset)  &  wire4415  &  wire17154 ) ;
 assign wire5389 = ( (~ preset)  &  wire4400  &  (~ wire17102) ) | ( (~ preset)  &  wire4400  &  wire17154 ) ;
 assign wire5398 = ( (~ preset)  &  wire4370  &  (~ wire17453) ) | ( (~ preset)  &  wire4370  &  wire18246 ) ;
 assign wire5403 = ( (~ preset)  &  wire4355  &  (~ wire17453) ) | ( (~ preset)  &  wire4355  &  wire18246 ) ;
 assign wire5407 = ( ppeaka_10_10_  &  wire5413 ) | ( ppeaka_10_10_  &  wire17694 ) ;
 assign wire5409 = ( wire12140  &  n_n3081  &  wire4266 ) ;
 assign wire5410 = ( ppeakp_10_10_  &  wire17696 ) | ( ppeakp_10_10_  &  wire17698 ) | ( ppeakp_10_10_  &  wire17703 ) ;
 assign wire5411 = ( ppeakb_10_10_  &  wire4199  &  wire3744 ) ;
 assign wire5413 = ( wire4199  &  wire3720  &  wire4024 ) ;
 assign wire5418 = ( wire4199  &  wire3720  &  (~ wire4024) ) ;
 assign wire5426 = ( wire6995  &  wire4199  &  wire3754  &  n_n2772 ) ;
 assign wire5427 = ( wire11885  &  n_n2772  &  n_n3081  &  wire4266 ) ;
 assign wire5428 = ( wire13505  &  wire4199  &  wire3750  &  n_n2772 ) ;
 assign wire5430 = ( wire11465  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire5431 = ( wire9545  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire5432 = ( wire13430  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire5433 = ( wire6185  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire5434 = ( wire13055  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire5436 = ( wire7445  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire5437 = ( wire5420  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire5438 = ( wire10895  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire5440 = ( wire15395  &  wire4226  &  n_n2772 ) ;
 assign wire5441 = ( wire10280  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire5443 = ( ppeaks_5_5_  &  wire17660 ) | ( ppeaks_5_5_  &  wire17662 ) ;
 assign wire5451 = ( wire8525  &  wire4199  &  wire3744 ) ;
 assign wire5452 = ( wire4310  &  wire4515 ) | ( wire4310  &  wire17649 ) | ( wire4310  &  wire17650 ) ;
 assign wire5453 = ( wire14225  &  n_n3925  &  wire5513 ) | ( wire14225  &  n_n3925  &  wire5514 ) ;
 assign wire5455 = ( wire8540  &  wire4199  &  wire3744 ) ;
 assign wire5456 = ( wire4295  &  wire4515 ) | ( wire4295  &  wire17649 ) | ( wire4295  &  wire17650 ) ;
 assign wire5457 = ( wire8825  &  n_n3925  &  wire5513 ) | ( wire8825  &  n_n3925  &  wire5514 ) ;
 assign wire5464 = ( wire4955  &  wire4199  &  wire3746  &  n_n2772 ) ;
 assign wire5467 = ( wire5870  &  wire4199  &  wire3727  &  n_n2772 ) ;
 assign wire5468 = ( wire7685  &  wire4199  &  n_n2772  &  wire4207 ) ;
 assign wire5471 = ( wire11690  &  wire4199  &  wire3715  &  n_n2772 ) ;
 assign wire5472 = ( wire15200  &  wire4199  &  wire3740  &  n_n2772 ) ;
 assign wire5473 = ( wire10745  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire5476 = ( wire15935  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire5479 = ( ppeaka_6_6_  &  wire4515 ) | ( ppeaka_6_6_  &  wire4199  &  wire3744 ) ;
 assign wire5483 = ( ppeaka_1_1_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire5484 = ( wire15650  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire5485 = ( wire5285  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire5486 = ( wire13310  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire5487 = ( wire13295  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire5488 = ( wire8480  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire5490 = ( wire14510  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire5492 = ( wire5030  &  wire4226  &  n_n2772 ) ;
 assign wire5493 = ( wire5150  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire5496 = ( ppeakb_1_1_  &  wire4515 ) | ( ppeakb_1_1_  &  wire4199  &  wire4211 ) ;
 assign wire5497 = ( ppeaka_12_12_  &  wire4199  &  n_n2772  &  wire4224 ) ;
 assign wire5498 = ( wire5945  &  wire4199  &  wire3747  &  n_n2772 ) ;
 assign wire5499 = ( wire9230  &  wire4199  &  wire3744  &  n_n2772 ) ;
 assign wire5500 = ( wire13325  &  wire4199  &  n_n2772  &  wire3720 ) ;
 assign wire5501 = ( wire15260  &  wire4199  &  wire3711  &  n_n2772 ) ;
 assign wire5502 = ( wire8495  &  wire4199  &  wire3738  &  n_n2772 ) ;
 assign wire5503 = ( wire7955  &  wire4199  &  wire3718  &  n_n2772 ) ;
 assign wire5506 = ( wire15845  &  wire4226  &  n_n2772 ) ;
 assign wire5507 = ( wire6545  &  wire4199  &  wire3723  &  n_n2772 ) ;
 assign wire5509 = ( ppeakb_12_12_  &  wire4515 ) | ( ppeakb_12_12_  &  wire4199  &  wire4211 ) ;
 assign wire5513 = ( (~ preset)  &  pdn  &  (~ wire17089)  &  (~ wire4202) ) ;
 assign wire5514 = ( (~ preset)  &  (~ wire17596)  &  wire4513 ) ;
 assign wire5520 = ( nrq1_4  &  wire17610 ) | ( (~ wire17596)  &  wire4513  &  wire17610 ) ;
 assign wire5522 = ( pdn  &  (~ wire17089)  &  wire4202 ) ;
 assign wire5528 = ( (~ wire17856)  &  wire18207 ) ;
 assign wire5582 = ( (~ preset)  &  ndout  &  (~ wire17791) ) | ( (~ preset)  &  ndout  &  wire17843 ) ;
 assign wire17517 = ( (~ ppeaki_6_6_)  &  (~ ppeaki_7_7_)  &  (~ wire17752) ) ;
 assign wire17519 = ( (~ wire17544)  &  wire17713  &  wire17752 ) ;
 assign wire17520 = ( wire17674  &  wire17609 ) ;
 assign wire17521 = ( wire17544  &  wire17713  &  wire17752 ) ;
 assign wire17522 = ( ppeaki_6_6_  &  (~ ppeaki_4_4_) ) ;
 assign wire17523 = ( (~ wire17713)  &  (~ wire17674) ) ;
 assign wire17524 = ( (~ ppeaki_5_5_)  &  ppeaki_4_4_ ) ;
 assign wire17525 = ( wire17713  &  wire17609 ) ;
 assign wire17527 = ( (~ wire17609)  &  wire17674  &  wire17713 ) ;
 assign wire17528 = ( ppeaki_6_6_  &  (~ ppeaki_7_7_)  &  (~ wire17752) ) ;
 assign wire17529 = ( (~ wire17713)  &  wire17674 ) ;
 assign wire17530 = ( (~ ppeaki_5_5_)  &  (~ ppeaki_4_4_) ) ;
 assign wire17532 = ( (~ wire17713)  &  wire17609 ) ;
 assign wire17533 = ( wire17674  &  wire17609 ) ;
 assign wire17534 = ( wire17544  &  (~ wire17713)  &  wire17752 ) ;
 assign wire17535 = ( (~ ppeaki_5_5_)  &  (~ ppeaki_4_4_) ) ;
 assign wire17536 = ( (~ wire17713)  &  (~ wire17609) ) ;
 assign wire17537 = ( ppeaki_6_6_  &  ppeaki_4_4_ ) ;
 assign wire17538 = ( wire17713  &  (~ wire17674) ) ;
 assign wire17540 = ( (~ ppeaki_5_5_)  &  ppeaki_4_4_ ) ;
 assign wire17541 = ( wire17713  &  (~ wire17609) ) ;
 assign wire17542 = ( ppeaki_6_6_  &  (~ ppeaki_7_7_)  &  (~ wire17752) ) ;
 assign wire17543 = ( wire17713  &  wire17674 ) ;
 assign wire17545 = ( (~ wire17609)  &  wire17674  &  (~ wire17713) ) ;
 assign wire17546 = ( (~ ppeaki_6_6_)  &  (~ ppeaki_7_7_)  &  (~ wire17752) ) ;
 assign wire17547 = ( (~ wire17544)  &  (~ wire17713)  &  wire17752 ) ;
 assign wire17555 = ( wire3784 ) | ( n_n2319 ) ;
 assign wire17556 = ( n_n2326 ) | ( n_n2314 ) | ( n_n2325 ) | ( n_n2316 ) ;
 assign wire17557 = ( n_n2318 ) | ( n_n2323 ) | ( n_n2317 ) | ( n_n2315 ) ;
 assign wire17558 = ( n_n2321 ) | ( n_n2324 ) | ( n_n2320 ) | ( n_n2322 ) ;
 assign wire17562 = ( wire17596  &  (~ wire17661)  &  (~ wire18597)  &  (~ wire18636) ) ;
 assign wire17564 = ( (~ n_n2333)  &  n_n3714  &  wire17562 ) | ( (~ n_n2333)  &  n_n3713  &  wire17562 ) ;
 assign wire17566 = ( wire17596  &  (~ wire17661)  &  (~ wire18597)  &  (~ wire18636) ) ;
 assign wire17568 = ( n_n3714  &  wire17566 ) | ( n_n3713  &  wire17566 ) ;
 assign wire17572 = ( wire17596  &  (~ wire17661)  &  (~ wire18597)  &  (~ wire18636) ) ;
 assign wire17574 = ( (~ n_n2333)  &  n_n3712  &  wire17572 ) | ( (~ n_n2333)  &  n_n3711  &  wire17572 ) ;
 assign wire17576 = ( wire17596  &  (~ wire17661)  &  (~ wire18597)  &  (~ wire18636) ) ;
 assign wire17577 = ( n_n3712  &  wire17576 ) | ( n_n3711  &  wire17576 ) ;
 assign wire17580 = ( (~ n_n2344)  &  (~ n_n2333)  &  wire17568 ) | ( (~ n_n2344)  &  (~ n_n2333)  &  wire17577 ) ;
 assign wire17582 = ( wire17596  &  (~ wire17661)  &  (~ wire18597) ) ;
 assign wire17593 = ( (~ wire10805)  &  (~ wire10820)  &  (~ wire18207) ) ;
 assign wire17594 = ( (~ wire11090)  &  (~ wire11345)  &  (~ wire11585)  &  (~ wire11600) ) ;
 assign wire17595 = ( (~ wire11810)  &  (~ wire11930)  &  (~ wire12065)  &  (~ wire12080) ) ;
 assign wire17597 = ( (~ wire12185)  &  (~ wire12200)  &  (~ wire12275)  &  (~ wire12485) ) ;
 assign wire17599 = ( wire17595  &  wire17594 ) ;
 assign wire17600 = ( (~ wire12695)  &  (~ wire12935)  &  wire17593  &  wire17597 ) ;
 assign wire17601 = ( wire17986  &  (~ wire17804) ) ;
 assign wire17602 = ( (~ wire17674)  &  (~ wire17609) ) ;
 assign wire17603 = ( (~ wire17544)  &  wire17713  &  wire17752 ) ;
 assign wire17605 = ( (~ ppeaki_6_6_)  &  ppeaki_4_4_ ) ;
 assign wire17606 = ( (~ wire17674)  &  (~ wire17609) ) ;
 assign wire17607 = ( (~ wire17544)  &  (~ wire17713)  &  wire17752 ) ;
 assign wire17608 = ( (~ ppeaki_6_6_)  &  (~ ppeaki_4_4_) ) ;
 assign wire17610 = ( (~ pirq_0_0_)  &  (~ preset)  &  (~ wire18064) ) | ( (~ pirq_0_0_)  &  (~ preset)  &  (~ wire18129) ) | ( (~ preset)  &  wire18064  &  (~ wire18129) ) ;
 assign wire17615 = ( wire5507 ) | ( wire15545  &  wire4269 ) ;
 assign wire17616 = ( wire5497 ) | ( wire5506 ) | ( wire6470  &  wire4260 ) ;
 assign wire17617 = ( wire5498 ) | ( wire5499 ) | ( wire5500 ) | ( wire5501 ) ;
 assign wire17621 = ( wire5502 ) | ( wire5503 ) | ( wire5509 ) | ( wire17617 ) ;
 assign wire17626 = ( wire5493 ) | ( wire9065  &  wire4269 ) ;
 assign wire17627 = ( wire5483 ) | ( wire5492 ) | ( wire5075  &  wire4260 ) ;
 assign wire17628 = ( wire5484 ) | ( wire5485 ) | ( wire5486 ) | ( wire5487 ) ;
 assign wire17631 = ( wire5488 ) | ( wire5490 ) | ( wire5496 ) | ( wire17628 ) ;
 assign wire17638 = ( wire5476 ) | ( wire5473 ) ;
 assign wire17639 = ( ppeakp_6_6_  &  wire4298 ) | ( ppeaka_7_7_  &  wire4392 ) ;
 assign wire17640 = ( (~ ppeaka_6_6_)  &  wire4260 ) | ( wire12560  &  wire4269 ) ;
 assign wire17641 = ( wire5464 ) | ( (~ ppeakb_6_6_)  &  wire4260 ) | ( ppeakb_6_6_  &  wire4397 ) ;
 assign wire17642 = ( wire5467 ) | ( wire5468 ) | ( wire5471 ) | ( wire5472 ) ;
 assign wire17647 = ( wire5479 ) | ( wire17638 ) | ( wire17639 ) | ( wire17640 ) ;
 assign wire17649 = ( wire4199  &  wire4219 ) | ( wire4199  &  wire4225 ) ;
 assign wire17650 = ( wire4199  &  wire3750 ) | ( wire4199  &  wire4212 ) ;
 assign wire17652 = ( wire5457 ) | ( wire7655  &  wire4199  &  wire3754 ) ;
 assign wire17654 = ( wire5453 ) | ( wire7640  &  wire4199  &  wire3754 ) ;
 assign wire17657 = ( (~ preset)  &  pdn  &  (~ wire17089)  &  (~ n_n3081) ) ;
 assign wire17658 = ( (~ wire5528)  &  (~ wire17599)  &  wire17657 ) | ( (~ wire5528)  &  (~ wire17600)  &  wire17657 ) ;
 assign wire17659 = ( (~ n_n3925)  &  wire5514 ) | ( (~ n_n3925)  &  (~ wire4202)  &  wire4266 ) ;
 assign wire17660 = ( n_n2772  &  wire17658 ) | ( n_n2772  &  wire17659 ) ;
 assign wire17662 = ( (~ preset)  &  (~ ndn7_2)  &  (~ wire4205) ) | ( (~ preset)  &  ndn7_2  &  wire4211 ) ;
 assign wire17668 = ( wire5438 ) | ( wire5437 ) ;
 assign wire17670 = ( wire5427 ) | ( wire5440 ) | ( wire5441 ) ;
 assign wire17671 = ( wire13700  &  wire4260 ) | ( wire14555  &  wire4269 ) ;
 assign wire17672 = ( wire5426 ) | ( wire5428 ) | ( wire5430 ) | ( wire5431 ) ;
 assign wire17673 = ( wire5432 ) | ( wire5433 ) | ( wire5434 ) | ( wire5436 ) ;
 assign wire17678 = ( wire5443 ) | ( wire17668 ) | ( wire17670 ) | ( wire17671 ) ;
 assign wire17688 = ( ppeakb_7_7_ ) | ( ppeakb_14_14_ ) | ( ppeakb_10_10_ ) | ( ppeakb_8_8_ ) ;
 assign wire17689 = ( ppeakb_9_9_ ) | ( ppeakb_15_15_ ) | ( ppeakb_11_11_ ) | ( ppeakb_0_0_ ) ;
 assign wire17690 = ( ppeakb_1_1_ ) | ( ppeakb_12_12_ ) | ( ppeakb_2_2_ ) | ( ppeakb_3_3_ ) ;
 assign wire17691 = ( ppeakb_13_13_ ) | ( ppeakb_4_4_ ) | ( ppeakb_5_5_ ) | ( ppeakb_6_6_ ) ;
 assign wire17694 = ( wire4199  &  wire3711 ) | ( wire4199  &  n_n2333 ) ;
 assign wire17695 = ( (~ preset_0_0_)  &  (~ wire17024)  &  wire4266 ) | ( wire17024  &  (~ wire18545)  &  wire4266 ) ;
 assign wire17696 = ( wire4199  &  wire3715 ) | ( wire4202  &  wire17695 ) ;
 assign wire17698 = ( wire4199  &  wire4207 ) | ( wire4199  &  wire4219 ) ;
 assign wire17699 = ( wire4199  &  wire4204 ) | ( wire4199  &  wire4208 ) ;
 assign wire17703 = ( wire5418 ) | ( wire17699 ) | ( (~ preset)  &  (~ n_n2772) ) ;
 assign wire17704 = ( wire5409 ) | ( wire4850  &  wire5513 ) | ( wire4850  &  wire5514 ) ;
 assign wire17705 = ( wire17704 ) | ( wire6965  &  wire4199  &  wire3740 ) ;
 assign wire17709 = ( n_n2344  &  (~ wire18610) ) ;
 assign wire17710 = ( (~ wire18610)  &  n_n2344  &  (~ nsl8_2) ) ;
 assign wire17711 = ( wire3770  &  (~ wire18168) ) ;
 assign wire17712 = ( wire3711  &  (~ wire18493) ) ;
 assign wire17714 = ( wire3720  &  (~ wire16920) ) ;
 assign wire17715 = ( wire3747  &  (~ wire17297) ) ;
 assign wire17716 = ( wire3775  &  (~ wire17453) ) ;
 assign wire17717 = ( nrq7_2  &  wire17715 ) | ( (~ wire16920)  &  nrq7_2  &  wire3720 ) ;
 assign wire17718 = ( nrq7_2  &  wire17712 ) | ( nrq7_2  &  wire17710  &  wire17716 ) ;
 assign wire17719 = ( ndn_latch24_2 ) | ( (~ wire17284)  &  nrq7_2  &  wire3738 ) ;
 assign wire17720 = ( wire18285  &  (~ wire18363) ) | ( (~ wire18311)  &  wire18506 ) ;
 assign wire17722 = ( nrq23_3 ) | ( nrq14_3 ) | ( wire5313 ) | ( wire17720 ) ;
 assign wire17724 = ( wire5320 ) | ( wire10025  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17727 = ( wire5322 ) | ( wire5323 ) | ( wire5325 ) | ( wire17724 ) ;
 assign wire17728 = ( wire5327 ) | ( wire10310  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17731 = ( wire5329 ) | ( wire5331 ) | ( wire5332 ) | ( wire17728 ) ;
 assign wire17738 = ( wire5295 ) | ( wire6860  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17742 = ( wire5297 ) | ( wire5298 ) | ( wire5299 ) | ( wire17738 ) ;
 assign wire17743 = ( (~ wire4507)  &  (~ ppeaka_1_1_) ) ;
 assign wire17745 = ( (~ ppeaka_3_3_)  &  (~ ppeaka_2_2_) ) ;
 assign wire17746 = ( (~ wire4508)  &  (~ ppeaka_4_4_) ) ;
 assign wire17748 = ( wire5287 ) | ( wire5288  &  wire17746 ) | ( wire5289  &  wire17746 ) ;
 assign wire17749 = ( (~ ppeaka_6_6_)  &  (~ ppeaka_5_5_) ) ;
 assign wire17753 = ( (~ ppeaka_9_9_)  &  (~ ppeaka_8_8_) ) ;
 assign wire17754 = ( (~ wire4509)  &  (~ ppeaka_10_10_) ) ;
 assign wire17756 = ( (~ ppeaka_12_12_)  &  (~ ppeaka_11_11_) ) ;
 assign wire17757 = ( (~ ppeaka_10_10_)  &  (~ ppeaka_11_11_)  &  wire18861 ) | ( (~ ppeaka_11_11_)  &  (~ nrq10_4)  &  wire18861 ) ;
 assign wire17758 = ( (~ nrq10_4)  &  (~ wire18861) ) | ( nrq10_4  &  (~ wire5271)  &  wire17757 ) | ( (~ wire18861)  &  (~ wire5271)  &  wire17757 ) ;
 assign wire17759 = ( wire5182 ) | ( wire4760  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17763 = ( wire5184 ) | ( wire5185 ) | ( wire5186 ) | ( wire17759 ) ;
 assign wire17764 = ( wire5192 ) | ( wire6845  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17768 = ( wire5194 ) | ( wire5196 ) | ( wire5197 ) | ( wire17764 ) ;
 assign wire17769 = ( (~ ppeaka_1_1_)  &  (~ ppeaka_2_2_)  &  (~ n_n2471) ) | ( (~ ppeaka_2_2_)  &  (~ nrq10_4)  &  (~ n_n2471) ) ;
 assign wire17770 = ( (~ nrq10_4)  &  wire19749  &  (~ wire5288) ) | ( nrq10_4  &  (~ wire5288)  &  wire17769 ) | ( wire19749  &  (~ wire5288)  &  wire17769 ) ;
 assign wire17771 = ( wire5201 ) | ( wire6170  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17774 = ( wire5203 ) | ( wire5205 ) | ( wire5206 ) | ( wire17771 ) ;
 assign wire17776 = ( wire5208 ) | ( wire8105  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17780 = ( wire5211 ) | ( wire5212 ) | ( wire5213 ) | ( wire17776 ) ;
 assign wire17781 = ( wire5218 ) | ( wire7475  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17784 = ( wire5221 ) | ( wire5222 ) | ( wire5223 ) | ( wire17781 ) ;
 assign wire17785 = ( (~ ppeaka_5_5_)  &  (~ wire5286)  &  (~ wire17748) ) ;
 assign wire17787 = ( wire5228 ) | ( wire9410  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17792 = ( wire5230 ) | ( wire5231 ) | ( wire5232 ) | ( wire17787 ) ;
 assign wire17793 = ( wire5235 ) | ( wire8750  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17796 = ( wire5237 ) | ( wire5238 ) | ( wire5239 ) | ( wire17793 ) ;
 assign wire17797 = ( wire5245 ) | ( wire10040  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17801 = ( wire5247 ) | ( wire5248 ) | ( wire5250 ) | ( wire17797 ) ;
 assign wire17805 = ( wire5254 ) | ( wire9770  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17808 = ( wire5257 ) | ( wire5258 ) | ( wire5259 ) | ( wire17805 ) ;
 assign wire17809 = ( wire5261 ) | ( wire10595  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17813 = ( wire5263 ) | ( wire5265 ) | ( wire5266 ) | ( wire17809 ) ;
 assign wire17826 = ( wire5113 ) | ( wire4775  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17829 = ( wire5116 ) | ( wire5117 ) | ( wire5118 ) | ( wire17826 ) ;
 assign wire17830 = ( wire5121 ) | ( wire5480  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17833 = ( wire5123 ) | ( wire5124 ) | ( wire5125 ) | ( wire17830 ) ;
 assign wire17834 = ( (~ ppeaka_13_13_)  &  ppeaka_14_14_ ) ;
 assign wire17836 = ( (~ nrq10_4)  &  (~ wire18861)  &  (~ wire5271) ) | ( nrq10_4  &  wire5271  &  wire17834 ) ;
 assign wire17837 = ( wire5094 ) | ( wire8765  &  (~ wire18311)  &  wire18506 ) ;
 assign wire17841 = ( wire5096 ) | ( wire5097 ) | ( wire5098 ) | ( wire17837 ) ;
 assign wire17842 = ( ppeaka_15_15_  &  (~ ppeaka_14_14_) ) ;
 assign wire17844 = ( nrq7_2  &  wire17710  &  wire17711  &  wire17842 ) ;
 assign wire17845 = ( (~ ppeaka_15_15_)  &  ppeaka_14_14_ ) ;
 assign wire17846 = ( nrq10_4  &  wire17845 ) | ( (~ nrq10_4)  &  (~ wire18861)  &  (~ wire5271) ) ;
 assign wire17865 = ( nrq4_2 ) | ( (~ wire18025)  &  nrq7_2  &  wire3740 ) ;
 assign wire17868 = ( wire5043 ) | ( wire5044 ) | ( wire5046 ) ;
 assign wire17871 = ( wire5040 ) | ( wire5042 ) | ( wire17868 ) ;
 assign wire17873 = ( wire5045 ) | ( wire5047 ) | ( wire17871 ) ;
 assign wire17875 = ( wire5034 ) | ( wire5035 ) | ( wire5037 ) ;
 assign wire17877 = ( wire5031 ) | ( wire5033 ) | ( wire17875 ) ;
 assign wire17880 = ( wire5036 ) | ( wire5038 ) | ( wire17877 ) ;
 assign wire17883 = ( wire5025 ) | ( wire5026 ) | ( wire5028 ) ;
 assign wire17885 = ( wire5021 ) | ( wire5023 ) | ( wire17883 ) ;
 assign wire17887 = ( wire5027 ) | ( wire5029 ) | ( wire17885 ) ;
 assign wire17889 = ( wire5016 ) | ( wire5017 ) | ( wire5019 ) ;
 assign wire17891 = ( wire5012 ) | ( wire5014 ) | ( wire17889 ) ;
 assign wire17894 = ( wire5018 ) | ( wire5020 ) | ( wire17891 ) ;
 assign wire17896 = ( wire5006 ) | ( wire5007 ) | ( wire5010 ) ;
 assign wire17898 = ( wire5003 ) | ( wire5005 ) | ( wire17896 ) ;
 assign wire17900 = ( wire5008 ) | ( wire5011 ) | ( wire17898 ) ;
 assign wire17901 = ( wire17635  &  (~ wire17986) ) | ( (~ wire17037)  &  wire18025 ) ;
 assign wire17902 = ( wire17427  &  (~ wire17648) ) | ( (~ wire17999)  &  wire18077 ) ;
 assign wire17903 = ( wire17902 ) | ( wire17901 ) ;
 assign wire17904 = ( wire17903 ) | ( (~ wire17245)  &  nrq7_2  &  wire3746 ) ;
 assign wire17906 = ( wire17904 ) | ( wire4978 ) ;
 assign wire17909 = ( wire4989 ) | ( wire4990 ) | ( wire4992 ) ;
 assign wire17911 = ( wire4986 ) | ( wire4988 ) | ( wire17909 ) ;
 assign wire17913 = ( wire4991 ) | ( wire4993 ) | ( wire17911 ) ;
 assign wire17915 = ( wire4998 ) | ( wire4999 ) | ( wire5001 ) ;
 assign wire17917 = ( wire4995 ) | ( wire4997 ) | ( wire17915 ) ;
 assign wire17920 = ( wire5000 ) | ( wire5002 ) | ( wire17917 ) ;
 assign wire17924 = ( ppeaks_0_0_  &  wire4273 ) | ( wire4273  &  wire17913 ) | ( wire17906  &  wire17913 ) ;
 assign wire17925 = ( ppeaka_2_2_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17926 = ( ppeaka_3_3_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17927 = ( ppeaka_4_4_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17928 = ( ppeaka_5_5_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17932 = ( ppeaka_6_6_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17937 = ( wire4947 ) | ( wire4948 ) | ( wire4951 ) ;
 assign wire17939 = ( wire4944 ) | ( wire4946 ) | ( wire17937 ) ;
 assign wire17941 = ( wire4950 ) | ( wire4952 ) | ( wire17939 ) ;
 assign wire17943 = ( wire4938 ) | ( wire4939 ) | ( wire4942 ) ;
 assign wire17946 = ( wire4935 ) | ( wire4937 ) | ( wire17943 ) ;
 assign wire17949 = ( wire4941 ) | ( wire4943 ) | ( wire17946 ) ;
 assign wire17951 = ( wire4929 ) | ( wire4930 ) | ( wire4932 ) ;
 assign wire17953 = ( wire4926 ) | ( wire4928 ) | ( wire17951 ) ;
 assign wire17955 = ( wire4931 ) | ( wire4933 ) | ( wire17953 ) ;
 assign wire17958 = ( wire4920 ) | ( wire4921 ) | ( wire4923 ) ;
 assign wire17961 = ( wire4916 ) | ( wire4918 ) | ( wire17958 ) ;
 assign wire17963 = ( wire4922 ) | ( wire4924 ) | ( wire17961 ) ;
 assign wire17964 = ( ppeaka_7_7_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17965 = ( ppeaka_8_8_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17966 = ( ppeaka_9_9_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17969 = ( ppeaka_10_10_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire17979 = ( wire4890 ) | ( wire4891 ) | ( wire4893 ) ;
 assign wire17981 = ( wire4886 ) | ( wire4888 ) | ( wire17979 ) ;
 assign wire17984 = ( wire4892 ) | ( wire4894 ) | ( wire17981 ) ;
 assign wire17987 = ( wire4881 ) | ( wire4882 ) | ( wire4884 ) ;
 assign wire17989 = ( wire4877 ) | ( wire4879 ) | ( wire17987 ) ;
 assign wire17991 = ( wire4883 ) | ( wire4885 ) | ( wire17989 ) ;
 assign wire17993 = ( wire4871 ) | ( wire4872 ) | ( wire4875 ) ;
 assign wire17996 = ( wire4868 ) | ( wire4870 ) | ( wire17993 ) ;
 assign wire17998 = ( wire4873 ) | ( wire4876 ) | ( wire17996 ) ;
 assign wire18001 = ( wire4862 ) | ( wire4863 ) | ( wire4866 ) ;
 assign wire18003 = ( wire4858 ) | ( wire4861 ) | ( wire18001 ) ;
 assign wire18005 = ( wire4864 ) | ( wire4867 ) | ( wire18003 ) ;
 assign wire18008 = ( wire4853 ) | ( wire4854 ) | ( wire4856 ) ;
 assign wire18010 = ( wire4849 ) | ( wire4852 ) | ( wire18008 ) ;
 assign wire18013 = ( wire4855 ) | ( wire4857 ) | ( wire18010 ) ;
 assign wire18014 = ( ppeaka_11_11_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire18015 = ( ppeaka_12_12_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire18016 = ( ppeaka_13_13_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire18017 = ( ppeaka_14_14_  &  (~ wire16933)  &  nrq7_2  &  wire3718 ) ;
 assign wire18037 = ( wire4803 ) | ( wire8405  &  wire4269 ) ;
 assign wire18039 = ( wire4793 ) | ( wire4802 ) | ( wire4355  &  wire4260 ) ;
 assign wire18040 = ( wire4794 ) | ( wire4795 ) | ( wire4796 ) | ( wire4797 ) ;
 assign wire18043 = ( wire4798 ) | ( wire4800 ) | ( wire4806 ) | ( wire18040 ) ;
 assign wire18047 = ( wire4788 ) | ( wire4786 ) ;
 assign wire18049 = ( ppeakp_7_7_  &  wire4298 ) | ( ppeaka_8_8_  &  wire4392 ) ;
 assign wire18050 = ( (~ ppeaka_7_7_)  &  wire4260 ) | ( wire12335  &  wire4269 ) ;
 assign wire18051 = ( wire4777 ) | ( (~ ppeakb_7_7_)  &  wire4260 ) | ( ppeakb_7_7_  &  wire4397 ) ;
 assign wire18052 = ( wire4779 ) | ( wire4780 ) | ( wire4783 ) | ( wire4785 ) ;
 assign wire18056 = ( wire4792 ) | ( wire18047 ) | ( wire18049 ) | ( wire18050 ) ;
 assign wire18057 = ( wire4776 ) | ( wire9620  &  wire4199  &  wire3754 ) ;
 assign wire18060 = ( wire4771 ) | ( wire9605  &  wire4199  &  wire3754 ) ;
 assign wire18068 = ( wire4761 ) | ( wire4759 ) ;
 assign wire18069 = ( wire4750 ) | ( wire4763 ) | ( wire4764 ) ;
 assign wire18070 = ( wire11120  &  wire4260 ) | ( wire14975  &  wire4269 ) ;
 assign wire18071 = ( wire4749 ) | ( wire4751 ) | ( wire4752 ) | ( wire4753 ) ;
 assign wire18073 = ( wire4755 ) | ( wire4756 ) | ( wire4757 ) | ( wire4758 ) ;
 assign wire18078 = ( wire4766 ) | ( wire18068 ) | ( wire18069 ) | ( wire18070 ) ;
 assign wire18079 = ( wire4744 ) | ( wire5555  &  wire5513 ) | ( wire5555  &  wire5514 ) ;
 assign wire18080 = ( wire18079 ) | ( wire6290  &  wire4199  &  wire3740 ) ;
 assign wire18114 = ( wire4626 ) | ( wire14810  &  wire4269 ) ;
 assign wire18115 = ( wire4615 ) | ( wire4624 ) | ( wire5090  &  wire4260 ) ;
 assign wire18117 = ( wire4616 ) | ( wire4617 ) | ( wire4618 ) | ( wire4620 ) ;
 assign wire18120 = ( wire4621 ) | ( wire4622 ) | ( wire4628 ) | ( wire18117 ) ;
 assign wire18124 = ( wire4611 ) | ( wire4608 ) ;
 assign wire18125 = ( ppeakp_8_8_  &  wire4298 ) | ( ppeaka_9_9_  &  wire4392 ) ;
 assign wire18127 = ( (~ ppeaka_8_8_)  &  wire4260 ) | ( wire15695  &  wire4269 ) ;
 assign wire18128 = ( wire4599 ) | ( (~ ppeakb_8_8_)  &  wire4260 ) | ( ppeakb_8_8_  &  wire4397 ) ;
 assign wire18130 = ( wire4601 ) | ( wire4602 ) | ( wire4606 ) | ( wire4607 ) ;
 assign wire18134 = ( wire4614 ) | ( wire18124 ) | ( wire18125 ) | ( wire18127 ) ;
 assign wire18135 = ( wire4598 ) | ( wire8945  &  wire4199  &  wire3754 ) ;
 assign wire18144 = ( wire4587 ) | ( wire4586 ) ;
 assign wire18145 = ( wire4577 ) | ( wire4590 ) | ( wire4591 ) ;
 assign wire18146 = ( wire11375  &  wire4260 ) | ( wire6725  &  wire4269 ) ;
 assign wire18147 = ( wire4576 ) | ( wire4578 ) | ( wire4579 ) | ( wire4581 ) ;
 assign wire18148 = ( wire4582 ) | ( wire4583 ) | ( wire4584 ) | ( wire4585 ) ;
 assign wire18153 = ( wire4593 ) | ( wire18144 ) | ( wire18145 ) | ( wire18146 ) ;
 assign wire18160 = ( wire4569 ) | ( wire4568 ) ;
 assign wire18161 = ( wire4558 ) | ( wire4571 ) | ( wire4572 ) ;
 assign wire18162 = ( wire9275  &  wire4260 ) | ( wire13745  &  wire4269 ) ;
 assign wire18163 = ( wire4557 ) | ( wire4560 ) | ( wire4561 ) | ( wire4562 ) ;
 assign wire18164 = ( wire4563 ) | ( wire4564 ) | ( wire4566 ) | ( wire4567 ) ;
 assign wire18170 = ( wire4575 ) | ( wire18160 ) | ( wire18161 ) | ( wire18162 ) ;
 assign wire18171 = ( wire4553 ) | ( wire8855  &  wire5513 ) | ( wire8855  &  wire5514 ) ;
 assign wire18172 = ( wire18171 ) | ( wire11210  &  wire4199  &  wire3740 ) ;
 assign wire18189 = ( wire4184 ) | ( wire15890  &  wire4269 ) ;
 assign wire18190 = ( wire4175 ) | ( wire4183 ) | ( wire4370  &  wire4260 ) ;
 assign wire18192 = ( wire4176 ) | ( wire4177 ) | ( wire4178 ) | ( wire4179 ) ;
 assign wire18196 = ( wire4180 ) | ( wire4181 ) | ( wire4186 ) | ( wire18192 ) ;
 assign wire18201 = ( wire4172 ) | ( wire7130  &  wire4269 ) ;
 assign wire18202 = ( wire4163 ) | ( wire4171 ) | ( wire5780  &  wire4260 ) ;
 assign wire18203 = ( wire4164 ) | ( wire4165 ) | ( wire4166 ) | ( wire4167 ) ;
 assign wire18208 = ( wire4168 ) | ( wire4169 ) | ( wire4174 ) | ( wire18203 ) ;
 assign wire18209 = ( wire4162 ) | ( wire5630  &  wire4199  &  wire3754 ) ;
 assign wire18217 = ( wire4153 ) | ( wire4152 ) ;
 assign wire18218 = ( wire4144 ) | ( wire4155 ) | ( wire4156 ) ;
 assign wire18219 = ( wire15320  &  wire4260 ) | ( wire7355  &  wire4269 ) ;
 assign wire18221 = ( wire4143 ) | ( wire4145 ) | ( wire4146 ) | ( wire4147 ) ;
 assign wire18222 = ( wire4148 ) | ( wire4149 ) | ( wire4150 ) | ( wire4151 ) ;
 assign wire18226 = ( wire4158 ) | ( wire18217 ) | ( wire18218 ) | ( wire18219 ) ;
 assign wire18234 = ( wire4137 ) | ( wire4136 ) ;
 assign wire18235 = ( wire4128 ) | ( wire4139 ) | ( wire4140 ) ;
 assign wire18236 = ( wire8615  &  wire4260 ) | ( wire14135  &  wire4269 ) ;
 assign wire18237 = ( wire4127 ) | ( wire4129 ) | ( wire4130 ) | ( wire4131 ) ;
 assign wire18238 = ( wire4132 ) | ( wire4133 ) | ( wire4134 ) | ( wire4135 ) ;
 assign wire18242 = ( wire4142 ) | ( wire18234 ) | ( wire18235 ) | ( wire18236 ) ;
 assign wire18244 = ( wire4123 ) | ( wire9530  &  wire5513 ) | ( wire9530  &  wire5514 ) ;
 assign wire18245 = ( wire18244 ) | ( wire10955  &  wire4199  &  wire3740 ) ;
 assign wire18253 = ( wire4043 ) | ( wire11240  &  wire4199  &  wire3754 ) ;
 assign wire18261 = ( wire4034 ) | ( wire4033 ) ;
 assign wire18262 = ( wire4025 ) | ( wire4036 ) | ( wire4037 ) ;
 assign wire18263 = ( wire4640  &  wire4260 ) | ( wire5360  &  wire4269 ) ;
 assign wire18264 = ( wire4023 ) | ( wire4026 ) | ( wire4027 ) | ( wire4028 ) ;
 assign wire18265 = ( wire4029 ) | ( wire4030 ) | ( wire4031 ) | ( wire4032 ) ;
 assign wire18270 = ( wire4039 ) | ( wire18261 ) | ( wire18262 ) | ( wire18263 ) ;
 assign wire18276 = ( wire4017 ) | ( wire4016 ) ;
 assign wire18277 = ( wire4008 ) | ( wire4019 ) | ( wire4020 ) ;
 assign wire18278 = ( wire4625  &  wire4260 ) | ( wire16055  &  wire4269 ) ;
 assign wire18279 = ( wire4007 ) | ( wire4009 ) | ( wire4010 ) | ( wire4011 ) ;
 assign wire18280 = ( wire4012 ) | ( wire4013 ) | ( wire4014 ) | ( wire4015 ) ;
 assign wire18286 = ( wire4022 ) | ( wire18276 ) | ( wire18277 ) | ( wire18278 ) ;
 assign wire18287 = ( wire4003 ) | ( wire7565  &  wire5513 ) | ( wire7565  &  wire5514 ) ;
 assign wire18288 = ( wire18287 ) | ( wire11195  &  wire4199  &  wire3740 ) ;
 assign wire18291 = ( wire3926 ) | ( wire10430  &  wire4199  &  wire3754 ) ;
 assign wire18300 = ( wire3917 ) | ( wire3916 ) ;
 assign wire18301 = ( wire3908 ) | ( wire3919 ) | ( wire3920 ) ;
 assign wire18302 = ( wire5345  &  wire4260 ) | ( wire6050  &  wire4269 ) ;
 assign wire18303 = ( wire3907 ) | ( wire3909 ) | ( wire3910 ) | ( wire3911 ) ;
 assign wire18304 = ( wire3912 ) | ( wire3913 ) | ( wire3914 ) | ( wire3915 ) ;
 assign wire18309 = ( wire3922 ) | ( wire18300 ) | ( wire18301 ) | ( wire18302 ) ;
 assign wire18310 = ( wire3903 ) | ( wire9815  &  wire5513 ) | ( wire9815  &  wire5514 ) ;
 assign wire18312 = ( wire18310 ) | ( wire8900  &  wire4199  &  wire3740 ) ;
 assign wire18315 = ( wire3897 ) | ( wire8195  &  wire5513 ) | ( wire8195  &  wire5514 ) ;
 assign wire18316 = ( wire18315 ) | ( wire10940  &  wire4199  &  wire3740 ) ;
 assign wire18320 = ( wire3820 ) | ( wire10715  &  wire4199  &  wire3754 ) ;
 assign wire18327 = ( wire3811 ) | ( wire3810 ) ;
 assign wire18328 = ( wire3802 ) | ( wire3813 ) | ( wire3814 ) ;
 assign wire18329 = ( wire6020  &  wire4260 ) | ( wire15350  &  wire4269 ) ;
 assign wire18330 = ( wire3801 ) | ( wire3803 ) | ( wire3804 ) | ( wire3805 ) ;
 assign wire18331 = ( wire3806 ) | ( wire3807 ) | ( wire3808 ) | ( wire3809 ) ;
 assign wire18336 = ( wire3816 ) | ( wire18327 ) | ( wire18328 ) | ( wire18329 ) ;
 assign wire18338 = ( wire3797 ) | ( wire10655  &  wire5513 ) | ( wire10655  &  wire5514 ) ;
 assign wire18339 = ( wire18338 ) | ( wire5600  &  wire4199  &  wire3740 ) ;
 assign wire18342 = ( wire3791 ) | ( wire6260  &  wire5513 ) | ( wire6260  &  wire5514 ) ;
 assign wire18343 = ( wire18342 ) | ( wire6950  &  wire4199  &  wire3740 ) ;
 assign wire18353 = ( wire3689 ) | ( wire3688 ) ;
 assign wire18354 = ( wire3680 ) | ( wire3691 ) | ( wire3692 ) ;
 assign wire18355 = ( wire6710  &  wire4260 ) | ( wire4655  &  wire4269 ) ;
 assign wire18356 = ( wire3679 ) | ( wire3681 ) | ( wire3682 ) | ( wire3683 ) ;
 assign wire18357 = ( wire3684 ) | ( wire3685 ) | ( wire3686 ) | ( wire3687 ) ;
 assign wire18362 = ( wire3694 ) | ( wire18353 ) | ( wire18354 ) | ( wire18355 ) ;
 assign wire18369 = ( wire3673 ) | ( wire3672 ) ;
 assign wire18370 = ( wire3664 ) | ( wire3675 ) | ( wire3676 ) ;
 assign wire18372 = ( wire6695  &  wire4260 ) | ( wire15710  &  wire4269 ) ;
 assign wire18373 = ( wire3663 ) | ( wire3665 ) | ( wire3666 ) | ( wire3667 ) ;
 assign wire18374 = ( wire3668 ) | ( wire3669 ) | ( wire3670 ) | ( wire3671 ) ;
 assign wire18379 = ( wire3678 ) | ( wire18369 ) | ( wire18370 ) | ( wire18372 ) ;
 assign wire18380 = ( wire3659 ) | ( wire10370  &  wire5513 ) | ( wire10370  &  wire5514 ) ;
 assign wire18381 = ( wire18380 ) | ( wire4895  &  wire4199  &  wire3740 ) ;
 assign wire18385 = ( wire3653 ) | ( wire6935  &  wire5513 ) | ( wire6935  &  wire5514 ) ;
 assign wire18386 = ( wire18385 ) | ( wire6275  &  wire4199  &  wire3740 ) ;
 assign wire18401 = ( wire3290 ) | ( wire13250  &  wire4269 ) ;
 assign wire18402 = ( wire3281 ) | ( wire3289 ) | ( wire13235  &  wire4260 ) ;
 assign wire18403 = ( wire3282 ) | ( wire3283 ) | ( wire3284 ) | ( wire3285 ) ;
 assign wire18406 = ( wire3286 ) | ( wire3287 ) | ( wire3292 ) | ( wire18403 ) ;
 assign wire18408 = ( wire3269 ) | ( wire7880  &  wire4199  &  wire3747 ) ;
 assign wire18414 = ( wire18408 ) | ( wire3266 ) ;
 assign wire18416 = ( wire3259 ) | ( wire3260 ) | ( wire3261 ) | ( wire3262 ) ;
 assign wire18417 = ( wire3263 ) | ( wire3264 ) | ( wire3265 ) | ( wire3267 ) ;
 assign wire18421 = ( wire3228 ) | ( wire6620  &  wire4199  &  wire3747 ) ;
 assign wire18427 = ( wire18421 ) | ( wire3225 ) ;
 assign wire18429 = ( wire3218 ) | ( wire3219 ) | ( wire3220 ) | ( wire3221 ) ;
 assign wire18430 = ( wire3222 ) | ( wire3223 ) | ( wire3224 ) | ( wire3226 ) ;
 assign wire18445 = ( wire3090 ) | ( wire5795  &  wire4269 ) ;
 assign wire18446 = ( wire3081 ) | ( wire3089 ) | ( wire14360  &  wire4260 ) ;
 assign wire18447 = ( wire3082 ) | ( wire3083 ) | ( wire3084 ) | ( wire3085 ) ;
 assign wire18451 = ( wire3086 ) | ( wire3087 ) | ( wire3092 ) | ( wire18447 ) ;
 assign wire18455 = ( wire3077 ) | ( wire3075 ) ;
 assign wire18456 = ( ppeakp_9_9_  &  wire4298 ) | ( ppeaka_10_10_  &  wire4392 ) ;
 assign wire18457 = ( (~ ppeaka_9_9_)  &  wire4260 ) | ( wire16040  &  wire4269 ) ;
 assign wire18458 = ( wire3067 ) | ( (~ ppeakb_9_9_)  &  wire4260 ) | ( ppeakb_9_9_  &  wire4397 ) ;
 assign wire18459 = ( wire3069 ) | ( wire3070 ) | ( wire3073 ) | ( wire3074 ) ;
 assign wire18463 = ( wire3080 ) | ( wire18455 ) | ( wire18456 ) | ( wire18457 ) ;
 assign wire18470 = ( wire3024 ) | ( wire6485  &  wire4269 ) ;
 assign wire18471 = ( wire3015 ) | ( wire3023 ) | ( wire13955  &  wire4260 ) ;
 assign wire18472 = ( wire3016 ) | ( wire3017 ) | ( wire3018 ) | ( wire3019 ) ;
 assign wire18476 = ( wire3020 ) | ( wire3021 ) | ( wire3026 ) | ( wire18472 ) ;
 assign wire18477 = ( wire3014 ) | ( wire9890  &  wire4199  &  wire3754 ) ;
 assign wire18479 = ( wire3007 ) | ( wire10085  &  wire5513 ) | ( wire10085  &  wire5514 ) ;
 assign wire18481 = ( wire18479 ) | ( wire9575  &  wire4199  &  wire3740 ) ;
 assign wire18487 = ( wire2959 ) | ( wire2957 ) ;
 assign wire18489 = ( ppeakp_11_11_  &  wire4298 ) | ( ppeaka_12_12_  &  wire4392 ) ;
 assign wire18490 = ( (~ ppeakb_11_11_)  &  wire4260 ) | ( wire15335  &  wire4269 ) ;
 assign wire18491 = ( wire2949 ) | ( wire2950 ) | ( (~ ppeaka_11_11_)  &  wire4260 ) ;
 assign wire18492 = ( wire2951 ) | ( wire2952 ) | ( wire2955 ) | ( wire2956 ) ;
 assign wire18497 = ( wire2962 ) | ( wire18487 ) | ( wire18489 ) | ( wire18490 ) ;
 assign wire18505 = ( wire2934 ) | ( wire2935 ) | ( wire2944 ) ;
 assign wire18507 = ( wire2936 ) | ( wire2937 ) | ( wire2938 ) | ( wire2939 ) ;
 assign wire18508 = ( wire2933 ) | ( wire2940 ) | ( wire2941 ) | ( wire2945 ) ;
 assign wire18511 = ( wire2942 ) | ( wire2943 ) | ( wire18505 ) | ( wire18508 ) ;
 assign wire18512 = ( wire2929 ) | ( wire8840  &  wire5513 ) | ( wire8840  &  wire5514 ) ;
 assign wire18513 = ( wire18512 ) | ( wire11660  &  wire4199  &  wire3740 ) ;
 assign wire18517 = ( wire2882 ) | ( wire14915  &  wire4199  &  wire3747 ) ;
 assign wire18522 = ( wire18517 ) | ( wire2879 ) ;
 assign wire18523 = ( wire2872 ) | ( wire2873 ) | ( wire2874 ) | ( wire2875 ) ;
 assign wire18524 = ( wire2876 ) | ( wire2877 ) | ( wire2878 ) | ( wire2880 ) ;
 assign wire18534 = ( wire2858 ) | ( wire2859 ) | ( wire2868 ) ;
 assign wire18535 = ( wire2860 ) | ( wire2861 ) | ( wire2862 ) | ( wire2863 ) ;
 assign wire18536 = ( wire2857 ) | ( wire2864 ) | ( wire2865 ) | ( wire2869 ) ;
 assign wire18539 = ( wire2866 ) | ( wire2867 ) | ( wire18534 ) | ( wire18536 ) ;
 assign wire18548 = ( wire2844 ) | ( wire2845 ) | ( wire2854 ) ;
 assign wire18549 = ( wire2846 ) | ( wire2847 ) | ( wire2848 ) | ( wire2849 ) ;
 assign wire18550 = ( wire2843 ) | ( wire2850 ) | ( wire2851 ) | ( wire2855 ) ;
 assign wire18553 = ( wire2852 ) | ( wire2853 ) | ( wire18548 ) | ( wire18550 ) ;
 assign wire18554 = ( wire2839 ) | ( wire9515  &  wire5513 ) | ( wire9515  &  wire5514 ) ;
 assign wire18556 = ( wire18554 ) | ( wire11435  &  wire4199  &  wire3740 ) ;
 assign wire18559 = ( wire2790 ) | ( wire13010  &  wire4199  &  wire3747 ) ;
 assign wire18564 = ( wire18559 ) | ( wire2787 ) ;
 assign wire18565 = ( wire2780 ) | ( wire2781 ) | ( wire2782 ) | ( wire2783 ) ;
 assign wire18566 = ( wire2784 ) | ( wire2785 ) | ( wire2786 ) | ( wire2788 ) ;
 assign wire18574 = ( wire2775 ) | ( wire2773 ) ;
 assign wire18575 = ( ppeakp_13_13_  &  wire4298 ) | ( ppeaka_14_14_  &  wire4392 ) ;
 assign wire18576 = ( (~ ppeakb_13_13_)  &  wire4260 ) | ( wire14540  &  wire4269 ) ;
 assign wire18577 = ( wire2765 ) | ( wire2766 ) | ( (~ ppeaka_13_13_)  &  wire4260 ) ;
 assign wire18578 = ( wire2767 ) | ( wire2768 ) | ( wire2771 ) | ( wire2772 ) ;
 assign wire18583 = ( wire2778 ) | ( wire18574 ) | ( wire18575 ) | ( wire18576 ) ;
 assign wire18591 = ( wire2752 ) | ( wire2753 ) | ( wire2762 ) ;
 assign wire18592 = ( wire2754 ) | ( wire2755 ) | ( wire2756 ) | ( wire2757 ) ;
 assign wire18593 = ( wire2751 ) | ( wire2758 ) | ( wire2759 ) | ( wire2763 ) ;
 assign wire18598 = ( wire2760 ) | ( wire2761 ) | ( wire18591 ) | ( wire18593 ) ;
 assign wire18599 = ( wire2750 ) | ( wire9875  &  wire4199  &  wire3754 ) ;
 assign wire18607 = ( wire2741 ) | ( wire2740 ) ;
 assign wire18608 = ( wire2732 ) | ( wire2743 ) | ( wire2744 ) ;
 assign wire18609 = ( wire7970  &  wire4260 ) | ( wire13040  &  wire4269 ) ;
 assign wire18611 = ( wire2731 ) | ( wire2733 ) | ( wire2734 ) | ( wire2735 ) ;
 assign wire18612 = ( wire2736 ) | ( wire2737 ) | ( wire2738 ) | ( wire2739 ) ;
 assign wire18616 = ( wire2746 ) | ( wire18607 ) | ( wire18608 ) | ( wire18609 ) ;
 assign wire18617 = ( wire2727 ) | ( wire7580  &  wire5513 ) | ( wire7580  &  wire5514 ) ;
 assign wire18619 = ( wire18617 ) | ( wire11675  &  wire4199  &  wire3740 ) ;
 assign wire18622 = ( wire2688 ) | ( wire16010  &  wire4199  &  wire3747 ) ;
 assign wire18627 = ( wire18622 ) | ( wire2685 ) ;
 assign wire18628 = ( wire2678 ) | ( wire2679 ) | ( wire2680 ) | ( wire2681 ) ;
 assign wire18629 = ( wire2682 ) | ( wire2683 ) | ( wire2684 ) | ( wire2686 ) ;
 assign wire18637 = ( wire2673 ) | ( wire2671 ) ;
 assign wire18638 = ( ppeakp_12_12_  &  wire4298 ) | ( ppeaka_13_13_  &  wire4392 ) ;
 assign wire18639 = ( (~ ppeaka_12_12_)  &  wire4260 ) | ( wire14120  &  wire4269 ) ;
 assign wire18640 = ( wire2663 ) | ( (~ ppeakb_12_12_)  &  wire4260 ) | ( ppeakb_12_12_  &  wire4397 ) ;
 assign wire18641 = ( wire2665 ) | ( wire2666 ) | ( wire2669 ) | ( wire2670 ) ;
 assign wire18646 = ( wire2676 ) | ( wire18637 ) | ( wire18638 ) | ( wire18639 ) ;
 assign wire18653 = ( wire2650 ) | ( wire2651 ) | ( wire2660 ) ;
 assign wire18654 = ( wire2652 ) | ( wire2653 ) | ( wire2654 ) | ( wire2655 ) ;
 assign wire18655 = ( wire2649 ) | ( wire2656 ) | ( wire2657 ) | ( wire2661 ) ;
 assign wire18658 = ( wire2658 ) | ( wire2659 ) | ( wire18653 ) | ( wire18655 ) ;
 assign wire18659 = ( wire2648 ) | ( wire10730  &  wire4199  &  wire3754 ) ;
 assign wire18666 = ( wire2639 ) | ( wire2638 ) ;
 assign wire18667 = ( wire2630 ) | ( wire2641 ) | ( wire2642 ) ;
 assign wire18668 = ( wire7340  &  wire4260 ) | ( wire13385  &  wire4269 ) ;
 assign wire18669 = ( wire2629 ) | ( wire2631 ) | ( wire2632 ) | ( wire2633 ) ;
 assign wire18670 = ( wire2634 ) | ( wire2635 ) | ( wire2636 ) | ( wire2637 ) ;
 assign wire18674 = ( wire2644 ) | ( wire18666 ) | ( wire18667 ) | ( wire18668 ) ;
 assign wire18675 = ( wire2625 ) | ( wire8210  &  wire5513 ) | ( wire8210  &  wire5514 ) ;
 assign wire18676 = ( wire18675 ) | ( wire11450  &  wire4199  &  wire3740 ) ;
 assign wire18679 = ( wire2586 ) | ( wire13685  &  wire4199  &  wire3747 ) ;
 assign wire18684 = ( wire18679 ) | ( wire2583 ) ;
 assign wire18685 = ( wire2576 ) | ( wire2577 ) | ( wire2578 ) | ( wire2579 ) ;
 assign wire18686 = ( wire2580 ) | ( wire2581 ) | ( wire2582 ) | ( wire2584 ) ;
 assign wire18695 = ( wire2562 ) | ( wire2563 ) | ( wire2564 ) | ( wire2565 ) ;
 assign wire18696 = ( wire2566 ) | ( wire2567 ) | ( wire2569 ) | ( wire2573 ) ;
 assign wire18697 = ( wire2568 ) | ( wire2570 ) | ( wire2571 ) | ( wire2572 ) ;
 assign wire18706 = ( wire2549 ) | ( wire2550 ) | ( wire2559 ) ;
 assign wire18707 = ( wire2551 ) | ( wire2552 ) | ( wire2553 ) | ( wire2554 ) ;
 assign wire18708 = ( wire2548 ) | ( wire2555 ) | ( wire2556 ) | ( wire2560 ) ;
 assign wire18711 = ( wire2557 ) | ( wire2558 ) | ( wire18706 ) | ( wire18708 ) ;
 assign wire18712 = ( wire2547 ) | ( wire10445  &  wire4199  &  wire3754 ) ;
 assign wire18714 = ( wire2543 ) | ( wire8930  &  wire4199  &  wire3754 ) ;
 assign wire18721 = ( wire2534 ) | ( wire2533 ) ;
 assign wire18722 = ( wire2525 ) | ( wire2536 ) | ( wire2537 ) ;
 assign wire18723 = ( wire5330  &  wire4260 ) | ( wire13025  &  wire4269 ) ;
 assign wire18724 = ( wire2524 ) | ( wire2526 ) | ( wire2527 ) | ( wire2528 ) ;
 assign wire18725 = ( wire2529 ) | ( wire2530 ) | ( wire2531 ) | ( wire2532 ) ;
 assign wire18729 = ( wire2539 ) | ( wire18721 ) | ( wire18722 ) | ( wire18723 ) ;
 assign wire18734 = ( wire2489 ) | ( wire6500  &  wire4269 ) ;
 assign wire18735 = ( wire2480 ) | ( wire2488 ) | ( wire7115  &  wire4260 ) ;
 assign wire18736 = ( wire2481 ) | ( wire2482 ) | ( wire2483 ) | ( wire2484 ) ;
 assign wire18739 = ( wire2485 ) | ( wire2486 ) | ( wire2491 ) | ( wire18736 ) ;
 assign wire18743 = ( wire2476 ) | ( wire2474 ) ;
 assign wire18744 = ( ppeakp_14_14_  &  wire4298 ) | ( ppeaka_15_15_  &  wire4392 ) ;
 assign wire18745 = ( (~ ppeaka_14_14_)  &  wire4260 ) | ( wire13370  &  wire4269 ) ;
 assign wire18746 = ( wire2466 ) | ( (~ ppeakb_14_14_)  &  wire4260 ) | ( ppeakb_14_14_  &  wire4397 ) ;
 assign wire18747 = ( wire2468 ) | ( wire2469 ) | ( wire2472 ) | ( wire2473 ) ;
 assign wire18751 = ( wire2479 ) | ( wire18743 ) | ( wire18744 ) | ( wire18745 ) ;
 assign wire18758 = ( wire2453 ) | ( wire2454 ) | ( wire2463 ) ;
 assign wire18759 = ( wire2455 ) | ( wire2456 ) | ( wire2457 ) | ( wire2458 ) ;
 assign wire18760 = ( wire2452 ) | ( wire2459 ) | ( wire2460 ) | ( wire2464 ) ;
 assign wire18763 = ( wire2461 ) | ( wire2462 ) | ( wire18758 ) | ( wire18760 ) ;
 assign wire18764 = ( wire2451 ) | ( wire8285  &  wire4199  &  wire3754 ) ;
 assign wire18766 = ( wire2447 ) | ( wire10145  &  wire4199  &  wire3754 ) ;
 assign wire18773 = ( wire2438 ) | ( wire2437 ) ;
 assign wire18774 = ( wire2429 ) | ( wire2440 ) | ( wire2441 ) ;
 assign wire18775 = ( wire6035  &  wire4260 ) | ( wire12800  &  wire4269 ) ;
 assign wire18776 = ( wire2428 ) | ( wire2430 ) | ( wire2431 ) | ( wire2432 ) ;
 assign wire18777 = ( wire2433 ) | ( wire2434 ) | ( wire2435 ) | ( wire2436 ) ;
 assign wire18781 = ( wire2443 ) | ( wire18773 ) | ( wire18774 ) | ( wire18775 ) ;
 assign wire18783 = ( wire17999  &  (~ wire18220) ) | ( (~ wire17791)  &  nen2_3 ) ;
 assign wire18784 = ( (~ wire17050)  &  wire17115 ) | ( wire17180  &  (~ wire17232) ) ;
 assign wire18785 = ( wire17206  &  (~ wire17271) ) | ( wire16933  &  (~ wire17388) ) ;
 assign wire18786 = ( (~ wire17414)  &  wire17843 ) | ( wire18311  &  (~ wire18389) ) ;
 assign wire18789 = ( wire18786 ) | ( wire18785 ) ;
 assign wire18790 = ( wire4235 ) | ( nrq14_8 ) | ( wire4488 ) | ( wire18784 ) ;
 assign wire18792 = ( nrq3_5 ) | ( wire18783 ) | ( wire18789 ) | ( wire18790 ) ;
 assign wire18793 = ( wire18792 ) | ( (~ wire17167)  &  nrq7_2  &  wire3727 ) ;
 assign wire18795 = ( nrq23_3 ) | ( nrq14_3 ) | ( wire4234 ) ;
 assign wire18796 = ( nrq10_4 ) | ( wire17717 ) | ( wire17718 ) | ( wire18793 ) ;
 assign wire18797 = ( wire17396 ) | ( (~ preset)  &  wire17284  &  (~ wire18376) ) ;
 assign wire18798 = ( wire18797 ) | ( (~ preset)  &  nrq7_2  &  wire17714 ) ;
 assign wire18799 = ( (~ preset)  &  nrq7_2  &  wire17712 ) | ( (~ preset)  &  nrq7_2  &  wire17715 ) ;
 assign wire18804 = ( wire2386 ) | ( wire2383 ) ;
 assign wire18805 = ( wire2387 ) | ( ppeakb_8_8_  &  wire4382 ) ;
 assign wire18806 = ( wire13460  &  wire4369 ) | ( wire7595  &  wire4378 ) ;
 assign wire18807 = ( wire11420  &  wire4341 ) | ( wire6410  &  wire4351 ) ;
 assign wire18808 = ( wire2378 ) | ( wire2380 ) | ( wire2381 ) | ( wire2382 ) ;
 assign wire18813 = ( wire2388 ) | ( wire2389 ) | ( wire18804 ) | ( wire18805 ) ;
 assign wire18814 = ( wire2390 ) | ( wire18806 ) | ( wire18807 ) | ( wire18808 ) ;
 assign wire18815 = ( wire2375 ) | ( (~ preset)  &  ppeakb_7_7_  &  wire4242 ) ;
 assign wire18816 = ( (~ wire17388)  &  (~ preset) ) ;
 assign wire18819 = ( wire2366 ) | ( wire2363 ) ;
 assign wire18820 = ( wire2367 ) | ( ppeakb_9_9_  &  wire4382 ) ;
 assign wire18821 = ( wire13820  &  wire4369 ) | ( wire10685  &  wire4378 ) ;
 assign wire18822 = ( wire11645  &  wire4341 ) | ( wire5720  &  wire4351 ) ;
 assign wire18823 = ( wire2358 ) | ( wire2360 ) | ( wire2361 ) | ( wire2362 ) ;
 assign wire18828 = ( wire2368 ) | ( wire2369 ) | ( wire18819 ) | ( wire18820 ) ;
 assign wire18829 = ( wire2370 ) | ( wire18821 ) | ( wire18822 ) | ( wire18823 ) ;
 assign wire18830 = ( wire2355 ) | ( (~ preset)  &  ppeakb_8_8_  &  wire4242 ) ;
 assign wire18832 = ( wire2352 ) | ( (~ preset)  &  ppeakb_5_5_  &  wire4242 ) ;
 assign wire18833 = ( wire2345 ) | ( (~ preset)  &  ppeakb_6_6_  &  wire4242 ) ;
 assign wire18834 = ( wire2342 ) | ( (~ preset)  &  ppeakb_15_15_  &  wire4242 ) ;
 assign wire18835 = ( (~ wire17050)  &  (~ preset) ) ;
 assign wire18836 = ( wire2337 ) | ( (~ preset)  &  ppeakb_3_3_  &  wire4242 ) ;
 assign wire18837 = ( (~ wire17232)  &  (~ preset) ) ;
 assign wire18838 = ( wire2330 ) | ( (~ preset)  &  ppeakb_4_4_  &  wire4242 ) ;
 assign wire18839 = ( (~ wire17271)  &  (~ preset) ) ;
 assign wire18842 = ( wire2325 ) | ( (~ preset)  &  ppeakb_1_1_  &  wire4242 ) ;
 assign wire18843 = ( (~ wire18376)  &  (~ preset) ) ;
 assign wire18845 = ( wire2320 ) | ( (~ preset)  &  ppeakb_2_2_  &  wire4242 ) ;
 assign wire18851 = ( wire2311 ) | ( wire2308 ) ;
 assign wire18852 = ( wire2312 ) | ( ppeakb_11_11_  &  wire4382 ) ;
 assign wire18853 = ( wire13115  &  wire4369 ) | ( wire10115  &  wire4378 ) ;
 assign wire18854 = ( wire16100  &  wire4341 ) | ( wire4295  &  wire4351 ) ;
 assign wire18855 = ( wire2303 ) | ( wire2305 ) | ( wire2306 ) | ( wire2307 ) ;
 assign wire18860 = ( wire2313 ) | ( wire2314 ) | ( wire18851 ) | ( wire18852 ) ;
 assign wire18862 = ( wire2315 ) | ( wire18853 ) | ( wire18854 ) | ( wire18855 ) ;
 assign wire18865 = ( wire2294 ) | ( wire2291 ) ;
 assign wire18866 = ( wire2295 ) | ( ppeakb_10_10_  &  wire4382 ) ;
 assign wire18867 = ( wire12860  &  wire4369 ) | ( wire10400  &  wire4378 ) ;
 assign wire18868 = ( wire10925  &  wire4341 ) | ( wire5015  &  wire4351 ) ;
 assign wire18869 = ( wire2286 ) | ( wire2288 ) | ( wire2289 ) | ( wire2290 ) ;
 assign wire18874 = ( wire2296 ) | ( wire2297 ) | ( wire18865 ) | ( wire18866 ) ;
 assign wire18875 = ( wire2298 ) | ( wire18867 ) | ( wire18868 ) | ( wire18869 ) ;
 assign wire18876 = ( wire2281 ) | ( (~ preset)  &  ppeakb_13_13_  &  wire4242 ) ;
 assign wire18880 = ( wire2268 ) | ( wire2265 ) ;
 assign wire18881 = ( wire2269 ) | ( ppeakb_13_13_  &  wire4382 ) ;
 assign wire18882 = ( wire12620  &  wire4369 ) | ( wire8885  &  wire4378 ) ;
 assign wire18883 = ( wire13805  &  wire4341 ) | ( wire15500  &  wire4351 ) ;
 assign wire18884 = ( wire2260 ) | ( wire2262 ) | ( wire2263 ) | ( wire2264 ) ;
 assign wire18889 = ( wire2270 ) | ( wire2271 ) | ( wire18880 ) | ( wire18881 ) ;
 assign wire18890 = ( wire2272 ) | ( wire18882 ) | ( wire18883 ) | ( wire18884 ) ;
 assign wire18891 = ( (~ wire4292) ) | ( (~ ppeaki_13_13_)  &  (~ ppeaki_12_12_) ) ;
 assign wire18892 = ( (~ wire4292) ) | ( (~ ppeaki_15_15_)  &  (~ ppeaki_14_14_) ) ;
 assign wire18897 = ( (~ wire4292)  &  wire18891 ) | ( (~ ppeaki_15_15_)  &  (~ ppeaki_14_14_)  &  wire18891 ) ;
 assign wire18898 = ( (~ wire1427)  &  (~ wire1342)  &  (~ wire1353)  &  (~ wire1439) ) ;
 assign wire18899 = ( (~ wire1368)  &  (~ wire1386)  &  (~ wire1398)  &  (~ wire1413) ) ;
 assign wire18900 = ( wire18891  &  wire18892  &  wire18898 ) ;
 assign wire18901 = ( wire18636  &  wire18899 ) | ( (~ nrq7_2)  &  wire17582  &  wire18899 ) ;
 assign wire18902 = ( wire17986  &  wire17596 ) ;
 assign wire18904 = ( wire17804 ) | ( wire2255 ) | ( wire17986  &  wire18597 ) ;
 assign wire18905 = ( (~ preset)  &  wire17596  &  (~ wire18597) ) ;
 assign wire18906 = ( (~ preset)  &  (~ wire17596)  &  wire4513 ) ;
 assign wire18909 = ( wire2239 ) | ( wire2236 ) ;
 assign wire18910 = ( wire2240 ) | ( ppeakb_12_12_  &  wire4382 ) ;
 assign wire18911 = ( wire12395  &  wire4369 ) | ( wire9845  &  wire4378 ) ;
 assign wire18912 = ( wire15755  &  wire4341 ) | ( wire15845  &  wire4351 ) ;
 assign wire18914 = ( wire2231 ) | ( wire2233 ) | ( wire2234 ) | ( wire2235 ) ;
 assign wire18919 = ( wire2241 ) | ( wire2242 ) | ( wire18909 ) | ( wire18910 ) ;
 assign wire18920 = ( wire2243 ) | ( wire18911 ) | ( wire18912 ) | ( wire18914 ) ;
 assign wire18923 = ( wire2218 ) | ( wire2215 ) ;
 assign wire18924 = ( wire2219 ) | ( ppeakb_15_15_  &  wire4382 ) ;
 assign wire18925 = ( wire15050  &  wire4369 ) | ( wire4880  &  wire4378 ) ;
 assign wire18926 = ( wire14615  &  wire4341 ) | ( wire13550  &  wire4351 ) ;
 assign wire18927 = ( wire2210 ) | ( wire2212 ) | ( wire2213 ) | ( wire2214 ) ;
 assign wire18932 = ( wire2220 ) | ( wire2221 ) | ( wire18923 ) | ( wire18924 ) ;
 assign wire18933 = ( wire2222 ) | ( wire18925 ) | ( wire18926 ) | ( wire18927 ) ;
 assign wire18936 = ( wire2201 ) | ( wire2198 ) ;
 assign wire18937 = ( wire2202 ) | ( ppeakb_14_14_  &  wire4382 ) ;
 assign wire18938 = ( wire15410  &  wire4369 ) | ( wire9560  &  wire4378 ) ;
 assign wire18939 = ( wire13445  &  wire4341 ) | ( wire15140  &  wire4351 ) ;
 assign wire18940 = ( wire2193 ) | ( wire2195 ) | ( wire2196 ) | ( wire2197 ) ;
 assign wire18945 = ( wire2203 ) | ( wire2204 ) | ( wire18936 ) | ( wire18937 ) ;
 assign wire18946 = ( wire2205 ) | ( wire18938 ) | ( wire18939 ) | ( wire18940 ) ;
 assign wire18947 = ( wire2188 ) | ( (~ preset)  &  ppeakb_9_9_  &  wire4242 ) ;
 assign wire18948 = ( wire2185 ) | ( (~ preset)  &  ppeakb_14_14_  &  wire4242 ) ;
 assign wire18951 = ( (~ wire17050)  &  wire17115 ) | ( wire17180  &  (~ wire17232) ) ;
 assign wire18952 = ( wire17206  &  (~ wire17271) ) | ( wire17232  &  (~ wire18441) ) ;
 assign wire18953 = ( (~ wire17427)  &  wire17518 ) | ( wire17583  &  (~ wire18077) ) ;
 assign wire18954 = ( wire17050  &  (~ wire17219) ) | ( wire17271  &  (~ wire17349) ) ;
 assign wire18958 = ( wire4235 ) | ( wire4488 ) | ( wire18951 ) | ( wire18952 ) ;
 assign wire18959 = ( wire18953 ) | ( wire18954 ) | ( wire18958 ) ;
 assign wire18960 = ( wire4235  &  (~ preset) ) ;
 assign wire18961 = ( pwr_0_0_  &  (~ preset) ) ;
 assign wire18962 = ( wire4234  &  wire18960 ) | ( wire18959  &  wire18960 ) | ( (~ wire4234)  &  (~ wire18959)  &  wire18961 ) ;
 assign wire18963 = ( (~ preset)  &  wire4234 ) | ( (~ preset)  &  nrq13_4  &  wire18959 ) ;
 assign wire18964 = ( wire17058  &  wire4234 ) | ( wire17240  &  wire4234 ) | ( wire17058  &  wire18959 ) | ( wire17240  &  wire18959 ) ;
 assign wire18966 = ( wire16933  &  (~ wire17388) ) | ( (~ wire17414)  &  wire17843 ) ;
 assign wire18967 = ( wire18311  &  (~ wire18389) ) | ( wire18363  &  (~ wire18415) ) ;
 assign wire18968 = ( wire17791  &  (~ wire17843) ) | ( wire17453  &  (~ wire18246) ) ;
 assign wire18969 = ( wire17102  &  (~ wire17154) ) | ( wire17167  &  (~ wire17362) ) ;
 assign wire18970 = ( (~ wire17310)  &  wire17388 ) | ( wire17414  &  (~ wire17505) ) ;
 assign wire18971 = ( (~ wire18142)  &  wire18220 ) | ( (~ wire18311)  &  wire18506 ) ;
 assign wire18972 = ( wire17570  &  (~ wire17635) ) | ( wire18285  &  (~ wire18363) ) ;
 assign wire18973 = ( wire18415  &  (~ wire18480) ) | ( (~ wire18428)  &  wire18493 ) ;
 assign wire18974 = ( (~ wire18298)  &  wire18376 ) | ( (~ wire16985)  &  wire18389 ) ;
 assign wire18975 = ( wire16920  &  (~ wire16972) ) | ( wire17297  &  (~ wire17375) ) ;
 assign wire18981 = ( wire4488 ) | ( wire18966 ) | ( wire18975 ) ;
 assign wire18982 = ( wire18967 ) | ( wire18968 ) | ( wire18969 ) | ( wire18970 ) ;
 assign wire18983 = ( wire18971 ) | ( wire18972 ) | ( wire18973 ) | ( wire18974 ) ;
 assign wire18985 = ( wire18981 ) | ( wire18982 ) | ( wire18983 ) ;
 assign wire18986 = ( nrq3_5 ) | ( wire18783 ) | ( wire18985 ) ;
 assign wire18987 = ( wire18986 ) | ( (~ wire17167)  &  nrq7_2  &  wire3727 ) ;
 assign wire18989 = ( nrq10_4 ) | ( nrq23_3 ) | ( nrq14_3 ) | ( wire18987 ) ;
 assign wire18990 = ( (~ preset)  &  nrq3_5 ) | ( (~ preset)  &  wire18783 ) ;
 assign wire18991 = ( prd_0_0_  &  (~ preset) ) ;
 assign wire18992 = ( wire4265  &  wire18990 ) | ( wire18989  &  wire18990 ) | ( (~ wire4265)  &  (~ wire18989)  &  wire18991 ) ;
 assign wire18993 = ( wire4243  &  wire4265 ) | ( wire4245  &  wire4265 ) | ( wire4243  &  wire18989 ) | ( wire4245  &  wire18989 ) ;
 assign wire18994 = ( wire18423  &  wire4265 ) | ( wire4241  &  wire4265 ) | ( wire18423  &  wire18989 ) | ( wire4241  &  wire18989 ) ;
 assign wire18995 = ( wire17422  &  wire4265 ) | ( wire18397  &  wire4265 ) | ( wire17422  &  wire18989 ) | ( wire18397  &  wire18989 ) ;
 assign wire18996 = ( wire17110  &  wire4265 ) | ( wire17175  &  wire4265 ) | ( wire17110  &  wire18989 ) | ( wire17175  &  wire18989 ) ;
 assign wire18999 = ( wire18992 ) | ( wire18993 ) | ( wire18996 ) ;
 assign wire19000 = ( wire2117 ) | ( (~ preset)  &  ppeakb_10_10_  &  wire4242 ) ;
 assign wire19001 = ( wire2108 ) | ( (~ preset)  &  ppeakb_12_12_  &  wire4242 ) ;
 assign wire19003 = ( wire18129  &  (~ preset) ) ;
 assign wire19004 = ( wire2077 ) | ( (~ preset)  &  ppeakb_11_11_  &  wire4242 ) ;
 assign wire19009 = ( wire2064 ) | ( wire2063 ) ;
 assign wire19010 = ( wire10670  &  wire4378 ) | ( ppeakb_0_0_  &  wire4382 ) ;
 assign wire19011 = ( wire4310  &  wire4351 ) | ( wire12605  &  wire4369 ) ;
 assign wire19012 = ( wire2055 ) | ( wire2068 ) | ( wire11630  &  wire4341 ) ;
 assign wire19013 = ( wire2057 ) | ( wire2058 ) | ( wire2059 ) | ( wire2060 ) ;
 assign wire19018 = ( wire2065 ) | ( wire2066 ) | ( wire19009 ) | ( wire19010 ) ;
 assign wire19019 = ( wire2067 ) | ( wire19011 ) | ( wire19012 ) | ( wire19013 ) ;
 assign wire19022 = ( (~ wire18415)  &  (~ preset) ) ;
 assign wire19028 = ( wire2045 ) | ( wire2041 ) ;
 assign wire19029 = ( wire9830  &  wire4378 ) | ( ppeakb_1_1_  &  wire4382 ) ;
 assign wire19030 = ( wire5030  &  wire4351 ) | ( wire12380  &  wire4369 ) ;
 assign wire19031 = ( wire2032 ) | ( wire2034 ) | ( wire9485  &  wire4341 ) ;
 assign wire19032 = ( wire2035 ) | ( wire2036 ) | ( wire2037 ) | ( wire2040 ) ;
 assign wire19037 = ( wire2042 ) | ( wire2043 ) | ( wire19028 ) | ( wire19029 ) ;
 assign wire19038 = ( wire2044 ) | ( wire19030 ) | ( wire19031 ) | ( wire19032 ) ;
 assign wire19039 = ( wire2029 ) | ( (~ preset)  &  ppeakb_0_0_  &  wire4242 ) ;
 assign wire19042 = ( wire2018 ) | ( wire2015 ) ;
 assign wire19043 = ( wire2019 ) | ( ppeakb_2_2_  &  wire4382 ) ;
 assign wire19044 = ( wire13100  &  wire4369 ) | ( wire10100  &  wire4378 ) ;
 assign wire19045 = ( wire7535  &  wire4341 ) | ( wire15515  &  wire4351 ) ;
 assign wire19046 = ( wire2010 ) | ( wire2012 ) | ( wire2013 ) | ( wire2014 ) ;
 assign wire19051 = ( wire2020 ) | ( wire2021 ) | ( wire19042 ) | ( wire19043 ) ;
 assign wire19052 = ( wire2022 ) | ( wire19044 ) | ( wire19045 ) | ( wire19046 ) ;
 assign wire19057 = ( wire2003 ) | ( wire2000 ) ;
 assign wire19058 = ( wire2004 ) | ( ppeakb_3_3_  &  wire4382 ) ;
 assign wire19059 = ( wire12845  &  wire4369 ) | ( wire5570  &  wire4378 ) ;
 assign wire19062 = ( wire8165  &  wire4341 ) | ( wire15860  &  wire4351 ) ;
 assign wire19063 = ( wire1995 ) | ( wire1997 ) | ( wire1998 ) | ( wire1999 ) ;
 assign wire19074 = ( wire2005 ) | ( wire2006 ) | ( wire19057 ) | ( wire19058 ) ;
 assign wire19075 = ( wire2007 ) | ( wire19059 ) | ( wire19062 ) | ( wire19063 ) ;
 assign wire19076 = ( (~ preset)  &  (~ pdn)  &  wire17700 ) ;
 assign wire19080 = ( wire1984 ) | ( wire1981 ) ;
 assign wire19081 = ( wire1985 ) | ( ppeakb_4_4_  &  wire4382 ) ;
 assign wire19083 = ( wire15035  &  wire4369 ) | ( wire4865  &  wire4378 ) ;
 assign wire19084 = ( wire6230  &  wire4341 ) | ( wire14765  &  wire4351 ) ;
 assign wire19085 = ( wire1976 ) | ( wire1978 ) | ( wire1979 ) | ( wire1980 ) ;
 assign wire19094 = ( wire1986 ) | ( wire1987 ) | ( wire19080 ) | ( wire19081 ) ;
 assign wire19095 = ( wire1988 ) | ( wire19083 ) | ( wire19084 ) | ( wire19085 ) ;
 assign wire19100 = ( wire1969 ) | ( wire1966 ) ;
 assign wire19101 = ( wire1970 ) | ( ppeakb_5_5_  &  wire4382 ) ;
 assign wire19102 = ( wire15395  &  wire4369 ) | ( wire9545  &  wire4378 ) ;
 assign wire19104 = ( wire6905  &  wire4341 ) | ( wire8330  &  wire4351 ) ;
 assign wire19105 = ( wire1961 ) | ( wire1963 ) | ( wire1964 ) | ( wire1965 ) ;
 assign wire19110 = ( wire1971 ) | ( wire1972 ) | ( wire19100 ) | ( wire19101 ) ;
 assign wire19111 = ( wire1973 ) | ( wire19102 ) | ( wire19104 ) | ( wire19105 ) ;
 assign wire19115 = ( wire1952 ) | ( wire1949 ) ;
 assign wire19116 = ( wire1953 ) | ( ppeakb_6_6_  &  wire4382 ) ;
 assign wire19117 = ( wire14210  &  wire4369 ) | ( wire8870  &  wire4378 ) ;
 assign wire19118 = ( wire4835  &  wire4341 ) | ( wire7685  &  wire4351 ) ;
 assign wire19119 = ( wire1944 ) | ( wire1946 ) | ( wire1947 ) | ( wire1948 ) ;
 assign wire19124 = ( wire1954 ) | ( wire1955 ) | ( wire19115 ) | ( wire19116 ) ;
 assign wire19125 = ( wire1956 ) | ( wire19117 ) | ( wire19118 ) | ( wire19119 ) ;
 assign wire19126 = ( (~ preset)  &  (~ pdn)  &  wire17596 ) ;
 assign wire19127 = ( (~ preset)  &  n_n2344  &  nrq7_2 ) ;
 assign wire19130 = ( (~ preset)  &  n_n2344  &  nsl8_2  &  nrq7_2 ) ;
 assign wire19132 = ( (~ preset)  &  wire18168  &  n_n2344  &  nrq7_2 ) ;
 assign wire19134 = ( (~ preset)  &  wire17453  &  n_n2344  &  nrq7_2 ) ;
 assign wire19135 = ( (~ ndn7_2)  &  wire19130 ) | ( (~ ndn7_2)  &  wire19132 ) ;
 assign wire19136 = ( (~ ndn7_2)  &  wire19134 ) | ( (~ ndn7_2)  &  (~ nrq8_2)  &  wire19127 ) ;
 assign wire19140 = ( wire1926 ) | ( wire1923 ) ;
 assign wire19141 = ( wire1927 ) | ( ppeakb_7_7_  &  wire4382 ) ;
 assign wire19142 = ( wire14630  &  wire4369 ) | ( wire8225  &  wire4378 ) ;
 assign wire19144 = ( wire5540  &  wire4341 ) | ( wire7055  &  wire4351 ) ;
 assign wire19145 = ( wire1918 ) | ( wire1920 ) | ( wire1921 ) | ( wire1922 ) ;
 assign wire19150 = ( wire1928 ) | ( wire1929 ) | ( wire19140 ) | ( wire19141 ) ;
 assign wire19151 = ( wire1930 ) | ( wire19142 ) | ( wire19144 ) | ( wire19145 ) ;
 assign wire19152 = ( (~ preset)  &  wire18493  &  nrq7_2 ) | ( (~ preset)  &  nrq7_2  &  wire3746 ) ;
 assign wire19154 = ( (~ preset)  &  wire18389  &  nrq7_2 ) | ( (~ preset)  &  wire18415  &  nrq7_2 ) ;
 assign wire19155 = ( (~ preset)  &  wire17388  &  nrq7_2 ) | ( (~ preset)  &  wire18376  &  nrq7_2 ) ;
 assign wire19156 = ( (~ preset)  &  wire17271  &  nrq7_2 ) | ( (~ preset)  &  wire17297  &  nrq7_2 ) ;
 assign wire19158 = ( (~ preset)  &  wire17167  &  nrq7_2 ) | ( (~ preset)  &  wire17232  &  nrq7_2 ) ;
 assign wire19159 = ( (~ preset)  &  wire17050  &  nrq7_2 ) | ( (~ preset)  &  wire17102  &  nrq7_2 ) ;
 assign wire19163 = ( wire1914 ) | ( wire19152 ) | ( wire19159 ) ;
 assign wire19164 = ( wire19154 ) | ( wire19155 ) | ( wire19156 ) | ( wire19158 ) ;


endmodule

