module alu4 (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, 
	i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, o_1_, o_2_, o_0_, o_7_, 
	o_5_, o_6_, o_3_, o_4_);

input i_9_;
input i_10_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_3_;
input i_13_;
input i_4_;
input i_12_;
input i_1_;
input i_11_;
input i_2_;
input i_0_;
output o_1_;
output o_2_;
output o_0_;
output o_7_;
output o_5_;
output o_6_;
output o_3_;
output o_4_;
wire n_n637;
wire n_n860;
wire n_n861;
wire wire8;
wire wire21;
wire wire23;
wire wire414;
wire n_n877;
wire n_n876;
wire n_n878;
wire n_n874;
wire wire18;
wire wire55;
wire wire126;
wire wire278;
wire wire283;
wire wire327;
wire wire343;
wire wire348;
wire wire386;
wire n_n1240;
wire n_n1241;
wire n_n1221;
wire n_n1236;
wire n_n1222;
wire n_n1121;
wire n_n1120;
wire n_n1108;
wire n_n1189;
wire n_n1187;
wire n_n658;
wire n_n741;
wire n_n566;
wire n_n764;
wire n_n701;
wire wire323;
wire wire325;
wire wire326;
wire n_n970;
wire n_n972;
wire n_n978;
wire n_n976;
wire n_n962;
wire n_n955;
wire n_n957;
wire n_n816;
wire n_n853;
wire n_n779;
wire n_n795;
wire wire17;
wire wire33;
wire wire35;
wire wire37;
wire wire68;
wire wire288;
wire wire313;
wire wire322;
wire wire336;
wire wire420;
wire n_n833;
wire n_n538;
wire n_n850;
wire n_n498;
wire n_n838;
wire n_n835;
wire n_n748;
wire n_n725;
wire wire341;
wire n_n665;
wire wire425;
wire wire337;
wire wire430;
wire n_n1245;
wire wire435;
wire wire434;
wire n_n716;
wire n_n849;
wire n_n36;
wire wire438;
wire n_n545;
wire n_n675;
wire wire29;
wire wire289;
wire wire443;
wire wire442;
wire n_n570;
wire n_n787;
wire n_n769;
wire n_n819;
wire n_n273;
wire wire381;
wire wire12;
wire wire377;
wire n_n847;
wire wire27;
wire n_n581;
wire wire264;
wire n_n638;
wire wire15;
wire n_n814;
wire n_n541;
wire wire28;
wire n_n746;
wire wire333;
wire n_n830;
wire n_n453;
wire n_n761;
wire n_n213;
wire n_n421;
wire n_n415;
wire wire344;
wire n_n369;
wire wire25;
wire n_n358;
wire wire14;
wire n_n412;
wire wire279;
wire n_n773;
wire n_n844;
wire wire13;
wire n_n639;
wire wire286;
wire n_n185;
wire n_n432;
wire n_n826;
wire n_n183;
wire wire96;
wire n_n818;
wire n_n153;
wire n_n316;
wire n_n197;
wire n_n843;
wire n_n699;
wire wire293;
wire n_n678;
wire n_n671;
wire wire26;
wire n_n176;
wire n_n712;
wire n_n751;
wire wire265;
wire n_n719;
wire wire31;
wire n_n687;
wire wire34;
wire n_n827;
wire n_n685;
wire wire309;
wire wire267;
wire n_n683;
wire n_n275;
wire n_n792;
wire n_n35;
wire wire69;
wire wire70;
wire wire106;
wire wire450;
wire n_n1261;
wire wire454;
wire wire453;
wire n_n1248;
wire n_n752;
wire wire307;
wire n_n635;
wire n_n592;
wire n_n832;
wire n_n852;
wire n_n1243;
wire n_n609;
wire wire465;
wire n_n598;
wire n_n575;
wire wire19;
wire wire9;
wire n_n672;
wire n_n810;
wire wire32;
wire wire370;
wire wire371;
wire wire295;
wire wire301;
wire wire346;
wire wire11;
wire n_n633;
wire n_n653;
wire n_n526;
wire n_n534;
wire n_n242;
wire n_n656;
wire n_n194;
wire n_n346;
wire n_n842;
wire wire281;
wire n_n791;
wire n_n755;
wire n_n846;
wire n_n1258;
wire n_n670;
wire wire113;
wire n_n756;
wire n_n550;
wire n_n732;
wire wire284;
wire wire483;
wire wire482;
wire wire118;
wire wire487;
wire wire486;
wire wire485;
wire n_n1126;
wire wire22;
wire wire38;
wire wire297;
wire n_n1127;
wire wire493;
wire wire491;
wire n_n1112;
wire wire268;
wire n_n274;
wire n_n837;
wire n_n240;
wire wire330;
wire n_n771;
wire n_n606;
wire n_n813;
wire wire290;
wire wire308;
wire wire318;
wire wire494;
wire wire360;
wire wire497;
wire n_n1250;
wire wire294;
wire wire296;
wire wire502;
wire wire501;
wire wire272;
wire wire298;
wire wire311;
wire wire363;
wire n_n1129;
wire wire104;
wire wire270;
wire wire379;
wire wire507;
wire n_n1123;
wire n_n623;
wire wire181;
wire wire364;
wire wire512;
wire wire516;
wire wire513;
wire wire300;
wire wire269;
wire n_n822;
wire n_n840;
wire n_n631;
wire n_n710;
wire n_n729;
wire wire519;
wire wire518;
wire wire517;
wire n_n1256;
wire n_n735;
wire wire523;
wire wire521;
wire n_n1231;
wire wire350;
wire wire529;
wire wire16;
wire wire533;
wire wire536;
wire wire277;
wire n_n597;
wire n_n651;
wire n_n1255;
wire wire405;
wire wire545;
wire wire544;
wire wire543;
wire n_n1253;
wire wire120;
wire n_n1229;
wire wire553;
wire wire552;
wire n_n1128;
wire wire30;
wire wire352;
wire wire557;
wire wire338;
wire wire560;
wire wire558;
wire n_n1000;
wire wire565;
wire wire564;
wire n_n503;
wire wire73;
wire wire121;
wire wire571;
wire n_n1233;
wire wire574;
wire n_n624;
wire wire20;
wire wire579;
wire wire578;
wire n_n619;
wire wire583;
wire wire581;
wire n_n1234;
wire wire591;
wire n_n851;
wire wire594;
wire wire593;
wire wire123;
wire wire276;
wire wire291;
wire wire354;
wire wire596;
wire n_n277;
wire wire115;
wire wire410;
wire wire604;
wire wire606;
wire n_n1264;
wire n_n1265;
wire wire292;
wire wire340;
wire wire359;
wire wire402;
wire wire612;
wire n_n1191;
wire n_n1185;
wire wire351;
wire wire369;
wire wire617;
wire wire616;
wire wire314;
wire wire365;
wire wire619;
wire n_n612;
wire wire275;
wire wire626;
wire wire628;
wire n_n768;
wire wire632;
wire wire639;
wire wire638;
wire wire637;
wire wire41;
wire wire382;
wire wire641;
wire wire324;
wire n_n910;
wire wire648;
wire wire299;
wire wire316;
wire wire376;
wire wire395;
wire wire36;
wire wire304;
wire wire384;
wire wire385;
wire wire347;
wire wire356;
wire wire655;
wire n_n991;
wire wire660;
wire n_n879;
wire wire287;
wire wire388;
wire n_n881;
wire wire668;
wire wire667;
wire wire666;
wire wire669;
wire wire671;
wire wire406;
wire wire676;
wire wire403;
wire wire334;
wire wire380;
wire wire686;
wire wire685;
wire n_n993;
wire n_n913;
wire wire696;
wire n_n906;
wire wire397;
wire wire701;
wire wire700;
wire wire321;
wire wire704;
wire wire703;
wire wire706;
wire wire705;
wire wire708;
wire n_n987;
wire wire366;
wire wire717;
wire wire716;
wire n_n965;
wire n_n981;
wire n_n984;
wire n_n983;
wire wire725;
wire wire724;
wire wire723;
wire wire374;
wire n_n986;
wire wire24;
wire wire735;
wire wire737;
wire wire736;
wire wire342;
wire wire738;
wire wire744;
wire wire747;
wire wire746;
wire wire751;
wire wire752;
wire wire263;
wire wire762;
wire wire761;
wire wire54;
wire wire10;
wire wire42;
wire wire51;
wire wire317;
wire wire319;
wire wire329;
wire wire335;
wire wire375;
wire wire393;
wire wire424;
wire wire423;
wire wire427;
wire wire426;
wire wire429;
wire wire428;
wire wire436;
wire wire440;
wire wire439;
wire wire447;
wire wire451;
wire wire452;
wire wire459;
wire wire469;
wire wire468;
wire wire479;
wire wire484;
wire wire503;
wire wire515;
wire wire520;
wire wire525;
wire wire524;
wire wire530;
wire wire531;
wire wire541;
wire wire546;
wire wire551;
wire wire562;
wire wire561;
wire wire569;
wire wire573;
wire wire572;
wire wire576;
wire wire584;
wire wire615;
wire wire622;
wire wire633;
wire wire636;
wire wire635;
wire wire644;
wire wire643;
wire wire646;
wire wire649;
wire wire653;
wire wire657;
wire wire673;
wire wire677;
wire wire680;
wire wire683;
wire wire684;
wire wire689;
wire wire698;
wire wire707;
wire wire712;
wire wire719;
wire wire718;
wire wire726;
wire wire728;
wire wire734;
wire wire741;
wire wire763;
wire wire40;
wire wire50;
wire wire52;
wire wire57;
wire wire59;
wire wire60;
wire wire62;
wire wire63;
wire wire64;
wire wire65;
wire wire80;
wire wire81;
wire wire82;
wire wire83;
wire wire84;
wire wire86;
wire wire89;
wire wire95;
wire wire97;
wire wire98;
wire wire103;
wire wire107;
wire wire112;
wire wire127;
wire wire128;
wire wire129;
wire wire130;
wire wire136;
wire wire139;
wire wire141;
wire wire142;
wire wire143;
wire wire144;
wire wire145;
wire wire150;
wire wire154;
wire wire156;
wire wire163;
wire wire166;
wire wire170;
wire wire171;
wire wire172;
wire wire176;
wire wire180;
wire wire182;
wire wire190;
wire wire192;
wire wire194;
wire wire198;
wire wire200;
wire wire201;
wire wire206;
wire wire207;
wire wire208;
wire wire212;
wire wire213;
wire wire215;
wire wire222;
wire wire223;
wire wire224;
wire wire225;
wire wire230;
wire wire231;
wire wire235;
wire wire236;
wire wire237;
wire wire238;
wire wire241;
wire wire245;
wire wire246;
wire wire247;
wire wire249;
wire wire252;
wire wire253;
wire wire255;
wire wire256;
wire wire258;
wire wire362;
wire wire373;
wire wire411;
wire wire768;
wire wire769;
wire wire772;
wire wire773;
wire wire777;
wire wire779;
wire wire784;
wire wire785;
wire wire788;
wire wire790;
wire wire791;
wire wire795;
wire wire798;
wire wire800;
wire wire801;
wire wire802;
wire wire808;
wire wire809;
wire wire814;
wire wire824;
wire wire825;
wire wire834;
wire wire835;
wire wire836;
wire wire837;
wire wire840;
wire wire841;
wire wire842;
wire wire843;
wire wire844;
wire wire845;
wire wire846;
wire wire850;
wire wire852;
wire wire853;
wire wire854;
wire wire855;
wire wire856;
wire wire857;
wire wire859;
wire wire863;
wire wire864;
wire wire879;
wire wire881;
wire wire882;
wire wire883;
wire wire884;
wire wire885;
wire wire887;
wire wire891;
wire wire895;
wire wire896;
wire wire901;
wire wire903;
wire wire905;
wire wire907;
wire wire909;
wire wire912;
wire wire917;
wire wire925;
wire wire927;
wire wire931;
wire wire932;
wire wire934;
wire wire937;
wire wire939;
wire wire947;
wire wire948;
wire wire949;
wire wire951;
wire wire954;
wire wire957;
wire wire958;
wire wire960;
wire wire961;
wire wire962;
wire wire970;
wire wire971;
wire wire972;
wire wire979;
wire wire981;
wire wire987;
wire wire988;
wire wire993;
wire wire995;
wire wire1003;
wire wire1005;
wire wire1009;
wire wire1011;
wire wire1012;
wire wire1017;
wire wire1019;
wire wire1021;
wire wire1023;
wire wire1024;
wire wire1026;
wire wire1027;
wire wire1030;
wire wire1033;
wire wire1040;
wire wire1041;
wire wire1042;
wire wire1043;
wire wire1044;
wire wire1047;
wire wire1064;
wire wire1067;
wire wire1074;
wire wire1076;
wire wire1082;
wire wire1083;
wire wire1087;
wire wire1089;
wire wire1092;
wire wire1093;
wire wire1094;
wire wire1096;
wire wire1097;
wire wire1103;
wire wire1108;
wire wire1109;
wire wire1110;
wire wire1115;
wire wire1116;
wire wire1117;
wire wire1119;
wire wire1121;
wire wire1122;
wire wire1123;
wire wire1130;
wire wire1132;
wire wire1133;
wire wire1134;
wire wire1135;
wire wire1139;
wire wire1143;
wire wire1152;
wire wire1154;
wire wire1156;
wire wire1160;
wire wire1162;
wire wire1165;
wire wire1166;
wire wire1168;
wire wire1169;
wire wire1171;
wire wire1173;
wire wire1175;
wire wire1180;
wire wire1181;
wire wire1182;
wire wire1183;
wire wire1186;
wire wire1194;
wire wire1195;
wire wire1196;
wire wire1198;
wire wire1199;
wire wire1200;
wire wire1202;
wire wire1203;
wire wire1204;
wire wire1213;
wire wire1214;
wire wire1215;
wire wire1216;
wire wire1217;
wire wire1218;
wire wire1221;
wire wire1228;
wire wire1229;
wire wire1230;
wire wire1234;
wire wire1235;
wire wire1239;
wire wire1245;
wire wire1246;
wire wire1247;
wire wire1248;
wire wire1249;
wire wire1250;
wire wire1252;
wire wire1255;
wire wire1263;
wire wire1266;
wire wire1267;
wire wire1272;
wire wire1274;
wire wire1277;
wire wire1279;
wire wire1283;
wire wire1290;
wire wire1293;
wire wire1294;
wire wire1295;
wire wire1296;
wire wire1297;
wire wire1298;
wire wire1299;
wire wire1300;
wire wire1301;
wire wire1302;
wire wire1307;
wire wire1308;
wire wire1314;
wire wire1315;
wire wire1316;
wire wire1317;
wire wire1321;
wire wire1324;
wire wire1326;
wire wire1327;
wire wire1328;
wire wire1329;
wire wire1331;
wire wire1332;
wire wire1333;
wire wire1334;
wire wire1336;
wire wire1337;
wire wire1338;
wire wire1339;
wire wire1340;
wire wire1341;
wire wire1343;
wire wire1344;
wire wire1346;
wire wire1348;
wire wire1350;
wire wire1351;
wire wire1352;
wire wire1353;
wire wire1354;
wire wire1355;
wire wire1361;
wire wire1362;
wire wire1363;
wire wire1366;
wire wire1372;
wire wire1373;
wire wire1375;
wire wire1376;
wire wire1377;
wire wire1383;
wire wire1385;
wire wire1388;
wire wire1390;
wire wire1391;
wire wire1392;
wire wire1393;
wire wire1394;
wire wire1396;
wire wire1397;
wire wire1400;
wire wire1402;
wire wire1403;
wire wire1406;
wire wire1408;
wire wire1409;
wire wire1410;
wire wire1412;
wire wire1414;
wire wire1416;
wire wire1418;
wire wire1419;
wire wire1423;
wire wire1425;
wire wire1432;
wire wire1433;
wire wire1436;
wire wire1437;
wire wire1438;
wire wire1440;
wire wire1441;
wire wire1444;
wire wire1446;
wire wire1447;
wire wire1450;
wire wire1453;
wire wire1454;
wire wire1462;
wire wire1463;
wire wire1464;
wire wire1466;
wire wire1472;
wire wire1474;
wire wire1480;
wire wire1481;
wire wire1488;
wire wire1490;
wire wire1493;
wire wire1500;
wire wire1501;
wire wire1502;
wire wire1503;
wire wire1504;
wire wire1506;
wire wire1511;
wire wire1517;
wire wire1524;
wire wire1525;
wire wire1526;
wire wire1527;
wire wire1528;
wire wire1529;
wire wire1530;
wire wire1534;
wire wire1535;
wire wire1537;
wire wire1538;
wire wire1539;
wire wire1542;
wire wire1543;
wire wire1547;
wire wire1552;
wire wire1553;
wire wire1554;
wire wire1555;
wire wire1558;
wire wire1562;
wire wire1563;
wire wire1564;
wire wire1565;
wire wire1569;
wire wire1571;
wire wire1572;
wire wire1574;
wire wire1575;
wire wire1582;
wire wire1583;
wire wire1584;
wire wire1585;
wire wire1587;
wire wire1588;
wire wire1596;
wire wire1603;
wire wire1605;
wire wire1609;
wire wire1610;
wire wire1611;
wire wire1612;
wire wire1613;
wire wire1614;
wire wire1620;
wire wire1624;
wire wire1629;
wire wire1630;
wire wire1634;
wire wire1635;
wire wire1637;
wire wire1639;
wire wire1640;
wire wire1643;
wire wire1644;
wire wire1647;
wire wire1648;
wire wire1652;
wire wire1656;
wire wire1661;
wire wire1663;
wire wire1669;
wire wire1672;
wire wire1673;
wire wire1675;
wire wire1679;
wire wire1681;
wire wire1684;
wire wire1685;
wire wire1686;
wire wire1689;
wire wire1691;
wire wire1692;
wire wire1694;
wire wire1699;
wire wire1702;
wire wire1703;
wire wire1704;
wire wire1705;
wire wire1708;
wire wire1709;
wire wire1712;
wire wire1713;
wire wire1720;
wire wire1721;
wire wire1722;
wire wire1723;
wire wire1724;
wire wire1725;
wire wire1726;
wire wire1729;
wire wire1732;
wire wire1740;
wire wire1741;
wire wire1744;
wire wire1746;
wire wire1748;
wire wire1750;
wire wire1756;
wire wire1763;
wire wire1764;
wire wire1765;
wire wire1766;
wire wire1767;
wire wire1768;
wire wire1770;
wire wire1776;
wire wire1778;
wire wire1779;
wire wire1780;
wire wire1781;
wire wire1789;
wire wire1792;
wire wire1794;
wire wire1796;
wire wire1797;
wire wire1798;
wire wire1799;
wire wire1803;
wire wire1804;
wire wire1805;
wire wire1806;
wire wire1808;
wire wire1810;
wire wire1814;
wire wire1816;
wire wire1817;
wire wire1820;
wire wire1821;
wire wire1823;
wire wire1825;
wire wire1829;
wire wire1832;
wire wire1833;
wire wire1838;
wire wire1839;
wire wire1841;
wire wire1844;
wire wire1845;
wire wire1848;
wire wire1849;
wire wire1850;
wire wire1852;
wire wire1853;
wire wire1856;
wire wire1857;
wire wire1861;
wire wire1863;
wire wire1867;
wire wire1869;
wire wire6473;
wire wire6474;
wire wire6475;
wire wire6478;
wire wire6479;
wire wire6485;
wire wire6488;
wire wire6491;
wire wire6493;
wire wire6494;
wire wire6495;
wire wire6496;
wire wire6499;
wire wire6500;
wire wire6501;
wire wire6504;
wire wire6506;
wire wire6507;
wire wire6509;
wire wire6510;
wire wire6512;
wire wire6515;
wire wire6516;
wire wire6517;
wire wire6520;
wire wire6522;
wire wire6523;
wire wire6524;
wire wire6526;
wire wire6527;
wire wire6528;
wire wire6530;
wire wire6536;
wire wire6537;
wire wire6538;
wire wire6549;
wire wire6550;
wire wire6551;
wire wire6553;
wire wire6554;
wire wire6555;
wire wire6557;
wire wire6558;
wire wire6559;
wire wire6561;
wire wire6562;
wire wire6563;
wire wire6567;
wire wire6573;
wire wire6575;
wire wire6577;
wire wire6578;
wire wire6579;
wire wire6582;
wire wire6584;
wire wire6585;
wire wire6587;
wire wire6588;
wire wire6589;
wire wire6591;
wire wire6593;
wire wire6594;
wire wire6595;
wire wire6598;
wire wire6600;
wire wire6603;
wire wire6604;
wire wire6605;
wire wire6615;
wire wire6616;
wire wire6618;
wire wire6620;
wire wire6621;
wire wire6622;
wire wire6623;
wire wire6624;
wire wire6627;
wire wire6628;
wire wire6629;
wire wire6630;
wire wire6631;
wire wire6632;
wire wire6633;
wire wire6636;
wire wire6637;
wire wire6638;
wire wire6640;
wire wire6642;
wire wire6643;
wire wire6644;
wire wire6645;
wire wire6647;
wire wire6651;
wire wire6653;
wire wire6654;
wire wire6658;
wire wire6660;
wire wire6661;
wire wire6665;
wire wire6667;
wire wire6669;
wire wire6670;
wire wire6672;
wire wire6673;
wire wire6674;
wire wire6675;
wire wire6678;
wire wire6683;
wire wire6686;
wire wire6687;
wire wire6688;
wire wire6693;
wire wire6694;
wire wire6698;
wire wire6702;
wire wire6704;
wire wire6708;
wire wire6709;
wire wire6712;
wire wire6713;
wire wire6714;
wire wire6715;
wire wire6719;
wire wire6725;
wire wire6730;
wire wire6731;
wire wire6735;
wire wire6737;
wire wire6745;
wire wire6748;
wire wire6749;
wire wire6750;
wire wire6752;
wire wire6755;
wire wire6756;
wire wire6757;
wire wire6759;
wire wire6762;
wire wire6763;
wire wire6764;
wire wire6766;
wire wire6770;
wire wire6771;
wire wire6772;
wire wire6773;
wire wire6775;
wire wire6776;
wire wire6777;
wire wire6780;
wire wire6782;
wire wire6785;
wire wire6787;
wire wire6788;
wire wire6789;
wire wire6791;
wire wire6794;
wire wire6799;
wire wire6803;
wire wire6805;
wire wire6806;
wire wire6807;
wire wire6811;
wire wire6812;
wire wire6814;
wire wire6816;
wire wire6819;
wire wire6820;
wire wire6821;
wire wire6823;
wire wire6824;
wire wire6825;
wire wire6827;
wire wire6828;
wire wire6831;
wire wire6834;
wire wire6835;
wire wire6837;
wire wire6838;
wire wire6840;
wire wire6842;
wire wire6843;
wire wire6846;
wire wire6848;
wire wire6850;
wire wire6852;
wire wire6853;
wire wire6854;
wire wire6857;
wire wire6858;
wire wire6860;
wire wire6864;
wire wire6865;
wire wire6868;
wire wire6869;
wire wire6870;
wire wire6871;
wire wire6872;
wire wire6873;
wire wire6875;
wire wire6876;
wire wire6879;
wire wire6884;
wire wire6885;
wire wire6886;
wire wire6887;
wire wire6888;
wire wire6890;
wire wire6893;
wire wire6894;
wire wire6896;
wire wire6897;
wire wire6899;
wire wire6900;
wire wire6901;
wire wire6902;
wire wire6904;
wire wire6905;
wire wire6906;
wire wire6908;
wire wire6911;
wire wire6913;
wire wire6914;
wire wire6915;
wire wire6916;
wire wire6918;
wire wire6919;
wire wire6920;
wire wire6921;
wire wire6922;
wire wire6923;
wire wire6924;
wire wire6925;
wire wire6926;
wire wire6929;
wire wire6930;
wire wire6931;
wire wire6934;
wire wire6937;
wire wire6938;
wire wire6941;
wire wire6942;
wire wire6943;
wire wire6944;
wire wire6945;
wire wire6946;
wire wire6949;
wire wire6950;
wire wire6952;
wire wire6954;
wire wire6955;
wire wire6956;
wire wire6958;
wire wire6959;
wire wire6961;
wire wire6963;
wire wire6964;
wire wire6965;
wire wire6966;
wire wire6967;
wire wire6968;
wire wire6969;
wire wire6970;
wire wire6972;
wire wire6973;
wire wire6975;
wire wire6976;
wire wire6978;
wire wire6979;
wire wire6982;
wire wire6983;
wire wire6984;
wire wire6985;
wire wire6987;
wire wire6991;
wire wire6992;
wire wire6994;
wire wire6995;
wire wire6996;
wire wire6997;
wire wire6999;
wire wire7001;
wire wire7003;
wire wire7004;
wire wire7005;
wire wire7007;
wire wire7008;
wire wire7009;
wire wire7010;
wire wire7011;
wire wire7013;
wire wire7015;
wire wire7017;
wire wire7018;
wire wire7019;
wire wire7021;
wire wire7022;
wire wire7023;
wire wire7024;
wire wire7027;
wire wire7028;
wire wire7029;
wire wire7030;
wire wire7032;
wire wire7033;
wire wire7035;
wire wire7037;
wire wire7038;
wire wire7039;
wire wire7040;
wire wire7041;
wire wire7042;
wire wire7043;
wire wire7045;
wire wire7046;
wire wire7047;
wire wire7050;
wire wire7051;
wire wire7054;
wire wire7057;
wire wire7058;
wire wire7059;
wire wire7060;
wire wire7062;
wire wire7063;
wire wire7065;
wire wire7066;
wire wire7067;
wire wire7068;
wire wire7070;
wire wire7071;
wire wire7074;
wire wire7076;
wire wire7077;
wire wire7078;
wire wire7079;
wire wire7080;
wire wire7082;
wire wire7083;
wire wire7084;
wire wire7085;
wire wire7086;
wire wire7087;
wire wire7088;
wire wire7091;
wire wire7092;
wire wire7093;
wire wire7094;
wire wire7100;
wire wire7102;
wire wire7104;
wire wire7105;
wire wire7107;
wire wire7108;
wire wire7109;
wire wire7110;
wire wire7111;
wire wire7113;
wire wire7114;
wire wire7115;
wire wire7117;
wire wire7118;
wire wire7119;
wire wire7121;
wire wire7122;
wire wire7126;
wire wire7127;
wire wire7128;
wire wire7129;
wire wire7130;
wire wire7132;
wire wire7133;
wire wire7134;
wire wire7136;
wire wire7138;
wire wire7140;
wire wire7144;
wire wire7146;
wire wire7149;
wire wire7151;
wire wire7155;
wire wire7157;
wire wire7161;
wire wire7163;
wire wire7164;
wire wire7165;
wire wire7167;
wire wire7168;
wire wire7174;
wire wire7175;
wire wire7177;
wire wire7178;
wire wire7181;
wire wire7182;
wire wire7183;
wire wire7184;
wire wire7185;
wire wire7188;
wire wire7190;
wire wire7191;
wire wire7194;
wire wire7196;
wire wire7199;
wire wire7200;
wire wire7202;
wire wire7203;
wire wire7205;
wire wire7208;
wire wire7211;
wire wire7214;
wire wire7215;
wire wire7218;
wire wire7219;
wire wire7222;
wire wire7223;
wire wire7226;
wire wire7227;
wire wire7228;
wire wire7229;
wire wire7231;
wire wire7232;
wire wire7233;
wire wire7234;
wire wire7235;
wire wire7237;
wire wire7239;
wire wire7241;
wire wire7244;
wire wire7246;
wire wire7248;
wire wire7249;
wire wire7250;
wire wire7251;
wire wire7253;
wire wire7254;
wire wire7255;
wire wire7257;
wire wire7260;
wire wire7261;
wire wire7262;
wire wire7263;
wire wire7264;
wire wire7266;
wire wire7267;
wire wire7268;
wire wire7269;
wire wire7271;
wire wire7272;
wire wire7273;
wire wire7275;
wire wire7277;
wire wire7278;
wire wire7279;
wire wire7280;
wire wire7282;
wire wire7286;
wire wire7287;
wire wire7288;
wire wire7289;
wire wire7292;
wire wire7293;
wire wire7294;
wire wire7295;
wire wire7296;
wire wire7297;
wire wire7300;
wire wire7302;
wire wire7303;
wire wire7304;
wire wire7307;
wire wire7308;
wire wire7309;
wire wire7310;
wire wire7311;
wire wire7312;
wire wire7313;
wire wire7314;
wire wire7317;
wire wire7318;
wire wire7319;
wire wire7321;
wire wire7322;
wire wire7324;
wire wire7325;
wire wire7326;
wire wire7327;
wire wire7329;
wire wire7335;
wire wire7336;
wire wire7337;
wire wire7338;
wire wire7339;
assign o_1_ = ( n_n860 ) | ( n_n861 ) | ( wire1852 ) | ( wire6485 ) ;
 assign o_2_ = ( n_n874 ) | ( wire1789 ) | ( wire6528 ) | ( wire6530 ) ;
 assign o_0_ = ( wire6536 ) | ( wire6537 ) | ( wire6538 ) ;
 assign o_7_ = ( n_n1221 ) | ( n_n1222 ) | ( wire6827 ) | ( wire6828 ) ;
 assign o_5_ = ( wire6937 ) | ( wire6938 ) | ( wire6949 ) | ( wire6950 ) ;
 assign o_6_ = ( n_n1185 ) | ( wire6975 ) | ( wire7001 ) ;
 assign o_3_ = ( n_n906 ) | ( wire7065 ) | ( wire7076 ) ;
 assign o_4_ = ( n_n955 ) | ( wire7337 ) | ( wire7338 ) | ( wire7339 ) ;
 assign n_n637 = ( i_13_  &  (~ i_11_) ) ;
 assign n_n860 = ( wire1867 ) | ( wire1869 ) | ( wire6474 ) | ( wire6475 ) ;
 assign n_n861 = ( wire1861 ) | ( wire6479 ) | ( (~ i_3_)  &  wire747 ) ;
 assign wire8 = ( i_9_  &  i_10_ ) ;
 assign wire21 = ( i_3_  &  (~ i_4_) ) ;
 assign wire23 = ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire414 = ( i_9_  &  i_10_ ) | ( i_9_  &  i_8_ ) | ( i_10_  &  (~ i_8_) ) ;
 assign n_n877 = ( wire1841 ) | ( wire6491 ) | ( (~ i_5_)  &  wire648 ) ;
 assign n_n876 = ( wire1832 ) | ( wire1833 ) | ( wire6495 ) | ( wire6496 ) ;
 assign n_n878 = ( wire1823 ) | ( wire1825 ) | ( wire6500 ) | ( wire6501 ) ;
 assign n_n874 = ( n_n879 ) | ( n_n881 ) | ( wire6520 ) ;
 assign wire18 = ( i_9_  &  i_8_ ) ;
 assign wire55 = ( i_3_ ) | ( i_2_ ) ;
 assign wire126 = ( i_10_  &  (~ i_8_)  &  i_3_ ) ;
 assign wire278 = ( i_10_  &  (~ i_8_) ) ;
 assign wire283 = ( i_9_  &  i_1_ ) ;
 assign wire327 = ( (~ i_6_)  &  i_3_  &  i_2_  &  i_0_ ) ;
 assign wire343 = ( i_9_  &  i_5_  &  i_0_ ) ;
 assign wire348 = ( i_10_  &  (~ i_5_)  &  i_0_ ) ;
 assign wire386 = ( i_9_  &  i_7_  &  i_2_ ) ;
 assign n_n1240 = ( wire6615 ) | ( wire6616 ) | ( wire284  &  wire483 ) ;
 assign n_n1241 = ( wire6627 ) | ( wire344  &  wire502  &  wire6594 ) ;
 assign n_n1221 = ( n_n1248 ) | ( n_n1229 ) | ( wire1547 ) | ( wire6704 ) ;
 assign n_n1236 = ( wire1535 ) | ( wire1537 ) | ( wire6715 ) ;
 assign n_n1222 = ( n_n1261 ) | ( n_n1231 ) | ( n_n1233 ) | ( wire6791 ) ;
 assign n_n1121 = ( wire1375 ) | ( wire1376 ) | ( wire6834 ) ;
 assign n_n1120 = ( wire1362 ) | ( wire1363 ) | ( wire1366 ) | ( wire6840 ) ;
 assign n_n1108 = ( wire1186 ) | ( wire1195 ) | ( wire6941 ) | ( wire6946 ) ;
 assign n_n1189 = ( wire6956 ) | ( wire14  &  wire6954 ) | ( wire14  &  wire6955 ) ;
 assign n_n1187 = ( wire1096 ) | ( wire1097 ) | ( wire6997 ) ;
 assign n_n658 = ( i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign n_n741 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n566 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_12_) ) ;
 assign n_n764 = ( (~ i_9_)  &  i_7_  &  i_8_ ) ;
 assign n_n701 = ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire323 = ( (~ i_5_)  &  (~ i_1_) ) ;
 assign wire325 = ( i_6_  &  (~ i_1_) ) ;
 assign wire326 = ( (~ i_6_)  &  (~ i_1_) ) ;
 assign n_n970 = ( wire947 ) | ( wire949 ) | ( wire7088 ) ;
 assign n_n972 = ( wire937 ) | ( i_0_  &  wire939 ) | ( i_0_  &  wire7093 ) ;
 assign n_n978 = ( wire925 ) | ( wire7102 ) | ( wire20  &  wire578 ) ;
 assign n_n976 = ( wire881 ) | ( wire882 ) | ( wire883 ) | ( wire884 ) ;
 assign n_n962 = ( n_n984 ) | ( n_n983 ) | ( wire7167 ) | ( wire7168 ) ;
 assign n_n955 = ( n_n965 ) | ( wire7232 ) | ( wire7233 ) | ( wire7244 ) ;
 assign n_n957 = ( wire40 ) | ( wire50 ) | ( wire52 ) | ( wire7329 ) ;
 assign n_n816 = ( (~ i_10_)  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n853 = ( (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign n_n779 = ( i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n795 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire17 = ( (~ i_13_)  &  i_4_  &  i_12_  &  i_11_ ) ;
 assign wire33 = ( i_1_  &  i_2_ ) ;
 assign wire35 = ( (~ i_5_)  &  i_4_ ) ;
 assign wire37 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign wire68 = ( (~ i_10_)  &  (~ i_8_)  &  wire17  &  n_n835 ) ;
 assign wire288 = ( (~ i_8_)  &  (~ i_5_) ) ;
 assign wire313 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign wire322 = ( (~ i_9_)  &  i_8_  &  i_5_  &  i_6_ ) ;
 assign wire336 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire420 = ( (~ i_6_)  &  (~ i_2_)  &  i_0_ ) | ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n833 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n538 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n850 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n498 = ( i_10_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign n_n838 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n835 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n748 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n725 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire341 = ( i_9_  &  (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign n_n665 = ( i_13_  &  (~ i_12_) ) ;
 assign wire425 = ( wire1756 ) | ( wire6555 ) | ( i_7_  &  wire427 ) ;
 assign wire337 = ( i_9_  &  i_10_  &  wire6557 ) ;
 assign wire430 = ( wire1746 ) | ( n_n609  &  wire6561 ) | ( n_n609  &  wire6562 ) ;
 assign n_n1245 = ( wire1744 ) | ( i_13_  &  (~ i_12_)  &  wire430 ) ;
 assign wire435 = ( n_n619  &  wire376 ) | ( n_n623  &  wire436 ) ;
 assign wire434 = ( n_n833  &  n_n633 ) | ( n_n830  &  n_n631 ) ;
 assign n_n716 = ( (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign n_n849 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n36 = ( (~ i_8_)  &  i_11_ ) ;
 assign wire438 = ( n_n779  &  wire309 ) | ( n_n685  &  wire439 ) ;
 assign n_n545 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign n_n675 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire29 = ( i_7_  &  (~ i_2_) ) ;
 assign wire289 = ( (~ i_8_)  &  i_6_ ) ;
 assign wire443 = ( n_n675  &  wire295 ) | ( n_n792  &  wire6837 ) ;
 assign wire442 = ( n_n779  &  wire289 ) | ( n_n685  &  wire269 ) ;
 assign n_n570 = ( (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n787 = ( (~ i_13_)  &  i_11_ ) ;
 assign n_n769 = ( (~ i_9_)  &  i_8_  &  i_6_ ) ;
 assign n_n819 = ( (~ i_9_)  &  i_7_  &  i_6_ ) ;
 assign n_n273 = ( (~ i_3_)  &  i_1_  &  (~ i_2_) ) ;
 assign wire381 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire12 = ( i_5_  &  i_6_ ) ;
 assign wire377 = ( (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n847 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire27 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n581 = ( i_9_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire264 = ( i_1_  &  i_0_ ) ;
 assign n_n638 = ( i_9_  &  i_7_  &  i_8_ ) ;
 assign wire15 = ( i_3_  &  i_1_ ) ;
 assign n_n814 = ( i_3_  &  i_1_  &  i_2_ ) ;
 assign n_n541 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire28 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n746 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire333 = ( i_1_  &  (~ i_0_) ) ;
 assign n_n830 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n453 = ( i_10_  &  (~ i_11_) ) ;
 assign n_n761 = ( (~ i_13_)  &  i_12_ ) ;
 assign n_n213 = ( i_10_  &  i_11_ ) ;
 assign n_n421 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign n_n415 = ( i_10_  &  i_12_  &  i_11_ ) ;
 assign wire344 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign n_n369 = ( i_3_  &  (~ i_4_)  &  i_1_ ) ;
 assign wire25 = ( i_9_  &  i_7_ ) ;
 assign n_n358 = ( i_9_  &  i_7_  &  i_6_ ) ;
 assign wire14 = ( (~ i_4_)  &  i_2_ ) ;
 assign n_n412 = ( i_3_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire279 = ( (~ i_10_)  &  (~ i_6_) ) ;
 assign n_n773 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n844 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire13 = ( i_5_  &  (~ i_6_) ) ;
 assign n_n639 = ( i_5_  &  (~ i_6_)  &  i_3_ ) ;
 assign wire286 = ( i_7_  &  i_8_ ) ;
 assign n_n185 = ( i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign n_n432 = ( i_9_  &  i_10_  &  i_12_ ) ;
 assign n_n826 = ( i_3_  &  i_1_  &  i_0_ ) ;
 assign n_n183 = ( i_9_  &  i_12_ ) ;
 assign wire96 = ( (~ i_3_) ) | ( (~ i_2_) ) ;
 assign n_n818 = ( i_3_  &  i_2_  &  i_0_ ) ;
 assign n_n153 = ( i_3_  &  (~ i_4_)  &  i_0_ ) ;
 assign n_n316 = ( i_12_  &  (~ i_11_) ) ;
 assign n_n197 = ( i_9_  &  i_11_ ) ;
 assign n_n843 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n699 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_6_) ) ;
 assign wire293 = ( (~ i_3_)  &  i_4_ ) ;
 assign n_n678 = ( (~ i_3_)  &  i_4_  &  (~ i_0_) ) ;
 assign n_n671 = ( (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire26 = ( (~ i_5_)  &  i_6_ ) ;
 assign n_n176 = ( i_8_  &  (~ i_5_)  &  i_6_ ) ;
 assign n_n712 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n751 = ( (~ i_9_)  &  (~ i_13_) ) ;
 assign wire265 = ( (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n719 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire31 = ( (~ i_3_)  &  (~ i_1_) ) ;
 assign n_n687 = ( (~ i_3_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire34 = ( i_7_  &  i_5_ ) ;
 assign n_n827 = ( (~ i_9_)  &  i_7_  &  i_5_ ) ;
 assign n_n685 = ( (~ i_3_)  &  i_4_  &  (~ i_1_) ) ;
 assign wire309 = ( (~ i_9_)  &  i_8_ ) ;
 assign wire267 = ( (~ i_9_)  &  i_7_ ) ;
 assign n_n683 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n275 = ( (~ i_9_)  &  i_7_  &  (~ i_8_) ) ;
 assign n_n792 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n35 = ( i_8_  &  i_12_ ) ;
 assign wire69 = ( (~ i_6_)  &  (~ i_0_)  &  wire17  &  n_n792 ) ;
 assign wire70 = ( (~ i_5_)  &  (~ i_6_)  &  n_n792  &  wire370 ) ;
 assign wire106 = ( n_n853  &  n_n792  &  n_n791 ) ;
 assign wire450 = ( n_n853  &  wire6735 ) | ( i_4_  &  wire323  &  n_n853 ) ;
 assign n_n1261 = ( wire1511 ) | ( wire6737 ) | ( n_n792  &  wire450 ) ;
 assign wire454 = ( wire1652 ) | ( n_n637  &  wire1656 ) | ( n_n637  &  wire6633 ) ;
 assign wire453 = ( i_0_  &  n_n639  &  wire265 ) | ( (~ i_0_)  &  wire265  &  n_n635 ) ;
 assign n_n1248 = ( wire1647 ) | ( wire1648 ) | ( n_n638  &  wire454 ) ;
 assign n_n752 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign wire307 = ( i_9_  &  i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n635 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_ ) ;
 assign n_n592 = ( i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n832 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n852 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n1243 = ( wire6587 ) | ( n_n665  &  wire1712 ) | ( n_n665  &  wire1713 ) ;
 assign n_n609 = ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire465 = ( wire388 ) | ( wire42 ) | ( wire6591 ) ;
 assign n_n598 = ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign n_n575 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire19 = ( i_8_  &  (~ i_3_) ) ;
 assign wire9 = ( (~ i_9_)  &  i_4_ ) ;
 assign n_n672 = ( (~ i_3_)  &  i_4_  &  (~ i_2_) ) ;
 assign n_n810 = ( (~ i_9_)  &  i_6_  &  i_4_ ) ;
 assign wire32 = ( (~ i_13_)  &  i_1_ ) ;
 assign wire370 = ( (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire371 = ( (~ i_13_)  &  i_4_  &  i_1_ ) ;
 assign wire295 = ( (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign wire301 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_  &  (~ i_2_) ) ;
 assign wire346 = ( (~ i_9_)  &  (~ i_3_)  &  i_4_  &  (~ i_2_) ) ;
 assign wire11 = ( (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n633 = ( i_5_  &  i_6_  &  i_3_ ) ;
 assign n_n653 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign n_n526 = ( (~ i_12_)  &  (~ i_11_) ) ;
 assign n_n534 = ( i_3_  &  (~ i_1_)  &  i_2_ ) ;
 assign n_n242 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign n_n656 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign n_n194 = ( i_9_  &  i_7_  &  i_11_ ) ;
 assign n_n346 = ( (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign n_n842 = ( (~ i_10_)  &  (~ i_13_) ) ;
 assign wire281 = ( i_4_  &  (~ i_1_) ) ;
 assign n_n791 = ( i_4_  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n755 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n846 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n1258 = ( wire1503 ) | ( wire1504 ) | ( wire6745 ) ;
 assign n_n670 = ( (~ i_3_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire113 = ( wire17  &  wire6669 ) ;
 assign n_n756 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n550 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n732 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire284 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire483 = ( wire1679 ) | ( wire1681 ) | ( n_n748  &  wire484 ) ;
 assign wire482 = ( n_n752  &  n_n575 ) | ( n_n756  &  n_n729 ) ;
 assign wire118 = ( i_13_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire487 = ( i_9_  &  i_13_  &  (~ i_12_) ) | ( i_9_  &  i_13_  &  i_1_ ) ;
 assign wire486 = ( i_9_  &  i_10_  &  i_13_ ) | ( i_10_  &  (~ i_6_)  &  i_13_ ) ;
 assign wire485 = ( i_10_  &  (~ i_6_) ) | ( (~ i_6_)  &  (~ i_1_) ) ;
 assign n_n1126 = ( wire6871 ) | ( wire6872 ) | ( wire6873 ) ;
 assign wire22 = ( (~ i_4_)  &  i_1_ ) ;
 assign wire38 = ( i_9_ ) | ( (~ i_1_) ) ;
 assign wire297 = ( (~ i_4_)  &  (~ i_12_)  &  i_11_ ) ;
 assign n_n1127 = ( wire1293 ) | ( wire1294 ) | ( wire1295 ) | ( wire1296 ) ;
 assign wire493 = ( i_10_  &  (~ i_7_)  &  i_6_ ) | ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire491 = ( n_n748  &  wire342 ) | ( n_n183  &  wire393 ) ;
 assign n_n1112 = ( n_n1126 ) | ( n_n1127 ) | ( wire1283 ) | ( wire6890 ) ;
 assign wire268 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n274 = ( (~ i_13_)  &  (~ i_11_) ) ;
 assign n_n837 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n240 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) ;
 assign wire330 = ( i_4_  &  (~ i_2_) ) ;
 assign n_n771 = ( i_4_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n606 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign n_n813 = ( (~ i_9_)  &  i_5_  &  i_4_ ) ;
 assign wire290 = ( (~ i_6_)  &  i_0_ ) ;
 assign wire308 = ( i_9_  &  i_13_  &  (~ i_12_) ) ;
 assign wire318 = ( (~ i_9_)  &  i_8_  &  i_4_ ) ;
 assign wire494 = ( wire33  &  n_n768 ) | ( n_n769  &  wire6748 ) ;
 assign wire360 = ( i_10_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire497 = ( wire1637 ) | ( n_n665  &  wire1643 ) | ( n_n665  &  wire6640 ) ;
 assign n_n1250 = ( wire1634 ) | ( wire1635 ) | ( (~ i_11_)  &  wire497 ) ;
 assign wire294 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire296 = ( (~ i_4_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire502 = ( wire1669 ) | ( wire6624 ) | ( (~ i_7_)  &  wire503 ) ;
 assign wire501 = ( (~ i_5_)  &  n_n847  &  wire277 ) | ( i_5_  &  n_n852  &  wire277 ) ;
 assign wire272 = ( i_3_  &  (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign wire298 = ( i_3_  &  (~ i_4_)  &  (~ i_1_)  &  i_2_ ) ;
 assign wire311 = ( i_10_  &  (~ i_6_) ) ;
 assign wire363 = ( i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign n_n1129 = ( wire6896 ) | ( i_6_  &  wire1274 ) | ( i_6_  &  wire6893 ) ;
 assign wire104 = ( i_9_  &  i_10_  &  i_12_  &  i_11_ ) ;
 assign wire270 = ( i_9_  &  i_8_  &  i_12_ ) ;
 assign wire379 = ( i_3_  &  i_1_  &  i_11_ ) ;
 assign wire507 = ( i_10_  &  (~ i_8_)  &  i_6_ ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign n_n1123 = ( wire6905 ) | ( (~ i_6_)  &  wire1263 ) | ( (~ i_6_)  &  wire6902 ) ;
 assign n_n623 = ( i_9_  &  i_8_  &  (~ i_11_) ) ;
 assign wire181 = ( (~ i_6_) ) | ( (~ i_12_) ) ;
 assign wire364 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire512 = ( i_3_  &  (~ i_12_)  &  i_2_ ) | ( i_3_  &  i_1_  &  i_2_ ) ;
 assign wire516 = ( (~ i_6_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire513 = ( (~ i_12_)  &  i_2_ ) | ( i_1_  &  i_2_ ) ;
 assign wire300 = ( (~ i_1_)  &  i_0_ ) ;
 assign wire269 = ( (~ i_7_)  &  i_6_ ) ;
 assign n_n822 = ( (~ i_10_)  &  i_12_  &  i_11_ ) ;
 assign n_n840 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n631 = ( (~ i_5_)  &  i_6_  &  i_3_ ) ;
 assign n_n710 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n729 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire519 = ( wire1629 ) | ( wire1630 ) | ( n_n725  &  wire520 ) ;
 assign wire518 = ( n_n837  &  wire277 ) | ( wire22  &  wire6644 ) ;
 assign wire517 = ( n_n843  &  n_n735 ) | ( n_n795  &  wire6642 ) ;
 assign n_n1256 = ( wire1624 ) | ( wire6651 ) | ( n_n732  &  wire519 ) ;
 assign n_n735 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire523 = ( n_n746  &  wire525 ) | ( n_n748  &  wire524 ) ;
 assign wire521 = ( (~ i_13_)  &  wire296 ) | ( n_n346  &  wire6756 ) ;
 assign n_n1231 = ( n_n1258 ) | ( wire1490 ) | ( wire6752 ) | ( wire6759 ) ;
 assign wire350 = ( i_7_  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire529 = ( (~ i_6_)  &  i_0_  &  n_n741 ) | ( i_6_  &  i_0_  &  n_n566 ) ;
 assign wire16 = ( (~ i_5_)  &  i_0_ ) ;
 assign wire533 = ( n_n746  &  n_n575 ) | ( n_n843  &  n_n729 ) ;
 assign wire536 = ( (~ i_8_)  &  (~ i_3_) ) | ( (~ i_7_)  &  (~ i_2_) ) ;
 assign wire277 = ( (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n597 = ( i_10_  &  i_7_  &  (~ i_8_) ) ;
 assign n_n651 = ( i_10_  &  i_7_  &  i_8_ ) ;
 assign n_n1255 = ( wire1609 ) | ( wire1610 ) | ( wire6658 ) ;
 assign wire405 = ( (~ i_13_)  &  i_11_  &  n_n835  &  n_n710 ) ;
 assign wire545 = ( wire1603 ) | ( wire1605 ) | ( wire381  &  wire546 ) ;
 assign wire544 = ( n_n833  &  n_n712 ) | ( n_n830  &  n_n710 ) ;
 assign wire543 = ( n_n847  &  n_n712 ) | ( n_n852  &  n_n710 ) ;
 assign n_n1253 = ( wire6683 ) | ( n_n849  &  wire571 ) ;
 assign wire120 = ( n_n853  &  n_n699  &  n_n678 ) ;
 assign n_n1229 = ( n_n1253 ) | ( wire1584 ) | ( wire6678 ) | ( wire6694 ) ;
 assign wire553 = ( n_n35  &  wire393 ) | ( n_n756  &  wire6922 ) ;
 assign wire552 = ( n_n638  &  (~ wire181) ) | ( n_n619  &  wire6921 ) ;
 assign n_n1128 = ( wire1221 ) | ( wire6926 ) | ( (~ i_4_)  &  wire553 ) ;
 assign wire30 = ( (~ i_7_)  &  (~ i_5_) ) ;
 assign wire352 = ( (~ i_7_)  &  i_2_ ) ;
 assign wire557 = ( n_n844  &  wire30 ) | ( wire7249  &  wire7250 ) ;
 assign wire338 = ( i_10_  &  (~ i_5_)  &  i_12_  &  i_0_ ) ;
 assign wire560 = ( n_n840  &  wire562 ) | ( wire333  &  wire561 ) ;
 assign wire558 = ( i_10_  &  i_1_  &  (~ i_11_) ) | ( i_10_  &  i_1_  &  i_0_ ) ;
 assign n_n1000 = ( wire176 ) | ( wire7255 ) | ( (~ i_12_)  &  wire560 ) ;
 assign wire565 = ( wire375 ) | ( wire170 ) | ( wire171 ) | ( wire172 ) ;
 assign wire564 = ( n_n432  &  wire36 ) | ( wire26  &  wire7257 ) ;
 assign n_n503 = ( (~ i_9_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire73 = ( (~ i_10_)  &  (~ i_7_)  &  wire17  &  n_n683 ) ;
 assign wire121 = ( (~ i_13_)  &  i_12_  &  n_n835  &  n_n712 ) ;
 assign wire571 = ( n_n712  &  wire573 ) | ( n_n710  &  wire572 ) ;
 assign n_n1233 = ( n_n1264 ) | ( n_n1265 ) | ( wire6782 ) ;
 assign wire574 = ( n_n826  &  wire9 ) | ( (~ wire38)  &  n_n851 ) ;
 assign n_n624 = ( i_5_  &  i_6_  &  (~ i_2_) ) ;
 assign wire20 = ( i_5_  &  i_0_ ) ;
 assign wire579 = ( wire24 ) | ( wire931 ) | ( wire932 ) ;
 assign wire578 = ( n_n752  &  wire24 ) | ( n_n819  &  wire6848 ) ;
 assign n_n619 = ( i_9_  &  i_10_  &  i_8_ ) ;
 assign wire583 = ( wire1418 ) | ( wire1419 ) | ( n_n843  &  wire584 ) ;
 assign wire581 = ( wire1414 ) | ( n_n832  &  wire410 ) | ( n_n832  &  wire1416 ) ;
 assign n_n1234 = ( wire115 ) | ( wire1400 ) | ( wire1402 ) | ( wire6814 ) ;
 assign wire591 = ( i_9_  &  i_7_  &  i_6_ ) | ( i_7_  &  (~ i_5_)  &  i_6_ ) ;
 assign n_n851 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire594 = ( i_9_  &  i_7_ ) | ( i_7_  &  (~ i_2_) ) ;
 assign wire593 = ( i_9_  &  i_10_ ) | ( i_10_  &  (~ i_7_) ) ;
 assign wire123 = ( (~ i_7_)  &  (~ i_6_)  &  i_3_  &  i_0_ ) ;
 assign wire276 = ( i_5_  &  (~ i_12_) ) ;
 assign wire291 = ( i_3_  &  i_0_ ) ;
 assign wire354 = ( (~ i_7_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire596 = ( n_n818  &  wire7287 ) | ( n_n415  &  wire7288 ) ;
 assign n_n277 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire115 = ( i_1_  &  i_2_  &  i_0_  &  wire6807 ) ;
 assign wire410 = ( (~ i_13_)  &  (~ i_12_)  &  n_n835  &  n_n541 ) ;
 assign wire604 = ( wire1214 ) | ( wire1215 ) | ( wire1216 ) | ( wire1217 ) ;
 assign wire606 = ( wire15  &  n_n827 ) | ( n_n819  &  wire291 ) ;
 assign n_n1264 = ( wire1462 ) | ( wire1463 ) | ( wire1466 ) | ( wire6766 ) ;
 assign n_n1265 = ( wire6773 ) | ( n_n849  &  wire1453 ) | ( n_n849  &  wire1454 ) ;
 assign wire292 = ( i_3_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire340 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire359 = ( (~ i_5_)  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire402 = ( (~ i_9_)  &  (~ i_13_)  &  n_n846  &  n_n822 ) ;
 assign wire612 = ( n_n818  &  n_n810 ) | ( n_n633  &  wire6777 ) ;
 assign n_n1191 = ( wire1132 ) | ( wire1134 ) | ( wire6978 ) | ( wire6979 ) ;
 assign n_n1185 = ( wire1154 ) | ( i_2_  &  wire6965 ) | ( i_2_  &  wire6966 ) ;
 assign wire351 = ( (~ i_9_)  &  i_7_  &  i_4_ ) ;
 assign wire369 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire617 = ( n_n816  &  wire9 ) | ( wire19  &  wire294 ) ;
 assign wire616 = ( n_n761  &  wire351 ) | ( (~ i_11_)  &  n_n761  &  n_n275 ) ;
 assign wire314 = ( i_9_  &  i_10_  &  i_7_ ) ;
 assign wire365 = ( i_3_  &  (~ i_12_) ) ;
 assign wire619 = ( n_n35  &  n_n656 ) | ( wire275  &  wire356 ) ;
 assign n_n612 = ( i_5_  &  i_1_  &  i_2_ ) ;
 assign wire275 = ( (~ i_7_)  &  (~ i_2_) ) ;
 assign wire626 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) | ( i_10_  &  (~ i_7_)  &  i_2_ ) ;
 assign wire628 = ( (~ i_8_)  &  wire37 ) | ( (~ i_8_)  &  (~ i_3_)  &  n_n716 ) ;
 assign n_n768 = ( (~ i_9_)  &  i_8_  &  i_5_ ) ;
 assign wire632 = ( n_n566  &  wire19 ) | ( n_n741  &  wire633 ) ;
 assign wire639 = ( wire7129 ) | ( i_5_  &  wire879 ) | ( i_5_  &  wire7128 ) ;
 assign wire638 = ( n_n545  &  wire377 ) | ( n_n755  &  wire7127 ) ;
 assign wire637 = ( n_n185  &  n_n683 ) | ( n_n752  &  wire7126 ) ;
 assign wire41 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_0_) ) | ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire382 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire641 = ( (~ i_6_)  &  (~ i_0_)  &  n_n242 ) | ( i_6_  &  (~ i_0_)  &  n_n277 ) ;
 assign wire324 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign n_n910 = ( wire1064 ) | ( wire7019 ) | ( wire382  &  wire324 ) ;
 assign wire648 = ( wire1848 ) | ( wire1849 ) | ( wire33  &  wire649 ) ;
 assign wire299 = ( i_12_  &  i_2_ ) ;
 assign wire316 = ( i_10_  &  (~ i_7_)  &  i_12_ ) ;
 assign wire376 = ( i_7_  &  i_5_  &  i_1_ ) ;
 assign wire395 = ( i_9_  &  i_5_  &  i_6_  &  i_12_ ) ;
 assign wire36 = ( i_6_  &  i_0_ ) ;
 assign wire304 = ( i_10_  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire384 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  i_2_ ) ;
 assign wire385 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) ;
 assign wire347 = ( i_10_  &  (~ i_5_) ) ;
 assign wire356 = ( i_8_  &  i_12_  &  (~ i_11_) ) ;
 assign wire655 = ( wire777 ) | ( wire7185 ) | ( i_8_  &  wire657 ) ;
 assign n_n991 = ( wire772 ) | ( wire773 ) | ( (~ i_4_)  &  wire655 ) ;
 assign wire660 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign n_n879 = ( wire1814 ) | ( wire6506 ) | ( wire6507 ) ;
 assign wire287 = ( i_7_  &  i_3_  &  i_1_  &  i_0_ ) ;
 assign wire388 = ( (~ i_7_)  &  (~ i_6_)  &  i_0_ ) ;
 assign n_n881 = ( wire1805 ) | ( wire1806 ) | ( wire1808 ) | ( wire6512 ) ;
 assign wire668 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire667 = ( n_n779  &  wire288 ) | ( n_n685  &  wire30 ) ;
 assign wire666 = ( n_n699  &  n_n710 ) | ( n_n792  &  wire7066 ) ;
 assign wire669 = ( wire1074 ) | ( n_n658  &  n_n275 ) | ( n_n275  &  wire7013 ) ;
 assign wire671 = ( wire35  &  n_n675 ) | ( n_n672  &  wire11 ) ;
 assign wire406 = ( i_4_  &  (~ i_1_)  &  (~ i_2_)  &  n_n768 ) ;
 assign wire676 = ( wire279  &  n_n671 ) | ( n_n792  &  wire677 ) ;
 assign wire403 = ( (~ i_9_)  &  i_7_  &  i_5_  &  n_n685 ) ;
 assign wire334 = ( i_9_  &  i_12_  &  i_11_ ) ;
 assign wire380 = ( (~ i_11_)  &  (~ i_0_) ) ;
 assign wire686 = ( n_n432  &  n_n176 ) | ( wire12  &  wire270 ) ;
 assign wire685 = ( i_5_  &  wire292 ) | ( i_5_  &  (~ i_12_)  &  n_n814 ) ;
 assign n_n993 = ( wire373 ) | ( wire7191 ) | ( wire18  &  wire685 ) ;
 assign n_n913 = ( wire1011 ) | ( wire1012 ) | ( wire7046 ) | ( wire7047 ) ;
 assign wire696 = ( wire1003 ) | ( wire1005 ) | ( wire7050 ) | ( wire7051 ) ;
 assign n_n906 = ( n_n913 ) | ( wire7054 ) | ( (~ i_12_)  &  wire696 ) ;
 assign wire397 = ( i_9_  &  i_5_  &  (~ i_6_)  &  i_11_ ) ;
 assign wire701 = ( i_9_  &  i_7_  &  i_6_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire700 = ( n_n432  &  n_n826 ) | ( wire380  &  wire7269 ) ;
 assign wire321 = ( i_5_  &  (~ i_0_) ) ;
 assign wire704 = ( i_5_  &  (~ i_6_)  &  i_3_ ) | ( i_5_  &  i_3_  &  i_1_ ) ;
 assign wire703 = ( n_n746  &  wire366 ) | ( n_n826  &  wire7275 ) ;
 assign wire706 = ( i_10_  &  (~ i_5_) ) | ( (~ i_5_)  &  (~ i_0_) ) ;
 assign wire705 = ( wire7294  &  wire7295 ) | ( wire707  &  wire7296 ) ;
 assign wire708 = ( n_n538  &  wire333 ) | ( n_n369  &  wire7178 ) ;
 assign n_n987 = ( wire784 ) | ( wire785 ) | ( wire354  &  wire708 ) ;
 assign wire366 = ( i_5_  &  i_3_  &  i_0_ ) ;
 assign wire717 = ( wire20  &  wire334 ) | ( n_n415  &  wire718 ) ;
 assign wire716 = ( n_n176  &  wire719 ) | ( wire270  &  wire7194 ) ;
 assign n_n965 = ( n_n991 ) | ( n_n993 ) | ( wire256 ) | ( wire7196 ) ;
 assign n_n981 = ( wire857 ) | ( wire7140 ) | ( i_5_  &  wire762 ) ;
 assign n_n984 = ( wire836 ) | ( wire837 ) | ( wire7155 ) ;
 assign n_n983 = ( wire73 ) | ( wire824 ) | ( wire825 ) | ( wire7161 ) ;
 assign wire725 = ( n_n773  &  n_n671 ) | ( n_n835  &  wire726 ) ;
 assign wire724 = ( wire37 ) | ( (~ i_3_)  &  n_n725 ) ;
 assign wire723 = ( wire37  &  n_n671 ) | ( n_n771  &  wire7165 ) ;
 assign wire374 = ( i_9_  &  (~ i_4_)  &  i_11_ ) ;
 assign n_n986 = ( wire246 ) | ( wire247 ) | ( wire249 ) | ( wire7205 ) ;
 assign wire24 = ( (~ i_9_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire735 = ( wire24 ) | ( wire808 ) | ( wire809 ) ;
 assign wire737 = ( wire395 ) | ( wire397 ) | ( i_6_  &  wire10 ) ;
 assign wire736 = ( wire230 ) | ( wire231 ) | ( wire263  &  wire7219 ) ;
 assign wire342 = ( i_9_  &  (~ i_12_)  &  i_11_ ) ;
 assign wire738 = ( n_n818  &  wire304 ) | ( n_n752  &  wire7226 ) ;
 assign wire744 = ( n_n581  &  wire290 ) | ( i_2_  &  wire288  &  wire290 ) ;
 assign wire747 = ( i_13_  &  (~ i_12_)  &  (~ i_11_) ) | ( (~ i_13_)  &  i_4_  &  i_12_  &  i_11_ ) ;
 assign wire746 = ( i_13_  &  (~ i_12_) ) | ( (~ i_13_)  &  i_4_  &  i_12_ ) ;
 assign wire751 = ( (~ i_5_)  &  i_6_  &  i_3_ ) | ( (~ i_5_)  &  i_3_  &  i_1_ ) ;
 assign wire752 = ( wire80 ) | ( wire81 ) | ( n_n840  &  wire54 ) ;
 assign wire263 = ( i_6_  &  (~ i_0_) ) ;
 assign wire762 = ( wire863 ) | ( wire864 ) | ( n_n716  &  wire763 ) ;
 assign wire761 = ( n_n678  &  wire7132 ) | ( n_n716  &  wire7133 ) ;
 assign wire54 = ( (~ i_5_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire10 = ( i_9_  &  i_10_  &  i_12_ ) | ( i_10_  &  (~ i_5_)  &  i_12_ ) ;
 assign wire42 = ( (~ i_5_)  &  i_1_  &  i_2_ ) | ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire51 = ( n_n769  &  n_n771 ) | ( n_n835  &  wire318 ) ;
 assign wire317 = ( i_8_  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire319 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  i_4_ ) ;
 assign wire329 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire335 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire375 = ( i_5_  &  i_6_  &  (~ i_12_) ) ;
 assign wire393 = ( i_10_  &  i_7_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire424 = ( n_n850  &  n_n751 ) | ( n_n570  &  n_n503 ) ;
 assign wire423 = ( wire329  &  wire6549 ) | ( n_n729  &  wire6550 ) ;
 assign wire427 = ( n_n623  &  wire429 ) | ( n_n619  &  wire428 ) ;
 assign wire426 = ( i_5_  &  i_1_  &  i_2_ ) | ( i_1_  &  i_2_  &  i_0_ ) ;
 assign wire429 = ( i_6_  &  (~ i_0_) ) | ( (~ i_1_)  &  (~ i_0_) ) ;
 assign wire428 = ( i_6_  &  i_0_ ) | ( i_1_  &  i_0_ ) ;
 assign wire436 = ( n_n835 ) | ( n_n624 ) | ( wire1740 ) | ( wire1741 ) ;
 assign wire440 = ( (~ i_9_)  &  i_7_  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire439 = ( (~ i_9_)  &  i_7_ ) | ( (~ i_10_)  &  (~ i_7_) ) ;
 assign wire447 = ( i_1_  &  wire335 ) | ( (~ i_13_)  &  i_1_  &  n_n277 ) ;
 assign wire451 = ( n_n816  &  wire264 ) | ( n_n822  &  wire452 ) ;
 assign wire452 = ( i_5_  &  (~ i_6_)  &  (~ i_13_) ) | ( i_5_  &  (~ i_13_)  &  i_1_ ) ;
 assign wire459 = ( wire279  &  wire301 ) | ( n_n852  &  wire329 ) ;
 assign wire469 = ( n_n658  &  n_n844 ) | ( n_n847  &  n_n653 ) ;
 assign wire468 = ( i_5_  &  (~ i_6_)  &  n_n838 ) | ( (~ i_5_)  &  i_6_  &  n_n830 ) ;
 assign wire479 = ( n_n852  &  n_n846 ) | ( n_n847  &  n_n851 ) ;
 assign wire484 = ( i_5_  &  n_n833  &  wire277 ) | ( (~ i_5_)  &  n_n830  &  wire277 ) ;
 assign wire503 = ( wire22  &  wire6622 ) | ( n_n735  &  wire6623 ) ;
 assign wire515 = ( i_6_  &  (~ i_12_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire520 = ( i_6_  &  n_n847  &  wire27 ) | ( (~ i_6_)  &  wire27  &  n_n840 ) ;
 assign wire525 = ( i_0_  &  wire265  &  n_n846 ) | ( (~ i_0_)  &  wire265  &  n_n851 ) ;
 assign wire524 = ( n_n833  &  n_n846 ) | ( n_n830  &  n_n851 ) ;
 assign wire530 = ( wire23  &  n_n729 ) | ( n_n575  &  wire531 ) ;
 assign wire531 = ( i_7_ ) | ( i_8_  &  (~ i_3_) ) ;
 assign wire541 = ( (~ i_5_)  &  n_n833  &  wire277 ) | ( i_5_  &  n_n830  &  wire277 ) ;
 assign wire546 = ( i_5_  &  n_n819  &  wire277 ) | ( (~ i_5_)  &  n_n699  &  wire277 ) ;
 assign wire551 = ( (~ i_5_)  &  i_6_  &  n_n838 ) | ( i_5_  &  (~ i_6_)  &  n_n830 ) ;
 assign wire562 = ( i_10_  &  (~ i_7_)  &  i_5_ ) | ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire561 = ( i_10_  &  i_5_  &  (~ i_6_) ) | ( i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire569 = ( n_n795  &  n_n570 ) | ( n_n843  &  n_n751 ) ;
 assign wire573 = ( n_n830  &  n_n756 ) | ( n_n746  &  n_n840 ) ;
 assign wire572 = ( n_n838  &  n_n752 ) | ( n_n833  &  n_n756 ) ;
 assign wire576 = ( i_5_  &  (~ i_6_)  &  i_2_ ) | ( i_5_  &  i_1_  &  i_2_ ) ;
 assign wire584 = ( i_0_  &  wire33  &  n_n541 ) | ( (~ i_0_)  &  wire33  &  wire6803 ) ;
 assign wire615 = ( i_10_  &  i_7_  &  (~ i_8_) ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire622 = ( i_2_ ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire633 = ( (~ i_8_)  &  (~ i_3_) ) | ( (~ i_7_)  &  (~ i_2_) ) ;
 assign wire636 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) | ( (~ i_10_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire635 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire644 = ( (~ i_9_)  &  (~ i_8_)  &  i_6_ ) | ( (~ i_10_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire643 = ( (~ i_7_) ) | ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire646 = ( i_6_  &  (~ i_3_)  &  (~ i_0_) ) | ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire649 = ( (~ i_8_)  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire653 = ( i_8_  &  i_12_ ) | ( i_10_  &  (~ i_7_)  &  i_12_ ) ;
 assign wire657 = ( i_0_  &  wire33  &  wire10 ) | ( (~ i_0_)  &  wire33  &  wire7184 ) ;
 assign wire673 = ( i_8_  &  (~ i_3_) ) | ( i_7_  &  (~ i_2_) ) ;
 assign wire677 = ( (~ i_5_)  &  (~ i_6_) ) | ( (~ i_6_)  &  (~ i_0_) ) ;
 assign wire680 = ( (~ i_9_)  &  i_7_  &  i_8_ ) | ( (~ i_10_)  &  (~ i_7_)  &  i_8_ ) ;
 assign wire683 = ( n_n814 ) | ( wire1794 ) | ( i_1_  &  wire684 ) ;
 assign wire684 = ( i_9_  &  i_7_  &  i_8_ ) | ( i_9_  &  i_7_  &  i_6_ ) ;
 assign wire689 = ( (~ i_5_)  &  i_0_  &  n_n432 ) | ( (~ i_5_)  &  (~ i_0_)  &  wire7190 ) ;
 assign wire698 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire707 = ( (~ i_5_)  &  i_0_ ) | ( i_5_  &  (~ i_12_)  &  (~ i_0_) ) ;
 assign wire712 = ( n_n541  &  wire333 ) | ( n_n369  &  wire347 ) ;
 assign wire719 = ( i_10_  &  i_12_  &  (~ i_11_) ) | ( i_10_  &  i_12_  &  i_0_ ) | ( i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire718 = ( i_9_  &  i_0_ ) | ( (~ i_5_)  &  i_0_ ) ;
 assign wire726 = ( (~ i_7_) ) | ( (~ i_8_)  &  (~ i_3_) ) ;
 assign wire728 = ( (~ i_9_)  &  i_4_ ) | ( (~ i_8_)  &  i_4_ ) ;
 assign wire734 = ( n_n819  &  wire381 ) | ( n_n752  &  n_n550 ) ;
 assign wire741 = ( i_9_  &  i_7_  &  i_8_ ) | ( i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign wire763 = ( n_n683  &  n_n792 ) | ( n_n699  &  wire7136 ) ;
 assign wire40 = ( (~ i_10_)  &  (~ i_13_)  &  n_n838  &  wire7322 ) ;
 assign wire50 = ( n_n687  &  wire57 ) | ( n_n687  &  n_n729  &  wire7325 ) ;
 assign wire52 = ( wire16  &  wire59 ) | ( wire16  &  wire60 ) | ( wire16  &  wire7327 ) ;
 assign wire57 = ( (~ i_7_)  &  (~ i_5_)  &  wire1202 ) | ( (~ i_7_)  &  (~ i_5_)  &  wire1203 ) ;
 assign wire59 = ( n_n699  &  wire62 ) | ( n_n699  &  wire63 ) ;
 assign wire60 = ( (~ i_1_)  &  wire329 ) ;
 assign wire62 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire63 = ( (~ i_13_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire64 = ( wire82  &  wire7312 ) | ( wire83  &  wire7312 ) ;
 assign wire65 = ( wire338  &  wire7313 ) | ( wire84  &  wire7313 ) ;
 assign wire80 = ( i_5_  &  (~ i_12_)  &  i_1_  &  i_2_ ) ;
 assign wire81 = ( i_5_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire82 = ( i_7_  &  i_12_  &  i_2_ ) ;
 assign wire83 = ( i_8_  &  i_3_  &  i_12_ ) ;
 assign wire84 = ( (~ i_5_)  &  i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire86 = ( i_12_  &  (~ i_11_)  &  n_n597  &  wire751 ) ;
 assign wire89 = ( wire126  &  wire95 ) | ( wire126  &  n_n526  &  n_n840 ) ;
 assign wire95 = ( (~ i_5_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire97 = ( (~ i_12_)  &  i_2_  &  n_n639  &  wire7304 ) ;
 assign wire98 = ( i_3_  &  i_2_  &  i_0_  &  wire304 ) ;
 assign wire103 = ( i_9_  &  i_10_  &  i_13_  &  i_0_ ) ;
 assign wire107 = ( i_10_  &  (~ i_5_)  &  i_13_  &  i_0_ ) ;
 assign wire112 = ( i_9_  &  i_5_  &  i_13_  &  (~ i_12_) ) ;
 assign wire127 = ( i_5_  &  (~ i_12_)  &  n_n840  &  wire7280 ) ;
 assign wire128 = ( i_10_  &  i_11_  &  n_n826  &  wire7282 ) ;
 assign wire129 = ( n_n316  &  n_n631  &  wire314 ) | ( n_n316  &  n_n631  &  wire136 ) ;
 assign wire130 = ( i_9_  &  i_10_  &  n_n639  &  wire354 ) ;
 assign wire136 = ( i_10_  &  (~ i_8_)  &  i_2_ ) ;
 assign wire139 = ( n_n194  &  wire144 ) | ( n_n194  &  wire145 ) ;
 assign wire141 = ( i_9_  &  i_5_  &  i_13_  &  i_0_ ) ;
 assign wire142 = ( i_5_  &  i_13_  &  (~ i_12_)  &  (~ i_0_) ) ;
 assign wire143 = ( i_13_  &  (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire144 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire145 = ( i_5_  &  (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire150 = ( (~ i_12_)  &  i_11_  &  n_n639  &  wire7264 ) ;
 assign wire154 = ( wire270  &  wire156 ) | ( n_n826  &  wire34  &  wire270 ) ;
 assign wire156 = ( i_5_  &  i_3_  &  i_11_  &  i_0_ ) ;
 assign wire163 = ( i_9_  &  i_10_  &  i_1_  &  i_0_ ) ;
 assign wire166 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire170 = ( (~ i_5_)  &  i_6_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire171 = ( i_6_  &  (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire172 = ( i_5_  &  i_6_  &  i_0_ ) ;
 assign wire176 = ( n_n656  &  wire180 ) | ( n_n656  &  wire182 ) ;
 assign wire180 = ( (~ i_5_)  &  i_6_  &  i_12_  &  i_2_ ) ;
 assign wire182 = ( (~ i_5_)  &  i_1_  &  i_2_ ) ;
 assign wire190 = ( i_3_  &  i_0_  &  wire104 ) | ( i_2_  &  i_0_  &  wire104 ) ;
 assign wire192 = ( i_1_  &  wire194 ) | ( i_1_  &  wire1408 ) | ( i_1_  &  wire1409 ) ;
 assign wire194 = ( i_9_  &  i_10_  &  i_5_  &  (~ i_12_) ) ;
 assign wire198 = ( i_9_  &  wire7234  &  wire7235 ) | ( (~ i_0_)  &  wire7234  &  wire7235 ) ;
 assign wire200 = ( (~ i_8_)  &  i_5_  &  n_n598  &  wire374 ) ;
 assign wire201 = ( (~ i_4_)  &  i_1_  &  wire206 ) | ( (~ i_4_)  &  i_1_  &  wire207 ) ;
 assign wire206 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  wire7239 ) ;
 assign wire207 = ( wire27  &  wire208 ) | ( wire27  &  wire841 ) | ( wire27  &  wire842 ) ;
 assign wire208 = ( i_9_  &  i_5_  &  i_11_  &  i_0_ ) ;
 assign wire212 = ( (~ i_6_)  &  (~ i_0_)  &  n_n538  &  wire7223 ) ;
 assign wire213 = ( i_5_  &  (~ i_6_)  &  n_n412  &  wire342 ) ;
 assign wire215 = ( (~ i_4_)  &  i_1_  &  wire222 ) | ( (~ i_4_)  &  i_1_  &  wire7229 ) ;
 assign wire222 = ( i_12_  &  (~ i_11_)  &  wire223 ) | ( i_12_  &  (~ i_11_)  &  wire224 ) ;
 assign wire223 = ( i_10_  &  i_7_  &  i_8_  &  (~ i_5_) ) ;
 assign wire224 = ( i_7_  &  i_8_  &  (~ i_5_)  &  (~ i_0_) ) ;
 assign wire225 = ( (~ i_5_)  &  i_6_  &  n_n412  &  wire7215 ) ;
 assign wire230 = ( i_1_  &  (~ i_11_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire231 = ( i_10_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire235 = ( i_7_  &  i_6_  &  n_n541  &  wire7208 ) ;
 assign wire236 = ( i_10_  &  i_12_  &  n_n153  &  wire591 ) ;
 assign wire237 = ( wire360  &  wire272 ) | ( wire272  &  wire241 ) ;
 assign wire238 = ( i_1_  &  i_2_  &  i_0_  &  wire307 ) ;
 assign wire241 = ( i_9_  &  i_5_  &  (~ i_12_) ) ;
 assign wire245 = ( wire307  &  wire7199 ) | ( wire253  &  wire7199 ) ;
 assign wire246 = ( wire304  &  wire7200 ) | ( wire397  &  wire7200 ) ;
 assign wire247 = ( (~ i_7_)  &  i_5_  &  n_n826  &  wire374 ) ;
 assign wire249 = ( (~ i_8_)  &  i_5_  &  wire252 ) | ( (~ i_8_)  &  i_5_  &  wire7203 ) ;
 assign wire252 = ( i_9_  &  i_11_  &  wire296 ) ;
 assign wire253 = ( i_5_  &  i_3_  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire255 = ( i_9_  &  i_12_  &  n_n752  &  wire366 ) ;
 assign wire256 = ( (~ i_4_)  &  i_2_  &  wire716 ) ;
 assign wire258 = ( i_6_  &  i_0_  &  n_n432  &  wire6976 ) ;
 assign wire362 = ( (~ i_11_)  &  (~ i_0_)  &  n_n176  &  wire7188 ) ;
 assign wire373 = ( i_3_  &  wire411 ) | ( i_3_  &  n_n752  &  wire689 ) ;
 assign wire411 = ( n_n840  &  wire768 ) | ( n_n840  &  wire769 ) ;
 assign wire768 = ( i_9_  &  i_8_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire769 = ( i_9_  &  i_8_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire772 = ( i_10_  &  (~ i_5_)  &  n_n346  &  wire356 ) ;
 assign wire773 = ( wire296  &  wire7181 ) ;
 assign wire777 = ( n_n752  &  wire338 ) | ( n_n752  &  wire779 ) ;
 assign wire779 = ( i_9_  &  i_5_  &  i_12_  &  i_0_ ) ;
 assign wire784 = ( (~ i_4_)  &  wire788 ) | ( (~ i_4_)  &  wire287  &  wire10 ) ;
 assign wire785 = ( i_7_  &  wire795 ) | ( i_7_  &  n_n316  &  wire712 ) ;
 assign wire788 = ( n_n826  &  wire790 ) | ( n_n826  &  wire791 ) ;
 assign wire790 = ( i_9_  &  i_7_  &  i_5_  &  i_12_ ) ;
 assign wire791 = ( i_10_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire795 = ( i_3_  &  (~ i_4_)  &  i_0_  &  wire395 ) ;
 assign wire798 = ( i_7_  &  i_0_  &  n_n658  &  wire24 ) ;
 assign wire800 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_)  &  wire7175 ) ;
 assign wire801 = ( wire20  &  wire802 ) | ( (~ i_3_)  &  wire20  &  wire734 ) ;
 assign wire802 = ( (~ i_1_)  &  wire335 ) | ( (~ i_1_)  &  wire286  &  wire24 ) ;
 assign wire808 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire809 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire814 = ( n_n853  &  n_n819  &  n_n678 ) ;
 assign wire824 = ( n_n853  &  wire7157 ) | ( n_n764  &  n_n853  &  n_n791 ) ;
 assign wire825 = ( (~ i_10_)  &  (~ i_6_)  &  wire17  &  n_n671 ) ;
 assign wire834 = ( i_5_  &  (~ i_6_)  &  n_n581  &  wire297 ) ;
 assign wire835 = ( i_6_  &  (~ i_0_)  &  n_n764  &  wire17 ) ;
 assign wire836 = ( n_n853  &  wire51 ) | ( n_n853  &  n_n671  &  n_n810 ) ;
 assign wire837 = ( n_n843  &  wire840 ) | ( n_n843  &  wire20  &  wire374 ) ;
 assign wire840 = ( (~ i_4_)  &  wire841 ) | ( (~ i_4_)  &  wire842 ) ;
 assign wire841 = ( i_5_  &  (~ i_12_)  &  i_11_  &  (~ i_0_) ) ;
 assign wire842 = ( i_10_  &  (~ i_5_)  &  i_11_  &  i_0_ ) ;
 assign wire843 = ( (~ i_5_)  &  (~ i_0_)  &  n_n819  &  wire301 ) ;
 assign wire844 = ( n_n671  &  n_n176  &  wire284 ) ;
 assign wire845 = ( n_n755  &  wire850 ) | ( n_n755  &  wire852 ) | ( n_n755  &  wire7146 ) ;
 assign wire846 = ( i_7_  &  n_n545  &  wire7138 ) ;
 assign wire850 = ( wire35  &  wire853 ) | ( wire35  &  wire854 ) | ( wire35  &  wire855 ) ;
 assign wire852 = ( i_7_  &  i_8_  &  (~ i_5_)  &  n_n791 ) ;
 assign wire853 = ( i_8_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire854 = ( i_7_  &  i_8_  &  i_6_  &  (~ i_0_) ) ;
 assign wire855 = ( i_7_  &  (~ i_3_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire856 = ( (~ i_7_)  &  i_5_  &  wire37  &  n_n683 ) ;
 assign wire857 = ( i_5_  &  (~ i_6_)  &  wire761 ) ;
 assign wire859 = ( i_8_  &  (~ i_3_)  &  n_n545  &  wire7138 ) ;
 assign wire863 = ( wire37  &  wire7134 ) ;
 assign wire864 = ( (~ i_7_)  &  (~ i_8_)  &  n_n849  &  n_n791 ) ;
 assign wire879 = ( i_8_  &  (~ i_3_)  &  n_n550 ) ;
 assign wire881 = ( n_n719  &  n_n837  &  wire7119 ) ;
 assign wire882 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  wire7121 ) ;
 assign wire883 = ( n_n716  &  wire885 ) | ( n_n716  &  n_n675  &  wire7015 ) ;
 assign wire884 = ( n_n761  &  wire406 ) | ( n_n761  &  wire887 ) | ( n_n761  &  wire7122 ) ;
 assign wire885 = ( i_5_  &  (~ i_3_)  &  (~ i_2_)  &  n_n503 ) ;
 assign wire887 = ( i_5_  &  i_6_  &  wire346 ) | ( i_5_  &  i_6_  &  wire891 ) ;
 assign wire891 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_4_ ) ;
 assign wire895 = ( (~ i_5_)  &  wire901 ) | ( (~ i_5_)  &  n_n816  &  wire9 ) ;
 assign wire896 = ( (~ i_10_)  &  wire903 ) | ( (~ i_10_)  &  wire301  &  wire317 ) ;
 assign wire901 = ( (~ i_9_)  &  (~ i_10_)  &  wire673  &  wire6594 ) ;
 assign wire903 = ( n_n545  &  wire350 ) | ( n_n545  &  wire905 ) ;
 assign wire905 = ( i_7_  &  (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire907 = ( (~ i_10_)  &  (~ i_5_)  &  n_n675  &  wire7109 ) ;
 assign wire909 = ( n_n761  &  wire912 ) | ( n_n761  &  wire7110 ) | ( n_n761  &  wire7111 ) ;
 assign wire912 = ( i_4_  &  (~ i_2_)  &  wire322 ) ;
 assign wire917 = ( n_n545  &  n_n240  &  wire668 ) ;
 assign wire925 = ( (~ i_7_)  &  i_5_  &  n_n838  &  wire7094 ) ;
 assign wire927 = ( wire319  &  wire7100 ) | ( wire335  &  wire7100 ) | ( wire934  &  wire7100 ) ;
 assign wire931 = ( (~ i_9_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire932 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire934 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire937 = ( i_5_  &  n_n741  &  n_n761  &  wire536 ) ;
 assign wire939 = ( (~ i_13_)  &  wire7091 ) | ( (~ i_13_)  &  n_n741  &  wire275 ) ;
 assign wire947 = ( wire954  &  wire7085 ) | ( wire7084  &  wire7085 ) ;
 assign wire948 = ( (~ i_5_)  &  (~ i_6_)  &  n_n670  &  wire7086 ) ;
 assign wire949 = ( n_n575  &  wire951 ) | ( n_n575  &  n_n606  &  wire7087 ) ;
 assign wire951 = ( i_8_  &  (~ i_5_)  &  (~ i_6_)  &  n_n670 ) ;
 assign wire954 = ( i_0_  &  wire957 ) | ( i_0_  &  wire958 ) ;
 assign wire957 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_2_) ) ;
 assign wire958 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire960 = ( wire350  &  wire7078 ) ;
 assign wire961 = ( n_n838  &  wire7080 ) | ( (~ i_5_)  &  n_n838  &  wire530 ) ;
 assign wire962 = ( (~ i_9_)  &  (~ i_13_)  &  n_n701  &  wire300 ) ;
 assign wire970 = ( (~ i_10_)  &  (~ i_5_)  &  n_n675  &  wire7067 ) ;
 assign wire971 = ( (~ i_9_)  &  i_7_  &  i_8_  &  wire7068 ) ;
 assign wire972 = ( (~ i_9_)  &  wire979 ) | ( (~ i_9_)  &  n_n526  &  n_n624 ) ;
 assign wire979 = ( (~ i_1_)  &  n_n701 ) | ( (~ i_1_)  &  wire375 ) | ( (~ i_1_)  &  wire981 ) ;
 assign wire981 = ( i_5_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire987 = ( n_n653  &  wire382 ) | ( n_n653  &  wire995 ) ;
 assign wire988 = ( (~ i_5_)  &  (~ i_11_)  &  (~ i_0_) ) | ( (~ i_12_)  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire993 = ( (~ i_9_)  &  (~ i_3_) ) | ( (~ i_9_)  &  (~ i_2_) ) ;
 assign wire995 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1003 = ( i_6_  &  (~ i_1_)  &  (~ i_0_) ) | ( i_6_  &  (~ i_0_)  &  wire1009 ) ;
 assign wire1005 = ( (~ i_10_)  &  i_8_  &  (~ i_6_)  &  n_n671 ) ;
 assign wire1009 = ( (~ i_9_)  &  i_7_  &  i_8_  &  (~ i_3_) ) ;
 assign wire1011 = ( (~ i_11_)  &  wire1017 ) | ( (~ i_11_)  &  n_n658  &  n_n275 ) ;
 assign wire1012 = ( (~ i_12_)  &  wire1019 ) | ( (~ i_12_)  &  wire265  &  n_n827 ) ;
 assign wire1017 = ( i_5_  &  (~ i_3_)  &  (~ i_2_)  &  n_n503 ) ;
 assign wire1019 = ( (~ i_10_)  &  wire350 ) | ( (~ i_10_)  &  wire1021 ) ;
 assign wire1021 = ( i_7_  &  (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1023 = ( n_n764  &  wire1026 ) | ( n_n764  &  wire1027 ) ;
 assign wire1024 = ( (~ i_12_)  &  wire1030 ) | ( (~ i_12_)  &  wire7042 ) | ( (~ i_12_)  &  wire7043 ) ;
 assign wire1026 = ( i_5_  &  i_6_  &  i_4_ ) | ( i_6_  &  i_4_  &  (~ i_0_) ) ;
 assign wire1027 = ( i_5_  &  (~ i_3_)  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1030 = ( (~ i_10_)  &  i_8_  &  (~ i_5_)  &  n_n675 ) ;
 assign wire1033 = ( (~ i_12_)  &  wire1040 ) | ( (~ i_12_)  &  wire1041 ) | ( (~ i_12_)  &  wire7035 ) ;
 assign wire1040 = ( (~ i_6_)  &  (~ i_0_)  &  wire1043 ) | ( (~ i_6_)  &  (~ i_0_)  &  wire1044 ) ;
 assign wire1041 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_0_)  &  wire680 ) ;
 assign wire1042 = ( i_7_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1043 = ( (~ i_10_)  &  i_7_  &  (~ i_2_) ) ;
 assign wire1044 = ( (~ i_10_)  &  (~ i_7_)  &  i_8_  &  (~ i_3_) ) ;
 assign wire1047 = ( (~ i_9_)  &  (~ i_10_)  &  i_4_ ) ;
 assign wire1064 = ( (~ i_11_)  &  wire7017 ) | ( (~ i_11_)  &  wire7018 ) ;
 assign wire1067 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_1_) ) ;
 assign wire1074 = ( (~ i_9_)  &  i_5_  &  (~ i_6_)  &  (~ i_1_) ) ;
 assign wire1076 = ( (~ i_11_)  &  wire7009 ) | ( (~ i_11_)  &  n_n671  &  wire644 ) ;
 assign wire1082 = ( (~ i_6_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire1083 = ( (~ i_10_)  &  wire1089 ) | ( (~ i_10_)  &  wire7004 ) | ( (~ i_10_)  &  wire7005 ) ;
 assign wire1087 = ( (~ i_5_)  &  i_6_  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1089 = ( (~ i_8_)  &  wire1092 ) | ( (~ i_8_)  &  wire1093 ) ;
 assign wire1092 = ( i_4_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1093 = ( (~ i_5_)  &  i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1094 = ( (~ i_9_)  &  i_7_  &  i_8_  &  wire6994 ) ;
 assign wire1096 = ( (~ i_7_)  &  wire6996 ) | ( (~ i_7_)  &  wire19  &  wire301 ) ;
 assign wire1097 = ( i_7_  &  wire1103 ) | ( i_7_  &  n_n761  &  n_n672 ) ;
 assign wire1103 = ( i_2_  &  wire319 ) | ( (~ i_3_)  &  i_2_  &  wire335 ) ;
 assign wire1108 = ( wire14  &  wire1115 ) | ( wire14  &  wire1116 ) | ( wire14  &  wire1117 ) ;
 assign wire1109 = ( i_3_  &  wire1119 ) | ( i_3_  &  wire8  &  wire622 ) ;
 assign wire1110 = ( i_3_  &  (~ i_12_)  &  wire314 ) ;
 assign wire1115 = ( i_10_  &  (~ i_7_)  &  i_8_  &  i_12_ ) ;
 assign wire1116 = ( i_9_  &  i_10_  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1117 = ( i_9_  &  i_7_  &  i_8_  &  i_12_ ) ;
 assign wire1119 = ( i_9_  &  i_10_  &  (~ i_7_)  &  (~ i_11_) ) ;
 assign wire1121 = ( i_3_  &  wire1130 ) | ( i_3_  &  wire6983 ) ;
 assign wire1122 = ( i_9_  &  i_10_  &  i_13_  &  i_2_ ) ;
 assign wire1123 = ( (~ i_7_)  &  i_13_  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire1130 = ( i_9_  &  i_7_  &  i_8_  &  (~ i_12_) ) ;
 assign wire1132 = ( (~ i_2_)  &  wire118 ) | ( (~ i_2_)  &  wire365  &  wire615 ) ;
 assign wire1133 = ( i_9_  &  i_7_  &  i_13_  &  i_2_ ) ;
 assign wire1134 = ( i_3_  &  i_2_  &  n_n592 ) ;
 assign wire1135 = ( i_7_  &  i_13_  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire1139 = ( wire1152  &  wire6967 ) | ( wire23  &  n_n719  &  wire6967 ) ;
 assign wire1143 = ( (~ i_7_)  &  (~ i_8_)  &  wire369 ) ;
 assign wire1152 = ( (~ i_9_)  &  (~ i_3_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire1154 = ( (~ i_10_)  &  (~ i_13_)  &  i_11_  &  wire6963 ) ;
 assign wire1156 = ( (~ i_13_)  &  wire1160 ) | ( (~ i_13_)  &  n_n566  &  wire19 ) ;
 assign wire1160 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  i_4_ ) ;
 assign wire1162 = ( (~ i_7_)  &  wire329 ) ;
 assign wire1165 = ( (~ i_8_)  &  (~ i_3_)  &  (~ i_13_)  &  n_n741 ) ;
 assign wire1166 = ( (~ i_9_)  &  (~ i_3_)  &  (~ i_13_)  &  n_n701 ) ;
 assign wire1168 = ( n_n853  &  n_n672 ) | ( n_n853  &  wire1171 ) ;
 assign wire1169 = ( wire21  &  wire1173 ) | ( wire21  &  wire1175 ) | ( wire21  &  wire6959 ) ;
 assign wire1171 = ( (~ i_9_)  &  i_8_  &  i_4_  &  (~ i_2_) ) ;
 assign wire1173 = ( i_9_  &  i_7_  &  (~ i_12_) ) | ( i_7_  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire1175 = ( (~ i_12_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire1180 = ( i_9_  &  i_7_  &  i_12_  &  i_11_ ) ;
 assign wire1181 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1182 = ( i_9_  &  i_7_  &  (~ i_8_)  &  i_11_ ) ;
 assign wire1183 = ( i_10_  &  (~ i_7_)  &  i_12_  &  i_11_ ) ;
 assign wire1186 = ( (~ i_6_)  &  wire6945 ) | ( (~ i_6_)  &  wire636  &  wire6943 ) ;
 assign wire1194 = ( (~ i_13_)  &  (~ i_11_)  &  n_n273  &  n_n773 ) ;
 assign wire1195 = ( (~ i_6_)  &  wire1198 ) | ( (~ i_6_)  &  wire1199 ) ;
 assign wire1196 = ( wire336  &  wire371 ) | ( wire371  &  wire1348 ) ;
 assign wire1198 = ( n_n792  &  wire371 ) | ( n_n792  &  wire1200 ) ;
 assign wire1199 = ( n_n273  &  wire1202 ) | ( n_n273  &  wire1203 ) ;
 assign wire1200 = ( (~ i_3_)  &  (~ i_13_)  &  i_1_  &  (~ i_11_) ) ;
 assign wire1202 = ( (~ i_10_)  &  i_8_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1203 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire1204 = ( (~ i_6_)  &  (~ i_11_)  &  wire298 ) ;
 assign wire1213 = ( i_12_  &  wire393 ) ;
 assign wire1214 = ( i_9_  &  (~ i_7_)  &  i_6_  &  i_11_ ) ;
 assign wire1215 = ( i_10_  &  i_7_  &  (~ i_6_)  &  i_12_ ) ;
 assign wire1216 = ( i_10_  &  (~ i_7_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1217 = ( i_9_  &  i_7_  &  i_6_  &  i_12_ ) ;
 assign wire1218 = ( i_9_  &  i_8_  &  i_12_  &  wire6920 ) ;
 assign wire1221 = ( (~ i_6_)  &  wire1228 ) | ( (~ i_6_)  &  wire6925 ) ;
 assign wire1228 = ( (~ i_4_)  &  i_2_  &  wire1229 ) | ( (~ i_4_)  &  i_2_  &  wire1230 ) ;
 assign wire1229 = ( i_8_  &  i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire1230 = ( i_10_  &  i_8_  &  i_12_  &  (~ i_11_) ) ;
 assign wire1234 = ( i_2_  &  wire1239 ) | ( i_2_  &  wire8  &  wire515 ) ;
 assign wire1235 = ( i_9_  &  i_10_  &  i_1_  &  i_2_ ) ;
 assign wire1239 = ( i_9_  &  i_10_  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire1245 = ( (~ i_6_)  &  n_n534  &  n_n623 ) | ( (~ i_12_)  &  n_n534  &  n_n623 ) ;
 assign wire1246 = ( n_n421  &  wire1249 ) | ( n_n421  &  wire1250 ) ;
 assign wire1247 = ( n_n638  &  wire1252 ) | ( n_n638  &  n_n316  &  wire6908 ) ;
 assign wire1248 = ( i_3_  &  i_1_  &  i_11_  &  wire364 ) ;
 assign wire1249 = ( (~ i_7_)  &  i_6_  &  i_3_  &  (~ i_12_) ) ;
 assign wire1250 = ( (~ i_7_)  &  i_3_  &  i_1_ ) ;
 assign wire1252 = ( i_6_  &  i_3_  &  i_12_  &  i_1_ ) ;
 assign wire1255 = ( (~ i_12_)  &  i_11_  &  n_n592  &  wire6897 ) ;
 assign wire1263 = ( (~ i_8_)  &  wire1266 ) | ( (~ i_8_)  &  wire15  &  n_n415 ) ;
 assign wire1266 = ( i_10_  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire1267 = ( (~ i_4_)  &  i_1_  &  wire104 ) | ( (~ i_4_)  &  i_1_  &  wire1272 ) ;
 assign wire1272 = ( i_10_  &  (~ i_6_)  &  i_12_  &  i_11_ ) ;
 assign wire1274 = ( i_9_  &  wire272 ) | ( i_9_  &  wire1277 ) ;
 assign wire1277 = ( i_3_  &  (~ i_4_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire1279 = ( (~ i_12_)  &  (~ i_1_)  &  i_2_  &  wire493 ) ;
 assign wire1283 = ( i_3_  &  i_1_  &  wire1290 ) | ( i_3_  &  i_1_  &  wire6887 ) ;
 assign wire1290 = ( i_9_  &  i_10_  &  i_7_  &  i_12_ ) ;
 assign wire1293 = ( wire6875  &  wire6876 ) ;
 assign wire1294 = ( wire364  &  wire6879 ) | ( wire1301  &  wire6879 ) | ( wire1302  &  wire6879 ) ;
 assign wire1295 = ( wire297  &  wire1297 ) | ( wire297  &  wire1298 ) ;
 assign wire1296 = ( n_n346  &  wire1299 ) | ( n_n346  &  wire1300 ) ;
 assign wire1297 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  (~ i_1_) ) ;
 assign wire1298 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire1299 = ( i_10_  &  (~ i_8_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1300 = ( i_9_  &  (~ i_8_)  &  i_6_  &  i_11_ ) ;
 assign wire1301 = ( i_9_  &  i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire1302 = ( i_9_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire1307 = ( i_6_  &  i_13_  &  (~ i_12_)  &  (~ i_1_) ) ;
 assign wire1308 = ( i_13_  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire1314 = ( (~ i_10_)  &  (~ i_3_)  &  n_n545  &  n_n746 ) ;
 assign wire1315 = ( i_6_  &  (~ i_13_)  &  i_12_  &  wire346 ) ;
 assign wire1316 = ( wire301  &  wire6864 ) ;
 assign wire1317 = ( wire295  &  wire1321 ) | ( wire295  &  wire1338 ) | ( wire295  &  wire1339 ) ;
 assign wire1321 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_6_ ) ;
 assign wire1324 = ( (~ i_9_)  &  (~ i_10_)  &  wire19  &  wire6594 ) ;
 assign wire1326 = ( n_n273  &  wire1331 ) | ( n_n273  &  n_n274  &  n_n503 ) ;
 assign wire1327 = ( i_6_  &  wire1332 ) | ( i_6_  &  wire1333 ) ;
 assign wire1328 = ( (~ i_3_)  &  (~ i_2_)  &  n_n716  &  n_n503 ) ;
 assign wire1329 = ( wire371  &  wire1338 ) | ( wire371  &  wire1339 ) ;
 assign wire1331 = ( (~ i_9_)  &  i_6_  &  (~ i_13_)  &  i_4_ ) ;
 assign wire1332 = ( n_n764  &  wire371 ) | ( n_n764  &  wire1334 ) ;
 assign wire1333 = ( n_n716  &  wire1336 ) | ( n_n716  &  wire1337 ) ;
 assign wire1334 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_1_ ) ;
 assign wire1336 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_2_) ) ;
 assign wire1337 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign wire1338 = ( (~ i_9_)  &  i_7_  &  i_6_  &  (~ i_3_) ) ;
 assign wire1339 = ( (~ i_9_)  &  i_8_  &  i_6_  &  (~ i_2_) ) ;
 assign wire1340 = ( (~ i_9_)  &  (~ i_13_)  &  n_n701  &  wire6852 ) ;
 assign wire1341 = ( (~ i_13_)  &  i_12_  &  n_n741  &  wire6853 ) ;
 assign wire1343 = ( wire336  &  wire370 ) | ( wire370  &  wire1346 ) | ( wire370  &  wire1348 ) ;
 assign wire1344 = ( i_7_  &  (~ i_2_)  &  n_n566  &  wire32 ) ;
 assign wire1346 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire1348 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire1350 = ( wire1361  &  wire6843 ) | ( wire6842  &  wire6843 ) ;
 assign wire1351 = ( (~ i_3_)  &  i_1_  &  n_n819  &  wire381 ) ;
 assign wire1352 = ( (~ i_13_)  &  (~ i_12_)  &  n_n769  &  n_n273 ) ;
 assign wire1353 = ( i_6_  &  wire1355 ) | ( i_6_  &  (~ i_2_)  &  wire447 ) ;
 assign wire1354 = ( i_1_  &  n_n819  &  wire6848 ) ;
 assign wire1355 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  wire6846 ) ;
 assign wire1361 = ( (~ i_3_)  &  i_4_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1362 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_  &  wire6835 ) ;
 assign wire1363 = ( (~ i_8_)  &  i_6_  &  n_n716  &  n_n675 ) ;
 assign wire1366 = ( (~ i_6_)  &  wire1372 ) | ( (~ i_6_)  &  n_n675  &  wire6838 ) ;
 assign wire1372 = ( n_n764  &  wire1373 ) | ( n_n764  &  n_n545  &  wire31 ) ;
 assign wire1373 = ( (~ i_13_)  &  i_4_  &  (~ i_1_)  &  i_11_ ) ;
 assign wire1375 = ( wire1383  &  wire6831 ) | ( wire31  &  n_n792  &  wire6831 ) ;
 assign wire1376 = ( (~ i_8_)  &  i_11_  &  n_n779  &  n_n849 ) ;
 assign wire1377 = ( wire17  &  n_n675 ) | ( (~ i_1_)  &  wire17  &  wire440 ) ;
 assign wire1383 = ( (~ i_7_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1385 = ( i_9_  &  i_10_  &  wire6820 ) | ( i_9_  &  i_10_  &  wire6821 ) ;
 assign wire1388 = ( n_n665  &  wire287 ) | ( n_n665  &  wire1393 ) | ( n_n665  &  wire1394 ) ;
 assign wire1390 = ( i_13_  &  wire292 ) ;
 assign wire1391 = ( (~ i_5_)  &  i_3_  &  (~ i_4_)  &  wire6816 ) ;
 assign wire1392 = ( (~ i_6_)  &  n_n538  &  n_n716 ) ;
 assign wire1393 = ( i_5_  &  i_6_  &  i_3_  &  i_2_ ) ;
 assign wire1394 = ( i_5_  &  i_3_  &  i_1_  &  i_2_ ) ;
 assign wire1396 = ( (~ i_7_)  &  n_n826 ) | ( (~ i_7_)  &  n_n635 ) ;
 assign wire1397 = ( (~ i_7_)  &  (~ i_5_)  &  i_3_  &  i_1_ ) ;
 assign wire1400 = ( n_n498  &  n_n835  &  wire307  &  wire269 ) ;
 assign wire1402 = ( i_9_  &  i_10_  &  wire1406 ) | ( i_9_  &  i_10_  &  wire6812 ) ;
 assign wire1403 = ( wire272  &  wire1408 ) | ( wire272  &  wire1409 ) ;
 assign wire1406 = ( i_13_  &  (~ i_11_)  &  wire327 ) | ( i_13_  &  (~ i_11_)  &  wire384 ) ;
 assign wire1408 = ( i_9_  &  i_10_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire1409 = ( i_9_  &  i_10_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1410 = ( n_n592  &  wire272  &  wire6794 ) ;
 assign wire1412 = ( i_10_  &  wire583 ) ;
 assign wire1414 = ( n_n541  &  n_n830  &  n_n550  &  n_n837 ) ;
 assign wire1416 = ( n_n538  &  n_n838  &  n_n550 ) ;
 assign wire1418 = ( n_n538  &  n_n850  &  n_n716  &  wire6799 ) ;
 assign wire1419 = ( n_n833  &  n_n538  &  n_n550  &  n_n837 ) ;
 assign wire1423 = ( n_n795  &  n_n822  &  wire6785 ) ;
 assign wire1425 = ( (~ i_8_)  &  wire1432 ) | ( (~ i_8_)  &  wire1433 ) ;
 assign wire1432 = ( n_n822  &  wire24  &  wire576 ) ;
 assign wire1433 = ( n_n816  &  wire9  &  wire42 ) | ( n_n816  &  wire9  &  wire6788 ) ;
 assign wire1436 = ( n_n751  &  n_n846  &  n_n822  &  wire6775 ) ;
 assign wire1437 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6776 ) ;
 assign wire1438 = ( (~ i_7_)  &  (~ i_6_)  &  wire402 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire1444 ) ;
 assign wire1440 = ( (~ i_9_)  &  i_4_  &  n_n816  &  wire359 ) ;
 assign wire1441 = ( wire292  &  wire340 ) ;
 assign wire1444 = ( n_n816  &  wire1446 ) | ( n_n816  &  wire1447 ) ;
 assign wire1446 = ( (~ i_9_)  &  i_3_  &  i_4_  &  i_0_ ) ;
 assign wire1447 = ( (~ i_9_)  &  (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire1450 = ( n_n844  &  n_n843  &  n_n842  &  n_n851 ) ;
 assign wire1453 = ( n_n851  &  wire6770 ) | ( n_n833  &  n_n832  &  n_n851 ) ;
 assign wire1454 = ( n_n846  &  wire6771 ) | ( n_n846  &  wire6772 ) ;
 assign wire1462 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6762 ) ;
 assign wire1463 = ( n_n822  &  wire24  &  wire6763 ) ;
 assign wire1464 = ( wire327  &  n_n816  &  wire9 ) | ( n_n816  &  wire9  &  wire384 ) ;
 assign wire1466 = ( n_n849  &  wire6764 ) | ( n_n849  &  wire9  &  wire287 ) ;
 assign wire1472 = ( n_n850  &  n_n725  &  n_n852  &  n_n735 ) ;
 assign wire1474 = ( (~ i_8_)  &  (~ i_3_)  &  n_n741  &  wire521 ) ;
 assign wire1480 = ( (~ i_8_)  &  i_6_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire1481 = ( (~ i_8_)  &  i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign wire1488 = ( n_n849  &  n_n844  &  wire318 ) ;
 assign wire1490 = ( n_n764  &  wire1493 ) | ( n_n764  &  wire6749 ) | ( n_n764  &  wire6750 ) ;
 assign wire1493 = ( i_5_  &  (~ i_1_)  &  wire17 ) | ( i_5_  &  i_1_  &  wire37 ) ;
 assign wire1500 = ( n_n844  &  n_n751  &  n_n752  &  n_n846 ) ;
 assign wire1501 = ( (~ i_2_)  &  wire17  &  wire322 ) ;
 assign wire1502 = ( i_1_  &  i_0_  &  n_n764  &  wire37 ) ;
 assign wire1503 = ( n_n755  &  wire1506 ) | ( n_n755  &  n_n756  &  wire479 ) ;
 assign wire1504 = ( n_n853  &  wire51 ) | ( n_n853  &  n_n779  &  n_n768 ) ;
 assign wire1506 = ( n_n752  &  n_n840  &  n_n851 ) ;
 assign wire1511 = ( n_n795  &  wire1517 ) | ( i_4_  &  n_n795  &  wire451 ) ;
 assign wire1517 = ( (~ i_6_)  &  i_0_  &  wire369 ) ;
 assign wire1524 = ( n_n816  &  n_n795  &  wire6719 ) ;
 assign wire1525 = ( (~ i_8_)  &  wire420  &  n_n822  &  wire24 ) ;
 assign wire1526 = ( (~ i_5_)  &  wire17  &  wire336 ) ;
 assign wire1527 = ( i_2_  &  wire37  &  wire322 ) ;
 assign wire1528 = ( (~ i_8_)  &  (~ i_5_)  &  n_n779  &  wire313 ) ;
 assign wire1529 = ( (~ i_9_)  &  i_4_  &  wire313  &  wire6725 ) ;
 assign wire1530 = ( n_n853  &  n_n773  &  n_n771 ) ;
 assign wire1534 = ( n_n795  &  n_n498  &  wire13  &  wire298 ) ;
 assign wire1535 = ( wire1543  &  wire6709 ) | ( n_n453  &  wire569  &  wire6709 ) ;
 assign wire1537 = ( i_13_  &  (~ i_12_)  &  wire1542 ) | ( i_13_  &  (~ i_12_)  &  wire6714 ) ;
 assign wire1538 = ( n_n850  &  n_n570  &  n_n541  &  n_n213 ) ;
 assign wire1539 = ( n_n538  &  n_n498  &  n_n843 ) ;
 assign wire1542 = ( i_5_  &  i_6_  &  i_3_  &  wire314 ) ;
 assign wire1543 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_12_)  &  wire6708 ) ;
 assign wire1547 = ( i_13_  &  (~ i_12_)  &  wire1555 ) | ( i_13_  &  (~ i_12_)  &  wire6702 ) ;
 assign wire1552 = ( i_7_  &  i_8_  &  n_n658  &  n_n835 ) ;
 assign wire1553 = ( n_n833  &  n_n653  &  n_n651 ) ;
 assign wire1554 = ( n_n656  &  wire41 ) | ( n_n656  &  wire6698 ) ;
 assign wire1555 = ( (~ i_3_)  &  wire1558 ) | ( (~ i_3_)  &  n_n651  &  wire551 ) ;
 assign wire1558 = ( i_10_  &  i_5_  &  n_n746  &  n_n840 ) ;
 assign wire1562 = ( (~ i_9_)  &  i_7_  &  wire313  &  n_n685 ) ;
 assign wire1563 = ( n_n822  &  wire24  &  wire6686 ) ;
 assign wire1564 = ( n_n853  &  wire403 ) | ( n_n853  &  wire6687 ) | ( n_n853  &  wire6688 ) ;
 assign wire1565 = ( (~ i_10_)  &  (~ i_5_)  &  wire17  &  n_n675 ) ;
 assign wire1569 = ( n_n822  &  wire24  &  wire1574 ) | ( n_n822  &  wire24  &  wire1575 ) ;
 assign wire1571 = ( (~ i_7_)  &  (~ i_5_)  &  wire313  &  n_n685 ) ;
 assign wire1572 = ( n_n835  &  n_n761  &  n_n712  &  n_n752 ) ;
 assign wire1574 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_3_)  &  i_0_ ) ;
 assign wire1575 = ( (~ i_7_)  &  (~ i_3_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire1582 = ( wire1587  &  wire6670 ) | ( wire1588  &  wire6670 ) ;
 assign wire1583 = ( n_n822  &  wire24  &  wire6672 ) ;
 assign wire1584 = ( n_n853  &  wire6674 ) | ( n_n853  &  wire6675 ) ;
 assign wire1585 = ( (~ i_10_)  &  (~ i_6_)  &  wire17  &  n_n671 ) ;
 assign wire1587 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign wire1588 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1596 = ( n_n835  &  n_n787  &  n_n843  &  n_n710 ) ;
 assign wire1603 = ( n_n849  &  n_n746  &  n_n710 ) ;
 assign wire1605 = ( (~ i_9_)  &  (~ i_13_)  &  n_n701  &  wire277 ) ;
 assign wire1609 = ( n_n837  &  wire1612 ) | ( n_n837  &  wire1613 ) ;
 assign wire1610 = ( n_n832  &  wire1614 ) | ( n_n725  &  n_n832  &  wire541 ) ;
 assign wire1611 = ( n_n835  &  n_n716  &  n_n732  &  n_n837 ) ;
 assign wire1612 = ( n_n838  &  n_n725  &  n_n735 ) ;
 assign wire1613 = ( n_n755  &  n_n840  &  n_n710 ) ;
 assign wire1614 = ( n_n847  &  n_n755  &  n_n710 ) ;
 assign wire1620 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  n_n843 ) ;
 assign wire1624 = ( (~ i_9_)  &  n_n716  &  n_n732  &  n_n837 ) ;
 assign wire1629 = ( (~ i_13_)  &  i_12_  &  n_n741  &  wire6647 ) ;
 assign wire1630 = ( n_n844  &  n_n719  &  n_n837 ) ;
 assign wire1634 = ( i_13_  &  (~ i_12_)  &  n_n675  &  wire360 ) ;
 assign wire1635 = ( i_13_  &  (~ i_12_)  &  (~ i_11_)  &  wire6636 ) ;
 assign wire1637 = ( wire308  &  wire1639 ) | ( wire308  &  wire1640 ) ;
 assign wire1639 = ( i_6_  &  (~ i_3_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1640 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_2_) ) ;
 assign wire1643 = ( n_n658  &  wire25 ) | ( wire25  &  n_n683 ) | ( wire25  &  wire1644 ) ;
 assign wire1644 = ( i_5_  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire1647 = ( wire6630  &  wire6631 ) | ( n_n844  &  wire317  &  wire6631 ) ;
 assign wire1648 = ( i_9_  &  i_8_  &  wire453  &  wire6563 ) ;
 assign wire1652 = ( i_5_  &  i_6_  &  i_3_  &  wire6632 ) ;
 assign wire1656 = ( (~ i_1_)  &  i_2_  &  (~ i_0_)  &  n_n635 ) ;
 assign wire1661 = ( (~ i_13_)  &  n_n566  &  wire19  &  wire296 ) ;
 assign wire1663 = ( n_n746  &  wire294  &  n_n735 ) ;
 assign wire1669 = ( (~ i_4_)  &  i_2_  &  wire317 ) ;
 assign wire1672 = ( n_n716  &  n_n847  &  wire307  &  n_n756 ) ;
 assign wire1673 = ( n_n844  &  n_n752  &  n_n550  &  n_n732 ) ;
 assign wire1675 = ( n_n835  &  n_n545  &  n_n746  &  n_n735 ) ;
 assign wire1679 = ( n_n838  &  n_n746  &  n_n732 ) ;
 assign wire1681 = ( n_n752  &  n_n840  &  n_n735 ) ;
 assign wire1684 = ( wire344  &  n_n598  &  wire6594  &  wire6595 ) ;
 assign wire1685 = ( n_n746  &  n_n844  &  n_n575  &  n_n735 ) ;
 assign wire1686 = ( i_13_  &  (~ i_11_)  &  wire1692 ) | ( i_13_  &  (~ i_11_)  &  wire6603 ) ;
 assign wire1689 = ( n_n358  &  n_n840  &  wire6598 ) ;
 assign wire1691 = ( (~ i_7_)  &  (~ i_8_)  &  n_n835  &  n_n653 ) ;
 assign wire1692 = ( n_n581  &  wire1694 ) | ( (~ i_3_)  &  n_n581  &  wire468 ) ;
 assign wire1694 = ( i_5_  &  i_6_  &  (~ i_3_)  &  n_n833 ) ;
 assign wire1699 = ( wire1704  &  wire6588 ) | ( wire1705  &  wire6588 ) ;
 assign wire1702 = ( i_10_  &  (~ i_8_)  &  (~ i_11_)  &  wire6589 ) ;
 assign wire1703 = ( n_n830  &  n_n639  &  n_n597 ) ;
 assign wire1704 = ( i_13_  &  (~ i_12_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign wire1705 = ( (~ i_5_)  &  (~ i_6_)  &  i_13_ ) ;
 assign wire1708 = ( n_n832  &  n_n852  &  wire6578  &  wire6579 ) ;
 assign wire1709 = ( n_n635  &  n_n592  &  wire6582 ) ;
 assign wire1712 = ( n_n597  &  wire6584 ) | ( n_n833  &  n_n635  &  n_n597 ) ;
 assign wire1713 = ( n_n592  &  wire6585 ) | ( n_n847  &  n_n592  &  n_n633 ) ;
 assign wire1720 = ( (~ i_11_)  &  wire341  &  n_n752  &  n_n840 ) ;
 assign wire1721 = ( n_n844  &  n_n752  &  wire307 ) ;
 assign wire1722 = ( i_9_  &  i_11_  &  wire1724 ) | ( i_9_  &  i_11_  &  wire1725 ) ;
 assign wire1723 = ( n_n638  &  wire6575 ) | ( n_n638  &  n_n541  &  wire459 ) ;
 assign wire1724 = ( n_n570  &  n_n847  &  n_n541  &  n_n752 ) ;
 assign wire1725 = ( n_n835  &  n_n570  &  n_n541  &  n_n756 ) ;
 assign wire1726 = ( (~ i_5_)  &  i_6_  &  wire294  &  wire298 ) ;
 assign wire1729 = ( i_6_  &  n_n840  &  wire6573 ) ;
 assign wire1732 = ( i_9_  &  i_8_  &  wire434  &  wire6563 ) ;
 assign wire1740 = ( i_5_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire1741 = ( i_6_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1744 = ( i_9_  &  i_10_  &  wire6557  &  wire6558 ) ;
 assign wire1746 = ( i_5_  &  i_6_  &  wire6559 ) | ( i_6_  &  i_0_  &  wire6559 ) ;
 assign wire1748 = ( (~ i_6_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire1750 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_0_) ) ;
 assign wire1756 = ( i_9_  &  i_10_  &  i_8_  &  wire426 ) ;
 assign wire1763 = ( n_n838  &  n_n748  &  n_n725  &  wire341 ) ;
 assign wire1764 = ( n_n538  &  n_n850  &  n_n498  &  n_n835 ) ;
 assign wire1765 = ( i_9_  &  wire1767 ) | ( i_9_  &  wire1768 ) ;
 assign wire1766 = ( n_n833  &  wire6551 ) | ( n_n833  &  n_n541  &  wire423 ) ;
 assign wire1767 = ( n_n538  &  n_n725  &  n_n746  &  n_n830 ) ;
 assign wire1768 = ( n_n538  &  n_n835  &  n_n748  &  n_n716 ) ;
 assign wire1770 = ( wire341  &  n_n575  &  n_n756 ) ;
 assign wire1776 = ( i_9_  &  i_10_  &  i_1_ ) | ( i_10_  &  (~ i_6_)  &  i_1_ ) ;
 assign wire1778 = ( i_10_  &  (~ i_7_)  &  i_2_ ) ;
 assign wire1779 = ( i_9_  &  i_6_  &  i_1_ ) ;
 assign wire1780 = ( i_9_  &  i_10_  &  i_3_ ) | ( i_9_  &  i_10_  &  i_2_ ) ;
 assign wire1781 = ( i_9_  &  i_8_  &  i_3_ ) ;
 assign wire1789 = ( i_5_  &  wire1792 ) | ( i_5_  &  i_12_  &  wire683 ) ;
 assign wire1792 = ( i_9_  &  i_10_  &  i_12_  &  i_1_ ) ;
 assign wire1794 = ( i_9_  &  i_7_  &  i_6_  &  i_2_ ) ;
 assign wire1796 = ( (~ i_7_)  &  wire1803 ) | ( (~ i_7_)  &  wire1804 ) ;
 assign wire1797 = ( n_n844  &  wire6515 ) | ( n_n844  &  wire6516 ) ;
 assign wire1798 = ( i_10_  &  (~ i_6_)  &  i_1_  &  i_0_ ) ;
 assign wire1799 = ( i_8_  &  i_12_  &  i_11_  &  wire6509 ) ;
 assign wire1803 = ( (~ i_8_)  &  i_1_  &  i_11_  &  i_0_ ) ;
 assign wire1804 = ( i_3_  &  i_1_  &  i_11_  &  i_0_ ) ;
 assign wire1805 = ( n_n598  &  wire1810 ) | ( n_n598  &  wire6510 ) ;
 assign wire1806 = ( i_12_  &  i_11_ ) | ( i_11_  &  wire327 ) | ( i_11_  &  wire123 ) ;
 assign wire1808 = ( i_12_  &  wire287 ) ;
 assign wire1810 = ( i_10_  &  (~ i_7_)  &  i_11_ ) ;
 assign wire1814 = ( (~ i_7_)  &  wire1820 ) | ( (~ i_7_)  &  wire1821 ) ;
 assign wire1816 = ( i_9_  &  i_6_  &  i_1_  &  i_0_ ) ;
 assign wire1817 = ( i_9_  &  i_10_  &  i_0_ ) ;
 assign wire1820 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire1821 = ( (~ i_5_)  &  (~ i_6_)  &  i_3_  &  i_11_ ) ;
 assign wire1823 = ( wire36  &  wire1829 ) | ( i_2_  &  wire36  &  wire653 ) ;
 assign wire1825 = ( i_11_  &  wire384 ) ;
 assign wire1829 = ( i_7_  &  i_8_  &  i_12_ ) | ( i_7_  &  i_3_  &  i_12_ ) ;
 assign wire1832 = ( wire316  &  wire6494 ) | ( wire6493  &  wire6494 ) ;
 assign wire1833 = ( i_7_  &  wire1838 ) | ( i_7_  &  wire1839 ) ;
 assign wire1838 = ( i_8_  &  i_5_  &  i_6_  &  i_12_ ) ;
 assign wire1839 = ( i_5_  &  i_6_  &  i_3_  &  i_12_ ) ;
 assign wire1841 = ( wire379  &  wire30 ) | ( wire30  &  wire1844 ) | ( wire30  &  wire1845 ) ;
 assign wire1844 = ( i_10_  &  i_1_  &  i_11_  &  i_2_ ) ;
 assign wire1845 = ( (~ i_8_)  &  i_1_  &  i_11_ ) ;
 assign wire1848 = ( i_9_  &  i_10_  &  i_1_  &  i_11_ ) ;
 assign wire1849 = ( i_3_  &  i_1_  &  i_11_  &  i_2_ ) ;
 assign wire1850 = ( i_9_  &  i_10_  &  i_3_  &  i_13_ ) ;
 assign wire1852 = ( (~ i_4_)  &  n_n609 ) | ( (~ i_4_)  &  wire1856 ) | ( (~ i_4_)  &  wire1857 ) ;
 assign wire1853 = ( (~ i_8_)  &  (~ i_3_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire1856 = ( i_9_  &  i_8_  &  (~ i_12_) ) | ( i_8_  &  (~ i_3_)  &  (~ i_12_) ) ;
 assign wire1857 = ( i_9_  &  i_10_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire1861 = ( i_13_  &  wire1863 ) | ( i_13_  &  wire6478 ) ;
 assign wire1863 = ( i_9_  &  i_8_  &  i_3_ ) ;
 assign wire1867 = ( i_3_  &  wire319 ) | ( i_3_  &  n_n842  &  wire728 ) ;
 assign wire1869 = ( (~ i_8_)  &  wire369 ) ;
 assign wire6473 = ( (~ i_8_)  &  (~ i_11_) ) | ( (~ i_12_)  &  (~ i_11_) ) ;
 assign wire6474 = ( wire23  &  wire370 ) | ( wire277  &  wire6473 ) ;
 assign wire6475 = ( wire313  &  wire9 ) | ( i_8_  &  n_n761  &  wire9 ) ;
 assign wire6478 = ( i_10_  &  (~ i_8_)  &  i_3_ ) | ( i_10_  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire6479 = ( n_n453  &  wire308 ) | ( wire19  &  wire746 ) ;
 assign wire6485 = ( wire1850 ) | ( wire1853 ) | ( wire21  &  wire414 ) ;
 assign wire6488 = ( i_9_  &  i_1_  &  i_11_ ) ;
 assign wire6491 = ( n_n35  &  n_n612 ) | ( wire26  &  wire6488 ) ;
 assign wire6493 = ( i_8_  &  i_12_ ) | ( i_9_  &  i_10_  &  i_12_ ) ;
 assign wire6494 = ( i_5_  &  i_6_  &  i_2_ ) ;
 assign wire6495 = ( i_1_  &  wire395 ) | ( i_1_  &  wire34  &  n_n35 ) ;
 assign wire6496 = ( n_n633  &  wire299 ) | ( n_n612  &  wire316 ) ;
 assign wire6499 = ( i_12_  &  i_2_  &  i_0_ ) ;
 assign wire6500 = ( n_n36  &  wire385 ) | ( n_n358  &  wire6499 ) ;
 assign wire6501 = ( n_n818  &  (~ wire181) ) | ( i_1_  &  wire304 ) ;
 assign wire6504 = ( i_9_  &  i_5_  &  i_0_ ) | ( i_10_  &  (~ i_5_)  &  i_0_ ) ;
 assign wire6506 = ( wire6504 ) | ( (~ i_7_)  &  i_2_  &  wire304 ) ;
 assign wire6507 = ( wire1816 ) | ( wire1817 ) | ( wire385  &  wire660 ) ;
 assign wire6509 = ( i_7_  &  i_1_  &  i_0_ ) ;
 assign wire6510 = ( (~ i_8_)  &  i_11_ ) | ( i_9_  &  i_7_  &  i_11_ ) ;
 assign wire6512 = ( n_n36  &  wire388 ) | ( n_n35  &  wire6509 ) ;
 assign wire6515 = ( i_10_  &  (~ i_7_) ) | ( (~ i_8_)  &  i_11_ ) ;
 assign wire6516 = ( i_9_  &  i_7_ ) | ( i_8_  &  i_12_ ) ;
 assign wire6517 = ( wire292 ) | ( wire1798 ) ;
 assign wire6520 = ( wire1796 ) | ( wire1797 ) | ( wire1799 ) | ( wire6517 ) ;
 assign wire6522 = ( i_7_  &  i_5_  &  i_3_  &  i_1_ ) ;
 assign wire6523 = ( i_5_  &  (~ i_6_)  &  i_1_ ) ;
 assign wire6524 = ( i_9_  &  i_7_  &  i_12_ ) ;
 assign wire6526 = ( i_12_  &  wire6522 ) | ( i_10_  &  i_12_  &  wire6523 ) ;
 assign wire6527 = ( wire376  &  wire334 ) | ( n_n612  &  wire6524 ) ;
 assign wire6528 = ( wire6527 ) | ( wire6526 ) ;
 assign wire6530 = ( n_n877 ) | ( n_n876 ) | ( n_n878 ) ;
 assign wire6536 = ( wire126 ) | ( wire343 ) | ( wire1776 ) ;
 assign wire6537 = ( wire348 ) | ( wire386 ) | ( wire1778 ) | ( wire1779 ) ;
 assign wire6538 = ( wire1780 ) | ( wire1781 ) | ( wire278  &  wire327 ) ;
 assign wire6549 = ( i_9_  &  i_8_  &  (~ i_6_) ) ;
 assign wire6550 = ( i_9_  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire6551 = ( wire1770 ) | ( n_n538  &  n_n453  &  wire424 ) ;
 assign wire6553 = ( wire1763 ) | ( wire1764 ) | ( wire1765 ) ;
 assign wire6554 = ( i_7_  &  i_5_  &  (~ i_1_) ) ;
 assign wire6555 = ( wire12  &  n_n638 ) | ( n_n623  &  wire6554 ) ;
 assign wire6557 = ( (~ i_8_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire6558 = ( (~ i_7_)  &  (~ i_5_)  &  i_1_ ) | ( (~ i_7_)  &  i_1_  &  i_0_ ) ;
 assign wire6559 = ( i_9_  &  i_10_  &  i_8_  &  i_2_ ) ;
 assign wire6561 = ( wire1748 ) | ( (~ i_5_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire6562 = ( n_n835 ) | ( n_n606 ) | ( wire1750 ) ;
 assign wire6563 = ( (~ i_7_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire6567 = ( wire1732 ) | ( n_n665  &  wire425 ) | ( n_n665  &  wire435 ) ;
 assign wire6573 = ( i_3_  &  (~ i_4_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire6575 = ( wire1726 ) | ( wire1729 ) | ( wire272  &  wire375 ) ;
 assign wire6577 = ( wire1720 ) | ( wire1721 ) | ( wire1722 ) ;
 assign wire6578 = ( i_5_  &  i_9_ ) ;
 assign wire6579 = ( (~ i_3_)  &  i_13_  &  (~ i_11_) ) ;
 assign wire6582 = ( i_13_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire6584 = ( (~ i_0_)  &  wire265  &  n_n633 ) | ( i_0_  &  wire265  &  n_n631 ) ;
 assign wire6585 = ( n_n639  &  n_n840 ) | ( n_n852  &  n_n631 ) ;
 assign wire6587 = ( wire1708 ) | ( wire1709 ) | ( n_n453  &  wire308 ) ;
 assign wire6588 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_11_) ) ;
 assign wire6589 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_1_) ) ;
 assign wire6591 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) | ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire6593 = ( wire1699 ) | ( n_n665  &  wire1702 ) | ( n_n665  &  wire1703 ) ;
 assign wire6594 = ( (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6595 = ( i_8_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire6598 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_3_) ) ;
 assign wire6600 = ( i_9_  &  i_7_  &  (~ i_8_) ) ;
 assign wire6603 = ( wire1689 ) | ( wire1691 ) | ( wire469  &  wire6600 ) ;
 assign wire6604 = ( wire1685 ) | ( wire1684 ) ;
 assign wire6605 = ( wire6593 ) | ( wire6604 ) | ( wire337  &  wire465 ) ;
 assign wire6615 = ( wire1675 ) | ( wire1673 ) ;
 assign wire6616 = ( wire1672 ) | ( wire341  &  n_n852  &  wire482 ) ;
 assign wire6618 = ( i_7_  &  i_8_  &  (~ i_6_)  &  wire284 ) ;
 assign wire6620 = ( (~ i_3_)  &  (~ i_4_)  &  i_0_ ) ;
 assign wire6621 = ( i_8_  &  (~ i_5_)  &  (~ i_3_) ) ;
 assign wire6622 = ( i_8_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire6623 = ( i_1_  &  i_8_ ) ;
 assign wire6624 = ( n_n746  &  wire6620 ) | ( n_n346  &  wire6621 ) ;
 assign wire6627 = ( wire1661 ) | ( wire1663 ) | ( wire501  &  wire6618 ) ;
 assign wire6628 = ( i_8_  &  (~ i_5_)  &  i_6_  &  (~ i_3_) ) ;
 assign wire6629 = ( i_8_  &  i_5_  &  i_6_  &  (~ i_3_) ) ;
 assign wire6630 = ( n_n852  &  wire6628 ) | ( n_n847  &  wire6629 ) ;
 assign wire6631 = ( i_10_  &  (~ i_7_)  &  i_13_  &  (~ i_12_) ) ;
 assign wire6632 = ( i_13_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire6633 = ( n_n639  &  n_n852 ) | ( n_n840  &  n_n631 ) ;
 assign wire6636 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire6637 = ( i_5_  &  i_9_ ) ;
 assign wire6638 = ( (~ i_0_)  &  (~ i_3_) ) ;
 assign wire6640 = ( n_n675  &  wire6637 ) | ( n_n358  &  wire6638 ) ;
 assign wire6642 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire6643 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_)  &  n_n844 ) ;
 assign wire6644 = ( i_7_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign wire6645 = ( (~ i_13_)  &  i_12_  &  i_0_  &  n_n741 ) ;
 assign wire6647 = ( i_7_  &  (~ i_8_)  &  i_1_ ) ;
 assign wire6651 = ( wire517  &  wire6643 ) | ( wire518  &  wire6645 ) ;
 assign wire6653 = ( n_n832  &  n_n852 ) | ( n_n844  &  n_n837 ) ;
 assign wire6654 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_  &  n_n712 ) ;
 assign wire6658 = ( wire1611 ) | ( wire1620  &  wire6654 ) | ( wire6653  &  wire6654 ) ;
 assign wire6660 = ( (~ i_10_)  &  (~ i_13_)  &  i_12_  &  n_n748 ) ;
 assign wire6661 = ( (~ i_9_)  &  (~ i_13_)  &  i_11_  &  n_n850 ) ;
 assign wire6665 = ( wire543  &  wire6660 ) | ( wire544  &  wire6661 ) ;
 assign wire6667 = ( wire1596 ) | ( wire6665 ) | ( n_n844  &  wire545 ) ;
 assign wire6669 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire6670 = ( i_10_  &  i_13_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire6672 = ( (~ i_6_)  &  (~ i_3_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire6673 = ( (~ i_10_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire6674 = ( n_n671  &  n_n810 ) | ( n_n675  &  n_n813 ) ;
 assign wire6675 = ( n_n672  &  wire6673 ) | ( (~ i_9_)  &  wire12  &  n_n672 ) ;
 assign wire6678 = ( wire113 ) | ( wire1582 ) | ( wire1583 ) | ( wire1585 ) ;
 assign wire6683 = ( wire73 ) | ( wire1569 ) | ( wire1571 ) | ( wire1572 ) ;
 assign wire6686 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire6687 = ( n_n819  &  n_n678 ) | ( n_n819  &  n_n712 ) ;
 assign wire6688 = ( n_n699  &  n_n710 ) | ( n_n683  &  wire351 ) ;
 assign wire6693 = ( wire120 ) | ( wire1562 ) | ( wire1563 ) | ( wire1565 ) ;
 assign wire6694 = ( wire1564 ) | ( wire6693 ) ;
 assign wire6698 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_3_) ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire6702 = ( wire1552 ) | ( wire1553 ) | ( wire1554 ) ;
 assign wire6704 = ( n_n1250 ) | ( n_n1256 ) | ( n_n1255 ) | ( wire6667 ) ;
 assign wire6708 = ( i_10_  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign wire6709 = ( (~ i_1_)  &  i_2_  &  i_0_  &  n_n538 ) ;
 assign wire6712 = ( i_10_  &  i_3_  &  i_0_ ) ;
 assign wire6713 = ( i_9_  &  i_10_  &  i_3_  &  i_1_ ) ;
 assign wire6714 = ( n_n358  &  wire6712 ) | ( wire34  &  wire6713 ) ;
 assign wire6715 = ( wire1534 ) | ( n_n847  &  wire1538 ) | ( n_n847  &  wire1539 ) ;
 assign wire6719 = ( (~ i_5_)  &  i_4_  &  i_1_ ) ;
 assign wire6725 = ( i_8_  &  i_1_  &  i_2_ ) ;
 assign wire6730 = ( wire68 ) | ( wire1524 ) | ( wire1528 ) | ( wire1530 ) ;
 assign wire6731 = ( wire1525 ) | ( wire1526 ) | ( wire1527 ) | ( wire1529 ) ;
 assign wire6735 = ( (~ i_9_)  &  i_4_  &  i_1_ ) ;
 assign wire6737 = ( wire69 ) | ( wire70 ) | ( wire106 ) ;
 assign wire6745 = ( wire1500 ) | ( wire1501 ) | ( wire1502 ) ;
 assign wire6748 = ( i_0_  &  i_2_ ) ;
 assign wire6749 = ( wire12  &  wire295 ) | ( n_n853  &  n_n791 ) ;
 assign wire6750 = ( i_6_  &  (~ i_0_)  &  wire17 ) | ( i_6_  &  i_0_  &  wire37 ) ;
 assign wire6752 = ( wire1488 ) | ( wire37  &  wire494 ) ;
 assign wire6755 = ( (~ i_13_)  &  i_12_  &  n_n741  &  wire14 ) ;
 assign wire6756 = ( i_5_  &  (~ i_13_)  &  i_12_ ) ;
 assign wire6757 = ( wire1472 ) | ( wire1480  &  wire6755 ) | ( wire1481  &  wire6755 ) ;
 assign wire6759 = ( wire1474 ) | ( wire6757 ) | ( n_n755  &  wire523 ) ;
 assign wire6762 = ( i_7_  &  i_6_  &  i_3_ ) ;
 assign wire6763 = ( i_5_  &  (~ i_6_)  &  i_3_  &  i_2_ ) ;
 assign wire6764 = ( n_n819  &  n_n846 ) | ( n_n814  &  n_n813 ) ;
 assign wire6766 = ( wire1464 ) | ( wire37  &  wire606 ) ;
 assign wire6770 = ( n_n850  &  n_n852 ) | ( n_n838  &  n_n837 ) ;
 assign wire6771 = ( n_n835  &  n_n837 ) | ( n_n843  &  n_n840 ) ;
 assign wire6772 = ( n_n850  &  n_n847 ) | ( n_n830  &  n_n832 ) ;
 assign wire6773 = ( wire1450 ) | ( (~ i_9_)  &  i_4_  &  wire313 ) ;
 assign wire6775 = ( i_1_  &  (~ i_7_) ) ;
 assign wire6776 = ( i_6_  &  i_3_  &  i_2_ ) ;
 assign wire6777 = ( (~ i_9_)  &  i_4_  &  i_2_ ) ;
 assign wire6780 = ( wire1440 ) | ( wire1441 ) | ( n_n849  &  wire612 ) ;
 assign wire6782 = ( wire1436 ) | ( wire1437 ) | ( wire1438 ) | ( wire6780 ) ;
 assign wire6785 = ( (~ i_13_)  &  i_4_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire6787 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire6788 = ( (~ i_5_)  &  (~ i_6_)  &  i_2_ ) | ( (~ i_6_)  &  i_2_  &  i_0_ ) ;
 assign wire6789 = ( wire1423 ) | ( wire574  &  wire6787 ) ;
 assign wire6791 = ( wire1425 ) | ( wire6730 ) | ( wire6731 ) | ( wire6789 ) ;
 assign wire6794 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_11_) ) ;
 assign wire6799 = ( (~ i_2_)  &  (~ i_9_) ) ;
 assign wire6803 = ( i_5_  &  i_3_  &  (~ i_4_)  &  (~ i_12_) ) ;
 assign wire6805 = ( wire1410 ) | ( wire364  &  n_n840  &  wire6573 ) ;
 assign wire6806 = ( wire6805 ) | ( i_10_  &  i_11_  &  wire581 ) ;
 assign wire6807 = ( i_9_  &  i_10_  &  i_3_  &  (~ i_4_) ) ;
 assign wire6811 = ( i_6_  &  i_13_  &  (~ i_12_) ) ;
 assign wire6812 = ( wire272  &  wire276 ) | ( n_n818  &  wire6811 ) ;
 assign wire6814 = ( wire1403 ) | ( n_n421  &  wire268  &  wire410 ) ;
 assign wire6816 = ( i_6_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6819 = ( wire123 ) | ( wire359 ) | ( wire1397 ) ;
 assign wire6820 = ( wire1390 ) | ( n_n847  &  wire1391 ) | ( n_n847  &  wire1392 ) ;
 assign wire6821 = ( wire1388 ) | ( n_n637  &  wire1396 ) | ( n_n637  &  wire6819 ) ;
 assign wire6823 = ( wire1723 ) | ( wire1766 ) | ( wire6553 ) | ( wire6577 ) ;
 assign wire6824 = ( n_n1240 ) | ( n_n1241 ) | ( n_n1236 ) ;
 assign wire6825 = ( n_n1245 ) | ( wire1412 ) | ( wire6567 ) | ( wire6806 ) ;
 assign wire6827 = ( n_n1243 ) | ( wire1686 ) | ( wire6605 ) | ( wire6824 ) ;
 assign wire6828 = ( n_n1234 ) | ( wire1385 ) | ( wire6823 ) | ( wire6825 ) ;
 assign wire6831 = ( i_6_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire6834 = ( wire1377 ) | ( n_n853  &  wire438 ) ;
 assign wire6835 = ( i_7_  &  (~ i_6_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire6837 = ( (~ i_13_)  &  i_4_  &  i_12_  &  (~ i_1_) ) ;
 assign wire6838 = ( i_8_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6840 = ( i_6_  &  wire443 ) | ( n_n849  &  wire442 ) ;
 assign wire6842 = ( n_n779  &  wire309 ) | ( n_n685  &  wire267 ) ;
 assign wire6843 = ( (~ i_6_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire6846 = ( (~ i_3_)  &  (~ i_13_)  &  i_1_  &  (~ i_11_) ) ;
 assign wire6848 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire6850 = ( wire1351 ) | ( wire1352 ) | ( wire1354 ) ;
 assign wire6852 = ( (~ i_3_)  &  i_1_ ) | ( i_1_  &  (~ i_2_) ) ;
 assign wire6853 = ( (~ i_8_)  &  i_6_  &  (~ i_3_) ) ;
 assign wire6854 = ( (~ i_10_)  &  (~ i_6_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire6857 = ( wire1340 ) | ( wire1344 ) | ( n_n849  &  n_n810 ) ;
 assign wire6858 = ( wire1341 ) | ( wire1343 ) | ( n_n672  &  wire6854 ) ;
 assign wire6860 = ( wire1326 ) | ( wire1328 ) | ( wire1329 ) ;
 assign wire6864 = ( (~ i_10_)  &  i_8_  &  (~ i_6_)  &  (~ i_3_) ) ;
 assign wire6865 = ( n_n816  &  wire9 ) | ( wire29  &  wire294 ) ;
 assign wire6868 = ( wire1317 ) | ( (~ i_6_)  &  wire1324 ) | ( (~ i_6_)  &  wire6865 ) ;
 assign wire6869 = ( wire1314 ) | ( wire1315 ) | ( wire1316 ) | ( wire6868 ) ;
 assign wire6870 = ( wire1327 ) | ( wire6857 ) | ( wire6858 ) | ( wire6860 ) ;
 assign wire6871 = ( wire1307 ) | ( i_10_  &  (~ i_11_)  &  wire308 ) ;
 assign wire6872 = ( wire1308 ) | ( i_13_  &  (~ i_11_)  &  wire485 ) ;
 assign wire6873 = ( i_6_  &  wire487 ) | ( i_1_  &  wire486 ) ;
 assign wire6875 = ( (~ i_8_)  &  i_6_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire6876 = ( i_9_  &  (~ i_12_)  &  i_11_ ) | ( (~ i_12_)  &  (~ i_1_)  &  i_11_ ) ;
 assign wire6879 = ( (~ i_4_)  &  i_1_  &  i_11_ ) ;
 assign wire6884 = ( i_10_  &  i_1_  &  i_2_ ) ;
 assign wire6885 = ( i_2_  &  (~ i_6_) ) ;
 assign wire6886 = ( i_10_  &  (~ i_6_)  &  i_12_ ) ;
 assign wire6887 = ( n_n748  &  n_n197 ) | ( n_n638  &  wire6886 ) ;
 assign wire6888 = ( wire28  &  wire6884 ) | ( n_n656  &  wire6885 ) ;
 assign wire6890 = ( wire1279 ) | ( wire6888 ) | ( i_3_  &  wire491 ) ;
 assign wire6893 = ( (~ i_12_)  &  wire298 ) | ( wire22  &  wire334 ) ;
 assign wire6894 = ( wire272  &  wire311 ) | ( n_n412  &  wire363 ) ;
 assign wire6896 = ( wire1267 ) | ( wire6894 ) | ( n_n526  &  wire298 ) ;
 assign wire6897 = ( i_6_  &  i_3_  &  (~ i_1_) ) ;
 assign wire6899 = ( i_3_  &  (~ i_12_)  &  (~ i_1_)  &  i_2_ ) ;
 assign wire6900 = ( i_9_  &  i_8_  &  i_6_  &  i_12_ ) ;
 assign wire6901 = ( i_3_  &  i_12_  &  i_1_ ) ;
 assign wire6902 = ( (~ wire96)  &  n_n609 ) | ( n_n597  &  wire6901 ) ;
 assign wire6904 = ( wire15  &  wire104 ) | ( i_11_  &  wire15  &  wire6900 ) ;
 assign wire6905 = ( wire1255 ) | ( wire6904 ) | ( wire507  &  wire6899 ) ;
 assign wire6906 = ( i_9_  &  i_8_  &  i_6_ ) ;
 assign wire6908 = ( (~ i_6_)  &  i_3_  &  (~ i_1_) ) ;
 assign wire6911 = ( wire1245 ) | ( wire1247 ) | ( wire512  &  wire6906 ) ;
 assign wire6913 = ( i_7_  &  (~ i_6_)  &  i_3_  &  i_12_ ) ;
 assign wire6914 = ( i_9_  &  i_7_  &  (~ i_1_)  &  i_2_ ) ;
 assign wire6915 = ( wire1235 ) | ( n_n609  &  wire6913 ) ;
 assign wire6916 = ( n_n358  &  wire513 ) | ( wire516  &  wire6914 ) ;
 assign wire6918 = ( wire1234 ) | ( wire6915 ) | ( wire6916 ) ;
 assign wire6919 = ( wire1246 ) | ( wire1248 ) | ( wire6911 ) | ( wire6918 ) ;
 assign wire6920 = ( i_6_  &  (~ i_4_)  &  i_1_  &  i_2_ ) ;
 assign wire6921 = ( i_12_  &  i_7_ ) ;
 assign wire6922 = ( i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire6923 = ( (~ i_4_)  &  i_12_  &  i_1_ ) ;
 assign wire6924 = ( i_10_  &  i_8_  &  i_12_ ) ;
 assign wire6925 = ( n_n651  &  wire6923 ) | ( n_n346  &  wire6924 ) ;
 assign wire6926 = ( wire1218 ) | ( (~ i_4_)  &  i_1_  &  wire552 ) ;
 assign wire6929 = ( i_9_  &  (~ i_12_)  &  i_11_ ) | ( (~ i_12_)  &  (~ i_1_)  &  i_11_ ) ;
 assign wire6930 = ( i_12_  &  (~ i_1_)  &  (~ i_11_) ) ;
 assign wire6931 = ( (~ i_7_)  &  i_6_  &  wire6929 ) | ( i_7_  &  (~ i_6_)  &  wire6930 ) ;
 assign wire6934 = ( wire1204 ) | ( wire21  &  wire1213 ) | ( wire21  &  wire6931 ) ;
 assign wire6937 = ( n_n1112 ) | ( wire6934 ) | ( n_n369  &  wire604 ) ;
 assign wire6938 = ( n_n1129 ) | ( n_n1123 ) | ( n_n1128 ) | ( wire6919 ) ;
 assign wire6941 = ( wire1194 ) | ( wire1196 ) | ( wire313  &  wire9 ) ;
 assign wire6942 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_1_ ) ;
 assign wire6943 = ( (~ i_13_)  &  i_1_  &  (~ i_2_) ) ;
 assign wire6944 = ( i_7_  &  i_1_  &  (~ i_2_) ) ;
 assign wire6945 = ( wire635  &  wire6942 ) | ( n_n575  &  wire6944 ) ;
 assign wire6946 = ( i_1_  &  wire340 ) | ( (~ i_13_)  &  i_1_  &  wire632 ) ;
 assign wire6949 = ( n_n1108 ) | ( wire1350 ) | ( wire1353 ) | ( wire6850 ) ;
 assign wire6950 = ( n_n1121 ) | ( n_n1120 ) | ( wire6869 ) | ( wire6870 ) ;
 assign wire6952 = ( (~ i_8_)  &  (~ i_4_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire6954 = ( wire1182 ) | ( wire1180 ) ;
 assign wire6955 = ( wire104 ) | ( wire1181 ) | ( wire1183 ) ;
 assign wire6956 = ( n_n412  &  wire593 ) | ( wire594  &  wire6952 ) ;
 assign wire6958 = ( (~ i_8_)  &  (~ i_13_)  &  i_4_  &  (~ i_2_) ) ;
 assign wire6959 = ( i_10_  &  (~ i_7_)  &  (~ i_11_) ) | ( (~ i_7_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire6961 = ( wire25  &  n_n412 ) | ( n_n822  &  wire6958 ) ;
 assign wire6963 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_ ) ;
 assign wire6964 = ( n_n792  &  n_n274 ) | ( n_n570  &  n_n240 ) ;
 assign wire6965 = ( wire340 ) | ( wire1165 ) | ( wire1166 ) ;
 assign wire6966 = ( wire1156 ) | ( (~ i_3_)  &  wire1162 ) | ( (~ i_3_)  &  wire6964 ) ;
 assign wire6967 = ( i_2_  &  i_7_ ) ;
 assign wire6968 = ( (~ i_10_)  &  (~ i_3_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire6969 = ( n_n849  &  wire351 ) | ( wire352  &  wire6968 ) ;
 assign wire6970 = ( wire313  &  wire9 ) | ( n_n764  &  wire295 ) ;
 assign wire6972 = ( wire1139 ) | ( (~ i_3_)  &  wire616 ) ;
 assign wire6973 = ( wire6970 ) | ( (~ i_7_)  &  wire617 ) ;
 assign wire6975 = ( wire1143 ) | ( wire6969 ) | ( wire6972 ) | ( wire6973 ) ;
 assign wire6976 = ( i_8_  &  (~ i_4_)  &  i_2_ ) ;
 assign wire6978 = ( wire1135 ) | ( n_n432  &  wire6976 ) ;
 assign wire6979 = ( wire1133 ) | ( (~ i_8_)  &  i_3_  &  n_n656 ) ;
 assign wire6982 = ( i_9_  &  i_8_  &  (~ i_2_) ) ;
 assign wire6983 = ( n_n623  &  wire275 ) | ( n_n526  &  wire6982 ) ;
 assign wire6984 = ( wire1123 ) | ( i_10_  &  (~ i_11_)  &  wire308 ) ;
 assign wire6985 = ( wire1122 ) | ( i_3_  &  i_2_  &  n_n638 ) ;
 assign wire6987 = ( wire6984 ) | ( wire6985 ) | ( i_13_  &  wire626 ) ;
 assign wire6991 = ( n_n1191 ) | ( wire1110 ) | ( (~ i_4_)  &  wire619 ) ;
 assign wire6992 = ( wire1108 ) | ( wire1109 ) | ( wire1121 ) | ( wire6987 ) ;
 assign wire6994 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_)  &  i_2_ ) ;
 assign wire6995 = ( i_8_  &  i_4_  &  (~ i_2_) ) ;
 assign wire6996 = ( n_n787  &  n_n672 ) | ( n_n755  &  wire6995 ) ;
 assign wire6997 = ( wire1094 ) | ( i_7_  &  (~ i_2_)  &  wire628 ) ;
 assign wire6999 = ( n_n1189 ) | ( wire1168 ) | ( wire1169 ) | ( wire6961 ) ;
 assign wire7001 = ( n_n1187 ) | ( wire6991 ) | ( wire6992 ) | ( wire6999 ) ;
 assign wire7003 = ( i_4_  &  (~ i_7_) ) ;
 assign wire7004 = ( wire1087 ) | ( (~ i_7_)  &  (~ i_5_)  &  n_n685 ) ;
 assign wire7005 = ( wire35  &  n_n675 ) | ( n_n683  &  wire7003 ) ;
 assign wire7007 = ( n_n835  &  wire293 ) | ( n_n675  &  n_n813 ) ;
 assign wire7008 = ( wire7007 ) | ( n_n792  &  n_n791 ) ;
 assign wire7009 = ( wire1082 ) | ( n_n835  &  wire643 ) ;
 assign wire7010 = ( wire41  &  wire382 ) | ( (~ i_2_)  &  wire641 ) ;
 assign wire7011 = ( i_5_  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire7013 = ( i_5_  &  (~ i_3_)  &  (~ i_1_) ) ;
 assign wire7015 = ( (~ i_9_)  &  (~ i_8_)  &  i_5_ ) ;
 assign wire7017 = ( wire1067 ) | ( n_n675  &  wire7015 ) ;
 assign wire7018 = ( wire1074 ) | ( n_n275  &  wire646 ) | ( n_n275  &  wire7013 ) ;
 assign wire7019 = ( (~ i_5_)  &  wire265  &  n_n242 ) | ( i_5_  &  wire265  &  n_n277 ) ;
 assign wire7021 = ( n_n819  &  n_n678 ) | ( n_n671  &  n_n810 ) ;
 assign wire7022 = ( n_n819  &  n_n712 ) | ( n_n779  &  n_n768 ) ;
 assign wire7023 = ( n_n769  &  n_n771 ) | ( n_n835  &  wire318 ) ;
 assign wire7024 = ( wire12  &  wire346 ) | ( n_n764  &  n_n791 ) ;
 assign wire7027 = ( wire7021 ) | ( wire7024 ) | ( wire322  &  wire330 ) ;
 assign wire7028 = ( wire1047 ) | ( n_n773  &  n_n771 ) ;
 assign wire7029 = ( n_n699  &  n_n710 ) | ( n_n672  &  wire6673 ) ;
 assign wire7030 = ( wire35  &  wire336 ) | ( n_n699  &  n_n678 ) ;
 assign wire7032 = ( wire7030 ) | ( i_4_  &  wire676 ) ;
 assign wire7033 = ( i_5_  &  i_4_  &  (~ i_1_) ) ;
 assign wire7035 = ( wire1042 ) | ( (~ i_2_)  &  (~ i_0_)  &  n_n819 ) ;
 assign wire7037 = ( n_n683  &  wire351 ) | ( n_n764  &  wire7033 ) ;
 assign wire7038 = ( wire7037 ) | ( n_n827  &  n_n685 ) ;
 assign wire7039 = ( wire7022 ) | ( wire7023 ) | ( wire7027 ) | ( wire7038 ) ;
 assign wire7040 = ( wire1033 ) | ( wire7028 ) | ( wire7029 ) | ( wire7032 ) ;
 assign wire7041 = ( (~ i_2_)  &  (~ i_10_) ) ;
 assign wire7042 = ( wire267  &  n_n624 ) | ( n_n675  &  n_n768 ) ;
 assign wire7043 = ( (~ wire55)  &  wire322 ) | ( wire317  &  wire7041 ) ;
 assign wire7045 = ( wire1023 ) | ( i_7_  &  (~ i_2_)  &  n_n566 ) ;
 assign wire7046 = ( n_n741  &  wire275 ) | ( (~ i_8_)  &  (~ i_3_)  &  n_n741 ) ;
 assign wire7047 = ( n_n242  &  n_n606 ) | ( n_n624  &  n_n277 ) ;
 assign wire7050 = ( wire321 ) | ( i_8_  &  (~ i_3_)  &  n_n835 ) ;
 assign wire7051 = ( n_n769  &  n_n671 ) | ( n_n240  &  wire698 ) ;
 assign wire7054 = ( wire1024 ) | ( wire7045 ) | ( n_n566  &  wire19 ) ;
 assign wire7057 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_11_)  &  (~ i_2_) ) ;
 assign wire7058 = ( (~ i_9_)  &  i_7_  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire7059 = ( n_n773  &  wire7057 ) | ( n_n658  &  wire7058 ) ;
 assign wire7060 = ( wire988 ) | ( n_n701  &  n_n606 ) | ( n_n701  &  wire993 ) ;
 assign wire7062 = ( wire987 ) | ( wire7059 ) | ( wire7060 ) ;
 assign wire7063 = ( wire1076 ) | ( wire7010 ) | ( wire7062 ) ;
 assign wire7065 = ( n_n910 ) | ( wire7039 ) | ( wire7040 ) | ( wire7063 ) ;
 assign wire7066 = ( (~ i_5_)  &  i_4_  &  (~ i_1_) ) ;
 assign wire7067 = ( (~ i_11_)  &  (~ i_8_) ) ;
 assign wire7068 = ( i_5_  &  i_6_  &  (~ i_3_)  &  (~ i_12_) ) ;
 assign wire7070 = ( n_n741  &  wire326 ) | ( n_n792  &  wire7066 ) ;
 assign wire7071 = ( n_n701  &  wire323 ) | ( n_n566  &  wire325 ) ;
 assign wire7074 = ( wire970 ) | ( wire971 ) | ( wire7070 ) | ( wire7071 ) ;
 assign wire7076 = ( wire972 ) | ( wire1083 ) | ( wire7008 ) | ( wire7074 ) ;
 assign wire7077 = ( (~ i_1_)  &  (~ i_13_) ) ;
 assign wire7078 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_12_)  &  i_0_ ) ;
 assign wire7079 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire7080 = ( n_n842  &  n_n710 ) | ( wire30  &  wire7079 ) ;
 assign wire7082 = ( wire960 ) | ( wire962 ) | ( wire529  &  wire7077 ) ;
 assign wire7083 = ( (~ i_5_)  &  (~ i_3_)  &  i_0_ ) ;
 assign wire7084 = ( wire11  &  n_n670 ) | ( n_n843  &  wire16 ) ;
 assign wire7085 = ( (~ i_10_)  &  (~ i_13_)  &  i_4_ ) ;
 assign wire7086 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire7087 = ( i_0_  &  (~ i_11_) ) ;
 assign wire7088 = ( wire948 ) | ( wire533  &  wire7083 ) ;
 assign wire7091 = ( n_n566  &  wire19 ) | ( i_7_  &  (~ i_2_)  &  n_n566 ) ;
 assign wire7092 = ( wire340 ) | ( (~ i_2_)  &  n_n701  &  n_n751 ) ;
 assign wire7093 = ( wire1165 ) | ( wire1166 ) | ( wire7092 ) ;
 assign wire7094 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_11_) ) ;
 assign wire7100 = ( i_5_  &  i_6_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire7102 = ( wire927 ) | ( wire12  &  n_n670  &  wire579 ) ;
 assign wire7104 = ( (~ i_5_)  &  i_6_  &  (~ i_1_) ) ;
 assign wire7105 = ( n_n849  &  n_n813 ) | ( wire294  &  wire7104 ) ;
 assign wire7107 = ( wire7105 ) | ( (~ i_13_)  &  i_11_  &  wire666 ) ;
 assign wire7108 = ( wire70 ) | ( wire917 ) | ( n_n816  &  wire667 ) ;
 assign wire7109 = ( i_8_  &  (~ i_13_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire7110 = ( n_n819  &  n_n712 ) | ( n_n764  &  wire7033 ) ;
 assign wire7111 = ( n_n827  &  n_n685 ) | ( n_n624  &  n_n277 ) ;
 assign wire7113 = ( wire907 ) | ( n_n716  &  wire669 ) ;
 assign wire7114 = ( (~ i_5_)  &  (~ i_13_)  &  i_4_  &  i_11_ ) ;
 assign wire7115 = ( n_n816  &  wire671 ) | ( wire336  &  wire7114 ) ;
 assign wire7117 = ( wire896 ) | ( wire7107 ) | ( wire7108 ) ;
 assign wire7118 = ( wire895 ) | ( wire909 ) | ( wire7113 ) | ( wire7115 ) ;
 assign wire7119 = ( i_5_  &  (~ i_3_)  &  i_0_ ) ;
 assign wire7121 = ( i_5_  &  i_6_  &  (~ i_1_)  &  i_0_ ) ;
 assign wire7122 = ( n_n675  &  n_n813 ) | ( n_n277  &  wire7011 ) ;
 assign wire7126 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_0_) ) ;
 assign wire7127 = ( i_7_  &  (~ i_3_)  &  i_4_  &  (~ i_0_) ) ;
 assign wire7128 = ( wire319 ) | ( (~ i_8_)  &  (~ i_3_)  &  n_n719 ) ;
 assign wire7129 = ( n_n712  &  n_n751 ) | ( n_n570  &  n_n827 ) ;
 assign wire7130 = ( wire26  &  wire638 ) | ( wire284  &  wire637 ) ;
 assign wire7132 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire7133 = ( (~ i_0_)  &  (~ i_1_) ) ;
 assign wire7134 = ( (~ i_8_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire7136 = ( (~ i_0_)  &  (~ i_2_) ) ;
 assign wire7138 = ( (~ i_5_)  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire7140 = ( wire405 ) | ( wire856 ) | ( wire859 ) ;
 assign wire7144 = ( (~ i_5_)  &  i_6_  &  i_4_ ) ;
 assign wire7146 = ( n_n176  &  n_n771 ) | ( n_n671  &  wire7144 ) ;
 assign wire7149 = ( wire843 ) | ( wire844 ) | ( wire846 ) ;
 assign wire7151 = ( wire845 ) | ( wire7130 ) | ( n_n838  &  wire639 ) ;
 assign wire7155 = ( wire834 ) | ( wire835 ) | ( wire17  &  wire6669 ) ;
 assign wire7157 = ( n_n773  &  n_n771 ) | ( n_n683  &  wire351 ) ;
 assign wire7161 = ( wire68 ) | ( wire69 ) | ( wire106 ) | ( wire120 ) ;
 assign wire7163 = ( i_5_  &  (~ i_0_)  &  n_n843 ) ;
 assign wire7164 = ( i_5_  &  (~ i_13_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire7165 = ( (~ i_10_)  &  (~ i_8_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire7167 = ( wire121 ) | ( wire814 ) | ( wire725  &  wire7164 ) ;
 assign wire7168 = ( wire13  &  wire723 ) | ( wire724  &  wire7163 ) ;
 assign wire7174 = ( i_7_  &  i_5_  &  n_n687 ) ;
 assign wire7175 = ( i_5_  &  (~ i_6_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire7177 = ( wire798 ) | ( wire800 ) | ( wire735  &  wire7174 ) ;
 assign wire7178 = ( i_5_  &  i_9_ ) ;
 assign wire7181 = ( i_9_  &  i_8_  &  i_5_  &  i_12_ ) ;
 assign wire7182 = ( i_10_  &  i_6_  &  i_12_  &  i_0_ ) ;
 assign wire7183 = ( (~ i_5_)  &  i_6_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7184 = ( (~ i_5_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire7185 = ( n_n638  &  wire7182 ) | ( n_n651  &  wire7183 ) ;
 assign wire7188 = ( i_9_  &  i_3_  &  i_12_  &  i_2_ ) ;
 assign wire7190 = ( i_9_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7191 = ( wire362 ) | ( n_n818  &  wire686 ) ;
 assign wire7194 = ( i_5_  &  i_6_  &  i_0_ ) ;
 assign wire7196 = ( wire255 ) | ( wire258 ) | ( (~ i_4_)  &  wire717 ) ;
 assign wire7199 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire7200 = ( (~ i_7_)  &  i_3_  &  (~ i_4_)  &  i_0_ ) ;
 assign wire7202 = ( i_10_  &  (~ i_8_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire7203 = ( wire297  &  n_n840 ) | ( n_n346  &  wire342 ) ;
 assign wire7205 = ( wire245 ) | ( wire296  &  wire7202 ) ;
 assign wire7208 = ( i_10_  &  i_12_  &  (~ i_11_) ) | ( i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire7211 = ( n_n840  &  wire6573 ) | ( n_n840  &  wire6803 ) ;
 assign wire7214 = ( wire235 ) | ( wire236 ) | ( wire7211 ) ;
 assign wire7215 = ( i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7218 = ( i_3_  &  (~ i_4_)  &  i_2_  &  i_0_ ) ;
 assign wire7219 = ( i_12_  &  (~ i_11_)  &  i_2_ ) ;
 assign wire7222 = ( wire115 ) | ( wire225 ) | ( wire737  &  wire7218 ) ;
 assign wire7223 = ( (~ i_12_)  &  i_11_  &  i_2_ ) ;
 assign wire7226 = ( (~ i_5_)  &  i_12_  &  (~ i_11_)  &  (~ i_0_) ) ;
 assign wire7227 = ( i_10_  &  i_12_  &  i_0_ ) ;
 assign wire7228 = ( i_7_  &  i_5_  &  i_0_ ) ;
 assign wire7229 = ( wire741  &  wire7227 ) | ( wire270  &  wire7228 ) ;
 assign wire7231 = ( wire212 ) | ( wire213 ) | ( (~ i_4_)  &  wire738 ) ;
 assign wire7232 = ( wire237 ) | ( wire238 ) | ( wire7214 ) | ( wire7231 ) ;
 assign wire7233 = ( wire215 ) | ( wire7222 ) | ( n_n541  &  wire736 ) ;
 assign wire7234 = ( (~ i_8_)  &  (~ i_4_)  &  i_2_ ) ;
 assign wire7235 = ( i_5_  &  (~ i_6_)  &  (~ i_12_)  &  i_11_ ) ;
 assign wire7237 = ( i_10_  &  (~ i_4_)  &  i_11_ ) ;
 assign wire7239 = ( i_5_  &  (~ i_12_)  &  i_11_ ) ;
 assign wire7241 = ( wire198 ) | ( wire200 ) | ( wire744  &  wire7237 ) ;
 assign wire7244 = ( n_n987 ) | ( n_n986 ) | ( wire201 ) | ( wire7241 ) ;
 assign wire7246 = ( (~ i_7_)  &  (~ i_5_)  &  i_2_  &  i_0_ ) ;
 assign wire7248 = ( i_10_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire7249 = ( (~ i_12_)  &  i_11_  &  (~ i_0_) ) ;
 assign wire7250 = ( (~ i_7_)  &  i_5_  &  (~ i_6_)  &  i_2_ ) ;
 assign wire7251 = ( n_n415  &  wire7246 ) | ( n_n598  &  wire7248 ) ;
 assign wire7253 = ( wire190 ) | ( wire7251 ) | ( i_10_  &  wire557 ) ;
 assign wire7254 = ( (~ i_7_)  &  i_6_  &  i_2_ ) ;
 assign wire7255 = ( wire11  &  wire558 ) | ( wire338  &  wire7254 ) ;
 assign wire7257 = ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7260 = ( wire163 ) | ( n_n421  &  n_n598 ) | ( n_n421  &  wire166 ) ;
 assign wire7261 = ( wire283  &  wire565 ) | ( i_2_  &  wire564 ) ;
 assign wire7262 = ( wire7261 ) | ( wire7260 ) ;
 assign wire7263 = ( n_n1000 ) | ( wire192 ) | ( wire7253 ) ;
 assign wire7264 = ( i_9_  &  i_8_  &  i_2_ ) ;
 assign wire7266 = ( i_5_  &  i_12_  &  i_2_  &  i_0_ ) ;
 assign wire7267 = ( i_8_  &  i_3_  &  i_2_  &  i_0_ ) ;
 assign wire7268 = ( i_9_  &  i_10_  &  i_8_  &  (~ i_5_) ) ;
 assign wire7269 = ( i_9_  &  i_3_  &  i_12_  &  i_1_ ) ;
 assign wire7271 = ( wire397  &  wire7267 ) | ( wire292  &  wire7268 ) ;
 assign wire7272 = ( wire154 ) | ( n_n185  &  wire700 ) ;
 assign wire7273 = ( wire150 ) | ( wire7271 ) | ( wire701  &  wire7266 ) ;
 assign wire7275 = ( (~ i_7_)  &  i_8_  &  i_5_ ) ;
 assign wire7277 = ( wire143 ) | ( wire18  &  wire354  &  wire704 ) ;
 assign wire7278 = ( wire139 ) | ( wire141 ) | ( wire142 ) ;
 assign wire7279 = ( wire7277 ) | ( i_9_  &  i_11_  &  wire703 ) ;
 assign wire7280 = ( i_10_  &  (~ i_8_)  &  i_3_ ) ;
 assign wire7282 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_) ) ;
 assign wire7286 = ( i_10_  &  i_3_  &  i_12_  &  i_0_ ) ;
 assign wire7287 = ( i_10_  &  (~ i_5_)  &  i_6_  &  i_12_ ) ;
 assign wire7288 = ( (~ i_5_)  &  i_3_  &  i_0_ ) ;
 assign wire7289 = ( n_n421  &  wire123 ) | ( n_n358  &  wire7286 ) ;
 assign wire7292 = ( wire7289 ) | ( (~ i_8_)  &  wire596 ) ;
 assign wire7293 = ( wire127 ) | ( wire128 ) | ( wire129 ) | ( wire130 ) ;
 assign wire7294 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_0_) ) ;
 assign wire7295 = ( i_5_  &  i_3_  &  (~ i_12_)  &  i_1_ ) ;
 assign wire7296 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_)  &  i_3_ ) ;
 assign wire7297 = ( n_n453  &  wire308 ) | ( n_n637  &  wire706 ) ;
 assign wire7300 = ( wire103 ) | ( wire107 ) | ( wire112 ) | ( wire7297 ) ;
 assign wire7302 = ( i_7_  &  (~ i_8_)  &  i_6_  &  i_3_ ) ;
 assign wire7303 = ( i_10_  &  (~ i_8_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire7304 = ( i_10_  &  i_11_  &  (~ i_0_) ) ;
 assign wire7307 = ( n_n609  &  wire359 ) | ( wire287  &  wire7303 ) ;
 assign wire7308 = ( wire86 ) | ( wire89 ) | ( wire338  &  wire7302 ) ;
 assign wire7309 = ( wire7307 ) | ( (~ i_8_)  &  wire97 ) | ( (~ i_8_)  &  wire98 ) ;
 assign wire7310 = ( wire7292 ) | ( wire7293 ) | ( wire7308 ) ;
 assign wire7311 = ( wire7300 ) | ( wire7309 ) | ( n_n213  &  wire705 ) ;
 assign wire7312 = ( i_9_  &  i_10_  &  i_11_  &  i_0_ ) ;
 assign wire7313 = ( i_9_  &  i_7_  &  i_6_  &  i_2_ ) ;
 assign wire7314 = ( (~ i_5_)  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign wire7317 = ( wire64 ) | ( wire65 ) | ( wire314  &  wire7314 ) ;
 assign wire7318 = ( wire7317 ) | ( i_9_  &  i_7_  &  wire752 ) ;
 assign wire7319 = ( wire7272 ) | ( wire7273 ) | ( wire7278 ) | ( wire7279 ) ;
 assign wire7321 = ( wire7262 ) | ( wire7263 ) | ( wire7310 ) | ( wire7311 ) ;
 assign wire7322 = ( (~ i_8_)  &  (~ i_5_)  &  i_4_ ) ;
 assign wire7324 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire7325 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_5_) ) ;
 assign wire7326 = ( (~ i_10_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire7327 = ( wire325  &  n_n575 ) | ( wire281  &  wire7326 ) ;
 assign wire7329 = ( wire313  &  wire9 ) | ( n_n729  &  wire7324 ) ;
 assign wire7335 = ( n_n970 ) | ( n_n957 ) | ( wire961 ) | ( wire7082 ) ;
 assign wire7336 = ( n_n978 ) | ( n_n976 ) | ( wire7117 ) | ( wire7118 ) ;
 assign wire7337 = ( n_n972 ) | ( n_n962 ) | ( wire801 ) | ( wire7177 ) ;
 assign wire7338 = ( n_n981 ) | ( wire7149 ) | ( wire7151 ) | ( wire7335 ) ;
 assign wire7339 = ( wire7318 ) | ( wire7319 ) | ( wire7321 ) | ( wire7336 ) ;


endmodule

