module ex1010 (
	i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, 
	i_2_, i_0_, o_1_, o_2_, o_0_, o_9_, o_7_, o_8_, o_5_, o_6_, 
	o_3_, o_4_);

input i_9_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_3_;
input i_4_;
input i_1_;
input i_2_;
input i_0_;
output o_1_;
output o_2_;
output o_0_;
output o_9_;
output o_7_;
output o_8_;
output o_5_;
output o_6_;
output o_3_;
output o_4_;
wire n_n1014;
wire n_n4309;
wire n_n1005;
wire n_n1004;
wire n_n1396;
wire n_n1397;
wire n_n1398;
wire n_n5305;
wire n_n5293;
wire n_n5296;
wire n_n5284;
wire n_n543;
wire n_n562;
wire n_n561;
wire n_n563;
wire n_n5297;
wire n_n3936;
wire n_n3920;
wire n_n3937;
wire n_n3187;
wire n_n3192;
wire n_n3191;
wire n_n3622;
wire n_n3624;
wire n_n3625;
wire n_n3626;
wire wire148;
wire n_n2530;
wire n_n2531;
wire n_n2525;
wire n_n2523;
wire n_n2845;
wire n_n2846;
wire n_n2827;
wire n_n2821;
wire n_n2826;
wire n_n2907;
wire n_n2906;
wire n_n2908;
wire n_n2898;
wire n_n1793;
wire n_n1792;
wire n_n1794;
wire n_n1784;
wire n_n1787;
wire n_n1786;
wire n_n2104;
wire n_n2087;
wire n_n2086;
wire n_n2166;
wire n_n2105;
wire n_n2155;
wire wire16;
wire n_n4338;
wire wire21;
wire n_n4339;
wire wire22;
wire n_n4337;
wire n_n4401;
wire n_n4403;
wire n_n4400;
wire wire13;
wire n_n4464;
wire n_n4467;
wire wire11;
wire n_n4463;
wire wire10;
wire n_n4666;
wire wire24;
wire n_n4667;
wire n_n4664;
wire n_n4737;
wire wire14;
wire n_n4738;
wire n_n4735;
wire n_n4782;
wire n_n4784;
wire n_n4779;
wire wire17;
wire n_n4830;
wire n_n4831;
wire n_n4900;
wire n_n4902;
wire n_n4898;
wire wire18;
wire n_n4976;
wire n_n4977;
wire n_n4975;
wire n_n5038;
wire n_n5040;
wire n_n5034;
wire wire12;
wire n_n5092;
wire wire20;
wire n_n5093;
wire n_n5091;
wire n_n4440;
wire n_n4434;
wire n_n4432;
wire wire98;
wire wire233;
wire wire236;
wire n_n4720;
wire n_n4216;
wire n_n4857;
wire n_n4862;
wire n_n4856;
wire wire40;
wire wire102;
wire wire245;
wire n_n4991;
wire n_n4996;
wire n_n4992;
wire n_n4995;
wire n_n4990;
wire n_n4998;
wire n_n4999;
wire wire103;
wire wire25;
wire n_n4617;
wire wire15;
wire n_n4637;
wire n_n4613;
wire n_n4927;
wire n_n4958;
wire n_n4920;
wire n_n4325;
wire wire23;
wire n_n4327;
wire n_n4324;
wire n_n4382;
wire n_n4383;
wire n_n4380;
wire n_n4923;
wire n_n4924;
wire n_n4921;
wire n_n4982;
wire n_n4983;
wire n_n4981;
wire n_n5035;
wire n_n5032;
wire n_n5111;
wire n_n5112;
wire n_n5109;
wire n_n5171;
wire n_n5174;
wire n_n5167;
wire n_n4597;
wire n_n4598;
wire n_n4602;
wire n_n4593;
wire n_n4601;
wire wire108;
wire n_n4744;
wire n_n4754;
wire n_n4757;
wire n_n4749;
wire n_n4756;
wire wire109;
wire n_n4887;
wire n_n4888;
wire n_n4885;
wire n_n3450;
wire n_n4882;
wire n_n3451;
wire n_n5026;
wire n_n5027;
wire n_n5025;
wire wire114;
wire n_n5181;
wire n_n5184;
wire n_n5183;
wire wire112;
wire n_n5310;
wire n_n5318;
wire n_n5314;
wire n_n5320;
wire wire459;
wire n_n4615;
wire n_n4616;
wire n_n4607;
wire wire396;
wire n_n3346;
wire n_n4641;
wire n_n4634;
wire n_n4648;
wire n_n4618;
wire n_n4628;
wire wire26;
wire wire118;
wire wire309;
wire n_n3281;
wire n_n5050;
wire n_n5060;
wire n_n5055;
wire n_n5054;
wire n_n5059;
wire n_n5048;
wire n_n5028;
wire n_n5036;
wire wire50;
wire wire230;
wire wire231;
wire wire356;
wire n_n4571;
wire n_n4578;
wire n_n4570;
wire n_n4849;
wire n_n4853;
wire n_n4847;
wire n_n5096;
wire n_n5099;
wire n_n5085;
wire n_n4314;
wire n_n4389;
wire n_n4369;
wire n_n4381;
wire n_n4340;
wire wire280;
wire n_n5101;
wire n_n5110;
wire n_n5142;
wire n_n5107;
wire n_n5130;
wire n_n5123;
wire n_n5129;
wire n_n5156;
wire n_n4317;
wire n_n4318;
wire n_n4388;
wire n_n4459;
wire n_n4461;
wire n_n4455;
wire n_n4513;
wire n_n4515;
wire n_n4512;
wire n_n4790;
wire n_n4791;
wire n_n4787;
wire n_n4859;
wire n_n4860;
wire n_n4858;
wire n_n4926;
wire n_n4928;
wire n_n4925;
wire n_n4988;
wire n_n4987;
wire n_n5041;
wire n_n5042;
wire n_n5100;
wire n_n4724;
wire n_n4727;
wire n_n4739;
wire wire95;
wire wire244;
wire n_n4864;
wire n_n4868;
wire n_n5018;
wire n_n5022;
wire n_n5017;
wire wire135;
wire wire296;
wire n_n4993;
wire n_n1576;
wire wire134;
wire wire252;
wire n_n5005;
wire n_n5004;
wire n_n5000;
wire wire136;
wire wire393;
wire n_n4907;
wire n_n4913;
wire n_n4922;
wire n_n4934;
wire n_n2451;
wire n_n2462;
wire n_n2464;
wire wire31;
wire n_n4453;
wire n_n4420;
wire n_n4407;
wire n_n2455;
wire n_n2454;
wire n_n2472;
wire n_n2473;
wire wire234;
wire n_n4372;
wire n_n4373;
wire n_n4371;
wire n_n4431;
wire n_n4433;
wire n_n4430;
wire n_n4494;
wire n_n4491;
wire n_n4834;
wire n_n4835;
wire n_n4832;
wire n_n4909;
wire n_n4911;
wire n_n4903;
wire n_n4979;
wire n_n5049;
wire n_n5179;
wire n_n5239;
wire wire19;
wire n_n5240;
wire n_n5238;
wire n_n4514;
wire n_n4247;
wire n_n4646;
wire n_n4644;
wire n_n4651;
wire n_n4649;
wire wire311;
wire n_n4951;
wire n_n4952;
wire n_n4950;
wire n_n3803;
wire n_n4942;
wire n_n4943;
wire wire59;
wire n_n4945;
wire n_n4946;
wire n_n4949;
wire n_n2222;
wire n_n5244;
wire n_n5245;
wire wire318;
wire n_n2200;
wire n_n4450;
wire n_n4445;
wire n_n4444;
wire n_n4442;
wire n_n4441;
wire wire368;
wire n_n4470;
wire n_n4460;
wire n_n4473;
wire n_n4466;
wire n_n4895;
wire n_n4890;
wire wire260;
wire n_n2226;
wire n_n4850;
wire wire277;
wire wire295;
wire n_n2228;
wire n_n4881;
wire n_n4878;
wire n_n4880;
wire n_n4869;
wire n_n4877;
wire wire174;
wire n_n2178;
wire n_n5321;
wire n_n2274;
wire n_n5307;
wire n_n5326;
wire n_n5325;
wire n_n5332;
wire n_n5329;
wire wire117;
wire wire269;
wire n_n2179;
wire n_n4776;
wire n_n4774;
wire n_n4786;
wire wire131;
wire wire313;
wire n_n2162;
wire n_n4755;
wire n_n4759;
wire n_n4760;
wire n_n4758;
wire n_n2182;
wire n_n2183;
wire n_n2163;
wire n_n4963;
wire n_n4959;
wire n_n4960;
wire n_n4964;
wire n_n2177;
wire wire250;
wire n_n4817;
wire n_n4827;
wire n_n4816;
wire n_n5097;
wire n_n5019;
wire n_n4404;
wire n_n4413;
wire n_n4416;
wire n_n4523;
wire n_n4547;
wire n_n4539;
wire n_n4521;
wire n_n4544;
wire n_n4557;
wire n_n4560;
wire n_n4553;
wire n_n4800;
wire n_n2130;
wire n_n4803;
wire n_n4783;
wire n_n4812;
wire n_n4811;
wire n_n4781;
wire n_n2099;
wire n_n4361;
wire n_n4363;
wire n_n4359;
wire n_n4438;
wire n_n4439;
wire n_n4437;
wire n_n4825;
wire n_n4828;
wire n_n4824;
wire n_n4879;
wire n_n4937;
wire n_n4938;
wire n_n4936;
wire n_n5010;
wire n_n5037;
wire n_n1570;
wire n_n5043;
wire n_n5045;
wire n_n5302;
wire n_n5294;
wire n_n4894;
wire n_n4916;
wire n_n4930;
wire n_n4947;
wire wire96;
wire n_n5131;
wire n_n5137;
wire n_n5136;
wire n_n5200;
wire n_n5206;
wire n_n5146;
wire n_n5204;
wire n_n5191;
wire n_n5113;
wire n_n5081;
wire n_n5089;
wire n_n5124;
wire wire335;
wire n_n5258;
wire n_n5274;
wire n_n5232;
wire n_n5255;
wire n_n5267;
wire n_n5222;
wire n_n5212;
wire n_n4344;
wire n_n4345;
wire n_n4343;
wire n_n4392;
wire n_n4393;
wire n_n4391;
wire n_n4612;
wire n_n4611;
wire n_n4669;
wire n_n4673;
wire n_n4668;
wire n_n4734;
wire n_n4733;
wire n_n4792;
wire n_n4854;
wire n_n4855;
wire n_n4912;
wire n_n4908;
wire n_n4966;
wire n_n4968;
wire n_n5014;
wire n_n5015;
wire n_n5012;
wire n_n5067;
wire n_n5069;
wire n_n5066;
wire n_n5241;
wire n_n5243;
wire n_n5300;
wire n_n5299;
wire n_n4364;
wire n_n4362;
wire n_n3533;
wire n_n4366;
wire n_n4367;
wire n_n4365;
wire n_n1308;
wire n_n4770;
wire n_n4769;
wire n_n4767;
wire n_n4764;
wire n_n4905;
wire wire352;
wire n_n5046;
wire n_n5056;
wire n_n5057;
wire wire166;
wire wire292;
wire n_n4843;
wire n_n4845;
wire n_n4846;
wire n_n4848;
wire n_n3820;
wire n_n4384;
wire n_n4390;
wire n_n4374;
wire n_n4638;
wire n_n4633;
wire n_n5155;
wire n_n5161;
wire n_n509;
wire n_n522;
wire n_n536;
wire n_n473;
wire n_n524;
wire n_n4425;
wire n_n464;
wire n_n526;
wire n_n455;
wire n_n535;
wire n_n528;
wire n_n4482;
wire n_n4489;
wire n_n500;
wire n_n4504;
wire n_n4511;
wire n_n491;
wire n_n520;
wire n_n4526;
wire n_n4533;
wire n_n4554;
wire n_n4561;
wire n_n4568;
wire n_n4575;
wire n_n390;
wire n_n4590;
wire n_n530;
wire n_n4640;
wire n_n4647;
wire n_n482;
wire n_n4662;
wire n_n532;
wire n_n4690;
wire n_n534;
wire n_n325;
wire n_n4704;
wire n_n4711;
wire n_n518;
wire n_n4748;
wire n_n4777;
wire n_n4821;
wire n_n260;
wire n_n4901;
wire n_n195;
wire n_n4974;
wire n_n5003;
wire n_n5047;
wire n_n130;
wire n_n5098;
wire n_n5105;
wire n_n5120;
wire n_n5127;
wire n_n5186;
wire n_n5193;
wire n_n65;
wire n_n5251;
wire n_n5266;
wire n_n5273;
wire n_n4347;
wire n_n4397;
wire n_n4398;
wire n_n4396;
wire n_n4524;
wire n_n4522;
wire wire170;
wire n_n4246;
wire n_n4670;
wire n_n4732;
wire n_n4789;
wire n_n4906;
wire n_n4967;
wire n_n5086;
wire n_n5087;
wire n_n4589;
wire n_n4587;
wire n_n881;
wire n_n4594;
wire n_n4083;
wire n_n4639;
wire n_n4904;
wire n_n4319;
wire n_n4320;
wire n_n4451;
wire n_n4918;
wire n_n4919;
wire n_n4917;
wire n_n4985;
wire n_n4984;
wire n_n5031;
wire n_n5114;
wire n_n5116;
wire n_n5162;
wire n_n4582;
wire n_n4584;
wire n_n4586;
wire wire365;
wire n_n3348;
wire n_n4876;
wire wire461;
wire n_n3326;
wire n_n5327;
wire n_n2643;
wire n_n5323;
wire n_n5324;
wire n_n5322;
wire n_n4577;
wire n_n4576;
wire n_n4569;
wire n_n4574;
wire n_n4581;
wire n_n4572;
wire n_n4573;
wire n_n4579;
wire n_n3282;
wire n_n4538;
wire n_n4525;
wire n_n4531;
wire n_n3871;
wire wire202;
wire n_n3260;
wire n_n4629;
wire n_n4583;
wire n_n4842;
wire n_n4844;
wire n_n4839;
wire n_n5303;
wire n_n5182;
wire n_n5173;
wire n_n5165;
wire n_n5230;
wire n_n5166;
wire n_n5163;
wire n_n5214;
wire n_n4994;
wire n_n5002;
wire n_n5053;
wire n_n5033;
wire n_n5051;
wire n_n5006;
wire n_n4454;
wire n_n4518;
wire n_n4517;
wire n_n3152;
wire n_n4725;
wire n_n4726;
wire n_n4861;
wire n_n5039;
wire n_n5103;
wire n_n5104;
wire n_n5102;
wire n_n4395;
wire n_n2638;
wire wire425;
wire n_n2560;
wire n_n4426;
wire n_n2635;
wire wire37;
wire n_n2559;
wire n_n4315;
wire n_n4312;
wire n_n4360;
wire n_n4487;
wire n_n4483;
wire n_n4840;
wire n_n4837;
wire n_n4899;
wire n_n4986;
wire n_n5044;
wire n_n5115;
wire n_n5175;
wire n_n5177;
wire n_n5311;
wire n_n4798;
wire n_n4804;
wire n_n4794;
wire n_n4795;
wire n_n4793;
wire n_n4796;
wire n_n4797;
wire n_n4801;
wire n_n4933;
wire n_n4935;
wire wire249;
wire n_n2223;
wire wire289;
wire n_n4497;
wire wire65;
wire wire66;
wire n_n4478;
wire n_n4254;
wire wire70;
wire wire184;
wire n_n2258;
wire wire388;
wire n_n2230;
wire wire176;
wire n_n2229;
wire n_n4822;
wire n_n4823;
wire n_n4806;
wire n_n4820;
wire n_n4818;
wire n_n4810;
wire wire186;
wire n_n2263;
wire n_n2190;
wire n_n2446;
wire n_n4336;
wire n_n2443;
wire n_n2445;
wire wire171;
wire wire198;
wire wire283;
wire n_n4379;
wire n_n2435;
wire wire54;
wire wire282;
wire wire423;
wire n_n4503;
wire n_n4502;
wire n_n4500;
wire n_n4546;
wire n_n4555;
wire wire212;
wire wire213;
wire n_n4656;
wire n_n4659;
wire n_n5106;
wire n_n4341;
wire n_n5117;
wire n_n5223;
wire n_n5328;
wire n_n5254;
wire n_n5249;
wire n_n5233;
wire n_n5236;
wire n_n5262;
wire n_n5278;
wire wire449;
wire n_n2083;
wire n_n4375;
wire n_n4436;
wire n_n4833;
wire n_n4875;
wire n_n4940;
wire n_n4939;
wire n_n4729;
wire n_n4728;
wire wire373;
wire wire374;
wire n_n5132;
wire n_n5128;
wire n_n5016;
wire n_n4129;
wire n_n5306;
wire n_n3019;
wire n_n5009;
wire n_n5335;
wire n_n4562;
wire n_n4506;
wire n_n4492;
wire n_n1338;
wire n_n4496;
wire n_n4535;
wire n_n1326;
wire n_n1336;
wire n_n4788;
wire n_n1325;
wire n_n4342;
wire n_n4608;
wire n_n4610;
wire n_n4606;
wire n_n4675;
wire n_n4676;
wire n_n4674;
wire n_n4730;
wire n_n4802;
wire n_n4851;
wire n_n4852;
wire n_n4914;
wire n_n4962;
wire n_n4956;
wire n_n5020;
wire n_n5064;
wire n_n5189;
wire n_n5190;
wire n_n5188;
wire n_n4352;
wire n_n4351;
wire n_n4356;
wire wire67;
wire n_n1120;
wire n_n4507;
wire n_n4509;
wire n_n4508;
wire wire129;
wire wire308;
wire n_n4622;
wire n_n4621;
wire wire75;
wire n_n3861;
wire n_n5073;
wire n_n5074;
wire n_n5072;
wire n_n4152;
wire n_n4931;
wire wire180;
wire wire382;
wire n_n4978;
wire n_n4980;
wire n_n4897;
wire n_n1077;
wire wire264;
wire n_n4349;
wire n_n4350;
wire n_n4348;
wire n_n1002;
wire n_n5172;
wire n_n4580;
wire n_n4357;
wire n_n4419;
wire n_n4605;
wire n_n4655;
wire n_n4661;
wire n_n4683;
wire n_n4689;
wire n_n4697;
wire n_n4703;
wire n_n4712;
wire n_n4718;
wire n_n4763;
wire n_n4778;
wire n_n4886;
wire n_n4915;
wire n_n4989;
wire n_n5011;
wire n_n5061;
wire n_n5070;
wire n_n5076;
wire n_n5135;
wire n_n5157;
wire n_n5201;
wire n_n5207;
wire n_n5237;
wire n_n5252;
wire n_n4353;
wire n_n4456;
wire n_n4458;
wire n_n4671;
wire n_n4747;
wire n_n4772;
wire n_n4773;
wire n_n4771;
wire n_n4205;
wire n_n5023;
wire n_n5024;
wire n_n5082;
wire n_n5084;
wire n_n5275;
wire n_n5276;
wire n_n4600;
wire wire45;
wire n_n4204;
wire n_n4010;
wire n_n4009;
wire n_n3990;
wire n_n4753;
wire n_n4752;
wire n_n4013;
wire wire47;
wire n_n3992;
wire n_n4457;
wire n_n5075;
wire n_n5079;
wire n_n5088;
wire n_n5078;
wire n_n5083;
wire wire123;
wire wire122;
wire wire232;
wire n_n5063;
wire n_n5058;
wire wire160;
wire n_n3558;
wire n_n3557;
wire n_n4409;
wire n_n4399;
wire n_n4370;
wire n_n3548;
wire n_n4505;
wire n_n5095;
wire n_n5158;
wire n_n5154;
wire n_n4775;
wire n_n4780;
wire n_n3469;
wire n_n5013;
wire n_n5150;
wire n_n5147;
wire wire76;
wire wire196;
wire wire57;
wire wire251;
wire n_n4948;
wire n_n4957;
wire n_n4971;
wire wire342;
wire n_n4488;
wire n_n4471;
wire n_n4490;
wire n_n901;
wire n_n3358;
wire n_n3285;
wire n_n4423;
wire n_n4421;
wire wire84;
wire wire470;
wire n_n4635;
wire n_n4630;
wire n_n5065;
wire n_n5287;
wire n_n5281;
wire n_n5268;
wire n_n5261;
wire n_n3194;
wire n_n4331;
wire n_n4332;
wire n_n4329;
wire n_n4448;
wire n_n4449;
wire n_n4447;
wire n_n4870;
wire n_n5029;
wire n_n3162;
wire n_n4472;
wire n_n4469;
wire n_n4477;
wire n_n4475;
wire n_n4479;
wire n_n4474;
wire n_n3001;
wire wire465;
wire n_n4620;
wire n_n5001;
wire n_n2548;
wire n_n4867;
wire n_n4866;
wire n_n2597;
wire n_n4863;
wire n_n2727;
wire n_n2549;
wire n_n4965;
wire wire228;
wire n_n2551;
wire wire315;
wire n_n4321;
wire n_n4417;
wire n_n4415;
wire n_n4972;
wire n_n5118;
wire n_n5119;
wire n_n5229;
wire n_n5228;
wire n_n5295;
wire n_n4540;
wire n_n4536;
wire n_n4532;
wire n_n4541;
wire wire416;
wire n_n4681;
wire n_n4679;
wire n_n4677;
wire n_n4678;
wire wire81;
wire n_n2242;
wire wire414;
wire wire345;
wire wire164;
wire n_n4465;
wire n_n4443;
wire n_n5121;
wire n_n5122;
wire n_n4486;
wire n_n4484;
wire wire199;
wire n_n4865;
wire n_n4893;
wire wire154;
wire n_n2095;
wire n_n5168;
wire n_n2091;
wire n_n4973;
wire n_n2084;
wire n_n4378;
wire n_n4377;
wire n_n4710;
wire n_n4709;
wire n_n4765;
wire n_n4603;
wire n_n4604;
wire n_n2037;
wire n_n4588;
wire n_n4595;
wire n_n1877;
wire n_n1450;
wire n_n5152;
wire n_n5149;
wire wire195;
wire wire358;
wire wire406;
wire n_n5288;
wire n_n4743;
wire n_n4751;
wire n_n1333;
wire n_n4386;
wire n_n4435;
wire n_n4626;
wire n_n4627;
wire n_n4625;
wire n_n4660;
wire n_n4719;
wire n_n4717;
wire n_n4954;
wire n_n4955;
wire n_n5133;
wire n_n5138;
wire n_n5139;
wire n_n5309;
wire n_n5308;
wire n_n1128;
wire n_n4387;
wire wire420;
wire n_n4619;
wire wire179;
wire n_n4750;
wire n_n4745;
wire n_n4736;
wire wire293;
wire wire457;
wire n_n5159;
wire n_n5160;
wire wire287;
wire n_n5169;
wire wire33;
wire wire107;
wire wire113;
wire wire254;
wire n_n4658;
wire n_n5108;
wire n_n4510;
wire n_n4355;
wire n_n4424;
wire n_n4498;
wire n_n4591;
wire n_n4663;
wire n_n4698;
wire n_n4705;
wire n_n4805;
wire n_n4841;
wire n_n4944;
wire n_n5068;
wire n_n5187;
wire n_n5199;
wire n_n5260;
wire n_n5272;
wire n_n4405;
wire n_n4406;
wire n_n4462;
wire n_n4501;
wire n_n4684;
wire n_n4222;
wire n_n4741;
wire n_n4740;
wire n_n4819;
wire n_n5077;
wire n_n5221;
wire n_n5220;
wire n_n834;
wire n_n5134;
wire n_n5125;
wire wire336;
wire n_n3988;
wire n_n5290;
wire n_n5291;
wire n_n5292;
wire n_n4026;
wire n_n3998;
wire wire441;
wire n_n3987;
wire n_n4410;
wire n_n4652;
wire n_n4650;
wire n_n3681;
wire wire97;
wire n_n3639;
wire wire159;
wire n_n5226;
wire n_n5218;
wire wire435;
wire n_n5153;
wire n_n5021;
wire n_n4654;
wire wire140;
wire wire391;
wire n_n4665;
wire wire72;
wire wire418;
wire wire248;
wire n_n4368;
wire n_n4394;
wire n_n3363;
wire n_n3362;
wire n_n3287;
wire n_n3369;
wire n_n3370;
wire wire156;
wire n_n3262;
wire n_n4891;
wire n_n4896;
wire n_n4428;
wire wire403;
wire n_n4499;
wire n_n4545;
wire wire471;
wire n_n4326;
wire n_n4328;
wire n_n4376;
wire n_n3176;
wire n_n4585;
wire n_n4873;
wire n_n4932;
wire n_n4592;
wire n_n5052;
wire n_n2956;
wire n_n5235;
wire n_n5234;
wire n_n5286;
wire n_n5285;
wire n_n1764;
wire n_n3810;
wire n_n2304;
wire n_n5256;
wire n_n5253;
wire n_n1139;
wire n_n4408;
wire n_n4414;
wire wire215;
wire n_n2169;
wire n_n5170;
wire wire168;
wire n_n2159;
wire n_n2214;
wire n_n2168;
wire n_n5333;
wire n_n4429;
wire n_n4813;
wire n_n4815;
wire n_n4838;
wire wire85;
wire n_n2096;
wire n_n4715;
wire n_n4714;
wire n_n5225;
wire n_n5224;
wire n_n1530;
wire wire437;
wire n_n5279;
wire n_n5277;
wire n_n4708;
wire n_n4706;
wire wire366;
wire n_n4427;
wire n_n4716;
wire n_n4807;
wire n_n1162;
wire n_n5312;
wire n_n5313;
wire n_n4596;
wire wire256;
wire n_n1059;
wire wire28;
wire n_n4672;
wire n_n4468;
wire n_n4418;
wire n_n4446;
wire n_n4688;
wire n_n4836;
wire n_n4871;
wire n_n4961;
wire n_n5140;
wire n_n5194;
wire n_n5259;
wire n_n5271;
wire n_n4537;
wire n_n4614;
wire n_n4058;
wire n_n3993;
wire n_n3995;
wire wire55;
wire n_n3986;
wire n_n4707;
wire n_n4701;
wire n_n4643;
wire n_n4642;
wire n_n3716;
wire n_n3650;
wire n_n4556;
wire n_n4550;
wire n_n3870;
wire wire91;
wire wire430;
wire n_n4609;
wire n_n3718;
wire n_n3629;
wire n_n4358;
wire n_n4493;
wire n_n5148;
wire n_n3461;
wire n_n3329;
wire n_n5126;
wire n_n3307;
wire n_n3277;
wire n_n4808;
wire n_n3330;
wire n_n3275;
wire n_n2710;
wire n_n3274;
wire wire58;
wire n_n3257;
wire wire456;
wire n_n4799;
wire n_n3202;
wire n_n3204;
wire n_n4685;
wire n_n4520;
wire n_n4884;
wire n_n5008;
wire n_n4623;
wire wire304;
wire n_n2601;
wire n_n2602;
wire wire433;
wire n_n5242;
wire wire320;
wire n_n5264;
wire n_n5270;
wire wire77;
wire wire334;
wire wire149;
wire wire267;
wire n_n2564;
wire n_n2566;
wire wire218;
wire wire385;
wire wire399;
wire wire125;
wire n_n2196;
wire wire44;
wire wire332;
wire wire90;
wire wire144;
wire wire239;
wire n_n4335;
wire n_n4411;
wire n_n4279;
wire n_n5219;
wire n_n1456;
wire n_n1521;
wire n_n4528;
wire n_n4529;
wire n_n5319;
wire wire328;
wire n_n4542;
wire wire201;
wire n_n4543;
wire n_n4549;
wire n_n4551;
wire n_n4691;
wire n_n3849;
wire n_n4692;
wire n_n1093;
wire wire299;
wire n_n1050;
wire n_n5269;
wire n_n5257;
wire wire62;
wire wire92;
wire wire409;
wire n_n1049;
wire n_n1048;
wire wire63;
wire wire200;
wire n_n1017;
wire n_n1045;
wire n_n1900;
wire wire115;
wire wire175;
wire n_n1007;
wire n_n4476;
wire n_n4686;
wire n_n4354;
wire n_n4889;
wire n_n5196;
wire n_n5203;
wire n_n5210;
wire n_n5217;
wire n_n3996;
wire n_n4929;
wire n_n4766;
wire wire447;
wire n_n1592;
wire n_n4742;
wire n_n4527;
wire n_n4713;
wire n_n3708;
wire n_n3648;
wire n_n4657;
wire n_n3711;
wire n_n3649;
wire n_n3653;
wire n_n3655;
wire n_n5090;
wire n_n5144;
wire n_n5143;
wire n_n2685;
wire n_n3308;
wire n_n5007;
wire wire211;
wire n_n3251;
wire n_n4953;
wire n_n3201;
wire n_n4334;
wire wire158;
wire wire380;
wire n_n4874;
wire wire49;
wire wire87;
wire wire182;
wire n_n5215;
wire wire220;
wire wire384;
wire wire454;
wire n_n4534;
wire n_n2558;
wire n_n2626;
wire n_n2533;
wire wire82;
wire wire224;
wire n_n5248;
wire n_n4412;
wire n_n2651;
wire n_n5195;
wire n_n5197;
wire n_n2291;
wire wire451;
wire n_n4316;
wire n_n4313;
wire n_n4723;
wire n_n4722;
wire n_n4892;
wire n_n5213;
wire n_n5209;
wire n_n1532;
wire wire288;
wire n_n5247;
wire wire446;
wire n_n1435;
wire n_n1103;
wire wire181;
wire wire452;
wire n_n5208;
wire n_n5211;
wire n_n1038;
wire wire79;
wire n_n3875;
wire n_n1040;
wire n_n4322;
wire n_n1041;
wire n_n4695;
wire n_n4826;
wire n_n5151;
wire n_n4197;
wire n_n4883;
wire wire330;
wire n_n5071;
wire n_n1167;
wire n_n3253;
wire n_n2997;
wire n_n5198;
wire n_n3037;
wire wire183;
wire wire453;
wire n_n5246;
wire n_n5176;
wire wire80;
wire wire157;
wire n_n2579;
wire wire88;
wire n_n2541;
wire wire297;
wire wire394;
wire n_n2528;
wire n_n2470;
wire n_n2467;
wire wire361;
wire wire378;
wire wire341;
wire wire362;
wire wire203;
wire wire205;
wire wire438;
wire n_n4699;
wire n_n4687;
wire wire340;
wire n_n5250;
wire n_n5205;
wire n_n801;
wire n_n1454;
wire n_n1436;
wire n_n5330;
wire n_n5331;
wire wire421;
wire wire432;
wire n_n1985;
wire n_n3815;
wire wire253;
wire n_n1061;
wire n_n1022;
wire wire104;
wire n_n1009;
wire n_n4323;
wire wire128;
wire n_n910;
wire n_n4631;
wire n_n559;
wire n_n4761;
wire n_n4680;
wire wire343;
wire wire379;
wire n_n2996;
wire wire431;
wire n_n2670;
wire n_n4402;
wire wire455;
wire wire238;
wire wire276;
wire n_n4702;
wire n_n1455;
wire n_n4599;
wire wire364;
wire n_n5283;
wire wire333;
wire n_n4632;
wire wire139;
wire n_n953;
wire wire99;
wire n_n942;
wire n_n725;
wire wire52;
wire wire150;
wire n_n4645;
wire wire310;
wire n_n4696;
wire n_n4762;
wire n_n5315;
wire n_n1952;
wire wire363;
wire wire407;
wire n_n4056;
wire wire42;
wire n_n814;
wire wire141;
wire wire317;
wire n_n5192;
wire wire106;
wire wire375;
wire n_n4558;
wire wire417;
wire wire27;
wire n_n1472;
wire n_n763;
wire wire286;
wire n_n667;
wire n_n761;
wire n_n635;
wire n_n777;
wire n_n3772;
wire n_n637;
wire n_n4552;
wire n_n4559;
wire n_n5227;
wire n_n5304;
wire n_n4694;
wire n_n4700;
wire n_n4219;
wire wire221;
wire n_n4075;
wire wire30;
wire wire173;
wire wire243;
wire n_n4065;
wire wire390;
wire n_n3926;
wire n_n3924;
wire n_n3923;
wire n_n3928;
wire n_n3124;
wire n_n2378;
wire n_n4693;
wire n_n3051;
wire n_n3007;
wire n_n3003;
wire n_n2604;
wire n_n4910;
wire wire190;
wire n_n1501;
wire n_n1426;
wire n_n1409;
wire n_n1448;
wire n_n1408;
wire wire347;
wire n_n5280;
wire n_n5080;
wire n_n680;
wire wire209;
wire n_n639;
wire n_n625;
wire n_n4721;
wire n_n4548;
wire n_n4099;
wire n_n4021;
wire n_n789;
wire wire445;
wire wire422;
wire wire442;
wire wire386;
wire n_n3879;
wire n_n2058;
wire wire324;
wire wire305;
wire wire291;
wire n_n1111;
wire n_n554;
wire wire279;
wire n_n4016;
wire wire401;
wire n_n3560;
wire wire434;
wire n_n3009;
wire n_n4330;
wire n_n3889;
wire n_n2238;
wire n_n4872;
wire n_n1677;
wire n_n1496;
wire n_n1467;
wire n_n1415;
wire n_n1091;
wire n_n4030;
wire wire124;
wire n_n1402;
wire wire204;
wire n_n956;
wire n_n941;
wire n_n937;
wire n_n4031;
wire wire600;
wire n_n1418;
wire n_n5289;
wire wire255;
wire n_n1712;
wire n_n1730;
wire n_n1729;
wire n_n1711;
wire n_n5282;
wire wire225;
wire n_n5298;
wire n_n3931;
wire n_n3929;
wire wire261;
wire n_n3694;
wire n_n2761;
wire n_n2982;
wire wire466;
wire n_n2953;
wire n_n2955;
wire n_n2915;
wire wire265;
wire n_n2902;
wire n_n2839;
wire n_n2630;
wire n_n1840;
wire n_n1801;
wire n_n1837;
wire n_n1800;
wire n_n1842;
wire n_n1725;
wire n_n707;
wire n_n691;
wire n_n632;
wire n_n646;
wire n_n627;
wire n_n856;
wire n_n648;
wire n_n628;
wire n_n621;
wire n_n1760;
wire n_n2841;
wire wire53;
wire n_n1852;
wire n_n1805;
wire n_n1789;
wire wire444;
wire n_n1724;
wire n_n1478;
wire n_n662;
wire n_n661;
wire n_n620;
wire n_n3736;
wire n_n2837;
wire n_n2611;
wire n_n1894;
wire n_n1862;
wire n_n1808;
wire n_n1856;
wire n_n1790;
wire n_n1727;
wire n_n1722;
wire n_n1721;
wire n_n722;
wire n_n653;
wire n_n630;
wire n_n3664;
wire n_n3012;
wire n_n2934;
wire n_n2985;
wire n_n2925;
wire n_n2824;
wire n_n2835;
wire n_n1892;
wire n_n1818;
wire n_n1865;
wire n_n1476;
wire n_n732;
wire n_n656;
wire n_n631;
wire n_n651;
wire n_n629;
wire n_n3561;
wire n_n2939;
wire n_n2832;
wire n_n2834;
wire n_n1032;
wire n_n948;
wire n_n700;
wire n_n3689;
wire n_n3724;
wire n_n949;
wire n_n715;
wire n_n3670;
wire n_n2937;
wire n_n2929;
wire n_n1718;
wire n_n1717;
wire n_n951;
wire n_n1824;
wire n_n1826;
wire n_n1885;
wire n_n1886;
wire n_n1879;
wire n_n1813;
wire n_n1812;
wire n_n1012;
wire n_n3729;
wire n_n3699;
wire n_n3701;
wire n_n3645;
wire n_n1872;
wire n_n1828;
wire n_n1797;
wire n_n3646;
wire n_n3635;
wire n_n3641;
wire n_n2905;
wire wire266;
wire wire606;
wire wire617;
wire wire636;
wire wire656;
wire wire664;
wire wire669;
wire wire671;
wire wire675;
wire wire677;
wire wire679;
wire wire683;
wire wire686;
wire wire693;
wire wire695;
wire wire706;
wire wire724;
wire wire732;
wire wire735;
wire wire743;
wire wire745;
wire wire755;
wire wire761;
wire wire765;
wire wire767;
wire wire771;
wire wire772;
wire wire773;
wire wire775;
wire wire783;
wire wire787;
wire wire789;
wire wire791;
wire wire11482;
wire wire11483;
wire wire11488;
wire wire11489;
wire wire11491;
wire wire11492;
wire wire11495;
wire wire11496;
wire wire11497;
wire wire11498;
wire wire11501;
wire wire11502;
wire wire11505;
wire wire11507;
wire wire11508;
wire wire11511;
wire wire11512;
wire wire11513;
wire wire11515;
wire wire11516;
wire wire11518;
wire wire11520;
wire wire11521;
wire wire11522;
wire wire11523;
wire wire11524;
wire wire11527;
wire wire11529;
wire wire11530;
wire wire11532;
wire wire11534;
wire wire11535;
wire wire11536;
wire wire11537;
wire wire11539;
wire wire11541;
wire wire11543;
wire wire11547;
wire wire11548;
wire wire11549;
wire wire11553;
wire wire11554;
wire wire11555;
wire wire11558;
wire wire11559;
wire wire11560;
wire wire11562;
wire wire11563;
wire wire11564;
wire wire11566;
wire wire11567;
wire wire11568;
wire wire11570;
wire wire11571;
wire wire11574;
wire wire11575;
wire wire11578;
wire wire11579;
wire wire11581;
wire wire11582;
wire wire11583;
wire wire11584;
wire wire11585;
wire wire11586;
wire wire11587;
wire wire11588;
wire wire11589;
wire wire11591;
wire wire11592;
wire wire11593;
wire wire11597;
wire wire11598;
wire wire11599;
wire wire11600;
wire wire11601;
wire wire11602;
wire wire11605;
wire wire11607;
wire wire11610;
wire wire11611;
wire wire11613;
wire wire11614;
wire wire11618;
wire wire11620;
wire wire11625;
wire wire11626;
wire wire11628;
wire wire11630;
wire wire11631;
wire wire11633;
wire wire11634;
wire wire11638;
wire wire11641;
wire wire11642;
wire wire11646;
wire wire11647;
wire wire11653;
wire wire11654;
wire wire11655;
wire wire11658;
wire wire11660;
wire wire11661;
wire wire11666;
wire wire11667;
wire wire11671;
wire wire11675;
wire wire11676;
wire wire11677;
wire wire11680;
wire wire11681;
wire wire11687;
wire wire11688;
wire wire11690;
wire wire11693;
wire wire11694;
wire wire11698;
wire wire11699;
wire wire11703;
wire wire11705;
wire wire11706;
wire wire11707;
wire wire11710;
wire wire11712;
wire wire11713;
wire wire11715;
wire wire11718;
wire wire11719;
wire wire11725;
wire wire11726;
wire wire11731;
wire wire11732;
wire wire11734;
wire wire11735;
wire wire11738;
wire wire11739;
wire wire11741;
wire wire11743;
wire wire11745;
wire wire11748;
wire wire11751;
wire wire11752;
wire wire11753;
wire wire11754;
wire wire11756;
wire wire11757;
wire wire11759;
wire wire11761;
wire wire11762;
wire wire11765;
wire wire11766;
wire wire11767;
wire wire11768;
wire wire11769;
wire wire11772;
wire wire11773;
wire wire11774;
wire wire11776;
wire wire11777;
wire wire11778;
wire wire11781;
wire wire11782;
wire wire11783;
wire wire11785;
wire wire11786;
wire wire11788;
wire wire11790;
wire wire11791;
wire wire11795;
wire wire11796;
wire wire11797;
wire wire11801;
wire wire11802;
wire wire11803;
wire wire11804;
wire wire11805;
wire wire11807;
wire wire11808;
wire wire11809;
wire wire11810;
wire wire11811;
wire wire11812;
wire wire11814;
wire wire11815;
wire wire11816;
wire wire11818;
wire wire11823;
wire wire11824;
wire wire11825;
wire wire11826;
wire wire11829;
wire wire11830;
wire wire11832;
wire wire11833;
wire wire11834;
wire wire11836;
wire wire11837;
wire wire11839;
wire wire11841;
wire wire11842;
wire wire11846;
wire wire11847;
wire wire11848;
wire wire11851;
wire wire11852;
wire wire11855;
wire wire11856;
wire wire11859;
wire wire11862;
wire wire11866;
wire wire11867;
wire wire11870;
wire wire11873;
wire wire11874;
wire wire11877;
wire wire11880;
wire wire11881;
wire wire11882;
wire wire11884;
wire wire11886;
wire wire11888;
wire wire11889;
wire wire11891;
wire wire11893;
wire wire11894;
wire wire11899;
wire wire11900;
wire wire11902;
wire wire11906;
wire wire11907;
wire wire11908;
wire wire11909;
wire wire11912;
wire wire11914;
wire wire11916;
wire wire11917;
wire wire11918;
wire wire11921;
wire wire11923;
wire wire11924;
wire wire11927;
wire wire11928;
wire wire11929;
wire wire11930;
wire wire11933;
wire wire11939;
wire wire11940;
wire wire11944;
wire wire11946;
wire wire11947;
wire wire11951;
wire wire11952;
wire wire11955;
wire wire11959;
wire wire11960;
wire wire11962;
wire wire11964;
wire wire11967;
wire wire11968;
wire wire11970;
wire wire11971;
wire wire11972;
wire wire11973;
wire wire11975;
wire wire11977;
wire wire11978;
wire wire11981;
wire wire11982;
wire wire11986;
wire wire11987;
wire wire11992;
wire wire11993;
wire wire11994;
wire wire11995;
wire wire11996;
wire wire11997;
wire wire11999;
wire wire12001;
wire wire12003;
wire wire12004;
wire wire12007;
wire wire12009;
wire wire12014;
wire wire12015;
wire wire12018;
wire wire12020;
wire wire12022;
wire wire12023;
wire wire12024;
wire wire12027;
wire wire12028;
wire wire12033;
wire wire12034;
wire wire12036;
wire wire12037;
wire wire12040;
wire wire12041;
wire wire12047;
wire wire12048;
wire wire12053;
wire wire12054;
wire wire12058;
wire wire12060;
wire wire12061;
wire wire12062;
wire wire12067;
wire wire12068;
wire wire12074;
wire wire12075;
wire wire12080;
wire wire12081;
wire wire12083;
wire wire12089;
wire wire12090;
wire wire12091;
wire wire12092;
wire wire12093;
wire wire12096;
wire wire12097;
wire wire12099;
wire wire12101;
wire wire12102;
wire wire12106;
wire wire12108;
wire wire12109;
wire wire12110;
wire wire12111;
wire wire12113;
wire wire12114;
wire wire12115;
wire wire12117;
wire wire12118;
wire wire12120;
wire wire12122;
wire wire12123;
wire wire12126;
wire wire12128;
wire wire12129;
wire wire12131;
wire wire12134;
wire wire12136;
wire wire12137;
wire wire12141;
wire wire12142;
wire wire12146;
wire wire12147;
wire wire12149;
wire wire12150;
wire wire12152;
wire wire12156;
wire wire12159;
wire wire12162;
wire wire12164;
wire wire12165;
wire wire12166;
wire wire12167;
wire wire12168;
wire wire12169;
wire wire12170;
wire wire12171;
wire wire12172;
wire wire12175;
wire wire12176;
wire wire12177;
wire wire12179;
wire wire12181;
wire wire12182;
wire wire12183;
wire wire12186;
wire wire12187;
wire wire12188;
wire wire12191;
wire wire12192;
wire wire12196;
wire wire12197;
wire wire12200;
wire wire12202;
wire wire12204;
wire wire12205;
wire wire12207;
wire wire12208;
wire wire12210;
wire wire12213;
wire wire12214;
wire wire12217;
wire wire12218;
wire wire12219;
wire wire12220;
wire wire12223;
wire wire12224;
wire wire12225;
wire wire12226;
wire wire12230;
wire wire12231;
wire wire12232;
wire wire12234;
wire wire12235;
wire wire12239;
wire wire12240;
wire wire12243;
wire wire12245;
wire wire12247;
wire wire12252;
wire wire12253;
wire wire12255;
wire wire12256;
wire wire12257;
wire wire12261;
wire wire12262;
wire wire12265;
wire wire12266;
wire wire12268;
wire wire12269;
wire wire12271;
wire wire12272;
wire wire12276;
wire wire12277;
wire wire12278;
wire wire12282;
wire wire12283;
wire wire12285;
wire wire12287;
wire wire12288;
wire wire12290;
wire wire12291;
wire wire12292;
wire wire12293;
wire wire12296;
wire wire12297;
wire wire12299;
wire wire12300;
wire wire12301;
wire wire12304;
wire wire12305;
wire wire12306;
wire wire12309;
wire wire12310;
wire wire12315;
wire wire12316;
wire wire12317;
wire wire12318;
wire wire12319;
wire wire12323;
wire wire12324;
wire wire12326;
wire wire12327;
wire wire12328;
wire wire12332;
wire wire12333;
wire wire12335;
wire wire12337;
wire wire12338;
wire wire12340;
wire wire12342;
wire wire12344;
wire wire12345;
wire wire12349;
wire wire12352;
wire wire12353;
wire wire12355;
wire wire12356;
wire wire12358;
wire wire12359;
wire wire12361;
wire wire12363;
wire wire12364;
wire wire12366;
wire wire12368;
wire wire12369;
wire wire12371;
wire wire12372;
wire wire12374;
wire wire12375;
wire wire12376;
wire wire12380;
wire wire12381;
wire wire12382;
wire wire12384;
wire wire12386;
wire wire12387;
wire wire12389;
wire wire12391;
wire wire12392;
wire wire12393;
wire wire12395;
wire wire12398;
wire wire12399;
wire wire12400;
wire wire12401;
wire wire12403;
wire wire12404;
wire wire12408;
wire wire12409;
wire wire12413;
wire wire12414;
wire wire12416;
wire wire12420;
wire wire12421;
wire wire12422;
wire wire12425;
wire wire12426;
wire wire12428;
wire wire12429;
wire wire12431;
wire wire12432;
wire wire12434;
wire wire12435;
wire wire12436;
wire wire12439;
wire wire12440;
wire wire12442;
wire wire12445;
wire wire12446;
wire wire12447;
wire wire12448;
wire wire12449;
wire wire12451;
wire wire12453;
wire wire12455;
wire wire12456;
wire wire12458;
wire wire12459;
wire wire12461;
wire wire12464;
wire wire12465;
wire wire12467;
wire wire12469;
wire wire12471;
wire wire12472;
wire wire12475;
wire wire12476;
wire wire12478;
wire wire12479;
wire wire12480;
wire wire12481;
wire wire12485;
wire wire12486;
wire wire12488;
wire wire12489;
wire wire12490;
wire wire12492;
wire wire12493;
wire wire12497;
wire wire12498;
wire wire12499;
wire wire12500;
wire wire12501;
wire wire12502;
wire wire12503;
wire wire12507;
wire wire12508;
wire wire12510;
wire wire12514;
wire wire12515;
wire wire12517;
wire wire12518;
wire wire12519;
wire wire12520;
wire wire12521;
wire wire12524;
wire wire12525;
wire wire12529;
wire wire12530;
wire wire12531;
wire wire12534;
wire wire12535;
wire wire12539;
wire wire12540;
wire wire12541;
wire wire12543;
wire wire12544;
wire wire12545;
wire wire12546;
wire wire12547;
wire wire12551;
wire wire12552;
wire wire12554;
wire wire12555;
wire wire12556;
wire wire12557;
wire wire12559;
wire wire12560;
wire wire12561;
wire wire12564;
wire wire12566;
wire wire12567;
wire wire12568;
wire wire12569;
wire wire12570;
wire wire12572;
wire wire12573;
wire wire12574;
wire wire12576;
wire wire12577;
wire wire12578;
wire wire12579;
wire wire12580;
wire wire12582;
wire wire12583;
wire wire12585;
wire wire12586;
wire wire12588;
wire wire12589;
wire wire12595;
wire wire12596;
wire wire12600;
wire wire12601;
wire wire12602;
wire wire12607;
wire wire12608;
wire wire12609;
wire wire12613;
wire wire12614;
wire wire12615;
wire wire12620;
wire wire12621;
wire wire12626;
wire wire12627;
wire wire12629;
wire wire12630;
wire wire12634;
wire wire12635;
wire wire12638;
wire wire12640;
wire wire12641;
wire wire12642;
wire wire12643;
wire wire12648;
wire wire12649;
wire wire12650;
wire wire12651;
wire wire12653;
wire wire12656;
wire wire12657;
wire wire12658;
wire wire12659;
wire wire12663;
wire wire12664;
wire wire12669;
wire wire12670;
wire wire12672;
wire wire12673;
wire wire12675;
wire wire12678;
wire wire12679;
wire wire12682;
wire wire12683;
wire wire12688;
wire wire12689;
wire wire12691;
wire wire12693;
wire wire12694;
wire wire12699;
wire wire12700;
wire wire12706;
wire wire12707;
wire wire12710;
wire wire12713;
wire wire12714;
wire wire12718;
wire wire12722;
wire wire12724;
wire wire12725;
wire wire12729;
wire wire12730;
wire wire12732;
wire wire12735;
wire wire12736;
wire wire12740;
wire wire12742;
wire wire12743;
wire wire12744;
wire wire12745;
wire wire12747;
wire wire12748;
wire wire12749;
wire wire12752;
wire wire12753;
wire wire12756;
wire wire12757;
wire wire12759;
wire wire12760;
wire wire12762;
wire wire12763;
wire wire12766;
wire wire12767;
wire wire12769;
wire wire12770;
wire wire12771;
wire wire12774;
wire wire12775;
wire wire12778;
wire wire12783;
wire wire12784;
wire wire12787;
wire wire12788;
wire wire12790;
wire wire12791;
wire wire12792;
wire wire12794;
wire wire12796;
wire wire12799;
wire wire12800;
wire wire12801;
wire wire12802;
wire wire12804;
wire wire12805;
wire wire12810;
wire wire12811;
wire wire12813;
wire wire12814;
wire wire12815;
wire wire12819;
wire wire12820;
wire wire12822;
wire wire12826;
wire wire12827;
wire wire12831;
wire wire12832;
wire wire12833;
wire wire12834;
wire wire12835;
wire wire12838;
wire wire12839;
wire wire12841;
wire wire12843;
wire wire12844;
wire wire12845;
wire wire12848;
wire wire12849;
wire wire12852;
wire wire12853;
wire wire12854;
wire wire12857;
wire wire12858;
wire wire12859;
wire wire12862;
wire wire12863;
wire wire12865;
wire wire12866;
wire wire12871;
wire wire12872;
wire wire12874;
wire wire12875;
wire wire12876;
wire wire12877;
wire wire12881;
wire wire12883;
wire wire12884;
wire wire12888;
wire wire12889;
wire wire12892;
wire wire12893;
wire wire12894;
wire wire12898;
wire wire12902;
wire wire12904;
wire wire12907;
wire wire12908;
wire wire12909;
wire wire12914;
wire wire12915;
wire wire12917;
wire wire12921;
wire wire12922;
wire wire12924;
wire wire12925;
wire wire12926;
wire wire12929;
wire wire12930;
wire wire12931;
wire wire12933;
wire wire12934;
wire wire12935;
wire wire12936;
wire wire12938;
wire wire12939;
wire wire12940;
wire wire12941;
wire wire12943;
wire wire12944;
wire wire12946;
wire wire12947;
wire wire12949;
wire wire12952;
wire wire12953;
wire wire12954;
wire wire12958;
wire wire12960;
wire wire12961;
wire wire12962;
wire wire12963;
wire wire12966;
wire wire12967;
wire wire12969;
wire wire12970;
wire wire12971;
wire wire12972;
wire wire12975;
wire wire12976;
wire wire12978;
wire wire12979;
wire wire12981;
wire wire12984;
wire wire12985;
wire wire12986;
wire wire12988;
wire wire12989;
wire wire12991;
wire wire12992;
wire wire12995;
wire wire12996;
wire wire12998;
wire wire12999;
wire wire13001;
wire wire13003;
wire wire13005;
wire wire13006;
wire wire13008;
wire wire13013;
wire wire13015;
wire wire13016;
wire wire13017;
wire wire13020;
wire wire13022;
wire wire13025;
wire wire13026;
wire wire13027;
wire wire13028;
wire wire13029;
wire wire13034;
wire wire13035;
wire wire13036;
wire wire13039;
wire wire13042;
wire wire13044;
wire wire13046;
wire wire13048;
wire wire13049;
wire wire13050;
wire wire13053;
wire wire13054;
wire wire13055;
wire wire13056;
wire wire13057;
wire wire13059;
wire wire13060;
wire wire13062;
wire wire13063;
wire wire13065;
wire wire13066;
wire wire13067;
wire wire13069;
wire wire13070;
wire wire13073;
wire wire13074;
wire wire13077;
wire wire13078;
wire wire13080;
wire wire13084;
wire wire13085;
wire wire13087;
wire wire13088;
wire wire13090;
wire wire13091;
wire wire13093;
wire wire13095;
wire wire13096;
wire wire13100;
wire wire13101;
wire wire13104;
wire wire13105;
wire wire13106;
wire wire13107;
wire wire13108;
wire wire13111;
wire wire13113;
wire wire13114;
wire wire13117;
wire wire13118;
wire wire13119;
wire wire13120;
wire wire13123;
wire wire13124;
wire wire13126;
wire wire13127;
wire wire13128;
wire wire13132;
wire wire13133;
wire wire13136;
wire wire13140;
wire wire13141;
wire wire13144;
wire wire13146;
wire wire13147;
wire wire13149;
wire wire13151;
wire wire13153;
wire wire13154;
wire wire13156;
wire wire13162;
wire wire13163;
wire wire13166;
wire wire13170;
wire wire13171;
wire wire13172;
wire wire13173;
wire wire13174;
wire wire13176;
wire wire13177;
wire wire13178;
wire wire13181;
wire wire13182;
wire wire13183;
wire wire13185;
wire wire13187;
wire wire13188;
wire wire13193;
wire wire13194;
wire wire13198;
wire wire13199;
wire wire13202;
wire wire13203;
wire wire13208;
wire wire13209;
wire wire13211;
wire wire13213;
wire wire13215;
wire wire13216;
wire wire13217;
wire wire13218;
wire wire13222;
wire wire13223;
wire wire13224;
wire wire13225;
wire wire13228;
wire wire13229;
wire wire13231;
wire wire13233;
wire wire13234;
wire wire13236;
wire wire13237;
wire wire13239;
wire wire13240;
wire wire13244;
wire wire13246;
wire wire13248;
wire wire13249;
wire wire13250;
wire wire13251;
wire wire13254;
wire wire13256;
wire wire13259;
wire wire13260;
wire wire13261;
wire wire13263;
wire wire13264;
wire wire13265;
wire wire13266;
wire wire13268;
wire wire13269;
wire wire13270;
wire wire13272;
wire wire13274;
wire wire13275;
wire wire13277;
wire wire13278;
wire wire13283;
wire wire13284;
wire wire13285;
wire wire13287;
wire wire13288;
wire wire13291;
wire wire13292;
wire wire13293;
wire wire13294;
wire wire13296;
wire wire13297;
wire wire13298;
wire wire13301;
wire wire13303;
wire wire13304;
wire wire13305;
wire wire13306;
wire wire13308;
wire wire13310;
wire wire13311;
wire wire13313;
wire wire13314;
wire wire13317;
wire wire13318;
wire wire13320;
wire wire13322;
wire wire13323;
wire wire13325;
wire wire13327;
wire wire13329;
wire wire13333;
wire wire13334;
wire wire13337;
wire wire13338;
wire wire13341;
wire wire13342;
wire wire13346;
wire wire13347;
wire wire13350;
wire wire13351;
wire wire13352;
wire wire13354;
wire wire13355;
wire wire13359;
wire wire13360;
wire wire13361;
wire wire13364;
wire wire13365;
wire wire13368;
wire wire13370;
wire wire13372;
wire wire13374;
wire wire13378;
wire wire13380;
wire wire13381;
wire wire13384;
wire wire13385;
wire wire13390;
wire wire13391;
wire wire13392;
wire wire13393;
wire wire13394;
wire wire13397;
wire wire13398;
wire wire13399;
wire wire13400;
wire wire13401;
wire wire13404;
wire wire13405;
wire wire13406;
wire wire13408;
wire wire13409;
wire wire13410;
wire wire13411;
wire wire13413;
wire wire13414;
wire wire13415;
wire wire13417;
wire wire13419;
wire wire13421;
wire wire13422;
wire wire13424;
wire wire13425;
wire wire13428;
wire wire13429;
wire wire13430;
wire wire13431;
wire wire13432;
wire wire13436;
wire wire13437;
wire wire13438;
wire wire13439;
wire wire13441;
wire wire13443;
wire wire13445;
wire wire13446;
wire wire13448;
wire wire13450;
wire wire13452;
wire wire13454;
wire wire13455;
wire wire13457;
wire wire13458;
wire wire13459;
wire wire13461;
wire wire13462;
wire wire13463;
wire wire13465;
wire wire13467;
wire wire13468;
wire wire13470;
wire wire13471;
wire wire13473;
wire wire13474;
wire wire13475;
wire wire13478;
wire wire13479;
wire wire13481;
wire wire13482;
wire wire13487;
wire wire13488;
wire wire13493;
wire wire13494;
wire wire13495;
wire wire13496;
wire wire13497;
wire wire13501;
wire wire13502;
wire wire13503;
wire wire13504;
wire wire13505;
wire wire13506;
wire wire13508;
wire wire13509;
wire wire13510;
wire wire13512;
wire wire13513;
wire wire13515;
wire wire13516;
wire wire13519;
wire wire13520;
wire wire13521;
wire wire13522;
wire wire13523;
wire wire13524;
wire wire13525;
wire wire13526;
wire wire13528;
wire wire13529;
wire wire13531;
wire wire13532;
wire wire13534;
wire wire13535;
wire wire13538;
wire wire13539;
wire wire13541;
wire wire13542;
wire wire13543;
wire wire13544;
wire wire13546;
wire wire13547;
wire wire13550;
wire wire13552;
wire wire13553;
wire wire13554;
wire wire13557;
wire wire13559;
wire wire13560;
wire wire13561;
wire wire13562;
wire wire13566;
wire wire13567;
wire wire13569;
wire wire13572;
wire wire13573;
wire wire13576;
wire wire13577;
wire wire13580;
wire wire13585;
wire wire13586;
wire wire13591;
wire wire13592;
wire wire13598;
wire wire13599;
wire wire13601;
wire wire13606;
wire wire13607;
wire wire13611;
wire wire13612;
wire wire13616;
wire wire13617;
wire wire13622;
wire wire13623;
wire wire13629;
wire wire13630;
wire wire13635;
wire wire13636;
wire wire13638;
wire wire13643;
wire wire13644;
wire wire13648;
wire wire13650;
wire wire13651;
wire wire13656;
wire wire13657;
wire wire13660;
wire wire13662;
wire wire13663;
wire wire13665;
wire wire13666;
wire wire13670;
wire wire13672;
wire wire13673;
wire wire13674;
wire wire13679;
wire wire13681;
wire wire13683;
wire wire13684;
wire wire13689;
wire wire13690;
wire wire13694;
wire wire13696;
wire wire13697;
wire wire13698;
wire wire13703;
wire wire13704;
wire wire13709;
wire wire13710;
wire wire13713;
wire wire13714;
wire wire13717;
wire wire13719;
wire wire13720;
wire wire13725;
wire wire13726;
wire wire13728;
wire wire13729;
wire wire13735;
wire wire13736;
wire wire13741;
wire wire13742;
wire wire13746;
wire wire13747;
wire wire13752;
wire wire13753;
wire wire13755;
wire wire13756;
wire wire13759;
wire wire13760;
wire wire13765;
wire wire13767;
wire wire13768;
wire wire13772;
wire wire13773;
wire wire13776;
wire wire13777;
wire wire13779;
wire wire13780;
wire wire13782;
wire wire13788;
wire wire13789;
wire wire13790;
wire wire13791;
wire wire13792;
wire wire13796;
wire wire13797;
wire wire13798;
wire wire13800;
wire wire13801;
wire wire13803;
wire wire13804;
wire wire13807;
wire wire13808;
wire wire13810;
wire wire13812;
wire wire13813;
wire wire13815;
wire wire13816;
wire wire13818;
wire wire13820;
wire wire13823;
wire wire13824;
wire wire13825;
wire wire13827;
wire wire13833;
wire wire13834;
wire wire13836;
wire wire13837;
wire wire13840;
wire wire13841;
wire wire13843;
wire wire13844;
wire wire13850;
wire wire13854;
wire wire13855;
wire wire13856;
wire wire13857;
wire wire13860;
wire wire13865;
wire wire13866;
wire wire13867;
wire wire13869;
wire wire13870;
wire wire13872;
wire wire13873;
wire wire13874;
wire wire13877;
wire wire13878;
wire wire13880;
wire wire13881;
wire wire13883;
wire wire13884;
wire wire13885;
wire wire13887;
wire wire13888;
wire wire13891;
wire wire13892;
wire wire13893;
wire wire13895;
wire wire13896;
wire wire13897;
wire wire13900;
wire wire13902;
wire wire13903;
wire wire13904;
wire wire13905;
wire wire13906;
wire wire13910;
wire wire13911;
wire wire13913;
wire wire13914;
wire wire13915;
wire wire13918;
wire wire13919;
wire wire13920;
wire wire13923;
wire wire13924;
wire wire13929;
wire wire13931;
wire wire13932;
wire wire13934;
wire wire13935;
wire wire13938;
wire wire13940;
wire wire13942;
wire wire13943;
wire wire13944;
wire wire13947;
wire wire13948;
wire wire13951;
wire wire13952;
wire wire13954;
wire wire13955;
wire wire13957;
wire wire13960;
wire wire13961;
wire wire13962;
wire wire13963;
wire wire13964;
wire wire13966;
wire wire13967;
wire wire13968;
wire wire13969;
wire wire13970;
wire wire13971;
wire wire13972;
wire wire13975;
wire wire13976;
wire wire13977;
wire wire13978;
wire wire13979;
wire wire13981;
wire wire13982;
wire wire13983;
wire wire13985;
wire wire13989;
wire wire13990;
wire wire13991;
wire wire13992;
wire wire13995;
wire wire13996;
wire wire13997;
wire wire13999;
wire wire14000;
wire wire14001;
wire wire14003;
wire wire14006;
wire wire14007;
wire wire14009;
wire wire14010;
wire wire14011;
wire wire14012;
wire wire14015;
wire wire14016;
wire wire14018;
wire wire14020;
wire wire14021;
wire wire14023;
wire wire14024;
wire wire14025;
wire wire14027;
wire wire14028;
wire wire14029;
wire wire14031;
wire wire14033;
wire wire14034;
wire wire14036;
wire wire14037;
wire wire14040;
wire wire14041;
wire wire14042;
wire wire14043;
wire wire14045;
wire wire14046;
wire wire14047;
wire wire14049;
wire wire14050;
wire wire14055;
wire wire14056;
wire wire14057;
wire wire14058;
wire wire14061;
wire wire14062;
wire wire14065;
wire wire14066;
wire wire14068;
wire wire14071;
wire wire14072;
wire wire14077;
wire wire14078;
wire wire14079;
wire wire14080;
wire wire14082;
wire wire14087;
wire wire14088;
wire wire14091;
wire wire14092;
wire wire14094;
wire wire14097;
wire wire14099;
wire wire14101;
wire wire14103;
wire wire14105;
wire wire14106;
wire wire14107;
wire wire14111;
wire wire14112;
wire wire14115;
wire wire14116;
wire wire14120;
wire wire14121;
wire wire14126;
wire wire14127;
wire wire14128;
wire wire14131;
wire wire14133;
wire wire14134;
wire wire14138;
wire wire14139;
wire wire14141;
wire wire14142;
wire wire14143;
wire wire14144;
wire wire14147;
wire wire14148;
wire wire14149;
wire wire14150;
wire wire14153;
wire wire14154;
wire wire14155;
wire wire14157;
wire wire14158;
wire wire14159;
wire wire14160;
wire wire14161;
wire wire14163;
wire wire14164;
wire wire14168;
wire wire14169;
wire wire14171;
wire wire14173;
wire wire14174;
wire wire14177;
wire wire14178;
wire wire14179;
wire wire14183;
wire wire14186;
wire wire14191;
wire wire14192;
wire wire14195;
wire wire14198;
wire wire14199;
wire wire14200;
wire wire14202;
wire wire14203;
wire wire14205;
wire wire14208;
wire wire14209;
wire wire14211;
wire wire14213;
wire wire14214;
wire wire14216;
wire wire14218;
wire wire14219;
wire wire14222;
wire wire14226;
wire wire14227;
wire wire14232;
wire wire14233;
wire wire14238;
wire wire14239;
wire wire14240;
wire wire14241;
wire wire14245;
wire wire14246;
wire wire14252;
wire wire14253;
wire wire14254;
wire wire14256;
wire wire14260;
wire wire14261;
wire wire14267;
wire wire14268;
wire wire14272;
wire wire14273;
wire wire14275;
wire wire14277;
wire wire14278;
wire wire14280;
wire wire14281;
wire wire14283;
wire wire14284;
wire wire14285;
wire wire14290;
wire wire14291;
wire wire14293;
wire wire14295;
wire wire14296;
wire wire14301;
wire wire14302;
wire wire14307;
wire wire14308;
wire wire14310;
wire wire14311;
wire wire14316;
wire wire14317;
wire wire14320;
wire wire14322;
wire wire14323;
wire wire14329;
wire wire14330;
wire wire14332;
wire wire14334;
wire wire14337;
wire wire14338;
wire wire14340;
wire wire14341;
wire wire14343;
wire wire14344;
wire wire14346;
wire wire14347;
wire wire14349;
wire wire14350;
wire wire14351;
wire wire14355;
wire wire14356;
wire wire14357;
wire wire14361;
wire wire14362;
wire wire14363;
wire wire14365;
wire wire14367;
wire wire14369;
wire wire14371;
wire wire14373;
wire wire14375;
wire wire14376;
wire wire14377;
wire wire14378;
wire wire14380;
wire wire14381;
wire wire14384;
wire wire14385;
wire wire14387;
wire wire14388;
wire wire14393;
wire wire14396;
wire wire14397;
wire wire14398;
wire wire14401;
wire wire14403;
wire wire14404;
wire wire14405;
wire wire14408;
wire wire14409;
wire wire14410;
wire wire14413;
wire wire14414;
wire wire14415;
wire wire14416;
wire wire14419;
wire wire14420;
wire wire14422;
wire wire14423;
wire wire14426;
wire wire14428;
wire wire14429;
wire wire14430;
wire wire14432;
wire wire14434;
wire wire14436;
wire wire14438;
wire wire14439;
wire wire14440;
wire wire14441;
wire wire14442;
wire wire14443;
wire wire14444;
wire wire14445;
wire wire14446;
wire wire14448;
wire wire14452;
wire wire14453;
wire wire14454;
wire wire14455;
wire wire14458;
wire wire14460;
wire wire14461;
wire wire14464;
wire wire14466;
wire wire14467;
wire wire14468;
wire wire14470;
wire wire14471;
wire wire14473;
wire wire14476;
wire wire14479;
wire wire14480;
wire wire14484;
wire wire14485;
wire wire14486;
wire wire14489;
wire wire14490;
wire wire14492;
wire wire14493;
wire wire14495;
wire wire14496;
wire wire14498;
wire wire14499;
wire wire14500;
wire wire14503;
wire wire14505;
wire wire14507;
wire wire14508;
wire wire14510;
wire wire14511;
wire wire14513;
wire wire14514;
wire wire14517;
wire wire14518;
wire wire14519;
wire wire14520;
wire wire14521;
wire wire14522;
wire wire14523;
wire wire14524;
wire wire14526;
wire wire14528;
wire wire14530;
wire wire14533;
wire wire14534;
wire wire14536;
wire wire14537;
wire wire14540;
wire wire14542;
wire wire14544;
wire wire14545;
wire wire14549;
wire wire14550;
wire wire14551;
wire wire14552;
wire wire14554;
wire wire14555;
wire wire14557;
wire wire14558;
wire wire14560;
wire wire14561;
wire wire14563;
wire wire14564;
wire wire14566;
wire wire14567;
wire wire14570;
wire wire14572;
wire wire14573;
wire wire14577;
wire wire14578;
wire wire14579;
wire wire14580;
wire wire14582;
wire wire14583;
wire wire14587;
wire wire14588;
wire wire14589;
wire wire14591;
wire wire14592;
wire wire14594;
wire wire14595;
wire wire14598;
wire wire14599;
wire wire14601;
wire wire14603;
wire wire14605;
wire wire14606;
wire wire14609;
wire wire14610;
wire wire14613;
wire wire14614;
wire wire14615;
wire wire14618;
wire wire14619;
wire wire14621;
wire wire14622;
wire wire14623;
wire wire14624;
wire wire14625;
wire wire14629;
wire wire14631;
wire wire14635;
wire wire14637;
wire wire14638;
wire wire14641;
wire wire14644;
wire wire14645;
wire wire14646;
wire wire14648;
wire wire14649;
wire wire14652;
wire wire14654;
wire wire14655;
wire wire14656;
wire wire14658;
wire wire14659;
wire wire14661;
wire wire14662;
wire wire14664;
wire wire14665;
wire wire14667;
wire wire14669;
wire wire14671;
wire wire14672;
wire wire14673;
wire wire14674;
wire wire14675;
wire wire14678;
wire wire14680;
wire wire14681;
wire wire14683;
wire wire14684;
wire wire14689;
wire wire14690;
wire wire14691;
wire wire14692;
wire wire14694;
wire wire14695;
wire wire14697;
wire wire14701;
wire wire14702;
wire wire14706;
wire wire14708;
wire wire14709;
wire wire14714;
wire wire14715;
wire wire14717;
wire wire14718;
wire wire14719;
wire wire14723;
wire wire14724;
wire wire14725;
wire wire14726;
wire wire14729;
wire wire14730;
wire wire14733;
wire wire14735;
wire wire14738;
wire wire14739;
wire wire14740;
wire wire14742;
wire wire14743;
wire wire14745;
wire wire14747;
wire wire14748;
wire wire14750;
wire wire14751;
wire wire14752;
wire wire14754;
wire wire14756;
wire wire14759;
wire wire14760;
wire wire14761;
wire wire14762;
wire wire14764;
wire wire14766;
wire wire14768;
wire wire14770;
wire wire14772;
wire wire14774;
wire wire14775;
wire wire14777;
wire wire14778;
wire wire14779;
wire wire14782;
wire wire14784;
wire wire14785;
wire wire14790;
wire wire14791;
wire wire14795;
wire wire14796;
wire wire14797;
wire wire14801;
wire wire14802;
wire wire14803;
wire wire14807;
wire wire14808;
wire wire14810;
wire wire14814;
wire wire14816;
wire wire14817;
wire wire14819;
wire wire14820;
wire wire14825;
wire wire14826;
wire wire14829;
wire wire14830;
wire wire14831;
wire wire14833;
wire wire14834;
wire wire14836;
wire wire14838;
wire wire14839;
wire wire14843;
wire wire14845;
wire wire14846;
wire wire14848;
wire wire14854;
wire wire14855;
wire wire14859;
wire wire14861;
wire wire14862;
wire wire14867;
wire wire14868;
wire wire14870;
wire wire14873;
wire wire14875;
wire wire14876;
wire wire14881;
wire wire14882;
wire wire14886;
wire wire14887;
wire wire14890;
wire wire14892;
wire wire14894;
wire wire14896;
wire wire14898;
wire wire14899;
wire wire14903;
wire wire14904;
wire wire14905;
wire wire14909;
wire wire14910;
wire wire14911;
wire wire14912;
wire wire14914;
wire wire14915;
wire wire14917;
wire wire14918;
wire wire14920;
wire wire14922;
wire wire14923;
wire wire14924;
wire wire14927;
wire wire14931;
wire wire14933;
wire wire14935;
wire wire14937;
wire wire14938;
wire wire14939;
wire wire14940;
wire wire14942;
wire wire14943;
wire wire14944;
wire wire14946;
wire wire14948;
wire wire14949;
wire wire14954;
wire wire14955;
wire wire14956;
wire wire14957;
wire wire14958;
wire wire14960;
wire wire14961;
wire wire14962;
wire wire14964;
wire wire14965;
wire wire14967;
wire wire14969;
wire wire14970;
wire wire14971;
wire wire14974;
wire wire14975;
wire wire14978;
wire wire14979;
wire wire14980;
wire wire14982;
wire wire14983;
wire wire14985;
wire wire14986;
wire wire14987;
wire wire14988;
wire wire14990;
wire wire14991;
wire wire14992;
wire wire14993;
wire wire14995;
wire wire14996;
wire wire14999;
wire wire15000;
wire wire15001;
wire wire15002;
wire wire15005;
wire wire15006;
wire wire15007;
wire wire15008;
wire wire15010;
wire wire15011;
wire wire15012;
wire wire15016;
wire wire15019;
wire wire15020;
wire wire15021;
wire wire15024;
wire wire15025;
wire wire15028;
wire wire15029;
wire wire15032;
wire wire15033;
wire wire15035;
wire wire15037;
wire wire15038;
wire wire15040;
wire wire15042;
wire wire15043;
wire wire15044;
wire wire15045;
wire wire15046;
wire wire15048;
wire wire15049;
wire wire15052;
wire wire15053;
wire wire15055;
wire wire15057;
wire wire15058;
wire wire15059;
wire wire15061;
wire wire15062;
wire wire15063;
wire wire15065;
wire wire15066;
wire wire15069;
wire wire15071;
wire wire15073;
wire wire15075;
wire wire15077;
wire wire15079;
wire wire15080;
wire wire15082;
wire wire15083;
wire wire15084;
wire wire15085;
wire wire15089;
wire wire15090;
wire wire15091;
wire wire15094;
wire wire15095;
wire wire15097;
wire wire15099;
wire wire15101;
wire wire15103;
wire wire15108;
wire wire15109;
wire wire15111;
wire wire15112;
wire wire15113;
wire wire15115;
wire wire15117;
wire wire15120;
wire wire15121;
wire wire15122;
wire wire15123;
wire wire15125;
wire wire15126;
wire wire15127;
wire wire15130;
wire wire15131;
wire wire15132;
wire wire15133;
wire wire15135;
wire wire15136;
wire wire15137;
wire wire15140;
wire wire15141;
wire wire15142;
wire wire15143;
wire wire15144;
wire wire15145;
wire wire15149;
wire wire15150;
wire wire15151;
wire wire15153;
wire wire15154;
wire wire15155;
wire wire15159;
wire wire15160;
wire wire15162;
wire wire15163;
wire wire15165;
wire wire15166;
wire wire15169;
wire wire15174;
wire wire15175;
wire wire15178;
wire wire15179;
wire wire15180;
wire wire15182;
wire wire15184;
wire wire15185;
wire wire15186;
wire wire15188;
wire wire15189;
wire wire15192;
wire wire15194;
wire wire15195;
wire wire15198;
wire wire15200;
wire wire15203;
wire wire15204;
wire wire15206;
wire wire15207;
wire wire15208;
wire wire15211;
wire wire15212;
wire wire15216;
wire wire15217;
wire wire15218;
wire wire15219;
wire wire15221;
wire wire15222;
wire wire15223;
wire wire15224;
wire wire15226;
wire wire15227;
wire wire15230;
wire wire15231;
wire wire15234;
wire wire15235;
wire wire15239;
wire wire15241;
wire wire15243;
wire wire15245;
wire wire15246;
wire wire15247;
wire wire15249;
wire wire15252;
wire wire15254;
wire wire15255;
wire wire15257;
wire wire15258;
wire wire15261;
wire wire15263;
wire wire15264;
wire wire15266;
wire wire15269;
wire wire15270;
wire wire15273;
wire wire15274;
wire wire15275;
wire wire15278;
wire wire15279;
wire wire15280;
wire wire15283;
wire wire15284;
wire wire15285;
wire wire15287;
wire wire15288;
wire wire15289;
wire wire15290;
wire wire15291;
wire wire15292;
wire wire15294;
wire wire15296;
wire wire15297;
wire wire15299;
wire wire15300;
wire wire15304;
wire wire15307;
wire wire15308;
wire wire15310;
wire wire15312;
wire wire15315;
wire wire15316;
wire wire15321;
wire wire15322;
wire wire15326;
wire wire15328;
wire wire15329;
wire wire15333;
wire wire15334;
wire wire15340;
wire wire15341;
wire wire15342;
wire wire15348;
wire wire15349;
wire wire15354;
wire wire15355;
wire wire15360;
wire wire15361;
wire wire15367;
wire wire15368;
wire wire15374;
wire wire15375;
wire wire15376;
wire wire15382;
wire wire15383;
wire wire15385;
wire wire15389;
wire wire15390;
wire wire15396;
wire wire15397;
wire wire15398;
wire wire15400;
wire wire15405;
wire wire15406;
wire wire15412;
wire wire15413;
wire wire15416;
wire wire15418;
wire wire15421;
wire wire15423;
wire wire15426;
wire wire15428;
wire wire15431;
wire wire15432;
wire wire15434;
wire wire15435;
wire wire15437;
wire wire15438;
wire wire15440;
wire wire15444;
wire wire15445;
wire wire15448;
wire wire15451;
wire wire15452;
wire wire15456;
wire wire15459;
wire wire15460;
wire wire15463;
wire wire15467;
wire wire15468;
wire wire15469;
wire wire15471;
wire wire15472;
wire wire15474;
wire wire15475;
wire wire15478;
wire wire15479;
wire wire15481;
wire wire15482;
wire wire15483;
wire wire15485;
wire wire15488;
wire wire15489;
wire wire15490;
wire wire15493;
wire wire15494;
wire wire15495;
wire wire15498;
wire wire15499;
wire wire15501;
wire wire15502;
wire wire15504;
wire wire15506;
wire wire15507;
wire wire15509;
wire wire15511;
wire wire15512;
wire wire15517;
wire wire15518;
wire wire15521;
wire wire15525;
wire wire15526;
wire wire15527;
wire wire15529;
wire wire15532;
wire wire15533;
wire wire15534;
wire wire15536;
wire wire15537;
wire wire15538;
wire wire15539;
wire wire15542;
wire wire15543;
wire wire15544;
wire wire15545;
wire wire15546;
wire wire15549;
wire wire15551;
wire wire15554;
wire wire15555;
wire wire15557;
wire wire15559;
wire wire15560;
wire wire15562;
wire wire15564;
wire wire15565;
wire wire15569;
wire wire15570;
wire wire15573;
wire wire15574;
wire wire15575;
wire wire15576;
wire wire15578;
wire wire15579;
wire wire15582;
wire wire15583;
wire wire15586;
wire wire15587;
wire wire15589;
wire wire15590;
wire wire15591;
wire wire15593;
wire wire15594;
wire wire15595;
wire wire15596;
wire wire15597;
wire wire15598;
wire wire15601;
wire wire15602;
wire wire15605;
wire wire15606;
wire wire15609;
wire wire15610;
wire wire15612;
wire wire15614;
wire wire15616;
wire wire15617;
wire wire15620;
wire wire15621;
wire wire15623;
wire wire15624;
wire wire15626;
wire wire15627;
wire wire15628;
wire wire15629;
wire wire15633;
wire wire15634;
wire wire15639;
wire wire15640;
wire wire15642;
wire wire15647;
wire wire15648;
wire wire15649;
wire wire15651;
wire wire15653;
wire wire15654;
wire wire15658;
wire wire15659;
wire wire15660;
wire wire15663;
wire wire15665;
wire wire15666;
wire wire15667;
wire wire15671;
wire wire15672;
wire wire15674;
wire wire15675;
wire wire15677;
wire wire15678;
wire wire15680;
wire wire15681;
wire wire15683;
wire wire15684;
wire wire15685;
wire wire15686;
wire wire15688;
wire wire15689;
wire wire15693;
wire wire15695;
wire wire15696;
wire wire15697;
wire wire15698;
wire wire15700;
wire wire15701;
wire wire15702;
wire wire15704;
wire wire15705;
wire wire15707;
wire wire15709;
wire wire15710;
wire wire15712;
wire wire15714;
wire wire15715;
wire wire15718;
wire wire15719;
wire wire15721;
wire wire15723;
wire wire15724;
wire wire15725;
wire wire15726;
wire wire15728;
wire wire15729;
wire wire15733;
wire wire15734;
wire wire15738;
wire wire15739;
wire wire15741;
wire wire15742;
wire wire15743;
wire wire15746;
wire wire15747;
wire wire15748;
wire wire15750;
wire wire15754;
wire wire15756;
wire wire15757;
wire wire15758;
wire wire15760;
wire wire15761;
wire wire15763;
wire wire15764;
wire wire15766;
wire wire15767;
wire wire15769;
wire wire15770;
wire wire15773;
wire wire15774;
wire wire15775;
wire wire15776;
wire wire15778;
wire wire15781;
wire wire15782;
wire wire15784;
wire wire15786;
wire wire15790;
wire wire15791;
wire wire15792;
wire wire15794;
wire wire15795;
wire wire15798;
wire wire15799;
wire wire15800;
wire wire15802;
wire wire15804;
wire wire15805;
wire wire15807;
wire wire15808;
wire wire15811;
wire wire15813;
wire wire15816;
wire wire15817;
wire wire15819;
wire wire15822;
wire wire15823;
wire wire15829;
wire wire15830;
wire wire15834;
wire wire15836;
wire wire15837;
wire wire15838;
wire wire15841;
wire wire15842;
wire wire15843;
wire wire15844;
wire wire15845;
wire wire15848;
wire wire15851;
wire wire15852;
wire wire15858;
wire wire15859;
wire wire15864;
wire wire15865;
wire wire15870;
wire wire15871;
wire wire15873;
wire wire15875;
wire wire15876;
wire wire15879;
wire wire15880;
wire wire15885;
wire wire15886;
wire wire15887;
wire wire15892;
wire wire15894;
wire wire15895;
wire wire15897;
wire wire15898;
wire wire15899;
wire wire15901;
wire wire15902;
wire wire15903;
wire wire15908;
wire wire15909;
wire wire15914;
wire wire15915;
wire wire15920;
wire wire15922;
wire wire15924;
wire wire15927;
wire wire15930;
wire wire15931;
wire wire15937;
wire wire15938;
wire wire15941;
wire wire15943;
wire wire15945;
wire wire15947;
wire wire15950;
wire wire15951;
wire wire15952;
wire wire15954;
wire wire15955;
wire wire15957;
wire wire15961;
wire wire15962;
wire wire15964;
wire wire15967;
wire wire15968;
wire wire15970;
wire wire15972;
wire wire15973;
wire wire15975;
wire wire15977;
wire wire15978;
wire wire15980;
wire wire15982;
wire wire15983;
wire wire15985;
wire wire15987;
wire wire15989;
wire wire15991;
wire wire15993;
wire wire15995;
wire wire15996;
wire wire15999;
wire wire16001;
wire wire16002;
wire wire16003;
wire wire16004;
wire wire16007;
wire wire16008;
wire wire16009;
wire wire16011;
wire wire16012;
wire wire16014;
wire wire16015;
wire wire16016;
wire wire16018;
wire wire16019;
wire wire16020;
wire wire16022;
wire wire16023;
wire wire16025;
wire wire16028;
wire wire16030;
wire wire16031;
wire wire16032;
wire wire16034;
wire wire16035;
wire wire16038;
wire wire16040;
wire wire16041;
wire wire16045;
wire wire16046;
wire wire16048;
wire wire16052;
wire wire16053;
wire wire16056;
wire wire16057;
wire wire16059;
wire wire16060;
wire wire16064;
wire wire16065;
wire wire16069;
wire wire16070;
wire wire16072;
wire wire16075;
wire wire16077;
wire wire16078;
wire wire16081;
wire wire16082;
wire wire16083;
wire wire16086;
wire wire16087;
wire wire16088;
wire wire16089;
wire wire16091;
wire wire16093;
wire wire16094;
wire wire16095;
wire wire16098;
wire wire16099;
wire wire16102;
wire wire16103;
wire wire16105;
wire wire16109;
wire wire16110;
wire wire16112;
wire wire16114;
wire wire16119;
wire wire16120;
wire wire16121;
wire wire16124;
wire wire16125;
wire wire16127;
wire wire16128;
wire wire16130;
wire wire16131;
wire wire16132;
wire wire16134;
wire wire16135;
wire wire16138;
wire wire16139;
wire wire16140;
wire wire16141;
wire wire16144;
wire wire16145;
wire wire16146;
wire wire16148;
wire wire16149;
wire wire16152;
wire wire16153;
wire wire16155;
wire wire16157;
wire wire16158;
wire wire16159;
wire wire16164;
wire wire16165;
wire wire16166;
wire wire16168;
wire wire16170;
wire wire16171;
wire wire16173;
wire wire16174;
wire wire16175;
wire wire16176;
wire wire16179;
wire wire16180;
wire wire16182;
wire wire16184;
wire wire16185;
wire wire16186;
wire wire16188;
wire wire16189;
wire wire16192;
wire wire16193;
wire wire16194;
wire wire16195;
wire wire16198;
wire wire16201;
wire wire16203;
wire wire16204;
wire wire16206;
wire wire16207;
wire wire16211;
wire wire16212;
wire wire16213;
wire wire16214;
wire wire16215;
wire wire16217;
wire wire16220;
wire wire16222;
wire wire16224;
wire wire16228;
wire wire16229;
wire wire16232;
wire wire16233;
wire wire16236;
wire wire16238;
wire wire16240;
wire wire16241;
wire wire16245;
wire wire16246;
wire wire16248;
wire wire16249;
wire wire16251;
wire wire16253;
wire wire16254;
wire wire16256;
wire wire16257;
wire wire16258;
wire wire16259;
wire wire16262;
wire wire16263;
wire wire16266;
wire wire16267;
wire wire16270;
wire wire16272;
wire wire16273;
wire wire16278;
wire wire16279;
wire wire16280;
wire wire16282;
wire wire16286;
wire wire16288;
wire wire16289;
wire wire16291;
wire wire16293;
wire wire16294;
wire wire16296;
wire wire16297;
wire wire16299;
wire wire16300;
wire wire16305;
wire wire16306;
wire wire16308;
wire wire16309;
wire wire16310;
wire wire16312;
wire wire16313;
wire wire16316;
wire wire16318;
wire wire16320;
wire wire16323;
wire wire16324;
wire wire16327;
wire wire16331;
wire wire16334;
wire wire16335;
wire wire16339;
wire wire16340;
wire wire16342;
wire wire16345;
wire wire16346;
wire wire16347;
wire wire16349;
wire wire16350;
wire wire16351;
wire wire16352;
wire wire16355;
wire wire16356;
wire wire16360;
wire wire16362;
wire wire16363;
wire wire16366;
wire wire16367;
wire wire16368;
wire wire16373;
wire wire16374;
wire wire16375;
wire wire16378;
wire wire16379;
wire wire16382;
wire wire16383;
wire wire16385;
wire wire16386;
wire wire16388;
wire wire16389;
wire wire16394;
wire wire16395;
wire wire16396;
wire wire16399;
wire wire16404;
wire wire16405;
wire wire16408;
wire wire16409;
wire wire16410;
wire wire16411;
wire wire16412;
wire wire16415;
wire wire16420;
wire wire16421;
wire wire16423;
wire wire16424;
wire wire16427;
wire wire16430;
wire wire16431;
wire wire16435;
wire wire16436;
wire wire16438;
wire wire16440;
wire wire16442;
wire wire16443;
wire wire16445;
wire wire16447;
wire wire16448;
wire wire16449;
wire wire16450;
wire wire16453;
wire wire16454;
wire wire16456;
wire wire16460;
wire wire16461;
wire wire16462;
wire wire16463;
wire wire16465;
wire wire16466;
wire wire16468;
wire wire16470;
wire wire16475;
wire wire16476;
wire wire16479;
wire wire16480;
wire wire16482;
wire wire16483;
wire wire16487;
wire wire16488;
wire wire16490;
wire wire16492;
wire wire16493;
wire wire16494;
wire wire16497;
wire wire16498;
wire wire16500;
wire wire16503;
wire wire16504;
wire wire16506;
wire wire16508;
wire wire16509;
wire wire16514;
wire wire16516;
wire wire16518;
wire wire16520;
wire wire16521;
wire wire16526;
wire wire16527;
wire wire16530;
wire wire16531;
wire wire16533;
wire wire16537;
wire wire16538;
wire wire16539;
wire wire16544;
wire wire16545;
wire wire16546;
wire wire16548;
wire wire16549;
wire wire16551;
wire wire16552;
wire wire16556;
wire wire16557;
wire wire16560;
wire wire16562;
wire wire16563;
wire wire16566;
wire wire16567;
wire wire16568;
wire wire16570;
wire wire16571;
wire wire16572;
wire wire16573;
wire wire16574;
wire wire16576;
wire wire16578;
wire wire16580;
wire wire16581;
wire wire16585;
wire wire16586;
wire wire16587;
wire wire16590;
wire wire16591;
wire wire16593;
wire wire16594;
wire wire16596;
wire wire16598;
wire wire16599;
wire wire16601;
wire wire16602;
wire wire16603;
wire wire16605;
wire wire16606;
wire wire16609;
wire wire16611;
wire wire16612;
wire wire16617;
wire wire16618;
wire wire16621;
wire wire16622;
wire wire16623;
wire wire16627;
wire wire16628;
wire wire16629;
wire wire16631;
wire wire16632;
wire wire16633;
wire wire16635;
wire wire16636;
wire wire16637;
wire wire16638;
wire wire16641;
wire wire16642;
wire wire16644;
wire wire16645;
wire wire16646;
wire wire16650;
wire wire16651;
wire wire16656;
wire wire16657;
wire wire16658;
wire wire16661;
wire wire16662;
wire wire16663;
wire wire16665;
wire wire16666;
wire wire16669;
wire wire16670;
wire wire16673;
wire wire16674;
wire wire16676;
wire wire16677;
wire wire16678;
wire wire16679;
wire wire16682;
wire wire16683;
wire wire16685;
wire wire16686;
wire wire16690;
wire wire16691;
wire wire16692;
wire wire16693;
wire wire16696;
wire wire16698;
wire wire16699;
wire wire16702;
wire wire16704;
wire wire16705;
wire wire16709;
wire wire16710;
wire wire16711;
wire wire16715;
wire wire16716;
wire wire16717;
wire wire16718;
wire wire16719;
wire wire16721;
wire wire16723;
wire wire16724;
wire wire16728;
wire wire16730;
wire wire16731;
wire wire16733;
wire wire16734;
wire wire16739;
wire wire16740;
wire wire16742;
wire wire16744;
wire wire16745;
wire wire16748;
wire wire16749;
wire wire16753;
wire wire16754;
wire wire16755;
wire wire16758;
wire wire16760;
wire wire16761;
wire wire16763;
wire wire16769;
wire wire16770;
wire wire16773;
wire wire16774;
wire wire16775;
wire wire16776;
wire wire16777;
wire wire16784;
wire wire16785;
wire wire16788;
wire wire16790;
wire wire16791;
wire wire16795;
wire wire16796;
wire wire16798;
wire wire16799;
wire wire16804;
wire wire16805;
wire wire16811;
wire wire16812;
wire wire16818;
wire wire16819;
wire wire16820;
wire wire16823;
wire wire16825;
wire wire16827;
wire wire16829;
wire wire16830;
wire wire16831;
assign o_1_ = ( n_n1005 ) | ( n_n1004 ) | ( wire12040 ) | ( wire12041 ) ;
 assign o_2_ = ( wire12585 ) | ( wire12586 ) | ( wire12588 ) | ( wire12589 ) ;
 assign o_0_ = ( n_n621 ) | ( n_n620 ) | ( wire13136 ) | ( wire13147 ) ;
 assign o_9_ = ( n_n3986 ) | ( wire13572 ) | ( wire13573 ) | ( wire13684 ) ;
 assign o_7_ = ( n_n3251 ) | ( n_n3253 ) | ( wire14216 ) | ( wire14222 ) ;
 assign o_8_ = ( n_n3622 ) | ( wire14777 ) | ( wire14778 ) | ( wire14779 ) ;
 assign o_5_ = ( n_n2525 ) | ( n_n2523 ) | ( wire15299 ) | ( wire15300 ) ;
 assign o_6_ = ( n_n2898 ) | ( wire15816 ) | ( wire15817 ) ;
 assign o_3_ = ( n_n1784 ) | ( wire16323 ) | ( wire16324 ) ;
 assign o_4_ = ( n_n2155 ) | ( wire16830 ) | ( wire16831 ) ;
 assign n_n1014 = ( n_n1038 ) | ( wire11501 ) | ( wire11502 ) | ( wire11530 ) ;
 assign n_n4309 = ( n_n942 ) | ( n_n941 ) | ( n_n937 ) | ( wire11745 ) ;
 assign n_n1005 = ( n_n1012 ) | ( wire11832 ) | ( wire11833 ) | ( wire11894 ) ;
 assign n_n1004 = ( n_n1007 ) | ( n_n1009 ) | ( wire12036 ) | ( wire12037 ) ;
 assign n_n1396 = ( n_n1456 ) | ( n_n1455 ) | ( wire12197 ) | ( wire12200 ) ;
 assign n_n1397 = ( n_n1415 ) | ( wire12223 ) | ( wire12224 ) | ( wire12247 ) ;
 assign n_n1398 = ( n_n1418 ) | ( wire12431 ) | ( wire12432 ) | ( wire12440 ) ;
 assign n_n5305 = ( wire25  &  n_n473  &  n_n65 ) ;
 assign n_n5293 = ( wire15  &  n_n482  &  n_n65 ) ;
 assign n_n5296 = ( wire19  &  n_n526  &  n_n482 ) ;
 assign n_n5284 = ( wire19  &  n_n522  &  n_n491 ) ;
 assign n_n543 = ( n_n559 ) | ( wire12600 ) | ( wire12601 ) | ( wire12609 ) ;
 assign n_n562 = ( n_n4379 ) | ( n_n4399 ) | ( wire12699 ) | ( wire12700 ) ;
 assign n_n561 = ( n_n4458 ) | ( n_n4488 ) | ( wire12706 ) | ( wire12707 ) ;
 assign n_n563 = ( n_n4350 ) | ( n_n4331 ) | ( wire12713 ) | ( wire12714 ) ;
 assign n_n5297 = ( wire22  &  n_n482  &  n_n65 ) ;
 assign n_n3936 = ( n_n4378 ) | ( n_n4408 ) | ( wire13622 ) | ( wire13623 ) ;
 assign n_n3920 = ( n_n3931 ) | ( n_n3929 ) | ( wire13643 ) | ( wire13644 ) ;
 assign n_n3937 = ( n_n4362 ) | ( n_n4312 ) | ( wire13674 ) | ( wire13679 ) ;
 assign n_n3187 = ( n_n3194 ) | ( wire13714 ) | ( wire13728 ) | ( wire13729 ) ;
 assign n_n3192 = ( n_n3202 ) | ( n_n3204 ) | ( wire13759 ) | ( wire13760 ) ;
 assign n_n3191 = ( n_n3201 ) | ( wire13767 ) | ( wire13768 ) | ( wire13782 ) ;
 assign n_n3622 = ( n_n3629 ) | ( wire14513 ) | ( wire14514 ) | ( wire14540 ) ;
 assign n_n3624 = ( n_n3635 ) | ( wire14613 ) | ( wire14614 ) | ( wire14638 ) ;
 assign n_n3625 = ( n_n3639 ) | ( wire14654 ) | ( wire14655 ) | ( wire14684 ) ;
 assign n_n3626 = ( n_n3641 ) | ( wire14750 ) | ( wire14751 ) | ( wire14772 ) ;
 assign wire148 = ( i_9_  &  n_n524  &  n_n464  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n65 ) ;
 assign n_n2530 = ( n_n2548 ) | ( n_n2549 ) | ( wire14935 ) ;
 assign n_n2531 = ( n_n2551 ) | ( wire15005 ) | ( wire15006 ) | ( wire15025 ) ;
 assign n_n2525 = ( n_n2533 ) | ( wire15150 ) | ( wire15151 ) | ( wire15169 ) ;
 assign n_n2523 = ( n_n2528 ) | ( wire15206 ) | ( wire15207 ) | ( wire15297 ) ;
 assign n_n2845 = ( n_n4436 ) | ( n_n4417 ) | ( wire15307 ) | ( wire15308 ) ;
 assign n_n2846 = ( n_n4355 ) | ( n_n4335 ) | ( wire15321 ) | ( wire15322 ) ;
 assign n_n2827 = ( n_n2841 ) | ( wire15328 ) | ( wire15329 ) | ( wire15342 ) ;
 assign n_n2821 = ( n_n2837 ) | ( n_n2824 ) | ( n_n2835 ) | ( wire15400 ) ;
 assign n_n2826 = ( n_n2839 ) | ( wire15412 ) | ( wire15413 ) | ( wire15418 ) ;
 assign n_n2907 = ( n_n2929 ) | ( wire15437 ) | ( wire15438 ) | ( wire15463 ) ;
 assign n_n2906 = ( wire15501 ) | ( wire15502 ) | ( wire15504 ) ;
 assign n_n2908 = ( n_n2934 ) | ( wire15543 ) | ( wire15544 ) | ( wire15549 ) ;
 assign n_n2898 = ( n_n2905 ) | ( wire15742 ) | ( wire15743 ) | ( wire15808 ) ;
 assign n_n1793 = ( n_n1885 ) | ( n_n1886 ) | ( wire16025 ) | ( wire16028 ) ;
 assign n_n1792 = ( n_n1813 ) | ( n_n1812 ) | ( wire16072 ) ;
 assign n_n1794 = ( n_n1818 ) | ( wire16086 ) | ( wire16087 ) | ( wire16114 ) ;
 assign n_n1784 = ( n_n1789 ) | ( n_n1790 ) | ( wire16240 ) | ( wire16241 ) ;
 assign n_n1787 = ( n_n1797 ) | ( wire16262 ) | ( wire16263 ) | ( wire16289 ) ;
 assign n_n1786 = ( n_n1824 ) | ( n_n1826 ) | ( wire16316 ) | ( wire16318 ) ;
 assign n_n2104 = ( n_n4404 ) | ( n_n4413 ) | ( wire16475 ) | ( wire16476 ) ;
 assign n_n2087 = ( wire16492 ) | ( wire16493 ) | ( wire16494 ) | ( wire16497 ) ;
 assign n_n2086 = ( n_n2099 ) | ( wire16503 ) | ( wire16504 ) | ( wire16516 ) ;
 assign n_n2166 = ( n_n2190 ) | ( wire16545 ) | ( wire16546 ) | ( wire16557 ) ;
 assign n_n2105 = ( n_n4367 ) | ( n_n4374 ) | ( wire16650 ) | ( wire16651 ) ;
 assign n_n2155 = ( n_n2159 ) | ( wire16744 ) | ( wire16745 ) | ( wire16763 ) ;
 assign wire16 = ( i_9_  &  i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n4338 = ( wire16  &  n_n524  &  n_n518 ) ;
 assign wire21 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4339 = ( wire21  &  n_n536  &  n_n518 ) ;
 assign wire22 = ( (~ i_9_)  &  i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n4337 = ( wire22  &  n_n536  &  n_n518 ) ;
 assign n_n4401 = ( wire22  &  n_n536  &  n_n482 ) ;
 assign n_n4403 = ( wire21  &  n_n536  &  n_n482 ) ;
 assign n_n4400 = ( wire16  &  n_n526  &  n_n482 ) ;
 assign wire13 = ( i_9_  &  i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4464 = ( wire13  &  n_n526  &  n_n518 ) ;
 assign n_n4467 = ( wire21  &  n_n455  &  n_n518 ) ;
 assign wire11 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4463 = ( wire11  &  n_n455  &  n_n518 ) ;
 assign wire10 = ( i_9_  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n4666 = ( wire10  &  n_n473  &  n_n532 ) ;
 assign wire24 = ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4667 = ( wire24  &  n_n473  &  n_n390 ) ;
 assign n_n4664 = ( wire10  &  n_n473  &  n_n534 ) ;
 assign n_n4737 = ( wire22  &  n_n509  &  n_n325 ) ;
 assign wire14 = ( i_9_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4738 = ( wire14  &  n_n509  &  n_n524 ) ;
 assign n_n4735 = ( wire11  &  n_n509  &  n_n325 ) ;
 assign n_n4782 = ( wire14  &  n_n528  &  n_n482 ) ;
 assign n_n4784 = ( wire14  &  n_n526  &  n_n482 ) ;
 assign n_n4779 = ( wire24  &  n_n482  &  n_n325 ) ;
 assign wire17 = ( i_9_  &  i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n4830 = ( wire17  &  n_n535  &  n_n528 ) ;
 assign n_n4831 = ( wire11  &  n_n535  &  n_n260 ) ;
 assign n_n4900 = ( wire17  &  n_n522  &  n_n491 ) ;
 assign n_n4902 = ( wire17  &  n_n491  &  n_n520 ) ;
 assign n_n4898 = ( wire17  &  n_n524  &  n_n491 ) ;
 assign wire18 = ( i_9_  &  i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n4976 = ( wire18  &  n_n526  &  n_n518 ) ;
 assign n_n4977 = ( wire22  &  n_n518  &  n_n195 ) ;
 assign n_n4975 = ( wire11  &  n_n518  &  n_n195 ) ;
 assign n_n5038 = ( wire18  &  n_n528  &  n_n482 ) ;
 assign n_n5040 = ( wire18  &  n_n526  &  n_n482 ) ;
 assign n_n5034 = ( wire18  &  n_n482  &  n_n532 ) ;
 assign wire12 = ( i_9_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n5092 = ( wire12  &  n_n522  &  n_n535 ) ;
 assign wire20 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n5093 = ( wire20  &  n_n535  &  n_n130 ) ;
 assign n_n5091 = ( wire21  &  n_n535  &  n_n130 ) ;
 assign n_n4440 = ( wire13  &  n_n535  &  n_n534 ) ;
 assign n_n4434 = ( wire16  &  n_n524  &  n_n464 ) ;
 assign n_n4432 = ( wire16  &  n_n464  &  n_n526 ) ;
 assign wire98 = ( wire22  &  n_n536  &  n_n464 ) | ( wire11  &  n_n536  &  n_n464 ) ;
 assign wire233 = ( i_9_  &  n_n536  &  n_n464  &  n_n520 ) | ( (~ i_9_)  &  n_n536  &  n_n464  &  n_n520 ) ;
 assign wire236 = ( i_9_  &  n_n522  &  n_n536  &  n_n464 ) | ( (~ i_9_)  &  n_n522  &  n_n536  &  n_n464 ) ;
 assign n_n4720 = ( wire14  &  n_n526  &  n_n518 ) ;
 assign n_n4216 = ( n_n4720 ) | ( n_n4718 ) | ( n_n4717 ) ;
 assign n_n4857 = ( wire25  &  n_n509  &  n_n260 ) ;
 assign n_n4862 = ( wire17  &  n_n509  &  n_n528 ) ;
 assign n_n4856 = ( wire17  &  n_n509  &  n_n534 ) ;
 assign wire40 = ( wire22  &  n_n509  &  n_n260 ) | ( wire11  &  n_n509  &  n_n260 ) ;
 assign wire102 = ( i_9_  &  n_n520  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n520  &  n_n518  &  n_n260 ) ;
 assign wire245 = ( i_9_  &  n_n509  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n509  &  n_n532  &  n_n260 ) ;
 assign n_n4991 = ( wire11  &  n_n509  &  n_n195 ) ;
 assign n_n4996 = ( wire18  &  n_n509  &  n_n522 ) ;
 assign n_n4992 = ( wire18  &  n_n509  &  n_n526 ) ;
 assign n_n4995 = ( wire21  &  n_n509  &  n_n195 ) ;
 assign n_n4990 = ( wire18  &  n_n509  &  n_n528 ) ;
 assign n_n4998 = ( wire18  &  n_n509  &  n_n520 ) ;
 assign n_n4999 = ( wire23  &  n_n509  &  n_n195 ) ;
 assign wire103 = ( i_9_  &  n_n500  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n534  &  n_n195 ) ;
 assign wire25 = ( (~ i_9_)  &  i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n4617 = ( wire25  &  n_n500  &  n_n390 ) ;
 assign wire15 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n4637 = ( wire15  &  n_n491  &  n_n390 ) ;
 assign n_n4613 = ( wire20  &  n_n509  &  n_n390 ) ;
 assign n_n4927 = ( wire11  &  n_n473  &  n_n260 ) ;
 assign n_n4958 = ( wire18  &  n_n535  &  n_n528 ) ;
 assign n_n4920 = ( wire17  &  n_n473  &  n_n534 ) ;
 assign n_n4325 = ( wire20  &  n_n536  &  n_n535 ) ;
 assign wire23 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4327 = ( wire23  &  n_n536  &  n_n535 ) ;
 assign n_n4324 = ( wire16  &  n_n522  &  n_n535 ) ;
 assign n_n4382 = ( wire16  &  n_n528  &  n_n491 ) ;
 assign n_n4383 = ( wire11  &  n_n536  &  n_n491 ) ;
 assign n_n4380 = ( wire16  &  n_n491  &  n_n530 ) ;
 assign n_n4923 = ( wire24  &  n_n473  &  n_n260 ) ;
 assign n_n4924 = ( wire17  &  n_n473  &  n_n530 ) ;
 assign n_n4921 = ( wire25  &  n_n473  &  n_n260 ) ;
 assign n_n4982 = ( wire18  &  n_n520  &  n_n518 ) ;
 assign n_n4983 = ( wire23  &  n_n518  &  n_n195 ) ;
 assign n_n4981 = ( wire20  &  n_n518  &  n_n195 ) ;
 assign n_n5035 = ( wire24  &  n_n482  &  n_n195 ) ;
 assign n_n5032 = ( wire18  &  n_n482  &  n_n534 ) ;
 assign n_n5111 = ( wire23  &  n_n518  &  n_n130 ) ;
 assign n_n5112 = ( wire12  &  n_n509  &  n_n534 ) ;
 assign n_n5109 = ( wire20  &  n_n518  &  n_n130 ) ;
 assign n_n5171 = ( wire21  &  n_n482  &  n_n130 ) ;
 assign n_n5174 = ( wire12  &  n_n520  &  n_n482 ) ;
 assign n_n5167 = ( wire11  &  n_n482  &  n_n130 ) ;
 assign n_n4597 = ( wire20  &  n_n390  &  n_n518 ) ;
 assign n_n4598 = ( wire10  &  n_n520  &  n_n518 ) ;
 assign n_n4602 = ( wire10  &  n_n509  &  n_n532 ) ;
 assign n_n4593 = ( wire22  &  n_n390  &  n_n518 ) ;
 assign n_n4601 = ( wire25  &  n_n509  &  n_n390 ) ;
 assign wire108 = ( i_9_  &  n_n509  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n509  &  n_n390  &  n_n530 ) ;
 assign n_n4744 = ( wire14  &  n_n500  &  n_n534 ) ;
 assign n_n4754 = ( wire14  &  n_n524  &  n_n500 ) ;
 assign n_n4757 = ( wire20  &  n_n500  &  n_n325 ) ;
 assign n_n4749 = ( wire15  &  n_n500  &  n_n325 ) ;
 assign n_n4756 = ( wire14  &  n_n522  &  n_n500 ) ;
 assign wire109 = ( i_9_  &  n_n528  &  n_n500  &  n_n325 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n325 ) ;
 assign n_n4887 = ( wire23  &  n_n500  &  n_n260 ) ;
 assign n_n4888 = ( wire17  &  n_n491  &  n_n534 ) ;
 assign n_n4885 = ( wire20  &  n_n500  &  n_n260 ) ;
 assign n_n3450 = ( n_n4887 ) | ( n_n4888 ) | ( n_n4885 ) ;
 assign n_n4882 = ( wire17  &  n_n524  &  n_n500 ) ;
 assign n_n3451 = ( n_n4882 ) | ( n_n4884 ) | ( n_n4883 ) ;
 assign n_n5026 = ( wire18  &  n_n524  &  n_n491 ) ;
 assign n_n5027 = ( wire21  &  n_n491  &  n_n195 ) ;
 assign n_n5025 = ( wire22  &  n_n491  &  n_n195 ) ;
 assign wire114 = ( i_9_  &  n_n473  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n130 ) ;
 assign n_n5181 = ( wire15  &  n_n473  &  n_n130 ) ;
 assign n_n5184 = ( wire12  &  n_n473  &  n_n526 ) ;
 assign n_n5183 = ( wire11  &  n_n473  &  n_n130 ) ;
 assign wire112 = ( i_9_  &  n_n473  &  n_n524  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n130 ) ;
 assign n_n5310 = ( wire19  &  n_n473  &  n_n528 ) ;
 assign n_n5318 = ( wire19  &  n_n473  &  n_n520 ) ;
 assign n_n5314 = ( wire19  &  n_n473  &  n_n524 ) ;
 assign n_n5320 = ( wire19  &  n_n464  &  n_n534 ) ;
 assign wire459 = ( i_9_  &  n_n473  &  n_n526  &  n_n65 ) | ( (~ i_9_)  &  n_n473  &  n_n526  &  n_n65 ) ;
 assign n_n4615 = ( wire23  &  n_n509  &  n_n390 ) ;
 assign n_n4616 = ( wire10  &  n_n500  &  n_n534 ) ;
 assign n_n4607 = ( wire11  &  n_n509  &  n_n390 ) ;
 assign wire396 = ( wire10  &  n_n509  &  n_n526 ) | ( wire10  &  n_n509  &  n_n528 ) ;
 assign n_n3346 = ( n_n4615 ) | ( n_n4616 ) | ( wire14071 ) | ( wire14072 ) ;
 assign n_n4641 = ( wire22  &  n_n491  &  n_n390 ) ;
 assign n_n4634 = ( wire10  &  n_n491  &  n_n532 ) ;
 assign n_n4648 = ( wire10  &  n_n482  &  n_n534 ) ;
 assign n_n4618 = ( wire10  &  n_n500  &  n_n532 ) ;
 assign n_n4628 = ( wire10  &  n_n522  &  n_n500 ) ;
 assign wire26 = ( i_9_  &  n_n491  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n491  &  n_n390  &  n_n530 ) ;
 assign wire118 = ( wire24  &  n_n500  &  n_n390 ) | ( wire15  &  n_n500  &  n_n390 ) ;
 assign wire309 = ( wire21  &  n_n491  &  n_n390 ) | ( wire20  &  n_n491  &  n_n390 ) ;
 assign n_n3281 = ( n_n3346 ) | ( wire14077 ) | ( wire14078 ) | ( wire14082 ) ;
 assign n_n5050 = ( wire18  &  n_n473  &  n_n532 ) ;
 assign n_n5060 = ( wire18  &  n_n522  &  n_n473 ) ;
 assign n_n5055 = ( wire11  &  n_n473  &  n_n195 ) ;
 assign n_n5054 = ( wire18  &  n_n473  &  n_n528 ) ;
 assign n_n5059 = ( wire21  &  n_n473  &  n_n195 ) ;
 assign n_n5048 = ( wire18  &  n_n473  &  n_n534 ) ;
 assign n_n5028 = ( wire18  &  n_n522  &  n_n491 ) ;
 assign n_n5036 = ( wire18  &  n_n530  &  n_n482 ) ;
 assign wire50 = ( i_9_  &  n_n491  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n195 ) ;
 assign wire230 = ( n_n5039 ) | ( wire97 ) | ( wire13983 ) ;
 assign wire231 = ( i_9_  &  n_n482  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n195 ) ;
 assign wire356 = ( wire18  &  n_n522  &  n_n482 ) | ( wire18  &  n_n520  &  n_n482 ) ;
 assign n_n4571 = ( wire24  &  n_n535  &  n_n390 ) ;
 assign n_n4578 = ( wire10  &  n_n524  &  n_n535 ) ;
 assign n_n4570 = ( wire10  &  n_n535  &  n_n532 ) ;
 assign n_n4849 = ( wire22  &  n_n518  &  n_n260 ) ;
 assign n_n4853 = ( wire20  &  n_n518  &  n_n260 ) ;
 assign n_n4847 = ( wire11  &  n_n518  &  n_n260 ) ;
 assign n_n5096 = ( wire12  &  n_n534  &  n_n518 ) ;
 assign n_n5099 = ( wire24  &  n_n518  &  n_n130 ) ;
 assign n_n5085 = ( wire15  &  n_n535  &  n_n130 ) ;
 assign n_n4314 = ( wire16  &  n_n535  &  n_n532 ) ;
 assign n_n4389 = ( wire20  &  n_n536  &  n_n491 ) ;
 assign n_n4369 = ( wire22  &  n_n536  &  n_n500 ) ;
 assign n_n4381 = ( wire15  &  n_n536  &  n_n491 ) ;
 assign n_n4340 = ( wire16  &  n_n522  &  n_n518 ) ;
 assign wire280 = ( i_9_  &  n_n536  &  n_n491  &  n_n532 ) | ( (~ i_9_)  &  n_n536  &  n_n491  &  n_n532 ) ;
 assign n_n5101 = ( wire15  &  n_n518  &  n_n130 ) ;
 assign n_n5110 = ( wire12  &  n_n520  &  n_n518 ) ;
 assign n_n5142 = ( wire12  &  n_n500  &  n_n520 ) ;
 assign n_n5107 = ( wire21  &  n_n518  &  n_n130 ) ;
 assign n_n5130 = ( wire12  &  n_n500  &  n_n532 ) ;
 assign n_n5123 = ( wire21  &  n_n509  &  n_n130 ) ;
 assign n_n5129 = ( wire25  &  n_n500  &  n_n130 ) ;
 assign n_n5156 = ( wire12  &  n_n522  &  n_n491 ) ;
 assign n_n4317 = ( wire15  &  n_n536  &  n_n535 ) ;
 assign n_n4318 = ( wire16  &  n_n535  &  n_n528 ) ;
 assign n_n4388 = ( wire16  &  n_n522  &  n_n491 ) ;
 assign n_n4459 = ( wire24  &  n_n455  &  n_n518 ) ;
 assign n_n4461 = ( wire15  &  n_n455  &  n_n518 ) ;
 assign n_n4455 = ( wire23  &  n_n455  &  n_n535 ) ;
 assign n_n4513 = ( wire22  &  n_n455  &  n_n491 ) ;
 assign n_n4515 = ( wire21  &  n_n455  &  n_n491 ) ;
 assign n_n4512 = ( wire13  &  n_n526  &  n_n491 ) ;
 assign n_n4790 = ( wire14  &  n_n520  &  n_n482 ) ;
 assign n_n4791 = ( wire23  &  n_n482  &  n_n325 ) ;
 assign n_n4787 = ( wire21  &  n_n482  &  n_n325 ) ;
 assign n_n4859 = ( wire24  &  n_n509  &  n_n260 ) ;
 assign n_n4860 = ( wire17  &  n_n509  &  n_n530 ) ;
 assign n_n4858 = ( wire17  &  n_n509  &  n_n532 ) ;
 assign n_n4926 = ( wire17  &  n_n473  &  n_n528 ) ;
 assign n_n4928 = ( wire17  &  n_n473  &  n_n526 ) ;
 assign n_n4925 = ( wire15  &  n_n473  &  n_n260 ) ;
 assign n_n4988 = ( wire18  &  n_n509  &  n_n530 ) ;
 assign n_n4987 = ( wire24  &  n_n509  &  n_n195 ) ;
 assign n_n5041 = ( wire22  &  n_n482  &  n_n195 ) ;
 assign n_n5042 = ( wire18  &  n_n524  &  n_n482 ) ;
 assign n_n5100 = ( wire12  &  n_n530  &  n_n518 ) ;
 assign n_n4724 = ( wire14  &  n_n522  &  n_n518 ) ;
 assign n_n4727 = ( wire23  &  n_n325  &  n_n518 ) ;
 assign n_n4739 = ( wire21  &  n_n509  &  n_n325 ) ;
 assign wire95 = ( i_9_  &  n_n509  &  n_n528  &  n_n325 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n325 ) ;
 assign wire244 = ( wire14  &  n_n509  &  n_n532 ) | ( wire14  &  n_n509  &  n_n534 ) ;
 assign n_n4864 = ( wire17  &  n_n509  &  n_n526 ) ;
 assign n_n4868 = ( wire17  &  n_n509  &  n_n522 ) ;
 assign n_n5018 = ( wire18  &  n_n491  &  n_n532 ) ;
 assign n_n5022 = ( wire18  &  n_n528  &  n_n491 ) ;
 assign n_n5017 = ( wire25  &  n_n491  &  n_n195 ) ;
 assign wire135 = ( i_9_  &  n_n500  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n520  &  n_n195 ) ;
 assign wire296 = ( wire11  &  n_n491  &  n_n195 ) | ( wire15  &  n_n491  &  n_n195 ) ;
 assign n_n4993 = ( wire22  &  n_n509  &  n_n195 ) ;
 assign n_n1576 = ( n_n4996 ) | ( n_n4995 ) | ( n_n4994 ) ;
 assign wire134 = ( i_9_  &  n_n509  &  n_n530  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n530  &  n_n195 ) ;
 assign wire252 = ( wire18  &  n_n522  &  n_n518 ) | ( wire18  &  n_n520  &  n_n518 ) ;
 assign n_n5005 = ( wire15  &  n_n500  &  n_n195 ) ;
 assign n_n5004 = ( wire18  &  n_n500  &  n_n530 ) ;
 assign n_n5000 = ( wire18  &  n_n500  &  n_n534 ) ;
 assign wire136 = ( i_9_  &  n_n528  &  n_n500  &  n_n195 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n195 ) ;
 assign wire393 = ( i_9_  &  n_n500  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n532  &  n_n195 ) ;
 assign n_n4907 = ( wire24  &  n_n482  &  n_n260 ) ;
 assign n_n4913 = ( wire22  &  n_n482  &  n_n260 ) ;
 assign n_n4922 = ( wire17  &  n_n473  &  n_n532 ) ;
 assign n_n4934 = ( wire17  &  n_n473  &  n_n520 ) ;
 assign n_n2451 = ( wire14801 ) | ( wire14802 ) | ( wire14803 ) | ( wire14807 ) ;
 assign n_n2462 = ( n_n4951 ) | ( n_n5010 ) | ( wire14810 ) | ( wire14814 ) ;
 assign n_n2464 = ( n_n4886 ) | ( n_n4865 ) | ( wire14819 ) | ( wire14820 ) ;
 assign wire31 = ( i_9_  &  n_n473  &  n_n526  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n526  &  n_n260 ) ;
 assign n_n4453 = ( wire20  &  n_n455  &  n_n535 ) ;
 assign n_n4420 = ( wire16  &  n_n522  &  n_n473 ) ;
 assign n_n4407 = ( wire23  &  n_n536  &  n_n482 ) ;
 assign n_n2455 = ( n_n2470 ) | ( wire14833 ) | ( wire14834 ) | ( wire14848 ) ;
 assign n_n2454 = ( n_n2467 ) | ( wire14861 ) | ( wire14862 ) | ( wire14870 ) ;
 assign n_n2472 = ( n_n4391 ) | ( n_n4362 ) | ( wire14875 ) | ( wire14876 ) ;
 assign n_n2473 = ( n_n4316 ) | ( n_n4313 ) | ( wire14881 ) | ( wire14882 ) ;
 assign wire234 = ( wire13  &  n_n535  &  n_n530 ) | ( wire13  &  n_n535  &  n_n534 ) ;
 assign n_n4372 = ( wire16  &  n_n522  &  n_n500 ) ;
 assign n_n4373 = ( wire20  &  n_n536  &  n_n500 ) ;
 assign n_n4371 = ( wire21  &  n_n536  &  n_n500 ) ;
 assign n_n4431 = ( wire11  &  n_n536  &  n_n464 ) ;
 assign n_n4433 = ( wire22  &  n_n536  &  n_n464 ) ;
 assign n_n4430 = ( wire16  &  n_n464  &  n_n528 ) ;
 assign n_n4494 = ( wire13  &  n_n528  &  n_n500 ) ;
 assign n_n4491 = ( wire24  &  n_n455  &  n_n500 ) ;
 assign n_n4834 = ( wire17  &  n_n524  &  n_n535 ) ;
 assign n_n4835 = ( wire21  &  n_n535  &  n_n260 ) ;
 assign n_n4832 = ( wire17  &  n_n526  &  n_n535 ) ;
 assign n_n4909 = ( wire15  &  n_n482  &  n_n260 ) ;
 assign n_n4911 = ( wire11  &  n_n482  &  n_n260 ) ;
 assign n_n4903 = ( wire23  &  n_n491  &  n_n260 ) ;
 assign n_n4979 = ( wire21  &  n_n518  &  n_n195 ) ;
 assign n_n5049 = ( wire25  &  n_n473  &  n_n195 ) ;
 assign n_n5179 = ( wire24  &  n_n473  &  n_n130 ) ;
 assign n_n5239 = ( wire23  &  n_n518  &  n_n65 ) ;
 assign wire19 = ( i_9_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n5240 = ( wire19  &  n_n509  &  n_n534 ) ;
 assign n_n5238 = ( wire19  &  n_n520  &  n_n518 ) ;
 assign n_n4514 = ( wire13  &  n_n524  &  n_n491 ) ;
 assign n_n4247 = ( n_n4515 ) | ( n_n4514 ) | ( wire791 ) ;
 assign n_n4646 = ( wire10  &  n_n491  &  n_n520 ) ;
 assign n_n4644 = ( wire10  &  n_n522  &  n_n491 ) ;
 assign n_n4651 = ( wire24  &  n_n390  &  n_n482 ) ;
 assign n_n4649 = ( wire25  &  n_n390  &  n_n482 ) ;
 assign wire311 = ( i_9_  &  n_n390  &  n_n530  &  n_n482 ) | ( (~ i_9_)  &  n_n390  &  n_n530  &  n_n482 ) ;
 assign n_n4951 = ( wire23  &  n_n464  &  n_n260 ) ;
 assign n_n4952 = ( wire18  &  n_n535  &  n_n534 ) ;
 assign n_n4950 = ( wire17  &  n_n464  &  n_n520 ) ;
 assign n_n3803 = ( n_n4951 ) | ( n_n4952 ) | ( n_n4950 ) ;
 assign n_n4942 = ( wire17  &  n_n464  &  n_n528 ) ;
 assign n_n4943 = ( wire11  &  n_n464  &  n_n260 ) ;
 assign wire59 = ( wire15  &  n_n464  &  n_n260 ) ;
 assign n_n4945 = ( wire22  &  n_n464  &  n_n260 ) ;
 assign n_n4946 = ( wire17  &  n_n524  &  n_n464 ) ;
 assign n_n4949 = ( wire20  &  n_n464  &  n_n260 ) ;
 assign n_n2222 = ( n_n3803 ) | ( wire59 ) | ( wire12166 ) | ( wire16327 ) ;
 assign n_n5244 = ( wire19  &  n_n509  &  n_n530 ) ;
 assign n_n5245 = ( wire15  &  n_n509  &  n_n65 ) ;
 assign wire318 = ( i_9_  &  n_n509  &  n_n528  &  n_n65 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n65 ) ;
 assign n_n2200 = ( n_n5238 ) | ( n_n5244 ) | ( wire16685 ) | ( wire16686 ) ;
 assign n_n4450 = ( wire13  &  n_n524  &  n_n535 ) ;
 assign n_n4445 = ( wire15  &  n_n455  &  n_n535 ) ;
 assign n_n4444 = ( wire13  &  n_n535  &  n_n530 ) ;
 assign n_n4442 = ( wire13  &  n_n535  &  n_n532 ) ;
 assign n_n4441 = ( wire25  &  n_n455  &  n_n535 ) ;
 assign wire368 = ( wire21  &  n_n455  &  n_n535 ) | ( wire22  &  n_n455  &  n_n535 ) ;
 assign n_n4470 = ( wire13  &  n_n520  &  n_n518 ) ;
 assign n_n4460 = ( wire13  &  n_n530  &  n_n518 ) ;
 assign n_n4473 = ( wire25  &  n_n509  &  n_n455 ) ;
 assign n_n4466 = ( wire13  &  n_n524  &  n_n518 ) ;
 assign n_n4895 = ( wire11  &  n_n491  &  n_n260 ) ;
 assign n_n4890 = ( wire17  &  n_n491  &  n_n532 ) ;
 assign wire260 = ( i_9_  &  n_n500  &  n_n520  &  n_n260 ) | ( (~ i_9_)  &  n_n500  &  n_n520  &  n_n260 ) ;
 assign n_n2226 = ( n_n3451 ) | ( n_n4895 ) | ( n_n4890 ) | ( wire16331 ) ;
 assign n_n4850 = ( wire17  &  n_n524  &  n_n518 ) ;
 assign wire277 = ( i_9_  &  n_n522  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n260 ) ;
 assign wire295 = ( wire17  &  n_n509  &  n_n522 ) | ( wire17  &  n_n509  &  n_n524 ) ;
 assign n_n2228 = ( n_n4859 ) | ( n_n4864 ) | ( wire16334 ) | ( wire16335 ) ;
 assign n_n4881 = ( wire22  &  n_n500  &  n_n260 ) ;
 assign n_n4878 = ( wire17  &  n_n528  &  n_n500 ) ;
 assign n_n4880 = ( wire17  &  n_n526  &  n_n500 ) ;
 assign n_n4869 = ( wire20  &  n_n509  &  n_n260 ) ;
 assign n_n4877 = ( wire15  &  n_n500  &  n_n260 ) ;
 assign wire174 = ( wire24  &  n_n500  &  n_n260 ) | ( wire25  &  n_n500  &  n_n260 ) ;
 assign n_n2178 = ( n_n2226 ) | ( n_n2228 ) | ( wire16342 ) ;
 assign n_n5321 = ( wire25  &  n_n464  &  n_n65 ) ;
 assign n_n2274 = ( n_n5323 ) | ( n_n5324 ) | ( n_n5322 ) ;
 assign n_n5307 = ( wire24  &  n_n473  &  n_n65 ) ;
 assign n_n5326 = ( wire19  &  n_n464  &  n_n528 ) ;
 assign n_n5325 = ( wire15  &  n_n464  &  n_n65 ) ;
 assign n_n5332 = ( wire19  &  n_n522  &  n_n464 ) ;
 assign n_n5329 = ( wire22  &  n_n464  &  n_n65 ) ;
 assign wire117 = ( wire459 ) | ( wire115 ) | ( wire16291 ) ;
 assign wire269 = ( i_9_  &  n_n473  &  n_n528  &  n_n65 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n65 ) ;
 assign n_n2179 = ( n_n2230 ) | ( n_n2229 ) | ( wire16362 ) | ( wire16363 ) ;
 assign n_n4776 = ( wire14  &  n_n482  &  n_n534 ) ;
 assign n_n4774 = ( wire14  &  n_n491  &  n_n520 ) ;
 assign n_n4786 = ( wire14  &  n_n524  &  n_n482 ) ;
 assign wire131 = ( wire21  &  n_n482  &  n_n325 ) | ( wire22  &  n_n482  &  n_n325 ) ;
 assign wire313 = ( i_9_  &  n_n522  &  n_n482  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n482  &  n_n325 ) ;
 assign n_n2162 = ( n_n2178 ) | ( n_n2179 ) | ( wire16374 ) | ( wire16375 ) ;
 assign n_n4755 = ( wire21  &  n_n500  &  n_n325 ) ;
 assign n_n4759 = ( wire23  &  n_n500  &  n_n325 ) ;
 assign n_n4760 = ( wire14  &  n_n491  &  n_n534 ) ;
 assign n_n4758 = ( wire14  &  n_n500  &  n_n520 ) ;
 assign n_n2182 = ( n_n2238 ) | ( wire16394 ) | ( wire16395 ) | ( wire16399 ) ;
 assign n_n2183 = ( n_n2242 ) | ( wire16410 ) | ( wire16411 ) | ( wire16415 ) ;
 assign n_n2163 = ( n_n2182 ) | ( n_n2183 ) | ( wire16423 ) | ( wire16424 ) ;
 assign n_n4963 = ( wire21  &  n_n535  &  n_n195 ) ;
 assign n_n4959 = ( wire11  &  n_n535  &  n_n195 ) ;
 assign n_n4960 = ( wire18  &  n_n526  &  n_n535 ) ;
 assign n_n4964 = ( wire18  &  n_n522  &  n_n535 ) ;
 assign n_n2177 = ( n_n2223 ) | ( wire16449 ) | ( wire16450 ) | ( wire16456 ) ;
 assign wire250 = ( wire18  &  n_n535  &  n_n528 ) | ( wire18  &  n_n535  &  n_n530 ) ;
 assign n_n4817 = ( wire22  &  n_n464  &  n_n325 ) ;
 assign n_n4827 = ( wire24  &  n_n535  &  n_n260 ) ;
 assign n_n4816 = ( wire14  &  n_n464  &  n_n526 ) ;
 assign n_n5097 = ( wire25  &  n_n518  &  n_n130 ) ;
 assign n_n5019 = ( wire24  &  n_n491  &  n_n195 ) ;
 assign n_n4404 = ( wire16  &  n_n522  &  n_n482 ) ;
 assign n_n4413 = ( wire15  &  n_n536  &  n_n473 ) ;
 assign n_n4416 = ( wire16  &  n_n473  &  n_n526 ) ;
 assign n_n4523 = ( wire24  &  n_n455  &  n_n482 ) ;
 assign n_n4547 = ( wire21  &  n_n473  &  n_n455 ) ;
 assign n_n4539 = ( wire24  &  n_n473  &  n_n455 ) ;
 assign n_n4521 = ( wire25  &  n_n455  &  n_n482 ) ;
 assign n_n4544 = ( wire13  &  n_n473  &  n_n526 ) ;
 assign n_n4557 = ( wire15  &  n_n464  &  n_n455 ) ;
 assign n_n4560 = ( wire13  &  n_n464  &  n_n526 ) ;
 assign n_n4553 = ( wire25  &  n_n464  &  n_n455 ) ;
 assign n_n4800 = ( wire14  &  n_n473  &  n_n526 ) ;
 assign n_n2130 = ( n_n4777 ) | ( n_n4778 ) | ( n_n4780 ) ;
 assign n_n4803 = ( wire21  &  n_n473  &  n_n325 ) ;
 assign n_n4783 = ( wire11  &  n_n482  &  n_n325 ) ;
 assign n_n4812 = ( wire14  &  n_n464  &  n_n530 ) ;
 assign n_n4811 = ( wire24  &  n_n464  &  n_n325 ) ;
 assign n_n4781 = ( wire15  &  n_n482  &  n_n325 ) ;
 assign n_n2099 = ( n_n4674 ) | ( n_n4661 ) | ( wire16508 ) | ( wire16509 ) ;
 assign n_n4361 = ( wire25  &  n_n536  &  n_n500 ) ;
 assign n_n4363 = ( wire24  &  n_n536  &  n_n500 ) ;
 assign n_n4359 = ( wire23  &  n_n509  &  n_n536 ) ;
 assign n_n4438 = ( wire16  &  n_n464  &  n_n520 ) ;
 assign n_n4439 = ( wire23  &  n_n536  &  n_n464 ) ;
 assign n_n4437 = ( wire20  &  n_n536  &  n_n464 ) ;
 assign n_n4825 = ( wire25  &  n_n535  &  n_n260 ) ;
 assign n_n4828 = ( wire17  &  n_n535  &  n_n530 ) ;
 assign n_n4824 = ( wire17  &  n_n535  &  n_n534 ) ;
 assign n_n4879 = ( wire11  &  n_n500  &  n_n260 ) ;
 assign n_n4937 = ( wire25  &  n_n464  &  n_n260 ) ;
 assign n_n4938 = ( wire17  &  n_n464  &  n_n532 ) ;
 assign n_n4936 = ( wire17  &  n_n464  &  n_n534 ) ;
 assign n_n5010 = ( wire18  &  n_n524  &  n_n500 ) ;
 assign n_n5037 = ( wire15  &  n_n482  &  n_n195 ) ;
 assign n_n1570 = ( n_n5038 ) | ( n_n5035 ) | ( n_n5037 ) ;
 assign n_n5043 = ( wire21  &  n_n482  &  n_n195 ) ;
 assign n_n5045 = ( wire20  &  n_n482  &  n_n195 ) ;
 assign n_n5302 = ( wire19  &  n_n520  &  n_n482 ) ;
 assign n_n5294 = ( wire19  &  n_n528  &  n_n482 ) ;
 assign n_n4894 = ( wire17  &  n_n528  &  n_n491 ) ;
 assign n_n4916 = ( wire17  &  n_n522  &  n_n482 ) ;
 assign n_n4930 = ( wire17  &  n_n473  &  n_n524 ) ;
 assign n_n4947 = ( wire21  &  n_n464  &  n_n260 ) ;
 assign wire96 = ( wire17  &  n_n522  &  n_n491 ) | ( wire17  &  n_n491  &  n_n520 ) ;
 assign n_n5131 = ( wire24  &  n_n500  &  n_n130 ) ;
 assign n_n5137 = ( wire22  &  n_n500  &  n_n130 ) ;
 assign n_n5136 = ( wire12  &  n_n526  &  n_n500 ) ;
 assign n_n5200 = ( wire12  &  n_n464  &  n_n526 ) ;
 assign n_n5206 = ( wire12  &  n_n464  &  n_n520 ) ;
 assign n_n5146 = ( wire12  &  n_n491  &  n_n532 ) ;
 assign n_n5204 = ( wire12  &  n_n522  &  n_n464 ) ;
 assign n_n5191 = ( wire23  &  n_n473  &  n_n130 ) ;
 assign n_n5113 = ( wire25  &  n_n509  &  n_n130 ) ;
 assign n_n5081 = ( wire25  &  n_n535  &  n_n130 ) ;
 assign n_n5089 = ( wire22  &  n_n535  &  n_n130 ) ;
 assign n_n5124 = ( wire12  &  n_n509  &  n_n522 ) ;
 assign wire335 = ( wire12  &  n_n509  &  n_n530 ) | ( wire12  &  n_n509  &  n_n532 ) ;
 assign n_n5258 = ( wire19  &  n_n500  &  n_n532 ) ;
 assign n_n5274 = ( wire19  &  n_n491  &  n_n532 ) ;
 assign n_n5232 = ( wire19  &  n_n526  &  n_n518 ) ;
 assign n_n5255 = ( wire23  &  n_n509  &  n_n65 ) ;
 assign n_n5267 = ( wire21  &  n_n500  &  n_n65 ) ;
 assign n_n5222 = ( wire19  &  n_n535  &  n_n520 ) ;
 assign n_n5212 = ( wire19  &  n_n535  &  n_n530 ) ;
 assign n_n4344 = ( wire16  &  n_n509  &  n_n534 ) ;
 assign n_n4345 = ( wire25  &  n_n509  &  n_n536 ) ;
 assign n_n4343 = ( wire23  &  n_n536  &  n_n518 ) ;
 assign n_n4392 = ( wire16  &  n_n482  &  n_n534 ) ;
 assign n_n4393 = ( wire25  &  n_n536  &  n_n482 ) ;
 assign n_n4391 = ( wire23  &  n_n536  &  n_n491 ) ;
 assign n_n4612 = ( wire10  &  n_n509  &  n_n522 ) ;
 assign n_n4611 = ( wire21  &  n_n509  &  n_n390 ) ;
 assign n_n4669 = ( wire15  &  n_n473  &  n_n390 ) ;
 assign n_n4673 = ( wire22  &  n_n473  &  n_n390 ) ;
 assign n_n4668 = ( wire10  &  n_n473  &  n_n530 ) ;
 assign n_n4734 = ( wire14  &  n_n509  &  n_n528 ) ;
 assign n_n4733 = ( wire15  &  n_n509  &  n_n325 ) ;
 assign n_n4792 = ( wire14  &  n_n473  &  n_n534 ) ;
 assign n_n4854 = ( wire17  &  n_n520  &  n_n518 ) ;
 assign n_n4855 = ( wire23  &  n_n518  &  n_n260 ) ;
 assign n_n4912 = ( wire17  &  n_n526  &  n_n482 ) ;
 assign n_n4908 = ( wire17  &  n_n530  &  n_n482 ) ;
 assign n_n4966 = ( wire18  &  n_n535  &  n_n520 ) ;
 assign n_n4968 = ( wire18  &  n_n534  &  n_n518 ) ;
 assign n_n5014 = ( wire18  &  n_n500  &  n_n520 ) ;
 assign n_n5015 = ( wire23  &  n_n500  &  n_n195 ) ;
 assign n_n5012 = ( wire18  &  n_n522  &  n_n500 ) ;
 assign n_n5067 = ( wire24  &  n_n464  &  n_n195 ) ;
 assign n_n5069 = ( wire15  &  n_n464  &  n_n195 ) ;
 assign n_n5066 = ( wire18  &  n_n464  &  n_n532 ) ;
 assign n_n5241 = ( wire25  &  n_n509  &  n_n65 ) ;
 assign n_n5243 = ( wire24  &  n_n509  &  n_n65 ) ;
 assign n_n5300 = ( wire19  &  n_n522  &  n_n482 ) ;
 assign n_n5299 = ( wire21  &  n_n482  &  n_n65 ) ;
 assign n_n4364 = ( wire16  &  n_n500  &  n_n530 ) ;
 assign n_n4362 = ( wire16  &  n_n500  &  n_n532 ) ;
 assign n_n3533 = ( n_n4363 ) | ( n_n4364 ) | ( n_n4362 ) ;
 assign n_n4366 = ( wire16  &  n_n528  &  n_n500 ) ;
 assign n_n4367 = ( wire11  &  n_n536  &  n_n500 ) ;
 assign n_n4365 = ( wire15  &  n_n536  &  n_n500 ) ;
 assign n_n1308 = ( wire11607 ) | ( wire15  &  n_n536  &  n_n500 ) ;
 assign n_n4770 = ( wire14  &  n_n524  &  n_n491 ) ;
 assign n_n4769 = ( wire22  &  n_n491  &  n_n325 ) ;
 assign n_n4767 = ( wire11  &  n_n491  &  n_n325 ) ;
 assign n_n4764 = ( wire14  &  n_n491  &  n_n530 ) ;
 assign n_n4905 = ( wire25  &  n_n482  &  n_n260 ) ;
 assign wire352 = ( wire17  &  n_n482  &  n_n532 ) | ( wire17  &  n_n482  &  n_n534 ) ;
 assign n_n5046 = ( wire18  &  n_n520  &  n_n482 ) ;
 assign n_n5056 = ( wire18  &  n_n473  &  n_n526 ) ;
 assign n_n5057 = ( wire22  &  n_n473  &  n_n195 ) ;
 assign wire166 = ( i_9_  &  n_n473  &  n_n530  &  n_n195 ) | ( (~ i_9_)  &  n_n473  &  n_n530  &  n_n195 ) ;
 assign wire292 = ( i_9_  &  n_n520  &  n_n482  &  n_n325 ) | ( (~ i_9_)  &  n_n520  &  n_n482  &  n_n325 ) ;
 assign n_n4843 = ( wire24  &  n_n518  &  n_n260 ) ;
 assign n_n4845 = ( wire15  &  n_n518  &  n_n260 ) ;
 assign n_n4846 = ( wire17  &  n_n528  &  n_n518 ) ;
 assign n_n4848 = ( wire17  &  n_n526  &  n_n518 ) ;
 assign n_n3820 = ( n_n4839 ) | ( n_n4840 ) | ( n_n4838 ) ;
 assign n_n4384 = ( wire16  &  n_n526  &  n_n491 ) ;
 assign n_n4390 = ( wire16  &  n_n491  &  n_n520 ) ;
 assign n_n4374 = ( wire16  &  n_n500  &  n_n520 ) ;
 assign n_n4638 = ( wire10  &  n_n528  &  n_n491 ) ;
 assign n_n4633 = ( wire25  &  n_n491  &  n_n390 ) ;
 assign n_n5155 = ( wire21  &  n_n491  &  n_n130 ) ;
 assign n_n5161 = ( wire25  &  n_n482  &  n_n130 ) ;
 assign n_n509 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n522 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n536 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n473 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n524 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4425 = ( wire25  &  n_n536  &  n_n464 ) ;
 assign n_n464 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n526 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n455 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n535 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n528 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4482 = ( wire13  &  n_n509  &  n_n524 ) ;
 assign n_n4489 = ( wire25  &  n_n455  &  n_n500 ) ;
 assign n_n500 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign n_n4504 = ( wire13  &  n_n491  &  n_n534 ) ;
 assign n_n4511 = ( wire11  &  n_n455  &  n_n491 ) ;
 assign n_n491 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n520 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n4526 = ( wire13  &  n_n528  &  n_n482 ) ;
 assign n_n4533 = ( wire20  &  n_n455  &  n_n482 ) ;
 assign n_n4554 = ( wire13  &  n_n464  &  n_n532 ) ;
 assign n_n4561 = ( wire22  &  n_n464  &  n_n455 ) ;
 assign n_n4568 = ( wire10  &  n_n535  &  n_n534 ) ;
 assign n_n4575 = ( wire11  &  n_n535  &  n_n390 ) ;
 assign n_n390 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n4590 = ( wire10  &  n_n528  &  n_n518 ) ;
 assign n_n530 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n4640 = ( wire10  &  n_n526  &  n_n491 ) ;
 assign n_n4647 = ( wire23  &  n_n491  &  n_n390 ) ;
 assign n_n482 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n4662 = ( wire10  &  n_n520  &  n_n482 ) ;
 assign n_n532 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n4690 = ( wire10  &  n_n524  &  n_n464 ) ;
 assign n_n534 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign n_n325 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n4704 = ( wire14  &  n_n526  &  n_n535 ) ;
 assign n_n4711 = ( wire23  &  n_n535  &  n_n325 ) ;
 assign n_n518 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n4748 = ( wire14  &  n_n500  &  n_n530 ) ;
 assign n_n4777 = ( wire25  &  n_n482  &  n_n325 ) ;
 assign n_n4821 = ( wire20  &  n_n464  &  n_n325 ) ;
 assign n_n260 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n4901 = ( wire20  &  n_n491  &  n_n260 ) ;
 assign n_n195 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n4974 = ( wire18  &  n_n528  &  n_n518 ) ;
 assign n_n5003 = ( wire24  &  n_n500  &  n_n195 ) ;
 assign n_n5047 = ( wire23  &  n_n482  &  n_n195 ) ;
 assign n_n130 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n5098 = ( wire12  &  n_n532  &  n_n518 ) ;
 assign n_n5105 = ( wire22  &  n_n518  &  n_n130 ) ;
 assign n_n5120 = ( wire12  &  n_n509  &  n_n526 ) ;
 assign n_n5127 = ( wire23  &  n_n509  &  n_n130 ) ;
 assign n_n5186 = ( wire12  &  n_n473  &  n_n524 ) ;
 assign n_n5193 = ( wire25  &  n_n464  &  n_n130 ) ;
 assign n_n65 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n5251 = ( wire21  &  n_n509  &  n_n65 ) ;
 assign n_n5266 = ( wire19  &  n_n524  &  n_n500 ) ;
 assign n_n5273 = ( wire25  &  n_n491  &  n_n65 ) ;
 assign n_n4347 = ( wire24  &  n_n509  &  n_n536 ) ;
 assign n_n4397 = ( wire15  &  n_n536  &  n_n482 ) ;
 assign n_n4398 = ( wire16  &  n_n528  &  n_n482 ) ;
 assign n_n4396 = ( wire16  &  n_n530  &  n_n482 ) ;
 assign n_n4524 = ( wire13  &  n_n530  &  n_n482 ) ;
 assign n_n4522 = ( wire13  &  n_n482  &  n_n532 ) ;
 assign wire170 = ( i_9_  &  n_n455  &  n_n482  &  n_n532 ) | ( (~ i_9_)  &  n_n455  &  n_n482  &  n_n532 ) ;
 assign n_n4246 = ( wire170 ) | ( wire13  &  n_n530  &  n_n482 ) ;
 assign n_n4670 = ( wire10  &  n_n473  &  n_n528 ) ;
 assign n_n4732 = ( wire14  &  n_n509  &  n_n530 ) ;
 assign n_n4789 = ( wire20  &  n_n482  &  n_n325 ) ;
 assign n_n4906 = ( wire17  &  n_n482  &  n_n532 ) ;
 assign n_n4967 = ( wire23  &  n_n535  &  n_n195 ) ;
 assign n_n5086 = ( wire12  &  n_n535  &  n_n528 ) ;
 assign n_n5087 = ( wire11  &  n_n535  &  n_n130 ) ;
 assign n_n4589 = ( wire15  &  n_n390  &  n_n518 ) ;
 assign n_n4587 = ( wire24  &  n_n390  &  n_n518 ) ;
 assign n_n881 = ( n_n4590 ) | ( n_n4589 ) | ( n_n4587 ) ;
 assign n_n4594 = ( wire10  &  n_n524  &  n_n518 ) ;
 assign n_n4083 = ( n_n4593 ) | ( n_n881 ) | ( n_n4594 ) | ( wire13441 ) ;
 assign n_n4639 = ( wire11  &  n_n491  &  n_n390 ) ;
 assign n_n4904 = ( wire17  &  n_n482  &  n_n534 ) ;
 assign n_n4319 = ( wire11  &  n_n536  &  n_n535 ) ;
 assign n_n4320 = ( wire16  &  n_n526  &  n_n535 ) ;
 assign n_n4451 = ( wire21  &  n_n455  &  n_n535 ) ;
 assign n_n4918 = ( wire17  &  n_n520  &  n_n482 ) ;
 assign n_n4919 = ( wire23  &  n_n482  &  n_n260 ) ;
 assign n_n4917 = ( wire20  &  n_n482  &  n_n260 ) ;
 assign n_n4985 = ( wire25  &  n_n509  &  n_n195 ) ;
 assign n_n4984 = ( wire18  &  n_n509  &  n_n534 ) ;
 assign n_n5031 = ( wire23  &  n_n491  &  n_n195 ) ;
 assign n_n5114 = ( wire12  &  n_n509  &  n_n532 ) ;
 assign n_n5116 = ( wire12  &  n_n509  &  n_n530 ) ;
 assign n_n5162 = ( wire12  &  n_n482  &  n_n532 ) ;
 assign n_n4582 = ( wire10  &  n_n535  &  n_n520 ) ;
 assign n_n4584 = ( wire10  &  n_n534  &  n_n518 ) ;
 assign n_n4586 = ( wire10  &  n_n532  &  n_n518 ) ;
 assign wire365 = ( i_9_  &  n_n390  &  n_n530  &  n_n518 ) | ( (~ i_9_)  &  n_n390  &  n_n530  &  n_n518 ) ;
 assign n_n3348 = ( n_n4582 ) | ( n_n4584 ) | ( wire14091 ) | ( wire14092 ) ;
 assign n_n4876 = ( wire17  &  n_n500  &  n_n530 ) ;
 assign wire461 = ( n_n4870 ) | ( n_n4871 ) | ( n_n4872 ) ;
 assign n_n3326 = ( n_n4879 ) | ( n_n4876 ) | ( wire461 ) | ( wire13850 ) ;
 assign n_n5327 = ( wire11  &  n_n464  &  n_n65 ) ;
 assign n_n2643 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5327 ) ;
 assign n_n5323 = ( wire24  &  n_n464  &  n_n65 ) ;
 assign n_n5324 = ( wire19  &  n_n464  &  n_n530 ) ;
 assign n_n5322 = ( wire19  &  n_n464  &  n_n532 ) ;
 assign n_n4577 = ( wire22  &  n_n535  &  n_n390 ) ;
 assign n_n4576 = ( wire10  &  n_n526  &  n_n535 ) ;
 assign n_n4569 = ( wire25  &  n_n535  &  n_n390 ) ;
 assign n_n4574 = ( wire10  &  n_n535  &  n_n528 ) ;
 assign n_n4581 = ( wire20  &  n_n535  &  n_n390 ) ;
 assign n_n4572 = ( wire10  &  n_n535  &  n_n530 ) ;
 assign n_n4573 = ( wire15  &  n_n535  &  n_n390 ) ;
 assign n_n4579 = ( wire21  &  n_n535  &  n_n390 ) ;
 assign n_n3282 = ( n_n3348 ) | ( wire14087 ) | ( wire14088 ) | ( wire14101 ) ;
 assign n_n4538 = ( wire13  &  n_n473  &  n_n532 ) ;
 assign n_n4525 = ( wire15  &  n_n455  &  n_n482 ) ;
 assign n_n4531 = ( wire21  &  n_n455  &  n_n482 ) ;
 assign n_n3871 = ( n_n4553 ) | ( n_n4551 ) | ( n_n4552 ) ;
 assign wire202 = ( wire212 ) | ( n_n4550 ) | ( n_n4543 ) | ( wire14107 ) ;
 assign n_n3260 = ( n_n3281 ) | ( n_n3282 ) | ( wire14115 ) | ( wire14116 ) ;
 assign n_n4629 = ( wire20  &  n_n500  &  n_n390 ) ;
 assign n_n4583 = ( wire23  &  n_n535  &  n_n390 ) ;
 assign n_n4842 = ( wire17  &  n_n532  &  n_n518 ) ;
 assign n_n4844 = ( wire17  &  n_n530  &  n_n518 ) ;
 assign n_n4839 = ( wire23  &  n_n535  &  n_n260 ) ;
 assign n_n5303 = ( wire23  &  n_n482  &  n_n65 ) ;
 assign n_n5182 = ( wire12  &  n_n473  &  n_n528 ) ;
 assign n_n5173 = ( wire20  &  n_n482  &  n_n130 ) ;
 assign n_n5165 = ( wire15  &  n_n482  &  n_n130 ) ;
 assign n_n5230 = ( wire19  &  n_n528  &  n_n518 ) ;
 assign n_n5166 = ( wire12  &  n_n528  &  n_n482 ) ;
 assign n_n5163 = ( wire24  &  n_n482  &  n_n130 ) ;
 assign n_n5214 = ( wire19  &  n_n535  &  n_n528 ) ;
 assign n_n4994 = ( wire18  &  n_n509  &  n_n524 ) ;
 assign n_n5002 = ( wire18  &  n_n500  &  n_n532 ) ;
 assign n_n5053 = ( wire15  &  n_n473  &  n_n195 ) ;
 assign n_n5033 = ( wire25  &  n_n482  &  n_n195 ) ;
 assign n_n5051 = ( wire24  &  n_n473  &  n_n195 ) ;
 assign n_n5006 = ( wire18  &  n_n528  &  n_n500 ) ;
 assign n_n4454 = ( wire13  &  n_n535  &  n_n520 ) ;
 assign n_n4518 = ( wire13  &  n_n491  &  n_n520 ) ;
 assign n_n4517 = ( wire20  &  n_n455  &  n_n491 ) ;
 assign n_n3152 = ( n_n4518 ) | ( n_n4517 ) | ( wire664 ) ;
 assign n_n4725 = ( wire20  &  n_n325  &  n_n518 ) ;
 assign n_n4726 = ( wire14  &  n_n520  &  n_n518 ) ;
 assign n_n4861 = ( wire15  &  n_n509  &  n_n260 ) ;
 assign n_n5039 = ( wire11  &  n_n482  &  n_n195 ) ;
 assign n_n5103 = ( wire11  &  n_n518  &  n_n130 ) ;
 assign n_n5104 = ( wire12  &  n_n526  &  n_n518 ) ;
 assign n_n5102 = ( wire12  &  n_n528  &  n_n518 ) ;
 assign n_n4395 = ( wire24  &  n_n536  &  n_n482 ) ;
 assign n_n2638 = ( n_n4366 ) | ( n_n4357 ) | ( wire15032 ) | ( wire15033 ) ;
 assign wire425 = ( i_9_  &  n_n536  &  n_n524  &  n_n491 ) | ( (~ i_9_)  &  n_n536  &  n_n524  &  n_n491 ) ;
 assign n_n2560 = ( n_n2638 ) | ( wire15028 ) | ( wire15029 ) | ( wire15040 ) ;
 assign n_n4426 = ( wire16  &  n_n464  &  n_n532 ) ;
 assign n_n2635 = ( n_n4404 ) | ( n_n4409 ) | ( wire15048 ) | ( wire15049 ) ;
 assign wire37 = ( i_9_  &  n_n536  &  n_n464  &  n_n534 ) | ( (~ i_9_)  &  n_n536  &  n_n464  &  n_n534 ) ;
 assign n_n2559 = ( n_n2635 ) | ( wire15044 ) | ( wire15045 ) | ( wire15055 ) ;
 assign n_n4315 = ( wire24  &  n_n536  &  n_n535 ) ;
 assign n_n4312 = ( wire16  &  n_n535  &  n_n534 ) ;
 assign n_n4360 = ( wire16  &  n_n500  &  n_n534 ) ;
 assign n_n4487 = ( wire23  &  n_n509  &  n_n455 ) ;
 assign n_n4483 = ( wire21  &  n_n509  &  n_n455 ) ;
 assign n_n4840 = ( wire17  &  n_n534  &  n_n518 ) ;
 assign n_n4837 = ( wire20  &  n_n535  &  n_n260 ) ;
 assign n_n4899 = ( wire21  &  n_n491  &  n_n260 ) ;
 assign n_n4986 = ( wire18  &  n_n509  &  n_n532 ) ;
 assign n_n5044 = ( wire18  &  n_n522  &  n_n482 ) ;
 assign n_n5115 = ( wire24  &  n_n509  &  n_n130 ) ;
 assign n_n5175 = ( wire23  &  n_n482  &  n_n130 ) ;
 assign n_n5177 = ( wire25  &  n_n473  &  n_n130 ) ;
 assign n_n5311 = ( wire11  &  n_n473  &  n_n65 ) ;
 assign n_n4798 = ( wire14  &  n_n473  &  n_n528 ) ;
 assign n_n4804 = ( wire14  &  n_n522  &  n_n473 ) ;
 assign n_n4794 = ( wire14  &  n_n473  &  n_n532 ) ;
 assign n_n4795 = ( wire24  &  n_n473  &  n_n325 ) ;
 assign n_n4793 = ( wire25  &  n_n473  &  n_n325 ) ;
 assign n_n4796 = ( wire14  &  n_n473  &  n_n530 ) ;
 assign n_n4797 = ( wire15  &  n_n473  &  n_n325 ) ;
 assign n_n4801 = ( wire22  &  n_n473  &  n_n325 ) ;
 assign n_n4933 = ( wire20  &  n_n473  &  n_n260 ) ;
 assign n_n4935 = ( wire23  &  n_n473  &  n_n260 ) ;
 assign wire249 = ( n_n4927 ) | ( n_n4924 ) | ( n_n4926 ) | ( n_n4925 ) ;
 assign n_n2223 = ( n_n4937 ) | ( n_n4933 ) | ( wire249 ) | ( wire16445 ) ;
 assign wire289 = ( wire22  &  n_n518  &  n_n130 ) | ( wire15  &  n_n518  &  n_n130 ) ;
 assign n_n4497 = ( wire22  &  n_n455  &  n_n500 ) ;
 assign wire65 = ( i_9_  &  n_n524  &  n_n455  &  n_n500 ) | ( (~ i_9_)  &  n_n524  &  n_n455  &  n_n500 ) ;
 assign wire66 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign n_n4478 = ( wire13  &  n_n509  &  n_n528 ) ;
 assign n_n4254 = ( n_n4477 ) | ( n_n4475 ) | ( n_n4476 ) ;
 assign wire70 = ( wire21  &  n_n509  &  n_n455 ) | ( wire20  &  n_n509  &  n_n455 ) ;
 assign wire184 = ( wire13  &  n_n509  &  n_n524 ) | ( wire13  &  n_n509  &  n_n526 ) ;
 assign n_n2258 = ( n_n4487 ) | ( n_n4478 ) | ( n_n4254 ) | ( wire16576 ) ;
 assign wire388 = ( n_n4830 ) | ( n_n4831 ) | ( n_n4828 ) | ( wire693 ) ;
 assign n_n2230 = ( wire388 ) | ( wire16351 ) | ( wire16352 ) ;
 assign wire176 = ( i_9_  &  n_n530  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n530  &  n_n518  &  n_n260 ) ;
 assign n_n2229 = ( n_n4843 ) | ( n_n4846 ) | ( wire16355 ) | ( wire16356 ) ;
 assign n_n4822 = ( wire14  &  n_n464  &  n_n520 ) ;
 assign n_n4823 = ( wire23  &  n_n464  &  n_n325 ) ;
 assign n_n4806 = ( wire14  &  n_n473  &  n_n520 ) ;
 assign n_n4820 = ( wire14  &  n_n522  &  n_n464 ) ;
 assign n_n4818 = ( wire14  &  n_n524  &  n_n464 ) ;
 assign n_n4810 = ( wire14  &  n_n464  &  n_n532 ) ;
 assign wire186 = ( wire21  &  n_n464  &  n_n325 ) | ( wire20  &  n_n464  &  n_n325 ) ;
 assign n_n2263 = ( n_n4415 ) | ( n_n4408 ) | ( wire16520 ) | ( wire16521 ) ;
 assign n_n2190 = ( n_n2263 ) | ( wire16526 ) | ( wire16527 ) | ( wire16533 ) ;
 assign n_n2446 = ( n_n4327 ) | ( n_n4324 ) | ( n_n4326 ) ;
 assign n_n4336 = ( wire16  &  n_n526  &  n_n518 ) ;
 assign n_n2443 = ( wire14473 ) | ( wire16  &  n_n522  &  n_n518 ) ;
 assign n_n2445 = ( n_n4331 ) | ( n_n4328 ) | ( n_n4330 ) ;
 assign wire171 = ( wire22  &  n_n536  &  n_n535 ) | ( wire11  &  n_n536  &  n_n535 ) ;
 assign wire198 = ( i_9_  &  n_n536  &  n_n530  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n530  &  n_n518 ) ;
 assign wire283 = ( i_9_  &  n_n536  &  n_n535  &  n_n532 ) | ( (~ i_9_)  &  n_n536  &  n_n535  &  n_n532 ) ;
 assign n_n4379 = ( wire24  &  n_n536  &  n_n491 ) ;
 assign n_n2435 = ( n_n4388 ) | ( n_n4391 ) | ( n_n4390 ) ;
 assign wire54 = ( n_n4386 ) | ( wire12447 ) | ( wire14460 ) ;
 assign wire282 = ( n_n4369 ) | ( n_n4370 ) | ( n_n4368 ) ;
 assign wire423 = ( i_9_  &  n_n536  &  n_n491  &  n_n534 ) | ( (~ i_9_)  &  n_n536  &  n_n491  &  n_n534 ) ;
 assign n_n4503 = ( wire23  &  n_n455  &  n_n500 ) ;
 assign n_n4502 = ( wire13  &  n_n500  &  n_n520 ) ;
 assign n_n4500 = ( wire13  &  n_n522  &  n_n500 ) ;
 assign n_n4546 = ( wire13  &  n_n473  &  n_n524 ) ;
 assign n_n4555 = ( wire24  &  n_n464  &  n_n455 ) ;
 assign wire212 = ( i_9_  &  n_n522  &  n_n473  &  n_n455 ) | ( (~ i_9_)  &  n_n522  &  n_n473  &  n_n455 ) ;
 assign wire213 = ( i_9_  &  n_n464  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n464  &  n_n455  &  n_n528 ) ;
 assign n_n4656 = ( wire10  &  n_n526  &  n_n482 ) ;
 assign n_n4659 = ( wire21  &  n_n390  &  n_n482 ) ;
 assign n_n5106 = ( wire12  &  n_n524  &  n_n518 ) ;
 assign n_n4341 = ( wire20  &  n_n536  &  n_n518 ) ;
 assign n_n5117 = ( wire15  &  n_n509  &  n_n130 ) ;
 assign n_n5223 = ( wire23  &  n_n535  &  n_n65 ) ;
 assign n_n5328 = ( wire19  &  n_n464  &  n_n526 ) ;
 assign n_n5254 = ( wire19  &  n_n509  &  n_n520 ) ;
 assign n_n5249 = ( wire22  &  n_n509  &  n_n65 ) ;
 assign n_n5233 = ( wire22  &  n_n518  &  n_n65 ) ;
 assign n_n5236 = ( wire19  &  n_n522  &  n_n518 ) ;
 assign n_n5262 = ( wire19  &  n_n528  &  n_n500 ) ;
 assign n_n5278 = ( wire19  &  n_n528  &  n_n491 ) ;
 assign wire449 = ( i_9_  &  n_n526  &  n_n535  &  n_n65 ) | ( (~ i_9_)  &  n_n526  &  n_n535  &  n_n65 ) ;
 assign n_n2083 = ( wire16774 ) | ( wire16775 ) | ( wire16776 ) | ( wire16777 ) ;
 assign n_n4375 = ( wire23  &  n_n536  &  n_n500 ) ;
 assign n_n4436 = ( wire16  &  n_n522  &  n_n464 ) ;
 assign n_n4833 = ( wire22  &  n_n535  &  n_n260 ) ;
 assign n_n4875 = ( wire24  &  n_n500  &  n_n260 ) ;
 assign n_n4940 = ( wire17  &  n_n464  &  n_n530 ) ;
 assign n_n4939 = ( wire24  &  n_n464  &  n_n260 ) ;
 assign n_n4729 = ( wire25  &  n_n509  &  n_n325 ) ;
 assign n_n4728 = ( wire14  &  n_n509  &  n_n534 ) ;
 assign wire373 = ( i_9_  &  n_n509  &  n_n520  &  n_n325 ) | ( (~ i_9_)  &  n_n509  &  n_n520  &  n_n325 ) ;
 assign wire374 = ( i_9_  &  n_n509  &  n_n522  &  n_n325 ) | ( (~ i_9_)  &  n_n509  &  n_n522  &  n_n325 ) ;
 assign n_n5132 = ( wire12  &  n_n500  &  n_n530 ) ;
 assign n_n5128 = ( wire12  &  n_n500  &  n_n534 ) ;
 assign n_n5016 = ( wire18  &  n_n491  &  n_n534 ) ;
 assign n_n4129 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) ;
 assign n_n5306 = ( wire19  &  n_n473  &  n_n532 ) ;
 assign n_n3019 = ( n_n5307 ) | ( n_n5306 ) | ( n_n5308 ) ;
 assign n_n5009 = ( wire22  &  n_n500  &  n_n195 ) ;
 assign n_n5335 = ( wire23  &  n_n464  &  n_n65 ) ;
 assign n_n4562 = ( wire13  &  n_n524  &  n_n464 ) ;
 assign n_n4506 = ( wire13  &  n_n491  &  n_n532 ) ;
 assign n_n4492 = ( wire13  &  n_n500  &  n_n530 ) ;
 assign n_n1338 = ( n_n4580 ) | ( n_n4635 ) | ( wire12047 ) | ( wire12048 ) ;
 assign n_n4496 = ( wire13  &  n_n526  &  n_n500 ) ;
 assign n_n4535 = ( wire23  &  n_n455  &  n_n482 ) ;
 assign n_n1326 = ( n_n1338 ) | ( wire12053 ) | ( wire12054 ) | ( wire12062 ) ;
 assign n_n1336 = ( n_n4732 ) | ( n_n4743 ) | ( wire12067 ) | ( wire12068 ) ;
 assign n_n4788 = ( wire14  &  n_n522  &  n_n482 ) ;
 assign n_n1325 = ( n_n1336 ) | ( wire12074 ) | ( wire12075 ) | ( wire12083 ) ;
 assign n_n4342 = ( wire16  &  n_n520  &  n_n518 ) ;
 assign n_n4608 = ( wire10  &  n_n509  &  n_n526 ) ;
 assign n_n4610 = ( wire10  &  n_n509  &  n_n524 ) ;
 assign n_n4606 = ( wire10  &  n_n509  &  n_n528 ) ;
 assign n_n4675 = ( wire21  &  n_n473  &  n_n390 ) ;
 assign n_n4676 = ( wire10  &  n_n522  &  n_n473 ) ;
 assign n_n4674 = ( wire10  &  n_n473  &  n_n524 ) ;
 assign n_n4730 = ( wire14  &  n_n509  &  n_n532 ) ;
 assign n_n4802 = ( wire14  &  n_n473  &  n_n524 ) ;
 assign n_n4851 = ( wire21  &  n_n518  &  n_n260 ) ;
 assign n_n4852 = ( wire17  &  n_n522  &  n_n518 ) ;
 assign n_n4914 = ( wire17  &  n_n524  &  n_n482 ) ;
 assign n_n4962 = ( wire18  &  n_n524  &  n_n535 ) ;
 assign n_n4956 = ( wire18  &  n_n535  &  n_n530 ) ;
 assign n_n5020 = ( wire18  &  n_n491  &  n_n530 ) ;
 assign n_n5064 = ( wire18  &  n_n464  &  n_n534 ) ;
 assign n_n5189 = ( wire20  &  n_n473  &  n_n130 ) ;
 assign n_n5190 = ( wire12  &  n_n473  &  n_n520 ) ;
 assign n_n5188 = ( wire12  &  n_n522  &  n_n473 ) ;
 assign n_n4352 = ( wire16  &  n_n509  &  n_n526 ) ;
 assign n_n4351 = ( wire11  &  n_n509  &  n_n536 ) ;
 assign n_n4356 = ( wire16  &  n_n509  &  n_n522 ) ;
 assign wire67 = ( i_9_  &  n_n509  &  n_n536  &  n_n532 ) | ( (~ i_9_)  &  n_n509  &  n_n536  &  n_n532 ) ;
 assign n_n1120 = ( n_n4352 ) | ( n_n4351 ) | ( wire11610 ) | ( wire11611 ) ;
 assign n_n4507 = ( wire24  &  n_n455  &  n_n491 ) ;
 assign n_n4509 = ( wire15  &  n_n455  &  n_n491 ) ;
 assign n_n4508 = ( wire13  &  n_n491  &  n_n530 ) ;
 assign wire129 = ( i_9_  &  n_n526  &  n_n455  &  n_n491 ) | ( (~ i_9_)  &  n_n526  &  n_n455  &  n_n491 ) ;
 assign wire308 = ( i_9_  &  n_n455  &  n_n528  &  n_n491 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n491 ) ;
 assign n_n4622 = ( wire10  &  n_n528  &  n_n500 ) ;
 assign n_n4621 = ( wire15  &  n_n500  &  n_n390 ) ;
 assign wire75 = ( wire10  &  n_n526  &  n_n500 ) ;
 assign n_n3861 = ( n_n4622 ) | ( n_n4621 ) | ( wire75 ) ;
 assign n_n5073 = ( wire22  &  n_n464  &  n_n195 ) ;
 assign n_n5074 = ( wire18  &  n_n524  &  n_n464 ) ;
 assign n_n5072 = ( wire18  &  n_n464  &  n_n526 ) ;
 assign n_n4152 = ( n_n5073 ) | ( n_n5074 ) | ( n_n5072 ) ;
 assign n_n4931 = ( wire21  &  n_n473  &  n_n260 ) ;
 assign wire180 = ( i_9_  &  n_n473  &  n_n520  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n520  &  n_n260 ) ;
 assign wire382 = ( i_9_  &  n_n522  &  n_n473  &  n_n260 ) | ( (~ i_9_)  &  n_n522  &  n_n473  &  n_n260 ) ;
 assign n_n4978 = ( wire18  &  n_n524  &  n_n518 ) ;
 assign n_n4980 = ( wire18  &  n_n522  &  n_n518 ) ;
 assign n_n4897 = ( wire22  &  n_n491  &  n_n260 ) ;
 assign n_n1077 = ( n_n4877 ) | ( n_n1985 ) | ( n_n3815 ) | ( wire11818 ) ;
 assign wire264 = ( wire17  &  n_n528  &  n_n491 ) | ( wire17  &  n_n491  &  n_n530 ) ;
 assign n_n4349 = ( wire15  &  n_n509  &  n_n536 ) ;
 assign n_n4350 = ( wire16  &  n_n509  &  n_n528 ) ;
 assign n_n4348 = ( wire16  &  n_n509  &  n_n530 ) ;
 assign n_n1002 = ( n_n4349 ) | ( n_n4350 ) | ( n_n4348 ) ;
 assign n_n5172 = ( wire12  &  n_n522  &  n_n482 ) ;
 assign n_n4580 = ( wire10  &  n_n522  &  n_n535 ) ;
 assign n_n4357 = ( wire20  &  n_n509  &  n_n536 ) ;
 assign n_n4419 = ( wire21  &  n_n536  &  n_n473 ) ;
 assign n_n4605 = ( wire15  &  n_n509  &  n_n390 ) ;
 assign n_n4655 = ( wire11  &  n_n390  &  n_n482 ) ;
 assign n_n4661 = ( wire20  &  n_n390  &  n_n482 ) ;
 assign n_n4683 = ( wire24  &  n_n464  &  n_n390 ) ;
 assign n_n4689 = ( wire22  &  n_n464  &  n_n390 ) ;
 assign n_n4697 = ( wire25  &  n_n535  &  n_n325 ) ;
 assign n_n4703 = ( wire11  &  n_n535  &  n_n325 ) ;
 assign n_n4712 = ( wire14  &  n_n534  &  n_n518 ) ;
 assign n_n4718 = ( wire14  &  n_n528  &  n_n518 ) ;
 assign n_n4763 = ( wire24  &  n_n491  &  n_n325 ) ;
 assign n_n4778 = ( wire14  &  n_n482  &  n_n532 ) ;
 assign n_n4886 = ( wire17  &  n_n500  &  n_n520 ) ;
 assign n_n4915 = ( wire21  &  n_n482  &  n_n260 ) ;
 assign n_n4989 = ( wire15  &  n_n509  &  n_n195 ) ;
 assign n_n5011 = ( wire21  &  n_n500  &  n_n195 ) ;
 assign n_n5061 = ( wire20  &  n_n473  &  n_n195 ) ;
 assign n_n5070 = ( wire18  &  n_n464  &  n_n528 ) ;
 assign n_n5076 = ( wire18  &  n_n522  &  n_n464 ) ;
 assign n_n5135 = ( wire11  &  n_n500  &  n_n130 ) ;
 assign n_n5157 = ( wire20  &  n_n491  &  n_n130 ) ;
 assign n_n5201 = ( wire22  &  n_n464  &  n_n130 ) ;
 assign n_n5207 = ( wire23  &  n_n464  &  n_n130 ) ;
 assign n_n5237 = ( wire20  &  n_n518  &  n_n65 ) ;
 assign n_n5252 = ( wire19  &  n_n509  &  n_n522 ) ;
 assign n_n4353 = ( wire22  &  n_n509  &  n_n536 ) ;
 assign n_n4456 = ( wire13  &  n_n534  &  n_n518 ) ;
 assign n_n4458 = ( wire13  &  n_n532  &  n_n518 ) ;
 assign n_n4671 = ( wire11  &  n_n473  &  n_n390 ) ;
 assign n_n4747 = ( wire24  &  n_n500  &  n_n325 ) ;
 assign n_n4772 = ( wire14  &  n_n522  &  n_n491 ) ;
 assign n_n4773 = ( wire20  &  n_n491  &  n_n325 ) ;
 assign n_n4771 = ( wire21  &  n_n491  &  n_n325 ) ;
 assign n_n4205 = ( wire12393 ) | ( wire21  &  n_n491  &  n_n325 ) ;
 assign n_n5023 = ( wire11  &  n_n491  &  n_n195 ) ;
 assign n_n5024 = ( wire18  &  n_n526  &  n_n491 ) ;
 assign n_n5082 = ( wire12  &  n_n535  &  n_n532 ) ;
 assign n_n5084 = ( wire12  &  n_n535  &  n_n530 ) ;
 assign n_n5275 = ( wire24  &  n_n491  &  n_n65 ) ;
 assign n_n5276 = ( wire19  &  n_n491  &  n_n530 ) ;
 assign n_n4600 = ( wire10  &  n_n509  &  n_n534 ) ;
 assign wire45 = ( i_9_  &  n_n520  &  n_n390  &  n_n518 ) | ( (~ i_9_)  &  n_n520  &  n_n390  &  n_n518 ) ;
 assign n_n4204 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4775 ) ;
 assign n_n4010 = ( n_n4065 ) | ( wire13162 ) | ( wire13163 ) | ( wire13166 ) ;
 assign n_n4009 = ( wire13176 ) | ( wire13177 ) | ( wire13178 ) | ( wire13181 ) ;
 assign n_n3990 = ( wire13228 ) | ( wire13229 ) | ( wire13233 ) | ( wire13236 ) ;
 assign n_n4753 = ( wire22  &  n_n500  &  n_n325 ) ;
 assign n_n4752 = ( wire14  &  n_n526  &  n_n500 ) ;
 assign n_n4013 = ( n_n4075 ) | ( wire13249 ) | ( wire13250 ) | ( wire13254 ) ;
 assign wire47 = ( wire14  &  n_n500  &  n_n532 ) | ( wire14  &  n_n500  &  n_n534 ) ;
 assign n_n3992 = ( n_n4013 ) | ( wire13269 ) | ( wire13270 ) | ( wire13278 ) ;
 assign n_n4457 = ( wire25  &  n_n455  &  n_n518 ) ;
 assign n_n5075 = ( wire21  &  n_n464  &  n_n195 ) ;
 assign n_n5079 = ( wire23  &  n_n464  &  n_n195 ) ;
 assign n_n5088 = ( wire12  &  n_n526  &  n_n535 ) ;
 assign n_n5078 = ( wire18  &  n_n464  &  n_n520 ) ;
 assign n_n5083 = ( wire24  &  n_n535  &  n_n130 ) ;
 assign wire123 = ( i_9_  &  n_n535  &  n_n530  &  n_n130 ) | ( (~ i_9_)  &  n_n535  &  n_n530  &  n_n130 ) ;
 assign wire122 = ( wire24  &  n_n518  &  n_n130 ) | ( wire15  &  n_n518  &  n_n130 ) ;
 assign wire232 = ( i_9_  &  n_n524  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n130 ) ;
 assign n_n5063 = ( wire23  &  n_n473  &  n_n195 ) ;
 assign n_n5058 = ( wire18  &  n_n473  &  n_n524 ) ;
 assign wire160 = ( wire18  &  n_n464  &  n_n530 ) | ( wire18  &  n_n464  &  n_n532 ) ;
 assign n_n3558 = ( n_n4891 ) | ( n_n4836 ) | ( wire14260 ) | ( wire14261 ) ;
 assign n_n3557 = ( wire14267 ) | ( wire14268 ) ;
 assign n_n4409 = ( wire25  &  n_n536  &  n_n473 ) ;
 assign n_n4399 = ( wire11  &  n_n536  &  n_n482 ) ;
 assign n_n4370 = ( wire16  &  n_n524  &  n_n500 ) ;
 assign n_n3548 = ( n_n3560 ) | ( n_n3561 ) | ( wire14332 ) ;
 assign n_n4505 = ( wire25  &  n_n455  &  n_n491 ) ;
 assign n_n5095 = ( wire23  &  n_n535  &  n_n130 ) ;
 assign n_n5158 = ( wire12  &  n_n491  &  n_n520 ) ;
 assign n_n5154 = ( wire12  &  n_n524  &  n_n491 ) ;
 assign n_n4775 = ( wire23  &  n_n491  &  n_n325 ) ;
 assign n_n4780 = ( wire14  &  n_n530  &  n_n482 ) ;
 assign n_n3469 = ( n_n4770 ) | ( n_n4773 ) | ( n_n4771 ) ;
 assign n_n5013 = ( wire20  &  n_n500  &  n_n195 ) ;
 assign n_n5150 = ( wire12  &  n_n528  &  n_n491 ) ;
 assign n_n5147 = ( wire24  &  n_n491  &  n_n130 ) ;
 assign wire76 = ( i_9_  &  n_n491  &  n_n530  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n530  &  n_n130 ) ;
 assign wire196 = ( i_9_  &  n_n526  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n130 ) ;
 assign wire57 = ( i_9_  &  n_n524  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n195 ) ;
 assign wire251 = ( i_9_  &  n_n520  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n520  &  n_n518  &  n_n195 ) ;
 assign n_n4948 = ( wire17  &  n_n522  &  n_n464 ) ;
 assign n_n4957 = ( wire15  &  n_n535  &  n_n195 ) ;
 assign n_n4971 = ( wire24  &  n_n518  &  n_n195 ) ;
 assign wire342 = ( i_9_  &  n_n524  &  n_n535  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n195 ) ;
 assign n_n4488 = ( wire13  &  n_n500  &  n_n534 ) ;
 assign n_n4471 = ( wire23  &  n_n455  &  n_n518 ) ;
 assign n_n4490 = ( wire13  &  n_n500  &  n_n532 ) ;
 assign n_n901 = ( n_n4478 ) | ( n_n4477 ) | ( n_n4479 ) ;
 assign n_n3358 = ( n_n4460 ) | ( n_n4457 ) | ( wire14120 ) | ( wire14121 ) ;
 assign n_n3285 = ( n_n3358 ) | ( wire14126 ) | ( wire14127 ) | ( wire14131 ) ;
 assign n_n4423 = ( wire23  &  n_n536  &  n_n473 ) ;
 assign n_n4421 = ( wire20  &  n_n536  &  n_n473 ) ;
 assign wire84 = ( i_9_  &  n_n536  &  n_n464  &  n_n532 ) | ( (~ i_9_)  &  n_n536  &  n_n464  &  n_n532 ) ;
 assign wire470 = ( n_n4445 ) | ( n_n4444 ) | ( n_n4446 ) ;
 assign n_n4635 = ( wire24  &  n_n491  &  n_n390 ) ;
 assign n_n4630 = ( wire10  &  n_n500  &  n_n520 ) ;
 assign n_n5065 = ( wire25  &  n_n464  &  n_n195 ) ;
 assign n_n5287 = ( wire23  &  n_n491  &  n_n65 ) ;
 assign n_n5281 = ( wire22  &  n_n491  &  n_n65 ) ;
 assign n_n5268 = ( wire19  &  n_n522  &  n_n500 ) ;
 assign n_n5261 = ( wire15  &  n_n500  &  n_n65 ) ;
 assign n_n3194 = ( n_n5281 ) | ( n_n5268 ) | ( wire13709 ) | ( wire13710 ) ;
 assign n_n4331 = ( wire24  &  n_n536  &  n_n518 ) ;
 assign n_n4332 = ( wire16  &  n_n530  &  n_n518 ) ;
 assign n_n4329 = ( wire25  &  n_n536  &  n_n518 ) ;
 assign n_n4448 = ( wire13  &  n_n526  &  n_n535 ) ;
 assign n_n4449 = ( wire22  &  n_n455  &  n_n535 ) ;
 assign n_n4447 = ( wire11  &  n_n455  &  n_n535 ) ;
 assign n_n4870 = ( wire17  &  n_n509  &  n_n520 ) ;
 assign n_n5029 = ( wire20  &  n_n491  &  n_n195 ) ;
 assign n_n3162 = ( n_n4467 ) | ( n_n4466 ) | ( n_n4468 ) ;
 assign n_n4472 = ( wire13  &  n_n509  &  n_n534 ) ;
 assign n_n4469 = ( wire20  &  n_n455  &  n_n518 ) ;
 assign n_n4477 = ( wire15  &  n_n509  &  n_n455 ) ;
 assign n_n4475 = ( wire24  &  n_n509  &  n_n455 ) ;
 assign n_n4479 = ( wire11  &  n_n509  &  n_n455 ) ;
 assign n_n4474 = ( wire13  &  n_n509  &  n_n532 ) ;
 assign n_n3001 = ( n_n3162 ) | ( n_n4479 ) | ( n_n4474 ) | ( wire15423 ) ;
 assign wire465 = ( i_9_  &  n_n509  &  n_n520  &  n_n390 ) | ( (~ i_9_)  &  n_n509  &  n_n520  &  n_n390 ) ;
 assign n_n4620 = ( wire10  &  n_n500  &  n_n530 ) ;
 assign n_n5001 = ( wire25  &  n_n500  &  n_n195 ) ;
 assign n_n2548 = ( n_n2601 ) | ( n_n2602 ) | ( wire14904 ) | ( wire14905 ) ;
 assign n_n4867 = ( wire21  &  n_n509  &  n_n260 ) ;
 assign n_n4866 = ( wire17  &  n_n509  &  n_n524 ) ;
 assign n_n2597 = ( n_n3450 ) | ( n_n4889 ) | ( wire12179 ) | ( wire14912 ) ;
 assign n_n4863 = ( wire11  &  n_n509  &  n_n260 ) ;
 assign n_n2727 = ( n_n4859 ) | ( n_n4860 ) | ( n_n4861 ) ;
 assign n_n2549 = ( n_n2604 ) | ( wire14922 ) | ( wire14923 ) | ( wire14927 ) ;
 assign n_n4965 = ( wire20  &  n_n535  &  n_n195 ) ;
 assign wire228 = ( i_9_  &  n_n526  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n195 ) ;
 assign n_n2551 = ( n_n2611 ) | ( wire15011 ) | ( wire15012 ) | ( wire15016 ) ;
 assign wire315 = ( i_9_  &  n_n482  &  n_n534  &  n_n325 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n325 ) ;
 assign n_n4321 = ( wire22  &  n_n536  &  n_n535 ) ;
 assign n_n4417 = ( wire22  &  n_n536  &  n_n473 ) ;
 assign n_n4415 = ( wire11  &  n_n536  &  n_n473 ) ;
 assign n_n4972 = ( wire18  &  n_n530  &  n_n518 ) ;
 assign n_n5118 = ( wire12  &  n_n509  &  n_n528 ) ;
 assign n_n5119 = ( wire11  &  n_n509  &  n_n130 ) ;
 assign n_n5229 = ( wire15  &  n_n518  &  n_n65 ) ;
 assign n_n5228 = ( wire19  &  n_n530  &  n_n518 ) ;
 assign n_n5295 = ( wire11  &  n_n482  &  n_n65 ) ;
 assign n_n4540 = ( wire13  &  n_n473  &  n_n530 ) ;
 assign n_n4536 = ( wire13  &  n_n473  &  n_n534 ) ;
 assign n_n4532 = ( wire13  &  n_n522  &  n_n482 ) ;
 assign n_n4541 = ( wire15  &  n_n473  &  n_n455 ) ;
 assign wire416 = ( i_9_  &  n_n473  &  n_n455  &  n_n528 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n528 ) ;
 assign n_n4681 = ( wire25  &  n_n464  &  n_n390 ) ;
 assign n_n4679 = ( wire23  &  n_n473  &  n_n390 ) ;
 assign n_n4677 = ( wire20  &  n_n473  &  n_n390 ) ;
 assign n_n4678 = ( wire10  &  n_n473  &  n_n520 ) ;
 assign wire81 = ( wire10  &  n_n464  &  n_n532 ) ;
 assign n_n2242 = ( n_n4677 ) | ( n_n4678 ) | ( wire16404 ) | ( wire16405 ) ;
 assign wire414 = ( i_9_  &  n_n509  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n130 ) ;
 assign wire345 = ( wire16  &  n_n500  &  n_n532 ) | ( wire16  &  n_n500  &  n_n534 ) ;
 assign wire164 = ( i_9_  &  n_n526  &  n_n491  &  n_n325 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n325 ) ;
 assign n_n4465 = ( wire22  &  n_n455  &  n_n518 ) ;
 assign n_n4443 = ( wire24  &  n_n455  &  n_n535 ) ;
 assign n_n5121 = ( wire22  &  n_n509  &  n_n130 ) ;
 assign n_n5122 = ( wire12  &  n_n509  &  n_n524 ) ;
 assign n_n4486 = ( wire13  &  n_n509  &  n_n520 ) ;
 assign n_n4484 = ( wire13  &  n_n509  &  n_n522 ) ;
 assign wire199 = ( wire22  &  n_n509  &  n_n455 ) | ( wire11  &  n_n509  &  n_n455 ) ;
 assign n_n4865 = ( wire22  &  n_n509  &  n_n260 ) ;
 assign n_n4893 = ( wire15  &  n_n491  &  n_n260 ) ;
 assign wire154 = ( i_9_  &  n_n482  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n260 ) ;
 assign n_n2095 = ( wire16784 ) | ( wire16785 ) ;
 assign n_n5168 = ( wire12  &  n_n526  &  n_n482 ) ;
 assign n_n2091 = ( n_n5193 ) | ( n_n5182 ) | ( wire16795 ) | ( wire16796 ) ;
 assign n_n4973 = ( wire15  &  n_n518  &  n_n195 ) ;
 assign n_n2084 = ( n_n2091 ) | ( wire16790 ) | ( wire16791 ) | ( wire16805 ) ;
 assign n_n4378 = ( wire16  &  n_n491  &  n_n532 ) ;
 assign n_n4377 = ( wire25  &  n_n536  &  n_n491 ) ;
 assign n_n4710 = ( wire14  &  n_n535  &  n_n520 ) ;
 assign n_n4709 = ( wire20  &  n_n535  &  n_n325 ) ;
 assign n_n4765 = ( wire15  &  n_n491  &  n_n325 ) ;
 assign n_n4603 = ( wire24  &  n_n509  &  n_n390 ) ;
 assign n_n4604 = ( wire10  &  n_n509  &  n_n530 ) ;
 assign n_n2037 = ( n_n4600 ) | ( n_n4603 ) | ( n_n4604 ) ;
 assign n_n4588 = ( wire10  &  n_n530  &  n_n518 ) ;
 assign n_n4595 = ( wire21  &  n_n390  &  n_n518 ) ;
 assign n_n1877 = ( n_n2037 ) | ( n_n4588 ) | ( n_n4595 ) | ( wire16038 ) ;
 assign n_n1450 = ( n_n5067 ) | ( n_n5061 ) | ( wire12309 ) | ( wire12310 ) ;
 assign n_n5152 = ( wire12  &  n_n526  &  n_n491 ) ;
 assign n_n5149 = ( wire15  &  n_n491  &  n_n130 ) ;
 assign wire195 = ( i_9_  &  n_n491  &  n_n520  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n130 ) ;
 assign wire358 = ( i_9_  &  n_n524  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n491  &  n_n130 ) ;
 assign wire406 = ( i_9_  &  n_n528  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n528  &  n_n491  &  n_n130 ) ;
 assign n_n5288 = ( wire19  &  n_n482  &  n_n534 ) ;
 assign n_n4743 = ( wire23  &  n_n509  &  n_n325 ) ;
 assign n_n4751 = ( wire11  &  n_n500  &  n_n325 ) ;
 assign n_n1333 = ( n_n4971 ) | ( n_n4972 ) | ( wire12122 ) | ( wire12123 ) ;
 assign n_n4386 = ( wire16  &  n_n524  &  n_n491 ) ;
 assign n_n4435 = ( wire21  &  n_n536  &  n_n464 ) ;
 assign n_n4626 = ( wire10  &  n_n524  &  n_n500 ) ;
 assign n_n4627 = ( wire21  &  n_n500  &  n_n390 ) ;
 assign n_n4625 = ( wire22  &  n_n500  &  n_n390 ) ;
 assign n_n4660 = ( wire10  &  n_n522  &  n_n482 ) ;
 assign n_n4719 = ( wire11  &  n_n325  &  n_n518 ) ;
 assign n_n4717 = ( wire15  &  n_n325  &  n_n518 ) ;
 assign n_n4954 = ( wire18  &  n_n535  &  n_n532 ) ;
 assign n_n4955 = ( wire24  &  n_n535  &  n_n195 ) ;
 assign n_n5133 = ( wire15  &  n_n500  &  n_n130 ) ;
 assign n_n5138 = ( wire12  &  n_n524  &  n_n500 ) ;
 assign n_n5139 = ( wire21  &  n_n500  &  n_n130 ) ;
 assign n_n5309 = ( wire15  &  n_n473  &  n_n65 ) ;
 assign n_n5308 = ( wire19  &  n_n473  &  n_n530 ) ;
 assign n_n1128 = ( n_n5310 ) | ( n_n5309 ) | ( n_n5308 ) ;
 assign n_n4387 = ( wire21  &  n_n536  &  n_n491 ) ;
 assign wire420 = ( wire22  &  n_n536  &  n_n491 ) | ( wire11  &  n_n536  &  n_n491 ) ;
 assign n_n4619 = ( wire24  &  n_n500  &  n_n390 ) ;
 assign wire179 = ( i_9_  &  n_n473  &  n_n532  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n325 ) ;
 assign n_n4750 = ( wire14  &  n_n528  &  n_n500 ) ;
 assign n_n4745 = ( wire25  &  n_n500  &  n_n325 ) ;
 assign n_n4736 = ( wire14  &  n_n509  &  n_n526 ) ;
 assign wire293 = ( wire21  &  n_n509  &  n_n325 ) | ( wire20  &  n_n509  &  n_n325 ) ;
 assign wire457 = ( n_n4720 ) | ( n_n4722 ) | ( n_n4721 ) ;
 assign n_n5159 = ( wire23  &  n_n491  &  n_n130 ) ;
 assign n_n5160 = ( wire12  &  n_n482  &  n_n534 ) ;
 assign wire287 = ( i_9_  &  n_n522  &  n_n491  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n491  &  n_n130 ) ;
 assign n_n5169 = ( wire22  &  n_n482  &  n_n130 ) ;
 assign wire33 = ( i_9_  &  n_n530  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n530  &  n_n482  &  n_n130 ) ;
 assign wire107 = ( i_9_  &  n_n524  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n482  &  n_n130 ) ;
 assign wire113 = ( i_9_  &  n_n473  &  n_n526  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n526  &  n_n130 ) ;
 assign wire254 = ( i_9_  &  n_n528  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n528  &  n_n482  &  n_n130 ) ;
 assign n_n4658 = ( wire10  &  n_n524  &  n_n482 ) ;
 assign n_n5108 = ( wire12  &  n_n522  &  n_n518 ) ;
 assign n_n4510 = ( wire13  &  n_n528  &  n_n491 ) ;
 assign n_n4355 = ( wire21  &  n_n509  &  n_n536 ) ;
 assign n_n4424 = ( wire16  &  n_n464  &  n_n534 ) ;
 assign n_n4498 = ( wire13  &  n_n524  &  n_n500 ) ;
 assign n_n4591 = ( wire11  &  n_n390  &  n_n518 ) ;
 assign n_n4663 = ( wire23  &  n_n390  &  n_n482 ) ;
 assign n_n4698 = ( wire14  &  n_n535  &  n_n532 ) ;
 assign n_n4705 = ( wire22  &  n_n535  &  n_n325 ) ;
 assign n_n4805 = ( wire20  &  n_n473  &  n_n325 ) ;
 assign n_n4841 = ( wire25  &  n_n518  &  n_n260 ) ;
 assign n_n4944 = ( wire17  &  n_n464  &  n_n526 ) ;
 assign n_n5068 = ( wire18  &  n_n464  &  n_n530 ) ;
 assign n_n5187 = ( wire21  &  n_n473  &  n_n130 ) ;
 assign n_n5199 = ( wire11  &  n_n464  &  n_n130 ) ;
 assign n_n5260 = ( wire19  &  n_n500  &  n_n530 ) ;
 assign n_n5272 = ( wire19  &  n_n491  &  n_n534 ) ;
 assign n_n4405 = ( wire20  &  n_n536  &  n_n482 ) ;
 assign n_n4406 = ( wire16  &  n_n520  &  n_n482 ) ;
 assign n_n4462 = ( wire13  &  n_n528  &  n_n518 ) ;
 assign n_n4501 = ( wire20  &  n_n455  &  n_n500 ) ;
 assign n_n4684 = ( wire10  &  n_n464  &  n_n530 ) ;
 assign n_n4222 = ( n_n4683 ) | ( wire81 ) | ( n_n4684 ) ;
 assign n_n4741 = ( wire20  &  n_n509  &  n_n325 ) ;
 assign n_n4740 = ( wire14  &  n_n509  &  n_n522 ) ;
 assign n_n4819 = ( wire21  &  n_n464  &  n_n325 ) ;
 assign n_n5077 = ( wire20  &  n_n464  &  n_n195 ) ;
 assign n_n5221 = ( wire20  &  n_n535  &  n_n65 ) ;
 assign n_n5220 = ( wire19  &  n_n522  &  n_n535 ) ;
 assign n_n834 = ( n_n4849 ) | ( n_n4850 ) | ( n_n4848 ) ;
 assign n_n5134 = ( wire12  &  n_n528  &  n_n500 ) ;
 assign n_n5125 = ( wire20  &  n_n509  &  n_n130 ) ;
 assign wire336 = ( wire12  &  n_n509  &  n_n522 ) | ( wire12  &  n_n509  &  n_n520 ) ;
 assign n_n3988 = ( wire13322 ) | ( wire13323 ) | ( wire13325 ) | ( wire13327 ) ;
 assign n_n5290 = ( wire19  &  n_n482  &  n_n532 ) ;
 assign n_n5291 = ( wire24  &  n_n482  &  n_n65 ) ;
 assign n_n5292 = ( wire19  &  n_n530  &  n_n482 ) ;
 assign n_n4026 = ( n_n5303 ) | ( n_n1128 ) | ( n_n5304 ) | ( wire13329 ) ;
 assign n_n3998 = ( n_n4030 ) | ( n_n4031 ) | ( wire13346 ) | ( wire13347 ) ;
 assign wire441 = ( i_9_  &  n_n522  &  n_n491  &  n_n65 ) | ( (~ i_9_)  &  n_n522  &  n_n491  &  n_n65 ) ;
 assign n_n3987 = ( n_n3998 ) | ( wire13364 ) | ( wire13365 ) | ( wire13374 ) ;
 assign n_n4410 = ( wire16  &  n_n473  &  n_n532 ) ;
 assign n_n4652 = ( wire10  &  n_n530  &  n_n482 ) ;
 assign n_n4650 = ( wire10  &  n_n482  &  n_n532 ) ;
 assign n_n3681 = ( n_n5045 ) | ( n_n5053 ) | ( wire14658 ) | ( wire14659 ) ;
 assign wire97 = ( i_9_  &  n_n526  &  n_n482  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n482  &  n_n195 ) ;
 assign n_n3639 = ( n_n3681 ) | ( wire14661 ) | ( wire14662 ) | ( wire14667 ) ;
 assign wire159 = ( wire11  &  n_n464  &  n_n195 ) | ( wire24  &  n_n464  &  n_n195 ) ;
 assign n_n5226 = ( wire19  &  n_n532  &  n_n518 ) ;
 assign n_n5218 = ( wire19  &  n_n524  &  n_n535 ) ;
 assign wire435 = ( wire19  &  n_n509  &  n_n522 ) | ( wire19  &  n_n509  &  n_n524 ) ;
 assign n_n5153 = ( wire22  &  n_n491  &  n_n130 ) ;
 assign n_n5021 = ( wire15  &  n_n491  &  n_n195 ) ;
 assign n_n4654 = ( wire10  &  n_n528  &  n_n482 ) ;
 assign wire140 = ( i_9_  &  n_n390  &  n_n482  &  n_n532 ) | ( (~ i_9_)  &  n_n390  &  n_n482  &  n_n532 ) ;
 assign wire391 = ( i_9_  &  n_n526  &  n_n390  &  n_n482 ) | ( (~ i_9_)  &  n_n526  &  n_n390  &  n_n482 ) ;
 assign n_n4665 = ( wire25  &  n_n473  &  n_n390 ) ;
 assign wire72 = ( wire21  &  n_n390  &  n_n482 ) | ( wire20  &  n_n390  &  n_n482 ) ;
 assign wire418 = ( i_9_  &  n_n464  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n464  &  n_n390  &  n_n534 ) ;
 assign wire248 = ( wire21  &  n_n509  &  n_n195 ) | ( wire20  &  n_n509  &  n_n195 ) ;
 assign n_n4368 = ( wire16  &  n_n526  &  n_n500 ) ;
 assign n_n4394 = ( wire16  &  n_n482  &  n_n532 ) ;
 assign n_n3363 = ( n_n4407 ) | ( n_n4404 ) | ( wire14168 ) | ( wire14169 ) ;
 assign n_n3362 = ( n_n4415 ) | ( n_n4408 ) | ( wire14173 ) | ( wire14174 ) ;
 assign n_n3287 = ( n_n3363 ) | ( n_n3362 ) | ( wire14178 ) | ( wire14179 ) ;
 assign n_n3369 = ( n_n4324 ) | ( n_n4335 ) | ( n_n4279 ) | ( wire14183 ) ;
 assign n_n3370 = ( n_n4319 ) | ( n_n4320 ) | ( wire363 ) | ( wire14186 ) ;
 assign wire156 = ( i_9_  &  n_n536  &  n_n520  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n520  &  n_n518 ) ;
 assign n_n3262 = ( n_n3287 ) | ( wire14163 ) | ( wire14164 ) | ( wire14195 ) ;
 assign n_n4891 = ( wire24  &  n_n491  &  n_n260 ) ;
 assign n_n4896 = ( wire17  &  n_n526  &  n_n491 ) ;
 assign n_n4428 = ( wire16  &  n_n464  &  n_n530 ) ;
 assign wire403 = ( wire13  &  n_n532  &  n_n518 ) | ( wire13  &  n_n534  &  n_n518 ) ;
 assign n_n4499 = ( wire21  &  n_n455  &  n_n500 ) ;
 assign n_n4545 = ( wire22  &  n_n473  &  n_n455 ) ;
 assign wire471 = ( i_9_  &  n_n522  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n455 ) ;
 assign n_n4326 = ( wire16  &  n_n535  &  n_n520 ) ;
 assign n_n4328 = ( wire16  &  n_n534  &  n_n518 ) ;
 assign n_n4376 = ( wire16  &  n_n491  &  n_n534 ) ;
 assign n_n3176 = ( wire423 ) | ( wire16  &  n_n491  &  n_n532 ) ;
 assign n_n4585 = ( wire25  &  n_n390  &  n_n518 ) ;
 assign n_n4873 = ( wire25  &  n_n500  &  n_n260 ) ;
 assign n_n4932 = ( wire17  &  n_n522  &  n_n473 ) ;
 assign n_n4592 = ( wire10  &  n_n526  &  n_n518 ) ;
 assign n_n5052 = ( wire18  &  n_n473  &  n_n530 ) ;
 assign n_n2956 = ( n_n5047 ) | ( n_n5051 ) | ( wire15601 ) | ( wire15602 ) ;
 assign n_n5235 = ( wire21  &  n_n518  &  n_n65 ) ;
 assign n_n5234 = ( wire19  &  n_n524  &  n_n518 ) ;
 assign n_n5286 = ( wire19  &  n_n491  &  n_n520 ) ;
 assign n_n5285 = ( wire20  &  n_n491  &  n_n65 ) ;
 assign n_n1764 = ( n_n4667 ) | ( n_n4664 ) | ( n_n4663 ) ;
 assign n_n3810 = ( n_n4898 ) | ( n_n4897 ) | ( n_n4896 ) ;
 assign n_n2304 = ( n_n5130 ) | ( n_n5133 ) | ( n_n5134 ) ;
 assign n_n5256 = ( wire19  &  n_n500  &  n_n534 ) ;
 assign n_n5253 = ( wire20  &  n_n509  &  n_n65 ) ;
 assign n_n1139 = ( n_n5255 ) | ( n_n5256 ) | ( n_n5253 ) ;
 assign n_n4408 = ( wire16  &  n_n473  &  n_n534 ) ;
 assign n_n4414 = ( wire16  &  n_n473  &  n_n528 ) ;
 assign wire215 = ( i_9_  &  n_n536  &  n_n473  &  n_n520 ) | ( (~ i_9_)  &  n_n536  &  n_n473  &  n_n520 ) ;
 assign n_n2169 = ( n_n2200 ) | ( wire16691 ) | ( wire16692 ) | ( wire16696 ) ;
 assign n_n5170 = ( wire12  &  n_n524  &  n_n482 ) ;
 assign wire168 = ( i_9_  &  n_n482  &  n_n534  &  n_n130 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n130 ) ;
 assign n_n2159 = ( n_n2169 ) | ( wire16682 ) | ( wire16683 ) | ( wire16705 ) ;
 assign n_n2214 = ( n_n5060 ) | ( n_n5055 ) | ( wire16733 ) | ( wire16734 ) ;
 assign n_n2168 = ( n_n2196 ) | ( wire16753 ) | ( wire16754 ) | ( wire16758 ) ;
 assign n_n5333 = ( wire20  &  n_n464  &  n_n65 ) ;
 assign n_n4429 = ( wire15  &  n_n536  &  n_n464 ) ;
 assign n_n4813 = ( wire15  &  n_n464  &  n_n325 ) ;
 assign n_n4815 = ( wire11  &  n_n464  &  n_n325 ) ;
 assign n_n4838 = ( wire17  &  n_n535  &  n_n520 ) ;
 assign wire85 = ( wire14  &  n_n464  &  n_n528 ) ;
 assign n_n2096 = ( n_n4815 ) | ( n_n4838 ) | ( wire16811 ) | ( wire16812 ) ;
 assign n_n4715 = ( wire24  &  n_n325  &  n_n518 ) ;
 assign n_n4714 = ( wire14  &  n_n532  &  n_n518 ) ;
 assign n_n5225 = ( wire25  &  n_n518  &  n_n65 ) ;
 assign n_n5224 = ( wire19  &  n_n534  &  n_n518 ) ;
 assign n_n1530 = ( n_n5226 ) | ( n_n5225 ) | ( n_n5224 ) ;
 assign wire437 = ( i_9_  &  n_n526  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n482  &  n_n130 ) ;
 assign n_n5279 = ( wire11  &  n_n491  &  n_n65 ) ;
 assign n_n5277 = ( wire15  &  n_n491  &  n_n65 ) ;
 assign n_n4708 = ( wire14  &  n_n522  &  n_n535 ) ;
 assign n_n4706 = ( wire14  &  n_n524  &  n_n535 ) ;
 assign wire366 = ( wire14  &  n_n532  &  n_n518 ) | ( wire14  &  n_n534  &  n_n518 ) ;
 assign n_n4427 = ( wire24  &  n_n536  &  n_n464 ) ;
 assign n_n4716 = ( wire14  &  n_n530  &  n_n518 ) ;
 assign n_n4807 = ( wire23  &  n_n473  &  n_n325 ) ;
 assign n_n1162 = ( n_n5136 ) | ( n_n5135 ) | ( n_n5134 ) ;
 assign n_n5312 = ( wire19  &  n_n473  &  n_n526 ) ;
 assign n_n5313 = ( wire22  &  n_n473  &  n_n65 ) ;
 assign n_n4596 = ( wire10  &  n_n522  &  n_n518 ) ;
 assign wire256 = ( wire10  &  n_n509  &  n_n530 ) | ( wire10  &  n_n509  &  n_n532 ) ;
 assign n_n1059 = ( n_n5128 ) | ( n_n5133 ) | ( n_n1162 ) | ( wire11912 ) ;
 assign wire28 = ( wire335 ) | ( n_n5115 ) | ( wire11914 ) ;
 assign n_n4672 = ( wire10  &  n_n473  &  n_n526 ) ;
 assign n_n4468 = ( wire13  &  n_n522  &  n_n518 ) ;
 assign n_n4418 = ( wire16  &  n_n473  &  n_n524 ) ;
 assign n_n4446 = ( wire13  &  n_n535  &  n_n528 ) ;
 assign n_n4688 = ( wire10  &  n_n464  &  n_n526 ) ;
 assign n_n4836 = ( wire17  &  n_n522  &  n_n535 ) ;
 assign n_n4871 = ( wire23  &  n_n509  &  n_n260 ) ;
 assign n_n4961 = ( wire22  &  n_n535  &  n_n195 ) ;
 assign n_n5140 = ( wire12  &  n_n522  &  n_n500 ) ;
 assign n_n5194 = ( wire12  &  n_n464  &  n_n532 ) ;
 assign n_n5259 = ( wire24  &  n_n500  &  n_n65 ) ;
 assign n_n5271 = ( wire23  &  n_n500  &  n_n65 ) ;
 assign n_n4537 = ( wire25  &  n_n473  &  n_n455 ) ;
 assign n_n4614 = ( wire10  &  n_n509  &  n_n520 ) ;
 assign n_n4058 = ( n_n4917 ) | ( n_n4914 ) | ( wire13202 ) | ( wire13203 ) ;
 assign n_n3993 = ( n_n4016 ) | ( wire13467 ) | ( wire13468 ) | ( wire13482 ) ;
 assign n_n3995 = ( n_n4021 ) | ( wire13519 ) | ( wire13520 ) | ( wire13547 ) ;
 assign wire55 = ( wire12471 ) | ( wire13  &  n_n528  &  n_n518 ) ;
 assign n_n3986 = ( n_n3993 ) | ( n_n3995 ) | ( wire13553 ) | ( wire13554 ) ;
 assign n_n4707 = ( wire21  &  n_n535  &  n_n325 ) ;
 assign n_n4701 = ( wire15  &  n_n535  &  n_n325 ) ;
 assign n_n4643 = ( wire21  &  n_n491  &  n_n390 ) ;
 assign n_n4642 = ( wire10  &  n_n524  &  n_n491 ) ;
 assign n_n3716 = ( n_n3861 ) | ( n_n4620 ) | ( n_n4625 ) | ( wire14393 ) ;
 assign n_n3650 = ( n_n3716 ) | ( wire14397 ) | ( wire14398 ) | ( wire14405 ) ;
 assign n_n4556 = ( wire13  &  n_n464  &  n_n530 ) ;
 assign n_n4550 = ( wire13  &  n_n473  &  n_n520 ) ;
 assign n_n3870 = ( wire455 ) | ( wire13  &  n_n522  &  n_n464 ) ;
 assign wire91 = ( wire13  &  n_n464  &  n_n520 ) ;
 assign wire430 = ( i_9_  &  n_n464  &  n_n455  &  n_n532 ) | ( (~ i_9_)  &  n_n464  &  n_n455  &  n_n532 ) ;
 assign n_n4609 = ( wire22  &  n_n509  &  n_n390 ) ;
 assign n_n3718 = ( n_n4597 ) | ( n_n4588 ) | ( wire14422 ) | ( wire14423 ) ;
 assign n_n3629 = ( n_n3650 ) | ( wire14419 ) | ( wire14420 ) | ( wire14436 ) ;
 assign n_n4358 = ( wire16  &  n_n509  &  n_n520 ) ;
 assign n_n4493 = ( wire15  &  n_n455  &  n_n500 ) ;
 assign n_n5148 = ( wire12  &  n_n491  &  n_n530 ) ;
 assign n_n3461 = ( n_n4831 ) | ( n_n4832 ) | ( n_n4833 ) ;
 assign n_n3329 = ( n_n4836 ) | ( n_n3461 ) | ( wire11769 ) | ( wire13808 ) ;
 assign n_n5126 = ( wire12  &  n_n509  &  n_n520 ) ;
 assign n_n3307 = ( n_n5128 ) | ( n_n5125 ) | ( wire13923 ) | ( wire13924 ) ;
 assign n_n3277 = ( wire13796 ) | ( wire13797 ) ;
 assign n_n4808 = ( wire14  &  n_n464  &  n_n534 ) ;
 assign n_n3330 = ( n_n4827 ) | ( n_n4822 ) | ( wire13803 ) | ( wire13804 ) ;
 assign n_n3275 = ( n_n3329 ) | ( wire13812 ) | ( wire13813 ) | ( wire13820 ) ;
 assign n_n2710 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) ;
 assign n_n3274 = ( n_n3326 ) | ( wire13855 ) | ( wire13856 ) | ( wire13860 ) ;
 assign wire58 = ( wire13867 ) | ( wire17  &  n_n464  &  n_n526 ) ;
 assign n_n3257 = ( n_n3274 ) | ( wire13843 ) | ( wire13844 ) | ( wire13878 ) ;
 assign wire456 = ( n_n4737 ) | ( n_n4738 ) | ( wire373 ) | ( wire12778 ) ;
 assign n_n4799 = ( wire11  &  n_n473  &  n_n325 ) ;
 assign n_n3202 = ( n_n4767 ) | ( n_n4752 ) | ( wire13746 ) | ( wire13747 ) ;
 assign n_n3204 = ( n_n4629 ) | ( n_n4583 ) | ( wire13752 ) | ( wire13753 ) ;
 assign n_n4685 = ( wire15  &  n_n464  &  n_n390 ) ;
 assign n_n4520 = ( wire13  &  n_n482  &  n_n534 ) ;
 assign n_n4884 = ( wire17  &  n_n522  &  n_n500 ) ;
 assign n_n5008 = ( wire18  &  n_n526  &  n_n500 ) ;
 assign n_n4623 = ( wire11  &  n_n500  &  n_n390 ) ;
 assign wire304 = ( wire17  &  n_n522  &  n_n535 ) | ( wire17  &  n_n524  &  n_n535 ) ;
 assign n_n2601 = ( n_n4837 ) | ( n_n4841 ) | ( n_n3461 ) | ( wire14894 ) ;
 assign n_n2602 = ( n_n4824 ) | ( n_n4823 ) | ( wire14898 ) | ( wire14899 ) ;
 assign wire433 = ( i_9_  &  n_n500  &  n_n534  &  n_n65 ) | ( (~ i_9_)  &  n_n500  &  n_n534  &  n_n65 ) ;
 assign n_n5242 = ( wire19  &  n_n509  &  n_n532 ) ;
 assign wire320 = ( wire20  &  n_n518  &  n_n65 ) | ( wire23  &  n_n518  &  n_n65 ) ;
 assign n_n5264 = ( wire19  &  n_n526  &  n_n500 ) ;
 assign n_n5270 = ( wire19  &  n_n500  &  n_n520 ) ;
 assign wire77 = ( i_9_  &  n_n522  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n522  &  n_n500  &  n_n65 ) ;
 assign wire334 = ( i_9_  &  n_n524  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n500  &  n_n65 ) ;
 assign wire149 = ( wire19  &  n_n522  &  n_n464 ) | ( wire19  &  n_n464  &  n_n520 ) ;
 assign wire267 = ( wire115 ) | ( n_n5315 ) | ( wire13557 ) ;
 assign n_n2564 = ( n_n5305 ) | ( n_n5302 ) | ( wire15194 ) | ( wire15195 ) ;
 assign n_n2566 = ( n_n5274 ) | ( n_n5271 ) | ( n_n2651 ) | ( wire15198 ) ;
 assign wire218 = ( i_9_  &  n_n524  &  n_n491  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n491  &  n_n65 ) ;
 assign wire385 = ( i_9_  &  n_n532  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n532  &  n_n518  &  n_n65 ) ;
 assign wire399 = ( i_9_  &  n_n509  &  n_n536  &  n_n528 ) | ( (~ i_9_)  &  n_n509  &  n_n536  &  n_n528 ) ;
 assign wire125 = ( wire24  &  n_n491  &  n_n130 ) | ( wire25  &  n_n491  &  n_n130 ) ;
 assign n_n2196 = ( n_n5294 ) | ( n_n5299 ) | ( wire16748 ) | ( wire16749 ) ;
 assign wire44 = ( i_9_  &  n_n520  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n520  &  n_n482  &  n_n130 ) ;
 assign wire332 = ( i_9_  &  n_n522  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n482  &  n_n130 ) ;
 assign wire90 = ( n_n5075 ) | ( n_n5078 ) | ( n_n5080 ) | ( wire209 ) ;
 assign wire144 = ( n_n5091 ) | ( n_n5090 ) | ( wire13305 ) | ( wire13306 ) ;
 assign wire239 = ( wire10  &  n_n535  &  n_n528 ) | ( wire10  &  n_n535  &  n_n530 ) ;
 assign n_n4335 = ( wire11  &  n_n536  &  n_n518 ) ;
 assign n_n4411 = ( wire24  &  n_n536  &  n_n473 ) ;
 assign n_n4279 = ( n_n4329 ) | ( n_n4328 ) | ( n_n4330 ) ;
 assign n_n5219 = ( wire21  &  n_n535  &  n_n65 ) ;
 assign n_n1456 = ( n_n4983 ) | ( n_n4984 ) | ( wire57 ) | ( wire12156 ) ;
 assign n_n1521 = ( n_n5272 ) | ( n_n5271 ) | ( n_n5270 ) ;
 assign n_n4528 = ( wire13  &  n_n526  &  n_n482 ) ;
 assign n_n4529 = ( wire22  &  n_n455  &  n_n482 ) ;
 assign n_n5319 = ( wire23  &  n_n473  &  n_n65 ) ;
 assign wire328 = ( i_9_  &  n_n536  &  n_n473  &  n_n530 ) | ( (~ i_9_)  &  n_n536  &  n_n473  &  n_n530 ) ;
 assign n_n4542 = ( wire13  &  n_n473  &  n_n528 ) ;
 assign wire201 = ( i_9_  &  n_n473  &  n_n455  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n530 ) ;
 assign n_n4543 = ( wire11  &  n_n473  &  n_n455 ) ;
 assign n_n4549 = ( wire20  &  n_n473  &  n_n455 ) ;
 assign n_n4551 = ( wire23  &  n_n473  &  n_n455 ) ;
 assign n_n4691 = ( wire21  &  n_n464  &  n_n390 ) ;
 assign n_n3849 = ( n_n4690 ) | ( n_n4689 ) | ( n_n4691 ) ;
 assign n_n4692 = ( wire10  &  n_n522  &  n_n464 ) ;
 assign n_n1093 = ( n_n4683 ) | ( n_n3849 ) | ( n_n4692 ) | ( wire11862 ) ;
 assign wire299 = ( i_9_  &  n_n500  &  n_n530  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n530  &  n_n195 ) ;
 assign n_n1050 = ( n_n5244 ) | ( n_n5249 ) | ( n_n1139 ) | ( wire11921 ) ;
 assign n_n5269 = ( wire20  &  n_n500  &  n_n65 ) ;
 assign n_n5257 = ( wire25  &  n_n500  &  n_n65 ) ;
 assign wire62 = ( i_9_  &  n_n500  &  n_n532  &  n_n65 ) | ( (~ i_9_)  &  n_n500  &  n_n532  &  n_n65 ) ;
 assign wire92 = ( wire11  &  n_n500  &  n_n65 ) ;
 assign wire409 = ( i_9_  &  n_n500  &  n_n530  &  n_n65 ) | ( (~ i_9_)  &  n_n500  &  n_n530  &  n_n65 ) ;
 assign n_n1049 = ( wire409 ) | ( wire11923 ) | ( wire11927 ) ;
 assign n_n1048 = ( n_n5273 ) | ( n_n5278 ) | ( n_n1521 ) | ( wire11933 ) ;
 assign wire63 = ( i_9_  &  n_n522  &  n_n482  &  n_n65 ) | ( (~ i_9_)  &  n_n522  &  n_n482  &  n_n65 ) ;
 assign wire200 = ( wire19  &  n_n524  &  n_n482 ) | ( wire19  &  n_n526  &  n_n482 ) ;
 assign n_n1017 = ( n_n1048 ) | ( wire11929 ) | ( wire11930 ) | ( wire11940 ) ;
 assign n_n1045 = ( n_n5303 ) | ( n_n5311 ) | ( n_n1128 ) | ( wire11944 ) ;
 assign n_n1900 = ( wire11946 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire115 = ( i_9_  &  n_n522  &  n_n473  &  n_n65 ) | ( (~ i_9_)  &  n_n522  &  n_n473  &  n_n65 ) ;
 assign wire175 = ( i_9_  &  n_n464  &  n_n530  &  n_n65 ) | ( (~ i_9_)  &  n_n464  &  n_n530  &  n_n65 ) ;
 assign n_n1007 = ( n_n1050 ) | ( n_n1049 ) | ( n_n1017 ) | ( wire11962 ) ;
 assign n_n4476 = ( wire13  &  n_n509  &  n_n530 ) ;
 assign n_n4686 = ( wire10  &  n_n464  &  n_n528 ) ;
 assign n_n4354 = ( wire16  &  n_n509  &  n_n524 ) ;
 assign n_n4889 = ( wire25  &  n_n491  &  n_n260 ) ;
 assign n_n5196 = ( wire12  &  n_n464  &  n_n530 ) ;
 assign n_n5203 = ( wire21  &  n_n464  &  n_n130 ) ;
 assign n_n5210 = ( wire19  &  n_n535  &  n_n532 ) ;
 assign n_n5217 = ( wire22  &  n_n535  &  n_n65 ) ;
 assign n_n3996 = ( wire267 ) | ( wire13566 ) | ( wire13567 ) ;
 assign n_n4929 = ( wire22  &  n_n473  &  n_n260 ) ;
 assign n_n4766 = ( wire14  &  n_n528  &  n_n491 ) ;
 assign wire447 = ( n_n4770 ) | ( n_n4771 ) | ( wire164 ) | ( wire12393 ) ;
 assign n_n1592 = ( n_n4921 ) | ( n_n4918 ) | ( n_n4919 ) ;
 assign n_n4742 = ( wire14  &  n_n509  &  n_n520 ) ;
 assign n_n4527 = ( wire11  &  n_n455  &  n_n482 ) ;
 assign n_n4713 = ( wire25  &  n_n325  &  n_n518 ) ;
 assign n_n3708 = ( n_n4715 ) | ( n_n4716 ) | ( wire14346 ) | ( wire14347 ) ;
 assign n_n3648 = ( n_n3708 ) | ( wire14350 ) | ( wire14351 ) | ( wire14357 ) ;
 assign n_n4657 = ( wire22  &  n_n390  &  n_n482 ) ;
 assign n_n3711 = ( n_n4222 ) | ( n_n3849 ) | ( wire14363 ) ;
 assign n_n3649 = ( n_n3711 ) | ( wire14361 ) | ( wire14362 ) | ( wire14371 ) ;
 assign n_n3653 = ( n_n3724 ) | ( wire14453 ) | ( wire14454 ) | ( wire14458 ) ;
 assign n_n3655 = ( n_n3729 ) | ( wire14521 ) | ( wire14522 ) | ( wire14530 ) ;
 assign n_n5090 = ( wire12  &  n_n524  &  n_n535 ) ;
 assign n_n5144 = ( wire12  &  n_n491  &  n_n534 ) ;
 assign n_n5143 = ( wire23  &  n_n500  &  n_n130 ) ;
 assign n_n2685 = ( n_n5120 ) | ( n_n5117 ) | ( n_n5119 ) ;
 assign n_n3308 = ( n_n5109 ) | ( n_n5113 ) | ( n_n2685 ) | ( wire13929 ) ;
 assign n_n5007 = ( wire11  &  n_n500  &  n_n195 ) ;
 assign wire211 = ( i_9_  &  n_n522  &  n_n500  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n500  &  n_n130 ) ;
 assign n_n3251 = ( wire14065 ) | ( wire14066 ) | ( wire14068 ) ;
 assign n_n4953 = ( wire25  &  n_n535  &  n_n195 ) ;
 assign n_n3201 = ( n_n4844 ) | ( n_n4839 ) | ( wire13772 ) | ( wire13773 ) ;
 assign n_n4334 = ( wire16  &  n_n528  &  n_n518 ) ;
 assign wire158 = ( i_9_  &  n_n473  &  n_n534  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n534  &  n_n325 ) ;
 assign wire380 = ( wire14  &  n_n473  &  n_n528 ) | ( wire14  &  n_n473  &  n_n530 ) ;
 assign n_n4874 = ( wire17  &  n_n500  &  n_n532 ) ;
 assign wire49 = ( i_9_  &  n_n491  &  n_n530  &  n_n260 ) | ( (~ i_9_)  &  n_n491  &  n_n530  &  n_n260 ) ;
 assign wire87 = ( wire11  &  n_n518  &  n_n65 ) ;
 assign wire182 = ( i_9_  &  n_n526  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n65 ) ;
 assign n_n5215 = ( wire11  &  n_n535  &  n_n65 ) ;
 assign wire220 = ( i_9_  &  n_n522  &  n_n464  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n130 ) ;
 assign wire384 = ( wire20  &  n_n535  &  n_n65 ) | ( wire23  &  n_n535  &  n_n65 ) ;
 assign wire454 = ( wire24  &  n_n535  &  n_n65 ) | ( wire15  &  n_n535  &  n_n65 ) ;
 assign n_n4534 = ( wire13  &  n_n520  &  n_n482 ) ;
 assign n_n2558 = ( n_n2630 ) | ( wire15065 ) | ( wire15066 ) | ( wire15075 ) ;
 assign n_n2626 = ( n_n4521 ) | ( n_n4511 ) | ( wire15079 ) | ( wire15080 ) ;
 assign n_n2533 = ( n_n2558 ) | ( wire15094 ) | ( wire15095 ) | ( wire15103 ) ;
 assign wire82 = ( n_n4553 ) | ( n_n4554 ) | ( n_n4552 ) ;
 assign wire224 = ( n_n4568 ) | ( wire471 ) | ( wire783 ) | ( wire11564 ) ;
 assign n_n5248 = ( wire19  &  n_n509  &  n_n526 ) ;
 assign n_n4412 = ( wire16  &  n_n473  &  n_n530 ) ;
 assign n_n2651 = ( n_n5281 ) | ( n_n5279 ) | ( n_n5280 ) ;
 assign n_n5195 = ( wire24  &  n_n464  &  n_n130 ) ;
 assign n_n5197 = ( wire15  &  n_n464  &  n_n130 ) ;
 assign n_n2291 = ( n_n5210 ) | ( n_n5209 ) | ( n_n5208 ) ;
 assign wire451 = ( wire12  &  n_n464  &  n_n530 ) | ( wire12  &  n_n464  &  n_n532 ) ;
 assign n_n4316 = ( wire16  &  n_n535  &  n_n530 ) ;
 assign n_n4313 = ( wire25  &  n_n536  &  n_n535 ) ;
 assign n_n4723 = ( wire21  &  n_n325  &  n_n518 ) ;
 assign n_n4722 = ( wire14  &  n_n524  &  n_n518 ) ;
 assign n_n4892 = ( wire17  &  n_n491  &  n_n530 ) ;
 assign n_n5213 = ( wire15  &  n_n535  &  n_n65 ) ;
 assign n_n5209 = ( wire25  &  n_n535  &  n_n65 ) ;
 assign n_n1532 = ( n_n5210 ) | ( n_n5213 ) | ( n_n5209 ) ;
 assign wire288 = ( i_9_  &  n_n500  &  n_n520  &  n_n130 ) | ( (~ i_9_)  &  n_n500  &  n_n520  &  n_n130 ) ;
 assign n_n5247 = ( wire11  &  n_n509  &  n_n65 ) ;
 assign wire446 = ( i_9_  &  n_n509  &  n_n526  &  n_n65 ) | ( (~ i_9_)  &  n_n509  &  n_n526  &  n_n65 ) ;
 assign n_n1435 = ( n_n5254 ) | ( n_n5259 ) | ( wire446 ) | ( wire12349 ) ;
 assign n_n1103 = ( n_n4555 ) | ( n_n4556 ) | ( wire82 ) | ( wire11541 ) ;
 assign wire181 = ( i_9_  &  n_n530  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n530  &  n_n518  &  n_n65 ) ;
 assign wire452 = ( wire12  &  n_n464  &  n_n528 ) | ( wire12  &  n_n464  &  n_n530 ) ;
 assign n_n5208 = ( wire19  &  n_n535  &  n_n534 ) ;
 assign n_n5211 = ( wire24  &  n_n535  &  n_n65 ) ;
 assign n_n1038 = ( n_n1111 ) | ( wire11511 ) | ( wire11512 ) | ( wire11518 ) ;
 assign wire79 = ( i_9_  &  n_n536  &  n_n473  &  n_n524 ) | ( (~ i_9_)  &  n_n536  &  n_n473  &  n_n524 ) ;
 assign n_n3875 = ( wire11543 ) | ( wire13  &  n_n520  &  n_n482 ) ;
 assign n_n1040 = ( wire11600 ) | ( wire11601 ) | ( wire11602 ) | ( wire11605 ) ;
 assign n_n4322 = ( wire16  &  n_n524  &  n_n535 ) ;
 assign n_n1041 = ( n_n1120 ) | ( n_n3176 ) | ( wire11614 ) | ( wire11618 ) ;
 assign n_n4695 = ( wire23  &  n_n464  &  n_n390 ) ;
 assign n_n4826 = ( wire17  &  n_n535  &  n_n532 ) ;
 assign n_n5151 = ( wire11  &  n_n491  &  n_n130 ) ;
 assign n_n4197 = ( n_n4811 ) | ( n_n4810 ) | ( wire773 ) ;
 assign n_n4883 = ( wire21  &  n_n500  &  n_n260 ) ;
 assign wire330 = ( i_9_  &  n_n528  &  n_n500  &  n_n260 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n260 ) ;
 assign n_n5071 = ( wire11  &  n_n464  &  n_n195 ) ;
 assign n_n1167 = ( n_n5100 ) | ( n_n5103 ) | ( n_n5102 ) ;
 assign n_n3253 = ( n_n3260 ) | ( n_n3262 ) | ( wire14211 ) ;
 assign n_n2997 = ( n_n4515 ) | ( n_n3152 ) | ( n_n4520 ) | ( wire15440 ) ;
 assign n_n5198 = ( wire12  &  n_n464  &  n_n528 ) ;
 assign n_n3037 = ( wire14615 ) | ( wire11  &  n_n535  &  n_n65 ) ;
 assign wire183 = ( wire21  &  n_n535  &  n_n65 ) | ( wire20  &  n_n535  &  n_n65 ) ;
 assign wire453 = ( wire24  &  n_n464  &  n_n130 ) | ( wire25  &  n_n464  &  n_n130 ) ;
 assign n_n5246 = ( wire19  &  n_n509  &  n_n528 ) ;
 assign n_n5176 = ( wire12  &  n_n473  &  n_n534 ) ;
 assign wire80 = ( wire21  &  n_n473  &  n_n390 ) | ( wire20  &  n_n473  &  n_n390 ) ;
 assign wire157 = ( i_9_  &  n_n473  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n530 ) ;
 assign n_n2579 = ( n_n5125 ) | ( n_n5126 ) | ( n_n2685 ) | ( wire15239 ) ;
 assign wire88 = ( wire12  &  n_n535  &  n_n520 ) ;
 assign n_n2541 = ( n_n2579 ) | ( wire15245 ) | ( wire15246 ) | ( wire15249 ) ;
 assign wire297 = ( wire25  &  n_n491  &  n_n195 ) | ( wire15  &  n_n491  &  n_n195 ) ;
 assign wire394 = ( i_9_  &  n_n526  &  n_n500  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n195 ) ;
 assign n_n2528 = ( n_n2541 ) | ( wire15234 ) | ( wire15235 ) | ( wire15264 ) ;
 assign n_n2470 = ( n_n4504 ) | ( n_n4525 ) | ( wire14838 ) | ( wire14839 ) ;
 assign n_n2467 = ( n_n4665 ) | ( n_n4708 ) | ( wire14854 ) | ( wire14855 ) ;
 assign wire361 = ( i_9_  &  n_n455  &  n_n530  &  n_n482 ) | ( (~ i_9_)  &  n_n455  &  n_n530  &  n_n482 ) ;
 assign wire378 = ( i_9_  &  n_n455  &  n_n528  &  n_n482 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n482 ) ;
 assign wire341 = ( i_9_  &  n_n534  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n534  &  n_n518  &  n_n195 ) ;
 assign wire362 = ( wire20  &  n_n535  &  n_n195 ) | ( wire23  &  n_n535  &  n_n195 ) ;
 assign wire203 = ( i_9_  &  n_n491  &  n_n534  &  n_n65 ) | ( (~ i_9_)  &  n_n491  &  n_n534  &  n_n65 ) ;
 assign wire205 = ( i_9_  &  n_n526  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n65 ) ;
 assign wire438 = ( i_9_  &  n_n491  &  n_n530  &  n_n65 ) | ( (~ i_9_)  &  n_n491  &  n_n530  &  n_n65 ) ;
 assign n_n4699 = ( wire24  &  n_n535  &  n_n325 ) ;
 assign n_n4687 = ( wire11  &  n_n464  &  n_n390 ) ;
 assign wire340 = ( wire17  &  n_n526  &  n_n482 ) | ( wire17  &  n_n528  &  n_n482 ) ;
 assign n_n5250 = ( wire19  &  n_n509  &  n_n524 ) ;
 assign n_n5205 = ( wire20  &  n_n464  &  n_n130 ) ;
 assign n_n801 = ( n_n5004 ) | ( n_n5003 ) | ( n_n5006 ) ;
 assign n_n1454 = ( n_n801 ) | ( wire12255 ) | ( wire12256 ) | ( wire12257 ) ;
 assign n_n1436 = ( n_n5243 ) | ( n_n5235 ) | ( wire12352 ) | ( wire12353 ) ;
 assign n_n5330 = ( wire19  &  n_n524  &  n_n464 ) ;
 assign n_n5331 = ( wire21  &  n_n464  &  n_n65 ) ;
 assign wire421 = ( i_9_  &  n_n455  &  n_n535  &  n_n532 ) | ( (~ i_9_)  &  n_n455  &  n_n535  &  n_n532 ) ;
 assign wire432 = ( n_n4663 ) | ( wire225 ) | ( wire11856 ) ;
 assign n_n1985 = ( n_n4885 ) | ( n_n4884 ) | ( n_n4883 ) ;
 assign n_n3815 = ( n_n4876 ) | ( n_n4875 ) | ( n_n4874 ) ;
 assign wire253 = ( i_9_  &  n_n482  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n482  &  n_n534  &  n_n195 ) ;
 assign n_n1061 = ( n_n5098 ) | ( n_n5105 ) | ( n_n1167 ) | ( wire12009 ) ;
 assign n_n1022 = ( n_n1061 ) | ( wire12014 ) | ( wire12015 ) | ( wire12020 ) ;
 assign wire104 = ( i_9_  &  n_n509  &  n_n526  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n526  &  n_n195 ) ;
 assign n_n1009 = ( n_n1022 ) | ( wire12003 ) | ( wire12004 ) | ( wire12028 ) ;
 assign n_n4323 = ( wire21  &  n_n536  &  n_n535 ) ;
 assign wire128 = ( i_9_  &  n_n455  &  n_n535  &  n_n520 ) | ( (~ i_9_)  &  n_n455  &  n_n535  &  n_n520 ) ;
 assign n_n910 = ( n_n4434 ) | ( n_n4433 ) | ( n_n4435 ) ;
 assign n_n4631 = ( wire23  &  n_n500  &  n_n390 ) ;
 assign n_n559 = ( n_n4585 ) | ( n_n4592 ) | ( wire12595 ) | ( wire12596 ) ;
 assign n_n4761 = ( wire25  &  n_n491  &  n_n325 ) ;
 assign n_n4680 = ( wire10  &  n_n464  &  n_n534 ) ;
 assign wire343 = ( wire18  &  n_n522  &  n_n500 ) | ( wire18  &  n_n524  &  n_n500 ) ;
 assign wire379 = ( wire13  &  n_n522  &  n_n482 ) | ( wire13  &  n_n524  &  n_n482 ) ;
 assign n_n2996 = ( n_n4524 ) | ( n_n4537 ) | ( wire15444 ) | ( wire15445 ) ;
 assign wire431 = ( i_9_  &  n_n528  &  n_n390  &  n_n482 ) | ( (~ i_9_)  &  n_n528  &  n_n390  &  n_n482 ) ;
 assign n_n2670 = ( n_n5200 ) | ( n_n5199 ) | ( n_n5198 ) ;
 assign n_n4402 = ( wire16  &  n_n524  &  n_n482 ) ;
 assign wire455 = ( i_9_  &  n_n524  &  n_n464  &  n_n455 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n455 ) ;
 assign wire238 = ( wire11  &  n_n535  &  n_n390 ) | ( wire15  &  n_n535  &  n_n390 ) ;
 assign wire276 = ( i_9_  &  n_n524  &  n_n535  &  n_n390 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n390 ) ;
 assign n_n4702 = ( wire14  &  n_n535  &  n_n528 ) ;
 assign n_n1455 = ( n_n4991 ) | ( n_n1576 ) | ( n_n5000 ) | ( wire12159 ) ;
 assign n_n4599 = ( wire23  &  n_n390  &  n_n518 ) ;
 assign wire364 = ( i_9_  &  n_n536  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n536  &  n_n535  &  n_n530 ) ;
 assign n_n5283 = ( wire21  &  n_n491  &  n_n65 ) ;
 assign wire333 = ( i_9_  &  n_n491  &  n_n532  &  n_n65 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n65 ) ;
 assign n_n4632 = ( wire10  &  n_n491  &  n_n534 ) ;
 assign wire139 = ( i_9_  &  n_n491  &  n_n520  &  n_n390 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n390 ) ;
 assign n_n953 = ( n_n4684 ) | ( n_n4708 ) | ( wire11646 ) | ( wire11647 ) ;
 assign wire99 = ( i_9_  &  n_n526  &  n_n535  &  n_n390 ) | ( (~ i_9_)  &  n_n526  &  n_n535  &  n_n390 ) ;
 assign n_n942 = ( n_n953 ) | ( wire11641 ) | ( wire11642 ) | ( wire11655 ) ;
 assign n_n725 = ( wire184 ) | ( n_n901 ) | ( wire787 ) | ( wire13020 ) ;
 assign wire52 = ( i_9_  &  n_n528  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n528  &  n_n518  &  n_n260 ) ;
 assign wire150 = ( wire22  &  n_n464  &  n_n325 ) | ( wire23  &  n_n464  &  n_n325 ) ;
 assign n_n4645 = ( wire20  &  n_n491  &  n_n390 ) ;
 assign wire310 = ( wire21  &  n_n491  &  n_n390 ) | ( wire22  &  n_n491  &  n_n390 ) ;
 assign n_n4696 = ( wire14  &  n_n535  &  n_n534 ) ;
 assign n_n4762 = ( wire14  &  n_n491  &  n_n532 ) ;
 assign n_n5315 = ( wire21  &  n_n473  &  n_n65 ) ;
 assign n_n1952 = ( n_n5069 ) | ( n_n5070 ) | ( n_n5071 ) ;
 assign wire363 = ( n_n4318 ) | ( n_n4321 ) | ( wire13512 ) ;
 assign wire407 = ( i_9_  &  n_n491  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n130 ) ;
 assign n_n4056 = ( wire13208 ) | ( wire13209 ) ;
 assign wire42 = ( i_9_  &  n_n473  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n260 ) ;
 assign n_n814 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4947 ) ;
 assign wire141 = ( wire18  &  n_n535  &  n_n532 ) | ( wire18  &  n_n535  &  n_n534 ) ;
 assign wire317 = ( wire20  &  n_n464  &  n_n260 ) | ( wire23  &  n_n464  &  n_n260 ) ;
 assign n_n5192 = ( wire12  &  n_n464  &  n_n534 ) ;
 assign wire106 = ( wire20  &  n_n536  &  n_n535 ) | ( wire23  &  n_n536  &  n_n535 ) ;
 assign wire375 = ( i_9_  &  n_n524  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n260 ) ;
 assign n_n4558 = ( wire13  &  n_n464  &  n_n528 ) ;
 assign wire417 = ( i_9_  &  n_n473  &  n_n520  &  n_n390 ) | ( (~ i_9_)  &  n_n473  &  n_n520  &  n_n390 ) ;
 assign wire27 = ( wire12449 ) | ( wire15  &  n_n536  &  n_n491 ) ;
 assign n_n1472 = ( n_n4783 ) | ( n_n4778 ) | ( wire12207 ) | ( wire12208 ) ;
 assign n_n763 = ( n_n5218 ) | ( n_n5217 ) | ( n_n5215 ) ;
 assign wire286 = ( wire21  &  n_n509  &  n_n130 ) | ( wire20  &  n_n509  &  n_n130 ) ;
 assign n_n667 = ( n_n5244 ) | ( n_n5243 ) | ( wire12871 ) | ( wire12872 ) ;
 assign n_n761 = ( wire12874 ) | ( wire19  &  n_n534  &  n_n518 ) ;
 assign n_n635 = ( n_n667 ) | ( wire12876 ) | ( wire12877 ) | ( wire12881 ) ;
 assign n_n777 = ( wire12884 ) | ( wire12  &  n_n522  &  n_n500 ) ;
 assign n_n3772 = ( n_n5130 ) | ( n_n5131 ) | ( n_n5132 ) ;
 assign n_n637 = ( n_n777 ) | ( n_n3772 ) | ( wire12894 ) | ( wire12898 ) ;
 assign n_n4552 = ( wire13  &  n_n464  &  n_n534 ) ;
 assign n_n4559 = ( wire11  &  n_n464  &  n_n455 ) ;
 assign n_n5227 = ( wire24  &  n_n518  &  n_n65 ) ;
 assign n_n5304 = ( wire19  &  n_n473  &  n_n534 ) ;
 assign n_n4694 = ( wire10  &  n_n464  &  n_n520 ) ;
 assign n_n4700 = ( wire14  &  n_n535  &  n_n530 ) ;
 assign n_n4219 = ( n_n4704 ) | ( n_n4703 ) | ( n_n4702 ) ;
 assign wire221 = ( i_9_  &  n_n535  &  n_n532  &  n_n325 ) | ( (~ i_9_)  &  n_n535  &  n_n532  &  n_n325 ) ;
 assign n_n4075 = ( n_n4694 ) | ( n_n4700 ) | ( n_n4219 ) | ( wire13244 ) ;
 assign wire30 = ( n_n4709 ) | ( wire14  &  n_n535  &  n_n520 ) ;
 assign wire173 = ( i_9_  &  n_n532  &  n_n325  &  n_n518 ) | ( (~ i_9_)  &  n_n532  &  n_n325  &  n_n518 ) ;
 assign wire243 = ( wire13246 ) | ( wire14  &  n_n509  &  n_n534 ) ;
 assign n_n4065 = ( n_n4827 ) | ( n_n4824 ) | ( wire388 ) | ( wire13156 ) ;
 assign wire390 = ( n_n4820 ) | ( n_n4819 ) | ( wire85 ) | ( wire12225 ) ;
 assign n_n3926 = ( n_n5112 ) | ( n_n5123 ) | ( wire13576 ) | ( wire13580 ) ;
 assign n_n3924 = ( n_n5219 ) | ( n_n5250 ) | ( wire13585 ) | ( wire13586 ) ;
 assign n_n3923 = ( n_n5333 ) | ( n_n5312 ) | ( wire13591 ) | ( wire13592 ) ;
 assign n_n3928 = ( n_n4994 ) | ( n_n5009 ) | ( wire13598 ) | ( wire13599 ) ;
 assign n_n3124 = ( wire13897 ) | ( wire21  &  n_n535  &  n_n325 ) ;
 assign n_n2378 = ( n_n4704 ) | ( n_n4703 ) | ( n_n4705 ) ;
 assign n_n4693 = ( wire20  &  n_n464  &  n_n390 ) ;
 assign n_n3051 = ( n_n5129 ) | ( n_n5127 ) | ( n_n5126 ) ;
 assign n_n3007 = ( n_n4388 ) | ( n_n4392 ) | ( wire15506 ) | ( wire15507 ) ;
 assign n_n3003 = ( n_n4440 ) | ( wire470 ) | ( n_n4449 ) | ( wire15426 ) ;
 assign n_n2604 = ( n_n4797 ) | ( n_n4802 ) | ( wire14917 ) | ( wire14918 ) ;
 assign n_n4910 = ( wire17  &  n_n528  &  n_n482 ) ;
 assign wire190 = ( wire21  &  n_n500  &  n_n390 ) | ( wire22  &  n_n500  &  n_n390 ) ;
 assign n_n1501 = ( n_n4403 ) | ( n_n4415 ) | ( wire12458 ) | ( wire12459 ) ;
 assign n_n1426 = ( n_n1501 ) | ( wire12464 ) | ( wire12465 ) | ( wire12469 ) ;
 assign n_n1409 = ( n_n1450 ) | ( wire12315 ) | ( wire12316 ) | ( wire12324 ) ;
 assign n_n1448 = ( n_n5078 ) | ( n_n5083 ) | ( wire12332 ) | ( wire12333 ) ;
 assign n_n1408 = ( n_n1448 ) | ( wire12327 ) | ( wire12328 ) | ( wire12340 ) ;
 assign wire347 = ( wire11  &  n_n455  &  n_n500 ) | ( wire15  &  n_n455  &  n_n500 ) ;
 assign n_n5280 = ( wire19  &  n_n526  &  n_n491 ) ;
 assign n_n5080 = ( wire12  &  n_n535  &  n_n534 ) ;
 assign n_n680 = ( n_n5061 ) | ( n_n5058 ) | ( n_n789 ) | ( wire12902 ) ;
 assign wire209 = ( i_9_  &  n_n522  &  n_n464  &  n_n195 ) | ( (~ i_9_)  &  n_n522  &  n_n464  &  n_n195 ) ;
 assign n_n639 = ( n_n680 ) | ( wire12907 ) | ( wire12908 ) | ( wire12915 ) ;
 assign n_n625 = ( n_n639 ) | ( wire12929 ) | ( wire12930 ) | ( wire12947 ) ;
 assign n_n4721 = ( wire22  &  n_n325  &  n_n518 ) ;
 assign n_n4548 = ( wire13  &  n_n522  &  n_n473 ) ;
 assign n_n4099 = ( n_n4389 ) | ( n_n4384 ) | ( wire13531 ) | ( wire13532 ) ;
 assign n_n4021 = ( n_n4099 ) | ( wire13528 ) | ( wire13529 ) | ( wire13539 ) ;
 assign n_n789 = ( n_n5064 ) | ( n_n5063 ) | ( n_n5065 ) ;
 assign wire445 = ( wire21  &  n_n464  &  n_n390 ) | ( wire20  &  n_n464  &  n_n390 ) ;
 assign wire422 = ( wire21  &  n_n500  &  n_n130 ) | ( wire22  &  n_n500  &  n_n130 ) ;
 assign wire442 = ( i_9_  &  n_n535  &  n_n530  &  n_n325 ) | ( (~ i_9_)  &  n_n535  &  n_n530  &  n_n325 ) ;
 assign wire386 = ( i_9_  &  n_n522  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n522  &  n_n518  &  n_n65 ) ;
 assign n_n3879 = ( n_n4518 ) | ( n_n4520 ) | ( wire789 ) ;
 assign n_n2058 = ( n_n4459 ) | ( n_n4456 ) | ( n_n4457 ) ;
 assign wire324 = ( i_9_  &  n_n500  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n500  &  n_n534  &  n_n260 ) ;
 assign wire305 = ( i_9_  &  n_n530  &  n_n482  &  n_n260 ) | ( (~ i_9_)  &  n_n530  &  n_n482  &  n_n260 ) ;
 assign wire291 = ( wire24  &  n_n455  &  n_n518 ) | ( wire15  &  n_n455  &  n_n518 ) ;
 assign n_n1111 = ( n_n4460 ) | ( n_n4457 ) | ( wire11507 ) | ( wire11508 ) ;
 assign n_n554 = ( n_n4870 ) | ( n_n4819 ) | ( wire12682 ) | ( wire12683 ) ;
 assign wire279 = ( i_9_  &  n_n534  &  n_n518  &  n_n130 ) | ( (~ i_9_)  &  n_n534  &  n_n518  &  n_n130 ) ;
 assign n_n4016 = ( n_n4083 ) | ( wire13445 ) | ( wire13446 ) | ( wire13452 ) ;
 assign wire401 = ( i_9_  &  n_n528  &  n_n500  &  n_n390 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n390 ) ;
 assign n_n3560 = ( n_n4708 ) | ( n_n4695 ) | ( wire14316 ) | ( wire14317 ) ;
 assign wire434 = ( wire21  &  n_n509  &  n_n65 ) | ( wire20  &  n_n509  &  n_n65 ) ;
 assign n_n3009 = ( n_n4365 ) | ( n_n4356 ) | ( wire15511 ) | ( wire15512 ) ;
 assign n_n4330 = ( wire16  &  n_n532  &  n_n518 ) ;
 assign n_n3889 = ( wire11520 ) | ( wire13  &  n_n535  &  n_n520 ) ;
 assign n_n2238 = ( n_n4724 ) | ( n_n4727 ) | ( wire16388 ) | ( wire16389 ) ;
 assign n_n4872 = ( wire17  &  n_n500  &  n_n534 ) ;
 assign n_n1677 = ( n_n4487 ) | ( n_n4488 ) | ( n_n4486 ) ;
 assign n_n1496 = ( n_n4471 ) | ( n_n4472 ) | ( wire12492 ) | ( wire12493 ) ;
 assign n_n1467 = ( n_n4848 ) | ( n_n4839 ) | ( wire12234 ) | ( wire12235 ) ;
 assign n_n1415 = ( n_n1467 ) | ( wire12230 ) | ( wire12231 ) | ( wire12240 ) ;
 assign n_n1091 = ( n_n4710 ) | ( n_n4719 ) | ( wire11866 ) | ( wire11867 ) ;
 assign n_n4030 = ( n_n5252 ) | ( n_n5261 ) | ( wire13337 ) | ( wire13338 ) ;
 assign wire124 = ( i_9_  &  n_n522  &  n_n536  &  n_n518 ) | ( (~ i_9_)  &  n_n522  &  n_n536  &  n_n518 ) ;
 assign n_n1402 = ( wire12363 ) | ( wire12364 ) | ( wire12368 ) | ( wire12369 ) ;
 assign wire204 = ( n_n5276 ) | ( n_n5277 ) | ( wire12371 ) | ( wire12372 ) ;
 assign n_n956 = ( n_n4479 ) | ( n_n4468 ) | ( wire11666 ) | ( wire11667 ) ;
 assign n_n941 = ( n_n951 ) | ( wire11675 ) | ( wire11676 ) | ( wire11690 ) ;
 assign n_n937 = ( n_n948 ) | ( n_n949 ) | ( wire11734 ) | ( wire11735 ) ;
 assign n_n4031 = ( n_n5239 ) | ( n_n5245 ) | ( wire13341 ) | ( wire13342 ) ;
 assign wire600 = ( (~ i_9_)  &  (~ i_7_)  &  i_8_  &  (~ i_6_) ) | ( (~ i_9_)  &  i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n1418 = ( n_n1478 ) | ( n_n1476 ) | ( wire12416 ) ;
 assign n_n5289 = ( wire25  &  n_n482  &  n_n65 ) ;
 assign wire255 = ( i_9_  &  n_n522  &  n_n390  &  n_n518 ) | ( (~ i_9_)  &  n_n522  &  n_n390  &  n_n518 ) ;
 assign n_n1712 = ( n_n1727 ) | ( wire15829 ) | ( wire15830 ) | ( wire15838 ) ;
 assign n_n1730 = ( n_n4394 ) | ( n_n4376 ) | ( wire15908 ) | ( wire15909 ) ;
 assign n_n1729 = ( n_n4451 ) | ( n_n4458 ) | ( wire15914 ) | ( wire15915 ) ;
 assign n_n1711 = ( n_n1725 ) | ( n_n1724 ) | ( wire15930 ) | ( wire15931 ) ;
 assign n_n5282 = ( wire19  &  n_n524  &  n_n491 ) ;
 assign wire225 = ( i_9_  &  n_n473  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n534 ) ;
 assign n_n5298 = ( wire19  &  n_n524  &  n_n482 ) ;
 assign n_n3931 = ( n_n4701 ) | ( n_n4692 ) | ( wire13629 ) | ( wire13630 ) ;
 assign n_n3929 = ( n_n4901 ) | ( n_n4904 ) | ( wire13635 ) | ( wire13636 ) ;
 assign wire261 = ( i_9_  &  n_n491  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n491  &  n_n534  &  n_n260 ) ;
 assign n_n3694 = ( n_n4885 ) | ( n_n4890 ) | ( n_n3810 ) | ( wire14733 ) ;
 assign n_n2761 = ( n_n4648 ) | ( n_n4647 ) | ( n_n4645 ) ;
 assign n_n2982 = ( wire457 ) | ( n_n4716 ) | ( n_n4713 ) | ( wire15750 ) ;
 assign wire466 = ( n_n5155 ) | ( wire195 ) | ( n_n5160 ) | ( wire287 ) ;
 assign n_n2953 = ( n_n5091 ) | ( n_n5100 ) | ( wire15605 ) | ( wire15606 ) ;
 assign n_n2955 = ( n_n5072 ) | ( n_n5061 ) | ( wire15609 ) | ( wire15610 ) ;
 assign n_n2915 = ( n_n2953 ) | ( n_n2955 ) | ( wire15616 ) | ( wire15617 ) ;
 assign wire265 = ( i_9_  &  n_n526  &  n_n491  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n195 ) ;
 assign n_n2902 = ( n_n2915 ) | ( wire15633 ) | ( wire15634 ) | ( wire15642 ) ;
 assign n_n2839 = ( n_n4778 ) | ( n_n4745 ) | ( wire15405 ) | ( wire15406 ) ;
 assign n_n2630 = ( n_n3162 ) | ( n_n4465 ) | ( n_n4462 ) | ( wire15069 ) ;
 assign n_n1840 = ( n_n5082 ) | ( n_n5079 ) | ( n_n1952 ) | ( wire15945 ) ;
 assign n_n1801 = ( n_n1840 ) | ( wire15950 ) | ( wire15951 ) | ( wire15957 ) ;
 assign n_n1837 = ( n_n5115 ) | ( n_n5128 ) | ( wire15961 ) | ( wire15962 ) ;
 assign n_n1800 = ( n_n1837 ) | ( wire15967 ) | ( wire15968 ) | ( wire15973 ) ;
 assign n_n1842 = ( n_n5045 ) | ( n_n5053 ) | ( wire15977 ) | ( wire15978 ) ;
 assign n_n1725 = ( n_n4678 ) | ( n_n1764 ) | ( n_n4687 ) | ( wire15920 ) ;
 assign n_n707 = ( n_n4708 ) | ( n_n4707 ) | ( wire12783 ) | ( wire12784 ) ;
 assign n_n691 = ( n_n4921 ) | ( wire249 ) | ( n_n4932 ) | ( wire12718 ) ;
 assign n_n632 = ( wire12966 ) | ( wire12967 ) ;
 assign n_n646 = ( n_n700 ) | ( wire12762 ) | ( wire12763 ) | ( wire12767 ) ;
 assign n_n627 = ( n_n646 ) | ( wire12752 ) | ( wire12753 ) | ( wire12775 ) ;
 assign n_n856 = ( n_n4734 ) | ( n_n4729 ) | ( wire683 ) ;
 assign n_n648 = ( n_n707 ) | ( wire12790 ) | ( wire12791 ) | ( wire12796 ) ;
 assign n_n628 = ( n_n648 ) | ( wire12813 ) | ( wire12814 ) | ( wire12827 ) ;
 assign n_n621 = ( n_n627 ) | ( n_n628 ) | ( wire12865 ) | ( wire12866 ) ;
 assign n_n1760 = ( n_n4738 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign n_n2841 = ( n_n4691 ) | ( n_n4686 ) | ( wire15333 ) | ( wire15334 ) ;
 assign wire53 = ( i_9_  &  n_n536  &  n_n524  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n524  &  n_n518 ) ;
 assign n_n1852 = ( wire249 ) | ( n_n4932 ) | ( wire42 ) | ( wire16159 ) ;
 assign n_n1805 = ( n_n1852 ) | ( wire16164 ) | ( wire16165 ) | ( wire16168 ) ;
 assign n_n1789 = ( n_n1805 ) | ( wire16157 ) | ( wire16158 ) | ( wire16180 ) ;
 assign wire444 = ( wire10  &  n_n524  &  n_n464 ) | ( wire10  &  n_n464  &  n_n526 ) ;
 assign n_n1724 = ( n_n4725 ) | ( n_n4700 ) | ( n_n1760 ) | ( wire15924 ) ;
 assign n_n1478 = ( n_n4701 ) | ( n_n4702 ) | ( wire12403 ) | ( wire12404 ) ;
 assign n_n662 = ( n_n5302 ) | ( n_n5306 ) | ( wire12969 ) | ( wire12970 ) ;
 assign n_n661 = ( wire269 ) | ( wire12971 ) | ( wire12975 ) ;
 assign n_n620 = ( n_n635 ) | ( n_n637 ) | ( n_n625 ) | ( wire13001 ) ;
 assign n_n3736 = ( n_n4366 ) | ( n_n4375 ) | ( wire14470 ) | ( wire14471 ) ;
 assign n_n2837 = ( wire15348 ) | ( wire15349 ) ;
 assign n_n2611 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4219 ) | ( wire15008 ) ;
 assign n_n1894 = ( n_n4365 ) | ( wire13055 ) | ( wire13056 ) | ( wire16089 ) ;
 assign n_n1862 = ( n_n4802 ) | ( n_n4805 ) | ( wire16188 ) | ( wire16189 ) ;
 assign n_n1808 = ( n_n1862 ) | ( wire16193 ) | ( wire16194 ) | ( wire16198 ) ;
 assign n_n1856 = ( n_n4876 ) | ( wire461 ) | ( n_n4875 ) | ( wire16217 ) ;
 assign n_n1790 = ( n_n1808 ) | ( wire16213 ) | ( wire16214 ) | ( wire16224 ) ;
 assign n_n1727 = ( n_n4572 ) | ( n_n4518 ) | ( wire15822 ) | ( wire15823 ) ;
 assign n_n1722 = ( n_n4801 ) | ( n_n4820 ) | ( wire15851 ) | ( wire15852 ) ;
 assign n_n1721 = ( n_n4915 ) | ( n_n4961 ) | ( wire15858 ) | ( wire15859 ) ;
 assign n_n722 = ( n_n4247 ) | ( n_n4508 ) | ( wire13028 ) | ( wire13029 ) ;
 assign n_n653 = ( n_n722 ) | ( wire13034 ) | ( wire13035 ) | ( wire13039 ) ;
 assign n_n630 = ( n_n653 ) | ( wire13016 ) | ( wire13017 ) | ( wire13046 ) ;
 assign n_n3664 = ( n_n5278 ) | ( n_n5275 ) | ( wire14544 ) | ( wire14545 ) ;
 assign n_n3012 = ( n_n4317 ) | ( n_n4326 ) | ( wire363 ) | ( wire15521 ) ;
 assign n_n2934 = ( n_n3012 ) | ( wire15517 ) | ( wire15518 ) | ( wire15527 ) ;
 assign n_n2985 = ( n_n4674 ) | ( n_n4681 ) | ( wire15769 ) | ( wire15770 ) ;
 assign n_n2925 = ( n_n2985 ) | ( wire15774 ) | ( wire15775 ) | ( wire15778 ) ;
 assign n_n2824 = ( n_n2832 ) | ( n_n2834 ) | ( wire15367 ) | ( wire15368 ) ;
 assign n_n2835 = ( n_n4986 ) | ( n_n4980 ) | ( wire15389 ) | ( wire15390 ) ;
 assign n_n1892 = ( n_n4391 ) | ( n_n4396 ) | ( wire16098 ) | ( wire16099 ) ;
 assign n_n1818 = ( n_n1892 ) | ( wire16094 ) | ( wire16095 ) | ( wire16105 ) ;
 assign n_n1865 = ( n_n4764 ) | ( n_n4763 ) | ( wire16232 ) | ( wire16233 ) ;
 assign n_n1476 = ( n_n4730 ) | ( n_n4722 ) | ( wire12408 ) | ( wire12409 ) ;
 assign n_n732 = ( n_n4393 ) | ( n_n4386 ) | ( wire13073 ) | ( wire13074 ) ;
 assign n_n656 = ( n_n732 ) | ( wire13069 ) | ( wire13070 ) | ( wire13080 ) ;
 assign n_n631 = ( n_n656 ) | ( wire13065 ) | ( wire13066 ) | ( wire13088 ) ;
 assign n_n651 = ( n_n715 ) | ( wire13106 ) | ( wire13107 ) | ( wire13111 ) ;
 assign n_n629 = ( n_n651 ) | ( wire13123 ) | ( wire13124 ) | ( wire13133 ) ;
 assign n_n3561 = ( n_n4660 ) | ( n_n4665 ) | ( wire14322 ) | ( wire14323 ) ;
 assign n_n2939 = ( n_n5281 ) | ( n_n5272 ) | ( wire15653 ) | ( wire15654 ) ;
 assign n_n2832 = ( n_n5140 ) | ( n_n5144 ) | ( wire15354 ) | ( wire15355 ) ;
 assign n_n2834 = ( n_n5033 ) | ( n_n4989 ) | ( wire15360 ) | ( wire15361 ) ;
 assign n_n1032 = ( n_n1093 ) | ( n_n1091 ) | ( wire11873 ) | ( wire11874 ) ;
 assign n_n948 = ( n_n5075 ) | ( n_n5063 ) | ( wire11718 ) | ( wire11719 ) ;
 assign n_n700 = ( n_n4808 ) | ( n_n4799 ) | ( wire12756 ) | ( wire12757 ) ;
 assign n_n3689 = ( n_n3803 ) | ( n_n4953 ) | ( wire14752 ) | ( wire14754 ) ;
 assign n_n3724 = ( n_n4524 ) | ( n_n4517 ) | ( n_n3879 ) | ( wire14448 ) ;
 assign n_n949 = ( n_n5044 ) | ( n_n5011 ) | ( wire11725 ) | ( wire11726 ) ;
 assign n_n715 = ( n_n4603 ) | ( n_n4591 ) | ( wire13100 ) | ( wire13101 ) ;
 assign n_n3670 = ( n_n5199 ) | ( n_n5194 ) | ( wire14618 ) | ( wire14619 ) ;
 assign n_n2937 = ( n_n5303 ) | ( n_n3019 ) | ( n_n5313 ) | ( wire15663 ) ;
 assign n_n2929 = ( n_n2997 ) | ( n_n2996 ) | ( wire15451 ) | ( wire15452 ) ;
 assign n_n1718 = ( n_n5078 ) | ( n_n5108 ) | ( wire15870 ) | ( wire15871 ) ;
 assign n_n1717 = ( n_n5131 ) | ( n_n5127 ) | ( wire15875 ) | ( wire15879 ) ;
 assign n_n951 = ( n_n4832 ) | ( n_n4850 ) | ( wire11680 ) | ( wire11681 ) ;
 assign n_n1824 = ( n_n5296 ) | ( n_n5299 ) | ( wire16299 ) | ( wire16300 ) ;
 assign n_n1826 = ( wire334 ) | ( wire203 ) | ( wire16305 ) ;
 assign n_n1885 = ( wire65 ) | ( wire347 ) | ( wire15995 ) ;
 assign n_n1886 = ( n_n4254 ) | ( n_n4484 ) | ( wire14438 ) | ( wire15996 ) ;
 assign n_n1879 = ( n_n4574 ) | ( n_n4573 ) | ( wire16034 ) | ( wire16035 ) ;
 assign n_n1813 = ( n_n1877 ) | ( wire16040 ) | ( wire16041 ) | ( wire16048 ) ;
 assign n_n1812 = ( n_n1872 ) | ( wire16059 ) | ( wire16060 ) | ( wire16065 ) ;
 assign n_n1012 = ( n_n1032 ) | ( wire11851 ) | ( wire11852 ) | ( wire11884 ) ;
 assign n_n3729 = ( n_n4454 ) | ( wire11520 ) | ( wire14517 ) | ( wire14518 ) ;
 assign n_n3699 = ( n_n4832 ) | ( n_n3820 ) | ( n_n4837 ) | ( wire14697 ) ;
 assign n_n3701 = ( n_n4810 ) | ( n_n4813 ) | ( wire14701 ) | ( wire14702 ) ;
 assign n_n3645 = ( n_n3699 ) | ( n_n3701 ) | ( wire14708 ) | ( wire14709 ) ;
 assign n_n1872 = ( n_n4674 ) | ( n_n4661 ) | ( wire16052 ) | ( wire16053 ) ;
 assign n_n1828 = ( n_n5234 ) | ( n_n5242 ) | ( wire16266 ) | ( wire16267 ) ;
 assign n_n1797 = ( n_n1828 ) | ( wire16272 ) | ( wire16273 ) | ( wire16280 ) ;
 assign n_n3646 = ( n_n4204 ) | ( wire447 ) | ( wire14717 ) | ( wire14723 ) ;
 assign n_n3635 = ( n_n3670 ) | ( wire14624 ) | ( wire14625 ) | ( wire14629 ) ;
 assign n_n3641 = ( n_n3689 ) | ( wire14760 ) | ( wire14761 ) | ( wire14764 ) ;
 assign n_n2905 = ( n_n2925 ) | ( wire15766 ) | ( wire15767 ) | ( wire15786 ) ;
 assign wire266 = ( wire23  &  n_n464  &  n_n455 ) ;
 assign wire606 = ( wire13  &  n_n522  &  n_n491 ) ;
 assign wire617 = ( wire20  &  n_n509  &  n_n455 ) ;
 assign wire636 = ( wire12  &  n_n524  &  n_n464 ) ;
 assign wire656 = ( wire20  &  n_n482  &  n_n65 ) ;
 assign wire664 = ( wire23  &  n_n455  &  n_n491 ) ;
 assign wire669 = ( wire18  &  n_n473  &  n_n520 ) ;
 assign wire671 = ( wire13  &  n_n522  &  n_n464 ) ;
 assign wire675 = ( wire16  &  n_n509  &  n_n532 ) ;
 assign wire677 = ( wire15  &  n_n536  &  n_n518 ) ;
 assign wire679 = ( wire20  &  n_n500  &  n_n130 ) ;
 assign wire683 = ( wire24  &  n_n509  &  n_n325 ) ;
 assign wire686 = ( wire25  &  n_n464  &  n_n325 ) ;
 assign wire693 = ( wire15  &  n_n535  &  n_n260 ) ;
 assign wire695 = ( wire18  &  n_n491  &  n_n520 ) ;
 assign wire706 = ( wire18  &  n_n532  &  n_n518 ) ;
 assign wire724 = ( wire13  &  n_n524  &  n_n482 ) ;
 assign wire732 = ( wire12  &  n_n473  &  n_n530 ) ;
 assign wire735 = ( wire15  &  n_n535  &  n_n260 ) ;
 assign wire743 = ( wire20  &  n_n509  &  n_n195 ) ;
 assign wire745 = ( wire10  &  n_n491  &  n_n530 ) ;
 assign wire755 = ( wire18  &  n_n473  &  n_n520 ) ;
 assign wire761 = ( wire12  &  n_n524  &  n_n464 ) ;
 assign wire765 = ( wire12  &  n_n473  &  n_n530 ) ;
 assign wire767 = ( wire24  &  n_n509  &  n_n325 ) ;
 assign wire771 = ( wire25  &  n_n518  &  n_n195 ) ;
 assign wire772 = ( wire18  &  n_n532  &  n_n518 ) ;
 assign wire773 = ( wire25  &  n_n464  &  n_n325 ) ;
 assign wire775 = ( wire15  &  n_n390  &  n_n482 ) ;
 assign wire783 = ( wire23  &  n_n464  &  n_n455 ) ;
 assign wire787 = ( wire22  &  n_n509  &  n_n455 ) ;
 assign wire789 = ( wire23  &  n_n455  &  n_n491 ) ;
 assign wire791 = ( wire13  &  n_n522  &  n_n491 ) ;
 assign wire11482 = ( n_n4432 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire11483 = ( n_n4440 ) | ( n_n4434 ) | ( wire236 ) | ( n_n4438 ) ;
 assign wire11488 = ( wire13  &  n_n524  &  n_n491 ) | ( wire13  &  n_n491  &  n_n532 ) ;
 assign wire11489 = ( wire24  &  n_n455  &  n_n491 ) | ( wire15  &  n_n455  &  n_n491 ) ;
 assign wire11491 = ( wire11488 ) | ( wire308 ) ;
 assign wire11492 = ( n_n4508 ) | ( wire129 ) | ( wire11489 ) ;
 assign wire11495 = ( n_n4515 ) | ( n_n4492 ) | ( wire791 ) ;
 assign wire11496 = ( wire65 ) | ( n_n4520 ) | ( wire789 ) ;
 assign wire11497 = ( n_n4502 ) | ( n_n4501 ) | ( wire347 ) ;
 assign wire11498 = ( n_n4521 ) | ( n_n4504 ) | ( n_n4517 ) | ( n_n4497 ) ;
 assign wire11501 = ( n_n4524 ) | ( wire170 ) | ( wire11495 ) | ( wire11498 ) ;
 assign wire11502 = ( wire11491 ) | ( wire11492 ) | ( wire11496 ) | ( wire11497 ) ;
 assign wire11505 = ( i_9_  &  n_n524  &  n_n455  &  n_n518 ) | ( (~ i_9_)  &  n_n524  &  n_n455  &  n_n518 ) ;
 assign wire11507 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4462 ) ;
 assign wire11508 = ( wire291 ) | ( wire403 ) ;
 assign wire11511 = ( wire70 ) | ( wire13  &  n_n509  &  n_n522 ) ;
 assign wire11512 = ( n_n4489 ) | ( wire184 ) | ( n_n4486 ) | ( wire787 ) ;
 assign wire11513 = ( wire25  &  n_n509  &  n_n455 ) | ( wire23  &  n_n509  &  n_n455 ) ;
 assign wire11515 = ( n_n4470 ) | ( n_n4469 ) | ( n_n4475 ) ;
 assign wire11516 = ( n_n4471 ) | ( n_n4472 ) | ( wire11513 ) ;
 assign wire11518 = ( n_n4465 ) | ( wire11505 ) | ( wire11515 ) | ( wire11516 ) ;
 assign wire11520 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign wire11521 = ( wire13  &  n_n524  &  n_n535 ) | ( wire13  &  n_n526  &  n_n535 ) ;
 assign wire11522 = ( n_n4445 ) | ( wire368 ) | ( n_n4446 ) ;
 assign wire11523 = ( n_n4454 ) | ( wire11520 ) | ( wire11521 ) ;
 assign wire11524 = ( wire20  &  n_n536  &  n_n473 ) | ( wire23  &  n_n536  &  n_n473 ) ;
 assign wire11527 = ( wire37 ) | ( n_n4428 ) | ( wire11524 ) ;
 assign wire11529 = ( wire11482 ) | ( wire11483 ) | ( wire11522 ) | ( wire11523 ) ;
 assign wire11530 = ( wire84 ) | ( wire79 ) | ( wire11527 ) | ( wire11529 ) ;
 assign wire11532 = ( i_9_  &  n_n473  &  n_n455  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n532 ) ;
 assign wire11534 = ( wire22  &  n_n473  &  n_n455 ) | ( wire11  &  n_n473  &  n_n455 ) ;
 assign wire11535 = ( wire20  &  n_n473  &  n_n455 ) | ( wire23  &  n_n473  &  n_n455 ) ;
 assign wire11536 = ( n_n4547 ) | ( n_n4544 ) | ( wire11534 ) ;
 assign wire11537 = ( n_n4542 ) | ( wire201 ) | ( wire11535 ) ;
 assign wire11539 = ( wire22  &  n_n464  &  n_n455 ) | ( wire15  &  n_n464  &  n_n455 ) ;
 assign wire11541 = ( wire11539 ) | ( wire213 ) ;
 assign wire11543 = ( wire20  &  n_n455  &  n_n482 ) | ( wire23  &  n_n455  &  n_n482 ) ;
 assign wire11547 = ( i_9_  &  n_n500  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n500  &  n_n390  &  n_n532 ) ;
 assign wire11548 = ( n_n4617 ) | ( n_n4613 ) | ( n_n4612 ) | ( n_n4611 ) ;
 assign wire11549 = ( n_n4616 ) | ( wire465 ) | ( wire11547 ) ;
 assign wire11553 = ( n_n4634 ) | ( n_n4639 ) | ( n_n4642 ) | ( n_n4631 ) ;
 assign wire11554 = ( n_n4629 ) | ( n_n4630 ) | ( wire190 ) ;
 assign wire11555 = ( n_n4637 ) | ( n_n4648 ) | ( n_n4628 ) | ( n_n4635 ) ;
 assign wire11558 = ( wire309 ) | ( n_n3861 ) | ( n_n4626 ) | ( wire11555 ) ;
 assign wire11559 = ( wire11548 ) | ( wire11549 ) | ( wire11553 ) | ( wire11554 ) ;
 assign wire11560 = ( wire10  &  n_n509  &  n_n524 ) | ( wire10  &  n_n509  &  n_n534 ) ;
 assign wire11562 = ( wire256 ) | ( wire45 ) ;
 assign wire11563 = ( wire396 ) | ( n_n4596 ) | ( wire11560 ) ;
 assign wire11564 = ( wire13  &  n_n524  &  n_n464 ) | ( wire13  &  n_n464  &  n_n520 ) ;
 assign wire11566 = ( wire10  &  n_n524  &  n_n535 ) | ( wire10  &  n_n535  &  n_n520 ) ;
 assign wire11567 = ( wire25  &  n_n535  &  n_n390 ) | ( wire15  &  n_n535  &  n_n390 ) ;
 assign wire11568 = ( wire21  &  n_n535  &  n_n390 ) | ( wire23  &  n_n535  &  n_n390 ) ;
 assign wire11570 = ( n_n4593 ) | ( n_n4594 ) | ( wire365 ) ;
 assign wire11571 = ( wire11567 ) | ( wire11566 ) ;
 assign wire11574 = ( n_n4591 ) | ( n_n4592 ) | ( wire224 ) | ( wire11568 ) ;
 assign wire11575 = ( wire11562 ) | ( wire11563 ) | ( wire11570 ) | ( wire11571 ) ;
 assign wire11578 = ( n_n4537 ) | ( n_n4534 ) | ( wire11532 ) | ( wire11543 ) ;
 assign wire11579 = ( n_n4525 ) | ( n_n4528 ) | ( n_n4529 ) | ( wire11578 ) ;
 assign wire11581 = ( n_n1103 ) | ( wire11536 ) | ( wire11537 ) | ( wire11579 ) ;
 assign wire11582 = ( wire11558 ) | ( wire11559 ) | ( wire11574 ) | ( wire11575 ) ;
 assign wire11583 = ( wire16  &  n_n535  &  n_n532 ) | ( wire16  &  n_n535  &  n_n534 ) ;
 assign wire11584 = ( wire16  &  n_n526  &  n_n535 ) | ( wire16  &  n_n535  &  n_n528 ) ;
 assign wire11585 = ( wire22  &  n_n536  &  n_n535 ) | ( wire24  &  n_n536  &  n_n535 ) ;
 assign wire11586 = ( wire11584 ) | ( wire364 ) ;
 assign wire11587 = ( n_n4313 ) | ( wire11583 ) | ( wire11585 ) ;
 assign wire11588 = ( wire20  &  n_n536  &  n_n491 ) | ( wire15  &  n_n536  &  n_n491 ) ;
 assign wire11589 = ( wire16  &  n_n522  &  n_n491 ) | ( wire16  &  n_n524  &  n_n491 ) ;
 assign wire11591 = ( wire11588 ) | ( wire420 ) ;
 assign wire11592 = ( n_n4380 ) | ( n_n4379 ) | ( n_n4387 ) | ( wire11589 ) ;
 assign wire11593 = ( wire21  &  n_n536  &  n_n482 ) | ( wire23  &  n_n536  &  n_n482 ) ;
 assign wire11597 = ( n_n4404 ) | ( n_n4415 ) | ( wire11593 ) ;
 assign wire11598 = ( n_n4406 ) | ( n_n4408 ) | ( n_n4411 ) | ( wire328 ) ;
 assign wire11599 = ( wire16  &  n_n526  &  n_n482 ) | ( wire16  &  n_n482  &  n_n534 ) ;
 assign wire11600 = ( n_n4393 ) | ( wire23  &  n_n536  &  n_n491 ) ;
 assign wire11601 = ( n_n4401 ) | ( n_n4397 ) | ( n_n4402 ) ;
 assign wire11602 = ( n_n4396 ) | ( n_n4399 ) | ( wire11599 ) ;
 assign wire11605 = ( wire11591 ) | ( wire11592 ) | ( wire11597 ) | ( wire11598 ) ;
 assign wire11607 = ( i_9_  &  n_n536  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n536  &  n_n528  &  n_n500 ) ;
 assign wire11610 = ( n_n4356 ) | ( n_n4357 ) | ( n_n4358 ) ;
 assign wire11611 = ( wire67 ) | ( n_n4353 ) | ( n_n4354 ) ;
 assign wire11613 = ( n_n4360 ) | ( wire23  &  n_n536  &  n_n500 ) ;
 assign wire11614 = ( n_n4372 ) | ( n_n4371 ) | ( n_n4361 ) | ( n_n4359 ) ;
 assign wire11618 = ( n_n3533 ) | ( n_n1308 ) | ( wire282 ) | ( wire11613 ) ;
 assign wire11620 = ( i_9_  &  n_n536  &  n_n524  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n524  &  n_n518 ) ;
 assign wire11625 = ( n_n4337 ) | ( n_n4344 ) | ( n_n4345 ) | ( n_n4343 ) ;
 assign wire11626 = ( n_n4341 ) | ( n_n4342 ) | ( n_n4335 ) | ( wire11620 ) ;
 assign wire11628 = ( wire16  &  n_n528  &  n_n518 ) | ( wire16  &  n_n534  &  n_n518 ) ;
 assign wire11630 = ( n_n4327 ) | ( n_n4331 ) | ( n_n4329 ) | ( n_n4330 ) ;
 assign wire11631 = ( wire198 ) | ( n_n4322 ) | ( wire11628 ) ;
 assign wire11633 = ( wire11586 ) | ( wire11587 ) | ( wire11625 ) | ( wire11626 ) ;
 assign wire11634 = ( wire11630 ) | ( wire11631 ) | ( wire11633 ) ;
 assign wire11638 = ( wire10  &  n_n522  &  n_n491 ) | ( wire10  &  n_n528  &  n_n491 ) ;
 assign wire11641 = ( n_n4607 ) | ( n_n4641 ) | ( wire11638 ) ;
 assign wire11642 = ( n_n4633 ) | ( n_n4605 ) | ( n_n4632 ) | ( wire139 ) ;
 assign wire11646 = ( n_n4671 ) | ( n_n4672 ) | ( n_n4723 ) ;
 assign wire11647 = ( n_n4667 ) | ( n_n4703 ) | ( n_n4658 ) | ( wire775 ) ;
 assign wire11653 = ( n_n4601 ) | ( n_n4571 ) | ( n_n4587 ) | ( n_n4584 ) ;
 assign wire11654 = ( n_n4574 ) | ( n_n4550 ) | ( n_n4527 ) | ( wire99 ) ;
 assign wire11655 = ( wire11654 ) | ( wire11653 ) ;
 assign wire11658 = ( wire22  &  n_n536  &  n_n464 ) | ( wire23  &  n_n536  &  n_n464 ) ;
 assign wire11660 = ( n_n4455 ) | ( n_n4420 ) | ( n_n4430 ) | ( n_n4429 ) ;
 assign wire11661 = ( n_n4409 ) | ( n_n4410 ) | ( n_n4394 ) | ( wire11658 ) ;
 assign wire11666 = ( n_n4518 ) | ( n_n4500 ) | ( n_n4476 ) ;
 assign wire11667 = ( n_n4496 ) | ( n_n4505 ) | ( n_n4490 ) | ( n_n4477 ) ;
 assign wire11671 = ( wire15  &  n_n473  &  n_n325 ) | ( wire15  &  n_n482  &  n_n325 ) ;
 assign wire11675 = ( n_n4801 ) | ( n_n4778 ) | ( wire11671 ) ;
 assign wire11676 = ( n_n4773 ) | ( n_n4813 ) | ( n_n4742 ) | ( wire150 ) ;
 assign wire11677 = ( i_9_  &  n_n535  &  n_n528  &  n_n260 ) | ( (~ i_9_)  &  n_n535  &  n_n528  &  n_n260 ) ;
 assign wire11680 = ( n_n4834 ) | ( n_n4844 ) | ( n_n4833 ) ;
 assign wire11681 = ( n_n4857 ) | ( n_n4847 ) | ( wire11677 ) ;
 assign wire11687 = ( n_n4998 ) | ( n_n4887 ) | ( n_n4915 ) ;
 assign wire11688 = ( n_n4907 ) | ( n_n4879 ) | ( n_n4936 ) | ( n_n4947 ) ;
 assign wire11690 = ( n_n4967 ) | ( n_n4986 ) | ( wire11687 ) | ( wire11688 ) ;
 assign wire11693 = ( wire19  &  n_n526  &  n_n535 ) | ( wire19  &  n_n526  &  n_n518 ) ;
 assign wire11694 = ( wire19  &  n_n535  &  n_n528 ) | ( wire19  &  n_n535  &  n_n520 ) ;
 assign wire11698 = ( n_n5254 ) | ( n_n5218 ) | ( wire11694 ) ;
 assign wire11699 = ( n_n5248 ) | ( n_n5213 ) | ( n_n5227 ) | ( wire11693 ) ;
 assign wire11703 = ( wire11  &  n_n464  &  n_n130 ) | ( wire15  &  n_n464  &  n_n130 ) ;
 assign wire11705 = ( n_n5206 ) | ( n_n5186 ) | ( n_n5182 ) | ( n_n5172 ) ;
 assign wire11706 = ( n_n5191 ) | ( n_n5209 ) | ( n_n5192 ) | ( wire11703 ) ;
 assign wire11707 = ( wire12  &  n_n500  &  n_n520 ) | ( wire12  &  n_n500  &  n_n532 ) ;
 assign wire11710 = ( i_9_  &  n_n509  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n130 ) ;
 assign wire11712 = ( n_n5113 ) | ( n_n5155 ) | ( n_n5161 ) | ( n_n5127 ) ;
 assign wire11713 = ( n_n5108 ) | ( wire11707 ) | ( wire11710 ) ;
 assign wire11715 = ( wire11  &  n_n535  &  n_n130 ) | ( wire15  &  n_n535  &  n_n130 ) ;
 assign wire11718 = ( n_n5093 ) | ( n_n5054 ) | ( n_n5068 ) ;
 assign wire11719 = ( n_n5106 ) | ( n_n5070 ) | ( wire11715 ) ;
 assign wire11725 = ( n_n5040 ) | ( n_n4999 ) | ( n_n5024 ) ;
 assign wire11726 = ( n_n5025 ) | ( n_n5049 ) | ( n_n5047 ) | ( n_n5051 ) ;
 assign wire11731 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5307 ) | ( n_n5329 ) ;
 assign wire11732 = ( n_n5302 ) | ( n_n5335 ) | ( n_n5304 ) | ( n_n5289 ) ;
 assign wire11734 = ( wire11698 ) | ( wire11699 ) | ( wire11731 ) | ( wire11732 ) ;
 assign wire11735 = ( wire11705 ) | ( wire11706 ) | ( wire11712 ) | ( wire11713 ) ;
 assign wire11738 = ( wire16  &  n_n522  &  n_n535 ) | ( wire16  &  n_n522  &  n_n518 ) ;
 assign wire11739 = ( wire16  &  n_n526  &  n_n491 ) | ( wire16  &  n_n491  &  n_n520 ) ;
 assign wire11741 = ( wire11739 ) | ( wire11738 ) ;
 assign wire11743 = ( n_n4374 ) | ( n_n1002 ) | ( n_n4323 ) | ( wire11741 ) ;
 assign wire11745 = ( n_n956 ) | ( wire11660 ) | ( wire11661 ) | ( wire11743 ) ;
 assign wire11748 = ( wire14  &  n_n522  &  n_n491 ) | ( wire14  &  n_n491  &  n_n520 ) ;
 assign wire11751 = ( n_n4770 ) | ( n_n4769 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire11752 = ( n_n4767 ) | ( n_n4764 ) | ( n_n4771 ) | ( wire11748 ) ;
 assign wire11753 = ( wire14  &  n_n473  &  n_n526 ) | ( wire14  &  n_n473  &  n_n528 ) ;
 assign wire11754 = ( wire14  &  n_n473  &  n_n524 ) | ( wire14  &  n_n473  &  n_n520 ) ;
 assign wire11756 = ( n_n4810 ) | ( wire773 ) | ( wire11753 ) ;
 assign wire11757 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( wire11754 ) ;
 assign wire11759 = ( wire14  &  n_n524  &  n_n464 ) | ( wire14  &  n_n464  &  n_n520 ) ;
 assign wire11761 = ( n_n4816 ) | ( n_n4812 ) | ( n_n4811 ) | ( n_n4815 ) ;
 assign wire11762 = ( wire186 ) | ( wire85 ) | ( wire11759 ) ;
 assign wire11765 = ( n_n4787 ) | ( n_n4792 ) | ( n_n4793 ) | ( wire179 ) ;
 assign wire11766 = ( wire313 ) | ( wire292 ) | ( wire11765 ) ;
 assign wire11767 = ( wire11756 ) | ( wire11757 ) | ( wire11761 ) | ( wire11762 ) ;
 assign wire11768 = ( wire21  &  n_n518  &  n_n260 ) | ( wire22  &  n_n518  &  n_n260 ) ;
 assign wire11769 = ( wire21  &  n_n535  &  n_n260 ) | ( wire20  &  n_n535  &  n_n260 ) ;
 assign wire11772 = ( n_n4862 ) | ( wire245 ) | ( n_n4861 ) ;
 assign wire11773 = ( n_n4856 ) | ( wire102 ) | ( n_n4853 ) | ( n_n4860 ) ;
 assign wire11774 = ( wire24  &  n_n535  &  n_n260 ) | ( wire24  &  n_n518  &  n_n260 ) ;
 assign wire11776 = ( n_n4825 ) | ( n_n4848 ) | ( n_n4826 ) ;
 assign wire11777 = ( n_n4842 ) | ( n_n4841 ) | ( wire11774 ) ;
 assign wire11778 = ( n_n4845 ) | ( n_n4846 ) | ( n_n4852 ) | ( wire11768 ) ;
 assign wire11781 = ( n_n3820 ) | ( n_n4836 ) | ( wire11769 ) | ( wire11778 ) ;
 assign wire11782 = ( wire11772 ) | ( wire11773 ) | ( wire11776 ) | ( wire11777 ) ;
 assign wire11783 = ( wire17  &  n_n522  &  n_n482 ) | ( wire17  &  n_n530  &  n_n482 ) ;
 assign wire11785 = ( n_n4913 ) | ( wire352 ) | ( n_n4914 ) ;
 assign wire11786 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4905 ) | ( wire11783 ) ;
 assign wire11788 = ( wire17  &  n_n473  &  n_n524 ) | ( wire17  &  n_n473  &  n_n532 ) ;
 assign wire11790 = ( n_n4924 ) | ( n_n4921 ) | ( n_n4926 ) | ( n_n4925 ) ;
 assign wire11791 = ( n_n4920 ) | ( n_n4918 ) | ( n_n4919 ) | ( wire11788 ) ;
 assign wire11795 = ( n_n4937 ) | ( n_n4938 ) | ( n_n4931 ) | ( wire180 ) ;
 assign wire11796 = ( n_n4940 ) | ( n_n4939 ) | ( wire382 ) | ( wire11795 ) ;
 assign wire11797 = ( wire11785 ) | ( wire11786 ) | ( wire11790 ) | ( wire11791 ) ;
 assign wire11801 = ( n_n4963 ) | ( n_n4966 ) | ( wire771 ) | ( wire772 ) ;
 assign wire11802 = ( wire250 ) | ( n_n4968 ) | ( n_n4962 ) | ( n_n4971 ) ;
 assign wire11803 = ( wire17  &  n_n464  &  n_n528 ) | ( wire17  &  n_n464  &  n_n520 ) ;
 assign wire11804 = ( wire22  &  n_n464  &  n_n260 ) | ( wire11  &  n_n464  &  n_n260 ) ;
 assign wire11805 = ( wire17  &  n_n522  &  n_n464 ) | ( wire17  &  n_n524  &  n_n464 ) ;
 assign wire11807 = ( wire11804 ) | ( wire11803 ) ;
 assign wire11808 = ( n_n4955 ) | ( wire141 ) | ( wire11805 ) ;
 assign wire11809 = ( wire18  &  n_n528  &  n_n518 ) | ( wire18  &  n_n530  &  n_n518 ) ;
 assign wire11810 = ( wire22  &  n_n518  &  n_n195 ) | ( wire11  &  n_n518  &  n_n195 ) ;
 assign wire11811 = ( wire21  &  n_n518  &  n_n195 ) | ( wire20  &  n_n518  &  n_n195 ) ;
 assign wire11812 = ( wire18  &  n_n522  &  n_n518 ) | ( wire18  &  n_n524  &  n_n518 ) ;
 assign wire11814 = ( n_n4973 ) | ( wire11809 ) | ( wire11812 ) ;
 assign wire11815 = ( wire11810 ) | ( wire11811 ) | ( wire11814 ) ;
 assign wire11816 = ( wire11801 ) | ( wire11802 ) | ( wire11807 ) | ( wire11808 ) ;
 assign wire11818 = ( wire17  &  n_n524  &  n_n500 ) | ( wire17  &  n_n526  &  n_n500 ) ;
 assign wire11823 = ( wire295 ) | ( n_n4869 ) | ( n_n4870 ) ;
 assign wire11824 = ( wire40 ) | ( n_n4864 ) | ( n_n4867 ) | ( n_n4873 ) ;
 assign wire11825 = ( wire17  &  n_n524  &  n_n491 ) | ( wire17  &  n_n491  &  n_n520 ) ;
 assign wire11826 = ( wire20  &  n_n491  &  n_n260 ) | ( wire23  &  n_n491  &  n_n260 ) ;
 assign wire11829 = ( n_n4900 ) | ( n_n4899 ) | ( n_n4897 ) | ( wire11826 ) ;
 assign wire11830 = ( wire264 ) | ( wire11825 ) | ( wire11829 ) ;
 assign wire11832 = ( n_n1077 ) | ( wire11823 ) | ( wire11824 ) | ( wire11830 ) ;
 assign wire11833 = ( wire11796 ) | ( wire11797 ) | ( wire11815 ) | ( wire11816 ) ;
 assign wire11834 = ( i_9_  &  n_n522  &  n_n500  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n500  &  n_n325 ) ;
 assign wire11836 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire11837 = ( n_n4755 ) | ( n_n4759 ) | ( n_n4763 ) | ( wire11834 ) ;
 assign wire11839 = ( i_9_  &  n_n528  &  n_n500  &  n_n325 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n325 ) ;
 assign wire11841 = ( n_n4754 ) | ( n_n4753 ) | ( wire47 ) ;
 assign wire11842 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4745 ) | ( wire11839 ) ;
 assign wire11846 = ( n_n4732 ) | ( n_n4725 ) | ( n_n4726 ) | ( wire767 ) ;
 assign wire11847 = ( n_n4737 ) | ( n_n4738 ) | ( wire293 ) ;
 assign wire11848 = ( n_n4733 ) | ( n_n4728 ) | ( n_n4730 ) | ( n_n4743 ) ;
 assign wire11851 = ( wire95 ) | ( n_n4736 ) | ( wire457 ) | ( wire11848 ) ;
 assign wire11852 = ( wire11841 ) | ( wire11842 ) | ( wire11846 ) | ( wire11847 ) ;
 assign wire11855 = ( n_n4675 ) | ( n_n4676 ) | ( wire417 ) ;
 assign wire11856 = ( i_9_  &  n_n522  &  n_n390  &  n_n482 ) | ( (~ i_9_)  &  n_n522  &  n_n390  &  n_n482 ) ;
 assign wire11859 = ( n_n4673 ) | ( n_n4662 ) | ( wire157 ) ;
 assign wire11862 = ( n_n4685 ) | ( n_n4686 ) | ( n_n4695 ) | ( n_n4696 ) ;
 assign wire11866 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4716 ) ;
 assign wire11867 = ( n_n4711 ) | ( n_n4712 ) | ( wire173 ) ;
 assign wire11870 = ( wire22  &  n_n535  &  n_n325 ) | ( wire20  &  n_n535  &  n_n325 ) ;
 assign wire11873 = ( n_n4704 ) | ( n_n4697 ) | ( wire11870 ) ;
 assign wire11874 = ( n_n4707 ) | ( n_n4702 ) | ( n_n4700 ) | ( wire221 ) ;
 assign wire11877 = ( wire21  &  n_n390  &  n_n482 ) | ( wire25  &  n_n390  &  n_n482 ) ;
 assign wire11880 = ( wire81 ) | ( wire418 ) | ( wire11877 ) ;
 assign wire11881 = ( n_n4652 ) | ( wire140 ) | ( wire391 ) | ( wire431 ) ;
 assign wire11882 = ( n_n4674 ) | ( n_n4677 ) | ( wire11855 ) | ( wire11880 ) ;
 assign wire11884 = ( wire432 ) | ( wire11859 ) | ( wire11881 ) | ( wire11882 ) ;
 assign wire11886 = ( wire14  &  n_n524  &  n_n482 ) | ( wire14  &  n_n528  &  n_n482 ) ;
 assign wire11888 = ( n_n4784 ) | ( n_n4783 ) | ( wire315 ) ;
 assign wire11889 = ( n_n4779 ) | ( n_n4775 ) | ( n_n4780 ) | ( wire11886 ) ;
 assign wire11891 = ( wire11751 ) | ( wire11752 ) | ( wire11836 ) | ( wire11837 ) ;
 assign wire11893 = ( wire11766 ) | ( wire11767 ) | ( wire11781 ) | ( wire11782 ) ;
 assign wire11894 = ( wire11888 ) | ( wire11889 ) | ( wire11891 ) | ( wire11893 ) ;
 assign wire11899 = ( n_n5162 ) | ( n_n5154 ) | ( wire287 ) ;
 assign wire11900 = ( n_n5152 ) | ( wire406 ) | ( n_n5159 ) | ( n_n5160 ) ;
 assign wire11902 = ( wire22  &  n_n482  &  n_n130 ) | ( wire24  &  n_n482  &  n_n130 ) ;
 assign wire11906 = ( wire114 ) | ( wire44 ) | ( n_n5176 ) | ( wire765 ) ;
 assign wire11907 = ( wire33 ) | ( wire107 ) | ( wire113 ) | ( wire254 ) ;
 assign wire11908 = ( n_n5181 ) | ( n_n5173 ) | ( wire11902 ) | ( wire11906 ) ;
 assign wire11909 = ( wire11899 ) | ( wire11900 ) | ( wire11907 ) ;
 assign wire11912 = ( n_n5131 ) | ( n_n5132 ) | ( wire336 ) ;
 assign wire11914 = ( i_9_  &  n_n520  &  n_n518  &  n_n130 ) | ( (~ i_9_)  &  n_n520  &  n_n518  &  n_n130 ) ;
 assign wire11916 = ( wire12  &  n_n509  &  n_n526 ) | ( wire12  &  n_n509  &  n_n534 ) ;
 assign wire11917 = ( wire22  &  n_n509  &  n_n130 ) | ( wire15  &  n_n509  &  n_n130 ) ;
 assign wire11918 = ( wire11917 ) | ( wire11916 ) ;
 assign wire11921 = ( wire435 ) | ( wire318 ) ;
 assign wire11923 = ( wire19  &  n_n524  &  n_n500 ) | ( wire19  &  n_n526  &  n_n500 ) ;
 assign wire11924 = ( wire20  &  n_n500  &  n_n65 ) | ( wire25  &  n_n500  &  n_n65 ) ;
 assign wire11927 = ( wire62 ) | ( wire92 ) | ( wire11924 ) ;
 assign wire11928 = ( wire21  &  n_n491  &  n_n65 ) | ( wire23  &  n_n491  &  n_n65 ) ;
 assign wire11929 = ( n_n5288 ) | ( wire441 ) | ( n_n5286 ) ;
 assign wire11930 = ( n_n5281 ) | ( n_n5279 ) | ( n_n5280 ) | ( wire11928 ) ;
 assign wire11933 = ( wire333 ) | ( wire438 ) ;
 assign wire11939 = ( n_n5299 ) | ( n_n5290 ) | ( n_n5291 ) | ( wire63 ) ;
 assign wire11940 = ( n_n5293 ) | ( n_n5294 ) | ( wire200 ) | ( wire11939 ) ;
 assign wire11944 = ( n_n5305 ) | ( wire459 ) | ( n_n5306 ) ;
 assign wire11946 = ( wire24  &  n_n464  &  n_n65 ) | ( wire25  &  n_n464  &  n_n65 ) ;
 assign wire11947 = ( i_9_  &  n_n464  &  n_n528  &  n_n65 ) | ( (~ i_9_)  &  n_n464  &  n_n528  &  n_n65 ) ;
 assign wire11951 = ( n_n5322 ) | ( n_n5333 ) | ( n_n5319 ) | ( wire11946 ) ;
 assign wire11952 = ( wire148 ) | ( wire115 ) | ( wire175 ) | ( wire11947 ) ;
 assign wire11955 = ( wire24  &  n_n509  &  n_n65 ) | ( wire25  &  n_n509  &  n_n65 ) ;
 assign wire11959 = ( n_n5230 ) | ( n_n5233 ) | ( n_n5236 ) | ( wire320 ) ;
 assign wire11960 = ( n_n5240 ) | ( n_n5238 ) | ( wire11955 ) | ( wire11959 ) ;
 assign wire11962 = ( n_n1045 ) | ( wire11951 ) | ( wire11952 ) | ( wire11960 ) ;
 assign wire11964 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n535  &  n_n530 ) ;
 assign wire11967 = ( wire11964 ) | ( wire181 ) ;
 assign wire11968 = ( n_n5226 ) | ( n_n5225 ) | ( n_n5215 ) | ( wire384 ) ;
 assign wire11970 = ( n_n5189 ) | ( n_n5190 ) | ( wire452 ) ;
 assign wire11971 = ( n_n5200 ) | ( n_n5188 ) | ( n_n5194 ) | ( wire453 ) ;
 assign wire11972 = ( wire21  &  n_n464  &  n_n130 ) | ( wire23  &  n_n464  &  n_n130 ) ;
 assign wire11973 = ( wire19  &  n_n535  &  n_n532 ) | ( wire19  &  n_n535  &  n_n534 ) ;
 assign wire11975 = ( n_n5201 ) | ( wire761 ) | ( wire11972 ) ;
 assign wire11977 = ( wire220 ) | ( n_n5211 ) | ( wire11973 ) | ( wire11975 ) ;
 assign wire11978 = ( wire11967 ) | ( wire11968 ) | ( wire11970 ) | ( wire11971 ) ;
 assign wire11981 = ( wire299 ) | ( wire248 ) ;
 assign wire11982 = ( wire103 ) | ( n_n5003 ) | ( n_n4994 ) | ( n_n5006 ) ;
 assign wire11986 = ( n_n5017 ) | ( n_n5019 ) | ( n_n5010 ) | ( n_n5020 ) ;
 assign wire11987 = ( wire135 ) | ( n_n5012 ) | ( n_n5009 ) | ( n_n5007 ) ;
 assign wire11992 = ( n_n5050 ) | ( n_n5055 ) | ( n_n5059 ) | ( n_n5045 ) ;
 assign wire11993 = ( n_n5046 ) | ( n_n5056 ) | ( n_n5057 ) | ( wire166 ) ;
 assign wire11994 = ( wire18  &  n_n524  &  n_n491 ) | ( wire18  &  n_n528  &  n_n491 ) ;
 assign wire11995 = ( n_n5027 ) | ( n_n5028 ) | ( wire296 ) ;
 assign wire11996 = ( wire50 ) | ( n_n5029 ) | ( wire11994 ) ;
 assign wire11997 = ( wire18  &  n_n528  &  n_n482 ) | ( wire18  &  n_n482  &  n_n532 ) ;
 assign wire11999 = ( wire21  &  n_n482  &  n_n195 ) | ( wire22  &  n_n482  &  n_n195 ) ;
 assign wire12001 = ( n_n5035 ) | ( n_n5036 ) | ( wire11997 ) ;
 assign wire12003 = ( n_n5039 ) | ( wire253 ) | ( wire11999 ) | ( wire12001 ) ;
 assign wire12004 = ( wire11992 ) | ( wire11993 ) | ( wire11995 ) | ( wire11996 ) ;
 assign wire12007 = ( wire21  &  n_n518  &  n_n130 ) | ( wire20  &  n_n518  &  n_n130 ) ;
 assign wire12009 = ( n_n5096 ) | ( n_n5099 ) | ( wire12007 ) ;
 assign wire12014 = ( n_n5081 ) | ( n_n5089 ) | ( n_n5082 ) | ( n_n5084 ) ;
 assign wire12015 = ( n_n5078 ) | ( n_n5083 ) | ( wire232 ) | ( n_n5095 ) ;
 assign wire12018 = ( n_n5060 ) | ( n_n5067 ) | ( n_n5064 ) | ( wire755 ) ;
 assign wire12020 = ( n_n5069 ) | ( n_n5066 ) | ( n_n4152 ) | ( wire12018 ) ;
 assign wire12022 = ( n_n4990 ) | ( wire18  &  n_n520  &  n_n518 ) ;
 assign wire12023 = ( n_n4983 ) | ( n_n4985 ) | ( n_n4984 ) ;
 assign wire12024 = ( n_n4988 ) | ( n_n4987 ) | ( wire104 ) ;
 assign wire12027 = ( wire11981 ) | ( wire11982 ) | ( wire11986 ) | ( wire11987 ) ;
 assign wire12028 = ( wire12022 ) | ( wire12023 ) | ( wire12024 ) | ( wire12027 ) ;
 assign wire12033 = ( n_n5149 ) | ( n_n5138 ) | ( wire125 ) | ( n_n5143 ) ;
 assign wire12034 = ( wire211 ) | ( wire422 ) | ( wire12033 ) ;
 assign wire12036 = ( n_n1059 ) | ( wire28 ) | ( wire11918 ) | ( wire12034 ) ;
 assign wire12037 = ( wire11908 ) | ( wire11909 ) | ( wire11977 ) | ( wire11978 ) ;
 assign wire12040 = ( n_n1014 ) | ( wire11581 ) | ( wire11582 ) ;
 assign wire12041 = ( n_n4309 ) | ( n_n1040 ) | ( n_n1041 ) | ( wire11634 ) ;
 assign wire12047 = ( n_n4591 ) | ( n_n4592 ) | ( wire745 ) ;
 assign wire12048 = ( n_n4617 ) | ( n_n4618 ) | ( n_n4576 ) | ( n_n4569 ) ;
 assign wire12053 = ( n_n4491 ) | ( n_n4438 ) | ( wire184 ) ;
 assign wire12054 = ( wire70 ) | ( n_n4436 ) | ( n_n4458 ) | ( n_n4474 ) ;
 assign wire12058 = ( wire13  &  n_n526  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire12060 = ( n_n4546 ) | ( n_n4555 ) | ( n_n4562 ) | ( n_n4506 ) ;
 assign wire12061 = ( n_n4512 ) | ( n_n4526 ) | ( n_n4535 ) | ( wire12058 ) ;
 assign wire12062 = ( wire12061 ) | ( wire12060 ) ;
 assign wire12067 = ( n_n4764 ) | ( n_n4763 ) | ( n_n4751 ) ;
 assign wire12068 = ( n_n4737 ) | ( n_n4756 ) | ( n_n4724 ) | ( n_n4759 ) ;
 assign wire12074 = ( n_n4666 ) | ( n_n4649 ) | ( n_n4638 ) | ( n_n4655 ) ;
 assign wire12075 = ( n_n4658 ) | ( n_n4708 ) | ( n_n4706 ) | ( wire366 ) ;
 assign wire12080 = ( n_n4790 ) | ( n_n4835 ) | ( n_n4788 ) ;
 assign wire12081 = ( n_n4774 ) | ( n_n4845 ) | ( n_n4796 ) | ( n_n4822 ) ;
 assign wire12083 = ( n_n4823 ) | ( n_n4806 ) | ( wire12080 ) | ( wire12081 ) ;
 assign wire12089 = ( n_n4920 ) | ( n_n4907 ) | ( n_n4950 ) | ( n_n4894 ) ;
 assign wire12090 = ( n_n4916 ) | ( n_n4930 ) | ( n_n4947 ) | ( wire96 ) ;
 assign wire12091 = ( wire24  &  n_n500  &  n_n130 ) | ( wire25  &  n_n500  &  n_n130 ) ;
 assign wire12092 = ( i_9_  &  n_n526  &  n_n500  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n130 ) ;
 assign wire12093 = ( wire12  &  n_n464  &  n_n526 ) | ( wire12  &  n_n464  &  n_n520 ) ;
 assign wire12096 = ( wire12093 ) | ( wire12092 ) ;
 assign wire12097 = ( n_n5146 ) | ( n_n5204 ) | ( n_n5191 ) | ( wire12091 ) ;
 assign wire12099 = ( wire22  &  n_n535  &  n_n130 ) | ( wire25  &  n_n535  &  n_n130 ) ;
 assign wire12101 = ( n_n5096 ) | ( n_n5113 ) | ( n_n5066 ) | ( n_n5063 ) ;
 assign wire12102 = ( n_n5124 ) | ( wire335 ) | ( wire12099 ) ;
 assign wire12106 = ( wire19  &  n_n526  &  n_n535 ) | ( wire19  &  n_n535  &  n_n520 ) ;
 assign wire12108 = ( n_n5274 ) | ( n_n5232 ) | ( n_n5255 ) | ( n_n5267 ) ;
 assign wire12109 = ( n_n5244 ) | ( n_n5258 ) | ( n_n5212 ) | ( wire12106 ) ;
 assign wire12110 = ( wire12109 ) | ( wire12108 ) ;
 assign wire12111 = ( wire12096 ) | ( wire12097 ) | ( wire12101 ) | ( wire12102 ) ;
 assign wire12113 = ( wire18  &  n_n522  &  n_n491 ) | ( wire18  &  n_n528  &  n_n491 ) ;
 assign wire12114 = ( wire21  &  n_n482  &  n_n195 ) | ( wire20  &  n_n482  &  n_n195 ) ;
 assign wire12115 = ( wire22  &  n_n473  &  n_n195 ) | ( wire15  &  n_n473  &  n_n195 ) ;
 assign wire12117 = ( wire12114 ) | ( wire12113 ) ;
 assign wire12118 = ( n_n5025 ) | ( n_n5048 ) | ( n_n5009 ) | ( wire12115 ) ;
 assign wire12120 = ( wire18  &  n_n522  &  n_n518 ) | ( wire18  &  n_n528  &  n_n518 ) ;
 assign wire12122 = ( n_n4954 ) | ( wire771 ) | ( wire772 ) ;
 assign wire12123 = ( n_n4987 ) | ( n_n5005 ) | ( wire12120 ) ;
 assign wire12126 = ( wire19  &  n_n528  &  n_n482 ) | ( wire19  &  n_n520  &  n_n482 ) ;
 assign wire12128 = ( n_n5321 ) | ( n_n5326 ) | ( n_n5335 ) | ( wire12126 ) ;
 assign wire12129 = ( wire12089 ) | ( wire12090 ) | ( wire12128 ) ;
 assign wire12131 = ( n_n1333 ) | ( wire12117 ) | ( wire12118 ) | ( wire12129 ) ;
 assign wire12134 = ( wire22  &  n_n536  &  n_n473 ) | ( wire25  &  n_n536  &  n_n473 ) ;
 assign wire12136 = ( n_n4420 ) | ( n_n4407 ) | ( n_n4430 ) | ( n_n4404 ) ;
 assign wire12137 = ( wire84 ) | ( n_n4410 ) | ( wire12134 ) ;
 assign wire12141 = ( n_n4340 ) | ( n_n4345 ) | ( wire399 ) ;
 assign wire12142 = ( n_n4312 ) | ( n_n4331 ) | ( wire156 ) | ( n_n4326 ) ;
 assign wire12146 = ( n_n4400 ) | ( n_n4383 ) | ( n_n4369 ) | ( n_n4372 ) ;
 assign wire12147 = ( n_n4397 ) | ( n_n4360 ) | ( wire423 ) | ( n_n4375 ) ;
 assign wire12149 = ( wire12136 ) | ( wire12137 ) | ( wire12141 ) | ( wire12142 ) ;
 assign wire12150 = ( wire12146 ) | ( wire12147 ) | ( wire12149 ) ;
 assign wire12152 = ( wire12110 ) | ( wire12111 ) | ( wire12131 ) | ( wire12150 ) ;
 assign wire12156 = ( n_n4982 ) | ( wire134 ) | ( n_n4985 ) | ( n_n4986 ) ;
 assign wire12159 = ( n_n4998 ) | ( wire104 ) | ( wire743 ) ;
 assign wire12162 = ( wire22  &  n_n535  &  n_n195 ) | ( wire15  &  n_n535  &  n_n195 ) ;
 assign wire12164 = ( n_n4951 ) | ( n_n4952 ) | ( n_n4959 ) | ( n_n4960 ) ;
 assign wire12165 = ( wire250 ) | ( n_n4953 ) | ( wire12162 ) ;
 assign wire12166 = ( i_9_  &  n_n464  &  n_n528  &  n_n260 ) | ( (~ i_9_)  &  n_n464  &  n_n528  &  n_n260 ) ;
 assign wire12167 = ( wire24  &  n_n464  &  n_n260 ) | ( wire20  &  n_n464  &  n_n260 ) ;
 assign wire12168 = ( n_n4937 ) | ( n_n4938 ) | ( n_n4944 ) ;
 assign wire12169 = ( wire59 ) | ( wire12166 ) | ( wire12167 ) ;
 assign wire12170 = ( wire17  &  n_n473  &  n_n528 ) | ( wire17  &  n_n473  &  n_n520 ) ;
 assign wire12171 = ( wire17  &  n_n524  &  n_n464 ) | ( wire17  &  n_n464  &  n_n534 ) ;
 assign wire12172 = ( wire21  &  n_n473  &  n_n260 ) | ( wire20  &  n_n473  &  n_n260 ) ;
 assign wire12175 = ( wire31 ) | ( wire42 ) | ( wire12172 ) ;
 assign wire12176 = ( wire12170 ) | ( wire12171 ) | ( wire12175 ) ;
 assign wire12177 = ( wire12164 ) | ( wire12165 ) | ( wire12168 ) | ( wire12169 ) ;
 assign wire12179 = ( i_9_  &  n_n491  &  n_n532  &  n_n260 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n260 ) ;
 assign wire12181 = ( wire49 ) | ( wire260 ) ;
 assign wire12182 = ( n_n4888 ) | ( n_n4895 ) | ( n_n4889 ) | ( wire12179 ) ;
 assign wire12183 = ( wire22  &  n_n482  &  n_n260 ) | ( wire25  &  n_n482  &  n_n260 ) ;
 assign wire12186 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4901 ) | ( n_n4904 ) ;
 assign wire12187 = ( wire12183 ) | ( wire305 ) ;
 assign wire12188 = ( n_n4917 ) | ( n_n4914 ) | ( n_n4915 ) | ( n_n4910 ) ;
 assign wire12191 = ( n_n3810 ) | ( n_n1592 ) | ( wire12188 ) ;
 assign wire12192 = ( wire12181 ) | ( wire12182 ) | ( wire12186 ) | ( wire12187 ) ;
 assign wire12196 = ( n_n4964 ) | ( n_n4968 ) | ( wire342 ) | ( n_n4973 ) ;
 assign wire12197 = ( wire228 ) | ( wire362 ) | ( wire12196 ) ;
 assign wire12200 = ( wire12176 ) | ( wire12177 ) | ( wire12191 ) | ( wire12192 ) ;
 assign wire12202 = ( wire21  &  n_n482  &  n_n325 ) | ( wire20  &  n_n482  &  n_n325 ) ;
 assign wire12204 = ( n_n4784 ) | ( n_n4791 ) | ( wire158 ) ;
 assign wire12205 = ( wire179 ) | ( n_n4799 ) | ( wire12202 ) ;
 assign wire12207 = ( n_n4779 ) | ( n_n4775 ) | ( n_n4780 ) ;
 assign wire12208 = ( n_n4782 ) | ( n_n4781 ) | ( wire315 ) ;
 assign wire12210 = ( wire17  &  n_n509  &  n_n530 ) | ( wire17  &  n_n509  &  n_n534 ) ;
 assign wire12213 = ( wire12210 ) | ( wire277 ) ;
 assign wire12214 = ( wire245 ) | ( n_n4864 ) | ( n_n4854 ) | ( n_n4865 ) ;
 assign wire12217 = ( wire21  &  n_n509  &  n_n260 ) | ( wire23  &  n_n509  &  n_n260 ) ;
 assign wire12218 = ( n_n4882 ) | ( n_n4881 ) | ( wire330 ) ;
 assign wire12219 = ( n_n4868 ) | ( n_n4880 ) | ( wire324 ) ;
 assign wire12220 = ( n_n4877 ) | ( n_n4870 ) | ( wire12217 ) ;
 assign wire12223 = ( n_n1985 ) | ( n_n3815 ) | ( wire12220 ) ;
 assign wire12224 = ( wire12213 ) | ( wire12214 ) | ( wire12218 ) | ( wire12219 ) ;
 assign wire12225 = ( i_9_  &  n_n464  &  n_n530  &  n_n325 ) | ( (~ i_9_)  &  n_n464  &  n_n530  &  n_n325 ) ;
 assign wire12226 = ( i_9_  &  n_n535  &  n_n528  &  n_n260 ) | ( (~ i_9_)  &  n_n535  &  n_n528  &  n_n260 ) ;
 assign wire12230 = ( n_n4827 ) | ( n_n4828 ) | ( wire12226 ) ;
 assign wire12231 = ( n_n4833 ) | ( n_n4838 ) | ( wire304 ) | ( wire735 ) ;
 assign wire12232 = ( wire22  &  n_n518  &  n_n260 ) | ( wire24  &  n_n518  &  n_n260 ) ;
 assign wire12234 = ( n_n4842 ) | ( n_n4851 ) | ( n_n4841 ) ;
 assign wire12235 = ( wire12232 ) | ( wire52 ) ;
 assign wire12239 = ( n_n4817 ) | ( n_n4824 ) | ( wire85 ) | ( wire12225 ) ;
 assign wire12240 = ( n_n4825 ) | ( wire186 ) | ( n_n4826 ) | ( wire12239 ) ;
 assign wire12243 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( n_n4808 ) ;
 assign wire12245 = ( n_n4802 ) | ( n_n4805 ) | ( n_n4197 ) | ( wire12243 ) ;
 assign wire12247 = ( n_n1472 ) | ( wire12204 ) | ( wire12205 ) | ( wire12245 ) ;
 assign wire12252 = ( wire296 ) | ( n_n5019 ) | ( n_n5020 ) ;
 assign wire12253 = ( n_n5026 ) | ( n_n5017 ) | ( wire135 ) | ( n_n5016 ) ;
 assign wire12255 = ( wire18  &  n_n522  &  n_n500 ) | ( wire18  &  n_n524  &  n_n500 ) ;
 assign wire12256 = ( wire21  &  n_n500  &  n_n195 ) | ( wire20  &  n_n500  &  n_n195 ) ;
 assign wire12257 = ( n_n5008 ) | ( wire11  &  n_n500  &  n_n195 ) ;
 assign wire12261 = ( wire406 ) | ( wire358 ) ;
 assign wire12262 = ( n_n5157 ) | ( n_n5152 ) | ( n_n5149 ) | ( wire195 ) ;
 assign wire12265 = ( wire288 ) | ( wire211 ) ;
 assign wire12266 = ( n_n5135 ) | ( n_n5148 ) | ( wire125 ) | ( n_n5144 ) ;
 assign wire12268 = ( wire22  &  n_n464  &  n_n130 ) | ( wire11  &  n_n464  &  n_n130 ) ;
 assign wire12269 = ( wire21  &  n_n464  &  n_n130 ) | ( wire15  &  n_n464  &  n_n130 ) ;
 assign wire12271 = ( wire12268 ) | ( wire453 ) ;
 assign wire12272 = ( wire452 ) | ( n_n5192 ) | ( wire12269 ) ;
 assign wire12276 = ( n_n5234 ) | ( wire21  &  n_n535  &  n_n65 ) ;
 assign wire12277 = ( n_n5207 ) | ( n_n5208 ) | ( n_n5205 ) ;
 assign wire12278 = ( n_n5230 ) | ( n_n5223 ) | ( n_n5233 ) | ( n_n5220 ) ;
 assign wire12282 = ( n_n1530 ) | ( n_n1532 ) | ( n_n763 ) | ( wire12276 ) ;
 assign wire12283 = ( wire12271 ) | ( wire12272 ) | ( wire12277 ) | ( wire12278 ) ;
 assign wire12285 = ( i_9_  &  n_n528  &  n_n482  &  n_n130 ) | ( (~ i_9_)  &  n_n528  &  n_n482  &  n_n130 ) ;
 assign wire12287 = ( wire437 ) | ( wire168 ) ;
 assign wire12288 = ( n_n5163 ) | ( wire33 ) | ( wire12285 ) ;
 assign wire12290 = ( wire21  &  n_n473  &  n_n130 ) | ( wire25  &  n_n473  &  n_n130 ) ;
 assign wire12291 = ( wire113 ) | ( wire114 ) ;
 assign wire12292 = ( n_n5189 ) | ( n_n5190 ) | ( wire332 ) ;
 assign wire12293 = ( n_n5171 ) | ( n_n5186 ) | ( wire12290 ) ;
 assign wire12296 = ( n_n4129 ) | ( wire44 ) | ( n_n5176 ) | ( wire12293 ) ;
 assign wire12297 = ( wire12287 ) | ( wire12288 ) | ( wire12291 ) | ( wire12292 ) ;
 assign wire12299 = ( n_n5127 ) | ( wire12  &  n_n500  &  n_n530 ) ;
 assign wire12300 = ( n_n5128 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire12301 = ( n_n5130 ) | ( n_n5120 ) | ( wire286 ) ;
 assign wire12304 = ( wire12261 ) | ( wire12262 ) | ( wire12265 ) | ( wire12266 ) ;
 assign wire12305 = ( wire12299 ) | ( wire12300 ) | ( wire12301 ) | ( wire12304 ) ;
 assign wire12306 = ( wire12282 ) | ( wire12283 ) | ( wire12296 ) | ( wire12297 ) ;
 assign wire12309 = ( n_n5064 ) | ( n_n5058 ) | ( wire755 ) ;
 assign wire12310 = ( n_n5060 ) | ( n_n5055 ) | ( n_n5059 ) | ( n_n5056 ) ;
 assign wire12315 = ( n_n5054 ) | ( n_n5042 ) | ( wire97 ) ;
 assign wire12316 = ( wire356 ) | ( n_n5049 ) | ( n_n5039 ) | ( n_n5052 ) ;
 assign wire12317 = ( wire22  &  n_n464  &  n_n195 ) | ( wire15  &  n_n464  &  n_n195 ) ;
 assign wire12318 = ( wire18  &  n_n524  &  n_n464 ) | ( wire18  &  n_n464  &  n_n526 ) ;
 assign wire12319 = ( wire18  &  n_n522  &  n_n464 ) | ( wire18  &  n_n464  &  n_n528 ) ;
 assign wire12323 = ( n_n5075 ) | ( n_n5068 ) | ( n_n5071 ) | ( wire12317 ) ;
 assign wire12324 = ( wire12318 ) | ( wire12319 ) | ( wire12323 ) ;
 assign wire12326 = ( wire24  &  n_n509  &  n_n130 ) | ( wire15  &  n_n509  &  n_n130 ) ;
 assign wire12327 = ( n_n5112 ) | ( n_n5110 ) | ( wire414 ) ;
 assign wire12328 = ( n_n5109 ) | ( n_n5107 ) | ( n_n5108 ) | ( wire12326 ) ;
 assign wire12332 = ( n_n5087 ) | ( n_n5088 ) | ( n_n5077 ) ;
 assign wire12333 = ( n_n5085 ) | ( n_n5082 ) | ( n_n5084 ) | ( n_n5079 ) ;
 assign wire12335 = ( wire21  &  n_n535  &  n_n130 ) | ( wire20  &  n_n535  &  n_n130 ) ;
 assign wire12337 = ( n_n5098 ) | ( n_n5095 ) | ( wire88 ) ;
 assign wire12338 = ( wire12335 ) | ( wire289 ) ;
 assign wire12340 = ( n_n5100 ) | ( n_n5103 ) | ( wire12337 ) | ( wire12338 ) ;
 assign wire12342 = ( wire11  &  n_n482  &  n_n65 ) | ( wire15  &  n_n482  &  n_n65 ) ;
 assign wire12344 = ( n_n5297 ) | ( n_n5291 ) | ( n_n5292 ) | ( n_n5298 ) ;
 assign wire12345 = ( n_n5288 ) | ( n_n5290 ) | ( n_n5289 ) | ( wire12342 ) ;
 assign wire12349 = ( n_n5251 ) | ( wire435 ) | ( n_n5257 ) | ( n_n5247 ) ;
 assign wire12352 = ( n_n5241 ) | ( n_n5242 ) | ( n_n5246 ) ;
 assign wire12353 = ( n_n5240 ) | ( n_n5245 ) | ( wire320 ) ;
 assign wire12355 = ( wire19  &  n_n528  &  n_n500 ) | ( wire19  &  n_n500  &  n_n530 ) ;
 assign wire12356 = ( i_9_  &  n_n526  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n65 ) ;
 assign wire12358 = ( n_n5272 ) | ( n_n5271 ) | ( n_n5270 ) | ( wire12356 ) ;
 assign wire12359 = ( wire77 ) | ( wire12355 ) | ( wire12358 ) ;
 assign wire12361 = ( wire11  &  n_n464  &  n_n65 ) | ( wire24  &  n_n464  &  n_n65 ) ;
 assign wire12363 = ( wire175 ) | ( wire149 ) ;
 assign wire12364 = ( n_n5333 ) | ( n_n5330 ) | ( wire12361 ) ;
 assign wire12366 = ( wire11  &  n_n473  &  n_n65 ) | ( wire15  &  n_n473  &  n_n65 ) ;
 assign wire12368 = ( n_n5314 ) | ( n_n5322 ) | ( wire115 ) ;
 assign wire12369 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5312 ) | ( wire12366 ) ;
 assign wire12371 = ( i_9_  &  n_n528  &  n_n491  &  n_n65 ) | ( (~ i_9_)  &  n_n528  &  n_n491  &  n_n65 ) ;
 assign wire12372 = ( wire24  &  n_n491  &  n_n65 ) | ( wire25  &  n_n491  &  n_n65 ) ;
 assign wire12374 = ( n_n5305 ) | ( wire21  &  n_n482  &  n_n65 ) ;
 assign wire12375 = ( wire218 ) | ( wire19  &  n_n491  &  n_n520 ) ;
 assign wire12376 = ( n_n5303 ) | ( wire63 ) | ( n_n5304 ) ;
 assign wire12380 = ( wire12344 ) | ( wire12345 ) | ( wire12375 ) | ( wire12376 ) ;
 assign wire12381 = ( n_n3019 ) | ( n_n1402 ) | ( wire204 ) | ( wire12374 ) ;
 assign wire12382 = ( n_n1435 ) | ( n_n1436 ) | ( wire12359 ) | ( wire12380 ) ;
 assign wire12384 = ( wire20  &  n_n491  &  n_n195 ) | ( wire23  &  n_n491  &  n_n195 ) ;
 assign wire12386 = ( n_n5038 ) | ( n_n5035 ) | ( n_n5037 ) | ( wire12384 ) ;
 assign wire12387 = ( n_n5034 ) | ( n_n5027 ) | ( wire253 ) | ( wire12386 ) ;
 assign wire12389 = ( n_n1454 ) | ( wire12252 ) | ( wire12253 ) | ( wire12387 ) ;
 assign wire12391 = ( n_n1409 ) | ( n_n1408 ) | ( wire12389 ) ;
 assign wire12392 = ( wire12305 ) | ( wire12306 ) | ( wire12381 ) | ( wire12382 ) ;
 assign wire12393 = ( i_9_  &  n_n522  &  n_n491  &  n_n325 ) | ( (~ i_9_)  &  n_n522  &  n_n491  &  n_n325 ) ;
 assign wire12395 = ( n_n4765 ) | ( n_n4766 ) | ( n_n4762 ) ;
 assign wire12398 = ( i_9_  &  n_n509  &  n_n522  &  n_n325 ) | ( (~ i_9_)  &  n_n509  &  n_n522  &  n_n325 ) ;
 assign wire12399 = ( n_n4738 ) | ( n_n4744 ) | ( n_n4739 ) | ( n_n4745 ) ;
 assign wire12400 = ( wire95 ) | ( n_n4736 ) | ( wire12398 ) ;
 assign wire12401 = ( wire11  &  n_n535  &  n_n325 ) | ( wire25  &  n_n535  &  n_n325 ) ;
 assign wire12403 = ( n_n4695 ) | ( n_n4696 ) | ( n_n4700 ) ;
 assign wire12404 = ( wire12401 ) | ( wire221 ) ;
 assign wire12408 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4721 ) ;
 assign wire12409 = ( n_n4720 ) | ( n_n4727 ) | ( n_n4729 ) | ( n_n4719 ) ;
 assign wire12413 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4713 ) ;
 assign wire12414 = ( n_n4704 ) | ( n_n4711 ) | ( n_n4710 ) | ( n_n4709 ) ;
 assign wire12416 = ( n_n4715 ) | ( n_n4716 ) | ( wire12413 ) | ( wire12414 ) ;
 assign wire12420 = ( n_n4673 ) | ( n_n4670 ) | ( wire417 ) ;
 assign wire12421 = ( n_n4674 ) | ( n_n4671 ) | ( wire81 ) | ( wire418 ) ;
 assign wire12422 = ( wire10  &  n_n522  &  n_n464 ) | ( wire10  &  n_n464  &  n_n520 ) ;
 assign wire12425 = ( wire225 ) | ( wire157 ) ;
 assign wire12426 = ( n_n4667 ) | ( n_n4662 ) | ( n_n4660 ) | ( wire72 ) ;
 assign wire12428 = ( wire11  &  n_n464  &  n_n390 ) | ( wire15  &  n_n464  &  n_n390 ) ;
 assign wire12429 = ( n_n4689 ) | ( n_n4684 ) | ( wire444 ) ;
 assign wire12431 = ( n_n4693 ) | ( wire12422 ) | ( wire12428 ) | ( wire12429 ) ;
 assign wire12432 = ( wire12420 ) | ( wire12421 ) | ( wire12425 ) | ( wire12426 ) ;
 assign wire12434 = ( n_n4755 ) | ( wire14  &  n_n526  &  n_n500 ) ;
 assign wire12435 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4761 ) ;
 assign wire12436 = ( n_n4754 ) | ( n_n4757 ) | ( n_n4749 ) | ( n_n4760 ) ;
 assign wire12439 = ( wire447 ) | ( wire12395 ) | ( wire12399 ) | ( wire12400 ) ;
 assign wire12440 = ( wire12434 ) | ( wire12435 ) | ( wire12436 ) | ( wire12439 ) ;
 assign wire12442 = ( wire21  &  n_n536  &  n_n500 ) | ( wire20  &  n_n536  &  n_n500 ) ;
 assign wire12445 = ( n_n4367 ) | ( n_n4368 ) | ( wire12442 ) ;
 assign wire12446 = ( wire280 ) | ( n_n4365 ) | ( n_n4374 ) | ( n_n4370 ) ;
 assign wire12447 = ( i_9_  &  n_n536  &  n_n526  &  n_n491 ) | ( (~ i_9_)  &  n_n536  &  n_n526  &  n_n491 ) ;
 assign wire12448 = ( wire16  &  n_n522  &  n_n491 ) | ( wire16  &  n_n491  &  n_n520 ) ;
 assign wire12449 = ( wire16  &  n_n528  &  n_n491 ) | ( wire16  &  n_n491  &  n_n530 ) ;
 assign wire12451 = ( n_n4356 ) | ( n_n4357 ) | ( n_n4355 ) | ( n_n4358 ) ;
 assign wire12453 = ( n_n4386 ) | ( n_n4387 ) | ( wire12447 ) | ( wire12448 ) ;
 assign wire12455 = ( n_n4361 ) | ( n_n3533 ) | ( n_n4348 ) | ( wire12453 ) ;
 assign wire12456 = ( wire27 ) | ( wire12445 ) | ( wire12446 ) | ( wire12451 ) ;
 assign wire12458 = ( n_n4405 ) | ( n_n4406 ) | ( n_n4408 ) ;
 assign wire12459 = ( n_n4411 ) | ( n_n4412 ) | ( wire79 ) ;
 assign wire12461 = ( wire16  &  n_n528  &  n_n482 ) | ( wire16  &  n_n482  &  n_n534 ) ;
 assign wire12464 = ( n_n4393 ) | ( wire37 ) | ( n_n4394 ) ;
 assign wire12465 = ( n_n4401 ) | ( n_n4396 ) | ( n_n4395 ) | ( n_n4402 ) ;
 assign wire12467 = ( wire98 ) | ( n_n4421 ) | ( wire215 ) | ( n_n4429 ) ;
 assign wire12469 = ( n_n4399 ) | ( n_n4428 ) | ( wire12461 ) | ( wire12467 ) ;
 assign wire12471 = ( i_9_  &  n_n455  &  n_n530  &  n_n518 ) | ( (~ i_9_)  &  n_n455  &  n_n530  &  n_n518 ) ;
 assign wire12472 = ( wire13  &  n_n535  &  n_n530 ) | ( wire13  &  n_n535  &  n_n534 ) ;
 assign wire12475 = ( n_n4445 ) | ( n_n4446 ) | ( wire12472 ) ;
 assign wire12476 = ( n_n4437 ) | ( n_n4447 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire12478 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign wire12479 = ( n_n4451 ) | ( wire13  &  n_n526  &  n_n535 ) ;
 assign wire12480 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4465 ) ;
 assign wire12481 = ( wire12478 ) | ( wire128 ) ;
 assign wire12485 = ( n_n3162 ) | ( wire55 ) | ( n_n2058 ) | ( wire12479 ) ;
 assign wire12486 = ( wire12475 ) | ( wire12476 ) | ( wire12480 ) | ( wire12481 ) ;
 assign wire12488 = ( wire22  &  n_n455  &  n_n500 ) | ( wire15  &  n_n455  &  n_n500 ) ;
 assign wire12489 = ( n_n4489 ) | ( wire66 ) | ( n_n4490 ) ;
 assign wire12490 = ( n_n4487 ) | ( n_n4488 ) | ( n_n4486 ) | ( wire12488 ) ;
 assign wire12492 = ( n_n4477 ) | ( n_n4475 ) | ( n_n4476 ) ;
 assign wire12493 = ( n_n4470 ) | ( n_n4469 ) | ( wire199 ) ;
 assign wire12497 = ( wire201 ) | ( wire416 ) ;
 assign wire12498 = ( n_n4547 ) | ( n_n4538 ) | ( wire212 ) | ( n_n4545 ) ;
 assign wire12499 = ( wire21  &  n_n455  &  n_n482 ) | ( wire25  &  n_n455  &  n_n482 ) ;
 assign wire12500 = ( i_9_  &  n_n473  &  n_n455  &  n_n534 ) | ( (~ i_9_)  &  n_n473  &  n_n455  &  n_n534 ) ;
 assign wire12501 = ( wire13  &  n_n526  &  n_n482 ) | ( wire13  &  n_n520  &  n_n482 ) ;
 assign wire12502 = ( wire170 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire12503 = ( wire12499 ) | ( wire361 ) ;
 assign wire12507 = ( n_n4247 ) | ( n_n3879 ) | ( wire12500 ) | ( wire12501 ) ;
 assign wire12508 = ( wire12497 ) | ( wire12498 ) | ( wire12502 ) | ( wire12503 ) ;
 assign wire12510 = ( wire24  &  n_n455  &  n_n491 ) | ( wire15  &  n_n455  &  n_n491 ) ;
 assign wire12514 = ( wire308 ) | ( n_n4505 ) | ( n_n4501 ) | ( n_n4499 ) ;
 assign wire12515 = ( n_n4504 ) | ( n_n4503 ) | ( wire12510 ) | ( wire12514 ) ;
 assign wire12517 = ( n_n1496 ) | ( wire12489 ) | ( wire12490 ) | ( wire12515 ) ;
 assign wire12518 = ( wire12485 ) | ( wire12486 ) | ( wire12507 ) | ( wire12508 ) ;
 assign wire12519 = ( i_9_  &  n_n509  &  n_n528  &  n_n390 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n390 ) ;
 assign wire12520 = ( i_9_  &  n_n390  &  n_n532  &  n_n518 ) | ( (~ i_9_)  &  n_n390  &  n_n532  &  n_n518 ) ;
 assign wire12521 = ( i_9_  &  n_n535  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n535  &  n_n390  &  n_n532 ) ;
 assign wire12524 = ( wire12521 ) | ( n_n464  &  n_n455  &  wire600 ) ;
 assign wire12525 = ( n_n4561 ) | ( n_n4568 ) | ( n_n4572 ) | ( wire238 ) ;
 assign wire12529 = ( wire276 ) | ( wire213 ) ;
 assign wire12530 = ( n_n4557 ) | ( n_n4560 ) | ( n_n4582 ) | ( n_n4581 ) ;
 assign wire12531 = ( n_n4554 ) | ( n_n4584 ) | ( n_n4577 ) | ( n_n4556 ) ;
 assign wire12534 = ( n_n3871 ) | ( n_n4585 ) | ( wire12520 ) | ( wire12531 ) ;
 assign wire12535 = ( wire12524 ) | ( wire12525 ) | ( wire12529 ) | ( wire12530 ) ;
 assign wire12539 = ( n_n4616 ) | ( n_n4612 ) | ( n_n4611 ) | ( n_n4619 ) ;
 assign wire12540 = ( n_n4608 ) | ( wire465 ) | ( n_n4620 ) | ( n_n4609 ) ;
 assign wire12541 = ( wire10  &  n_n528  &  n_n518 ) | ( wire10  &  n_n520  &  n_n518 ) ;
 assign wire12543 = ( n_n4593 ) | ( n_n4594 ) | ( wire255 ) ;
 assign wire12544 = ( wire365 ) | ( n_n4595 ) | ( wire12541 ) ;
 assign wire12545 = ( wire10  &  n_n524  &  n_n500 ) | ( wire10  &  n_n526  &  n_n500 ) ;
 assign wire12546 = ( i_9_  &  n_n522  &  n_n500  &  n_n390 ) | ( (~ i_9_)  &  n_n522  &  n_n500  &  n_n390 ) ;
 assign wire12547 = ( wire25  &  n_n491  &  n_n390 ) | ( wire15  &  n_n491  &  n_n390 ) ;
 assign wire12551 = ( n_n4648 ) | ( n_n4646 ) | ( wire391 ) ;
 assign wire12552 = ( n_n4644 ) | ( wire311 ) | ( n_n4650 ) | ( n_n4654 ) ;
 assign wire12554 = ( n_n4630 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign wire12555 = ( wire401 ) | ( wire310 ) ;
 assign wire12556 = ( n_n4640 ) | ( n_n4621 ) | ( n_n4625 ) | ( wire12545 ) ;
 assign wire12557 = ( n_n4639 ) | ( n_n4627 ) | ( wire12546 ) | ( wire12547 ) ;
 assign wire12559 = ( wire12557 ) | ( wire12556 ) ;
 assign wire12560 = ( wire12551 ) | ( wire12552 ) | ( wire12554 ) | ( wire12555 ) ;
 assign wire12561 = ( i_9_  &  n_n509  &  n_n390  &  n_n534 ) | ( (~ i_9_)  &  n_n509  &  n_n390  &  n_n534 ) ;
 assign wire12564 = ( n_n4605 ) | ( n_n4603 ) | ( n_n4599 ) | ( wire12519 ) ;
 assign wire12566 = ( wire12539 ) | ( wire12540 ) | ( wire12543 ) | ( wire12544 ) ;
 assign wire12567 = ( wire256 ) | ( wire12561 ) | ( wire12564 ) | ( wire12566 ) ;
 assign wire12568 = ( wire12534 ) | ( wire12535 ) | ( wire12559 ) | ( wire12560 ) ;
 assign wire12569 = ( wire16  &  n_n522  &  n_n535 ) | ( wire16  &  n_n524  &  n_n535 ) ;
 assign wire12570 = ( i_9_  &  n_n536  &  n_n526  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n526  &  n_n518 ) ;
 assign wire12572 = ( wire53 ) | ( wire67 ) ;
 assign wire12573 = ( n_n4344 ) | ( n_n4341 ) | ( n_n4335 ) | ( wire12570 ) ;
 assign wire12574 = ( wire16  &  n_n526  &  n_n535 ) | ( wire16  &  n_n535  &  n_n528 ) ;
 assign wire12576 = ( wire364 ) | ( wire283 ) ;
 assign wire12577 = ( wire171 ) | ( n_n4313 ) | ( wire12574 ) ;
 assign wire12578 = ( wire16  &  n_n530  &  n_n518 ) | ( wire16  &  n_n534  &  n_n518 ) ;
 assign wire12579 = ( n_n4329 ) | ( wire106 ) | ( n_n4330 ) ;
 assign wire12580 = ( n_n4323 ) | ( wire12569 ) | ( wire12578 ) ;
 assign wire12582 = ( wire12572 ) | ( wire12573 ) | ( wire12576 ) | ( wire12577 ) ;
 assign wire12583 = ( wire12579 ) | ( wire12580 ) | ( wire12582 ) ;
 assign wire12585 = ( n_n1426 ) | ( wire12455 ) | ( wire12456 ) | ( wire12583 ) ;
 assign wire12586 = ( wire12517 ) | ( wire12518 ) | ( wire12567 ) | ( wire12568 ) ;
 assign wire12588 = ( n_n1398 ) | ( n_n1326 ) | ( n_n1325 ) | ( wire12152 ) ;
 assign wire12589 = ( n_n1396 ) | ( n_n1397 ) | ( wire12391 ) | ( wire12392 ) ;
 assign wire12595 = ( n_n4597 ) | ( n_n4601 ) | ( n_n4631 ) ;
 assign wire12596 = ( n_n4578 ) | ( n_n4611 ) | ( n_n4633 ) | ( n_n4581 ) ;
 assign wire12600 = ( wire310 ) | ( wire139 ) ;
 assign wire12601 = ( n_n4648 ) | ( n_n4635 ) | ( wire140 ) | ( n_n4645 ) ;
 assign wire12602 = ( wire24  &  n_n473  &  n_n455 ) | ( wire24  &  n_n455  &  n_n482 ) ;
 assign wire12607 = ( n_n4557 ) | ( n_n4572 ) | ( n_n4531 ) | ( n_n4555 ) ;
 assign wire12608 = ( n_n4528 ) | ( n_n4549 ) | ( n_n4559 ) | ( wire12602 ) ;
 assign wire12609 = ( wire12608 ) | ( wire12607 ) ;
 assign wire12613 = ( n_n4756 ) | ( n_n4753 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire12614 = ( wire131 ) | ( n_n4792 ) | ( n_n4764 ) | ( n_n4763 ) ;
 assign wire12615 = ( wire10  &  n_n473  &  n_n528 ) | ( wire10  &  n_n473  &  n_n530 ) ;
 assign wire12620 = ( n_n4656 ) | ( n_n4676 ) | ( n_n4703 ) | ( n_n4698 ) ;
 assign wire12621 = ( n_n4672 ) | ( n_n4692 ) | ( n_n4686 ) | ( wire12615 ) ;
 assign wire12626 = ( n_n4735 ) | ( n_n4749 ) | ( n_n4740 ) ;
 assign wire12627 = ( n_n4727 ) | ( n_n4733 ) | ( n_n4730 ) | ( n_n4718 ) ;
 assign wire12629 = ( n_n4750 ) | ( n_n4736 ) | ( wire12626 ) | ( wire12627 ) ;
 assign wire12630 = ( wire12613 ) | ( wire12614 ) | ( wire12620 ) | ( wire12621 ) ;
 assign wire12634 = ( n_n5258 ) | ( n_n5212 ) | ( n_n5262 ) | ( n_n5259 ) ;
 assign wire12635 = ( n_n5266 ) | ( n_n5236 ) | ( n_n5235 ) | ( wire320 ) ;
 assign wire12638 = ( wire12  &  n_n526  &  n_n482 ) | ( wire12  &  n_n528  &  n_n482 ) ;
 assign wire12640 = ( n_n5183 ) | ( n_n5204 ) | ( n_n5182 ) | ( n_n5173 ) ;
 assign wire12641 = ( wire114 ) | ( n_n5211 ) | ( wire12638 ) ;
 assign wire12642 = ( wire21  &  n_n509  &  n_n130 ) | ( wire21  &  n_n491  &  n_n130 ) ;
 assign wire12643 = ( wire15  &  n_n509  &  n_n130 ) | ( wire15  &  n_n482  &  n_n130 ) ;
 assign wire12648 = ( n_n5121 ) | ( n_n5134 ) | ( n_n5151 ) | ( wire12642 ) ;
 assign wire12649 = ( n_n5135 ) | ( n_n5158 ) | ( wire12643 ) | ( wire12648 ) ;
 assign wire12650 = ( wire12634 ) | ( wire12635 ) | ( wire12640 ) | ( wire12641 ) ;
 assign wire12651 = ( wire12  &  n_n530  &  n_n518 ) | ( wire12  &  n_n534  &  n_n518 ) ;
 assign wire12653 = ( wire22  &  n_n518  &  n_n130 ) | ( wire11  &  n_n518  &  n_n130 ) ;
 assign wire12656 = ( n_n5089 ) | ( n_n5098 ) | ( wire12653 ) ;
 assign wire12657 = ( n_n5104 ) | ( n_n5078 ) | ( n_n5090 ) | ( wire12651 ) ;
 assign wire12658 = ( wire18  &  n_n509  &  n_n526 ) | ( wire18  &  n_n526  &  n_n518 ) ;
 assign wire12659 = ( wire24  &  n_n509  &  n_n195 ) | ( wire24  &  n_n491  &  n_n195 ) ;
 assign wire12663 = ( n_n5010 ) | ( n_n4966 ) | ( wire12659 ) ;
 assign wire12664 = ( n_n5011 ) | ( n_n4961 ) | ( wire706 ) | ( wire12658 ) ;
 assign wire12669 = ( n_n5027 ) | ( n_n5048 ) | ( wire695 ) ;
 assign wire12670 = ( n_n5042 ) | ( n_n5022 ) | ( n_n5067 ) | ( n_n5020 ) ;
 assign wire12672 = ( n_n5072 ) | ( n_n5075 ) | ( wire12669 ) | ( wire12670 ) ;
 assign wire12673 = ( wire12656 ) | ( wire12657 ) | ( wire12663 ) | ( wire12664 ) ;
 assign wire12675 = ( wire11  &  n_n491  &  n_n260 ) | ( wire23  &  n_n491  &  n_n260 ) ;
 assign wire12678 = ( n_n4885 ) | ( n_n4911 ) | ( wire12675 ) ;
 assign wire12679 = ( n_n4890 ) | ( n_n4886 ) | ( n_n4892 ) | ( wire324 ) ;
 assign wire12682 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4815 ) ;
 assign wire12683 = ( n_n4830 ) | ( n_n4800 ) | ( n_n4825 ) | ( wire693 ) ;
 assign wire12688 = ( n_n4918 ) | ( n_n4917 ) | ( n_n4954 ) ;
 assign wire12689 = ( n_n4928 ) | ( n_n4950 ) | ( n_n4936 ) | ( n_n4956 ) ;
 assign wire12691 = ( n_n4931 ) | ( n_n4948 ) | ( wire12688 ) | ( wire12689 ) ;
 assign wire12693 = ( n_n554 ) | ( wire12678 ) | ( wire12679 ) | ( wire12691 ) ;
 assign wire12694 = ( wire12649 ) | ( wire12650 ) | ( wire12672 ) | ( wire12673 ) ;
 assign wire12699 = ( n_n4371 ) | ( n_n4442 ) | ( n_n4417 ) ;
 assign wire12700 = ( n_n4441 ) | ( n_n4404 ) | ( n_n4437 ) | ( n_n4384 ) ;
 assign wire12706 = ( n_n4512 ) | ( n_n4453 ) | ( n_n4471 ) ;
 assign wire12707 = ( n_n4450 ) | ( n_n4460 ) | ( n_n4473 ) | ( n_n4506 ) ;
 assign wire12710 = ( wire24  &  n_n509  &  n_n536 ) | ( wire24  &  n_n536  &  n_n500 ) ;
 assign wire12713 = ( n_n4338 ) | ( n_n4327 ) | ( n_n4326 ) ;
 assign wire12714 = ( n_n4320 ) | ( n_n4315 ) | ( wire12710 ) ;
 assign wire12718 = ( wire42 ) | ( wire22  &  n_n473  &  n_n260 ) ;
 assign wire12722 = ( wire22  &  n_n491  &  n_n260 ) | ( wire15  &  n_n491  &  n_n260 ) ;
 assign wire12724 = ( n_n4898 ) | ( n_n4901 ) | ( n_n4904 ) | ( n_n4899 ) ;
 assign wire12725 = ( wire154 ) | ( n_n4896 ) | ( wire12722 ) ;
 assign wire12729 = ( n_n4869 ) | ( n_n4876 ) | ( wire330 ) ;
 assign wire12730 = ( wire295 ) | ( n_n4875 ) | ( n_n4871 ) | ( n_n4874 ) ;
 assign wire12732 = ( wire17  &  n_n509  &  n_n526 ) | ( wire17  &  n_n509  &  n_n530 ) ;
 assign wire12735 = ( n_n4857 ) | ( n_n4862 ) | ( wire12732 ) ;
 assign wire12736 = ( wire277 ) | ( n_n4861 ) | ( n_n4851 ) | ( n_n4863 ) ;
 assign wire12740 = ( wire22  &  n_n535  &  n_n260 ) | ( wire20  &  n_n535  &  n_n260 ) ;
 assign wire12742 = ( n_n4835 ) | ( n_n4832 ) | ( n_n4828 ) | ( n_n4839 ) ;
 assign wire12743 = ( n_n4838 ) | ( wire304 ) | ( wire12740 ) ;
 assign wire12744 = ( wire24  &  n_n518  &  n_n260 ) | ( wire15  &  n_n518  &  n_n260 ) ;
 assign wire12745 = ( wire17  &  n_n530  &  n_n518 ) | ( wire17  &  n_n534  &  n_n518 ) ;
 assign wire12747 = ( wire150 ) | ( wire52 ) ;
 assign wire12748 = ( n_n4827 ) | ( n_n4824 ) | ( wire12744 ) ;
 assign wire12749 = ( n_n4822 ) | ( n_n4826 ) | ( wire12745 ) ;
 assign wire12752 = ( n_n834 ) | ( wire85 ) | ( wire12225 ) | ( wire12749 ) ;
 assign wire12753 = ( wire12742 ) | ( wire12743 ) | ( wire12747 ) | ( wire12748 ) ;
 assign wire12756 = ( n_n4803 ) | ( n_n4804 ) | ( wire686 ) ;
 assign wire12757 = ( n_n4811 ) | ( n_n4801 ) | ( n_n4802 ) | ( n_n4807 ) ;
 assign wire12759 = ( wire24  &  n_n482  &  n_n325 ) | ( wire25  &  n_n482  &  n_n325 ) ;
 assign wire12760 = ( wire14  &  n_n522  &  n_n482 ) | ( wire14  &  n_n482  &  n_n532 ) ;
 assign wire12762 = ( n_n4782 ) | ( n_n4781 ) | ( wire12759 ) ;
 assign wire12763 = ( n_n4784 ) | ( n_n4783 ) | ( n_n4780 ) | ( wire12760 ) ;
 assign wire12766 = ( n_n4789 ) | ( n_n4793 ) | ( n_n4797 ) | ( wire179 ) ;
 assign wire12767 = ( wire292 ) | ( wire380 ) | ( wire12766 ) ;
 assign wire12769 = ( n_n4887 ) | ( wire17  &  n_n526  &  n_n500 ) ;
 assign wire12770 = ( n_n4891 ) | ( n_n4884 ) | ( n_n4883 ) ;
 assign wire12771 = ( n_n4882 ) | ( n_n4881 ) | ( wire261 ) ;
 assign wire12774 = ( wire12729 ) | ( wire12730 ) | ( wire12735 ) | ( wire12736 ) ;
 assign wire12775 = ( wire12769 ) | ( wire12770 ) | ( wire12771 ) | ( wire12774 ) ;
 assign wire12778 = ( wire21  &  n_n509  &  n_n325 ) | ( wire20  &  n_n509  &  n_n325 ) ;
 assign wire12783 = ( n_n4705 ) | ( n_n4706 ) | ( n_n4713 ) ;
 assign wire12784 = ( n_n4711 ) | ( n_n4712 ) | ( n_n4710 ) | ( n_n4709 ) ;
 assign wire12787 = ( wire11  &  n_n325  &  n_n518 ) | ( wire15  &  n_n325  &  n_n518 ) ;
 assign wire12788 = ( wire21  &  n_n325  &  n_n518 ) | ( wire24  &  n_n325  &  n_n518 ) ;
 assign wire12790 = ( n_n4720 ) | ( n_n4728 ) | ( wire12787 ) ;
 assign wire12791 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4721 ) | ( wire12788 ) ;
 assign wire12792 = ( wire24  &  n_n535  &  n_n325 ) | ( wire25  &  n_n535  &  n_n325 ) ;
 assign wire12794 = ( n_n4695 ) | ( n_n4696 ) | ( wire12792 ) ;
 assign wire12796 = ( n_n3849 ) | ( n_n4702 ) | ( n_n4694 ) | ( wire12794 ) ;
 assign wire12799 = ( n_n4683 ) | ( n_n4684 ) | ( wire417 ) ;
 assign wire12800 = ( n_n4677 ) | ( wire81 ) | ( wire418 ) | ( n_n4685 ) ;
 assign wire12801 = ( i_9_  &  n_n473  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n532 ) ;
 assign wire12802 = ( wire21  &  n_n473  &  n_n390 ) | ( wire15  &  n_n473  &  n_n390 ) ;
 assign wire12804 = ( wire12801 ) | ( wire225 ) ;
 assign wire12805 = ( n_n4673 ) | ( n_n4674 ) | ( n_n4671 ) | ( wire12802 ) ;
 assign wire12810 = ( n_n4644 ) | ( n_n4649 ) | ( n_n4657 ) ;
 assign wire12811 = ( n_n4662 ) | ( n_n4659 ) | ( n_n4655 ) | ( n_n4658 ) ;
 assign wire12813 = ( n_n4663 ) | ( n_n4652 ) | ( wire12810 ) | ( wire12811 ) ;
 assign wire12814 = ( wire12799 ) | ( wire12800 ) | ( wire12804 ) | ( wire12805 ) ;
 assign wire12815 = ( wire21  &  n_n500  &  n_n325 ) | ( wire20  &  n_n500  &  n_n325 ) ;
 assign wire12819 = ( n_n4758 ) | ( n_n4747 ) | ( wire12815 ) ;
 assign wire12820 = ( n_n4752 ) | ( wire47 ) | ( n_n4751 ) | ( n_n4745 ) ;
 assign wire12822 = ( n_n4760 ) | ( n_n4769 ) | ( n_n4762 ) ;
 assign wire12826 = ( n_n856 ) | ( wire12819 ) | ( wire12820 ) | ( wire12822 ) ;
 assign wire12827 = ( n_n4205 ) | ( n_n4204 ) | ( wire456 ) | ( wire12826 ) ;
 assign wire12831 = ( wire11  &  n_n535  &  n_n195 ) | ( wire15  &  n_n535  &  n_n195 ) ;
 assign wire12832 = ( wire24  &  n_n535  &  n_n195 ) | ( wire25  &  n_n535  &  n_n195 ) ;
 assign wire12833 = ( n_n4952 ) | ( n_n4949 ) | ( wire12831 ) ;
 assign wire12834 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4947 ) | ( wire12832 ) ;
 assign wire12835 = ( wire18  &  n_n522  &  n_n535 ) | ( wire18  &  n_n526  &  n_n535 ) ;
 assign wire12838 = ( n_n4940 ) | ( n_n4939 ) | ( wire342 ) ;
 assign wire12839 = ( wire362 ) | ( wire341 ) ;
 assign wire12841 = ( wire59 ) | ( wire180 ) | ( n_n4971 ) | ( wire12166 ) ;
 assign wire12843 = ( n_n4938 ) | ( n_n4933 ) | ( wire12835 ) | ( wire12841 ) ;
 assign wire12844 = ( wire12833 ) | ( wire12834 ) | ( wire12838 ) | ( wire12839 ) ;
 assign wire12845 = ( wire21  &  n_n509  &  n_n195 ) | ( wire11  &  n_n509  &  n_n195 ) ;
 assign wire12848 = ( n_n4983 ) | ( n_n4984 ) | ( wire12845 ) ;
 assign wire12849 = ( n_n4993 ) | ( wire134 ) | ( n_n4994 ) | ( n_n4986 ) ;
 assign wire12852 = ( wire252 ) | ( wire103 ) ;
 assign wire12853 = ( n_n4998 ) | ( wire57 ) | ( wire743 ) ;
 assign wire12854 = ( n_n4975 ) | ( n_n4999 ) | ( n_n4981 ) | ( n_n5002 ) ;
 assign wire12857 = ( n_n4973 ) | ( n_n801 ) | ( wire11809 ) | ( wire12854 ) ;
 assign wire12858 = ( wire12848 ) | ( wire12849 ) | ( wire12852 ) | ( wire12853 ) ;
 assign wire12859 = ( wire17  &  n_n522  &  n_n482 ) | ( wire17  &  n_n530  &  n_n482 ) ;
 assign wire12862 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4915 ) | ( wire12859 ) ;
 assign wire12863 = ( n_n4920 ) | ( n_n4919 ) | ( wire340 ) | ( wire12862 ) ;
 assign wire12865 = ( n_n691 ) | ( wire12724 ) | ( wire12725 ) | ( wire12863 ) ;
 assign wire12866 = ( wire12843 ) | ( wire12844 ) | ( wire12857 ) | ( wire12858 ) ;
 assign wire12871 = ( n_n5241 ) | ( n_n5234 ) | ( n_n5242 ) ;
 assign wire12872 = ( n_n5240 ) | ( n_n5238 ) | ( wire318 ) ;
 assign wire12874 = ( i_9_  &  n_n535  &  n_n520  &  n_n65 ) | ( (~ i_9_)  &  n_n535  &  n_n520  &  n_n65 ) ;
 assign wire12875 = ( n_n5229 ) | ( wire19  &  n_n522  &  n_n535 ) ;
 assign wire12876 = ( wire182 ) | ( wire19  &  n_n532  &  n_n518 ) ;
 assign wire12877 = ( n_n5228 ) | ( n_n5225 ) | ( wire183 ) ;
 assign wire12881 = ( n_n2291 ) | ( n_n763 ) | ( n_n761 ) | ( wire12875 ) ;
 assign wire12883 = ( i_9_  &  n_n526  &  n_n500  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n130 ) ;
 assign wire12884 = ( i_9_  &  n_n524  &  n_n500  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n500  &  n_n130 ) ;
 assign wire12888 = ( n_n5167 ) | ( n_n5162 ) | ( wire168 ) ;
 assign wire12889 = ( n_n5163 ) | ( n_n5159 ) | ( wire287 ) | ( n_n5169 ) ;
 assign wire12892 = ( n_n5142 ) | ( n_n5144 ) | ( wire679 ) ;
 assign wire12893 = ( n_n5150 ) | ( n_n5149 ) | ( wire407 ) ;
 assign wire12894 = ( n_n5133 ) | ( n_n5153 ) | ( n_n5148 ) | ( wire12883 ) ;
 assign wire12898 = ( wire12888 ) | ( wire12889 ) | ( wire12892 ) | ( wire12893 ) ;
 assign wire12902 = ( n_n5059 ) | ( n_n5073 ) | ( wire160 ) ;
 assign wire12904 = ( i_9_  &  n_n473  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n195 ) ;
 assign wire12907 = ( n_n5050 ) | ( n_n5049 ) | ( wire12904 ) ;
 assign wire12908 = ( n_n5057 ) | ( wire166 ) | ( n_n5047 ) | ( n_n5051 ) ;
 assign wire12909 = ( wire25  &  n_n535  &  n_n130 ) | ( wire15  &  n_n535  &  n_n130 ) ;
 assign wire12914 = ( n_n5079 ) | ( n_n5083 ) | ( n_n5080 ) | ( wire209 ) ;
 assign wire12915 = ( n_n5074 ) | ( n_n5082 ) | ( wire12909 ) | ( wire12914 ) ;
 assign wire12917 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire12921 = ( n_n5129 ) | ( n_n5120 ) | ( wire336 ) ;
 assign wire12922 = ( n_n5127 ) | ( n_n5128 ) | ( wire414 ) | ( n_n5122 ) ;
 assign wire12924 = ( wire12  &  n_n524  &  n_n518 ) | ( wire12  &  n_n528  &  n_n518 ) ;
 assign wire12925 = ( n_n5107 ) | ( wire122 ) | ( n_n5108 ) ;
 assign wire12926 = ( n_n5112 ) | ( n_n5086 ) | ( n_n5087 ) | ( n_n5088 ) ;
 assign wire12929 = ( wire28 ) | ( wire88 ) | ( wire12917 ) | ( wire12924 ) ;
 assign wire12930 = ( wire12921 ) | ( wire12922 ) | ( wire12925 ) | ( wire12926 ) ;
 assign wire12931 = ( wire18  &  n_n522  &  n_n500 ) | ( wire18  &  n_n500  &  n_n520 ) ;
 assign wire12933 = ( wire394 ) | ( wire297 ) ;
 assign wire12934 = ( n_n5016 ) | ( n_n5013 ) | ( n_n5007 ) | ( wire12931 ) ;
 assign wire12935 = ( wire18  &  n_n522  &  n_n491 ) | ( wire18  &  n_n524  &  n_n491 ) ;
 assign wire12936 = ( wire11  &  n_n491  &  n_n195 ) | ( wire23  &  n_n491  &  n_n195 ) ;
 assign wire12938 = ( wire12935 ) | ( wire265 ) ;
 assign wire12939 = ( n_n5029 ) | ( wire253 ) | ( wire12936 ) ;
 assign wire12940 = ( wire18  &  n_n526  &  n_n482 ) | ( wire18  &  n_n530  &  n_n482 ) ;
 assign wire12941 = ( wire22  &  n_n482  &  n_n195 ) | ( wire15  &  n_n482  &  n_n195 ) ;
 assign wire12943 = ( n_n5043 ) | ( n_n5044 ) | ( wire12940 ) ;
 assign wire12944 = ( wire231 ) | ( n_n5039 ) | ( wire12941 ) ;
 assign wire12946 = ( wire12933 ) | ( wire12934 ) | ( wire12938 ) | ( wire12939 ) ;
 assign wire12947 = ( wire12943 ) | ( wire12944 ) | ( wire12946 ) ;
 assign wire12949 = ( wire20  &  n_n491  &  n_n65 ) | ( wire25  &  n_n491  &  n_n65 ) ;
 assign wire12952 = ( n_n5277 ) | ( n_n5283 ) | ( n_n5280 ) | ( wire12371 ) ;
 assign wire12953 = ( wire21  &  n_n509  &  n_n65 ) | ( wire21  &  n_n500  &  n_n65 ) ;
 assign wire12954 = ( wire19  &  n_n509  &  n_n522 ) | ( wire19  &  n_n509  &  n_n520 ) ;
 assign wire12958 = ( n_n5260 ) | ( n_n5253 ) | ( wire12954 ) ;
 assign wire12960 = ( wire77 ) | ( wire446 ) | ( wire205 ) | ( wire12953 ) ;
 assign wire12961 = ( n_n5255 ) | ( wire433 ) | ( n_n1521 ) | ( wire12958 ) ;
 assign wire12962 = ( wire333 ) | ( wire12949 ) | ( wire12952 ) | ( wire12960 ) ;
 assign wire12963 = ( wire20  &  n_n464  &  n_n65 ) | ( wire23  &  n_n464  &  n_n65 ) ;
 assign wire12966 = ( n_n5327 ) | ( n_n5328 ) | ( wire149 ) | ( wire12963 ) ;
 assign wire12967 = ( wire148 ) | ( n_n5322 ) | ( wire175 ) | ( wire11946 ) ;
 assign wire12969 = ( n_n5303 ) | ( wire63 ) | ( n_n5304 ) ;
 assign wire12970 = ( n_n5307 ) | ( n_n5309 ) | ( n_n5308 ) ;
 assign wire12971 = ( wire19  &  n_n522  &  n_n473 ) | ( wire19  &  n_n473  &  n_n526 ) ;
 assign wire12972 = ( wire22  &  n_n473  &  n_n65 ) | ( wire23  &  n_n473  &  n_n65 ) ;
 assign wire12975 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5315 ) | ( wire12972 ) ;
 assign wire12976 = ( wire21  &  n_n482  &  n_n65 ) | ( wire11  &  n_n482  &  n_n65 ) ;
 assign wire12978 = ( n_n5291 ) | ( n_n5292 ) | ( n_n5298 ) ;
 assign wire12979 = ( n_n5288 ) | ( n_n5286 ) | ( wire12976 ) ;
 assign wire12981 = ( n_n5290 ) | ( n_n5289 ) | ( wire12978 ) | ( wire12979 ) ;
 assign wire12984 = ( n_n632 ) | ( n_n662 ) | ( n_n661 ) | ( wire12981 ) ;
 assign wire12985 = ( wire11  &  n_n464  &  n_n130 ) | ( wire23  &  n_n464  &  n_n130 ) ;
 assign wire12986 = ( wire21  &  n_n464  &  n_n130 ) | ( wire15  &  n_n464  &  n_n130 ) ;
 assign wire12988 = ( wire12985 ) | ( wire452 ) ;
 assign wire12989 = ( n_n5201 ) | ( n_n5205 ) | ( wire761 ) | ( wire12986 ) ;
 assign wire12991 = ( wire112 ) | ( n_n5189 ) | ( n_n5190 ) ;
 assign wire12992 = ( n_n5188 ) | ( n_n5194 ) | ( wire453 ) | ( n_n5192 ) ;
 assign wire12995 = ( n_n5181 ) | ( n_n5184 ) | ( wire107 ) ;
 assign wire12996 = ( n_n5177 ) | ( n_n5172 ) | ( wire44 ) | ( n_n5176 ) ;
 assign wire12998 = ( wire12988 ) | ( wire12989 ) | ( wire12991 ) | ( wire12992 ) ;
 assign wire12999 = ( wire12995 ) | ( wire12996 ) | ( wire12998 ) ;
 assign wire13001 = ( wire12961 ) | ( wire12962 ) | ( wire12984 ) | ( wire12999 ) ;
 assign wire13003 = ( wire13  &  n_n522  &  n_n535 ) | ( wire13  &  n_n526  &  n_n535 ) ;
 assign wire13005 = ( n_n4445 ) | ( n_n4446 ) | ( wire128 ) ;
 assign wire13006 = ( wire368 ) | ( n_n4447 ) | ( wire13003 ) ;
 assign wire13008 = ( wire16  &  n_n464  &  n_n528 ) | ( wire16  &  n_n464  &  n_n532 ) ;
 assign wire13013 = ( n_n4436 ) | ( n_n4443 ) | ( n_n4428 ) | ( n_n4427 ) ;
 assign wire13015 = ( wire233 ) | ( wire234 ) | ( wire37 ) | ( wire13008 ) ;
 assign wire13016 = ( n_n4421 ) | ( wire215 ) | ( n_n910 ) | ( wire13013 ) ;
 assign wire13017 = ( wire13005 ) | ( wire13006 ) | ( wire13015 ) ;
 assign wire13020 = ( n_n4470 ) | ( n_n4472 ) | ( n_n4476 ) ;
 assign wire13022 = ( wire24  &  n_n455  &  n_n500 ) | ( wire25  &  n_n455  &  n_n500 ) ;
 assign wire13025 = ( wire13022 ) | ( wire70 ) ;
 assign wire13026 = ( n_n4487 ) | ( wire66 ) | ( n_n4492 ) | ( n_n4486 ) ;
 assign wire13027 = ( i_9_  &  n_n526  &  n_n455  &  n_n500 ) | ( (~ i_9_)  &  n_n526  &  n_n455  &  n_n500 ) ;
 assign wire13028 = ( wire24  &  n_n455  &  n_n491 ) | ( wire15  &  n_n455  &  n_n491 ) ;
 assign wire13029 = ( wire308 ) | ( wire22  &  n_n455  &  n_n491 ) ;
 assign wire13034 = ( n_n4502 ) | ( n_n4501 ) | ( wire378 ) ;
 assign wire13035 = ( n_n4521 ) | ( n_n4504 ) | ( n_n4524 ) | ( n_n4503 ) ;
 assign wire13036 = ( n_n4522 ) | ( n_n4525 ) | ( n_n4505 ) | ( n_n4499 ) ;
 assign wire13039 = ( n_n4498 ) | ( n_n3879 ) | ( wire13027 ) | ( wire13036 ) ;
 assign wire13042 = ( n_n4467 ) | ( n_n4463 ) | ( n_n4466 ) | ( n_n4468 ) ;
 assign wire13044 = ( n_n4469 ) | ( n_n4462 ) | ( n_n2058 ) | ( wire13042 ) ;
 assign wire13046 = ( n_n725 ) | ( wire13025 ) | ( wire13026 ) | ( wire13044 ) ;
 assign wire13048 = ( wire16  &  n_n524  &  n_n535 ) | ( wire16  &  n_n535  &  n_n528 ) ;
 assign wire13049 = ( wire364 ) | ( wire171 ) ;
 assign wire13050 = ( n_n4313 ) | ( wire11583 ) | ( wire13048 ) ;
 assign wire13053 = ( n_n4325 ) | ( n_n4329 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire13054 = ( n_n4335 ) | ( n_n4323 ) | ( n_n4330 ) | ( wire12570 ) ;
 assign wire13055 = ( wire16  &  n_n528  &  n_n500 ) | ( wire16  &  n_n500  &  n_n530 ) ;
 assign wire13056 = ( n_n4369 ) | ( n_n4367 ) | ( n_n4368 ) ;
 assign wire13057 = ( wire15  &  n_n509  &  n_n536 ) | ( wire23  &  n_n509  &  n_n536 ) ;
 assign wire13059 = ( n_n4352 ) | ( n_n4351 ) | ( n_n4356 ) | ( n_n4355 ) ;
 assign wire13060 = ( n_n4357 ) | ( n_n4358 ) | ( n_n4354 ) | ( wire13057 ) ;
 assign wire13062 = ( n_n4373 ) | ( n_n4374 ) | ( wire345 ) ;
 assign wire13063 = ( n_n4361 ) | ( wire423 ) | ( n_n4370 ) | ( n_n4378 ) ;
 assign wire13065 = ( n_n4365 ) | ( wire13055 ) | ( wire13056 ) | ( wire13063 ) ;
 assign wire13066 = ( wire27 ) | ( wire13059 ) | ( wire13060 ) | ( wire13062 ) ;
 assign wire13067 = ( wire16  &  n_n522  &  n_n473 ) | ( wire16  &  n_n473  &  n_n532 ) ;
 assign wire13069 = ( wire79 ) | ( wire328 ) ;
 assign wire13070 = ( n_n4416 ) | ( n_n4415 ) | ( n_n4414 ) | ( wire13067 ) ;
 assign wire13073 = ( n_n4389 ) | ( n_n4390 ) | ( n_n4394 ) ;
 assign wire13074 = ( n_n4383 ) | ( n_n4388 ) | ( n_n4396 ) | ( n_n4395 ) ;
 assign wire13077 = ( n_n4401 ) | ( n_n4405 ) | ( n_n4402 ) ;
 assign wire13078 = ( n_n4397 ) | ( n_n4398 ) | ( n_n4406 ) | ( n_n4408 ) ;
 assign wire13080 = ( n_n4400 ) | ( n_n4407 ) | ( wire13077 ) | ( wire13078 ) ;
 assign wire13084 = ( n_n4345 ) | ( wire124 ) | ( wire675 ) ;
 assign wire13085 = ( n_n4339 ) | ( n_n4344 ) | ( n_n4348 ) | ( wire156 ) ;
 assign wire13087 = ( wire13049 ) | ( wire13050 ) | ( wire13053 ) | ( wire13054 ) ;
 assign wire13088 = ( wire13084 ) | ( wire13085 ) | ( wire13087 ) ;
 assign wire13090 = ( wire13  &  n_n473  &  n_n530 ) | ( wire13  &  n_n473  &  n_n532 ) ;
 assign wire13091 = ( i_9_  &  n_n473  &  n_n524  &  n_n455 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n455 ) ;
 assign wire13093 = ( wire13  &  n_n473  &  n_n528 ) | ( wire13  &  n_n473  &  n_n520 ) ;
 assign wire13095 = ( n_n4544 ) | ( n_n4541 ) | ( wire13093 ) ;
 assign wire13096 = ( n_n4545 ) | ( n_n4551 ) | ( n_n4548 ) | ( wire13091 ) ;
 assign wire13100 = ( n_n4595 ) | ( n_n4596 ) | ( n_n4599 ) ;
 assign wire13101 = ( n_n4598 ) | ( n_n4593 ) | ( n_n4594 ) | ( n_n4600 ) ;
 assign wire13104 = ( wire10  &  n_n522  &  n_n535 ) | ( wire10  &  n_n535  &  n_n528 ) ;
 assign wire13105 = ( n_n4570 ) | ( n_n4569 ) | ( wire91 ) ;
 assign wire13106 = ( n_n4584 ) | ( n_n4583 ) | ( wire238 ) ;
 assign wire13107 = ( n_n4568 ) | ( wire99 ) | ( wire783 ) ;
 assign wire13108 = ( n_n4571 ) | ( n_n4582 ) | ( wire13104 ) ;
 assign wire13111 = ( n_n881 ) | ( wire13105 ) | ( wire13108 ) ;
 assign wire13113 = ( n_n4612 ) | ( n_n4610 ) | ( n_n4609 ) ;
 assign wire13114 = ( n_n4613 ) | ( n_n4605 ) | ( wire465 ) | ( wire12519 ) ;
 assign wire13117 = ( n_n4639 ) | ( n_n4642 ) | ( n_n4632 ) ;
 assign wire13118 = ( n_n4637 ) | ( n_n4638 ) | ( wire190 ) ;
 assign wire13119 = ( n_n4616 ) | ( n_n4629 ) | ( n_n4630 ) | ( n_n4619 ) ;
 assign wire13120 = ( n_n4617 ) | ( n_n4634 ) | ( n_n4628 ) | ( n_n4640 ) ;
 assign wire13123 = ( n_n3861 ) | ( wire13117 ) | ( wire13120 ) ;
 assign wire13124 = ( wire13113 ) | ( wire13114 ) | ( wire13118 ) | ( wire13119 ) ;
 assign wire13126 = ( wire13  &  n_n464  &  n_n528 ) | ( wire13  &  n_n464  &  n_n530 ) ;
 assign wire13127 = ( n_n4561 ) | ( n_n4532 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire13128 = ( n_n4536 ) | ( wire13090 ) | ( wire13126 ) ;
 assign wire13132 = ( n_n3875 ) | ( wire13095 ) | ( wire13096 ) | ( wire13127 ) ;
 assign wire13133 = ( n_n3870 ) | ( wire82 ) | ( wire13128 ) | ( wire13132 ) ;
 assign wire13136 = ( n_n630 ) | ( n_n631 ) | ( n_n629 ) ;
 assign wire13140 = ( n_n5305 ) | ( n_n5293 ) | ( n_n5297 ) ;
 assign wire13141 = ( n_n5296 ) | ( n_n5284 ) | ( wire13140 ) ;
 assign wire13144 = ( n_n562 ) | ( n_n561 ) | ( n_n563 ) | ( wire13141 ) ;
 assign wire13146 = ( n_n543 ) | ( wire12629 ) | ( wire12630 ) | ( wire13144 ) ;
 assign wire13147 = ( wire12693 ) | ( wire12694 ) | ( wire13146 ) ;
 assign wire13149 = ( n_n4767 ) | ( n_n4764 ) | ( n_n4766 ) ;
 assign wire13151 = ( i_9_  &  n_n473  &  n_n530  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n530  &  n_n325 ) ;
 assign wire13153 = ( n_n4790 ) | ( n_n4798 ) | ( wire158 ) ;
 assign wire13154 = ( wire179 ) | ( n_n4799 ) | ( wire13151 ) ;
 assign wire13156 = ( n_n4821 ) | ( n_n4822 ) | ( n_n4823 ) ;
 assign wire13162 = ( n_n4816 ) | ( n_n4806 ) | ( n_n4805 ) | ( n_n4815 ) ;
 assign wire13163 = ( n_n4817 ) | ( n_n4800 ) | ( n_n4803 ) | ( n_n4804 ) ;
 assign wire13166 = ( n_n4801 ) | ( n_n4818 ) | ( n_n4197 ) | ( wire390 ) ;
 assign wire13170 = ( wire245 ) | ( wire102 ) ;
 assign wire13171 = ( n_n4857 ) | ( n_n4862 ) | ( n_n4856 ) | ( wire40 ) ;
 assign wire13172 = ( wire21  &  n_n518  &  n_n260 ) | ( wire11  &  n_n518  &  n_n260 ) ;
 assign wire13173 = ( wire176 ) | ( wire277 ) ;
 assign wire13174 = ( n_n4849 ) | ( n_n4850 ) | ( n_n4848 ) | ( wire13172 ) ;
 assign wire13176 = ( n_n4843 ) | ( wire20  &  n_n535  &  n_n260 ) ;
 assign wire13177 = ( n_n4839 ) | ( n_n4840 ) | ( n_n4838 ) ;
 assign wire13178 = ( n_n4834 ) | ( n_n4835 ) | ( n_n4832 ) | ( n_n4833 ) ;
 assign wire13181 = ( wire13170 ) | ( wire13171 ) | ( wire13173 ) | ( wire13174 ) ;
 assign wire13182 = ( wire14  &  n_n526  &  n_n482 ) | ( wire14  &  n_n528  &  n_n482 ) ;
 assign wire13183 = ( wire24  &  n_n482  &  n_n325 ) | ( wire20  &  n_n482  &  n_n325 ) ;
 assign wire13185 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4775 ) | ( wire13183 ) ;
 assign wire13187 = ( wire447 ) | ( wire13149 ) | ( wire13153 ) | ( wire13154 ) ;
 assign wire13188 = ( wire131 ) | ( wire13182 ) | ( wire13185 ) | ( wire13187 ) ;
 assign wire13193 = ( n_n4885 ) | ( n_n4882 ) | ( wire330 ) ;
 assign wire13194 = ( wire260 ) | ( n_n4880 ) | ( n_n4889 ) | ( n_n4883 ) ;
 assign wire13198 = ( n_n4898 ) | ( n_n4895 ) | ( wire49 ) ;
 assign wire13199 = ( n_n4894 ) | ( wire96 ) | ( n_n4897 ) | ( n_n4891 ) ;
 assign wire13202 = ( n_n4911 ) | ( n_n4912 ) | ( n_n4915 ) ;
 assign wire13203 = ( n_n4909 ) | ( n_n4916 ) | ( wire154 ) ;
 assign wire13208 = ( n_n4943 ) | ( n_n4937 ) | ( n_n4938 ) | ( n_n4936 ) ;
 assign wire13209 = ( n_n4930 ) | ( n_n4939 ) | ( wire180 ) | ( n_n4944 ) ;
 assign wire13211 = ( wire42 ) | ( wire31 ) ;
 assign wire13213 = ( n_n4926 ) | ( n_n4925 ) | ( n_n1592 ) | ( wire13211 ) ;
 assign wire13215 = ( wire18  &  n_n522  &  n_n535 ) | ( wire18  &  n_n535  &  n_n520 ) ;
 assign wire13216 = ( i_9_  &  n_n535  &  n_n530  &  n_n195 ) | ( (~ i_9_)  &  n_n535  &  n_n530  &  n_n195 ) ;
 assign wire13217 = ( wire11  &  n_n518  &  n_n195 ) | ( wire24  &  n_n518  &  n_n195 ) ;
 assign wire13218 = ( i_9_  &  n_n530  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n530  &  n_n518  &  n_n195 ) ;
 assign wire13222 = ( n_n4959 ) | ( n_n4960 ) | ( wire771 ) | ( wire772 ) ;
 assign wire13223 = ( wire317 ) | ( wire141 ) ;
 assign wire13224 = ( n_n4967 ) | ( n_n4962 ) | ( n_n4948 ) | ( n_n4953 ) ;
 assign wire13225 = ( n_n4965 ) | ( n_n4955 ) | ( wire13215 ) | ( wire13216 ) ;
 assign wire13228 = ( wire228 ) | ( wire13217 ) | ( wire13218 ) | ( wire13225 ) ;
 assign wire13229 = ( n_n814 ) | ( wire13222 ) | ( wire13223 ) | ( wire13224 ) ;
 assign wire13231 = ( wire174 ) | ( wire295 ) ;
 assign wire13233 = ( n_n4869 ) | ( n_n4876 ) | ( wire461 ) | ( wire13231 ) ;
 assign wire13234 = ( wire13193 ) | ( wire13194 ) | ( wire13198 ) | ( wire13199 ) ;
 assign wire13236 = ( n_n4058 ) | ( n_n4056 ) | ( wire13213 ) | ( wire13234 ) ;
 assign wire13237 = ( i_9_  &  n_n509  &  n_n528  &  n_n325 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n325 ) ;
 assign wire13239 = ( n_n4737 ) | ( n_n4738 ) | ( n_n4732 ) | ( wire767 ) ;
 assign wire13240 = ( wire374 ) | ( n_n4743 ) | ( wire13237 ) ;
 assign wire13244 = ( n_n4697 ) | ( n_n4695 ) | ( wire221 ) ;
 assign wire13246 = ( i_9_  &  n_n520  &  n_n325  &  n_n518 ) | ( (~ i_9_)  &  n_n520  &  n_n325  &  n_n518 ) ;
 assign wire13248 = ( wire21  &  n_n325  &  n_n518 ) | ( wire25  &  n_n325  &  n_n518 ) ;
 assign wire13249 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4705 ) | ( n_n4706 ) ;
 assign wire13250 = ( n_n4722 ) | ( wire173 ) | ( n_n4721 ) ;
 assign wire13251 = ( n_n4708 ) | ( n_n4716 ) | ( wire13248 ) ;
 assign wire13254 = ( n_n4216 ) | ( n_n4728 ) | ( wire13246 ) | ( wire13251 ) ;
 assign wire13256 = ( i_9_  &  n_n473  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n532 ) ;
 assign wire13259 = ( n_n4658 ) | ( wire775 ) | ( wire13256 ) ;
 assign wire13260 = ( n_n4664 ) | ( n_n4662 ) | ( wire72 ) | ( n_n4657 ) ;
 assign wire13261 = ( i_9_  &  n_n473  &  n_n528  &  n_n390 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n390 ) ;
 assign wire13263 = ( n_n4673 ) | ( n_n4674 ) | ( wire157 ) ;
 assign wire13264 = ( wire80 ) | ( n_n4680 ) | ( wire13261 ) ;
 assign wire13265 = ( wire10  &  n_n524  &  n_n464 ) | ( wire10  &  n_n464  &  n_n526 ) ;
 assign wire13266 = ( wire11  &  n_n464  &  n_n390 ) | ( wire15  &  n_n464  &  n_n390 ) ;
 assign wire13268 = ( n_n4683 ) | ( wire81 ) | ( n_n4684 ) | ( wire13266 ) ;
 assign wire13269 = ( wire445 ) | ( wire13265 ) | ( wire13268 ) ;
 assign wire13270 = ( wire13259 ) | ( wire13260 ) | ( wire13263 ) | ( wire13264 ) ;
 assign wire13272 = ( wire22  &  n_n500  &  n_n325 ) | ( wire24  &  n_n500  &  n_n325 ) ;
 assign wire13274 = ( n_n4754 ) | ( n_n4749 ) | ( wire47 ) ;
 assign wire13275 = ( wire109 ) | ( n_n4752 ) | ( wire13272 ) ;
 assign wire13277 = ( wire11836 ) | ( wire11837 ) | ( wire13239 ) | ( wire13240 ) ;
 assign wire13278 = ( wire13274 ) | ( wire13275 ) | ( wire13277 ) ;
 assign wire13283 = ( n_n5142 ) | ( n_n5135 ) | ( wire407 ) ;
 assign wire13284 = ( n_n5150 ) | ( wire76 ) | ( n_n5140 ) | ( n_n5143 ) ;
 assign wire13285 = ( wire20  &  n_n491  &  n_n130 ) | ( wire23  &  n_n491  &  n_n130 ) ;
 assign wire13287 = ( wire168 ) | ( wire358 ) ;
 assign wire13288 = ( wire196 ) | ( n_n5151 ) | ( wire13285 ) ;
 assign wire13291 = ( wire12  &  n_n473  &  n_n532 ) | ( wire12  &  n_n473  &  n_n534 ) ;
 assign wire13292 = ( n_n5174 ) | ( n_n5183 ) | ( wire113 ) ;
 assign wire13293 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) | ( wire13291 ) ;
 assign wire13294 = ( wire12  &  n_n526  &  n_n482 ) | ( wire12  &  n_n482  &  n_n532 ) ;
 assign wire13296 = ( wire332 ) | ( wire254 ) ;
 assign wire13297 = ( n_n5169 ) | ( wire33 ) | ( wire13294 ) ;
 assign wire13298 = ( i_9_  &  n_n522  &  n_n473  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n473  &  n_n130 ) ;
 assign wire13301 = ( n_n5187 ) | ( n_n5196 ) | ( wire13298 ) ;
 assign wire13303 = ( n_n5195 ) | ( n_n2670 ) | ( n_n5192 ) | ( wire13301 ) ;
 assign wire13304 = ( wire13292 ) | ( wire13293 ) | ( wire13296 ) | ( wire13297 ) ;
 assign wire13305 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire13306 = ( i_9_  &  n_n526  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n535  &  n_n130 ) ;
 assign wire13308 = ( n_n5109 ) | ( n_n5107 ) | ( n_n5113 ) | ( n_n5108 ) ;
 assign wire13310 = ( wire12  &  n_n530  &  n_n518 ) | ( wire12  &  n_n532  &  n_n518 ) ;
 assign wire13311 = ( i_9_  &  n_n535  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n535  &  n_n528  &  n_n130 ) ;
 assign wire13313 = ( wire279 ) | ( wire289 ) ;
 assign wire13314 = ( n_n5099 ) | ( n_n5085 ) | ( wire13310 ) ;
 assign wire13317 = ( n_n5106 ) | ( n_n5095 ) | ( wire144 ) | ( wire13311 ) ;
 assign wire13318 = ( wire28 ) | ( wire13308 ) | ( wire13313 ) | ( wire13314 ) ;
 assign wire13320 = ( wire12  &  n_n509  &  n_n528 ) | ( wire12  &  n_n528  &  n_n500 ) ;
 assign wire13322 = ( n_n5130 ) | ( n_n5127 ) | ( wire336 ) ;
 assign wire13323 = ( n_n5121 ) | ( n_n5122 ) | ( n_n5125 ) | ( wire13320 ) ;
 assign wire13325 = ( wire13283 ) | ( wire13284 ) | ( wire13287 ) | ( wire13288 ) ;
 assign wire13327 = ( wire13303 ) | ( wire13304 ) | ( wire13317 ) | ( wire13318 ) ;
 assign wire13329 = ( n_n5305 ) | ( n_n5306 ) | ( wire63 ) ;
 assign wire13333 = ( n_n5279 ) | ( wire333 ) | ( n_n5280 ) ;
 assign wire13334 = ( n_n5276 ) | ( n_n5281 ) | ( n_n5277 ) | ( wire218 ) ;
 assign wire13337 = ( n_n5262 ) | ( n_n5256 ) | ( n_n5259 ) ;
 assign wire13338 = ( n_n5258 ) | ( n_n5254 ) | ( wire434 ) ;
 assign wire13341 = ( n_n5241 ) | ( n_n5249 ) | ( n_n5242 ) ;
 assign wire13342 = ( n_n5244 ) | ( wire318 ) | ( n_n5243 ) ;
 assign wire13346 = ( wire205 ) | ( wire203 ) ;
 assign wire13347 = ( n_n5266 ) | ( n_n5271 ) | ( n_n5270 ) | ( wire77 ) ;
 assign wire13350 = ( wire19  &  n_n524  &  n_n535 ) | ( wire19  &  n_n535  &  n_n528 ) ;
 assign wire13351 = ( wire19  &  n_n528  &  n_n518 ) | ( wire19  &  n_n520  &  n_n518 ) ;
 assign wire13352 = ( wire21  &  n_n518  &  n_n65 ) | ( wire20  &  n_n518  &  n_n65 ) ;
 assign wire13354 = ( wire13351 ) | ( wire181 ) ;
 assign wire13355 = ( wire87 ) | ( wire182 ) | ( wire13352 ) ;
 assign wire13359 = ( n_n5210 ) | ( wire384 ) | ( n_n5209 ) ;
 assign wire13360 = ( n_n5204 ) | ( n_n5201 ) | ( n_n5207 ) | ( n_n5208 ) ;
 assign wire13361 = ( n_n5220 ) | ( n_n5203 ) | ( n_n5211 ) | ( n_n5205 ) ;
 assign wire13364 = ( n_n1530 ) | ( n_n5215 ) | ( wire13350 ) | ( wire13361 ) ;
 assign wire13365 = ( wire13354 ) | ( wire13355 ) | ( wire13359 ) | ( wire13360 ) ;
 assign wire13368 = ( i_9_  &  n_n482  &  n_n532  &  n_n65 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n65 ) ;
 assign wire13370 = ( n_n5294 ) | ( n_n5299 ) | ( n_n5287 ) | ( n_n5288 ) ;
 assign wire13372 = ( n_n5292 ) | ( wire441 ) | ( wire13368 ) | ( wire13370 ) ;
 assign wire13374 = ( n_n4026 ) | ( wire13333 ) | ( wire13334 ) | ( wire13372 ) ;
 assign wire13378 = ( wire18  &  n_n509  &  n_n528 ) | ( wire18  &  n_n509  &  n_n520 ) ;
 assign wire13380 = ( n_n4991 ) | ( n_n4996 ) | ( n_n4992 ) | ( n_n4995 ) ;
 assign wire13381 = ( n_n4999 ) | ( wire103 ) | ( wire13378 ) ;
 assign wire13384 = ( wire343 ) | ( wire393 ) ;
 assign wire13385 = ( n_n5004 ) | ( wire136 ) | ( n_n5013 ) | ( n_n5008 ) ;
 assign wire13390 = ( n_n5081 ) | ( n_n5082 ) | ( n_n5084 ) | ( n_n5079 ) ;
 assign wire13391 = ( wire21  &  n_n473  &  n_n195 ) | ( wire11  &  n_n473  &  n_n195 ) ;
 assign wire13392 = ( n_n5067 ) | ( n_n5057 ) | ( n_n5058 ) ;
 assign wire13393 = ( n_n5061 ) | ( wire160 ) | ( wire669 ) ;
 assign wire13394 = ( n_n5073 ) | ( n_n5074 ) | ( n_n5072 ) | ( wire13391 ) ;
 assign wire13397 = ( n_n1952 ) | ( n_n789 ) | ( wire13394 ) ;
 assign wire13398 = ( wire90 ) | ( wire13390 ) | ( wire13392 ) | ( wire13393 ) ;
 assign wire13399 = ( i_9_  &  n_n524  &  n_n491  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n491  &  n_n195 ) ;
 assign wire13400 = ( i_9_  &  n_n528  &  n_n491  &  n_n195 ) | ( (~ i_9_)  &  n_n528  &  n_n491  &  n_n195 ) ;
 assign wire13401 = ( wire18  &  n_n473  &  n_n528 ) | ( wire18  &  n_n473  &  n_n534 ) ;
 assign wire13404 = ( n_n5050 ) | ( n_n5049 ) | ( wire13401 ) ;
 assign wire13405 = ( n_n5045 ) | ( wire166 ) | ( n_n5051 ) | ( n_n5044 ) ;
 assign wire13406 = ( wire18  &  n_n526  &  n_n482 ) | ( wire18  &  n_n528  &  n_n482 ) ;
 assign wire13408 = ( i_9_  &  n_n524  &  n_n482  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n482  &  n_n195 ) ;
 assign wire13409 = ( n_n5034 ) | ( n_n5041 ) | ( wire13406 ) ;
 assign wire13410 = ( wire50 ) | ( n_n5029 ) | ( wire13408 ) ;
 assign wire13411 = ( i_9_  &  n_n491  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n491  &  n_n532  &  n_n195 ) ;
 assign wire13413 = ( n_n5025 ) | ( n_n5024 ) | ( wire13399 ) | ( wire13400 ) ;
 assign wire13414 = ( n_n5014 ) | ( wire13411 ) | ( wire13413 ) ;
 assign wire13415 = ( wire13404 ) | ( wire13405 ) | ( wire13409 ) | ( wire13410 ) ;
 assign wire13417 = ( i_9_  &  n_n509  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n534  &  n_n195 ) ;
 assign wire13419 = ( n_n4982 ) | ( n_n4981 ) | ( wire57 ) ;
 assign wire13421 = ( wire134 ) | ( n_n4980 ) | ( wire13417 ) | ( wire13419 ) ;
 assign wire13422 = ( wire13380 ) | ( wire13381 ) | ( wire13384 ) | ( wire13385 ) ;
 assign wire13424 = ( wire13397 ) | ( wire13398 ) | ( wire13414 ) | ( wire13415 ) ;
 assign wire13425 = ( i_9_  &  n_n522  &  n_n455  &  n_n535 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n535 ) ;
 assign wire13428 = ( wire236 ) | ( wire233 ) ;
 assign wire13429 = ( n_n4440 ) | ( n_n4434 ) | ( n_n4432 ) | ( wire98 ) ;
 assign wire13430 = ( wire22  &  n_n455  &  n_n535 ) | ( wire25  &  n_n455  &  n_n535 ) ;
 assign wire13431 = ( n_n4448 ) | ( n_n4447 ) | ( wire421 ) ;
 assign wire13432 = ( n_n4445 ) | ( n_n4444 ) | ( n_n4446 ) | ( wire13430 ) ;
 assign wire13436 = ( n_n4430 ) | ( n_n4425 ) | ( n_n4423 ) | ( n_n4429 ) ;
 assign wire13437 = ( n_n4421 ) | ( wire84 ) | ( n_n4424 ) | ( n_n4428 ) ;
 assign wire13438 = ( wire13437 ) | ( wire13436 ) ;
 assign wire13439 = ( wire13428 ) | ( wire13429 ) | ( wire13431 ) | ( wire13432 ) ;
 assign wire13441 = ( n_n4595 ) | ( n_n4591 ) | ( n_n4592 ) | ( n_n4596 ) ;
 assign wire13443 = ( wire10  &  n_n509  &  n_n524 ) | ( wire10  &  n_n509  &  n_n528 ) ;
 assign wire13445 = ( n_n4612 ) | ( wire45 ) | ( n_n4609 ) ;
 assign wire13446 = ( wire108 ) | ( n_n4600 ) | ( wire13443 ) ;
 assign wire13448 = ( wire22  &  n_n535  &  n_n390 ) | ( wire20  &  n_n535  &  n_n390 ) ;
 assign wire13450 = ( n_n4575 ) | ( n_n4584 ) | ( n_n4586 ) | ( n_n4583 ) ;
 assign wire13452 = ( n_n4573 ) | ( wire239 ) | ( wire13448 ) | ( wire13450 ) ;
 assign wire13454 = ( i_9_  &  n_n526  &  n_n491  &  n_n390 ) | ( (~ i_9_)  &  n_n526  &  n_n491  &  n_n390 ) ;
 assign wire13455 = ( i_9_  &  n_n390  &  n_n482  &  n_n534 ) | ( (~ i_9_)  &  n_n390  &  n_n482  &  n_n534 ) ;
 assign wire13457 = ( wire13455 ) | ( wire140 ) ;
 assign wire13458 = ( n_n4652 ) | ( n_n4643 ) | ( n_n4642 ) | ( wire13454 ) ;
 assign wire13459 = ( wire10  &  n_n528  &  n_n491 ) | ( wire10  &  n_n491  &  n_n532 ) ;
 assign wire13461 = ( wire22  &  n_n500  &  n_n390 ) | ( wire23  &  n_n500  &  n_n390 ) ;
 assign wire13462 = ( wire118 ) | ( n_n4633 ) | ( n_n4630 ) ;
 assign wire13463 = ( wire13459 ) | ( wire401 ) ;
 assign wire13465 = ( n_n4616 ) | ( wire465 ) | ( n_n4627 ) | ( wire12546 ) ;
 assign wire13467 = ( n_n4635 ) | ( n_n4620 ) | ( wire13461 ) | ( wire13465 ) ;
 assign wire13468 = ( wire13457 ) | ( wire13458 ) | ( wire13462 ) | ( wire13463 ) ;
 assign wire13470 = ( n_n4568 ) | ( wire455 ) | ( wire783 ) ;
 assign wire13471 = ( n_n4560 ) | ( n_n4569 ) | ( wire471 ) | ( wire91 ) ;
 assign wire13473 = ( wire13  &  n_n522  &  n_n473 ) | ( wire13  &  n_n473  &  n_n520 ) ;
 assign wire13474 = ( n_n4554 ) | ( n_n4541 ) | ( wire416 ) ;
 assign wire13475 = ( n_n4545 ) | ( wire13091 ) | ( wire13473 ) ;
 assign wire13478 = ( n_n4533 ) | ( n_n4536 ) | ( wire379 ) ;
 assign wire13479 = ( n_n4537 ) | ( n_n4527 ) | ( n_n4534 ) | ( wire11532 ) ;
 assign wire13481 = ( wire13470 ) | ( wire13471 ) | ( wire13474 ) | ( wire13475 ) ;
 assign wire13482 = ( wire13478 ) | ( wire13479 ) | ( wire13481 ) ;
 assign wire13487 = ( n_n4482 ) | ( n_n4489 ) | ( wire199 ) ;
 assign wire13488 = ( n_n4487 ) | ( n_n4478 ) | ( wire70 ) | ( n_n4486 ) ;
 assign wire13493 = ( n_n4491 ) | ( n_n4497 ) | ( n_n4500 ) | ( n_n4492 ) ;
 assign wire13494 = ( wire66 ) | ( n_n4496 ) | ( n_n4499 ) | ( n_n4493 ) ;
 assign wire13495 = ( n_n4512 ) | ( wire23  &  n_n455  &  n_n500 ) ;
 assign wire13496 = ( n_n4506 ) | ( n_n4508 ) | ( n_n4505 ) ;
 assign wire13497 = ( n_n4502 ) | ( wire308 ) | ( n_n4501 ) ;
 assign wire13501 = ( n_n4247 ) | ( n_n4246 ) | ( n_n3152 ) | ( wire13495 ) ;
 assign wire13502 = ( wire13493 ) | ( wire13494 ) | ( wire13496 ) | ( wire13497 ) ;
 assign wire13503 = ( wire21  &  n_n455  &  n_n518 ) | ( wire23  &  n_n455  &  n_n518 ) ;
 assign wire13504 = ( i_9_  &  n_n522  &  n_n455  &  n_n518 ) | ( (~ i_9_)  &  n_n522  &  n_n455  &  n_n518 ) ;
 assign wire13505 = ( n_n4464 ) | ( n_n4463 ) | ( wire13503 ) ;
 assign wire13506 = ( n_n4477 ) | ( n_n4475 ) | ( n_n4476 ) | ( wire13504 ) ;
 assign wire13508 = ( i_9_  &  n_n509  &  n_n536  &  n_n534 ) | ( (~ i_9_)  &  n_n509  &  n_n536  &  n_n534 ) ;
 assign wire13509 = ( wire156 ) | ( wire67 ) ;
 assign wire13510 = ( n_n4337 ) | ( wire53 ) | ( wire13508 ) ;
 assign wire13512 = ( i_9_  &  n_n536  &  n_n524  &  n_n535 ) | ( (~ i_9_)  &  n_n536  &  n_n524  &  n_n535 ) ;
 assign wire13513 = ( wire16  &  n_n526  &  n_n535 ) | ( wire16  &  n_n526  &  n_n518 ) ;
 assign wire13515 = ( wire283 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire13516 = ( n_n4316 ) | ( n_n4313 ) | ( wire13513 ) ;
 assign wire13519 = ( n_n2446 ) | ( n_n4279 ) | ( wire13516 ) ;
 assign wire13520 = ( wire363 ) | ( wire13509 ) | ( wire13510 ) | ( wire13515 ) ;
 assign wire13521 = ( n_n4372 ) | ( n_n4373 ) | ( n_n4374 ) ;
 assign wire13522 = ( n_n4381 ) | ( wire423 ) | ( n_n4375 ) | ( wire12449 ) ;
 assign wire13523 = ( wire22  &  n_n509  &  n_n536 ) | ( wire20  &  n_n509  &  n_n536 ) ;
 assign wire13524 = ( n_n4352 ) | ( n_n4351 ) | ( n_n4356 ) | ( n_n4355 ) ;
 assign wire13525 = ( n_n4349 ) | ( n_n4350 ) | ( n_n4348 ) | ( wire13523 ) ;
 assign wire13526 = ( wire22  &  n_n536  &  n_n473 ) | ( wire25  &  n_n536  &  n_n473 ) ;
 assign wire13528 = ( n_n4411 ) | ( n_n4412 ) | ( wire79 ) ;
 assign wire13529 = ( n_n4416 ) | ( n_n4415 ) | ( n_n4414 ) | ( wire13526 ) ;
 assign wire13531 = ( n_n4393 ) | ( n_n4390 ) | ( n_n4394 ) ;
 assign wire13532 = ( wire420 ) | ( wire425 ) ;
 assign wire13534 = ( wire21  &  n_n536  &  n_n482 ) | ( wire22  &  n_n536  &  n_n482 ) ;
 assign wire13535 = ( wire16  &  n_n522  &  n_n482 ) | ( wire16  &  n_n526  &  n_n482 ) ;
 assign wire13538 = ( n_n4396 ) | ( n_n4405 ) | ( n_n4406 ) | ( wire13535 ) ;
 assign wire13539 = ( n_n4397 ) | ( n_n4398 ) | ( wire13534 ) | ( wire13538 ) ;
 assign wire13541 = ( wire22  &  n_n536  &  n_n500 ) | ( wire11  &  n_n536  &  n_n500 ) ;
 assign wire13542 = ( wire16  &  n_n524  &  n_n500 ) | ( wire16  &  n_n500  &  n_n534 ) ;
 assign wire13543 = ( n_n4361 ) | ( n_n4359 ) | ( wire13541 ) ;
 assign wire13544 = ( n_n4365 ) | ( wire13055 ) | ( wire13542 ) ;
 assign wire13546 = ( wire13521 ) | ( wire13522 ) | ( wire13524 ) | ( wire13525 ) ;
 assign wire13547 = ( wire13543 ) | ( wire13544 ) | ( wire13546 ) ;
 assign wire13550 = ( n_n4451 ) | ( n_n4462 ) | ( wire12471 ) | ( wire13425 ) ;
 assign wire13552 = ( wire13487 ) | ( wire13488 ) | ( wire13505 ) | ( wire13506 ) ;
 assign wire13553 = ( n_n4455 ) | ( wire403 ) | ( wire13550 ) | ( wire13552 ) ;
 assign wire13554 = ( wire13438 ) | ( wire13439 ) | ( wire13501 ) | ( wire13502 ) ;
 assign wire13557 = ( wire19  &  n_n473  &  n_n524 ) | ( wire19  &  n_n473  &  n_n520 ) ;
 assign wire13559 = ( wire19  &  n_n464  &  n_n528 ) | ( wire19  &  n_n464  &  n_n534 ) ;
 assign wire13560 = ( wire22  &  n_n464  &  n_n65 ) | ( wire11  &  n_n464  &  n_n65 ) ;
 assign wire13561 = ( wire19  &  n_n464  &  n_n526 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire13562 = ( i_9_  &  n_n464  &  n_n520  &  n_n65 ) | ( (~ i_9_)  &  n_n464  &  n_n520  &  n_n65 ) ;
 assign wire13566 = ( n_n5321 ) | ( n_n5313 ) | ( n_n5319 ) | ( wire13562 ) ;
 assign wire13567 = ( wire175 ) | ( wire13559 ) | ( wire13560 ) | ( wire13561 ) ;
 assign wire13569 = ( n_n4010 ) | ( n_n4009 ) | ( n_n3996 ) | ( wire13188 ) ;
 assign wire13572 = ( wire13421 ) | ( wire13422 ) | ( wire13424 ) | ( wire13569 ) ;
 assign wire13573 = ( n_n3990 ) | ( n_n3992 ) | ( n_n3988 ) | ( n_n3987 ) ;
 assign wire13576 = ( wire12  &  n_n526  &  n_n500 ) | ( wire12  &  n_n526  &  n_n518 ) ;
 assign wire13577 = ( wire11  &  n_n509  &  n_n130 ) | ( wire15  &  n_n509  &  n_n130 ) ;
 assign wire13580 = ( n_n5144 ) | ( wire422 ) | ( wire13577 ) ;
 assign wire13585 = ( n_n5240 ) | ( n_n5222 ) | ( n_n5227 ) ;
 assign wire13586 = ( n_n5236 ) | ( n_n5278 ) | ( n_n5260 ) | ( n_n5286 ) ;
 assign wire13591 = ( n_n5297 ) | ( n_n5289 ) | ( n_n5298 ) ;
 assign wire13592 = ( n_n5293 ) | ( n_n5296 ) | ( n_n5323 ) | ( n_n5311 ) ;
 assign wire13598 = ( n_n4927 ) | ( n_n4958 ) | ( n_n4961 ) ;
 assign wire13599 = ( n_n4920 ) | ( n_n4987 ) | ( n_n4963 ) | ( n_n4974 ) ;
 assign wire13601 = ( wire18  &  n_n530  &  n_n482 ) | ( wire18  &  n_n482  &  n_n534 ) ;
 assign wire13606 = ( n_n5017 ) | ( n_n5037 ) | ( n_n5015 ) | ( n_n5056 ) ;
 assign wire13607 = ( n_n5047 ) | ( n_n5020 ) | ( n_n5021 ) | ( wire13601 ) ;
 assign wire13611 = ( n_n5156 ) | ( n_n5191 ) | ( n_n5175 ) | ( n_n5177 ) ;
 assign wire13612 = ( n_n5190 ) | ( wire107 ) | ( n_n5194 ) | ( n_n5213 ) ;
 assign wire13616 = ( wire13606 ) | ( wire13607 ) | ( wire13611 ) | ( wire13612 ) ;
 assign wire13617 = ( n_n3926 ) | ( n_n3924 ) | ( n_n3923 ) | ( n_n3928 ) ;
 assign wire13622 = ( n_n4388 ) | ( n_n4407 ) | ( n_n4402 ) ;
 assign wire13623 = ( n_n4371 ) | ( n_n4392 ) | ( n_n4391 ) | ( n_n4399 ) ;
 assign wire13629 = ( n_n4724 ) | ( n_n4679 ) | ( n_n4686 ) ;
 assign wire13630 = ( n_n4663 ) | ( n_n4665 ) | ( n_n4672 ) | ( n_n4707 ) ;
 assign wire13635 = ( n_n4842 ) | ( n_n4867 ) | ( n_n4841 ) ;
 assign wire13636 = ( n_n4913 ) | ( n_n4903 ) | ( n_n4905 ) | ( n_n4846 ) ;
 assign wire13638 = ( wire15  &  n_n509  &  n_n325 ) | ( wire15  &  n_n482  &  n_n325 ) ;
 assign wire13643 = ( n_n4748 ) | ( n_n4725 ) | ( n_n4788 ) | ( n_n4802 ) ;
 assign wire13644 = ( n_n4765 ) | ( n_n4808 ) | ( n_n4742 ) | ( wire13638 ) ;
 assign wire13648 = ( wire10  &  n_n522  &  n_n535 ) | ( wire10  &  n_n526  &  n_n535 ) ;
 assign wire13650 = ( n_n4570 ) | ( n_n4557 ) | ( n_n4553 ) | ( n_n4558 ) ;
 assign wire13651 = ( n_n4549 ) | ( n_n4551 ) | ( n_n4552 ) | ( wire13648 ) ;
 assign wire13656 = ( n_n4617 ) | ( n_n4637 ) | ( n_n4613 ) | ( n_n4602 ) ;
 assign wire13657 = ( n_n4611 ) | ( n_n4639 ) | ( n_n4608 ) | ( wire139 ) ;
 assign wire13660 = ( wire24  &  n_n455  &  n_n491 ) | ( wire15  &  n_n455  &  n_n491 ) ;
 assign wire13662 = ( n_n4521 ) | ( n_n4544 ) | ( n_n4520 ) ;
 assign wire13663 = ( n_n4504 ) | ( n_n4535 ) | ( wire13660 ) ;
 assign wire13665 = ( n_n4540 ) | ( n_n4498 ) | ( wire13662 ) | ( wire13663 ) ;
 assign wire13666 = ( wire13650 ) | ( wire13651 ) | ( wire13656 ) | ( wire13657 ) ;
 assign wire13670 = ( wire13  &  n_n509  &  n_n526 ) | ( wire13  &  n_n509  &  n_n534 ) ;
 assign wire13672 = ( n_n4470 ) | ( n_n4473 ) | ( n_n4413 ) | ( n_n4457 ) ;
 assign wire13673 = ( n_n4459 ) | ( n_n4420 ) | ( n_n4410 ) | ( wire13670 ) ;
 assign wire13674 = ( wire20  &  n_n536  &  n_n535 ) | ( wire15  &  n_n536  &  n_n535 ) ;
 assign wire13679 = ( n_n4368 ) | ( n_n4358 ) | ( n_n4354 ) | ( wire124 ) ;
 assign wire13681 = ( n_n3936 ) | ( n_n3937 ) | ( wire13672 ) | ( wire13673 ) ;
 assign wire13683 = ( wire13616 ) | ( wire13617 ) | ( wire13681 ) ;
 assign wire13684 = ( n_n3920 ) | ( wire13665 ) | ( wire13666 ) | ( wire13683 ) ;
 assign wire13689 = ( n_n4339 ) | ( n_n4401 ) | ( n_n4314 ) | ( n_n4389 ) ;
 assign wire13690 = ( n_n4369 ) | ( n_n4381 ) | ( n_n4340 ) | ( wire280 ) ;
 assign wire13694 = ( wire25  &  n_n500  &  n_n130 ) | ( wire25  &  n_n491  &  n_n130 ) ;
 assign wire13696 = ( n_n5142 ) | ( n_n5107 ) | ( n_n5130 ) | ( n_n5123 ) ;
 assign wire13697 = ( n_n5101 ) | ( n_n5110 ) | ( n_n5156 ) | ( wire13694 ) ;
 assign wire13698 = ( i_9_  &  n_n520  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n520  &  n_n518  &  n_n65 ) ;
 assign wire13703 = ( n_n5182 ) | ( n_n5173 ) | ( n_n5165 ) | ( n_n5230 ) ;
 assign wire13704 = ( n_n5166 ) | ( n_n5163 ) | ( n_n5214 ) | ( wire13698 ) ;
 assign wire13709 = ( n_n5293 ) | ( n_n5240 ) | ( n_n5261 ) ;
 assign wire13710 = ( n_n5274 ) | ( n_n5300 ) | ( n_n5254 ) | ( n_n5287 ) ;
 assign wire13713 = ( n_n5305 ) | ( n_n5302 ) | ( n_n5303 ) ;
 assign wire13714 = ( wire13703 ) | ( wire13704 ) | ( wire13713 ) ;
 assign wire13717 = ( wire23  &  n_n473  &  n_n195 ) | ( wire23  &  n_n464  &  n_n195 ) ;
 assign wire13719 = ( n_n5085 ) | ( n_n5072 ) | ( n_n5082 ) | ( n_n5075 ) ;
 assign wire13720 = ( n_n5096 ) | ( n_n5099 ) | ( n_n5065 ) | ( wire13717 ) ;
 assign wire13725 = ( n_n4996 ) | ( n_n4987 ) | ( n_n5006 ) ;
 assign wire13726 = ( n_n5056 ) | ( n_n4994 ) | ( n_n5002 ) | ( n_n5053 ) ;
 assign wire13728 = ( n_n5033 ) | ( n_n5051 ) | ( wire13725 ) | ( wire13726 ) ;
 assign wire13729 = ( wire13696 ) | ( wire13697 ) | ( wire13719 ) | ( wire13720 ) ;
 assign wire13735 = ( n_n4437 ) | ( n_n4487 ) | ( n_n4409 ) | ( n_n4472 ) ;
 assign wire13736 = ( n_n4484 ) | ( n_n4462 ) | ( n_n4428 ) | ( wire403 ) ;
 assign wire13741 = ( n_n4539 ) | ( n_n4544 ) | ( n_n4533 ) | ( n_n4507 ) ;
 assign wire13742 = ( n_n4532 ) | ( n_n4499 ) | ( n_n4545 ) | ( wire471 ) ;
 assign wire13746 = ( n_n4724 ) | ( n_n4799 ) | ( n_n4723 ) ;
 assign wire13747 = ( n_n4779 ) | ( n_n4786 ) | ( n_n4755 ) | ( n_n4781 ) ;
 assign wire13752 = ( n_n4633 ) | ( n_n4635 ) | ( n_n4630 ) ;
 assign wire13753 = ( n_n4571 ) | ( n_n4578 ) | ( n_n4570 ) | ( n_n4594 ) ;
 assign wire13755 = ( wire24  &  n_n535  &  n_n325 ) | ( wire25  &  n_n535  &  n_n325 ) ;
 assign wire13756 = ( wire10  &  n_n526  &  n_n491 ) | ( wire10  &  n_n528  &  n_n491 ) ;
 assign wire13759 = ( n_n4662 ) | ( n_n4683 ) | ( wire13756 ) ;
 assign wire13760 = ( n_n4663 ) | ( n_n4685 ) | ( n_n4696 ) | ( wire13755 ) ;
 assign wire13765 = ( wire18  &  n_n522  &  n_n518 ) | ( wire18  &  n_n530  &  n_n518 ) ;
 assign wire13767 = ( n_n4977 ) | ( n_n4920 ) | ( n_n4922 ) | ( n_n4959 ) ;
 assign wire13768 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4953 ) | ( wire13765 ) ;
 assign wire13772 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4818 ) ;
 assign wire13773 = ( n_n4816 ) | ( n_n4811 ) | ( n_n4828 ) | ( n_n4842 ) ;
 assign wire13776 = ( wire11  &  n_n518  &  n_n260 ) | ( wire20  &  n_n518  &  n_n260 ) ;
 assign wire13777 = ( wire17  &  n_n509  &  n_n526 ) | ( wire17  &  n_n526  &  n_n482 ) ;
 assign wire13779 = ( n_n4900 ) | ( n_n4849 ) | ( n_n4896 ) ;
 assign wire13780 = ( wire13777 ) | ( wire13776 ) ;
 assign wire13782 = ( n_n4908 ) | ( n_n4891 ) | ( wire13779 ) | ( wire13780 ) ;
 assign wire13788 = ( n_n4784 ) | ( n_n4783 ) | ( wire292 ) ;
 assign wire13789 = ( n_n4782 ) | ( wire131 ) | ( n_n4789 ) | ( n_n4788 ) ;
 assign wire13790 = ( n_n4759 ) | ( wire14  &  n_n491  &  n_n530 ) ;
 assign wire13791 = ( n_n4765 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire13792 = ( n_n4760 ) | ( n_n4758 ) | ( wire164 ) ;
 assign wire13796 = ( n_n2130 ) | ( n_n4204 ) | ( n_n3469 ) | ( wire13790 ) ;
 assign wire13797 = ( wire13788 ) | ( wire13789 ) | ( wire13791 ) | ( wire13792 ) ;
 assign wire13798 = ( wire14  &  n_n473  &  n_n526 ) | ( wire14  &  n_n473  &  n_n532 ) ;
 assign wire13800 = ( n_n4801 ) | ( n_n4802 ) | ( wire380 ) ;
 assign wire13801 = ( n_n4795 ) | ( wire158 ) | ( wire13798 ) ;
 assign wire13803 = ( n_n4825 ) | ( n_n4815 ) | ( n_n4826 ) ;
 assign wire13804 = ( n_n4830 ) | ( wire186 ) | ( wire693 ) ;
 assign wire13807 = ( i_9_  &  n_n534  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n534  &  n_n518  &  n_n260 ) ;
 assign wire13808 = ( wire13807 ) | ( wire17  &  n_n535  &  n_n520 ) ;
 assign wire13810 = ( wire21  &  n_n509  &  n_n260 ) | ( wire20  &  n_n509  &  n_n260 ) ;
 assign wire13812 = ( wire245 ) | ( wire40 ) ;
 assign wire13813 = ( n_n4857 ) | ( n_n4860 ) | ( n_n4866 ) | ( wire13810 ) ;
 assign wire13815 = ( wire24  &  n_n518  &  n_n260 ) | ( wire15  &  n_n518  &  n_n260 ) ;
 assign wire13816 = ( wire17  &  n_n526  &  n_n518 ) | ( wire17  &  n_n528  &  n_n518 ) ;
 assign wire13818 = ( n_n4856 ) | ( n_n4850 ) | ( wire13815 ) ;
 assign wire13820 = ( wire102 ) | ( n_n4852 ) | ( wire13816 ) | ( wire13818 ) ;
 assign wire13823 = ( n_n4806 ) | ( n_n4810 ) | ( n_n4805 ) | ( wire773 ) ;
 assign wire13824 = ( wire85 ) | ( n_n4807 ) | ( n_n4808 ) | ( wire12225 ) ;
 assign wire13825 = ( wire13824 ) | ( wire13823 ) ;
 assign wire13827 = ( n_n3330 ) | ( wire13800 ) | ( wire13801 ) | ( wire13825 ) ;
 assign wire13833 = ( n_n4976 ) | ( n_n4981 ) | ( wire251 ) ;
 assign wire13834 = ( n_n4988 ) | ( n_n4985 ) | ( n_n4984 ) | ( wire57 ) ;
 assign wire13836 = ( n_n4975 ) | ( n_n4968 ) | ( wire771 ) | ( wire772 ) ;
 assign wire13837 = ( wire21  &  n_n464  &  n_n260 ) | ( wire20  &  n_n464  &  n_n260 ) ;
 assign wire13840 = ( wire13837 ) | ( wire342 ) ;
 assign wire13841 = ( n_n4974 ) | ( n_n4948 ) | ( n_n4957 ) | ( n_n4971 ) ;
 assign wire13843 = ( n_n4965 ) | ( wire13215 ) | ( wire13836 ) | ( wire13841 ) ;
 assign wire13844 = ( n_n3803 ) | ( wire13833 ) | ( wire13834 ) | ( wire13840 ) ;
 assign wire13850 = ( n_n4881 ) | ( n_n4878 ) | ( n_n4880 ) | ( n_n4877 ) ;
 assign wire13854 = ( wire25  &  n_n491  &  n_n260 ) | ( wire25  &  n_n482  &  n_n260 ) ;
 assign wire13855 = ( n_n4898 ) | ( n_n4901 ) | ( n_n4904 ) | ( n_n4897 ) ;
 assign wire13856 = ( n_n4902 ) | ( n_n4907 ) | ( wire49 ) ;
 assign wire13857 = ( n_n4909 ) | ( n_n4894 ) | ( wire13854 ) ;
 assign wire13860 = ( n_n3450 ) | ( n_n3451 ) | ( wire13857 ) ;
 assign wire13865 = ( n_n4927 ) | ( n_n4926 ) | ( n_n4925 ) | ( n_n4934 ) ;
 assign wire13866 = ( wire31 ) | ( n_n4930 ) | ( n_n4933 ) | ( n_n4931 ) ;
 assign wire13867 = ( wire22  &  n_n464  &  n_n260 ) | ( wire11  &  n_n464  &  n_n260 ) ;
 assign wire13869 = ( n_n4919 ) | ( wire17  &  n_n528  &  n_n482 ) ;
 assign wire13870 = ( n_n4911 ) | ( n_n4916 ) | ( n_n4918 ) | ( n_n4917 ) ;
 assign wire13872 = ( wire25  &  n_n473  &  n_n260 ) | ( wire23  &  n_n473  &  n_n260 ) ;
 assign wire13873 = ( n_n4923 ) | ( n_n4924 ) | ( n_n4937 ) | ( n_n4938 ) ;
 assign wire13874 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) | ( wire13872 ) ;
 assign wire13877 = ( wire58 ) | ( wire13865 ) | ( wire13866 ) | ( wire13873 ) ;
 assign wire13878 = ( wire13869 ) | ( wire13870 ) | ( wire13874 ) | ( wire13877 ) ;
 assign wire13880 = ( wire14  &  n_n524  &  n_n500 ) | ( wire14  &  n_n500  &  n_n534 ) ;
 assign wire13881 = ( wire20  &  n_n500  &  n_n325 ) | ( wire15  &  n_n500  &  n_n325 ) ;
 assign wire13883 = ( n_n4748 ) | ( n_n4747 ) | ( wire13880 ) ;
 assign wire13884 = ( n_n4756 ) | ( wire109 ) | ( wire13881 ) ;
 assign wire13885 = ( wire11  &  n_n390  &  n_n482 ) | ( wire25  &  n_n390  &  n_n482 ) ;
 assign wire13887 = ( wire391 ) | ( wire140 ) ;
 assign wire13888 = ( wire311 ) | ( n_n4654 ) | ( wire13885 ) ;
 assign wire13891 = ( n_n4669 ) | ( n_n4670 ) | ( wire72 ) ;
 assign wire13892 = ( n_n4671 ) | ( wire418 ) | ( n_n4672 ) ;
 assign wire13893 = ( n_n4673 ) | ( n_n4658 ) | ( n_n4684 ) | ( n_n4665 ) ;
 assign wire13895 = ( n_n4674 ) | ( n_n4677 ) | ( wire11855 ) | ( wire13893 ) ;
 assign wire13896 = ( wire13887 ) | ( wire13888 ) | ( wire13891 ) | ( wire13892 ) ;
 assign wire13897 = ( wire14  &  n_n522  &  n_n535 ) | ( wire14  &  n_n524  &  n_n535 ) ;
 assign wire13900 = ( wire10  &  n_n464  &  n_n526 ) | ( wire10  &  n_n464  &  n_n528 ) ;
 assign wire13902 = ( n_n4690 ) | ( n_n4689 ) | ( wire442 ) ;
 assign wire13903 = ( n_n4694 ) | ( wire445 ) | ( wire13900 ) ;
 assign wire13904 = ( n_n4711 ) | ( wire11  &  n_n325  &  n_n518 ) ;
 assign wire13905 = ( n_n4718 ) | ( n_n4717 ) | ( n_n4716 ) ;
 assign wire13906 = ( n_n4710 ) | ( n_n4709 ) | ( wire366 ) ;
 assign wire13910 = ( wire457 ) | ( n_n3124 ) | ( n_n2378 ) | ( wire13904 ) ;
 assign wire13911 = ( wire13902 ) | ( wire13903 ) | ( wire13905 ) | ( wire13906 ) ;
 assign wire13913 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4729 ) ;
 assign wire13914 = ( wire244 ) | ( n_n4732 ) | ( wire767 ) ;
 assign wire13915 = ( n_n4727 ) | ( wire95 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign wire13918 = ( wire13883 ) | ( wire13884 ) | ( wire13913 ) | ( wire13914 ) ;
 assign wire13919 = ( wire456 ) | ( wire13915 ) | ( wire13918 ) ;
 assign wire13920 = ( wire13895 ) | ( wire13896 ) | ( wire13910 ) | ( wire13911 ) ;
 assign wire13923 = ( n_n5121 ) | ( n_n5122 ) | ( n_n5126 ) ;
 assign wire13924 = ( n_n5131 ) | ( n_n5124 ) | ( n_n5127 ) | ( n_n5132 ) ;
 assign wire13929 = ( n_n5111 ) | ( n_n5112 ) | ( wire335 ) ;
 assign wire13931 = ( wire19  &  n_n473  &  n_n528 ) | ( wire19  &  n_n473  &  n_n520 ) ;
 assign wire13932 = ( wire19  &  n_n522  &  n_n473 ) | ( wire19  &  n_n473  &  n_n524 ) ;
 assign wire13934 = ( wire13931 ) | ( wire459 ) ;
 assign wire13935 = ( n_n5320 ) | ( n_n5321 ) | ( n_n5319 ) | ( wire13932 ) ;
 assign wire13938 = ( wire21  &  n_n482  &  n_n65 ) | ( wire22  &  n_n482  &  n_n65 ) ;
 assign wire13940 = ( wire19  &  n_n473  &  n_n530 ) | ( wire19  &  n_n473  &  n_n534 ) ;
 assign wire13942 = ( n_n5306 ) | ( n_n5309 ) | ( wire13938 ) ;
 assign wire13943 = ( wire200 ) | ( wire656 ) | ( wire13940 ) ;
 assign wire13944 = ( i_9_  &  n_n464  &  n_n526  &  n_n65 ) | ( (~ i_9_)  &  n_n464  &  n_n526  &  n_n65 ) ;
 assign wire13947 = ( n_n2274 ) | ( n_n2643 ) | ( n_n5330 ) | ( wire13944 ) ;
 assign wire13948 = ( wire13934 ) | ( wire13935 ) | ( wire13942 ) | ( wire13943 ) ;
 assign wire13951 = ( wire181 ) | ( wire384 ) ;
 assign wire13952 = ( n_n5222 ) | ( n_n5225 ) | ( wire385 ) | ( wire87 ) ;
 assign wire13954 = ( wire434 ) | ( wire446 ) ;
 assign wire13955 = ( n_n5255 ) | ( wire433 ) | ( n_n5247 ) | ( n_n5250 ) ;
 assign wire13957 = ( i_9_  &  n_n524  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n65 ) ;
 assign wire13960 = ( n_n5244 ) | ( n_n5243 ) | ( n_n5246 ) | ( wire13957 ) ;
 assign wire13961 = ( n_n5232 ) | ( n_n5241 ) | ( wire386 ) | ( wire13960 ) ;
 assign wire13962 = ( wire13951 ) | ( wire13952 ) | ( wire13954 ) | ( wire13955 ) ;
 assign wire13963 = ( i_9_  &  n_n524  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n500  &  n_n65 ) ;
 assign wire13964 = ( wire19  &  n_n528  &  n_n500 ) | ( wire19  &  n_n500  &  n_n530 ) ;
 assign wire13966 = ( n_n5270 ) | ( n_n5269 ) | ( wire13963 ) ;
 assign wire13967 = ( wire62 ) | ( wire92 ) | ( wire13964 ) ;
 assign wire13968 = ( wire218 ) | ( wire19  &  n_n526  &  n_n491 ) ;
 assign wire13969 = ( i_9_  &  n_n528  &  n_n482  &  n_n65 ) | ( (~ i_9_)  &  n_n528  &  n_n482  &  n_n65 ) ;
 assign wire13970 = ( n_n5288 ) | ( wire24  &  n_n482  &  n_n65 ) ;
 assign wire13971 = ( n_n5290 ) | ( n_n5286 ) | ( n_n5289 ) ;
 assign wire13972 = ( wire13969 ) | ( wire441 ) ;
 assign wire13975 = ( wire204 ) | ( wire13966 ) | ( wire13967 ) | ( wire13968 ) ;
 assign wire13976 = ( wire13970 ) | ( wire13971 ) | ( wire13972 ) | ( wire13975 ) ;
 assign wire13977 = ( wire13947 ) | ( wire13948 ) | ( wire13961 ) | ( wire13962 ) ;
 assign wire13978 = ( wire18  &  n_n522  &  n_n473 ) | ( wire18  &  n_n473  &  n_n532 ) ;
 assign wire13979 = ( i_9_  &  n_n473  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n473  &  n_n528  &  n_n195 ) ;
 assign wire13981 = ( n_n5057 ) | ( n_n5058 ) | ( wire13978 ) ;
 assign wire13982 = ( n_n5059 ) | ( n_n5064 ) | ( wire755 ) | ( wire13979 ) ;
 assign wire13983 = ( wire18  &  n_n524  &  n_n482 ) | ( wire18  &  n_n528  &  n_n482 ) ;
 assign wire13985 = ( wire18  &  n_n473  &  n_n534 ) | ( wire18  &  n_n482  &  n_n534 ) ;
 assign wire13989 = ( n_n5025 ) | ( n_n5028 ) | ( n_n5036 ) | ( wire13399 ) ;
 assign wire13990 = ( wire50 ) | ( wire231 ) | ( wire356 ) | ( wire13985 ) ;
 assign wire13991 = ( n_n5039 ) | ( wire97 ) | ( wire13983 ) | ( wire13989 ) ;
 assign wire13992 = ( wire13981 ) | ( wire13982 ) | ( wire13990 ) ;
 assign wire13995 = ( n_n5018 ) | ( n_n5019 ) | ( n_n5015 ) | ( n_n5020 ) ;
 assign wire13996 = ( n_n5016 ) | ( n_n5024 ) | ( n_n5021 ) | ( wire13400 ) ;
 assign wire13997 = ( i_9_  &  n_n509  &  n_n528  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n195 ) ;
 assign wire13999 = ( wire248 ) | ( wire103 ) ;
 assign wire14000 = ( n_n4998 ) | ( n_n4993 ) | ( n_n4989 ) | ( wire13997 ) ;
 assign wire14001 = ( i_9_  &  n_n526  &  n_n518  &  n_n130 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n130 ) ;
 assign wire14003 = ( wire18  &  n_n522  &  n_n464 ) | ( wire18  &  n_n524  &  n_n464 ) ;
 assign wire14006 = ( n_n5081 ) | ( n_n5069 ) | ( wire14003 ) ;
 assign wire14007 = ( n_n5083 ) | ( wire160 ) | ( n_n5077 ) | ( n_n5071 ) ;
 assign wire14009 = ( i_9_  &  n_n535  &  n_n528  &  n_n130 ) | ( (~ i_9_)  &  n_n535  &  n_n528  &  n_n130 ) ;
 assign wire14010 = ( n_n5098 ) | ( n_n5084 ) | ( n_n5095 ) ;
 assign wire14011 = ( n_n5097 ) | ( n_n5089 ) | ( wire232 ) ;
 assign wire14012 = ( n_n5106 ) | ( wire14001 ) | ( wire14009 ) ;
 assign wire14015 = ( n_n1167 ) | ( wire88 ) | ( wire12917 ) | ( wire14012 ) ;
 assign wire14016 = ( wire14006 ) | ( wire14007 ) | ( wire14010 ) | ( wire14011 ) ;
 assign wire14018 = ( wire21  &  n_n500  &  n_n195 ) | ( wire24  &  n_n500  &  n_n195 ) ;
 assign wire14020 = ( n_n5005 ) | ( n_n5010 ) | ( wire14018 ) ;
 assign wire14021 = ( n_n5013 ) | ( n_n5008 ) | ( n_n5007 ) | ( wire12931 ) ;
 assign wire14023 = ( wire13995 ) | ( wire13996 ) | ( wire13999 ) | ( wire14000 ) ;
 assign wire14024 = ( wire14020 ) | ( wire14021 ) | ( wire14023 ) ;
 assign wire14025 = ( wire13991 ) | ( wire13992 ) | ( wire14015 ) | ( wire14016 ) ;
 assign wire14027 = ( wire22  &  n_n473  &  n_n130 ) | ( wire11  &  n_n473  &  n_n130 ) ;
 assign wire14028 = ( n_n5181 ) | ( n_n5184 ) | ( wire112 ) ;
 assign wire14029 = ( wire114 ) | ( wire765 ) | ( wire14027 ) ;
 assign wire14031 = ( wire12  &  n_n524  &  n_n491 ) | ( wire12  &  n_n528  &  n_n491 ) ;
 assign wire14033 = ( n_n5157 ) | ( n_n5158 ) | ( wire196 ) ;
 assign wire14034 = ( n_n5147 ) | ( wire76 ) | ( wire14031 ) ;
 assign wire14036 = ( wire11  &  n_n482  &  n_n130 ) | ( wire25  &  n_n482  &  n_n130 ) ;
 assign wire14037 = ( wire12  &  n_n530  &  n_n482 ) | ( wire12  &  n_n482  &  n_n532 ) ;
 assign wire14040 = ( n_n5175 ) | ( n_n5177 ) | ( n_n5176 ) | ( wire14037 ) ;
 assign wire14041 = ( n_n5171 ) | ( n_n5174 ) | ( wire14036 ) | ( wire14040 ) ;
 assign wire14042 = ( wire14028 ) | ( wire14029 ) | ( wire14033 ) | ( wire14034 ) ;
 assign wire14043 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n524  &  n_n535 ) ;
 assign wire14045 = ( wire449 ) | ( n_n5210 ) | ( n_n5209 ) ;
 assign wire14046 = ( n_n5212 ) | ( n_n5219 ) | ( n_n5211 ) | ( wire14043 ) ;
 assign wire14047 = ( wire12  &  n_n464  &  n_n526 ) | ( wire12  &  n_n464  &  n_n520 ) ;
 assign wire14049 = ( n_n5201 ) | ( n_n5207 ) | ( n_n5208 ) | ( wire761 ) ;
 assign wire14050 = ( n_n5203 ) | ( wire220 ) | ( wire14047 ) ;
 assign wire14055 = ( n_n5193 ) | ( n_n5189 ) | ( n_n5188 ) | ( n_n5199 ) ;
 assign wire14056 = ( n_n5197 ) | ( wire451 ) | ( n_n5198 ) | ( n_n5192 ) ;
 assign wire14057 = ( wire14056 ) | ( wire14055 ) ;
 assign wire14058 = ( wire14045 ) | ( wire14046 ) | ( wire14049 ) | ( wire14050 ) ;
 assign wire14061 = ( n_n5146 ) | ( n_n5138 ) | ( wire211 ) ;
 assign wire14062 = ( n_n5133 ) | ( n_n5144 ) | ( n_n5143 ) | ( wire12883 ) ;
 assign wire14065 = ( n_n3307 ) | ( n_n3308 ) | ( wire14061 ) | ( wire14062 ) ;
 assign wire14066 = ( wire14041 ) | ( wire14042 ) | ( wire14057 ) | ( wire14058 ) ;
 assign wire14068 = ( wire13976 ) | ( wire13977 ) | ( wire14024 ) | ( wire14025 ) ;
 assign wire14071 = ( n_n4607 ) | ( n_n4612 ) | ( n_n4609 ) ;
 assign wire14072 = ( n_n4617 ) | ( n_n4613 ) | ( wire396 ) ;
 assign wire14077 = ( wire309 ) | ( wire118 ) ;
 assign wire14078 = ( n_n4639 ) | ( n_n4642 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign wire14079 = ( n_n4641 ) | ( n_n4634 ) | ( n_n4648 ) | ( n_n4618 ) ;
 assign wire14080 = ( n_n4628 ) | ( wire26 ) | ( n_n4625 ) | ( wire12545 ) ;
 assign wire14082 = ( wire14080 ) | ( wire14079 ) ;
 assign wire14087 = ( n_n4597 ) | ( n_n4598 ) | ( n_n4595 ) | ( n_n4596 ) ;
 assign wire14088 = ( n_n4602 ) | ( n_n4593 ) | ( n_n4601 ) | ( wire108 ) ;
 assign wire14091 = ( n_n4586 ) | ( n_n4591 ) | ( n_n4592 ) ;
 assign wire14092 = ( n_n4590 ) | ( n_n4587 ) | ( wire365 ) ;
 assign wire14094 = ( wire22  &  n_n535  &  n_n390 ) | ( wire11  &  n_n535  &  n_n390 ) ;
 assign wire14097 = ( i_9_  &  n_n535  &  n_n390  &  n_n530 ) | ( (~ i_9_)  &  n_n535  &  n_n390  &  n_n530 ) ;
 assign wire14099 = ( n_n4576 ) | ( n_n4569 ) | ( n_n4574 ) | ( n_n4581 ) ;
 assign wire14101 = ( n_n4579 ) | ( wire14094 ) | ( wire14097 ) | ( wire14099 ) ;
 assign wire14103 = ( i_9_  &  n_n464  &  n_n526  &  n_n455 ) | ( (~ i_9_)  &  n_n464  &  n_n526  &  n_n455 ) ;
 assign wire14105 = ( n_n4568 ) | ( wire430 ) | ( wire783 ) ;
 assign wire14106 = ( wire213 ) | ( n_n4556 ) | ( wire14103 ) ;
 assign wire14107 = ( i_9_  &  n_n473  &  n_n524  &  n_n455 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n455 ) ;
 assign wire14111 = ( wire21  &  n_n455  &  n_n482 ) | ( wire15  &  n_n455  &  n_n482 ) ;
 assign wire14112 = ( n_n4526 ) | ( n_n4538 ) | ( n_n4535 ) | ( n_n4536 ) ;
 assign wire14115 = ( wire202 ) | ( n_n4542 ) | ( wire201 ) | ( wire14111 ) ;
 assign wire14116 = ( n_n3871 ) | ( wire14105 ) | ( wire14106 ) | ( wire14112 ) ;
 assign wire14120 = ( n_n4463 ) | ( n_n4466 ) | ( n_n4465 ) ;
 assign wire14121 = ( wire291 ) | ( wire128 ) ;
 assign wire14126 = ( n_n4491 ) | ( n_n4492 ) | ( n_n4475 ) | ( n_n4476 ) ;
 assign wire14127 = ( n_n4467 ) | ( n_n4470 ) | ( n_n4489 ) | ( n_n4469 ) ;
 assign wire14128 = ( n_n4483 ) | ( n_n4488 ) | ( n_n4471 ) | ( n_n4490 ) ;
 assign wire14131 = ( wire184 ) | ( n_n901 ) | ( wire787 ) | ( wire14128 ) ;
 assign wire14133 = ( wire13  &  n_n524  &  n_n535 ) | ( wire13  &  n_n526  &  n_n535 ) ;
 assign wire14134 = ( wire16  &  n_n524  &  n_n464 ) | ( wire16  &  n_n464  &  n_n526 ) ;
 assign wire14138 = ( n_n4431 ) | ( n_n4441 ) | ( wire14134 ) ;
 assign wire14139 = ( n_n4439 ) | ( n_n4436 ) | ( n_n4435 ) | ( wire421 ) ;
 assign wire14141 = ( wire20  &  n_n536  &  n_n473 ) | ( wire23  &  n_n536  &  n_n473 ) ;
 assign wire14142 = ( wire37 ) | ( wire16  &  n_n473  &  n_n520 ) ;
 assign wire14143 = ( n_n4420 ) | ( n_n4430 ) | ( wire84 ) ;
 assign wire14144 = ( n_n4451 ) | ( wire13425 ) | ( wire14141 ) ;
 assign wire14147 = ( wire470 ) | ( n_n4449 ) | ( wire14133 ) | ( wire14144 ) ;
 assign wire14148 = ( wire14138 ) | ( wire14139 ) | ( wire14142 ) | ( wire14143 ) ;
 assign wire14149 = ( i_9_  &  n_n536  &  n_n500  &  n_n534 ) | ( (~ i_9_)  &  n_n536  &  n_n500  &  n_n534 ) ;
 assign wire14150 = ( i_9_  &  n_n509  &  n_n522  &  n_n536 ) | ( (~ i_9_)  &  n_n509  &  n_n522  &  n_n536 ) ;
 assign wire14153 = ( wire14150 ) | ( wire14149 ) ;
 assign wire14154 = ( n_n4353 ) | ( n_n4358 ) | ( wire399 ) | ( n_n4354 ) ;
 assign wire14155 = ( i_9_  &  n_n536  &  n_n528  &  n_n491 ) | ( (~ i_9_)  &  n_n536  &  n_n528  &  n_n491 ) ;
 assign wire14157 = ( i_9_  &  n_n536  &  n_n524  &  n_n500 ) | ( (~ i_9_)  &  n_n536  &  n_n524  &  n_n500 ) ;
 assign wire14158 = ( n_n4373 ) | ( n_n4374 ) | ( n_n4368 ) ;
 assign wire14159 = ( n_n4380 ) | ( n_n4372 ) | ( wire14155 ) ;
 assign wire14160 = ( n_n4363 ) | ( n_n4364 ) | ( n_n4362 ) | ( wire14157 ) ;
 assign wire14161 = ( n_n4365 ) | ( wire423 ) | ( n_n4375 ) | ( wire11607 ) ;
 assign wire14163 = ( wire14161 ) | ( wire14160 ) ;
 assign wire14164 = ( wire14153 ) | ( wire14154 ) | ( wire14158 ) | ( wire14159 ) ;
 assign wire14168 = ( n_n4398 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign wire14169 = ( n_n4403 ) | ( n_n4400 ) | ( n_n4396 ) | ( n_n4399 ) ;
 assign wire14171 = ( wire22  &  n_n536  &  n_n473 ) | ( wire15  &  n_n536  &  n_n473 ) ;
 assign wire14173 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) ;
 assign wire14174 = ( wire14171 ) | ( wire79 ) ;
 assign wire14177 = ( i_9_  &  n_n536  &  n_n482  &  n_n532 ) | ( (~ i_9_)  &  n_n536  &  n_n482  &  n_n532 ) ;
 assign wire14178 = ( n_n4392 ) | ( n_n4384 ) | ( wire425 ) ;
 assign wire14179 = ( n_n4388 ) | ( n_n4391 ) | ( n_n4390 ) | ( wire14177 ) ;
 assign wire14183 = ( wire106 ) | ( wire198 ) ;
 assign wire14186 = ( wire364 ) | ( wire24  &  n_n536  &  n_n535 ) ;
 assign wire14191 = ( n_n4338 ) | ( n_n4337 ) | ( wire156 ) ;
 assign wire14192 = ( n_n4345 ) | ( n_n4341 ) | ( wire67 ) | ( n_n4348 ) ;
 assign wire14195 = ( n_n3369 ) | ( n_n3370 ) | ( wire14191 ) | ( wire14192 ) ;
 assign wire14198 = ( wire66 ) | ( n_n4502 ) | ( n_n4501 ) ;
 assign wire14199 = ( n_n4500 ) | ( n_n4498 ) | ( n_n4493 ) | ( wire13027 ) ;
 assign wire14200 = ( i_9_  &  n_n455  &  n_n491  &  n_n530 ) | ( (~ i_9_)  &  n_n455  &  n_n491  &  n_n530 ) ;
 assign wire14202 = ( n_n4506 ) | ( wire129 ) | ( n_n4505 ) ;
 assign wire14203 = ( n_n4511 ) | ( n_n4503 ) | ( n_n4510 ) | ( wire14200 ) ;
 assign wire14205 = ( n_n4521 ) | ( n_n4517 ) | ( n_n4520 ) ;
 assign wire14208 = ( wire14198 ) | ( wire14199 ) | ( wire14202 ) | ( wire14203 ) ;
 assign wire14209 = ( n_n4247 ) | ( n_n4246 ) | ( wire14205 ) | ( wire14208 ) ;
 assign wire14211 = ( n_n3285 ) | ( wire14147 ) | ( wire14148 ) | ( wire14209 ) ;
 assign wire14213 = ( wire149 ) | ( n_n5331 ) | ( wire12963 ) ;
 assign wire14214 = ( n_n3277 ) | ( n_n3275 ) | ( wire13827 ) | ( wire14213 ) ;
 assign wire14216 = ( n_n3257 ) | ( wire13919 ) | ( wire13920 ) | ( wire14214 ) ;
 assign wire14218 = ( wire13689 ) | ( wire13690 ) | ( wire13735 ) | ( wire13736 ) ;
 assign wire14219 = ( wire13741 ) | ( wire13742 ) | ( wire14218 ) ;
 assign wire14222 = ( n_n3187 ) | ( n_n3192 ) | ( n_n3191 ) | ( wire14219 ) ;
 assign wire14226 = ( n_n5124 ) | ( n_n5117 ) | ( wire125 ) ;
 assign wire14227 = ( n_n5135 ) | ( n_n5152 ) | ( n_n5153 ) | ( wire168 ) ;
 assign wire14232 = ( n_n5172 ) | ( n_n5207 ) | ( n_n5169 ) | ( n_n5197 ) ;
 assign wire14233 = ( wire254 ) | ( n_n5211 ) | ( n_n5176 ) | ( n_n5205 ) ;
 assign wire14238 = ( n_n5092 ) | ( n_n5110 ) | ( n_n5100 ) | ( n_n5097 ) ;
 assign wire14239 = ( n_n5087 ) | ( n_n5065 ) | ( n_n5077 ) | ( wire159 ) ;
 assign wire14240 = ( wire14239 ) | ( wire14238 ) ;
 assign wire14241 = ( wire14226 ) | ( wire14227 ) | ( wire14232 ) | ( wire14233 ) ;
 assign wire14245 = ( n_n5307 ) | ( n_n5266 ) | ( wire63 ) ;
 assign wire14246 = ( n_n5295 ) | ( n_n5290 ) | ( wire433 ) | ( n_n5283 ) ;
 assign wire14252 = ( n_n5320 ) | ( n_n5325 ) | ( wire435 ) ;
 assign wire14253 = ( n_n5232 ) | ( n_n5255 ) | ( n_n5212 ) | ( n_n5249 ) ;
 assign wire14254 = ( n_n5237 ) | ( n_n5308 ) | ( n_n5226 ) | ( n_n5218 ) ;
 assign wire14256 = ( wire14252 ) | ( wire14253 ) | ( wire14254 ) ;
 assign wire14260 = ( n_n4869 ) | ( n_n4870 ) | ( n_n4883 ) ;
 assign wire14261 = ( n_n4895 ) | ( n_n4825 ) | ( n_n4879 ) | ( n_n4841 ) ;
 assign wire14267 = ( n_n4958 ) | ( n_n4921 ) | ( n_n4963 ) | ( n_n4916 ) ;
 assign wire14268 = ( wire352 ) | ( n_n4933 ) | ( n_n4948 ) | ( n_n4973 ) ;
 assign wire14272 = ( n_n4994 ) | ( n_n5061 ) | ( wire669 ) ;
 assign wire14273 = ( n_n5034 ) | ( n_n4996 ) | ( n_n5026 ) | ( n_n4988 ) ;
 assign wire14275 = ( n_n5057 ) | ( n_n4974 ) | ( wire14272 ) | ( wire14273 ) ;
 assign wire14277 = ( wire14245 ) | ( wire14246 ) | ( wire14256 ) | ( wire14275 ) ;
 assign wire14278 = ( n_n3558 ) | ( n_n3557 ) | ( wire14240 ) | ( wire14241 ) ;
 assign wire14280 = ( wire21  &  n_n455  &  n_n535 ) | ( wire22  &  n_n455  &  n_n535 ) ;
 assign wire14281 = ( wire13  &  n_n509  &  n_n526 ) | ( wire13  &  n_n509  &  n_n520 ) ;
 assign wire14283 = ( n_n4464 ) | ( n_n4467 ) | ( wire14280 ) ;
 assign wire14284 = ( n_n4432 ) | ( n_n4435 ) | ( n_n4493 ) | ( wire14281 ) ;
 assign wire14285 = ( wire16  &  n_n522  &  n_n535 ) | ( wire16  &  n_n535  &  n_n532 ) ;
 assign wire14290 = ( n_n4317 ) | ( n_n4362 ) | ( n_n4319 ) | ( n_n4336 ) ;
 assign wire14291 = ( n_n4348 ) | ( n_n4321 ) | ( n_n4355 ) | ( wire14285 ) ;
 assign wire14293 = ( wire21  &  n_n500  &  n_n390 ) | ( wire24  &  n_n500  &  n_n390 ) ;
 assign wire14295 = ( n_n4617 ) | ( n_n4637 ) | ( n_n4638 ) | ( n_n4626 ) ;
 assign wire14296 = ( n_n4613 ) | ( n_n4610 ) | ( n_n4632 ) | ( wire14293 ) ;
 assign wire14301 = ( n_n4514 ) | ( n_n4544 ) | ( n_n4561 ) | ( n_n4522 ) ;
 assign wire14302 = ( n_n4525 ) | ( wire65 ) | ( n_n4542 ) | ( n_n4559 ) ;
 assign wire14307 = ( n_n4602 ) | ( n_n4601 ) | ( n_n4595 ) ;
 assign wire14308 = ( n_n4568 ) | ( n_n4590 ) | ( n_n4582 ) | ( n_n4581 ) ;
 assign wire14310 = ( n_n4579 ) | ( n_n4608 ) | ( wire14307 ) | ( wire14308 ) ;
 assign wire14311 = ( wire14295 ) | ( wire14296 ) | ( wire14301 ) | ( wire14302 ) ;
 assign wire14316 = ( n_n4744 ) | ( n_n4697 ) | ( n_n4721 ) ;
 assign wire14317 = ( n_n4703 ) | ( n_n4717 ) | ( n_n4736 ) | ( n_n4741 ) ;
 assign wire14320 = ( wire10  &  n_n473  &  n_n528 ) | ( wire10  &  n_n473  &  n_n520 ) ;
 assign wire14322 = ( n_n4658 ) | ( n_n4687 ) | ( wire775 ) ;
 assign wire14323 = ( n_n4646 ) | ( n_n4668 ) | ( wire14320 ) ;
 assign wire14329 = ( n_n4784 ) | ( n_n4787 ) | ( n_n4780 ) ;
 assign wire14330 = ( n_n4759 ) | ( n_n4811 ) | ( n_n4793 ) | ( n_n4778 ) ;
 assign wire14332 = ( n_n4747 ) | ( n_n4752 ) | ( wire14329 ) | ( wire14330 ) ;
 assign wire14334 = ( wire16  &  n_n500  &  n_n520 ) | ( wire16  &  n_n500  &  n_n530 ) ;
 assign wire14337 = ( n_n4406 ) | ( n_n4408 ) | ( wire14334 ) ;
 assign wire14338 = ( wire37 ) | ( n_n4409 ) | ( n_n4399 ) | ( n_n4370 ) ;
 assign wire14340 = ( wire14283 ) | ( wire14284 ) | ( wire14290 ) | ( wire14291 ) ;
 assign wire14341 = ( wire14337 ) | ( wire14338 ) | ( wire14340 ) ;
 assign wire14343 = ( n_n3548 ) | ( wire14310 ) | ( wire14311 ) | ( wire14341 ) ;
 assign wire14344 = ( wire14  &  n_n528  &  n_n518 ) | ( wire14  &  n_n520  &  n_n518 ) ;
 assign wire14346 = ( n_n4724 ) | ( n_n4723 ) | ( n_n4722 ) ;
 assign wire14347 = ( n_n4720 ) | ( n_n4719 ) | ( wire14344 ) ;
 assign wire14349 = ( wire14  &  n_n535  &  n_n528 ) | ( wire14  &  n_n535  &  n_n534 ) ;
 assign wire14350 = ( wire442 ) | ( wire221 ) ;
 assign wire14351 = ( n_n4693 ) | ( wire12422 ) | ( wire14349 ) ;
 assign wire14355 = ( n_n4704 ) | ( n_n4711 ) | ( n_n4705 ) | ( n_n4706 ) ;
 assign wire14356 = ( n_n4710 ) | ( wire366 ) | ( n_n4707 ) | ( n_n4713 ) ;
 assign wire14357 = ( wire14356 ) | ( wire14355 ) ;
 assign wire14361 = ( n_n4673 ) | ( n_n4674 ) | ( wire80 ) ;
 assign wire14362 = ( n_n4676 ) | ( n_n4679 ) | ( wire418 ) | ( n_n4672 ) ;
 assign wire14363 = ( n_n4688 ) | ( n_n4685 ) | ( n_n4686 ) ;
 assign wire14365 = ( i_9_  &  n_n473  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n473  &  n_n390  &  n_n532 ) ;
 assign wire14367 = ( i_9_  &  n_n520  &  n_n390  &  n_n482 ) | ( (~ i_9_)  &  n_n520  &  n_n390  &  n_n482 ) ;
 assign wire14369 = ( n_n4664 ) | ( n_n4669 ) | ( wire14365 ) ;
 assign wire14371 = ( wire72 ) | ( n_n4657 ) | ( wire14367 ) | ( wire14369 ) ;
 assign wire14373 = ( wire11  &  n_n491  &  n_n325 ) | ( wire25  &  n_n491  &  n_n325 ) ;
 assign wire14375 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4764 ) | ( n_n4763 ) ;
 assign wire14376 = ( n_n4765 ) | ( n_n4766 ) | ( n_n4762 ) | ( wire14373 ) ;
 assign wire14377 = ( wire21  &  n_n509  &  n_n325 ) | ( wire22  &  n_n509  &  n_n325 ) ;
 assign wire14378 = ( wire14  &  n_n509  &  n_n522 ) | ( wire14  &  n_n509  &  n_n530 ) ;
 assign wire14380 = ( wire14377 ) | ( wire244 ) ;
 assign wire14381 = ( wire95 ) | ( n_n4742 ) | ( wire14378 ) ;
 assign wire14384 = ( n_n4754 ) | ( n_n4749 ) | ( wire109 ) ;
 assign wire14385 = ( n_n4755 ) | ( n_n4743 ) | ( n_n4745 ) | ( wire11834 ) ;
 assign wire14387 = ( wire14375 ) | ( wire14376 ) | ( wire14380 ) | ( wire14381 ) ;
 assign wire14388 = ( wire14384 ) | ( wire14385 ) | ( wire14387 ) ;
 assign wire14393 = ( n_n4615 ) | ( n_n4618 ) | ( n_n4629 ) | ( n_n4630 ) ;
 assign wire14396 = ( wire10  &  n_n526  &  n_n482 ) | ( wire10  &  n_n530  &  n_n482 ) ;
 assign wire14397 = ( wire431 ) | ( wire140 ) ;
 assign wire14398 = ( n_n4648 ) | ( n_n4647 ) | ( n_n4645 ) | ( wire14396 ) ;
 assign wire14401 = ( wire21  &  n_n491  &  n_n390 ) | ( wire24  &  n_n491  &  n_n390 ) ;
 assign wire14403 = ( n_n4641 ) | ( n_n4644 ) | ( n_n4640 ) | ( n_n4639 ) ;
 assign wire14404 = ( n_n4634 ) | ( n_n4642 ) | ( n_n4631 ) | ( wire14401 ) ;
 assign wire14405 = ( wire14404 ) | ( wire14403 ) ;
 assign wire14408 = ( wire11  &  n_n473  &  n_n455 ) | ( wire25  &  n_n473  &  n_n455 ) ;
 assign wire14409 = ( n_n4539 ) | ( n_n4536 ) | ( wire201 ) ;
 assign wire14410 = ( n_n4545 ) | ( wire13091 ) | ( wire14408 ) ;
 assign wire14413 = ( wire13  &  n_n473  &  n_n520 ) | ( wire13  &  n_n464  &  n_n520 ) ;
 assign wire14414 = ( n_n4557 ) | ( wire212 ) | ( n_n4558 ) ;
 assign wire14415 = ( n_n4571 ) | ( n_n4560 ) | ( wire430 ) ;
 assign wire14416 = ( n_n4569 ) | ( n_n4556 ) | ( wire14413 ) ;
 assign wire14419 = ( n_n3871 ) | ( wire455 ) | ( wire671 ) | ( wire14416 ) ;
 assign wire14420 = ( wire14409 ) | ( wire14410 ) | ( wire14414 ) | ( wire14415 ) ;
 assign wire14422 = ( n_n4591 ) | ( n_n4592 ) | ( n_n4596 ) ;
 assign wire14423 = ( n_n4593 ) | ( n_n4594 ) | ( wire45 ) ;
 assign wire14426 = ( i_9_  &  n_n390  &  n_n532  &  n_n518 ) | ( (~ i_9_)  &  n_n390  &  n_n532  &  n_n518 ) ;
 assign wire14428 = ( n_n4578 ) | ( n_n4575 ) | ( wire99 ) ;
 assign wire14429 = ( n_n4583 ) | ( wire239 ) | ( wire14426 ) ;
 assign wire14430 = ( i_9_  &  n_n509  &  n_n528  &  n_n390 ) | ( (~ i_9_)  &  n_n509  &  n_n528  &  n_n390 ) ;
 assign wire14432 = ( n_n4612 ) | ( n_n4611 ) | ( wire14430 ) ;
 assign wire14434 = ( n_n2037 ) | ( n_n4614 ) | ( n_n4609 ) | ( wire14432 ) ;
 assign wire14436 = ( n_n3718 ) | ( wire14428 ) | ( wire14429 ) | ( wire14434 ) ;
 assign wire14438 = ( wire21  &  n_n509  &  n_n455 ) | ( wire23  &  n_n509  &  n_n455 ) ;
 assign wire14439 = ( wire13  &  n_n509  &  n_n524 ) | ( wire13  &  n_n509  &  n_n528 ) ;
 assign wire14440 = ( n_n4475 ) | ( wire199 ) | ( n_n4476 ) ;
 assign wire14441 = ( n_n4484 ) | ( wire14438 ) | ( wire14439 ) ;
 assign wire14442 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign wire14443 = ( wire13  &  n_n522  &  n_n500 ) | ( wire13  &  n_n526  &  n_n500 ) ;
 assign wire14444 = ( n_n4491 ) | ( n_n4492 ) | ( wire14442 ) ;
 assign wire14445 = ( n_n4489 ) | ( n_n4488 ) | ( n_n4490 ) | ( wire14443 ) ;
 assign wire14446 = ( wire24  &  n_n455  &  n_n482 ) | ( wire25  &  n_n455  &  n_n482 ) ;
 assign wire14448 = ( n_n4515 ) | ( wire791 ) | ( wire14446 ) ;
 assign wire14452 = ( n_n4506 ) | ( n_n4505 ) | ( n_n4529 ) ;
 assign wire14453 = ( wire378 ) | ( wire129 ) ;
 assign wire14454 = ( n_n4504 ) | ( n_n4503 ) | ( wire379 ) ;
 assign wire14455 = ( n_n4531 ) | ( n_n4507 ) | ( n_n4510 ) | ( n_n4501 ) ;
 assign wire14458 = ( n_n4534 ) | ( wire11543 ) | ( wire14452 ) | ( wire14455 ) ;
 assign wire14460 = ( wire11  &  n_n536  &  n_n491 ) | ( wire15  &  n_n536  &  n_n491 ) ;
 assign wire14461 = ( wire24  &  n_n536  &  n_n500 ) | ( wire25  &  n_n536  &  n_n500 ) ;
 assign wire14464 = ( wire16  &  n_n509  &  n_n522 ) | ( wire16  &  n_n509  &  n_n520 ) ;
 assign wire14466 = ( n_n4359 ) | ( n_n4365 ) | ( n_n4360 ) | ( n_n4352 ) ;
 assign wire14467 = ( n_n4354 ) | ( wire14461 ) | ( wire14464 ) ;
 assign wire14468 = ( wire22  &  n_n536  &  n_n500 ) | ( wire20  &  n_n536  &  n_n500 ) ;
 assign wire14470 = ( n_n4372 ) | ( n_n4371 ) | ( n_n4376 ) ;
 assign wire14471 = ( n_n4367 ) | ( n_n4368 ) | ( wire14468 ) ;
 assign wire14473 = ( wire21  &  n_n536  &  n_n518 ) | ( wire22  &  n_n536  &  n_n518 ) ;
 assign wire14476 = ( wire16  &  n_n535  &  n_n530 ) | ( wire16  &  n_n535  &  n_n534 ) ;
 assign wire14479 = ( n_n4320 ) | ( n_n4315 ) | ( wire14476 ) ;
 assign wire14480 = ( n_n4313 ) | ( n_n4322 ) | ( n_n4323 ) | ( wire106 ) ;
 assign wire14484 = ( wire156 ) | ( wire198 ) ;
 assign wire14485 = ( n_n4344 ) | ( n_n4345 ) | ( n_n4347 ) | ( wire675 ) ;
 assign wire14486 = ( n_n4341 ) | ( n_n4351 ) | ( n_n4349 ) | ( n_n4334 ) ;
 assign wire14489 = ( n_n4340 ) | ( n_n2445 ) | ( wire14473 ) | ( wire14486 ) ;
 assign wire14490 = ( wire14479 ) | ( wire14480 ) | ( wire14484 ) | ( wire14485 ) ;
 assign wire14492 = ( wire22  &  n_n536  &  n_n473 ) | ( wire20  &  n_n536  &  n_n473 ) ;
 assign wire14493 = ( i_9_  &  n_n536  &  n_n473  &  n_n528 ) | ( (~ i_9_)  &  n_n536  &  n_n473  &  n_n528 ) ;
 assign wire14495 = ( n_n4420 ) | ( n_n4419 ) | ( wire14492 ) ;
 assign wire14496 = ( n_n4418 ) | ( wire328 ) | ( wire14493 ) ;
 assign wire14498 = ( n_n4393 ) | ( n_n4396 ) | ( n_n4395 ) | ( n_n4394 ) ;
 assign wire14499 = ( n_n4391 ) | ( n_n4397 ) | ( n_n4387 ) | ( wire12448 ) ;
 assign wire14500 = ( wire21  &  n_n536  &  n_n482 ) | ( wire22  &  n_n536  &  n_n482 ) ;
 assign wire14503 = ( i_9_  &  n_n536  &  n_n473  &  n_n532 ) | ( (~ i_9_)  &  n_n536  &  n_n473  &  n_n532 ) ;
 assign wire14505 = ( n_n4400 ) | ( n_n4407 ) | ( n_n4398 ) | ( n_n4405 ) ;
 assign wire14507 = ( n_n4402 ) | ( wire14500 ) | ( wire14503 ) | ( wire14505 ) ;
 assign wire14508 = ( wire14495 ) | ( wire14496 ) | ( wire14498 ) | ( wire14499 ) ;
 assign wire14510 = ( n_n4382 ) | ( n_n4380 ) | ( n_n4379 ) | ( n_n4377 ) ;
 assign wire14511 = ( n_n4386 ) | ( wire12447 ) | ( wire14460 ) | ( wire14510 ) ;
 assign wire14513 = ( n_n3736 ) | ( wire14466 ) | ( wire14467 ) | ( wire14511 ) ;
 assign wire14514 = ( wire14489 ) | ( wire14490 ) | ( wire14507 ) | ( wire14508 ) ;
 assign wire14517 = ( n_n4455 ) | ( n_n4456 ) | ( n_n4457 ) | ( n_n4462 ) ;
 assign wire14518 = ( n_n4461 ) | ( wire13  &  n_n532  &  n_n518 ) ;
 assign wire14519 = ( i_9_  &  n_n536  &  n_n464  &  n_n530 ) | ( (~ i_9_)  &  n_n536  &  n_n464  &  n_n530 ) ;
 assign wire14520 = ( wire16  &  n_n524  &  n_n464 ) | ( wire16  &  n_n464  &  n_n532 ) ;
 assign wire14521 = ( wire215 ) | ( wire98 ) ;
 assign wire14522 = ( n_n4427 ) | ( wire14519 ) | ( wire14520 ) ;
 assign wire14523 = ( wire13  &  n_n524  &  n_n535 ) | ( wire13  &  n_n535  &  n_n534 ) ;
 assign wire14524 = ( i_9_  &  n_n455  &  n_n535  &  n_n530 ) | ( (~ i_9_)  &  n_n455  &  n_n535  &  n_n530 ) ;
 assign wire14526 = ( wire11  &  n_n455  &  n_n535 ) | ( wire24  &  n_n455  &  n_n535 ) ;
 assign wire14528 = ( n_n4442 ) | ( n_n4437 ) | ( wire14524 ) ;
 assign wire14530 = ( n_n4446 ) | ( wire14523 ) | ( wire14526 ) | ( wire14528 ) ;
 assign wire14533 = ( n_n4471 ) | ( n_n4472 ) | ( n_n4468 ) ;
 assign wire14534 = ( n_n4463 ) | ( n_n4470 ) | ( n_n4466 ) | ( n_n4469 ) ;
 assign wire14536 = ( n_n4474 ) | ( n_n4465 ) | ( wire14533 ) | ( wire14534 ) ;
 assign wire14537 = ( wire14440 ) | ( wire14441 ) | ( wire14444 ) | ( wire14445 ) ;
 assign wire14540 = ( n_n3653 ) | ( n_n3655 ) | ( wire14536 ) | ( wire14537 ) ;
 assign wire14542 = ( i_9_  &  n_n491  &  n_n520  &  n_n65 ) | ( (~ i_9_)  &  n_n491  &  n_n520  &  n_n65 ) ;
 assign wire14544 = ( n_n5279 ) | ( n_n5270 ) | ( n_n5280 ) ;
 assign wire14545 = ( wire438 ) | ( wire203 ) ;
 assign wire14549 = ( wire205 ) | ( wire409 ) ;
 assign wire14550 = ( n_n5267 ) | ( n_n5262 ) | ( wire77 ) | ( wire92 ) ;
 assign wire14551 = ( wire19  &  n_n473  &  n_n524 ) | ( wire19  &  n_n473  &  n_n528 ) ;
 assign wire14552 = ( wire11  &  n_n473  &  n_n65 ) | ( wire20  &  n_n473  &  n_n65 ) ;
 assign wire14554 = ( n_n5305 ) | ( n_n5306 ) | ( wire14551 ) ;
 assign wire14555 = ( wire459 ) | ( n_n5315 ) | ( wire14552 ) ;
 assign wire14557 = ( wire22  &  n_n464  &  n_n65 ) | ( wire11  &  n_n464  &  n_n65 ) ;
 assign wire14558 = ( wire19  &  n_n464  &  n_n530 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire14560 = ( n_n5318 ) | ( n_n5326 ) | ( wire14557 ) ;
 assign wire14561 = ( n_n5321 ) | ( n_n5328 ) | ( n_n5319 ) | ( wire14558 ) ;
 assign wire14563 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5292 ) ;
 assign wire14564 = ( n_n5303 ) | ( wire200 ) | ( n_n5304 ) ;
 assign wire14566 = ( n_n5302 ) | ( n_n5299 ) | ( wire14563 ) | ( wire14564 ) ;
 assign wire14567 = ( wire14554 ) | ( wire14555 ) | ( wire14560 ) | ( wire14561 ) ;
 assign wire14570 = ( wire21  &  n_n518  &  n_n65 ) | ( wire15  &  n_n518  &  n_n65 ) ;
 assign wire14572 = ( n_n5240 ) | ( n_n5238 ) | ( n_n5244 ) | ( n_n5233 ) ;
 assign wire14573 = ( n_n5241 ) | ( n_n5234 ) | ( n_n5242 ) | ( wire14570 ) ;
 assign wire14577 = ( n_n5228 ) | ( n_n5225 ) | ( wire62 ) ;
 assign wire14578 = ( wire434 ) | ( wire183 ) ;
 assign wire14579 = ( n_n5245 ) | ( n_n5254 ) | ( n_n5217 ) | ( n_n5248 ) ;
 assign wire14580 = ( wire318 ) | ( n_n5224 ) | ( n_n5227 ) | ( wire12874 ) ;
 assign wire14582 = ( wire14580 ) | ( wire14579 ) ;
 assign wire14583 = ( wire14572 ) | ( wire14573 ) | ( wire14577 ) | ( wire14578 ) ;
 assign wire14587 = ( n_n5284 ) | ( n_n5281 ) | ( n_n5288 ) | ( n_n5291 ) ;
 assign wire14588 = ( n_n5285 ) | ( n_n5289 ) | ( n_n5282 ) | ( wire14542 ) ;
 assign wire14589 = ( wire14588 ) | ( wire14587 ) ;
 assign wire14591 = ( n_n3664 ) | ( wire14549 ) | ( wire14550 ) | ( wire14589 ) ;
 assign wire14592 = ( wire14566 ) | ( wire14567 ) | ( wire14582 ) | ( wire14583 ) ;
 assign wire14594 = ( n_n5142 ) | ( wire76 ) | ( wire679 ) ;
 assign wire14595 = ( n_n5140 ) | ( n_n5144 ) | ( n_n5143 ) | ( wire12884 ) ;
 assign wire14598 = ( wire287 ) | ( wire406 ) ;
 assign wire14599 = ( n_n5155 ) | ( n_n5163 ) | ( n_n5154 ) | ( wire195 ) ;
 assign wire14601 = ( wire12  &  n_n509  &  n_n526 ) | ( wire12  &  n_n509  &  n_n530 ) ;
 assign wire14603 = ( wire22  &  n_n509  &  n_n130 ) | ( wire11  &  n_n509  &  n_n130 ) ;
 assign wire14605 = ( n_n5115 ) | ( n_n5118 ) | ( wire14601 ) ;
 assign wire14606 = ( n_n5122 ) | ( wire286 ) | ( wire14603 ) ;
 assign wire14609 = ( n_n5111 ) | ( n_n5112 ) | ( n_n5107 ) | ( n_n5108 ) ;
 assign wire14610 = ( n_n5113 ) | ( n_n5114 ) | ( n_n5106 ) | ( wire14001 ) ;
 assign wire14613 = ( n_n5133 ) | ( n_n3772 ) | ( wire12883 ) | ( wire14610 ) ;
 assign wire14614 = ( n_n3051 ) | ( wire14605 ) | ( wire14606 ) | ( wire14609 ) ;
 assign wire14615 = ( wire19  &  n_n526  &  n_n535 ) | ( wire19  &  n_n535  &  n_n528 ) ;
 assign wire14618 = ( n_n5201 ) | ( n_n5192 ) | ( wire761 ) ;
 assign wire14619 = ( n_n5200 ) | ( n_n5193 ) | ( wire452 ) ;
 assign wire14621 = ( wire22  &  n_n473  &  n_n130 ) | ( wire11  &  n_n473  &  n_n130 ) ;
 assign wire14622 = ( wire12  &  n_n522  &  n_n464 ) | ( wire12  &  n_n464  &  n_n520 ) ;
 assign wire14623 = ( n_n5191 ) | ( wire12  &  n_n522  &  n_n473 ) ;
 assign wire14624 = ( n_n5189 ) | ( n_n5190 ) | ( n_n5203 ) ;
 assign wire14625 = ( wire14622 ) | ( wire14621 ) ;
 assign wire14629 = ( n_n4129 ) | ( n_n1532 ) | ( n_n3037 ) | ( wire14623 ) ;
 assign wire14631 = ( wire21  &  n_n482  &  n_n130 ) | ( wire20  &  n_n482  &  n_n130 ) ;
 assign wire14635 = ( wire114 ) | ( n_n5175 ) | ( n_n5177 ) | ( n_n5170 ) ;
 assign wire14637 = ( wire14594 ) | ( wire14595 ) | ( wire14598 ) | ( wire14599 ) ;
 assign wire14638 = ( wire33 ) | ( wire14631 ) | ( wire14635 ) | ( wire14637 ) ;
 assign wire14641 = ( wire21  &  n_n464  &  n_n195 ) | ( wire23  &  n_n464  &  n_n195 ) ;
 assign wire14644 = ( n_n5081 ) | ( n_n5076 ) | ( wire14641 ) ;
 assign wire14645 = ( n_n5088 ) | ( n_n5078 ) | ( n_n5083 ) | ( wire123 ) ;
 assign wire14646 = ( wire22  &  n_n535  &  n_n130 ) | ( wire20  &  n_n535  &  n_n130 ) ;
 assign wire14648 = ( wire232 ) | ( wire122 ) ;
 assign wire14649 = ( n_n5098 ) | ( n_n5103 ) | ( n_n5095 ) | ( wire14646 ) ;
 assign wire14652 = ( n_n5060 ) | ( n_n5070 ) | ( wire160 ) ;
 assign wire14654 = ( n_n4152 ) | ( n_n5063 ) | ( n_n5058 ) | ( wire14652 ) ;
 assign wire14655 = ( wire14644 ) | ( wire14645 ) | ( wire14648 ) | ( wire14649 ) ;
 assign wire14656 = ( wire18  &  n_n473  &  n_n528 ) | ( wire18  &  n_n473  &  n_n532 ) ;
 assign wire14658 = ( n_n5055 ) | ( n_n5056 ) | ( n_n5051 ) ;
 assign wire14659 = ( n_n5048 ) | ( n_n5047 ) | ( wire14656 ) ;
 assign wire14661 = ( n_n5027 ) | ( n_n5028 ) | ( n_n5031 ) ;
 assign wire14662 = ( n_n5024 ) | ( wire253 ) | ( wire13400 ) ;
 assign wire14664 = ( n_n5043 ) | ( n_n5039 ) | ( n_n5044 ) ;
 assign wire14665 = ( n_n5025 ) | ( n_n5042 ) | ( wire97 ) ;
 assign wire14667 = ( n_n1570 ) | ( wire14664 ) | ( wire14665 ) ;
 assign wire14669 = ( i_9_  &  n_n500  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n532  &  n_n195 ) ;
 assign wire14671 = ( wire299 ) | ( wire136 ) ;
 assign wire14672 = ( wire103 ) | ( n_n5008 ) | ( wire14669 ) ;
 assign wire14673 = ( wire21  &  n_n509  &  n_n195 ) | ( wire23  &  n_n509  &  n_n195 ) ;
 assign wire14674 = ( n_n4998 ) | ( wire104 ) | ( wire743 ) ;
 assign wire14675 = ( n_n4989 ) | ( wire13997 ) | ( wire14673 ) ;
 assign wire14678 = ( wire21  &  n_n500  &  n_n195 ) | ( wire20  &  n_n500  &  n_n195 ) ;
 assign wire14680 = ( n_n5018 ) | ( n_n5017 ) | ( n_n5014 ) | ( n_n5020 ) ;
 assign wire14681 = ( n_n5021 ) | ( wire343 ) | ( wire14678 ) ;
 assign wire14683 = ( wire14671 ) | ( wire14672 ) | ( wire14674 ) | ( wire14675 ) ;
 assign wire14684 = ( wire14680 ) | ( wire14681 ) | ( wire14683 ) ;
 assign wire14689 = ( wire324 ) | ( wire295 ) ;
 assign wire14690 = ( n_n4862 ) | ( wire40 ) | ( n_n4867 ) | ( n_n4871 ) ;
 assign wire14691 = ( wire24  &  n_n518  &  n_n260 ) | ( wire15  &  n_n518  &  n_n260 ) ;
 assign wire14692 = ( wire17  &  n_n526  &  n_n518 ) | ( wire17  &  n_n532  &  n_n518 ) ;
 assign wire14694 = ( wire14691 ) | ( wire375 ) ;
 assign wire14695 = ( n_n4844 ) | ( wire52 ) | ( wire14692 ) ;
 assign wire14697 = ( n_n4830 ) | ( n_n4834 ) | ( n_n4833 ) | ( wire693 ) ;
 assign wire14701 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4808 ) ;
 assign wire14702 = ( n_n4816 ) | ( n_n4812 ) | ( n_n4804 ) | ( n_n4815 ) ;
 assign wire14706 = ( i_9_  &  n_n524  &  n_n464  &  n_n325 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n325 ) ;
 assign wire14708 = ( n_n4817 ) | ( n_n4828 ) | ( n_n4823 ) | ( n_n4820 ) ;
 assign wire14709 = ( n_n4821 ) | ( n_n4822 ) | ( n_n4826 ) | ( wire14706 ) ;
 assign wire14714 = ( n_n4801 ) | ( n_n4802 ) | ( wire380 ) ;
 assign wire14715 = ( n_n4791 ) | ( n_n4803 ) | ( wire179 ) | ( n_n4799 ) ;
 assign wire14717 = ( n_n4786 ) | ( wire11  &  n_n482  &  n_n325 ) ;
 assign wire14718 = ( wire313 ) | ( wire22  &  n_n482  &  n_n325 ) ;
 assign wire14719 = ( n_n4782 ) | ( n_n4779 ) | ( n_n4790 ) | ( n_n4781 ) ;
 assign wire14723 = ( wire14714 ) | ( wire14715 ) | ( wire14718 ) | ( wire14719 ) ;
 assign wire14724 = ( i_9_  &  n_n509  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n509  &  n_n534  &  n_n260 ) ;
 assign wire14725 = ( n_n4853 ) | ( wire17  &  n_n509  &  n_n532 ) ;
 assign wire14726 = ( wire14724 ) | ( wire102 ) ;
 assign wire14729 = ( wire14689 ) | ( wire14690 ) | ( wire14694 ) | ( wire14695 ) ;
 assign wire14730 = ( n_n2727 ) | ( wire14725 ) | ( wire14726 ) | ( wire14729 ) ;
 assign wire14733 = ( wire261 ) | ( wire264 ) ;
 assign wire14735 = ( wire11  &  n_n482  &  n_n260 ) | ( wire15  &  n_n482  &  n_n260 ) ;
 assign wire14738 = ( n_n4900 ) | ( n_n4903 ) | ( n_n4908 ) | ( n_n4899 ) ;
 assign wire14739 = ( n_n4905 ) | ( n_n4901 ) | ( n_n4910 ) | ( wire14735 ) ;
 assign wire14740 = ( wire21  &  n_n473  &  n_n260 ) | ( wire11  &  n_n473  &  n_n260 ) ;
 assign wire14742 = ( n_n4926 ) | ( n_n4925 ) | ( wire180 ) ;
 assign wire14743 = ( wire31 ) | ( n_n4932 ) | ( wire14740 ) ;
 assign wire14745 = ( wire17  &  n_n526  &  n_n482 ) | ( wire17  &  n_n520  &  n_n482 ) ;
 assign wire14747 = ( n_n4920 ) | ( n_n4919 ) | ( wire42 ) ;
 assign wire14748 = ( n_n4924 ) | ( n_n4947 ) | ( wire14745 ) ;
 assign wire14750 = ( n_n4917 ) | ( n_n4914 ) | ( wire14747 ) | ( wire14748 ) ;
 assign wire14751 = ( wire12168 ) | ( wire12169 ) | ( wire14742 ) | ( wire14743 ) ;
 assign wire14752 = ( i_9_  &  n_n535  &  n_n532  &  n_n195 ) | ( (~ i_9_)  &  n_n535  &  n_n532  &  n_n195 ) ;
 assign wire14754 = ( n_n4959 ) | ( n_n4962 ) | ( n_n4961 ) ;
 assign wire14756 = ( i_9_  &  n_n526  &  n_n518  &  n_n195 ) | ( (~ i_9_)  &  n_n526  &  n_n518  &  n_n195 ) ;
 assign wire14759 = ( wire18  &  n_n522  &  n_n518 ) | ( wire18  &  n_n524  &  n_n518 ) ;
 assign wire14760 = ( n_n4983 ) | ( n_n4984 ) | ( n_n4972 ) ;
 assign wire14761 = ( n_n4981 ) | ( n_n4987 ) | ( wire14756 ) ;
 assign wire14762 = ( n_n4985 ) | ( n_n4986 ) | ( wire14759 ) ;
 assign wire14764 = ( n_n4965 ) | ( wire13215 ) | ( wire13836 ) | ( wire14762 ) ;
 assign wire14766 = ( wire17  &  n_n526  &  n_n500 ) | ( wire17  &  n_n528  &  n_n500 ) ;
 assign wire14768 = ( n_n4882 ) | ( n_n4881 ) | ( wire14766 ) ;
 assign wire14770 = ( n_n4877 ) | ( n_n4884 ) | ( n_n3815 ) | ( wire14768 ) ;
 assign wire14772 = ( n_n3694 ) | ( wire14738 ) | ( wire14739 ) | ( wire14770 ) ;
 assign wire14774 = ( wire148 ) | ( wire149 ) | ( wire12963 ) ;
 assign wire14775 = ( n_n3648 ) | ( n_n3649 ) | ( wire14388 ) | ( wire14774 ) ;
 assign wire14777 = ( n_n3625 ) | ( n_n3645 ) | ( n_n3646 ) | ( wire14730 ) ;
 assign wire14778 = ( n_n3626 ) | ( wire14277 ) | ( wire14278 ) | ( wire14343 ) ;
 assign wire14779 = ( n_n3624 ) | ( wire14591 ) | ( wire14592 ) | ( wire14775 ) ;
 assign wire14782 = ( wire25  &  n_n509  &  n_n130 ) | ( wire25  &  n_n535  &  n_n130 ) ;
 assign wire14784 = ( n_n5131 ) | ( n_n5087 ) | ( n_n5132 ) | ( n_n5088 ) ;
 assign wire14785 = ( n_n5098 ) | ( n_n5104 ) | ( n_n5095 ) | ( wire14782 ) ;
 assign wire14790 = ( n_n5174 ) | ( n_n5184 ) | ( n_n5212 ) | ( n_n5172 ) ;
 assign wire14791 = ( n_n5234 ) | ( n_n5170 ) | ( n_n5148 ) | ( wire385 ) ;
 assign wire14795 = ( n_n5059 ) | ( wire231 ) | ( n_n5018 ) | ( n_n5045 ) ;
 assign wire14796 = ( n_n5048 ) | ( n_n5047 ) | ( wire97 ) | ( wire14795 ) ;
 assign wire14797 = ( wire14784 ) | ( wire14785 ) | ( wire14790 ) | ( wire14791 ) ;
 assign wire14801 = ( n_n5292 ) | ( wire21  &  n_n518  &  n_n65 ) ;
 assign wire14802 = ( n_n5284 ) | ( n_n5240 ) | ( n_n5248 ) ;
 assign wire14803 = ( n_n5245 ) | ( n_n5278 ) | ( n_n5287 ) | ( n_n5261 ) ;
 assign wire14807 = ( n_n5296 ) | ( n_n5320 ) | ( n_n5324 ) | ( n_n5335 ) ;
 assign wire14808 = ( wire11  &  n_n518  &  n_n195 ) | ( wire23  &  n_n518  &  n_n195 ) ;
 assign wire14810 = ( wire23  &  n_n535  &  n_n195 ) | ( wire23  &  n_n500  &  n_n195 ) ;
 assign wire14814 = ( n_n4985 ) | ( n_n4986 ) | ( n_n4962 ) | ( wire14808 ) ;
 assign wire14816 = ( wire17  &  n_n535  &  n_n530 ) | ( wire17  &  n_n530  &  n_n518 ) ;
 assign wire14817 = ( wire21  &  n_n491  &  n_n260 ) | ( wire22  &  n_n491  &  n_n260 ) ;
 assign wire14819 = ( n_n4847 ) | ( n_n4868 ) | ( n_n4871 ) ;
 assign wire14820 = ( wire14817 ) | ( wire14816 ) ;
 assign wire14825 = ( n_n4925 ) | ( n_n4907 ) | ( n_n4901 ) | ( n_n4904 ) ;
 assign wire14826 = ( n_n4913 ) | ( n_n4922 ) | ( n_n4934 ) | ( wire31 ) ;
 assign wire14829 = ( n_n2451 ) | ( wire14825 ) | ( wire14826 ) ;
 assign wire14830 = ( n_n2462 ) | ( n_n2464 ) | ( wire14796 ) | ( wire14797 ) ;
 assign wire14831 = ( wire10  &  n_n522  &  n_n500 ) | ( wire10  &  n_n500  &  n_n534 ) ;
 assign wire14833 = ( wire118 ) | ( n_n4631 ) | ( n_n4632 ) ;
 assign wire14834 = ( wire396 ) | ( n_n4629 ) | ( wire14831 ) ;
 assign wire14836 = ( wire13  &  n_n520  &  n_n518 ) | ( wire13  &  n_n530  &  n_n518 ) ;
 assign wire14838 = ( n_n4457 ) | ( n_n4475 ) | ( n_n4476 ) ;
 assign wire14839 = ( n_n4463 ) | ( n_n4494 ) | ( wire14836 ) ;
 assign wire14843 = ( wire24  &  n_n390  &  n_n518 ) | ( wire15  &  n_n390  &  n_n518 ) ;
 assign wire14845 = ( n_n4593 ) | ( n_n4571 ) | ( n_n4527 ) ;
 assign wire14846 = ( n_n4557 ) | ( n_n4533 ) | ( wire14843 ) ;
 assign wire14848 = ( n_n4592 ) | ( n_n4556 ) | ( wire14845 ) | ( wire14846 ) ;
 assign wire14854 = ( n_n4673 ) | ( n_n4690 ) | ( n_n4692 ) ;
 assign wire14855 = ( n_n4656 ) | ( n_n4697 ) | ( n_n4681 ) | ( n_n4660 ) ;
 assign wire14859 = ( wire24  &  n_n500  &  n_n325 ) | ( wire25  &  n_n500  &  n_n325 ) ;
 assign wire14861 = ( n_n4735 ) | ( n_n4724 ) | ( n_n4733 ) | ( n_n4725 ) ;
 assign wire14862 = ( n_n4760 ) | ( n_n4758 ) | ( n_n4714 ) | ( wire14859 ) ;
 assign wire14867 = ( n_n4790 ) | ( n_n4800 ) | ( n_n4826 ) ;
 assign wire14868 = ( n_n4803 ) | ( n_n4770 ) | ( n_n4772 ) | ( n_n4771 ) ;
 assign wire14870 = ( n_n4805 ) | ( n_n4766 ) | ( wire14867 ) | ( wire14868 ) ;
 assign wire14873 = ( wire21  &  n_n536  &  n_n500 ) | ( wire20  &  n_n536  &  n_n500 ) ;
 assign wire14875 = ( n_n4396 ) | ( n_n4375 ) | ( n_n4399 ) ;
 assign wire14876 = ( n_n4403 ) | ( n_n4382 ) | ( wire14873 ) ;
 assign wire14881 = ( n_n4352 ) | ( n_n4351 ) | ( n_n4330 ) ;
 assign wire14882 = ( n_n4318 ) | ( n_n4344 ) | ( n_n4320 ) | ( n_n4341 ) ;
 assign wire14886 = ( n_n4416 ) | ( n_n4448 ) | ( n_n4447 ) | ( n_n4415 ) ;
 assign wire14887 = ( n_n4453 ) | ( n_n4420 ) | ( n_n4407 ) | ( wire234 ) ;
 assign wire14890 = ( n_n2472 ) | ( n_n2473 ) | ( wire14886 ) | ( wire14887 ) ;
 assign wire14892 = ( n_n2455 ) | ( n_n2454 ) | ( wire14890 ) ;
 assign wire14894 = ( n_n4839 ) | ( n_n4840 ) | ( wire304 ) ;
 assign wire14896 = ( wire24  &  n_n535  &  n_n260 ) | ( wire25  &  n_n535  &  n_n260 ) ;
 assign wire14898 = ( n_n4830 ) | ( n_n4818 ) | ( wire693 ) ;
 assign wire14899 = ( n_n4821 ) | ( n_n4822 ) | ( wire14896 ) ;
 assign wire14903 = ( wire17  &  n_n526  &  n_n518 ) | ( wire17  &  n_n532  &  n_n518 ) ;
 assign wire14904 = ( n_n4856 ) | ( n_n4853 ) | ( n_n4858 ) | ( n_n4845 ) ;
 assign wire14905 = ( n_n4852 ) | ( wire11768 ) | ( wire14903 ) ;
 assign wire14909 = ( wire17  &  n_n500  &  n_n530 ) | ( wire17  &  n_n500  &  n_n532 ) ;
 assign wire14910 = ( n_n4880 ) | ( wire174 ) | ( n_n4879 ) ;
 assign wire14911 = ( n_n4882 ) | ( n_n4884 ) | ( n_n4883 ) | ( wire14909 ) ;
 assign wire14912 = ( wire49 ) | ( wire17  &  n_n528  &  n_n491 ) ;
 assign wire14914 = ( wire14  &  n_n522  &  n_n473 ) | ( wire14  &  n_n473  &  n_n528 ) ;
 assign wire14915 = ( wire24  &  n_n473  &  n_n325 ) | ( wire25  &  n_n473  &  n_n325 ) ;
 assign wire14917 = ( n_n4807 ) | ( n_n4808 ) | ( n_n4799 ) ;
 assign wire14918 = ( wire14915 ) | ( wire14914 ) ;
 assign wire14920 = ( wire14  &  n_n524  &  n_n482 ) | ( wire14  &  n_n528  &  n_n482 ) ;
 assign wire14922 = ( wire313 ) | ( wire131 ) ;
 assign wire14923 = ( n_n4784 ) | ( n_n4816 ) | ( n_n4783 ) | ( n_n4815 ) ;
 assign wire14924 = ( n_n4817 ) | ( n_n4792 ) | ( wire14920 ) ;
 assign wire14927 = ( wire85 ) | ( n_n4197 ) | ( wire12225 ) | ( wire14924 ) ;
 assign wire14931 = ( n_n4862 ) | ( n_n4870 ) | ( n_n4867 ) | ( n_n4872 ) ;
 assign wire14933 = ( n_n4866 ) | ( n_n4863 ) | ( n_n2727 ) | ( wire14931 ) ;
 assign wire14935 = ( n_n2597 ) | ( wire14910 ) | ( wire14911 ) | ( wire14933 ) ;
 assign wire14937 = ( wire22  &  n_n509  &  n_n195 ) | ( wire24  &  n_n509  &  n_n195 ) ;
 assign wire14938 = ( wire252 ) | ( wire134 ) ;
 assign wire14939 = ( n_n4996 ) | ( n_n4995 ) | ( n_n4994 ) | ( wire14937 ) ;
 assign wire14940 = ( i_9_  &  n_n500  &  n_n530  &  n_n195 ) | ( (~ i_9_)  &  n_n500  &  n_n530  &  n_n195 ) ;
 assign wire14942 = ( n_n4998 ) | ( wire393 ) | ( wire743 ) ;
 assign wire14943 = ( n_n5000 ) | ( wire136 ) | ( wire14940 ) ;
 assign wire14944 = ( wire11  &  n_n473  &  n_n260 ) | ( wire24  &  n_n473  &  n_n260 ) ;
 assign wire14946 = ( wire17  &  n_n473  &  n_n524 ) | ( wire17  &  n_n473  &  n_n528 ) ;
 assign wire14948 = ( n_n4924 ) | ( n_n4921 ) | ( wire14944 ) ;
 assign wire14949 = ( n_n4920 ) | ( n_n4919 ) | ( n_n4931 ) | ( wire14946 ) ;
 assign wire14954 = ( n_n4898 ) | ( n_n4903 ) | ( n_n4895 ) | ( n_n4908 ) ;
 assign wire14955 = ( wire96 ) | ( n_n4905 ) | ( n_n4906 ) | ( n_n4896 ) ;
 assign wire14956 = ( wire17  &  n_n522  &  n_n482 ) | ( wire17  &  n_n526  &  n_n482 ) ;
 assign wire14957 = ( i_9_  &  n_n524  &  n_n482  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n482  &  n_n260 ) ;
 assign wire14958 = ( n_n4918 ) | ( n_n4917 ) | ( wire14956 ) ;
 assign wire14960 = ( n_n4910 ) | ( wire14735 ) | ( wire14957 ) | ( wire14958 ) ;
 assign wire14961 = ( wire14948 ) | ( wire14949 ) | ( wire14954 ) | ( wire14955 ) ;
 assign wire14962 = ( i_9_  &  n_n524  &  n_n464  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n260 ) ;
 assign wire14964 = ( n_n4959 ) | ( n_n4960 ) | ( wire250 ) ;
 assign wire14965 = ( n_n4964 ) | ( n_n4957 ) | ( n_n4953 ) | ( wire14752 ) ;
 assign wire14967 = ( wire20  &  n_n464  &  n_n260 ) | ( wire25  &  n_n464  &  n_n260 ) ;
 assign wire14969 = ( wire382 ) | ( wire24  &  n_n464  &  n_n260 ) ;
 assign wire14970 = ( n_n4952 ) | ( n_n4950 ) | ( wire14967 ) ;
 assign wire14971 = ( n_n4936 ) | ( n_n4935 ) | ( n_n4948 ) | ( wire14962 ) ;
 assign wire14974 = ( n_n4944 ) | ( n_n2710 ) | ( wire13867 ) | ( wire14971 ) ;
 assign wire14975 = ( wire14964 ) | ( wire14965 ) | ( wire14969 ) | ( wire14970 ) ;
 assign wire14978 = ( n_n4978 ) | ( n_n4965 ) | ( n_n4973 ) | ( wire11809 ) ;
 assign wire14979 = ( wire228 ) | ( wire771 ) | ( wire772 ) | ( wire14978 ) ;
 assign wire14980 = ( wire14938 ) | ( wire14939 ) | ( wire14942 ) | ( wire14943 ) ;
 assign wire14982 = ( wire14960 ) | ( wire14961 ) | ( wire14974 ) | ( wire14975 ) ;
 assign wire14983 = ( wire22  &  n_n500  &  n_n325 ) | ( wire15  &  n_n500  &  n_n325 ) ;
 assign wire14985 = ( wire293 ) | ( wire47 ) ;
 assign wire14986 = ( wire109 ) | ( n_n4742 ) | ( wire14983 ) ;
 assign wire14987 = ( wire21  &  n_n500  &  n_n325 ) | ( wire23  &  n_n500  &  n_n325 ) ;
 assign wire14988 = ( wire11  &  n_n491  &  n_n325 ) | ( wire15  &  n_n491  &  n_n325 ) ;
 assign wire14990 = ( n_n4764 ) | ( n_n4763 ) | ( wire14987 ) ;
 assign wire14991 = ( wire164 ) | ( n_n4761 ) | ( wire14988 ) ;
 assign wire14992 = ( wire10  &  n_n473  &  n_n528 ) | ( wire10  &  n_n473  &  n_n532 ) ;
 assign wire14993 = ( wire10  &  n_n522  &  n_n473 ) | ( wire10  &  n_n473  &  n_n524 ) ;
 assign wire14995 = ( wire14992 ) | ( wire157 ) ;
 assign wire14996 = ( n_n4671 ) | ( wire80 ) | ( wire14993 ) ;
 assign wire14999 = ( n_n4695 ) | ( n_n4696 ) | ( n_n4694 ) ;
 assign wire15000 = ( n_n4685 ) | ( n_n4686 ) | ( wire417 ) ;
 assign wire15001 = ( wire442 ) | ( wire445 ) ;
 assign wire15002 = ( n_n4698 ) | ( n_n4688 ) | ( n_n4687 ) | ( n_n4680 ) ;
 assign wire15005 = ( n_n4222 ) | ( wire14999 ) | ( wire15002 ) ;
 assign wire15006 = ( wire14995 ) | ( wire14996 ) | ( wire15000 ) | ( wire15001 ) ;
 assign wire15007 = ( wire21  &  n_n535  &  n_n325 ) | ( wire23  &  n_n535  &  n_n325 ) ;
 assign wire15008 = ( n_n4705 ) | ( n_n4706 ) | ( wire15007 ) ;
 assign wire15010 = ( n_n4716 ) | ( wire25  &  n_n325  &  n_n518 ) ;
 assign wire15011 = ( n_n4737 ) | ( n_n4738 ) | ( n_n4723 ) ;
 assign wire15012 = ( n_n4712 ) | ( n_n4736 ) | ( n_n4722 ) | ( n_n4721 ) ;
 assign wire15016 = ( n_n4216 ) | ( wire243 ) | ( n_n856 ) | ( wire15010 ) ;
 assign wire15019 = ( n_n4778 ) | ( wire20  &  n_n491  &  n_n325 ) ;
 assign wire15020 = ( n_n4779 ) | ( n_n4775 ) | ( n_n4780 ) ;
 assign wire15021 = ( n_n4774 ) | ( n_n4781 ) | ( wire315 ) ;
 assign wire15024 = ( wire14985 ) | ( wire14986 ) | ( wire14990 ) | ( wire14991 ) ;
 assign wire15025 = ( wire15019 ) | ( wire15020 ) | ( wire15021 ) | ( wire15024 ) ;
 assign wire15028 = ( n_n4380 ) | ( n_n4367 ) | ( n_n4379 ) | ( n_n4368 ) ;
 assign wire15029 = ( n_n4384 ) | ( n_n4374 ) | ( wire423 ) | ( n_n4378 ) ;
 assign wire15032 = ( n_n4356 ) | ( n_n4355 ) | ( n_n4358 ) ;
 assign wire15033 = ( n_n4361 ) | ( n_n4363 ) | ( n_n4359 ) | ( n_n4364 ) ;
 assign wire15035 = ( wire22  &  n_n536  &  n_n491 ) | ( wire20  &  n_n536  &  n_n491 ) ;
 assign wire15037 = ( n_n4393 ) | ( n_n4395 ) | ( n_n4394 ) ;
 assign wire15038 = ( wire15035 ) | ( wire425 ) ;
 assign wire15040 = ( n_n4388 ) | ( n_n4392 ) | ( wire15037 ) | ( wire15038 ) ;
 assign wire15042 = ( wire21  &  n_n536  &  n_n473 ) | ( wire22  &  n_n536  &  n_n473 ) ;
 assign wire15043 = ( wire16  &  n_n473  &  n_n528 ) | ( wire16  &  n_n473  &  n_n532 ) ;
 assign wire15044 = ( n_n4411 ) | ( n_n4412 ) | ( wire15042 ) ;
 assign wire15045 = ( n_n4421 ) | ( wire215 ) | ( wire15043 ) ;
 assign wire15046 = ( i_9_  &  n_n536  &  n_n526  &  n_n482 ) | ( (~ i_9_)  &  n_n536  &  n_n526  &  n_n482 ) ;
 assign wire15048 = ( n_n4405 ) | ( n_n4406 ) | ( n_n4408 ) ;
 assign wire15049 = ( n_n4397 ) | ( n_n4398 ) | ( wire15046 ) ;
 assign wire15052 = ( wire16  &  n_n464  &  n_n528 ) | ( wire16  &  n_n464  &  n_n532 ) ;
 assign wire15053 = ( n_n4432 ) | ( n_n4431 ) | ( wire37 ) ;
 assign wire15055 = ( n_n4427 ) | ( wire14519 ) | ( wire15052 ) | ( wire15053 ) ;
 assign wire15057 = ( wire21  &  n_n473  &  n_n455 ) | ( wire24  &  n_n473  &  n_n455 ) ;
 assign wire15058 = ( wire13  &  n_n473  &  n_n526 ) | ( wire13  &  n_n473  &  n_n532 ) ;
 assign wire15059 = ( wire25  &  n_n473  &  n_n455 ) | ( wire15  &  n_n473  &  n_n455 ) ;
 assign wire15061 = ( wire15058 ) | ( wire15057 ) ;
 assign wire15062 = ( n_n4535 ) | ( n_n4536 ) | ( n_n4543 ) | ( wire15059 ) ;
 assign wire15063 = ( wire13  &  n_n532  &  n_n518 ) | ( wire13  &  n_n534  &  n_n518 ) ;
 assign wire15065 = ( wire291 ) | ( wire128 ) ;
 assign wire15066 = ( wire368 ) | ( n_n4446 ) | ( wire15063 ) ;
 assign wire15069 = ( n_n4464 ) | ( n_n4471 ) | ( n_n4472 ) | ( n_n4469 ) ;
 assign wire15071 = ( wire25  &  n_n455  &  n_n535 ) | ( wire15  &  n_n455  &  n_n535 ) ;
 assign wire15073 = ( wire15071 ) | ( wire236 ) ;
 assign wire15075 = ( n_n4439 ) | ( n_n4443 ) | ( n_n910 ) | ( wire15073 ) ;
 assign wire15077 = ( wire13  &  n_n524  &  n_n491 ) | ( wire13  &  n_n526  &  n_n491 ) ;
 assign wire15079 = ( n_n4515 ) | ( n_n4518 ) | ( wire791 ) ;
 assign wire15080 = ( n_n4520 ) | ( wire789 ) | ( wire15077 ) ;
 assign wire15082 = ( wire25  &  n_n509  &  n_n455 ) | ( wire15  &  n_n509  &  n_n455 ) ;
 assign wire15083 = ( wire13  &  n_n509  &  n_n522 ) | ( wire13  &  n_n509  &  n_n532 ) ;
 assign wire15084 = ( wire15082 ) | ( wire70 ) ;
 assign wire15085 = ( wire184 ) | ( wire787 ) | ( wire15083 ) ;
 assign wire15089 = ( n_n4489 ) | ( wire65 ) | ( n_n4490 ) ;
 assign wire15090 = ( n_n4497 ) | ( n_n4502 ) | ( wire347 ) ;
 assign wire15091 = ( n_n4492 ) | ( n_n4507 ) | ( n_n4505 ) | ( n_n4501 ) ;
 assign wire15094 = ( n_n4510 ) | ( n_n1677 ) | ( wire14200 ) | ( wire15091 ) ;
 assign wire15095 = ( wire15084 ) | ( wire15085 ) | ( wire15089 ) | ( wire15090 ) ;
 assign wire15097 = ( wire13  &  n_n522  &  n_n482 ) | ( wire13  &  n_n526  &  n_n482 ) ;
 assign wire15099 = ( n_n4526 ) | ( n_n4531 ) | ( n_n4529 ) | ( wire724 ) ;
 assign wire15101 = ( wire170 ) | ( n_n4534 ) | ( wire15097 ) | ( wire15099 ) ;
 assign wire15103 = ( n_n2626 ) | ( wire15061 ) | ( wire15062 ) | ( wire15101 ) ;
 assign wire15108 = ( n_n4602 ) | ( n_n4601 ) | ( wire45 ) ;
 assign wire15109 = ( wire108 ) | ( n_n4607 ) | ( n_n4600 ) | ( n_n4603 ) ;
 assign wire15111 = ( wire10  &  n_n528  &  n_n500 ) | ( wire10  &  n_n500  &  n_n530 ) ;
 assign wire15112 = ( n_n4617 ) | ( n_n4612 ) | ( n_n4611 ) | ( n_n4610 ) ;
 assign wire15113 = ( n_n4613 ) | ( wire465 ) | ( wire15111 ) ;
 assign wire15115 = ( wire10  &  n_n524  &  n_n518 ) | ( wire10  &  n_n532  &  n_n518 ) ;
 assign wire15117 = ( wire21  &  n_n390  &  n_n518 ) | ( wire11  &  n_n390  &  n_n518 ) ;
 assign wire15120 = ( n_n4597 ) | ( n_n4590 ) | ( n_n4585 ) | ( wire15117 ) ;
 assign wire15121 = ( n_n4583 ) | ( n_n4588 ) | ( wire15115 ) | ( wire15120 ) ;
 assign wire15122 = ( wire15108 ) | ( wire15109 ) | ( wire15112 ) | ( wire15113 ) ;
 assign wire15123 = ( wire10  &  n_n524  &  n_n535 ) | ( wire10  &  n_n535  &  n_n528 ) ;
 assign wire15125 = ( n_n4582 ) | ( n_n4581 ) | ( wire99 ) ;
 assign wire15126 = ( n_n4580 ) | ( wire238 ) | ( wire15123 ) ;
 assign wire15127 = ( wire24  &  n_n390  &  n_n482 ) | ( wire25  &  n_n390  &  n_n482 ) ;
 assign wire15130 = ( wire15127 ) | ( wire431 ) ;
 assign wire15131 = ( n_n4663 ) | ( n_n4652 ) | ( wire72 ) | ( n_n4657 ) ;
 assign wire15132 = ( wire10  &  n_n526  &  n_n491 ) | ( wire10  &  n_n528  &  n_n491 ) ;
 assign wire15133 = ( i_9_  &  n_n491  &  n_n390  &  n_n532 ) | ( (~ i_9_)  &  n_n491  &  n_n390  &  n_n532 ) ;
 assign wire15135 = ( wire26 ) | ( n_n4633 ) | ( n_n4630 ) ;
 assign wire15136 = ( wire190 ) | ( wire310 ) ;
 assign wire15137 = ( n_n4642 ) | ( n_n4623 ) | ( wire15133 ) ;
 assign wire15140 = ( n_n4639 ) | ( n_n2761 ) | ( wire15132 ) | ( wire15137 ) ;
 assign wire15141 = ( wire15130 ) | ( wire15131 ) | ( wire15135 ) | ( wire15136 ) ;
 assign wire15142 = ( i_9_  &  n_n464  &  n_n526  &  n_n455 ) | ( (~ i_9_)  &  n_n464  &  n_n526  &  n_n455 ) ;
 assign wire15143 = ( n_n4572 ) | ( wire24  &  n_n464  &  n_n455 ) ;
 assign wire15144 = ( wire212 ) | ( wire23  &  n_n473  &  n_n455 ) ;
 assign wire15145 = ( n_n4570 ) | ( n_n4569 ) | ( wire15142 ) ;
 assign wire15149 = ( wire15125 ) | ( wire15126 ) | ( wire15144 ) | ( wire15145 ) ;
 assign wire15150 = ( wire82 ) | ( wire224 ) | ( wire15143 ) | ( wire15149 ) ;
 assign wire15151 = ( wire15121 ) | ( wire15122 ) | ( wire15140 ) | ( wire15141 ) ;
 assign wire15153 = ( i_9_  &  n_n536  &  n_n528  &  n_n518 ) | ( (~ i_9_)  &  n_n536  &  n_n528  &  n_n518 ) ;
 assign wire15154 = ( n_n4336 ) | ( wire198 ) | ( n_n4329 ) ;
 assign wire15155 = ( n_n4337 ) | ( wire53 ) | ( wire15153 ) ;
 assign wire15159 = ( n_n4324 ) | ( n_n4319 ) | ( wire106 ) ;
 assign wire15160 = ( wire283 ) | ( n_n4321 ) | ( n_n4326 ) | ( n_n4322 ) ;
 assign wire15162 = ( n_n4348 ) | ( n_n4353 ) | ( n_n4354 ) ;
 assign wire15163 = ( n_n4345 ) | ( wire156 ) | ( wire675 ) ;
 assign wire15165 = ( n_n4340 ) | ( n_n4350 ) | ( wire15162 ) | ( wire15163 ) ;
 assign wire15166 = ( wire15154 ) | ( wire15155 ) | ( wire15159 ) | ( wire15160 ) ;
 assign wire15169 = ( n_n2560 ) | ( n_n2559 ) | ( wire15165 ) | ( wire15166 ) ;
 assign wire15174 = ( n_n5258 ) | ( n_n5255 ) | ( wire433 ) ;
 assign wire15175 = ( n_n5251 ) | ( n_n5254 ) | ( wire435 ) | ( n_n5253 ) ;
 assign wire15178 = ( n_n5244 ) | ( n_n5243 ) | ( wire320 ) ;
 assign wire15179 = ( n_n5238 ) | ( wire318 ) | ( n_n5249 ) | ( n_n5242 ) ;
 assign wire15180 = ( i_9_  &  n_n526  &  n_n500  &  n_n65 ) | ( (~ i_9_)  &  n_n526  &  n_n500  &  n_n65 ) ;
 assign wire15182 = ( n_n5262 ) | ( n_n5259 ) | ( wire334 ) ;
 assign wire15184 = ( n_n5270 ) | ( wire77 ) | ( wire15180 ) | ( wire15182 ) ;
 assign wire15185 = ( wire15174 ) | ( wire15175 ) | ( wire15178 ) | ( wire15179 ) ;
 assign wire15186 = ( wire19  &  n_n464  &  n_n526 ) | ( wire19  &  n_n464  &  n_n532 ) ;
 assign wire15188 = ( n_n5321 ) | ( wire149 ) | ( n_n5319 ) ;
 assign wire15189 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5327 ) | ( wire15186 ) ;
 assign wire15192 = ( wire148 ) | ( n_n3019 ) | ( n_n5312 ) | ( wire15189 ) ;
 assign wire15194 = ( n_n5297 ) | ( n_n5295 ) | ( n_n5298 ) ;
 assign wire15195 = ( n_n5303 ) | ( wire63 ) | ( n_n5304 ) ;
 assign wire15198 = ( wire438 ) | ( wire203 ) ;
 assign wire15200 = ( i_9_  &  n_n482  &  n_n532  &  n_n65 ) | ( (~ i_9_)  &  n_n482  &  n_n532  &  n_n65 ) ;
 assign wire15203 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5285 ) | ( wire15200 ) ;
 assign wire15204 = ( n_n5288 ) | ( n_n5286 ) | ( wire218 ) | ( wire15203 ) ;
 assign wire15206 = ( wire267 ) | ( wire15188 ) | ( wire15192 ) | ( wire15204 ) ;
 assign wire15207 = ( n_n2564 ) | ( n_n2566 ) | ( wire15184 ) | ( wire15185 ) ;
 assign wire15208 = ( wire19  &  n_n522  &  n_n518 ) | ( wire19  &  n_n528  &  n_n518 ) ;
 assign wire15211 = ( n_n5228 ) | ( n_n5225 ) | ( wire15208 ) ;
 assign wire15212 = ( n_n5229 ) | ( n_n5224 ) | ( wire87 ) | ( wire182 ) ;
 assign wire15216 = ( n_n5210 ) | ( wire220 ) | ( n_n5209 ) ;
 assign wire15217 = ( wire454 ) | ( wire384 ) ;
 assign wire15218 = ( n_n5206 ) | ( n_n5222 ) | ( n_n5214 ) | ( n_n5207 ) ;
 assign wire15219 = ( wire449 ) | ( n_n5219 ) | ( n_n5215 ) | ( wire14043 ) ;
 assign wire15221 = ( wire15219 ) | ( wire15218 ) ;
 assign wire15222 = ( wire15211 ) | ( wire15212 ) | ( wire15216 ) | ( wire15217 ) ;
 assign wire15223 = ( wire18  &  n_n522  &  n_n473 ) | ( wire18  &  n_n473  &  n_n532 ) ;
 assign wire15224 = ( wire22  &  n_n473  &  n_n195 ) | ( wire20  &  n_n473  &  n_n195 ) ;
 assign wire15226 = ( n_n5055 ) | ( n_n5056 ) | ( wire15223 ) ;
 assign wire15227 = ( wire166 ) | ( n_n5058 ) | ( wire15224 ) ;
 assign wire15230 = ( n_n5066 ) | ( wire123 ) | ( n_n5063 ) ;
 assign wire15231 = ( n_n5070 ) | ( n_n5082 ) | ( wire159 ) ;
 assign wire15234 = ( n_n4152 ) | ( n_n5065 ) | ( wire90 ) | ( n_n5090 ) ;
 assign wire15235 = ( wire15226 ) | ( wire15227 ) | ( wire15230 ) | ( wire15231 ) ;
 assign wire15239 = ( n_n5129 ) | ( n_n5124 ) | ( n_n5128 ) | ( n_n5122 ) ;
 assign wire15241 = ( wire21  &  n_n518  &  n_n130 ) | ( wire15  &  n_n518  &  n_n130 ) ;
 assign wire15243 = ( wire12  &  n_n524  &  n_n518 ) | ( wire12  &  n_n528  &  n_n518 ) ;
 assign wire15245 = ( n_n5096 ) | ( n_n5099 ) | ( wire15241 ) ;
 assign wire15246 = ( n_n5100 ) | ( n_n5103 ) | ( wire15243 ) ;
 assign wire15247 = ( n_n5091 ) | ( n_n5108 ) | ( wire88 ) | ( wire13305 ) ;
 assign wire15249 = ( wire335 ) | ( n_n5115 ) | ( wire11914 ) | ( wire15247 ) ;
 assign wire15252 = ( wire21  &  n_n482  &  n_n195 ) | ( wire15  &  n_n482  &  n_n195 ) ;
 assign wire15254 = ( n_n5036 ) | ( n_n5049 ) | ( wire253 ) ;
 assign wire15255 = ( wire356 ) | ( n_n5039 ) | ( wire15252 ) ;
 assign wire15257 = ( n_n5027 ) | ( n_n5028 ) | ( wire265 ) ;
 assign wire15258 = ( n_n5026 ) | ( wire50 ) | ( n_n5023 ) | ( n_n5029 ) ;
 assign wire15261 = ( n_n5022 ) | ( n_n5011 ) | ( n_n5013 ) | ( wire12931 ) ;
 assign wire15263 = ( wire15254 ) | ( wire15255 ) | ( wire15257 ) | ( wire15258 ) ;
 assign wire15264 = ( wire297 ) | ( wire394 ) | ( wire15261 ) | ( wire15263 ) ;
 assign wire15266 = ( wire22  &  n_n473  &  n_n130 ) | ( wire15  &  n_n473  &  n_n130 ) ;
 assign wire15269 = ( n_n5191 ) | ( n_n5192 ) | ( wire15266 ) ;
 assign wire15270 = ( wire112 ) | ( n_n5193 ) | ( n_n5182 ) | ( n_n5190 ) ;
 assign wire15273 = ( n_n5201 ) | ( wire437 ) | ( wire761 ) ;
 assign wire15274 = ( n_n5175 ) | ( n_n5177 ) | ( wire451 ) ;
 assign wire15275 = ( n_n5173 ) | ( n_n5203 ) | ( n_n5197 ) | ( n_n5176 ) ;
 assign wire15278 = ( wire114 ) | ( n_n2670 ) | ( wire765 ) | ( wire15275 ) ;
 assign wire15279 = ( wire15269 ) | ( wire15270 ) | ( wire15273 ) | ( wire15274 ) ;
 assign wire15280 = ( wire12  &  n_n530  &  n_n482 ) | ( wire12  &  n_n482  &  n_n532 ) ;
 assign wire15283 = ( wire15280 ) | ( wire254 ) ;
 assign wire15284 = ( n_n5163 ) | ( n_n5157 ) | ( wire195 ) | ( n_n5160 ) ;
 assign wire15285 = ( wire21  &  n_n491  &  n_n130 ) | ( wire25  &  n_n491  &  n_n130 ) ;
 assign wire15287 = ( wire407 ) | ( wire288 ) ;
 assign wire15288 = ( wire196 ) | ( n_n5149 ) | ( wire15285 ) ;
 assign wire15289 = ( wire22  &  n_n500  &  n_n130 ) | ( wire11  &  n_n500  &  n_n130 ) ;
 assign wire15290 = ( i_9_  &  n_n524  &  n_n500  &  n_n130 ) | ( (~ i_9_)  &  n_n524  &  n_n500  &  n_n130 ) ;
 assign wire15291 = ( wire15289 ) | ( wire211 ) ;
 assign wire15292 = ( n_n5130 ) | ( n_n5133 ) | ( n_n5134 ) | ( wire15290 ) ;
 assign wire15294 = ( wire15283 ) | ( wire15284 ) | ( wire15287 ) | ( wire15288 ) ;
 assign wire15296 = ( wire15221 ) | ( wire15222 ) | ( wire15278 ) | ( wire15279 ) ;
 assign wire15297 = ( wire15291 ) | ( wire15292 ) | ( wire15294 ) | ( wire15296 ) ;
 assign wire15299 = ( n_n2530 ) | ( wire14979 ) | ( wire14980 ) | ( wire14982 ) ;
 assign wire15300 = ( n_n2531 ) | ( wire14829 ) | ( wire14830 ) | ( wire14892 ) ;
 assign wire15304 = ( wire23  &  n_n509  &  n_n536 ) | ( wire23  &  n_n536  &  n_n491 ) ;
 assign wire15307 = ( n_n4371 ) | ( n_n4431 ) | ( n_n4424 ) ;
 assign wire15308 = ( n_n4384 ) | ( n_n4397 ) | ( wire15304 ) ;
 assign wire15310 = ( wire21  &  n_n455  &  n_n535 ) | ( wire20  &  n_n455  &  n_n535 ) ;
 assign wire15312 = ( wire13  &  n_n532  &  n_n518 ) | ( wire13  &  n_n534  &  n_n518 ) ;
 assign wire15315 = ( n_n4487 ) | ( n_n4478 ) | ( wire15312 ) ;
 assign wire15316 = ( n_n4457 ) | ( n_n4488 ) | ( n_n4476 ) | ( wire15310 ) ;
 assign wire15321 = ( n_n4345 ) | ( n_n4319 ) | ( n_n4316 ) ;
 assign wire15322 = ( n_n4320 ) | ( n_n4315 ) | ( n_n4348 ) | ( n_n4357 ) ;
 assign wire15326 = ( wire10  &  n_n509  &  n_n528 ) | ( wire10  &  n_n509  &  n_n534 ) ;
 assign wire15328 = ( n_n4598 ) | ( n_n4570 ) | ( n_n4612 ) | ( n_n4572 ) ;
 assign wire15329 = ( n_n4609 ) | ( wire401 ) | ( wire15326 ) ;
 assign wire15333 = ( n_n4634 ) | ( n_n4687 ) | ( n_n4631 ) ;
 assign wire15334 = ( n_n4659 ) | ( wire75 ) | ( n_n4689 ) | ( n_n4698 ) ;
 assign wire15340 = ( n_n4514 ) | ( n_n4511 ) | ( n_n4525 ) | ( n_n4528 ) ;
 assign wire15341 = ( wire416 ) | ( n_n4527 ) | ( n_n4534 ) | ( n_n4552 ) ;
 assign wire15342 = ( wire15341 ) | ( wire15340 ) ;
 assign wire15348 = ( n_n4898 ) | ( n_n4877 ) | ( n_n4876 ) | ( n_n4899 ) ;
 assign wire15349 = ( n_n4886 ) | ( n_n4915 ) | ( wire154 ) | ( n_n4874 ) ;
 assign wire15354 = ( n_n5111 ) | ( n_n5113 ) | ( n_n5143 ) ;
 assign wire15355 = ( n_n5161 ) | ( n_n5120 ) | ( n_n5135 ) | ( n_n5147 ) ;
 assign wire15360 = ( n_n5064 ) | ( n_n5001 ) | ( wire755 ) ;
 assign wire15361 = ( n_n4990 ) | ( n_n5027 ) | ( n_n5048 ) | ( n_n5053 ) ;
 assign wire15367 = ( n_n5092 ) | ( n_n5069 ) | ( n_n5084 ) | ( n_n5078 ) ;
 assign wire15368 = ( n_n5068 ) | ( n_n5090 ) | ( n_n5080 ) | ( wire279 ) ;
 assign wire15374 = ( n_n5230 ) | ( n_n5168 ) | ( wire107 ) ;
 assign wire15375 = ( n_n5169 ) | ( wire33 ) | ( n_n5235 ) | ( n_n5217 ) ;
 assign wire15376 = ( wire22  &  n_n464  &  n_n65 ) | ( wire15  &  n_n464  &  n_n65 ) ;
 assign wire15382 = ( n_n5302 ) | ( n_n5273 ) | ( n_n5327 ) | ( n_n5254 ) ;
 assign wire15383 = ( n_n5278 ) | ( n_n5319 ) | ( wire200 ) | ( n_n5282 ) ;
 assign wire15385 = ( wire386 ) | ( wire15376 ) | ( wire15382 ) | ( wire15383 ) ;
 assign wire15389 = ( n_n4959 ) | ( n_n4960 ) | ( n_n4961 ) ;
 assign wire15390 = ( n_n4963 ) | ( n_n4964 ) | ( n_n4974 ) | ( n_n4967 ) ;
 assign wire15396 = ( n_n4921 ) | ( n_n4938 ) | ( n_n4936 ) | ( n_n4917 ) ;
 assign wire15397 = ( n_n4931 ) | ( n_n4948 ) | ( n_n4957 ) | ( wire141 ) ;
 assign wire15398 = ( wire15397 ) | ( wire15396 ) ;
 assign wire15400 = ( wire15374 ) | ( wire15375 ) | ( wire15385 ) | ( wire15398 ) ;
 assign wire15405 = ( n_n4757 ) | ( n_n4760 ) | ( n_n4815 ) ;
 assign wire15406 = ( n_n4769 ) | ( n_n4794 ) | ( n_n4797 ) | ( n_n4788 ) ;
 assign wire15412 = ( n_n4854 ) | ( n_n4843 ) | ( wire150 ) ;
 assign wire15413 = ( wire40 ) | ( n_n4852 ) | ( n_n4826 ) | ( n_n4872 ) ;
 assign wire15416 = ( n_n4711 ) | ( n_n4732 ) | ( n_n4729 ) | ( wire767 ) ;
 assign wire15418 = ( n_n4718 ) | ( n_n4700 ) | ( n_n1760 ) | ( wire15416 ) ;
 assign wire15421 = ( wire24  &  n_n509  &  n_n455 ) | ( wire15  &  n_n509  &  n_n455 ) ;
 assign wire15423 = ( n_n4472 ) | ( n_n4469 ) | ( wire15421 ) ;
 assign wire15426 = ( n_n4448 ) | ( n_n4447 ) | ( wire421 ) ;
 assign wire15428 = ( i_9_  &  n_n455  &  n_n528  &  n_n500 ) | ( (~ i_9_)  &  n_n455  &  n_n528  &  n_n500 ) ;
 assign wire15431 = ( n_n4491 ) | ( n_n4492 ) | ( wire15428 ) ;
 assign wire15432 = ( n_n4497 ) | ( wire65 ) | ( n_n4500 ) | ( n_n4496 ) ;
 assign wire15434 = ( n_n4506 ) | ( n_n4505 ) | ( n_n4490 ) ;
 assign wire15435 = ( n_n4504 ) | ( n_n4502 ) | ( n_n4507 ) | ( n_n4501 ) ;
 assign wire15437 = ( n_n4510 ) | ( wire14200 ) | ( wire15434 ) | ( wire15435 ) ;
 assign wire15438 = ( wire11511 ) | ( wire11512 ) | ( wire15431 ) | ( wire15432 ) ;
 assign wire15440 = ( wire129 ) | ( wire170 ) ;
 assign wire15444 = ( n_n4535 ) | ( n_n4536 ) | ( n_n4529 ) ;
 assign wire15445 = ( n_n4526 ) | ( n_n4533 ) | ( wire379 ) ;
 assign wire15448 = ( wire13  &  n_n473  &  n_n524 ) | ( wire13  &  n_n473  &  n_n532 ) ;
 assign wire15451 = ( n_n4547 ) | ( n_n4544 ) | ( wire15448 ) ;
 assign wire15452 = ( n_n4545 ) | ( n_n4550 ) | ( wire201 ) | ( n_n4549 ) ;
 assign wire15456 = ( wire13  &  n_n522  &  n_n535 ) | ( wire13  &  n_n524  &  n_n535 ) ;
 assign wire15459 = ( n_n4463 ) | ( n_n4455 ) | ( wire15456 ) ;
 assign wire15460 = ( n_n4454 ) | ( n_n4465 ) | ( n_n4462 ) | ( wire291 ) ;
 assign wire15463 = ( n_n3001 ) | ( n_n3003 ) | ( wire15459 ) | ( wire15460 ) ;
 assign wire15467 = ( wire157 ) | ( wire309 ) ;
 assign wire15468 = ( n_n4666 ) | ( n_n4648 ) | ( wire139 ) ;
 assign wire15469 = ( n_n4644 ) | ( n_n4658 ) | ( n_n4642 ) | ( wire13454 ) ;
 assign wire15471 = ( n_n4663 ) | ( wire225 ) | ( wire11856 ) | ( wire15469 ) ;
 assign wire15472 = ( wire13887 ) | ( wire13888 ) | ( wire15467 ) | ( wire15468 ) ;
 assign wire15474 = ( n_n4568 ) | ( wire276 ) | ( wire783 ) ;
 assign wire15475 = ( n_n4574 ) | ( n_n4573 ) | ( wire455 ) | ( wire671 ) ;
 assign wire15478 = ( n_n4582 ) | ( n_n4584 ) | ( n_n4581 ) | ( n_n4583 ) ;
 assign wire15479 = ( n_n4587 ) | ( wire365 ) | ( n_n4580 ) | ( n_n4585 ) ;
 assign wire15481 = ( wire10  &  n_n500  &  n_n530 ) | ( wire10  &  n_n500  &  n_n532 ) ;
 assign wire15482 = ( n_n4617 ) | ( n_n4613 ) | ( n_n4607 ) | ( n_n4610 ) ;
 assign wire15483 = ( n_n4616 ) | ( wire465 ) | ( wire15481 ) ;
 assign wire15485 = ( wire10  &  n_n524  &  n_n518 ) | ( wire10  &  n_n528  &  n_n518 ) ;
 assign wire15488 = ( n_n4593 ) | ( n_n4601 ) | ( wire15485 ) ;
 assign wire15489 = ( wire108 ) | ( n_n4603 ) | ( n_n4595 ) | ( n_n4592 ) ;
 assign wire15490 = ( i_9_  &  n_n522  &  n_n500  &  n_n390 ) | ( (~ i_9_)  &  n_n522  &  n_n500  &  n_n390 ) ;
 assign wire15493 = ( n_n4639 ) | ( n_n4621 ) | ( n_n4632 ) | ( wire12547 ) ;
 assign wire15494 = ( wire190 ) | ( wire15490 ) | ( wire15493 ) ;
 assign wire15495 = ( wire15482 ) | ( wire15483 ) | ( wire15488 ) | ( wire15489 ) ;
 assign wire15498 = ( n_n4557 ) | ( n_n4558 ) | ( n_n4559 ) ;
 assign wire15499 = ( n_n4560 ) | ( n_n4553 ) | ( wire430 ) ;
 assign wire15501 = ( n_n4561 ) | ( n_n4556 ) | ( wire15498 ) | ( wire15499 ) ;
 assign wire15502 = ( wire15474 ) | ( wire15475 ) | ( wire15478 ) | ( wire15479 ) ;
 assign wire15504 = ( wire15471 ) | ( wire15472 ) | ( wire15494 ) | ( wire15495 ) ;
 assign wire15506 = ( n_n4393 ) | ( n_n4396 ) | ( n_n4399 ) ;
 assign wire15507 = ( n_n4389 ) | ( n_n4390 ) | ( wire420 ) ;
 assign wire15509 = ( wire16  &  n_n528  &  n_n500 ) | ( wire16  &  n_n500  &  n_n532 ) ;
 assign wire15511 = ( n_n4353 ) | ( n_n4358 ) | ( n_n4354 ) ;
 assign wire15512 = ( n_n4367 ) | ( n_n4368 ) | ( wire15509 ) ;
 assign wire15517 = ( n_n4344 ) | ( n_n4342 ) | ( wire124 ) ;
 assign wire15518 = ( n_n4352 ) | ( wire67 ) | ( n_n4349 ) | ( n_n4350 ) ;
 assign wire15521 = ( n_n4325 ) | ( n_n4314 ) | ( n_n4328 ) ;
 assign wire15525 = ( n_n4336 ) | ( n_n4331 ) | ( n_n4334 ) | ( wire677 ) ;
 assign wire15526 = ( n_n4337 ) | ( n_n4332 ) | ( n_n4329 ) | ( wire53 ) ;
 assign wire15527 = ( wire15526 ) | ( wire15525 ) ;
 assign wire15529 = ( wire16  &  n_n524  &  n_n464 ) | ( wire16  &  n_n464  &  n_n526 ) ;
 assign wire15532 = ( n_n4430 ) | ( n_n4429 ) | ( wire15529 ) ;
 assign wire15533 = ( n_n4433 ) | ( n_n4438 ) | ( n_n4425 ) | ( wire84 ) ;
 assign wire15534 = ( wire16  &  n_n522  &  n_n473 ) | ( wire16  &  n_n473  &  n_n526 ) ;
 assign wire15536 = ( wire79 ) | ( wire215 ) ;
 assign wire15537 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) | ( wire15534 ) ;
 assign wire15538 = ( wire21  &  n_n536  &  n_n482 ) | ( wire23  &  n_n536  &  n_n482 ) ;
 assign wire15539 = ( wire16  &  n_n522  &  n_n482 ) | ( wire16  &  n_n520  &  n_n482 ) ;
 assign wire15542 = ( n_n4401 ) | ( n_n4408 ) | ( n_n4402 ) | ( wire15539 ) ;
 assign wire15543 = ( n_n4409 ) | ( n_n4410 ) | ( wire15538 ) | ( wire15542 ) ;
 assign wire15544 = ( wire15532 ) | ( wire15533 ) | ( wire15536 ) | ( wire15537 ) ;
 assign wire15545 = ( n_n4369 ) | ( n_n4373 ) | ( n_n4374 ) ;
 assign wire15546 = ( n_n4381 ) | ( wire423 ) | ( n_n4378 ) | ( wire12449 ) ;
 assign wire15549 = ( n_n3007 ) | ( n_n3009 ) | ( wire15545 ) | ( wire15546 ) ;
 assign wire15551 = ( wire12  &  n_n464  &  n_n526 ) | ( wire12  &  n_n464  &  n_n520 ) ;
 assign wire15554 = ( n_n5207 ) | ( n_n5208 ) | ( wire15551 ) ;
 assign wire15555 = ( n_n5199 ) | ( wire220 ) | ( n_n5209 ) | ( wire636 ) ;
 assign wire15557 = ( wire19  &  n_n522  &  n_n535 ) | ( wire19  &  n_n535  &  n_n532 ) ;
 assign wire15559 = ( n_n5191 ) | ( wire454 ) | ( n_n5192 ) ;
 assign wire15560 = ( wire453 ) | ( wire183 ) ;
 assign wire15562 = ( wire112 ) | ( n_n5215 ) | ( n_n5198 ) | ( wire14615 ) ;
 assign wire15564 = ( n_n5183 ) | ( n_n5188 ) | ( wire15557 ) | ( wire15562 ) ;
 assign wire15565 = ( wire15554 ) | ( wire15555 ) | ( wire15559 ) | ( wire15560 ) ;
 assign wire15569 = ( n_n5223 ) | ( n_n5229 ) | ( wire182 ) ;
 assign wire15570 = ( n_n5228 ) | ( n_n5225 ) | ( n_n5224 ) | ( wire385 ) ;
 assign wire15573 = ( n_n5239 ) | ( n_n5240 ) | ( n_n5244 ) | ( n_n5243 ) ;
 assign wire15574 = ( wire446 ) | ( wire62 ) ;
 assign wire15575 = ( n_n5241 ) | ( n_n5262 ) | ( n_n5234 ) | ( n_n5246 ) ;
 assign wire15576 = ( n_n5255 ) | ( n_n5251 ) | ( wire435 ) | ( wire433 ) ;
 assign wire15578 = ( wire15576 ) | ( wire15575 ) ;
 assign wire15579 = ( wire15569 ) | ( wire15570 ) | ( wire15573 ) | ( wire15574 ) ;
 assign wire15582 = ( wire11  &  n_n482  &  n_n130 ) | ( wire24  &  n_n482  &  n_n130 ) ;
 assign wire15583 = ( wire15582 ) | ( wire12  &  n_n522  &  n_n482 ) ;
 assign wire15586 = ( n_n5142 ) | ( wire196 ) | ( wire679 ) ;
 assign wire15587 = ( n_n5146 ) | ( wire76 ) | ( n_n5139 ) | ( n_n5151 ) ;
 assign wire15589 = ( i_9_  &  n_n473  &  n_n534  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n534  &  n_n130 ) ;
 assign wire15590 = ( n_n5179 ) | ( n_n5173 ) | ( wire44 ) ;
 assign wire15591 = ( n_n5181 ) | ( n_n5182 ) | ( wire732 ) | ( wire15589 ) ;
 assign wire15593 = ( wire466 ) | ( wire15583 ) | ( wire15586 ) | ( wire15587 ) ;
 assign wire15594 = ( wire15590 ) | ( wire15591 ) | ( wire15593 ) ;
 assign wire15595 = ( wire15564 ) | ( wire15565 ) | ( wire15578 ) | ( wire15579 ) ;
 assign wire15596 = ( wire20  &  n_n482  &  n_n195 ) | ( wire15  &  n_n482  &  n_n195 ) ;
 assign wire15597 = ( n_n5043 ) | ( n_n5044 ) | ( wire15596 ) ;
 assign wire15598 = ( wire18  &  n_n473  &  n_n528 ) | ( wire18  &  n_n473  &  n_n532 ) ;
 assign wire15601 = ( n_n5055 ) | ( n_n5056 ) | ( n_n5052 ) ;
 assign wire15602 = ( n_n5049 ) | ( n_n5046 ) | ( wire15598 ) ;
 assign wire15605 = ( n_n5089 ) | ( n_n5098 ) | ( n_n5095 ) ;
 assign wire15606 = ( n_n5087 ) | ( n_n5088 ) | ( wire122 ) ;
 assign wire15609 = ( n_n5057 ) | ( n_n5058 ) | ( n_n5065 ) ;
 assign wire15610 = ( n_n5066 ) | ( n_n5063 ) | ( wire159 ) ;
 assign wire15612 = ( wire25  &  n_n535  &  n_n130 ) | ( wire15  &  n_n535  &  n_n130 ) ;
 assign wire15614 = ( i_9_  &  n_n524  &  n_n464  &  n_n195 ) | ( (~ i_9_)  &  n_n524  &  n_n464  &  n_n195 ) ;
 assign wire15616 = ( n_n5086 ) | ( n_n5073 ) | ( wire15612 ) ;
 assign wire15617 = ( n_n5079 ) | ( wire209 ) | ( wire15614 ) ;
 assign wire15620 = ( wire11  &  n_n518  &  n_n130 ) | ( wire20  &  n_n518  &  n_n130 ) ;
 assign wire15621 = ( wire12  &  n_n526  &  n_n518 ) | ( wire12  &  n_n528  &  n_n518 ) ;
 assign wire15623 = ( n_n5112 ) | ( n_n5110 ) | ( wire15620 ) ;
 assign wire15624 = ( n_n5107 ) | ( n_n5106 ) | ( n_n5108 ) | ( wire15621 ) ;
 assign wire15626 = ( wire11  &  n_n509  &  n_n130 ) | ( wire24  &  n_n509  &  n_n130 ) ;
 assign wire15627 = ( wire12  &  n_n524  &  n_n500 ) | ( wire12  &  n_n528  &  n_n500 ) ;
 assign wire15628 = ( wire335 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire15629 = ( n_n5136 ) | ( n_n5124 ) | ( wire286 ) ;
 assign wire15633 = ( n_n3772 ) | ( n_n3051 ) | ( wire15626 ) | ( wire15627 ) ;
 assign wire15634 = ( wire15623 ) | ( wire15624 ) | ( wire15628 ) | ( wire15629 ) ;
 assign wire15639 = ( n_n5036 ) | ( wire231 ) | ( n_n5031 ) | ( n_n5029 ) ;
 assign wire15640 = ( n_n5032 ) | ( n_n5028 ) | ( wire265 ) | ( wire15639 ) ;
 assign wire15642 = ( wire230 ) | ( n_n2956 ) | ( wire15597 ) | ( wire15640 ) ;
 assign wire15647 = ( n_n5322 ) | ( wire20  &  n_n473  &  n_n65 ) ;
 assign wire15648 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5315 ) ;
 assign wire15649 = ( n_n5321 ) | ( n_n5326 ) | ( n_n5323 ) | ( n_n5324 ) ;
 assign wire15651 = ( wire19  &  n_n522  &  n_n491 ) | ( wire19  &  n_n491  &  n_n530 ) ;
 assign wire15653 = ( n_n5279 ) | ( n_n5283 ) | ( n_n5280 ) ;
 assign wire15654 = ( wire15651 ) | ( wire333 ) ;
 assign wire15658 = ( n_n5270 ) | ( n_n5269 ) | ( wire205 ) ;
 assign wire15659 = ( n_n5268 ) | ( n_n5271 ) | ( wire334 ) | ( wire92 ) ;
 assign wire15660 = ( wire19  &  n_n473  &  n_n524 ) | ( wire19  &  n_n473  &  n_n528 ) ;
 assign wire15663 = ( n_n5300 ) | ( n_n5299 ) | ( wire15660 ) ;
 assign wire15665 = ( n_n5295 ) | ( wire20  &  n_n491  &  n_n65 ) ;
 assign wire15666 = ( n_n5291 ) | ( n_n5292 ) | ( n_n5289 ) ;
 assign wire15667 = ( n_n5293 ) | ( n_n5294 ) | ( n_n5288 ) | ( n_n5286 ) ;
 assign wire15671 = ( n_n5328 ) | ( n_n5335 ) | ( wire149 ) | ( n_n5331 ) ;
 assign wire15672 = ( wire15647 ) | ( wire15648 ) | ( wire15649 ) | ( wire15671 ) ;
 assign wire15674 = ( n_n2937 ) | ( wire15665 ) | ( wire15666 ) | ( wire15667 ) ;
 assign wire15675 = ( n_n2939 ) | ( wire15658 ) | ( wire15659 ) | ( wire15672 ) ;
 assign wire15677 = ( wire15594 ) | ( wire15595 ) | ( wire15674 ) | ( wire15675 ) ;
 assign wire15678 = ( wire17  &  n_n509  &  n_n526 ) | ( wire17  &  n_n509  &  n_n530 ) ;
 assign wire15680 = ( n_n4862 ) | ( n_n4869 ) | ( n_n4861 ) | ( n_n4870 ) ;
 assign wire15681 = ( wire245 ) | ( n_n4868 ) | ( wire15678 ) ;
 assign wire15683 = ( wire49 ) | ( wire96 ) ;
 assign wire15684 = ( n_n4903 ) | ( n_n4896 ) | ( n_n4889 ) | ( wire12179 ) ;
 assign wire15685 = ( n_n4828 ) | ( wire20  &  n_n464  &  n_n325 ) ;
 assign wire15686 = ( n_n4830 ) | ( n_n4827 ) | ( n_n4824 ) | ( wire693 ) ;
 assign wire15688 = ( i_9_  &  n_n509  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n509  &  n_n534  &  n_n260 ) ;
 assign wire15689 = ( wire22  &  n_n518  &  n_n260 ) | ( wire20  &  n_n518  &  n_n260 ) ;
 assign wire15693 = ( n_n4855 ) | ( n_n4842 ) | ( wire15689 ) ;
 assign wire15695 = ( wire176 ) | ( wire52 ) | ( wire375 ) | ( wire15688 ) ;
 assign wire15696 = ( n_n3820 ) | ( n_n4836 ) | ( wire11769 ) | ( wire15693 ) ;
 assign wire15697 = ( n_n3461 ) | ( wire15685 ) | ( wire15686 ) | ( wire15695 ) ;
 assign wire15698 = ( wire17  &  n_n473  &  n_n526 ) | ( wire17  &  n_n473  &  n_n532 ) ;
 assign wire15700 = ( n_n4920 ) | ( n_n4926 ) | ( n_n4925 ) | ( n_n4919 ) ;
 assign wire15701 = ( n_n4930 ) | ( wire382 ) | ( wire15698 ) ;
 assign wire15702 = ( wire18  &  n_n528  &  n_n491 ) | ( wire18  &  n_n491  &  n_n532 ) ;
 assign wire15704 = ( wire296 ) | ( n_n5019 ) | ( n_n5020 ) ;
 assign wire15705 = ( n_n5017 ) | ( wire135 ) | ( wire15702 ) ;
 assign wire15707 = ( wire18  &  n_n500  &  n_n530 ) | ( wire18  &  n_n500  &  n_n534 ) ;
 assign wire15709 = ( n_n4998 ) | ( wire136 ) | ( wire743 ) ;
 assign wire15710 = ( wire104 ) | ( wire394 ) ;
 assign wire15712 = ( n_n5003 ) | ( n_n4994 ) | ( wire12255 ) | ( wire12256 ) ;
 assign wire15714 = ( n_n4996 ) | ( n_n4999 ) | ( wire15707 ) | ( wire15712 ) ;
 assign wire15715 = ( wire15704 ) | ( wire15705 ) | ( wire15709 ) | ( wire15710 ) ;
 assign wire15718 = ( n_n4988 ) | ( n_n4987 ) | ( wire251 ) ;
 assign wire15719 = ( n_n4991 ) | ( n_n4981 ) | ( n_n4985 ) | ( wire57 ) ;
 assign wire15721 = ( wire18  &  n_n524  &  n_n535 ) | ( wire18  &  n_n535  &  n_n520 ) ;
 assign wire15723 = ( wire24  &  n_n535  &  n_n195 ) | ( wire25  &  n_n535  &  n_n195 ) ;
 assign wire15724 = ( wire317 ) | ( wire341 ) ;
 assign wire15725 = ( n_n4958 ) | ( n_n4947 ) | ( wire15721 ) ;
 assign wire15726 = ( n_n4956 ) | ( n_n4965 ) | ( wire15723 ) ;
 assign wire15728 = ( wire228 ) | ( wire13217 ) | ( wire13218 ) | ( wire15726 ) ;
 assign wire15729 = ( wire15718 ) | ( wire15719 ) | ( wire15724 ) | ( wire15725 ) ;
 assign wire15733 = ( n_n4942 ) | ( wire59 ) | ( n_n4940 ) | ( n_n4939 ) ;
 assign wire15734 = ( n_n4946 ) | ( n_n4937 ) | ( wire180 ) | ( n_n4944 ) ;
 assign wire15738 = ( n_n4913 ) | ( n_n4916 ) | ( wire305 ) ;
 assign wire15739 = ( n_n4905 ) | ( n_n4918 ) | ( n_n4914 ) | ( wire340 ) ;
 assign wire15741 = ( wire15700 ) | ( wire15701 ) | ( wire15733 ) | ( wire15734 ) ;
 assign wire15742 = ( wire15738 ) | ( wire15739 ) | ( wire15741 ) ;
 assign wire15743 = ( wire15714 ) | ( wire15715 ) | ( wire15728 ) | ( wire15729 ) ;
 assign wire15746 = ( wire244 ) | ( n_n4725 ) | ( n_n4726 ) ;
 assign wire15747 = ( n_n4724 ) | ( n_n4727 ) | ( n_n4739 ) | ( wire95 ) ;
 assign wire15748 = ( wire11  &  n_n325  &  n_n518 ) | ( wire15  &  n_n325  &  n_n518 ) ;
 assign wire15750 = ( wire15748 ) | ( wire173 ) ;
 assign wire15754 = ( wire22  &  n_n482  &  n_n325 ) | ( wire25  &  n_n482  &  n_n325 ) ;
 assign wire15756 = ( n_n4784 ) | ( n_n4779 ) | ( n_n4786 ) | ( n_n4783 ) ;
 assign wire15757 = ( n_n4782 ) | ( n_n4781 ) | ( n_n4775 ) | ( wire15754 ) ;
 assign wire15758 = ( i_9_  &  n_n500  &  n_n520  &  n_n325 ) | ( (~ i_9_)  &  n_n500  &  n_n520  &  n_n325 ) ;
 assign wire15760 = ( n_n4756 ) | ( n_n4753 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire15761 = ( wire109 ) | ( n_n4752 ) | ( wire15758 ) ;
 assign wire15763 = ( wire14  &  n_n526  &  n_n491 ) | ( wire14  &  n_n528  &  n_n491 ) ;
 assign wire15764 = ( n_n4770 ) | ( n_n4764 ) | ( n_n4763 ) | ( n_n4765 ) ;
 assign wire15766 = ( n_n4771 ) | ( wire11748 ) | ( wire15763 ) | ( wire15764 ) ;
 assign wire15767 = ( wire15756 ) | ( wire15757 ) | ( wire15760 ) | ( wire15761 ) ;
 assign wire15769 = ( n_n4683 ) | ( n_n4678 ) | ( n_n4684 ) ;
 assign wire15770 = ( n_n4671 ) | ( n_n4672 ) | ( wire80 ) ;
 assign wire15773 = ( i_9_  &  n_n464  &  n_n520  &  n_n390 ) | ( (~ i_9_)  &  n_n464  &  n_n520  &  n_n390 ) ;
 assign wire15774 = ( wire444 ) | ( wire20  &  n_n464  &  n_n390 ) ;
 assign wire15775 = ( n_n4712 ) | ( n_n4685 ) | ( wire15773 ) ;
 assign wire15776 = ( n_n4707 ) | ( n_n4696 ) | ( wire13755 ) | ( wire13897 ) ;
 assign wire15778 = ( n_n4710 ) | ( n_n4709 ) | ( n_n4219 ) | ( wire15776 ) ;
 assign wire15781 = ( n_n4748 ) | ( n_n4747 ) | ( n_n4742 ) ;
 assign wire15782 = ( wire47 ) | ( wire374 ) ;
 assign wire15784 = ( n_n4749 ) | ( n_n4743 ) | ( wire15781 ) | ( wire15782 ) ;
 assign wire15786 = ( n_n2982 ) | ( wire15746 ) | ( wire15747 ) | ( wire15784 ) ;
 assign wire15790 = ( wire380 ) | ( wire158 ) ;
 assign wire15791 = ( n_n4787 ) | ( wire292 ) | ( n_n4795 ) | ( n_n4799 ) ;
 assign wire15792 = ( wire14  &  n_n473  &  n_n526 ) | ( wire14  &  n_n464  &  n_n526 ) ;
 assign wire15794 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4807 ) | ( n_n4808 ) ;
 assign wire15795 = ( n_n4801 ) | ( n_n4802 ) | ( wire15792 ) ;
 assign wire15798 = ( n_n4806 ) | ( n_n4805 ) | ( n_n4197 ) | ( wire390 ) ;
 assign wire15799 = ( wire15790 ) | ( wire15791 ) | ( wire15794 ) | ( wire15795 ) ;
 assign wire15800 = ( wire17  &  n_n524  &  n_n500 ) | ( wire17  &  n_n528  &  n_n500 ) ;
 assign wire15802 = ( wire15800 ) | ( wire174 ) ;
 assign wire15804 = ( n_n3450 ) | ( n_n4879 ) | ( n_n4884 ) | ( wire15802 ) ;
 assign wire15805 = ( wire15680 ) | ( wire15681 ) | ( wire15683 ) | ( wire15684 ) ;
 assign wire15807 = ( wire15696 ) | ( wire15697 ) | ( wire15798 ) | ( wire15799 ) ;
 assign wire15808 = ( wire15804 ) | ( wire15805 ) | ( wire15807 ) ;
 assign wire15811 = ( n_n2845 ) | ( n_n2846 ) | ( wire15315 ) | ( wire15316 ) ;
 assign wire15813 = ( n_n2827 ) | ( n_n2826 ) | ( wire15811 ) ;
 assign wire15816 = ( n_n2821 ) | ( n_n2907 ) | ( wire15813 ) ;
 assign wire15817 = ( n_n2906 ) | ( n_n2908 ) | ( n_n2902 ) | ( wire15677 ) ;
 assign wire15819 = ( wire21  &  n_n455  &  n_n491 ) | ( wire22  &  n_n455  &  n_n491 ) ;
 assign wire15822 = ( n_n4593 ) | ( n_n4594 ) | ( n_n4552 ) ;
 assign wire15823 = ( n_n4511 ) | ( n_n4590 ) | ( wire15819 ) ;
 assign wire15829 = ( n_n4641 ) | ( n_n4648 ) | ( n_n4651 ) | ( n_n4622 ) ;
 assign wire15830 = ( n_n4620 ) | ( n_n4627 ) | ( n_n4631 ) | ( wire255 ) ;
 assign wire15834 = ( wire13  &  n_n509  &  n_n520 ) | ( wire13  &  n_n509  &  n_n532 ) ;
 assign wire15836 = ( n_n4478 ) | ( n_n4502 ) | ( n_n4509 ) | ( n_n4471 ) ;
 assign wire15837 = ( n_n4473 ) | ( n_n4497 ) | ( wire617 ) | ( wire15834 ) ;
 assign wire15838 = ( wire15837 ) | ( wire15836 ) ;
 assign wire15841 = ( wire19  &  n_n509  &  n_n520 ) | ( wire19  &  n_n520  &  n_n482 ) ;
 assign wire15842 = ( wire11  &  n_n482  &  n_n65 ) | ( wire24  &  n_n482  &  n_n65 ) ;
 assign wire15843 = ( n_n5253 ) | ( wire25  &  n_n500  &  n_n65 ) ;
 assign wire15844 = ( n_n5238 ) | ( n_n5245 ) | ( n_n5280 ) ;
 assign wire15845 = ( wire15842 ) | ( wire15841 ) ;
 assign wire15848 = ( wire17  &  n_n509  &  n_n522 ) | ( wire17  &  n_n509  &  n_n530 ) ;
 assign wire15851 = ( n_n4849 ) | ( n_n4790 ) | ( n_n4813 ) ;
 assign wire15852 = ( n_n4821 ) | ( n_n4842 ) | ( wire15848 ) ;
 assign wire15858 = ( n_n4887 ) | ( n_n4930 ) | ( n_n4929 ) ;
 assign wire15859 = ( n_n4912 ) | ( n_n4968 ) | ( n_n4967 ) | ( n_n4899 ) ;
 assign wire15864 = ( n_n4993 ) | ( n_n4994 ) | ( wire248 ) ;
 assign wire15865 = ( wire136 ) | ( n_n5009 ) | ( n_n4978 ) | ( n_n5001 ) ;
 assign wire15870 = ( n_n5111 ) | ( n_n5081 ) | ( n_n5080 ) ;
 assign wire15871 = ( n_n5098 ) | ( n_n5087 ) | ( n_n5116 ) | ( n_n5102 ) ;
 assign wire15873 = ( i_9_  &  n_n473  &  n_n532  &  n_n130 ) | ( (~ i_9_)  &  n_n473  &  n_n532  &  n_n130 ) ;
 assign wire15875 = ( wire12  &  n_n522  &  n_n473 ) | ( wire12  &  n_n473  &  n_n520 ) ;
 assign wire15876 = ( wire15  &  n_n500  &  n_n130 ) | ( wire15  &  n_n491  &  n_n130 ) ;
 assign wire15879 = ( n_n5138 ) | ( wire15873 ) | ( wire15876 ) ;
 assign wire15880 = ( wire18  &  n_n473  &  n_n532 ) | ( wire18  &  n_n482  &  n_n532 ) ;
 assign wire15885 = ( n_n5059 ) | ( n_n5018 ) | ( n_n5022 ) | ( n_n5046 ) ;
 assign wire15886 = ( n_n5033 ) | ( n_n5063 ) | ( n_n5052 ) | ( wire15880 ) ;
 assign wire15887 = ( wire15886 ) | ( wire15885 ) ;
 assign wire15892 = ( i_9_  &  n_n524  &  n_n535  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n65 ) ;
 assign wire15894 = ( n_n5214 ) | ( n_n5207 ) | ( n_n5229 ) | ( n_n5221 ) ;
 assign wire15895 = ( n_n5200 ) | ( n_n5222 ) | ( n_n5203 ) | ( wire15892 ) ;
 assign wire15897 = ( wire21  &  n_n464  &  n_n65 ) | ( wire20  &  n_n464  &  n_n65 ) ;
 assign wire15898 = ( n_n5325 ) | ( n_n5303 ) | ( wire15897 ) ;
 assign wire15899 = ( wire15843 ) | ( wire15844 ) | ( wire15845 ) | ( wire15898 ) ;
 assign wire15901 = ( wire15864 ) | ( wire15865 ) | ( wire15894 ) | ( wire15895 ) ;
 assign wire15902 = ( n_n1722 ) | ( n_n1721 ) | ( wire15899 ) ;
 assign wire15903 = ( n_n1718 ) | ( n_n1717 ) | ( wire15887 ) | ( wire15901 ) ;
 assign wire15908 = ( n_n4420 ) | ( n_n4407 ) | ( n_n4412 ) ;
 assign wire15909 = ( n_n4373 ) | ( n_n4392 ) | ( n_n4426 ) | ( n_n4419 ) ;
 assign wire15914 = ( n_n4432 ) | ( n_n4435 ) | ( n_n4468 ) ;
 assign wire15915 = ( n_n4464 ) | ( n_n4455 ) | ( n_n4433 ) | ( n_n4441 ) ;
 assign wire15920 = ( n_n4676 ) | ( n_n4655 ) | ( wire391 ) ;
 assign wire15922 = ( wire23  &  n_n535  &  n_n325 ) | ( wire23  &  n_n325  &  n_n518 ) ;
 assign wire15924 = ( wire15922 ) | ( wire444 ) ;
 assign wire15927 = ( wire21  &  n_n482  &  n_n325 ) | ( wire15  &  n_n482  &  n_n325 ) ;
 assign wire15930 = ( n_n4784 ) | ( n_n4754 ) | ( wire15927 ) ;
 assign wire15931 = ( n_n4748 ) | ( n_n4772 ) | ( wire164 ) | ( n_n4766 ) ;
 assign wire15937 = ( n_n4337 ) | ( n_n4314 ) | ( n_n4345 ) | ( wire675 ) ;
 assign wire15938 = ( n_n4371 ) | ( n_n4343 ) | ( n_n4320 ) | ( wire345 ) ;
 assign wire15941 = ( n_n1730 ) | ( n_n1729 ) | ( wire15937 ) | ( wire15938 ) ;
 assign wire15943 = ( n_n1712 ) | ( n_n1711 ) | ( wire15941 ) ;
 assign wire15945 = ( wire209 ) | ( wire123 ) ;
 assign wire15947 = ( i_9_  &  n_n522  &  n_n535  &  n_n130 ) | ( (~ i_9_)  &  n_n522  &  n_n535  &  n_n130 ) ;
 assign wire15950 = ( wire15947 ) | ( wire279 ) ;
 assign wire15951 = ( n_n5089 ) | ( n_n5086 ) | ( n_n5088 ) | ( wire232 ) ;
 assign wire15952 = ( wire18  &  n_n522  &  n_n473 ) | ( wire18  &  n_n473  &  n_n528 ) ;
 assign wire15954 = ( n_n5057 ) | ( n_n5058 ) | ( n_n5065 ) ;
 assign wire15955 = ( wire15952 ) | ( wire160 ) ;
 assign wire15957 = ( n_n5067 ) | ( n_n5064 ) | ( wire15954 ) | ( wire15955 ) ;
 assign wire15961 = ( n_n5118 ) | ( n_n5121 ) | ( n_n5122 ) ;
 assign wire15962 = ( n_n5123 ) | ( n_n5114 ) | ( wire336 ) ;
 assign wire15964 = ( wire21  &  n_n518  &  n_n130 ) | ( wire20  &  n_n518  &  n_n130 ) ;
 assign wire15967 = ( n_n5112 ) | ( n_n5110 ) | ( wire15964 ) ;
 assign wire15968 = ( n_n5113 ) | ( n_n5104 ) | ( n_n5106 ) | ( wire122 ) ;
 assign wire15970 = ( wire12  &  n_n522  &  n_n500 ) | ( wire12  &  n_n500  &  n_n530 ) ;
 assign wire15972 = ( n_n5136 ) | ( n_n5135 ) | ( n_n5134 ) | ( wire15970 ) ;
 assign wire15973 = ( n_n5130 ) | ( n_n5129 ) | ( wire422 ) | ( wire15972 ) ;
 assign wire15975 = ( wire18  &  n_n524  &  n_n482 ) | ( wire18  &  n_n528  &  n_n482 ) ;
 assign wire15977 = ( n_n5048 ) | ( n_n5047 ) | ( n_n5044 ) ;
 assign wire15978 = ( wire15975 ) | ( wire97 ) ;
 assign wire15980 = ( wire18  &  n_n524  &  n_n491 ) | ( wire18  &  n_n491  &  n_n534 ) ;
 assign wire15982 = ( wire265 ) | ( wire296 ) ;
 assign wire15983 = ( wire135 ) | ( n_n5020 ) | ( wire15980 ) ;
 assign wire15985 = ( i_9_  &  n_n530  &  n_n482  &  n_n195 ) | ( (~ i_9_)  &  n_n530  &  n_n482  &  n_n195 ) ;
 assign wire15987 = ( n_n5035 ) | ( n_n5032 ) | ( n_n5027 ) | ( n_n5028 ) ;
 assign wire15989 = ( wire50 ) | ( n_n5029 ) | ( wire15985 ) | ( wire15987 ) ;
 assign wire15991 = ( n_n1842 ) | ( wire15982 ) | ( wire15983 ) | ( wire15989 ) ;
 assign wire15993 = ( wire13  &  n_n526  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire15995 = ( n_n4489 ) | ( n_n4488 ) | ( n_n4490 ) | ( wire15993 ) ;
 assign wire15996 = ( wire184 ) | ( wire11  &  n_n509  &  n_n455 ) ;
 assign wire15999 = ( i_9_  &  n_n522  &  n_n536  &  n_n464 ) | ( (~ i_9_)  &  n_n522  &  n_n536  &  n_n464 ) ;
 assign wire16001 = ( n_n4434 ) | ( wire234 ) | ( n_n4431 ) ;
 assign wire16002 = ( wire233 ) | ( n_n4447 ) | ( wire15999 ) ;
 assign wire16003 = ( n_n4470 ) | ( n_n4472 ) | ( n_n4469 ) ;
 assign wire16004 = ( n_n4449 ) | ( n_n4465 ) | ( wire11505 ) | ( wire14133 ) ;
 assign wire16007 = ( n_n4462 ) | ( n_n2058 ) | ( wire12471 ) | ( wire16004 ) ;
 assign wire16008 = ( n_n3889 ) | ( wire16001 ) | ( wire16002 ) | ( wire16003 ) ;
 assign wire16009 = ( wire21  &  n_n455  &  n_n482 ) | ( wire20  &  n_n455  &  n_n482 ) ;
 assign wire16011 = ( n_n4535 ) | ( n_n4536 ) | ( wire16009 ) ;
 assign wire16012 = ( n_n4532 ) | ( n_n4537 ) | ( n_n4529 ) | ( wire11532 ) ;
 assign wire16014 = ( wire170 ) | ( wire20  &  n_n455  &  n_n491 ) ;
 assign wire16015 = ( n_n4520 ) | ( wire361 ) | ( wire789 ) ;
 assign wire16016 = ( n_n4521 ) | ( n_n4526 ) | ( n_n4542 ) | ( wire201 ) ;
 assign wire16018 = ( wire16016 ) | ( wire202 ) ;
 assign wire16019 = ( wire16011 ) | ( wire16012 ) | ( wire16014 ) | ( wire16015 ) ;
 assign wire16020 = ( wire13  &  n_n524  &  n_n491 ) | ( wire13  &  n_n526  &  n_n491 ) ;
 assign wire16022 = ( n_n4506 ) | ( n_n4505 ) | ( wire606 ) ;
 assign wire16023 = ( n_n4504 ) | ( n_n4503 ) | ( wire16020 ) ;
 assign wire16025 = ( n_n4500 ) | ( n_n4508 ) | ( wire16022 ) | ( wire16023 ) ;
 assign wire16028 = ( wire16007 ) | ( wire16008 ) | ( wire16018 ) | ( wire16019 ) ;
 assign wire16030 = ( n_n4582 ) | ( n_n4581 ) | ( wire276 ) ;
 assign wire16031 = ( n_n4584 ) | ( n_n4580 ) | ( n_n4585 ) | ( wire12520 ) ;
 assign wire16032 = ( wire11  &  n_n535  &  n_n390 ) | ( wire24  &  n_n535  &  n_n390 ) ;
 assign wire16034 = ( n_n4570 ) | ( n_n4569 ) | ( wire266 ) ;
 assign wire16035 = ( wire16032 ) | ( wire99 ) ;
 assign wire16038 = ( wire45 ) | ( n_n4591 ) | ( n_n4592 ) ;
 assign wire16040 = ( n_n4612 ) | ( n_n4608 ) | ( n_n4609 ) ;
 assign wire16041 = ( n_n4613 ) | ( n_n4605 ) | ( wire465 ) | ( wire12519 ) ;
 assign wire16045 = ( n_n4616 ) | ( n_n4619 ) | ( n_n4623 ) ;
 assign wire16046 = ( n_n4617 ) | ( n_n4628 ) | ( n_n4621 ) | ( n_n4630 ) ;
 assign wire16048 = ( n_n4626 ) | ( n_n4625 ) | ( wire16045 ) | ( wire16046 ) ;
 assign wire16052 = ( n_n4669 ) | ( n_n4670 ) | ( n_n4665 ) ;
 assign wire16053 = ( n_n4666 ) | ( n_n4662 ) | ( n_n4671 ) | ( n_n4672 ) ;
 assign wire16056 = ( wire10  &  n_n522  &  n_n482 ) | ( wire10  &  n_n530  &  n_n482 ) ;
 assign wire16057 = ( wire10  &  n_n528  &  n_n482 ) | ( wire10  &  n_n482  &  n_n532 ) ;
 assign wire16059 = ( n_n4646 ) | ( n_n4659 ) | ( wire16056 ) ;
 assign wire16060 = ( wire309 ) | ( n_n4642 ) | ( wire16057 ) ;
 assign wire16064 = ( n_n4639 ) | ( n_n4635 ) | ( n_n4632 ) | ( wire15132 ) ;
 assign wire16065 = ( n_n4634 ) | ( wire26 ) | ( n_n4633 ) | ( wire16064 ) ;
 assign wire16069 = ( n_n4560 ) | ( wire471 ) | ( wire91 ) | ( n_n4551 ) ;
 assign wire16070 = ( n_n4557 ) | ( wire430 ) | ( n_n4558 ) | ( wire16069 ) ;
 assign wire16072 = ( n_n1879 ) | ( wire16030 ) | ( wire16031 ) | ( wire16070 ) ;
 assign wire16075 = ( i_9_  &  n_n509  &  n_n536  &  n_n530 ) | ( (~ i_9_)  &  n_n509  &  n_n536  &  n_n530 ) ;
 assign wire16077 = ( n_n4344 ) | ( n_n4347 ) | ( wire53 ) ;
 assign wire16078 = ( n_n4335 ) | ( wire124 ) | ( wire16075 ) ;
 assign wire16081 = ( wire364 ) | ( wire171 ) ;
 assign wire16082 = ( n_n4334 ) | ( wire106 ) | ( wire677 ) ;
 assign wire16083 = ( n_n4318 ) | ( n_n4331 ) | ( n_n4326 ) | ( n_n4313 ) ;
 assign wire16086 = ( n_n4279 ) | ( n_n4323 ) | ( wire12569 ) | ( wire16083 ) ;
 assign wire16087 = ( wire16077 ) | ( wire16078 ) | ( wire16081 ) | ( wire16082 ) ;
 assign wire16088 = ( wire16  &  n_n522  &  n_n500 ) | ( wire16  &  n_n500  &  n_n520 ) ;
 assign wire16089 = ( wire16088 ) | ( wire23  &  n_n536  &  n_n500 ) ;
 assign wire16091 = ( n_n4380 ) | ( wire280 ) | ( n_n4377 ) ;
 assign wire16093 = ( wire16  &  n_n473  &  n_n524 ) | ( wire16  &  n_n473  &  n_n528 ) ;
 assign wire16094 = ( n_n4430 ) | ( n_n4416 ) | ( wire37 ) ;
 assign wire16095 = ( n_n4421 ) | ( wire215 ) | ( wire16093 ) ;
 assign wire16098 = ( n_n4397 ) | ( n_n4398 ) | ( n_n4399 ) ;
 assign wire16099 = ( n_n4389 ) | ( n_n4388 ) | ( n_n4393 ) | ( n_n4390 ) ;
 assign wire16102 = ( n_n4405 ) | ( n_n4406 ) | ( n_n4411 ) ;
 assign wire16103 = ( n_n4401 ) | ( n_n4409 ) | ( n_n4410 ) | ( n_n4402 ) ;
 assign wire16105 = ( n_n4403 ) | ( n_n4400 ) | ( wire16102 ) | ( wire16103 ) ;
 assign wire16109 = ( n_n4357 ) | ( n_n4358 ) | ( n_n4354 ) ;
 assign wire16110 = ( n_n4361 ) | ( n_n4363 ) | ( n_n4359 ) | ( n_n4356 ) ;
 assign wire16112 = ( n_n4350 ) | ( n_n4355 ) | ( wire16109 ) | ( wire16110 ) ;
 assign wire16114 = ( wire54 ) | ( n_n1894 ) | ( wire16091 ) | ( wire16112 ) ;
 assign wire16119 = ( n_n4735 ) | ( n_n4744 ) | ( wire374 ) ;
 assign wire16120 = ( n_n4734 ) | ( n_n4729 ) | ( n_n4728 ) | ( wire373 ) ;
 assign wire16121 = ( wire21  &  n_n500  &  n_n325 ) | ( wire15  &  n_n500  &  n_n325 ) ;
 assign wire16124 = ( n_n4756 ) | ( n_n4753 ) | ( wire16121 ) ;
 assign wire16125 = ( wire109 ) | ( n_n4747 ) | ( n_n4752 ) | ( n_n4745 ) ;
 assign wire16127 = ( n_n4724 ) | ( n_n4723 ) | ( n_n4722 ) ;
 assign wire16128 = ( n_n4720 ) | ( n_n4719 ) | ( wire173 ) ;
 assign wire16130 = ( n_n4718 ) | ( n_n4717 ) | ( wire16127 ) | ( wire16128 ) ;
 assign wire16131 = ( wire16119 ) | ( wire16120 ) | ( wire16124 ) | ( wire16125 ) ;
 assign wire16132 = ( wire25  &  n_n535  &  n_n325 ) | ( wire15  &  n_n535  &  n_n325 ) ;
 assign wire16134 = ( wire445 ) | ( wire221 ) ;
 assign wire16135 = ( n_n4692 ) | ( n_n4695 ) | ( n_n4696 ) | ( wire16132 ) ;
 assign wire16138 = ( n_n4708 ) | ( wire21  &  n_n535  &  n_n325 ) ;
 assign wire16139 = ( n_n4683 ) | ( n_n4684 ) | ( n_n4680 ) ;
 assign wire16140 = ( n_n4685 ) | ( n_n4686 ) | ( wire80 ) ;
 assign wire16141 = ( n_n4689 ) | ( n_n4712 ) | ( n_n4681 ) | ( n_n4705 ) ;
 assign wire16144 = ( n_n4219 ) | ( wire30 ) | ( wire16138 ) | ( wire16139 ) ;
 assign wire16145 = ( wire16134 ) | ( wire16135 ) | ( wire16140 ) | ( wire16141 ) ;
 assign wire16146 = ( wire18  &  n_n509  &  n_n522 ) | ( wire18  &  n_n509  &  n_n526 ) ;
 assign wire16148 = ( n_n4988 ) | ( n_n4987 ) | ( wire16146 ) ;
 assign wire16149 = ( n_n4999 ) | ( n_n4986 ) | ( n_n4989 ) | ( wire13997 ) ;
 assign wire16152 = ( wire393 ) | ( wire252 ) ;
 assign wire16153 = ( n_n4983 ) | ( n_n4984 ) | ( wire228 ) ;
 assign wire16155 = ( n_n4979 ) | ( n_n4985 ) | ( wire12255 ) | ( wire12256 ) ;
 assign wire16157 = ( n_n4975 ) | ( n_n5000 ) | ( wire299 ) | ( wire16155 ) ;
 assign wire16158 = ( wire16148 ) | ( wire16149 ) | ( wire16152 ) | ( wire16153 ) ;
 assign wire16159 = ( wire17  &  n_n473  &  n_n526 ) | ( wire17  &  n_n473  &  n_n534 ) ;
 assign wire16164 = ( n_n4940 ) | ( n_n4939 ) | ( wire180 ) ;
 assign wire16165 = ( n_n4937 ) | ( n_n4938 ) | ( wire305 ) ;
 assign wire16166 = ( n_n4907 ) | ( n_n4942 ) | ( n_n4936 ) | ( n_n4933 ) ;
 assign wire16168 = ( n_n4919 ) | ( n_n4910 ) | ( wire13870 ) | ( wire16166 ) ;
 assign wire16170 = ( wire317 ) | ( wire17  &  n_n464  &  n_n520 ) ;
 assign wire16171 = ( n_n4948 ) | ( n_n4944 ) | ( wire13867 ) | ( wire14962 ) ;
 assign wire16173 = ( n_n4953 ) | ( wire771 ) | ( wire772 ) ;
 assign wire16174 = ( n_n4959 ) | ( n_n4960 ) | ( wire141 ) ;
 assign wire16175 = ( n_n4962 ) | ( n_n4971 ) | ( n_n4973 ) | ( wire11809 ) ;
 assign wire16176 = ( n_n4965 ) | ( n_n4955 ) | ( wire13215 ) | ( wire13216 ) ;
 assign wire16179 = ( wire16170 ) | ( wire16171 ) | ( wire16173 ) | ( wire16174 ) ;
 assign wire16180 = ( wire16175 ) | ( wire16176 ) | ( wire16179 ) ;
 assign wire16182 = ( wire11  &  n_n491  &  n_n260 ) | ( wire23  &  n_n491  &  n_n260 ) ;
 assign wire16184 = ( n_n4898 ) | ( wire352 ) | ( n_n4897 ) ;
 assign wire16185 = ( wire96 ) | ( n_n4901 ) | ( wire16182 ) ;
 assign wire16186 = ( wire14  &  n_n473  &  n_n526 ) | ( wire14  &  n_n473  &  n_n520 ) ;
 assign wire16188 = ( n_n4803 ) | ( n_n4804 ) | ( n_n4799 ) ;
 assign wire16189 = ( n_n4807 ) | ( n_n4808 ) | ( wire16186 ) ;
 assign wire16192 = ( i_9_  &  n_n535  &  n_n534  &  n_n260 ) | ( (~ i_9_)  &  n_n535  &  n_n534  &  n_n260 ) ;
 assign wire16193 = ( n_n4816 ) | ( n_n4818 ) | ( n_n4815 ) ;
 assign wire16194 = ( n_n4834 ) | ( n_n4833 ) | ( wire150 ) ;
 assign wire16195 = ( n_n4832 ) | ( n_n4812 ) | ( wire16192 ) ;
 assign wire16198 = ( wire388 ) | ( n_n4197 ) | ( wire16195 ) ;
 assign wire16201 = ( i_9_  &  n_n520  &  n_n518  &  n_n260 ) | ( (~ i_9_)  &  n_n520  &  n_n518  &  n_n260 ) ;
 assign wire16203 = ( n_n4857 ) | ( n_n4858 ) | ( wire375 ) ;
 assign wire16204 = ( n_n4848 ) | ( wire52 ) | ( wire16201 ) ;
 assign wire16206 = ( n_n4862 ) | ( wire40 ) | ( n_n4861 ) ;
 assign wire16207 = ( n_n4859 ) | ( n_n4864 ) | ( n_n4866 ) | ( wire13810 ) ;
 assign wire16211 = ( n_n4835 ) | ( n_n4843 ) | ( n_n4839 ) | ( n_n4840 ) ;
 assign wire16212 = ( wire176 ) | ( n_n4841 ) | ( n_n4838 ) | ( n_n4836 ) ;
 assign wire16213 = ( wire16212 ) | ( wire16211 ) ;
 assign wire16214 = ( wire16203 ) | ( wire16204 ) | ( wire16206 ) | ( wire16207 ) ;
 assign wire16215 = ( i_9_  &  n_n528  &  n_n500  &  n_n260 ) | ( (~ i_9_)  &  n_n528  &  n_n500  &  n_n260 ) ;
 assign wire16217 = ( n_n4882 ) | ( n_n4881 ) | ( wire16215 ) ;
 assign wire16220 = ( wire261 ) | ( wire264 ) ;
 assign wire16222 = ( n_n4886 ) | ( n_n4891 ) | ( n_n1985 ) | ( wire16220 ) ;
 assign wire16224 = ( n_n1856 ) | ( wire16184 ) | ( wire16185 ) | ( wire16222 ) ;
 assign wire16228 = ( n_n4791 ) | ( n_n4792 ) | ( wire380 ) ;
 assign wire16229 = ( n_n4789 ) | ( n_n4793 ) | ( n_n4797 ) | ( wire179 ) ;
 assign wire16232 = ( n_n4765 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire16233 = ( n_n4757 ) | ( n_n4759 ) | ( n_n4760 ) | ( n_n4767 ) ;
 assign wire16236 = ( n_n4782 ) | ( n_n4777 ) | ( n_n4788 ) ;
 assign wire16238 = ( n_n4204 ) | ( n_n3469 ) | ( wire16236 ) ;
 assign wire16240 = ( n_n1865 ) | ( wire16228 ) | ( wire16229 ) | ( wire16238 ) ;
 assign wire16241 = ( wire16130 ) | ( wire16131 ) | ( wire16144 ) | ( wire16145 ) ;
 assign wire16245 = ( n_n5161 ) | ( n_n5162 ) | ( n_n5163 ) ;
 assign wire16246 = ( wire12  &  n_n520  &  n_n482 ) | ( wire12  &  n_n530  &  n_n482 ) ;
 assign wire16248 = ( wire332 ) | ( wire437 ) ;
 assign wire16249 = ( wire254 ) | ( n_n5170 ) | ( wire16246 ) ;
 assign wire16251 = ( wire22  &  n_n473  &  n_n130 ) | ( wire11  &  n_n473  &  n_n130 ) ;
 assign wire16253 = ( n_n5181 ) | ( n_n5184 ) | ( n_n5175 ) | ( n_n5177 ) ;
 assign wire16254 = ( wire112 ) | ( n_n5182 ) | ( wire16251 ) ;
 assign wire16256 = ( wire22  &  n_n464  &  n_n130 ) | ( wire11  &  n_n464  &  n_n130 ) ;
 assign wire16257 = ( wire454 ) | ( wire220 ) ;
 assign wire16258 = ( n_n5191 ) | ( wire452 ) | ( n_n5192 ) ;
 assign wire16259 = ( n_n5212 ) | ( n_n5189 ) | ( wire16256 ) ;
 assign wire16262 = ( n_n5194 ) | ( n_n2291 ) | ( wire453 ) | ( wire16259 ) ;
 assign wire16263 = ( wire16253 ) | ( wire16254 ) | ( wire16257 ) | ( wire16258 ) ;
 assign wire16266 = ( n_n5239 ) | ( n_n5240 ) | ( n_n5246 ) ;
 assign wire16267 = ( n_n5244 ) | ( n_n5241 ) | ( wire386 ) ;
 assign wire16270 = ( i_9_  &  n_n534  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n534  &  n_n518  &  n_n65 ) ;
 assign wire16272 = ( n_n5228 ) | ( n_n5220 ) | ( wire182 ) ;
 assign wire16273 = ( wire385 ) | ( n_n5215 ) | ( wire16270 ) ;
 assign wire16278 = ( n_n5258 ) | ( n_n5251 ) | ( n_n5249 ) | ( n_n5252 ) ;
 assign wire16279 = ( n_n5259 ) | ( wire409 ) | ( n_n5247 ) | ( n_n5250 ) ;
 assign wire16280 = ( wire16279 ) | ( wire16278 ) ;
 assign wire16282 = ( wire12  &  n_n524  &  n_n491 ) | ( wire12  &  n_n491  &  n_n532 ) ;
 assign wire16286 = ( n_n5150 ) | ( n_n5147 ) | ( wire196 ) | ( n_n5148 ) ;
 assign wire16288 = ( wire466 ) | ( wire16245 ) | ( wire16248 ) | ( wire16249 ) ;
 assign wire16289 = ( wire288 ) | ( wire16282 ) | ( wire16286 ) | ( wire16288 ) ;
 assign wire16291 = ( i_9_  &  n_n473  &  n_n524  &  n_n65 ) | ( (~ i_9_)  &  n_n473  &  n_n524  &  n_n65 ) ;
 assign wire16293 = ( wire19  &  n_n528  &  n_n491 ) | ( wire19  &  n_n491  &  n_n530 ) ;
 assign wire16294 = ( wire22  &  n_n491  &  n_n65 ) | ( wire23  &  n_n491  &  n_n65 ) ;
 assign wire16296 = ( wire16293 ) | ( wire218 ) ;
 assign wire16297 = ( wire441 ) | ( n_n5279 ) | ( wire16294 ) ;
 assign wire16299 = ( n_n5290 ) | ( n_n5292 ) | ( n_n5289 ) ;
 assign wire16300 = ( n_n5293 ) | ( n_n5297 ) | ( n_n5294 ) | ( n_n5298 ) ;
 assign wire16305 = ( n_n5275 ) | ( n_n5271 ) | ( n_n5264 ) | ( wire77 ) ;
 assign wire16306 = ( wire25  &  n_n473  &  n_n65 ) | ( wire15  &  n_n473  &  n_n65 ) ;
 assign wire16308 = ( n_n5307 ) | ( n_n5308 ) | ( wire63 ) ;
 assign wire16309 = ( wire269 ) | ( n_n5304 ) | ( wire16306 ) ;
 assign wire16310 = ( wire19  &  n_n522  &  n_n464 ) | ( wire19  &  n_n464  &  n_n528 ) ;
 assign wire16312 = ( n_n5318 ) | ( n_n5320 ) | ( n_n5330 ) ;
 assign wire16313 = ( n_n5329 ) | ( n_n5319 ) | ( wire16310 ) ;
 assign wire16316 = ( n_n1900 ) | ( wire16296 ) | ( wire16297 ) | ( wire16312 ) ;
 assign wire16318 = ( wire117 ) | ( wire16308 ) | ( wire16309 ) | ( wire16313 ) ;
 assign wire16320 = ( n_n1786 ) | ( n_n1801 ) | ( n_n1800 ) | ( wire15991 ) ;
 assign wire16323 = ( wire15902 ) | ( wire15903 ) | ( wire15943 ) | ( wire16320 ) ;
 assign wire16324 = ( n_n1793 ) | ( n_n1792 ) | ( n_n1794 ) | ( n_n1787 ) ;
 assign wire16327 = ( n_n4945 ) | ( n_n4946 ) | ( n_n4949 ) ;
 assign wire16331 = ( n_n4888 ) | ( n_n4885 ) | ( wire260 ) ;
 assign wire16334 = ( n_n4862 ) | ( n_n4850 ) | ( n_n4861 ) ;
 assign wire16335 = ( wire295 ) | ( wire277 ) ;
 assign wire16339 = ( n_n4877 ) | ( n_n4870 ) | ( n_n4872 ) ;
 assign wire16340 = ( n_n4881 ) | ( n_n4878 ) | ( wire174 ) ;
 assign wire16342 = ( n_n4880 ) | ( n_n4869 ) | ( wire16339 ) | ( wire16340 ) ;
 assign wire16345 = ( wire14  &  n_n522  &  n_n473 ) | ( wire14  &  n_n473  &  n_n532 ) ;
 assign wire16346 = ( wire24  &  n_n473  &  n_n325 ) | ( wire25  &  n_n473  &  n_n325 ) ;
 assign wire16347 = ( i_9_  &  n_n473  &  n_n530  &  n_n325 ) | ( (~ i_9_)  &  n_n473  &  n_n530  &  n_n325 ) ;
 assign wire16349 = ( wire16346 ) | ( wire16345 ) ;
 assign wire16350 = ( n_n4791 ) | ( n_n4798 ) | ( n_n4801 ) | ( wire16347 ) ;
 assign wire16351 = ( i_9_  &  n_n524  &  n_n535  &  n_n260 ) | ( (~ i_9_)  &  n_n524  &  n_n535  &  n_n260 ) ;
 assign wire16352 = ( n_n4832 ) | ( n_n4825 ) | ( n_n4826 ) ;
 assign wire16355 = ( n_n4842 ) | ( n_n4837 ) | ( n_n4841 ) ;
 assign wire16356 = ( n_n4839 ) | ( n_n4840 ) | ( wire176 ) ;
 assign wire16360 = ( wire14  &  n_n522  &  n_n464 ) | ( wire14  &  n_n524  &  n_n464 ) ;
 assign wire16362 = ( n_n4824 ) | ( n_n4822 ) | ( n_n4823 ) | ( n_n4806 ) ;
 assign wire16363 = ( n_n4810 ) | ( wire186 ) | ( wire16360 ) ;
 assign wire16366 = ( wire11  &  n_n491  &  n_n325 ) | ( wire24  &  n_n491  &  n_n325 ) ;
 assign wire16367 = ( wire164 ) | ( n_n4765 ) | ( n_n4766 ) ;
 assign wire16368 = ( n_n4770 ) | ( n_n4773 ) | ( n_n4771 ) | ( wire16366 ) ;
 assign wire16373 = ( n_n4776 ) | ( n_n4774 ) | ( n_n4786 ) | ( wire131 ) ;
 assign wire16374 = ( n_n4779 ) | ( n_n4790 ) | ( wire313 ) | ( wire16373 ) ;
 assign wire16375 = ( wire16349 ) | ( wire16350 ) | ( wire16367 ) | ( wire16368 ) ;
 assign wire16378 = ( i_9_  &  n_n500  &  n_n530  &  n_n325 ) | ( (~ i_9_)  &  n_n500  &  n_n530  &  n_n325 ) ;
 assign wire16379 = ( wire22  &  n_n500  &  n_n325 ) | ( wire24  &  n_n500  &  n_n325 ) ;
 assign wire16382 = ( wire16379 ) | ( wire16378 ) ;
 assign wire16383 = ( wire373 ) | ( n_n4752 ) | ( n_n4751 ) | ( n_n4750 ) ;
 assign wire16385 = ( n_n4732 ) | ( wire293 ) | ( wire767 ) ;
 assign wire16386 = ( n_n4738 ) | ( wire95 ) | ( n_n4733 ) | ( n_n4736 ) ;
 assign wire16388 = ( n_n4725 ) | ( n_n4726 ) | ( n_n4729 ) ;
 assign wire16389 = ( wire244 ) | ( n_n4722 ) | ( n_n4721 ) ;
 assign wire16394 = ( n_n4695 ) | ( n_n4696 ) | ( wire173 ) ;
 assign wire16395 = ( n_n4711 ) | ( n_n4712 ) | ( wire442 ) ;
 assign wire16396 = ( n_n4709 ) | ( n_n4698 ) | ( n_n4707 ) | ( n_n4702 ) ;
 assign wire16399 = ( n_n4216 ) | ( n_n2378 ) | ( wire16396 ) ;
 assign wire16404 = ( n_n4669 ) | ( n_n4670 ) | ( wire81 ) ;
 assign wire16405 = ( n_n4673 ) | ( n_n4676 ) | ( n_n4681 ) | ( n_n4679 ) ;
 assign wire16408 = ( wire10  &  n_n522  &  n_n482 ) | ( wire10  &  n_n524  &  n_n482 ) ;
 assign wire16409 = ( wire10  &  n_n464  &  n_n526 ) | ( wire10  &  n_n464  &  n_n528 ) ;
 assign wire16410 = ( wire431 ) | ( wire22  &  n_n390  &  n_n482 ) ;
 assign wire16411 = ( n_n4662 ) | ( n_n4683 ) | ( wire16408 ) ;
 assign wire16412 = ( n_n4667 ) | ( n_n4664 ) | ( n_n4663 ) | ( wire16409 ) ;
 assign wire16415 = ( n_n3849 ) | ( n_n4693 ) | ( wire12422 ) | ( wire16412 ) ;
 assign wire16420 = ( n_n4758 ) | ( n_n4761 ) | ( n_n4762 ) ;
 assign wire16421 = ( n_n4754 ) | ( n_n4757 ) | ( n_n4756 ) | ( n_n4755 ) ;
 assign wire16423 = ( n_n4759 ) | ( n_n4760 ) | ( wire16420 ) | ( wire16421 ) ;
 assign wire16424 = ( wire16382 ) | ( wire16383 ) | ( wire16385 ) | ( wire16386 ) ;
 assign wire16427 = ( i_9_  &  n_n509  &  n_n520  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n520  &  n_n195 ) ;
 assign wire16430 = ( wire16427 ) | ( wire393 ) ;
 assign wire16431 = ( n_n5004 ) | ( wire136 ) | ( n_n4994 ) | ( n_n5001 ) ;
 assign wire16435 = ( n_n5018 ) | ( n_n5015 ) | ( wire343 ) ;
 assign wire16436 = ( n_n5016 ) | ( n_n5009 ) | ( n_n5013 ) | ( wire297 ) ;
 assign wire16438 = ( i_9_  &  n_n509  &  n_n534  &  n_n195 ) | ( (~ i_9_)  &  n_n509  &  n_n534  &  n_n195 ) ;
 assign wire16440 = ( n_n4990 ) | ( n_n4988 ) | ( n_n4987 ) | ( n_n4979 ) ;
 assign wire16442 = ( n_n4986 ) | ( wire251 ) | ( wire16438 ) | ( wire16440 ) ;
 assign wire16443 = ( wire16430 ) | ( wire16431 ) | ( wire16435 ) | ( wire16436 ) ;
 assign wire16445 = ( wire31 ) | ( wire23  &  n_n473  &  n_n260 ) ;
 assign wire16447 = ( wire11  &  n_n482  &  n_n260 ) | ( wire15  &  n_n482  &  n_n260 ) ;
 assign wire16448 = ( wire20  &  n_n491  &  n_n260 ) | ( wire23  &  n_n491  &  n_n260 ) ;
 assign wire16449 = ( n_n4900 ) | ( n_n4899 ) | ( wire16447 ) ;
 assign wire16450 = ( n_n4898 ) | ( n_n4897 ) | ( n_n4896 ) | ( wire16448 ) ;
 assign wire16453 = ( n_n4913 ) | ( n_n4914 ) | ( n_n4915 ) ;
 assign wire16454 = ( n_n4920 ) | ( n_n4923 ) | ( n_n4918 ) | ( n_n4917 ) ;
 assign wire16456 = ( n_n4921 ) | ( n_n4919 ) | ( wire16453 ) | ( wire16454 ) ;
 assign wire16460 = ( wire362 ) | ( wire341 ) ;
 assign wire16461 = ( n_n4966 ) | ( n_n4978 ) | ( wire228 ) | ( n_n4972 ) ;
 assign wire16462 = ( wire21  &  n_n535  &  n_n195 ) | ( wire11  &  n_n535  &  n_n195 ) ;
 assign wire16463 = ( wire18  &  n_n522  &  n_n535 ) | ( wire18  &  n_n526  &  n_n535 ) ;
 assign wire16465 = ( n_n4953 ) | ( wire14752 ) | ( wire16463 ) ;
 assign wire16466 = ( wire250 ) | ( wire16462 ) | ( wire16465 ) ;
 assign wire16468 = ( n_n2222 ) | ( wire16460 ) | ( wire16461 ) | ( wire16466 ) ;
 assign wire16470 = ( n_n2177 ) | ( wire16442 ) | ( wire16443 ) | ( wire16468 ) ;
 assign wire16475 = ( n_n4416 ) | ( n_n4405 ) | ( n_n4406 ) ;
 assign wire16476 = ( n_n4400 ) | ( n_n4389 ) | ( n_n4420 ) | ( n_n4407 ) ;
 assign wire16479 = ( wire13  &  n_n526  &  n_n500 ) | ( wire13  &  n_n500  &  n_n530 ) ;
 assign wire16480 = ( wire13  &  n_n509  &  n_n520 ) | ( wire13  &  n_n509  &  n_n532 ) ;
 assign wire16482 = ( n_n4513 ) | ( n_n4518 ) | ( wire16479 ) ;
 assign wire16483 = ( n_n4484 ) | ( wire199 ) | ( wire16480 ) ;
 assign wire16487 = ( n_n4617 ) | ( n_n4612 ) | ( wire239 ) ;
 assign wire16488 = ( n_n4640 ) | ( n_n4581 ) | ( wire256 ) | ( n_n4623 ) ;
 assign wire16490 = ( wire21  &  n_n473  &  n_n455 ) | ( wire24  &  n_n473  &  n_n455 ) ;
 assign wire16492 = ( n_n4557 ) | ( wire13  &  n_n464  &  n_n526 ) ;
 assign wire16493 = ( n_n4571 ) | ( n_n4523 ) | ( n_n4553 ) ;
 assign wire16494 = ( n_n4521 ) | ( n_n4544 ) | ( wire16490 ) ;
 assign wire16497 = ( wire16482 ) | ( wire16483 ) | ( wire16487 ) | ( wire16488 ) ;
 assign wire16498 = ( wire14  &  n_n522  &  n_n491 ) | ( wire14  &  n_n491  &  n_n530 ) ;
 assign wire16500 = ( wire14  &  n_n509  &  n_n522 ) | ( wire14  &  n_n522  &  n_n535 ) ;
 assign wire16503 = ( n_n4710 ) | ( n_n4719 ) | ( wire16500 ) ;
 assign wire16504 = ( n_n4706 ) | ( n_n4699 ) | ( n_n4687 ) | ( wire16498 ) ;
 assign wire16506 = ( wire21  &  n_n473  &  n_n390 ) | ( wire21  &  n_n390  &  n_n482 ) ;
 assign wire16508 = ( n_n4671 ) | ( n_n4672 ) | ( n_n4685 ) ;
 assign wire16509 = ( n_n4647 ) | ( n_n4656 ) | ( wire16506 ) ;
 assign wire16514 = ( n_n4800 ) | ( n_n4803 ) | ( n_n4783 ) | ( n_n4812 ) ;
 assign wire16516 = ( n_n2130 ) | ( n_n4811 ) | ( n_n4781 ) | ( wire16514 ) ;
 assign wire16518 = ( wire21  &  n_n536  &  n_n473 ) | ( wire22  &  n_n536  &  n_n473 ) ;
 assign wire16520 = ( n_n4414 ) | ( n_n4411 ) | ( n_n4412 ) ;
 assign wire16521 = ( n_n4409 ) | ( n_n4410 ) | ( wire16518 ) ;
 assign wire16526 = ( n_n4440 ) | ( n_n4434 ) | ( wire215 ) ;
 assign wire16527 = ( wire98 ) | ( n_n4430 ) | ( n_n4439 ) | ( n_n4428 ) ;
 assign wire16530 = ( n_n4401 ) | ( n_n4395 ) | ( n_n4402 ) ;
 assign wire16531 = ( n_n4403 ) | ( n_n4392 ) | ( n_n4396 ) | ( n_n4399 ) ;
 assign wire16533 = ( n_n4393 ) | ( n_n4398 ) | ( wire16530 ) | ( wire16531 ) ;
 assign wire16537 = ( n_n4353 ) | ( wire399 ) | ( n_n4354 ) ;
 assign wire16538 = ( n_n4343 ) | ( n_n4352 ) | ( wire67 ) | ( n_n4349 ) ;
 assign wire16539 = ( n_n4317 ) | ( wire16  &  n_n535  &  n_n534 ) ;
 assign wire16544 = ( n_n4336 ) | ( wire171 ) | ( wire198 ) | ( wire283 ) ;
 assign wire16545 = ( n_n2446 ) | ( n_n2443 ) | ( n_n2445 ) | ( wire16539 ) ;
 assign wire16546 = ( wire16537 ) | ( wire16538 ) | ( wire16544 ) ;
 assign wire16548 = ( n_n4356 ) | ( wire345 ) | ( n_n4355 ) ;
 assign wire16549 = ( n_n4363 ) | ( n_n4359 ) | ( n_n4365 ) | ( wire13055 ) ;
 assign wire16551 = ( n_n4372 ) | ( n_n4371 ) | ( n_n4379 ) ;
 assign wire16552 = ( n_n4382 ) | ( n_n4373 ) | ( wire423 ) ;
 assign wire16556 = ( wire16548 ) | ( wire16549 ) | ( wire16551 ) | ( wire16552 ) ;
 assign wire16557 = ( n_n2435 ) | ( wire54 ) | ( wire282 ) | ( wire16556 ) ;
 assign wire16560 = ( wire13  &  n_n535  &  n_n530 ) | ( wire13  &  n_n535  &  n_n532 ) ;
 assign wire16562 = ( n_n4450 ) | ( n_n4445 ) | ( wire368 ) ;
 assign wire16563 = ( n_n4441 ) | ( n_n4448 ) | ( n_n4447 ) | ( wire16560 ) ;
 assign wire16566 = ( n_n4464 ) | ( n_n4463 ) | ( n_n4466 ) ;
 assign wire16567 = ( n_n4467 ) | ( n_n4471 ) | ( n_n4472 ) | ( n_n4468 ) ;
 assign wire16568 = ( n_n4459 ) | ( n_n4470 ) | ( n_n4460 ) | ( n_n4473 ) ;
 assign wire16570 = ( n_n4454 ) | ( wire11520 ) | ( wire14517 ) | ( wire16568 ) ;
 assign wire16571 = ( wire16562 ) | ( wire16563 ) | ( wire16566 ) | ( wire16567 ) ;
 assign wire16572 = ( wire22  &  n_n455  &  n_n500 ) | ( wire24  &  n_n455  &  n_n500 ) ;
 assign wire16573 = ( wire66 ) | ( wire65 ) ;
 assign wire16574 = ( n_n4489 ) | ( n_n4488 ) | ( n_n4490 ) | ( wire16572 ) ;
 assign wire16576 = ( wire184 ) | ( wire70 ) ;
 assign wire16578 = ( wire20  &  n_n455  &  n_n482 ) | ( wire23  &  n_n455  &  n_n482 ) ;
 assign wire16580 = ( wire16578 ) | ( wire416 ) ;
 assign wire16581 = ( n_n4536 ) | ( n_n4532 ) | ( n_n4541 ) | ( wire13090 ) ;
 assign wire16585 = ( n_n4520 ) | ( n_n4529 ) | ( wire724 ) | ( wire789 ) ;
 assign wire16586 = ( wire378 ) | ( wire361 ) ;
 assign wire16587 = ( n_n4512 ) | ( n_n4522 ) | ( n_n4531 ) | ( n_n4517 ) ;
 assign wire16590 = ( n_n4247 ) | ( wire308 ) | ( n_n4528 ) | ( wire16587 ) ;
 assign wire16591 = ( wire16580 ) | ( wire16581 ) | ( wire16585 ) | ( wire16586 ) ;
 assign wire16593 = ( wire13  &  n_n522  &  n_n500 ) | ( wire13  &  n_n500  &  n_n520 ) ;
 assign wire16594 = ( n_n4504 ) | ( n_n4503 ) | ( n_n4506 ) | ( n_n4505 ) ;
 assign wire16596 = ( n_n4508 ) | ( wire13028 ) | ( wire16593 ) | ( wire16594 ) ;
 assign wire16598 = ( n_n2258 ) | ( wire16573 ) | ( wire16574 ) | ( wire16596 ) ;
 assign wire16599 = ( wire16570 ) | ( wire16571 ) | ( wire16590 ) | ( wire16591 ) ;
 assign wire16601 = ( n_n4570 ) | ( n_n4569 ) | ( wire455 ) ;
 assign wire16602 = ( n_n4561 ) | ( n_n4568 ) | ( wire471 ) | ( wire91 ) ;
 assign wire16603 = ( i_9_  &  n_n526  &  n_n535  &  n_n390 ) | ( (~ i_9_)  &  n_n526  &  n_n535  &  n_n390 ) ;
 assign wire16605 = ( wire276 ) | ( wire238 ) ;
 assign wire16606 = ( n_n4584 ) | ( n_n4583 ) | ( n_n4580 ) | ( wire16603 ) ;
 assign wire16609 = ( wire10  &  n_n509  &  n_n526 ) | ( wire10  &  n_n509  &  n_n520 ) ;
 assign wire16611 = ( n_n4616 ) | ( n_n4607 ) | ( n_n4618 ) | ( n_n4611 ) ;
 assign wire16612 = ( n_n4613 ) | ( n_n4610 ) | ( n_n4609 ) | ( wire16609 ) ;
 assign wire16617 = ( n_n4598 ) | ( n_n4601 ) | ( n_n4594 ) | ( n_n4606 ) ;
 assign wire16618 = ( n_n4605 ) | ( n_n4600 ) | ( n_n4603 ) | ( wire255 ) ;
 assign wire16621 = ( n_n4593 ) | ( n_n4590 ) | ( n_n4585 ) | ( wire12520 ) ;
 assign wire16622 = ( wire365 ) | ( n_n4591 ) | ( n_n4592 ) | ( wire16621 ) ;
 assign wire16623 = ( wire16611 ) | ( wire16612 ) | ( wire16617 ) | ( wire16618 ) ;
 assign wire16627 = ( n_n4648 ) | ( n_n4646 ) | ( wire311 ) ;
 assign wire16628 = ( wire309 ) | ( n_n4644 ) | ( n_n4651 ) | ( n_n4649 ) ;
 assign wire16629 = ( wire10  &  n_n522  &  n_n500 ) | ( wire10  &  n_n500  &  n_n530 ) ;
 assign wire16631 = ( n_n4629 ) | ( n_n4630 ) | ( wire190 ) ;
 assign wire16632 = ( wire118 ) | ( n_n4626 ) | ( wire16629 ) ;
 assign wire16633 = ( wire22  &  n_n491  &  n_n390 ) | ( wire25  &  n_n491  &  n_n390 ) ;
 assign wire16635 = ( n_n4637 ) | ( n_n4634 ) | ( n_n4638 ) | ( n_n4631 ) ;
 assign wire16636 = ( n_n4639 ) | ( n_n4635 ) | ( n_n4642 ) | ( wire16633 ) ;
 assign wire16637 = ( wire16636 ) | ( wire16635 ) ;
 assign wire16638 = ( wire16627 ) | ( wire16628 ) | ( wire16631 ) | ( wire16632 ) ;
 assign wire16641 = ( wire213 ) | ( n_n4551 ) | ( n_n4552 ) ;
 assign wire16642 = ( n_n4554 ) | ( n_n4546 ) | ( n_n4555 ) | ( wire212 ) ;
 assign wire16644 = ( wire16601 ) | ( wire16602 ) | ( wire16605 ) | ( wire16606 ) ;
 assign wire16645 = ( wire16641 ) | ( wire16642 ) | ( wire16644 ) ;
 assign wire16646 = ( wire16622 ) | ( wire16623 ) | ( wire16637 ) | ( wire16638 ) ;
 assign wire16650 = ( n_n4341 ) | ( n_n4357 ) | ( n_n4358 ) ;
 assign wire16651 = ( n_n4338 ) | ( n_n4325 ) | ( n_n4380 ) | ( n_n4345 ) ;
 assign wire16656 = ( wire148 ) | ( n_n5318 ) | ( n_n5320 ) ;
 assign wire16657 = ( n_n5321 ) | ( n_n5307 ) | ( wire269 ) ;
 assign wire16658 = ( n_n5326 ) | ( n_n5325 ) | ( n_n5332 ) | ( n_n5329 ) ;
 assign wire16661 = ( wire117 ) | ( n_n5302 ) | ( n_n5306 ) | ( wire12969 ) ;
 assign wire16662 = ( n_n2274 ) | ( wire16656 ) | ( wire16657 ) | ( wire16658 ) ;
 assign wire16663 = ( wire12  &  n_n526  &  n_n491 ) | ( wire12  &  n_n491  &  n_n520 ) ;
 assign wire16665 = ( wire125 ) | ( wire358 ) ;
 assign wire16666 = ( wire76 ) | ( n_n5140 ) | ( wire16663 ) ;
 assign wire16669 = ( wire332 ) | ( wire44 ) ;
 assign wire16670 = ( n_n5171 ) | ( wire114 ) | ( n_n5181 ) | ( n_n5177 ) ;
 assign wire16673 = ( n_n5191 ) | ( wire113 ) | ( n_n5192 ) ;
 assign wire16674 = ( n_n5183 ) | ( wire112 ) | ( n_n5190 ) | ( n_n5188 ) ;
 assign wire16676 = ( wire24  &  n_n464  &  n_n130 ) | ( wire15  &  n_n464  &  n_n130 ) ;
 assign wire16677 = ( wire454 ) | ( wire220 ) ;
 assign wire16678 = ( n_n5201 ) | ( wire451 ) | ( wire761 ) ;
 assign wire16679 = ( n_n5212 ) | ( n_n5203 ) | ( wire16676 ) ;
 assign wire16682 = ( n_n5215 ) | ( n_n2291 ) | ( wire13350 ) | ( wire16679 ) ;
 assign wire16683 = ( wire16673 ) | ( wire16674 ) | ( wire16677 ) | ( wire16678 ) ;
 assign wire16685 = ( n_n5245 ) | ( n_n5241 ) | ( n_n5242 ) ;
 assign wire16686 = ( n_n5239 ) | ( n_n5240 ) | ( wire318 ) ;
 assign wire16690 = ( i_9_  &  n_n524  &  n_n518  &  n_n65 ) | ( (~ i_9_)  &  n_n524  &  n_n518  &  n_n65 ) ;
 assign wire16691 = ( wire181 ) | ( wire62 ) ;
 assign wire16692 = ( n_n5232 ) | ( n_n5237 ) | ( wire183 ) ;
 assign wire16693 = ( n_n5260 ) | ( n_n5226 ) | ( wire16690 ) ;
 assign wire16696 = ( n_n5251 ) | ( wire435 ) | ( n_n1139 ) | ( wire16693 ) ;
 assign wire16698 = ( wire12  &  n_n528  &  n_n482 ) | ( wire12  &  n_n482  &  n_n532 ) ;
 assign wire16699 = ( wire22  &  n_n482  &  n_n130 ) | ( wire24  &  n_n482  &  n_n130 ) ;
 assign wire16702 = ( wire33 ) | ( n_n5170 ) | ( wire16699 ) ;
 assign wire16704 = ( wire16665 ) | ( wire16666 ) | ( wire16669 ) | ( wire16670 ) ;
 assign wire16705 = ( wire168 ) | ( wire16698 ) | ( wire16702 ) | ( wire16704 ) ;
 assign wire16709 = ( n_n5066 ) | ( n_n5063 ) | ( n_n5068 ) ;
 assign wire16710 = ( wire159 ) | ( wire123 ) ;
 assign wire16711 = ( n_n5081 ) | ( n_n5087 ) | ( n_n5064 ) | ( n_n5082 ) ;
 assign wire16715 = ( n_n4152 ) | ( n_n5079 ) | ( n_n5083 ) | ( wire144 ) ;
 assign wire16716 = ( wire90 ) | ( wire16709 ) | ( wire16710 ) | ( wire16711 ) ;
 assign wire16717 = ( wire12  &  n_n530  &  n_n518 ) | ( wire12  &  n_n534  &  n_n518 ) ;
 assign wire16718 = ( n_n5098 ) | ( wire289 ) | ( n_n5095 ) ;
 assign wire16719 = ( n_n5109 ) | ( n_n5107 ) | ( n_n5108 ) | ( wire16717 ) ;
 assign wire16721 = ( wire12  &  n_n509  &  n_n530 ) | ( wire12  &  n_n509  &  n_n532 ) ;
 assign wire16723 = ( n_n5111 ) | ( n_n5113 ) | ( wire414 ) ;
 assign wire16724 = ( n_n5112 ) | ( n_n5110 ) | ( n_n5115 ) | ( wire16721 ) ;
 assign wire16728 = ( n_n5136 ) | ( n_n5127 ) | ( n_n5128 ) | ( n_n5135 ) ;
 assign wire16730 = ( n_n5139 ) | ( n_n5125 ) | ( n_n2304 ) | ( wire16728 ) ;
 assign wire16731 = ( wire16718 ) | ( wire16719 ) | ( wire16723 ) | ( wire16724 ) ;
 assign wire16733 = ( n_n5059 ) | ( n_n5057 ) | ( n_n5058 ) ;
 assign wire16734 = ( wire166 ) | ( n_n5061 ) | ( wire669 ) ;
 assign wire16739 = ( n_n5050 ) | ( n_n5049 ) | ( n_n5043 ) | ( n_n5044 ) ;
 assign wire16740 = ( n_n5040 ) | ( n_n5048 ) | ( n_n5036 ) | ( n_n5047 ) ;
 assign wire16742 = ( n_n5039 ) | ( n_n5029 ) | ( wire16739 ) | ( wire16740 ) ;
 assign wire16744 = ( n_n2214 ) | ( wire14661 ) | ( wire14662 ) | ( wire16742 ) ;
 assign wire16745 = ( wire16715 ) | ( wire16716 ) | ( wire16730 ) | ( wire16731 ) ;
 assign wire16748 = ( n_n5295 ) | ( n_n5291 ) | ( n_n5292 ) ;
 assign wire16749 = ( n_n5293 ) | ( n_n5296 ) | ( n_n5297 ) | ( n_n5298 ) ;
 assign wire16753 = ( wire205 ) | ( wire203 ) ;
 assign wire16754 = ( n_n5270 ) | ( n_n5269 ) | ( wire438 ) ;
 assign wire16755 = ( n_n5274 ) | ( n_n5266 ) | ( n_n5275 ) | ( n_n5261 ) ;
 assign wire16758 = ( n_n5285 ) | ( n_n2651 ) | ( wire14542 ) | ( wire16755 ) ;
 assign wire16760 = ( i_9_  &  n_n464  &  n_n520  &  n_n65 ) | ( (~ i_9_)  &  n_n464  &  n_n520  &  n_n65 ) ;
 assign wire16761 = ( wire16760 ) | ( wire20  &  n_n464  &  n_n65 ) ;
 assign wire16763 = ( n_n2168 ) | ( wire16661 ) | ( wire16662 ) | ( wire16761 ) ;
 assign wire16769 = ( n_n4432 ) | ( n_n4461 ) | ( n_n4438 ) | ( n_n4421 ) ;
 assign wire16770 = ( wire84 ) | ( n_n4465 ) | ( n_n4443 ) | ( n_n4429 ) ;
 assign wire16773 = ( wire22  &  n_n509  &  n_n65 ) | ( wire22  &  n_n518  &  n_n65 ) ;
 assign wire16774 = ( n_n5236 ) | ( wire19  &  n_n528  &  n_n500 ) ;
 assign wire16775 = ( n_n5278 ) | ( n_n5290 ) | ( n_n5289 ) ;
 assign wire16776 = ( n_n5206 ) | ( n_n5223 ) | ( wire449 ) ;
 assign wire16777 = ( n_n5328 ) | ( n_n5254 ) | ( wire16773 ) ;
 assign wire16784 = ( n_n4902 ) | ( n_n4856 ) | ( n_n4894 ) | ( n_n4854 ) ;
 assign wire16785 = ( n_n4905 ) | ( n_n4865 ) | ( n_n4893 ) | ( wire154 ) ;
 assign wire16788 = ( wire12  &  n_n524  &  n_n518 ) | ( wire12  &  n_n526  &  n_n518 ) ;
 assign wire16790 = ( n_n5034 ) | ( n_n5099 ) | ( n_n5097 ) | ( n_n5019 ) ;
 assign wire16791 = ( n_n5117 ) | ( n_n5121 ) | ( n_n5122 ) | ( wire16788 ) ;
 assign wire16795 = ( n_n5142 ) | ( n_n5168 ) | ( wire679 ) ;
 assign wire16796 = ( n_n5123 ) | ( n_n5131 ) | ( n_n5137 ) | ( n_n5146 ) ;
 assign wire16798 = ( wire11  &  n_n509  &  n_n195 ) | ( wire11  &  n_n518  &  n_n195 ) ;
 assign wire16799 = ( wire18  &  n_n509  &  n_n522 ) | ( wire18  &  n_n509  &  n_n526 ) ;
 assign wire16804 = ( n_n5000 ) | ( n_n4957 ) | ( n_n4973 ) | ( wire16798 ) ;
 assign wire16805 = ( n_n4981 ) | ( n_n5005 ) | ( wire16799 ) | ( wire16804 ) ;
 assign wire16811 = ( n_n4847 ) | ( n_n4817 ) | ( wire85 ) ;
 assign wire16812 = ( n_n4827 ) | ( n_n4816 ) | ( n_n4833 ) | ( n_n4813 ) ;
 assign wire16818 = ( n_n4934 ) | ( n_n4938 ) | ( n_n4947 ) | ( n_n4940 ) ;
 assign wire16819 = ( n_n4931 ) | ( n_n4944 ) | ( n_n4932 ) | ( wire340 ) ;
 assign wire16820 = ( wire16819 ) | ( wire16818 ) ;
 assign wire16823 = ( n_n2083 ) | ( n_n2095 ) | ( n_n2096 ) | ( wire16820 ) ;
 assign wire16825 = ( n_n2104 ) | ( n_n2105 ) | ( wire16769 ) | ( wire16770 ) ;
 assign wire16827 = ( n_n2084 ) | ( wire16823 ) | ( wire16825 ) ;
 assign wire16829 = ( wire16598 ) | ( wire16599 ) | ( wire16645 ) | ( wire16646 ) ;
 assign wire16830 = ( n_n2087 ) | ( n_n2086 ) | ( n_n2166 ) | ( wire16827 ) ;
 assign wire16831 = ( n_n2162 ) | ( n_n2163 ) | ( wire16470 ) | ( wire16829 ) ;


endmodule

