module tseng (
	tin_pv10_4_4_, tin_pv11_4_4_, tin_pv6_7_7_, tin_pv2_0_0_, tin_pv10_3_3_, tin_pv1_2_2_, tin_pv11_3_3_, tin_pv4_3_3_, 
	tin_pv10_2_2_, tin_pv11_2_2_, tin_pv6_0_0_, tin_pv2_1_1_, tin_pv10_1_1_, tin_pv1_3_3_, preset_0_0_, tin_pv11_1_1_, tin_pv4_4_4_, tin_pready_0_0_, 
	tin_pv10_0_0_, tin_pv11_0_0_, tin_pv6_1_1_, tin_pv2_2_2_, tin_pv1_4_4_, tin_pv4_5_5_, tin_pv6_2_2_, tin_pv2_3_3_, tin_pv1_5_5_, tin_pv4_6_6_, 
	tin_pv6_3_3_, tin_pv2_4_4_, tin_pv1_6_6_, pclk, tin_pv4_7_7_, tin_pv6_4_4_, tin_pv2_5_5_, tin_pv1_7_7_, tin_pv4_0_0_, tin_pv6_5_5_, 
	tin_pv2_6_6_, tin_pv10_7_7_, tin_pv1_0_0_, tin_pv11_7_7_, tin_pv4_1_1_, tin_pv10_6_6_, tin_pv11_6_6_, tin_pv6_6_6_, tin_pv2_7_7_, preset, 
	tin_pv10_5_5_, tin_pv1_1_1_, tin_pv11_5_5_, tin_pv4_2_2_, pv14_2_2_, pv12_3_3_, pv10_4_4_, pv7_5_5_, pv3_6_6_, pv15_2_2_, 
	pv13_3_3_, pv11_4_4_, pv6_7_7_, pv2_0_0_, pv14_1_1_, pv12_2_2_, pv10_3_3_, pv9_0_0_, pv5_1_1_, pv1_2_2_, 
	pv15_1_1_, pv13_2_2_, pv11_3_3_, pv8_2_2_, pv4_3_3_, pv14_0_0_, pv12_1_1_, pv10_2_2_, pv7_6_6_, pv3_7_7_, 
	pv15_0_0_, pv13_1_1_, pv11_2_2_, pv6_0_0_, pv2_1_1_, pv12_0_0_, pv10_1_1_, pv9_1_1_, pv5_2_2_, pv1_3_3_, 
	pv13_0_0_, pv11_1_1_, pv8_3_3_, pv4_4_4_, pready_0_0_, pv10_0_0_, pv7_7_7_, pv3_0_0_, pv11_0_0_, pv6_1_1_, 
	pv2_2_2_, pv9_2_2_, pv5_3_3_, pv1_4_4_, pv8_4_4_, pv4_5_5_, pv7_0_0_, pv3_1_1_, pv6_2_2_, pv2_3_3_, 
	pv9_3_3_, pv5_4_4_, pv1_5_5_, pv8_5_5_, pv4_6_6_, pv7_1_1_, pv3_2_2_, pv6_3_3_, pv2_4_4_, pv9_4_4_, 
	pv5_5_5_, pv1_6_6_, pv8_6_6_, pv4_7_7_, pv7_2_2_, pv3_3_3_, pv6_4_4_, pv2_5_5_, pv14_7_7_, pv9_5_5_, 
	pv5_6_6_, pv1_7_7_, pv15_7_7_, pv8_7_7_, pv4_0_0_, pv14_6_6_, pv12_7_7_, pv7_3_3_, pv3_4_4_, pv15_6_6_, 
	pv13_7_7_, pv6_5_5_, pv2_6_6_, pdn, pv14_5_5_, pv12_6_6_, pv10_7_7_, pv9_6_6_, pv5_7_7_, pv1_0_0_, 
	pv15_5_5_, pv13_6_6_, pv11_7_7_, pv8_0_0_, pv4_1_1_, pv14_4_4_, pv12_5_5_, pv10_6_6_, pv7_4_4_, pv3_5_5_, 
	pv15_4_4_, pv13_5_5_, pv11_6_6_, pv6_6_6_, pv2_7_7_, pv14_3_3_, pv12_4_4_, pv10_5_5_, pv9_7_7_, pv5_0_0_, 
	pv1_1_1_, pv15_3_3_, pv13_4_4_, pv11_5_5_, pv8_1_1_, pv4_2_2_);

input tin_pv10_4_4_;
input tin_pv11_4_4_;
input tin_pv6_7_7_;
input tin_pv2_0_0_;
input tin_pv10_3_3_;
input tin_pv1_2_2_;
input tin_pv11_3_3_;
input tin_pv4_3_3_;
input tin_pv10_2_2_;
input tin_pv11_2_2_;
input tin_pv6_0_0_;
input tin_pv2_1_1_;
input tin_pv10_1_1_;
input tin_pv1_3_3_;
input preset_0_0_;
input tin_pv11_1_1_;
input tin_pv4_4_4_;
input tin_pready_0_0_;
input tin_pv10_0_0_;
input tin_pv11_0_0_;
input tin_pv6_1_1_;
input tin_pv2_2_2_;
input tin_pv1_4_4_;
input tin_pv4_5_5_;
input tin_pv6_2_2_;
input tin_pv2_3_3_;
input tin_pv1_5_5_;
input tin_pv4_6_6_;
input tin_pv6_3_3_;
input tin_pv2_4_4_;
input tin_pv1_6_6_;
input pclk;
input tin_pv4_7_7_;
input tin_pv6_4_4_;
input tin_pv2_5_5_;
input tin_pv1_7_7_;
input tin_pv4_0_0_;
input tin_pv6_5_5_;
input tin_pv2_6_6_;
input tin_pv10_7_7_;
input tin_pv1_0_0_;
input tin_pv11_7_7_;
input tin_pv4_1_1_;
input tin_pv10_6_6_;
input tin_pv11_6_6_;
input tin_pv6_6_6_;
input tin_pv2_7_7_;
input preset;
input tin_pv10_5_5_;
input tin_pv1_1_1_;
input tin_pv11_5_5_;
input tin_pv4_2_2_;
output pv14_2_2_;
output pv12_3_3_;
output pv10_4_4_;
output pv7_5_5_;
output pv3_6_6_;
output pv15_2_2_;
output pv13_3_3_;
output pv11_4_4_;
output pv6_7_7_;
output pv2_0_0_;
output pv14_1_1_;
output pv12_2_2_;
output pv10_3_3_;
output pv9_0_0_;
output pv5_1_1_;
output pv1_2_2_;
output pv15_1_1_;
output pv13_2_2_;
output pv11_3_3_;
output pv8_2_2_;
output pv4_3_3_;
output pv14_0_0_;
output pv12_1_1_;
output pv10_2_2_;
output pv7_6_6_;
output pv3_7_7_;
output pv15_0_0_;
output pv13_1_1_;
output pv11_2_2_;
output pv6_0_0_;
output pv2_1_1_;
output pv12_0_0_;
output pv10_1_1_;
output pv9_1_1_;
output pv5_2_2_;
output pv1_3_3_;
output pv13_0_0_;
output pv11_1_1_;
output pv8_3_3_;
output pv4_4_4_;
output pready_0_0_;
output pv10_0_0_;
output pv7_7_7_;
output pv3_0_0_;
output pv11_0_0_;
output pv6_1_1_;
output pv2_2_2_;
output pv9_2_2_;
output pv5_3_3_;
output pv1_4_4_;
output pv8_4_4_;
output pv4_5_5_;
output pv7_0_0_;
output pv3_1_1_;
output pv6_2_2_;
output pv2_3_3_;
output pv9_3_3_;
output pv5_4_4_;
output pv1_5_5_;
output pv8_5_5_;
output pv4_6_6_;
output pv7_1_1_;
output pv3_2_2_;
output pv6_3_3_;
output pv2_4_4_;
output pv9_4_4_;
output pv5_5_5_;
output pv1_6_6_;
output pv8_6_6_;
output pv4_7_7_;
output pv7_2_2_;
output pv3_3_3_;
output pv6_4_4_;
output pv2_5_5_;
output pv14_7_7_;
output pv9_5_5_;
output pv5_6_6_;
output pv1_7_7_;
output pv15_7_7_;
output pv8_7_7_;
output pv4_0_0_;
output pv14_6_6_;
output pv12_7_7_;
output pv7_3_3_;
output pv3_4_4_;
output pv15_6_6_;
output pv13_7_7_;
output pv6_5_5_;
output pv2_6_6_;
output pdn;
output pv14_5_5_;
output pv12_6_6_;
output pv10_7_7_;
output pv9_6_6_;
output pv5_7_7_;
output pv1_0_0_;
output pv15_5_5_;
output pv13_6_6_;
output pv11_7_7_;
output pv8_0_0_;
output pv4_1_1_;
output pv14_4_4_;
output pv12_5_5_;
output pv10_6_6_;
output pv7_4_4_;
output pv3_5_5_;
output pv15_4_4_;
output pv13_5_5_;
output pv11_6_6_;
output pv6_6_6_;
output pv2_7_7_;
output pv14_3_3_;
output pv12_4_4_;
output pv10_5_5_;
output pv9_7_7_;
output pv5_0_0_;
output pv1_1_1_;
output pv15_3_3_;
output pv13_4_4_;
output pv11_5_5_;
output pv8_1_1_;
output pv4_2_2_;
wire n_n4140;
wire n_n3935;
wire n_n3444;
wire n_n3007;
wire n_n3725;
wire n_n3399;
wire n_n3143;
wire n_n3781;
wire n_n3066;
wire n_n3507;
wire n_n3224;
wire n_n3179;
wire n_n3273;
wire n_n3166;
wire n_n3686;
wire n_n3380;
wire n_n3096;
wire n_n4106;
wire n_n3496;
wire n_n3791;
wire n_n3518;
wire n_n4348;
wire n_n3028;
wire n_n3618;
wire n_n3263;
wire n_n3778;
wire n_n3227;
wire n_n4113;
wire n_n3145;
wire n_n3510;
wire n_n3151;
wire n_n129;
wire n_n4280;
wire n_n3304;
wire n_n3309;
wire n_n3490;
wire n_n3377;
wire n_n3203;
wire n_n3023;
wire n_n4137;
wire n_n3084;
wire n_n3131;
wire n_n4073;
wire n_n3269;
wire n_n3181;
wire n_n3455;
wire n_n3520;
wire n_n3080;
wire n_n3296;
wire n_n3668;
wire n_n4210;
wire n_n3076;
wire n_n3148;
wire n_n3226;
wire n_n3194;
wire n_n3523;
wire n_n3727;
wire n_n3875;
wire n_n3614;
wire n_n3547;
wire n_n3488;
wire n_n3762;
wire n_n3256;
wire n_n124;
wire n_n3515;
wire n_n3016;
wire n_n3168;
wire n_n3011;
wire n_n3373;
wire n_n3371;
wire n_n3343;
wire n_n3018;
wire n_n3077;
wire n_n3312;
wire n_n3410;
wire n_n3230;
wire n_n3395;
wire n_n3431;
wire n_n3605;
wire n_n3732;
wire n_n3063;
wire n_n3913;
wire n_n3119;
wire n_n3220;
wire n_n3172;
wire n_n3070;
wire n_n3112;
wire n_n3241;
wire n_n3117;
wire n_n3375;
wire n_n4088;
wire n_n3043;
wire n_n3625;
wire n_n3027;
wire n_n3110;
wire n_n3320;
wire n_n3442;
wire n_n3214;
wire n_n3751;
wire n_n4170;
wire n_n3982;
wire n_n3589;
wire n_n4109;
wire n_n3941;
wire n_n3575;
wire n_n4128;
wire n_n4186;
wire n_n4283;
wire n_n3022;
wire n_n3437;
wire n_n3566;
wire n_n3032;
wire n_n3074;
wire n_n3353;
wire n_n3464;
wire n_n4321;
wire n_n3616;
wire n_n4161;
wire n_n3206;
wire n_n4119;
wire n_n3064;
wire n_n4004;
wire n_n3265;
wire n_n3216;
wire n_n3599;
wire n_n3414;
wire n_n4242;
wire n_n3871;
wire n_n3647;
wire n_n3357;
wire n_n3349;
wire n_n3675;
wire n_n3115;
wire n_n3582;
wire n_n3904;
wire n_n4130;
wire n_n3314;
wire n_n3060;
wire n_n3047;
wire n_n3837;
wire n_n3508;
wire n_n3127;
wire n_n3235;
wire n_n4212;
wire n_n3759;
wire n_n4218;
wire n_n3251;
wire n_n3382;
wire n_n3327;
wire n_n3987;
wire n_n3347;
wire n_n3543;
wire n_n3100;
wire n_n4276;
wire n_n3895;
wire n_n3735;
wire n_n3049;
wire n_n3649;
wire n_n3306;
wire n_n4293;
wire n_n3907;
wire n_n3579;
wire n_n4163;
wire n_n3154;
wire n_n3748;
wire n_n3271;
wire n_n4346;
wire n_n3825;
wire n_n3359;
wire n_n3147;
wire n_n3092;
wire n_n3156;
wire n_n3505;
wire n_n3160;
wire n_n3318;
wire n_n3428;
wire n_n3969;
wire n_n3447;
wire n_n4081;
wire n_n3302;
wire n_n3182;
wire n_n3129;
wire n_n3430;
wire n_n4046;
wire n_n3123;
wire n_n3238;
wire n_n3972;
wire n_n3889;
wire n_n4001;
wire n_n3090;
wire n_n3983;
wire n_n3325;
wire n_n3540;
wire n_n125;
wire n_n3693;
wire n_n4373;
wire n_n3866;
wire n_n4289;
wire n_n3459;
wire n_n4121;
wire n_n3773;
wire n_n3013;
wire n_n4239;
wire n_n3950;
wire n_n3236;
wire n_n3530;
wire n_n3033;
wire n_n3550;
wire n_n3378;
wire n_n3009;
wire n_n3569;
wire n_n3853;
wire n_n131;
wire n_n3450;
wire n_n4036;
wire n_n3406;
wire n_n4228;
wire n_n3701;
wire n_n3338;
wire n_n4361;
wire n_n3466;
wire n_n3355;
wire n_n4184;
wire n_n3068;
wire n_n3642;
wire n_n3402;
wire n_n3056;
wire n_n3019;
wire n_n3827;
wire n_n3629;
wire n_n3137;
wire n_n126;
wire n_n4063;
wire n_n3677;
wire n_n3285;
wire n_n3308;
wire n_n4058;
wire n_n3435;
wire n_n3635;
wire n_n3460;
wire n_n4011;
wire n_n3050;
wire n_n3072;
wire n_n3775;
wire n_n3199;
wire n_n3025;
wire n_n3058;
wire n_n3258;
wire n_n3503;
wire n_n130;
wire n_n121;
wire n_n3134;
wire n_n4370;
wire n_n4234;
wire n_n3039;
wire n_n3873;
wire n_n3998;
wire n_n3222;
wire n_n3036;
wire n_n3062;
wire n_n3017;
wire n_n3212;
wire n_n3094;
wire n_n3662;
wire n_n3217;
wire n_n3037;
wire n_n3368;
wire n_n3030;
wire n_n3494;
wire n_n3711;
wire n_n3088;
wire n_n3210;
wire n_n3366;
wire n_n3433;
wire n_n3125;
wire n_n4190;
wire n_n4134;
wire n_n3052;
wire n_n3937;
wire n_n3632;
wire n_n4387;
wire n_n127;
wire n_n3902;
wire n_n3684;
wire n_n3046;
wire n_n3817;
wire n_n3374;
wire n_n3462;
wire n_n3174;
wire n_n3054;
wire n_n3200;
wire n_n3383;
wire n_n4076;
wire n_n3141;
wire n_n3289;
wire n_n3552;
wire n_n3821;
wire n_n3721;
wire n_n4307;
wire n_n3229;
wire n_n3021;
wire n_n3835;
wire n_n3469;
wire n_n3329;
wire n_n3881;
wire n_n3031;
wire n_n4156;
wire n_n4086;
wire n_n3045;
wire n_n3189;
wire n_n4028;
wire n_n3041;
wire n_n133;
wire n_n122;
wire n_n3187;
wire n_n4300;
wire n_n3249;
wire n_n3169;
wire n_n3757;
wire n_n3908;
wire n_n3106;
wire n_n3149;
wire n_n4317;
wire n_n4359;
wire n_n4245;
wire n_n4196;
wire n_n3964;
wire n_n3184;
wire n_n3010;
wire n_n3122;
wire n_n3512;
wire n_n3571;
wire n_n4165;
wire n_n3519;
wire n_n3392;
wire n_n4094;
wire n_n3862;
wire n_n3719;
wire n_n3810;
wire n_n3755;
wire n_n3665;
wire n_n3340;
wire n_n3528;
wire n_n4207;
wire n_n3585;
wire n_n3336;
wire n_n3026;
wire n_n4152;
wire n_n128;
wire n_n3232;
wire n_n4262;
wire n_n3412;
wire n_n3015;
wire n_n3526;
wire n_n3440;
wire n_n3140;
wire n_n4339;
wire n_n4100;
wire n_n3275;
wire n_n4178;
wire n_n3877;
wire n_n3538;
wire n_n3680;
wire n_n3104;
wire n_n3484;
wire n_n3473;
wire n_n3673;
wire n_n3592;
wire n_n3607;
wire n_n3292;
wire n_n4017;
wire n_n4352;
wire n_n3796;
wire n_n3737;
wire n_n3644;
wire n_n3059;
wire n_n3535;
wire n_n3804;
wire n_n3086;
wire n_n4104;
wire n_n3261;
wire n_n4124;
wire n_n3813;
wire n_n132;
wire n_n123;
wire wire988;
wire wire896;
wire wire1016;
wire wire992;
wire wire894;
wire wire916;
wire wire934;
wire wire1020;
wire n_n4069;
wire n_n4015;
wire wire1004;
wire wire990;
wire wire1021;
wire wire994;
wire n_n3563;
wire wire1022;
wire wire1002;
wire wire997;
wire wire1006;
wire wire999;
wire nak3_17;
wire n_n4038;
wire n_n3653;
wire wire944;
wire wire1028;
wire n_n4116;
wire n_n3689;
wire wire1014;
wire n_n4158;
wire wire973;
wire wire1041;
wire n_n4079;
wire wire1012;
wire wire1042;
wire n_n3745;
wire nrq1_3;
wire n_n3741;
wire wire982;
wire n_n4256;
wire wire947;
wire n_n4084;
wire n_n4133;
wire nrq3_12;
wire n_n3832;
wire wire1015;
wire wire1063;
wire wire1064;
wire wire1068;
wire wire923;
wire wire1069;
wire n_n4297;
wire n_n4126;
wire wire1070;
wire wire935;
wire n_n3765;
wire n_n4367;
wire wire984;
wire n_n4335;
wire wire899;
wire n_n3786;
wire wire1075;
wire wire1076;
wire n_n3788;
wire n_n4305;
wire n_n3656;
wire n_n3500;
wire wire1078;
wire wire1079;
wire wire1013;
wire nrq3_15;
wire n_n3363;
wire n_n3362;
wire n_n4078;
wire n_n3888;
wire n_n4345;
wire n_n4019;
wire n_n3884;
wire wire1086;
wire n_n4039;
wire n_n3622;
wire n_n3981;
wire wire1088;
wire n_n3294;
wire n_n3334;
wire n_n4296;
wire n_n3324;
wire n_n3243;
wire n_n3830;
wire n_n3869;
wire n_n3205;
wire wire901;
wire n_n3240;
wire n_n4181;
wire wire1094;
wire n_n3870;
wire wire1096;
wire n_n4144;
wire n_n4223;
wire n_n4034;
wire n_n4259;
wire n_n3900;
wire n_n3124;
wire n_n135;
wire n_n4315;
wire wire1104;
wire n_n4096;
wire wire904;
wire n_n3986;
wire n_n3994;
wire n_n3595;
wire n_n4357;
wire wire1109;
wire n_n4268;
wire n_n4006;
wire n_n3848;
wire n_n4098;
wire wire942;
wire wire1110;
wire n_n3852;
wire wire903;
wire n_n4082;
wire nrq3_2;
wire n_n4169;
wire n_n4168;
wire n_n4155;
wire wire905;
wire wire1116;
wire n_n3420;
wire wire902;
wire n_n4231;
wire wire907;
wire n_n3253;
wire wire1119;
wire wire900;
wire n_n3785;
wire n_n4097;
wire wire941;
wire n_n3975;
wire n_n3974;
wire wire1122;
wire n_n4267;
wire n_n3899;
wire wire906;
wire wire1128;
wire wire1129;
wire wire908;
wire n_n4254;
wire n_n3923;
wire wire1137;
wire wire1136;
wire n_n3927;
wire wire914;
wire wire936;
wire wire1155;
wire wire1008;
wire wire1019;
wire wire1034;
wire wire1038;
wire wire1051;
wire wire1062;
wire wire1082;
wire wire911;
wire wire921;
wire wire922;
wire wire937;
wire wire946;
wire wire971;
wire wire974;
wire wire976;
wire wire978;
wire wire983;
wire wire1165;
wire wire1166;
wire wire1167;
wire wire1168;
wire wire1171;
wire wire1172;
wire wire1173;
wire wire1179;
wire wire1182;
wire wire1184;
wire wire1187;
wire wire1189;
wire wire1191;
wire wire1195;
wire wire1199;
wire wire1201;
wire wire1204;
wire wire1206;
wire wire1208;
wire wire1212;
wire wire1213;
wire wire1214;
wire wire1218;
wire wire1225;
wire wire1230;
wire wire1232;
wire wire1242;
wire wire1246;
wire wire1248;
wire wire1251;
wire wire1259;
wire wire1260;
wire wire1261;
wire wire1263;
wire wire1265;
wire wire1267;
wire wire1270;
wire wire1271;
wire wire1275;
wire wire1280;
wire wire1282;
wire wire1283;
wire wire1285;
wire wire1287;
wire wire1291;
wire wire1295;
wire wire1298;
wire wire1301;
wire wire1303;
wire wire1307;
wire wire1312;
wire wire1315;
wire wire1316;
wire wire1318;
wire wire1323;
wire wire1325;
wire wire1329;
wire wire1333;
wire wire1335;
wire wire1339;
wire wire1341;
wire wire1347;
wire wire1351;
wire wire1355;
wire wire1357;
wire wire1360;
wire wire1362;
wire wire1363;
wire wire1365;
wire wire1375;
wire wire1378;
wire wire1381;
wire wire1385;
wire wire1387;
wire wire1391;
wire wire1392;
wire wire1393;
wire wire1400;
wire wire1402;
wire wire1412;
wire wire1414;
wire wire1416;
wire wire1425;
wire wire1427;
wire wire1429;
wire wire1433;
wire wire1437;
wire wire1447;
wire wire1449;
wire wire1451;
wire wire1455;
wire wire1463;
wire wire1465;
wire wire1468;
wire wire1470;
wire wire1472;
wire wire1477;
wire wire1482;
wire wire1486;
wire wire1487;
wire wire1488;
wire wire1492;
wire wire1494;
wire wire1497;
wire wire1500;
wire wire1504;
wire wire1508;
wire wire1509;
wire wire1510;
wire wire1513;
wire wire1514;
wire wire1518;
wire wire1520;
wire wire1524;
wire wire1527;
wire wire1529;
wire wire1534;
wire wire1538;
wire wire1539;
wire wire1541;
wire wire1547;
wire wire1551;
wire wire1552;
wire wire1557;
wire wire1561;
wire wire1565;
wire wire1574;
wire wire1580;
wire wire1582;
wire wire1584;
wire wire1586;
wire wire1588;
wire wire1594;
wire wire1598;
wire wire1602;
wire wire1604;
wire wire1612;
wire wire1613;
wire wire1614;
wire wire1621;
wire wire1623;
wire wire1630;
wire wire1632;
wire wire1633;
wire wire1638;
wire wire1640;
wire wire1642;
wire wire1647;
wire wire1648;
wire wire1655;
wire wire1659;
wire wire1671;
wire wire1673;
wire wire1679;
wire wire1683;
wire wire1686;
wire wire1687;
wire wire1689;
wire wire1693;
wire wire1699;
wire wire1707;
wire wire1708;
wire wire1711;
wire wire1716;
wire wire1719;
wire wire1724;
wire wire1726;
wire wire1728;
wire wire1736;
wire wire1740;
wire wire1742;
wire wire1745;
wire wire1752;
wire wire1753;
wire wire1754;
wire wire1755;
wire wire1767;
wire wire1771;
wire wire1772;
wire wire1773;
wire wire1774;
wire wire1776;
wire wire1780;
wire wire1784;
wire wire1786;
wire wire1788;
wire wire1792;
wire wire1795;
wire wire1800;
wire wire1806;
wire wire1812;
wire wire1825;
wire wire1830;
wire wire1833;
wire wire1837;
wire wire1843;
wire wire1847;
wire wire1849;
wire wire1853;
wire wire1859;
wire wire1868;
wire wire1870;
wire wire1874;
wire wire1876;
wire wire1881;
wire wire1882;
wire wire1884;
wire wire1885;
wire wire1892;
wire wire1893;
wire wire1894;
wire wire1896;
wire wire1898;
wire wire1899;
wire wire1901;
wire wire1903;
wire wire1904;
wire wire1905;
wire wire1908;
wire wire1909;
wire wire1910;
wire wire1912;
wire wire1914;
wire wire1919;
wire wire1921;
wire wire1925;
wire wire1926;
wire wire1927;
wire wire1928;
wire wire1932;
wire wire1940;
wire wire1944;
wire wire1946;
wire wire1949;
wire wire1953;
wire wire1957;
wire wire1961;
wire wire1963;
wire wire1965;
wire wire1969;
wire wire1971;
wire wire1976;
wire wire1980;
wire wire1984;
wire wire1986;
wire wire1990;
wire wire1992;
wire wire1996;
wire wire1998;
wire wire2000;
wire wire2005;
wire wire2007;
wire wire2009;
wire wire2011;
wire wire2023;
wire wire2027;
wire wire2029;
wire wire2035;
wire wire2036;
wire wire2037;
wire wire2039;
wire wire2044;
wire wire2045;
wire wire2046;
wire wire2047;
wire wire2048;
wire wire2049;
wire wire2050;
wire wire2051;
wire wire2060;
wire wire2061;
wire wire2122;
wire wire2126;
wire wire2141;
wire wire2153;
wire wire2162;
wire wire2166;
wire wire2173;
wire wire2174;
wire wire2175;
wire wire2176;
wire wire2177;
wire wire2182;
wire wire2183;
wire wire2184;
wire wire2185;
wire wire2187;
wire wire2188;
wire wire2189;
wire wire2190;
wire wire2191;
wire wire2192;
wire wire2195;
wire wire2198;
wire wire2202;
wire wire2224;
wire wire2226;
wire wire2240;
wire wire2241;
wire wire2242;
wire wire2259;
wire wire2261;
wire wire2262;
wire wire2263;
wire wire2264;
wire wire2270;
wire wire2275;
wire wire6250;
wire wire6251;
wire wire6252;
wire wire6254;
wire wire6255;
wire wire6257;
wire wire6259;
wire wire6265;
wire wire6266;
wire wire6268;
wire wire6270;
wire wire6272;
wire wire6275;
wire wire6278;
wire wire6281;
wire wire6284;
wire wire6287;
wire wire6289;
wire wire6290;
wire wire6291;
wire wire6295;
wire wire6296;
wire wire6299;
wire wire6300;
wire wire6302;
wire wire6303;
wire wire6306;
wire wire6309;
wire wire6310;
wire wire6312;
wire wire6317;
wire wire6318;
wire wire6321;
wire wire6322;
wire wire6324;
wire wire6325;
wire wire6330;
wire wire6332;
wire wire6333;
wire wire6337;
wire wire6338;
wire wire6342;
wire wire6343;
wire wire6346;
wire wire6349;
wire wire6350;
wire wire6354;
wire wire6355;
wire wire6356;
wire wire6357;
wire wire6358;
wire wire6361;
wire wire6366;
wire wire6370;
wire wire6374;
wire wire6376;
wire wire6379;
wire wire6380;
wire wire6385;
wire wire6386;
wire wire6387;
wire wire6389;
reg n_n4142;

reg n_n3936;

reg n_n3574;

reg n_n3008;

reg n_n3726;

reg n_n3604;

reg n_n3144;

reg n_n3782;

reg n_n3067;

reg n_n4258;

reg n_n3225;

reg n_n3180;

reg n_n3274;

reg n_n3475;

reg n_n3687;

reg n_n3381;

reg n_n3098;

reg n_n4108;

reg n_n3497;

reg n_n3793;

reg n_n4316;

reg n_n4349;

reg n_n3029;

reg n_n3619;

reg n_n3264;

reg n_n3780;

reg ndn3_4;

reg n_n4114;

reg n_n3146;

reg n_n3511;

reg n_n3152;

reg n_n3833;

reg n_n4282;

reg n_n3305;

reg n_n4392;

reg n_n4224;

reg n_n3198;

reg n_n3204;

reg n_n3024;

reg n_n4139;

reg ndn3_15;

reg n_n3133;

reg n_n4074;

reg n_n3270;

reg n_n3858;

reg n_n3456;

reg n_n3521;

reg n_n3081;

reg n_n4381;

reg n_n3670;

reg n_n4211;

reg n_n3493;

reg n_n3495;

reg n_n3916;

reg n_n3195;

reg n_n3525;

reg n_n3729;

reg n_n3876;

reg ndn3_5;

reg n_n3549;

reg n_n3489;

reg n_n3764;

reg n_n3281;

reg n_n3707;

reg n_n3517;

reg n_n4160;

reg n_n4222;

reg n_n3012;

reg n_n4071;

reg n_n3372;

reg n_n3344;

reg n_n3688;

reg n_n3079;

reg n_n3313;

reg n_n3411;

reg n_n3231;

reg n_n3396;

reg n_n3432;

reg n_n3606;

reg n_n3733;

reg n_n3556;

reg n_n4040;

reg n_n3120;

reg n_n3221;

reg n_n3173;

reg n_n3851;

reg n_n3113;

reg n_n3242;

reg n_n3118;

reg n_n3376;

reg n_n4089;

reg n_n3044;

reg n_n3627;

reg n_n3035;

reg n_n3111;

reg n_n3321;

reg n_n3443;

reg n_n3215;

reg ndn3_10;

reg n_n4172;

reg nlc1_2;

reg n_n3590;

reg n_n4110;

reg nlc3_3;

reg n_n3576;

reg n_n4129;

reg n_n4189;

reg n_n4286;

reg n_n4383;

reg pdn;

reg n_n3567;

reg n_n3892;

reg n_n3075;

reg n_n3354;

reg n_n3465;

reg ndn3_6;

reg n_n3617;

reg n_n4162;

reg n_n3207;

reg n_n4120;

reg n_n3065;

reg n_n4005;

reg n_n3266;

reg n_n4337;

reg n_n3600;

reg n_n3415;

reg n_n4243;

reg n_n3872;

reg n_n3648;

reg n_n3358;

reg n_n3350;

reg ndn3_7;

reg n_n3116;

reg n_n3583;

reg n_n3906;

reg n_n4131;

reg n_n3316;

reg n_n3061;

reg n_n3048;

reg n_n3886;

reg n_n3919;

reg n_n3128;

reg n_n3995;

reg n_n4213;

reg n_n3761;

reg ndn3_8;

reg n_n3252;

reg n_n4366;

reg n_n3328;

reg n_n3988;

reg n_n3348;

reg n_n3544;

reg n_n3101;

reg n_n4279;

reg n_n3896;

reg n_n3736;

reg n_n4251;

reg n_n3650;

reg n_n3307;

reg n_n4294;

reg n_n4334;

reg n_n3955;

reg n_n4164;

reg n_n3155;

reg n_n3749;

reg n_n4233;

reg n_n4347;

reg n_n3826;

reg n_n3360;

reg n_n3458;

reg n_n3093;

reg n_n3157;

reg n_n3506;

reg n_n3161;

reg n_n3319;

reg n_n3429;

reg n_n3971;

reg n_n3449;

reg n_n4270;

reg n_n4288;

reg n_n3183;

reg n_n3130;

reg nlak4_2;

reg n_n4047;

reg n_n3978;

reg n_n3239;

reg n_n4145;

reg n_n3890;

reg n_n4003;

reg n_n3091;

reg n_n3985;

reg n_n3326;

reg n_n4052;

reg nsr4_2;

reg n_n4099;

reg n_n4375;

reg n_n4067;

reg n_n4290;

reg n_n3898;

reg n_n4122;

reg n_n3774;

reg n_n3014;

reg n_n4241;

reg n_n3952;

reg n_n3237;

reg n_n3968;

reg n_n3922;

reg n_n3551;

reg n_n3379;

reg n_n4275;

reg n_n3570;

reg n_n3854;

reg n_n4057;

reg n_n3451;

reg n_n4037;

reg n_n3408;

reg n_n4229;

reg n_n4201;

reg n_n3339;

reg n_n4362;

reg n_n3483;

reg n_n3557;

reg n_n4185;

reg n_n3069;

reg n_n3643;

reg n_n3404;

reg n_n3057;

reg n_n3020;

reg n_n3828;

reg n_n3631;

reg n_n3138;

reg nsr1_2;

reg n_n4065;

reg n_n3679;

reg n_n3287;

reg n_n4351;

reg n_n4059;

reg n_n3436;

reg nen3_10;

reg n_n3461;

reg n_n4012;

reg n_n3051;

reg n_n3073;

reg n_n3777;

reg n_n3709;

reg n_n3946;

reg n_n3085;

reg n_n3259;

reg n_n3504;

reg n_n4045;

reg n_n3954;

reg n_n3136;

reg n_n4372;

reg n_n4236;

reg n_n3040;

reg n_n3874;

reg n_n3999;

reg n_n3223;

reg ndn1_34;

reg n_n3743;

reg n_n3657;

reg n_n3213;

reg n_n3095;

reg n_n3663;

reg n_n3724;

reg n_n3038;

reg n_n3370;

reg n_n3624;

reg n_n3578;

reg n_n3713;

reg n_n3089;

reg n_n3211;

reg n_n3367;

reg n_n3434;

reg n_n3126;

reg n_n4192;

reg n_n4136;

reg n_n3053;

reg n_n3938;

reg n_n3769;

reg n_n4390;

reg nsr3_17;

reg n_n3903;

reg n_n3658;

reg nrq3_11;

reg n_n3818;

reg n_n3533;

reg n_n3463;

reg n_n3175;

reg n_n3055;

reg n_n3202;

reg n_n3385;

reg n_n4077;

reg n_n3142;

reg n_n3901;

reg n_n3934;

reg n_n3823;

reg n_n3722;

reg n_n4309;

reg n_n4159;

reg n_n4330;

reg n_n3836;

reg n_n3470;

reg n_n3331;

reg n_n3883;

reg n_n4299;

reg n_n4157;

reg ndn3_9;

reg n_n3208;

reg n_n3190;

reg n_n4029;

reg n_n3042;

reg nsr3_14;

reg n_n4151;

reg n_n3188;

reg n_n4303;

reg n_n3250;

reg n_n3170;

reg n_n3758;

reg n_n3910;

reg n_n3108;

reg n_n3150;

reg n_n4320;

reg n_n4360;

reg n_n4247;

reg n_n4199;

reg n_n3966;

reg n_n3766;

reg n_n4021;

reg n_n4062;

reg n_n3514;

reg n_n3572;

reg n_n4166;

reg n_n3976;

reg n_n3394;

reg n_n4095;

reg n_n3863;

reg n_n3720;

reg ngfdn_3;

reg n_n3756;

reg n_n3667;

reg n_n3342;

reg n_n3529;

reg n_n4209;

reg n_n4324;

reg n_n3337;

reg n_n4227;

reg n_n4153;

reg n_n3831;

reg n_n3233;

reg n_n4263;

reg n_n3413;

reg n_n4182;

reg n_n3841;

reg n_n3441;

reg n_n4026;

reg n_n4342;

reg n_n4102;

reg n_n3277;

reg n_n4180;

reg n_n3878;

reg n_n3931;

reg n_n3845;

reg n_n3865;

reg n_n3486;

reg n_n4056;

reg n_n3674;

reg n_n3959;

reg n_n3608;

reg n_n4080;

reg n_n4018;

reg n_n4354;

reg n_n3797;

reg n_n3739;

reg n_n3646;

reg n_n3099;

reg n_n3537;

reg n_n3806;

reg n_n3087;

reg n_n4105;

reg n_n3262;

reg n_n4125;

reg n_n3814;

reg n_n4093;

reg nsr3_3;

always  @(posedge pclk)
	n_n4142<=n_n4140;

 always  @(posedge pclk)
	n_n3936<=n_n3935;

 always  @(posedge pclk)
	n_n3574<=n_n3444;

 always  @(posedge pclk)
	n_n3008<=n_n3007;

 always  @(posedge pclk)
	n_n3726<=n_n3725;

 always  @(posedge pclk)
	n_n3604<=n_n3399;

 always  @(posedge pclk)
	n_n3144<=n_n3143;

 always  @(posedge pclk)
	n_n3782<=n_n3781;

 always  @(posedge pclk)
	n_n3067<=n_n3066;

 always  @(posedge pclk)
	n_n4258<=n_n3507;

 always  @(posedge pclk)
	n_n3225<=n_n3224;

 always  @(posedge pclk)
	n_n3180<=n_n3179;

 always  @(posedge pclk)
	n_n3274<=n_n3273;

 always  @(posedge pclk)
	n_n3475<=n_n3166;

 always  @(posedge pclk)
	n_n3687<=n_n3686;

 always  @(posedge pclk)
	n_n3381<=n_n3380;

 always  @(posedge pclk)
	n_n3098<=n_n3096;

 always  @(posedge pclk)
	n_n4108<=n_n4106;

 always  @(posedge pclk)
	n_n3497<=n_n3496;

 always  @(posedge pclk)
	n_n3793<=n_n3791;

 always  @(posedge pclk)
	n_n4316<=n_n3518;

 always  @(posedge pclk)
	n_n4349<=n_n4348;

 always  @(posedge pclk)
	n_n3029<=n_n3028;

 always  @(posedge pclk)
	n_n3619<=n_n3618;

 always  @(posedge pclk)
	n_n3264<=n_n3263;

 always  @(posedge pclk)
	n_n3780<=n_n3778;

 always  @(posedge pclk)
	ndn3_4<=n_n3227;

 always  @(posedge pclk)
	n_n4114<=n_n4113;

 always  @(posedge pclk)
	n_n3146<=n_n3145;

 always  @(posedge pclk)
	n_n3511<=n_n3510;

 always  @(posedge pclk)
	n_n3152<=n_n3151;

 always  @(posedge pclk)
	n_n3833<=n_n129;

 always  @(posedge pclk)
	n_n4282<=n_n4280;

 always  @(posedge pclk)
	n_n3305<=n_n3304;

 always  @(posedge pclk)
	n_n4392<=n_n3309;

 always  @(posedge pclk)
	n_n4224<=n_n3490;

 always  @(posedge pclk)
	n_n3198<=n_n3377;

 always  @(posedge pclk)
	n_n3204<=n_n3203;

 always  @(posedge pclk)
	n_n3024<=n_n3023;

 always  @(posedge pclk)
	n_n4139<=n_n4137;

 always  @(posedge pclk)
	ndn3_15<=n_n3084;

 always  @(posedge pclk)
	n_n3133<=n_n3131;

 always  @(posedge pclk)
	n_n4074<=n_n4073;

 always  @(posedge pclk)
	n_n3270<=n_n3269;

 always  @(posedge pclk)
	n_n3858<=n_n3181;

 always  @(posedge pclk)
	n_n3456<=n_n3455;

 always  @(posedge pclk)
	n_n3521<=n_n3520;

 always  @(posedge pclk)
	n_n3081<=n_n3080;

 always  @(posedge pclk)
	n_n4381<=n_n3296;

 always  @(posedge pclk)
	n_n3670<=n_n3668;

 always  @(posedge pclk)
	n_n4211<=n_n4210;

 always  @(posedge pclk)
	n_n3493<=n_n3076;

 always  @(posedge pclk)
	n_n3495<=n_n3148;

 always  @(posedge pclk)
	n_n3916<=n_n3226;

 always  @(posedge pclk)
	n_n3195<=n_n3194;

 always  @(posedge pclk)
	n_n3525<=n_n3523;

 always  @(posedge pclk)
	n_n3729<=n_n3727;

 always  @(posedge pclk)
	n_n3876<=n_n3875;

 always  @(posedge pclk)
	ndn3_5<=n_n3614;

 always  @(posedge pclk)
	n_n3549<=n_n3547;

 always  @(posedge pclk)
	n_n3489<=n_n3488;

 always  @(posedge pclk)
	n_n3764<=n_n3762;

 always  @(posedge pclk)
	n_n3281<=n_n3256;

 always  @(posedge pclk)
	n_n3707<=n_n124;

 always  @(posedge pclk)
	n_n3517<=n_n3515;

 always  @(posedge pclk)
	n_n4160<=n_n3016;

 always  @(posedge pclk)
	n_n4222<=n_n3168;

 always  @(posedge pclk)
	n_n3012<=n_n3011;

 always  @(posedge pclk)
	n_n4071<=n_n3373;

 always  @(posedge pclk)
	n_n3372<=n_n3371;

 always  @(posedge pclk)
	n_n3344<=n_n3343;

 always  @(posedge pclk)
	n_n3688<=n_n3018;

 always  @(posedge pclk)
	n_n3079<=n_n3077;

 always  @(posedge pclk)
	n_n3313<=n_n3312;

 always  @(posedge pclk)
	n_n3411<=n_n3410;

 always  @(posedge pclk)
	n_n3231<=n_n3230;

 always  @(posedge pclk)
	n_n3396<=n_n3395;

 always  @(posedge pclk)
	n_n3432<=n_n3431;

 always  @(posedge pclk)
	n_n3606<=n_n3605;

 always  @(posedge pclk)
	n_n3733<=n_n3732;

 always  @(posedge pclk)
	n_n3556<=n_n3063;

 always  @(posedge pclk)
	n_n4040<=n_n3913;

 always  @(posedge pclk)
	n_n3120<=n_n3119;

 always  @(posedge pclk)
	n_n3221<=n_n3220;

 always  @(posedge pclk)
	n_n3173<=n_n3172;

 always  @(posedge pclk)
	n_n3851<=n_n3070;

 always  @(posedge pclk)
	n_n3113<=n_n3112;

 always  @(posedge pclk)
	n_n3242<=n_n3241;

 always  @(posedge pclk)
	n_n3118<=n_n3117;

 always  @(posedge pclk)
	n_n3376<=n_n3375;

 always  @(posedge pclk)
	n_n4089<=n_n4088;

 always  @(posedge pclk)
	n_n3044<=n_n3043;

 always  @(posedge pclk)
	n_n3627<=n_n3625;

 always  @(posedge pclk)
	n_n3035<=n_n3027;

 always  @(posedge pclk)
	n_n3111<=n_n3110;

 always  @(posedge pclk)
	n_n3321<=n_n3320;

 always  @(posedge pclk)
	n_n3443<=n_n3442;

 always  @(posedge pclk)
	n_n3215<=n_n3214;

 always  @(posedge pclk)
	ndn3_10<=n_n3751;

 always  @(posedge pclk)
	n_n4172<=n_n4170;

 always  @(posedge pclk)
	nlc1_2<=n_n3982;

 always  @(posedge pclk)
	n_n3590<=n_n3589;

 always  @(posedge pclk)
	n_n4110<=n_n4109;

 always  @(posedge pclk)
	nlc3_3<=n_n3941;

 always  @(posedge pclk)
	n_n3576<=n_n3575;

 always  @(posedge pclk)
	n_n4129<=n_n4128;

 always  @(posedge pclk)
	n_n4189<=n_n4186;

 always  @(posedge pclk)
	n_n4286<=n_n4283;

 always  @(posedge pclk)
	n_n4383<=n_n3022;

 always  @(posedge pclk)
	pdn<=n_n3437;

 always  @(posedge pclk)
	n_n3567<=n_n3566;

 always  @(posedge pclk)
	n_n3892<=n_n3032;

 always  @(posedge pclk)
	n_n3075<=n_n3074;

 always  @(posedge pclk)
	n_n3354<=n_n3353;

 always  @(posedge pclk)
	n_n3465<=n_n3464;

 always  @(posedge pclk)
	ndn3_6<=n_n4321;

 always  @(posedge pclk)
	n_n3617<=n_n3616;

 always  @(posedge pclk)
	n_n4162<=n_n4161;

 always  @(posedge pclk)
	n_n3207<=n_n3206;

 always  @(posedge pclk)
	n_n4120<=n_n4119;

 always  @(posedge pclk)
	n_n3065<=n_n3064;

 always  @(posedge pclk)
	n_n4005<=n_n4004;

 always  @(posedge pclk)
	n_n3266<=n_n3265;

 always  @(posedge pclk)
	n_n4337<=n_n3216;

 always  @(posedge pclk)
	n_n3600<=n_n3599;

 always  @(posedge pclk)
	n_n3415<=n_n3414;

 always  @(posedge pclk)
	n_n4243<=n_n4242;

 always  @(posedge pclk)
	n_n3872<=n_n3871;

 always  @(posedge pclk)
	n_n3648<=n_n3647;

 always  @(posedge pclk)
	n_n3358<=n_n3357;

 always  @(posedge pclk)
	n_n3350<=n_n3349;

 always  @(posedge pclk)
	ndn3_7<=n_n3675;

 always  @(posedge pclk)
	n_n3116<=n_n3115;

 always  @(posedge pclk)
	n_n3583<=n_n3582;

 always  @(posedge pclk)
	n_n3906<=n_n3904;

 always  @(posedge pclk)
	n_n4131<=n_n4130;

 always  @(posedge pclk)
	n_n3316<=n_n3314;

 always  @(posedge pclk)
	n_n3061<=n_n3060;

 always  @(posedge pclk)
	n_n3048<=n_n3047;

 always  @(posedge pclk)
	n_n3886<=n_n3837;

 always  @(posedge pclk)
	n_n3919<=n_n3508;

 always  @(posedge pclk)
	n_n3128<=n_n3127;

 always  @(posedge pclk)
	n_n3995<=n_n3235;

 always  @(posedge pclk)
	n_n4213<=n_n4212;

 always  @(posedge pclk)
	n_n3761<=n_n3759;

 always  @(posedge pclk)
	ndn3_8<=n_n4218;

 always  @(posedge pclk)
	n_n3252<=n_n3251;

 always  @(posedge pclk)
	n_n4366<=n_n3382;

 always  @(posedge pclk)
	n_n3328<=n_n3327;

 always  @(posedge pclk)
	n_n3988<=n_n3987;

 always  @(posedge pclk)
	n_n3348<=n_n3347;

 always  @(posedge pclk)
	n_n3544<=n_n3543;

 always  @(posedge pclk)
	n_n3101<=n_n3100;

 always  @(posedge pclk)
	n_n4279<=n_n4276;

 always  @(posedge pclk)
	n_n3896<=n_n3895;

 always  @(posedge pclk)
	n_n3736<=n_n3735;

 always  @(posedge pclk)
	n_n4251<=n_n3049;

 always  @(posedge pclk)
	n_n3650<=n_n3649;

 always  @(posedge pclk)
	n_n3307<=n_n3306;

 always  @(posedge pclk)
	n_n4294<=n_n4293;

 always  @(posedge pclk)
	n_n4334<=n_n3907;

 always  @(posedge pclk)
	n_n3955<=n_n3579;

 always  @(posedge pclk)
	n_n4164<=n_n4163;

 always  @(posedge pclk)
	n_n3155<=n_n3154;

 always  @(posedge pclk)
	n_n3749<=n_n3748;

 always  @(posedge pclk)
	n_n4233<=n_n3271;

 always  @(posedge pclk)
	n_n4347<=n_n4346;

 always  @(posedge pclk)
	n_n3826<=n_n3825;

 always  @(posedge pclk)
	n_n3360<=n_n3359;

 always  @(posedge pclk)
	n_n3458<=n_n3147;

 always  @(posedge pclk)
	n_n3093<=n_n3092;

 always  @(posedge pclk)
	n_n3157<=n_n3156;

 always  @(posedge pclk)
	n_n3506<=n_n3505;

 always  @(posedge pclk)
	n_n3161<=n_n3160;

 always  @(posedge pclk)
	n_n3319<=n_n3318;

 always  @(posedge pclk)
	n_n3429<=n_n3428;

 always  @(posedge pclk)
	n_n3971<=n_n3969;

 always  @(posedge pclk)
	n_n3449<=n_n3447;

 always  @(posedge pclk)
	n_n4270<=n_n4081;

 always  @(posedge pclk)
	n_n4288<=n_n3302;

 always  @(posedge pclk)
	n_n3183<=n_n3182;

 always  @(posedge pclk)
	n_n3130<=n_n3129;

 always  @(posedge pclk)
	nlak4_2<=n_n3430;

 always  @(posedge pclk)
	n_n4047<=n_n4046;

 always  @(posedge pclk)
	n_n3978<=n_n3123;

 always  @(posedge pclk)
	n_n3239<=n_n3238;

 always  @(posedge pclk)
	n_n4145<=n_n3972;

 always  @(posedge pclk)
	n_n3890<=n_n3889;

 always  @(posedge pclk)
	n_n4003<=n_n4001;

 always  @(posedge pclk)
	n_n3091<=n_n3090;

 always  @(posedge pclk)
	n_n3985<=n_n3983;

 always  @(posedge pclk)
	n_n3326<=n_n3325;

 always  @(posedge pclk)
	n_n4052<=n_n3540;

 always  @(posedge pclk)
	nsr4_2<=n_n125;

 always  @(posedge pclk)
	n_n4099<=n_n3693;

 always  @(posedge pclk)
	n_n4375<=n_n4373;

 always  @(posedge pclk)
	n_n4067<=n_n3866;

 always  @(posedge pclk)
	n_n4290<=n_n4289;

 always  @(posedge pclk)
	n_n3898<=n_n3459;

 always  @(posedge pclk)
	n_n4122<=n_n4121;

 always  @(posedge pclk)
	n_n3774<=n_n3773;

 always  @(posedge pclk)
	n_n3014<=n_n3013;

 always  @(posedge pclk)
	n_n4241<=n_n4239;

 always  @(posedge pclk)
	n_n3952<=n_n3950;

 always  @(posedge pclk)
	n_n3237<=n_n3236;

 always  @(posedge pclk)
	n_n3968<=n_n3530;

 always  @(posedge pclk)
	n_n3922<=n_n3033;

 always  @(posedge pclk)
	n_n3551<=n_n3550;

 always  @(posedge pclk)
	n_n3379<=n_n3378;

 always  @(posedge pclk)
	n_n4275<=n_n3009;

 always  @(posedge pclk)
	n_n3570<=n_n3569;

 always  @(posedge pclk)
	n_n3854<=n_n3853;

 always  @(posedge pclk)
	n_n4057<=n_n131;

 always  @(posedge pclk)
	n_n3451<=n_n3450;

 always  @(posedge pclk)
	n_n4037<=n_n4036;

 always  @(posedge pclk)
	n_n3408<=n_n3406;

 always  @(posedge pclk)
	n_n4229<=n_n4228;

 always  @(posedge pclk)
	n_n4201<=n_n3701;

 always  @(posedge pclk)
	n_n3339<=n_n3338;

 always  @(posedge pclk)
	n_n4362<=n_n4361;

 always  @(posedge pclk)
	n_n3483<=n_n3466;

 always  @(posedge pclk)
	n_n3557<=n_n3355;

 always  @(posedge pclk)
	n_n4185<=n_n4184;

 always  @(posedge pclk)
	n_n3069<=n_n3068;

 always  @(posedge pclk)
	n_n3643<=n_n3642;

 always  @(posedge pclk)
	n_n3404<=n_n3402;

 always  @(posedge pclk)
	n_n3057<=n_n3056;

 always  @(posedge pclk)
	n_n3020<=n_n3019;

 always  @(posedge pclk)
	n_n3828<=n_n3827;

 always  @(posedge pclk)
	n_n3631<=n_n3629;

 always  @(posedge pclk)
	n_n3138<=n_n3137;

 always  @(posedge pclk)
	nsr1_2<=n_n126;

 always  @(posedge pclk)
	n_n4065<=n_n4063;

 always  @(posedge pclk)
	n_n3679<=n_n3677;

 always  @(posedge pclk)
	n_n3287<=n_n3285;

 always  @(posedge pclk)
	n_n4351<=n_n3308;

 always  @(posedge pclk)
	n_n4059<=n_n4058;

 always  @(posedge pclk)
	n_n3436<=n_n3435;

 always  @(posedge pclk)
	nen3_10<=n_n3635;

 always  @(posedge pclk)
	n_n3461<=n_n3460;

 always  @(posedge pclk)
	n_n4012<=n_n4011;

 always  @(posedge pclk)
	n_n3051<=n_n3050;

 always  @(posedge pclk)
	n_n3073<=n_n3072;

 always  @(posedge pclk)
	n_n3777<=n_n3775;

 always  @(posedge pclk)
	n_n3709<=n_n3199;

 always  @(posedge pclk)
	n_n3946<=n_n3025;

 always  @(posedge pclk)
	n_n3085<=n_n3058;

 always  @(posedge pclk)
	n_n3259<=n_n3258;

 always  @(posedge pclk)
	n_n3504<=n_n3503;

 always  @(posedge pclk)
	n_n4045<=n_n130;

 always  @(posedge pclk)
	n_n3954<=n_n121;

 always  @(posedge pclk)
	n_n3136<=n_n3134;

 always  @(posedge pclk)
	n_n4372<=n_n4370;

 always  @(posedge pclk)
	n_n4236<=n_n4234;

 always  @(posedge pclk)
	n_n3040<=n_n3039;

 always  @(posedge pclk)
	n_n3874<=n_n3873;

 always  @(posedge pclk)
	n_n3999<=n_n3998;

 always  @(posedge pclk)
	n_n3223<=n_n3222;

 always  @(posedge pclk)
	ndn1_34<=n_n3036;

 always  @(posedge pclk)
	n_n3743<=n_n3062;

 always  @(posedge pclk)
	n_n3657<=n_n3017;

 always  @(posedge pclk)
	n_n3213<=n_n3212;

 always  @(posedge pclk)
	n_n3095<=n_n3094;

 always  @(posedge pclk)
	n_n3663<=n_n3662;

 always  @(posedge pclk)
	n_n3724<=n_n3217;

 always  @(posedge pclk)
	n_n3038<=n_n3037;

 always  @(posedge pclk)
	n_n3370<=n_n3368;

 always  @(posedge pclk)
	n_n3624<=n_n3030;

 always  @(posedge pclk)
	n_n3578<=n_n3494;

 always  @(posedge pclk)
	n_n3713<=n_n3711;

 always  @(posedge pclk)
	n_n3089<=n_n3088;

 always  @(posedge pclk)
	n_n3211<=n_n3210;

 always  @(posedge pclk)
	n_n3367<=n_n3366;

 always  @(posedge pclk)
	n_n3434<=n_n3433;

 always  @(posedge pclk)
	n_n3126<=n_n3125;

 always  @(posedge pclk)
	n_n4192<=n_n4190;

 always  @(posedge pclk)
	n_n4136<=n_n4134;

 always  @(posedge pclk)
	n_n3053<=n_n3052;

 always  @(posedge pclk)
	n_n3938<=n_n3937;

 always  @(posedge pclk)
	n_n3769<=n_n3632;

 always  @(posedge pclk)
	n_n4390<=n_n4387;

 always  @(posedge pclk)
	nsr3_17<=n_n127;

 always  @(posedge pclk)
	n_n3903<=n_n3902;

 always  @(posedge pclk)
	n_n3658<=n_n3684;

 always  @(posedge pclk)
	nrq3_11<=n_n3046;

 always  @(posedge pclk)
	n_n3818<=n_n3817;

 always  @(posedge pclk)
	n_n3533<=n_n3374;

 always  @(posedge pclk)
	n_n3463<=n_n3462;

 always  @(posedge pclk)
	n_n3175<=n_n3174;

 always  @(posedge pclk)
	n_n3055<=n_n3054;

 always  @(posedge pclk)
	n_n3202<=n_n3200;

 always  @(posedge pclk)
	n_n3385<=n_n3383;

 always  @(posedge pclk)
	n_n4077<=n_n4076;

 always  @(posedge pclk)
	n_n3142<=n_n3141;

 always  @(posedge pclk)
	n_n3901<=n_n3289;

 always  @(posedge pclk)
	n_n3934<=n_n3552;

 always  @(posedge pclk)
	n_n3823<=n_n3821;

 always  @(posedge pclk)
	n_n3722<=n_n3721;

 always  @(posedge pclk)
	n_n4309<=n_n4307;

 always  @(posedge pclk)
	n_n4159<=n_n3229;

 always  @(posedge pclk)
	n_n4330<=n_n3021;

 always  @(posedge pclk)
	n_n3836<=n_n3835;

 always  @(posedge pclk)
	n_n3470<=n_n3469;

 always  @(posedge pclk)
	n_n3331<=n_n3329;

 always  @(posedge pclk)
	n_n3883<=n_n3881;

 always  @(posedge pclk)
	n_n4299<=n_n3031;

 always  @(posedge pclk)
	n_n4157<=n_n4156;

 always  @(posedge pclk)
	ndn3_9<=n_n4086;

 always  @(posedge pclk)
	n_n3208<=n_n3045;

 always  @(posedge pclk)
	n_n3190<=n_n3189;

 always  @(posedge pclk)
	n_n4029<=n_n4028;

 always  @(posedge pclk)
	n_n3042<=n_n3041;

 always  @(posedge pclk)
	nsr3_14<=n_n133;

 always  @(posedge pclk)
	n_n4151<=n_n122;

 always  @(posedge pclk)
	n_n3188<=n_n3187;

 always  @(posedge pclk)
	n_n4303<=n_n4300;

 always  @(posedge pclk)
	n_n3250<=n_n3249;

 always  @(posedge pclk)
	n_n3170<=n_n3169;

 always  @(posedge pclk)
	n_n3758<=n_n3757;

 always  @(posedge pclk)
	n_n3910<=n_n3908;

 always  @(posedge pclk)
	n_n3108<=n_n3106;

 always  @(posedge pclk)
	n_n3150<=n_n3149;

 always  @(posedge pclk)
	n_n4320<=n_n4317;

 always  @(posedge pclk)
	n_n4360<=n_n4359;

 always  @(posedge pclk)
	n_n4247<=n_n4245;

 always  @(posedge pclk)
	n_n4199<=n_n4196;

 always  @(posedge pclk)
	n_n3966<=n_n3964;

 always  @(posedge pclk)
	n_n3766<=n_n3184;

 always  @(posedge pclk)
	n_n4021<=n_n3010;

 always  @(posedge pclk)
	n_n4062<=n_n3122;

 always  @(posedge pclk)
	n_n3514<=n_n3512;

 always  @(posedge pclk)
	n_n3572<=n_n3571;

 always  @(posedge pclk)
	n_n4166<=n_n4165;

 always  @(posedge pclk)
	n_n3976<=n_n3519;

 always  @(posedge pclk)
	n_n3394<=n_n3392;

 always  @(posedge pclk)
	n_n4095<=n_n4094;

 always  @(posedge pclk)
	n_n3863<=n_n3862;

 always  @(posedge pclk)
	n_n3720<=n_n3719;

 always  @(posedge pclk)
	ngfdn_3<=n_n3810;

 always  @(posedge pclk)
	n_n3756<=n_n3755;

 always  @(posedge pclk)
	n_n3667<=n_n3665;

 always  @(posedge pclk)
	n_n3342<=n_n3340;

 always  @(posedge pclk)
	n_n3529<=n_n3528;

 always  @(posedge pclk)
	n_n4209<=n_n4207;

 always  @(posedge pclk)
	n_n4324<=n_n3585;

 always  @(posedge pclk)
	n_n3337<=n_n3336;

 always  @(posedge pclk)
	n_n4227<=n_n3026;

 always  @(posedge pclk)
	n_n4153<=n_n4152;

 always  @(posedge pclk)
	n_n3831<=n_n128;

 always  @(posedge pclk)
	n_n3233<=n_n3232;

 always  @(posedge pclk)
	n_n4263<=n_n4262;

 always  @(posedge pclk)
	n_n3413<=n_n3412;

 always  @(posedge pclk)
	n_n4182<=n_n3015;

 always  @(posedge pclk)
	n_n3841<=n_n3526;

 always  @(posedge pclk)
	n_n3441<=n_n3440;

 always  @(posedge pclk)
	n_n4026<=n_n3140;

 always  @(posedge pclk)
	n_n4342<=n_n4339;

 always  @(posedge pclk)
	n_n4102<=n_n4100;

 always  @(posedge pclk)
	n_n3277<=n_n3275;

 always  @(posedge pclk)
	n_n4180<=n_n4178;

 always  @(posedge pclk)
	n_n3878<=n_n3877;

 always  @(posedge pclk)
	n_n3931<=n_n3538;

 always  @(posedge pclk)
	n_n3845<=n_n3680;

 always  @(posedge pclk)
	n_n3865<=n_n3104;

 always  @(posedge pclk)
	n_n3486<=n_n3484;

 always  @(posedge pclk)
	n_n4056<=n_n3473;

 always  @(posedge pclk)
	n_n3674<=n_n3673;

 always  @(posedge pclk)
	n_n3959<=n_n3592;

 always  @(posedge pclk)
	n_n3608<=n_n3607;

 always  @(posedge pclk)
	n_n4080<=n_n3292;

 always  @(posedge pclk)
	n_n4018<=n_n4017;

 always  @(posedge pclk)
	n_n4354<=n_n4352;

 always  @(posedge pclk)
	n_n3797<=n_n3796;

 always  @(posedge pclk)
	n_n3739<=n_n3737;

 always  @(posedge pclk)
	n_n3646<=n_n3644;

 always  @(posedge pclk)
	n_n3099<=n_n3059;

 always  @(posedge pclk)
	n_n3537<=n_n3535;

 always  @(posedge pclk)
	n_n3806<=n_n3804;

 always  @(posedge pclk)
	n_n3087<=n_n3086;

 always  @(posedge pclk)
	n_n4105<=n_n4104;

 always  @(posedge pclk)
	n_n3262<=n_n3261;

 always  @(posedge pclk)
	n_n4125<=n_n4124;

 always  @(posedge pclk)
	n_n3814<=n_n3813;

 always  @(posedge pclk)
	n_n4093<=n_n132;

 always  @(posedge pclk)
	nsr3_3<=n_n123;

 assign pv14_2_2_ = ( n_n3358  &  n_n4153 ) ;
 assign pv12_3_3_ = ( n_n3631  &  n_n3367 ) ;
 assign pv10_4_4_ = ( n_n4136  &  n_n3042 ) | ( tin_pv10_4_4_  &  (~ n_n3042) ) ;
 assign pv7_5_5_ = ( n_n3130  &  n_n3679 ) ;
 assign pv3_6_6_ = ( n_n3252  &  n_n3057 ) ;
 assign pv15_2_2_ = ( n_n3113  &  n_n4037 ) ;
 assign pv13_3_3_ = ( n_n3600  &  n_n3404 ) ;
 assign pv11_4_4_ = ( tin_pv11_4_4_  &  (~ n_n4120) ) | ( n_n4120  &  n_n3966 ) ;
 assign pv6_7_7_ = ( tin_pv6_7_7_  &  (~ n_n4164) ) | ( n_n4164  &  n_n3370 ) ;
 assign pv2_0_0_ = ( tin_pv2_0_0_  &  (~ n_n3211) ) | ( n_n3211  &  n_n3910 ) ;
 assign pv14_1_1_ = ( n_n3012  &  n_n3038 ) ;
 assign pv12_2_2_ = ( n_n3067  &  n_n3576 ) ;
 assign pv10_3_3_ = ( tin_pv10_3_3_  &  (~ n_n4129) ) | ( n_n4129  &  n_n3213 ) ;
 assign pv9_0_0_ = ( n_n3128  &  n_n3890 ) ;
 assign pv5_1_1_ = ( n_n3443  &  n_n3287 ) ;
 assign pv1_2_2_ = ( tin_pv1_2_2_  &  (~ n_n3470) ) | ( n_n3470  &  n_n3537 ) ;
 assign pv15_1_1_ = ( n_n3606  &  n_n3108 ) ;
 assign pv13_2_2_ = ( n_n3379  &  n_n3463 ) ;
 assign pv11_3_3_ = ( tin_pv11_3_3_  &  (~ n_n3432) ) | ( n_n3432  &  n_n3583 ) ;
 assign pv8_2_2_ = ( n_n3456  &  n_n3055 ) ;
 assign pv4_3_3_ = ( tin_pv4_3_3_  &  (~ n_n3489) ) | ( n_n3489  &  n_n4309 ) ;
 assign pv14_0_0_ = ( n_n3761  &  n_n3903 ) ;
 assign pv12_1_1_ = ( n_n3264  &  n_n4390 ) ;
 assign pv10_2_2_ = ( n_n3549  &  n_n3065 ) | ( tin_pv10_2_2_  &  (~ n_n3065) ) ;
 assign pv7_6_6_ = ( n_n3670  &  n_n3617 ) ;
 assign pv3_7_7_ = ( n_n3590  &  n_n4102 ) ;
 assign pv15_0_0_ = ( n_n4003  &  n_n3188 ) ;
 assign pv13_1_1_ = ( n_n3221  &  n_n3150 ) ;
 assign pv11_2_2_ = ( tin_pv11_2_2_  &  (~ n_n3152) ) | ( n_n3152  &  n_n3823 ) ;
 assign pv6_0_0_ = ( tin_pv6_0_0_  &  (~ n_n3029) ) | ( n_n3029  &  n_n3506 ) ;
 assign pv2_1_1_ = ( tin_pv2_1_1_  &  (~ n_n3999) ) | ( n_n3999  &  n_n3646 ) ;
 assign pv12_0_0_ = ( n_n3098  &  n_n3339 ) ;
 assign pv10_1_1_ = ( n_n3270  &  n_n3872 ) | ( tin_pv10_1_1_  &  (~ n_n3872) ) ;
 assign pv9_1_1_ = ( n_n3024  &  n_n3044 ) ;
 assign pv5_2_2_ = ( n_n4286  &  n_n3350 ) ;
 assign pv1_3_3_ = ( tin_pv1_3_3_  &  (~ n_n3441) ) | ( n_n3441  &  n_n4180 ) ;
 assign pv13_0_0_ = ( n_n3061  &  n_n3434 ) ;
 assign pv11_1_1_ = ( n_n4142  &  n_n4185 ) | ( tin_pv11_1_1_  &  (~ n_n4185) ) ;
 assign pv8_3_3_ = ( n_n3146  &  n_n3091 ) ;
 assign pv4_4_4_ = ( n_n3627  &  n_n4110 ) | ( tin_pv4_4_4_  &  (~ n_n4110) ) ;
 assign pready_0_0_ = ( tin_pready_0_0_  &  (~ n_n4108) ) | ( n_n4108  &  n_n3354 ) ;
 assign pv10_0_0_ = ( tin_pv10_0_0_  &  (~ n_n4282) ) | ( n_n4282  &  n_n4209 ) ;
 assign pv7_7_7_ = ( n_n3136  &  n_n4077 ) ;
 assign pv3_0_0_ = ( n_n3173  &  n_n3828 ) ;
 assign pv11_0_0_ = ( n_n3514  &  n_n3233 ) | ( tin_pv11_0_0_  &  (~ n_n3233) ) ;
 assign pv6_1_1_ = ( tin_pv6_1_1_  &  (~ n_n3144) ) | ( n_n3144  &  n_n3952 ) ;
 assign pv2_2_2_ = ( n_n3202  &  n_n4354 ) | ( tin_pv2_2_2_  &  (~ n_n4354) ) ;
 assign pv9_2_2_ = ( n_n3736  &  n_n3157 ) ;
 assign pv5_3_3_ = ( n_n3321  &  n_n4236 ) ;
 assign pv1_4_4_ = ( tin_pv1_4_4_  &  (~ n_n3863) ) | ( n_n3863  &  n_n3806 ) ;
 assign pv8_4_4_ = ( n_n3344  &  n_n3095 ) ;
 assign pv4_5_5_ = ( n_n3733  &  n_n3087 ) | ( tin_pv4_5_5_  &  (~ n_n3087) ) ;
 assign pv7_0_0_ = ( n_n3161  &  n_n3069 ) ;
 assign pv3_1_1_ = ( n_n3048  &  n_n3461 ) ;
 assign pv6_2_2_ = ( tin_pv6_2_2_  &  (~ n_n3307) ) | ( n_n3307  &  n_n3138 ) ;
 assign pv2_3_3_ = ( n_n3465  &  n_n3874 ) | ( tin_pv2_3_3_  &  (~ n_n3874) ) ;
 assign pv9_3_3_ = ( n_n3906  &  n_n3749 ) ;
 assign pv5_4_4_ = ( n_n3793  &  n_n4213 ) ;
 assign pv1_5_5_ = ( n_n3313  &  n_n3101 ) | ( tin_pv1_5_5_  &  (~ n_n3101) ) ;
 assign pv8_5_5_ = ( n_n3116  &  n_n3331 ) ;
 assign pv4_6_6_ = ( tin_pv4_6_6_  &  (~ n_n3774) ) | ( n_n3774  &  n_n3413 ) ;
 assign pv7_1_1_ = ( n_n3415  &  n_n3971 ) ;
 assign pv3_2_2_ = ( n_n3190  &  n_n3739 ) ;
 assign pv6_3_3_ = ( tin_pv6_3_3_  &  (~ n_n3204) ) | ( n_n3204  &  n_n3486 ) ;
 assign pv2_4_4_ = ( n_n3133  &  n_n3643 ) | ( tin_pv2_4_4_  &  (~ n_n3643) ) ;
 assign pv9_4_4_ = ( n_n3687  &  n_n3650 ) ;
 assign pv5_5_5_ = ( n_n3266  &  n_n3408 ) ;
 assign pv1_6_6_ = ( n_n3118  &  n_n4018 ) | ( tin_pv1_6_6_  &  (~ n_n4018) ) ;
 assign pv8_6_6_ = ( n_n3180  &  n_n3223 ) ;
 assign pv4_7_7_ = ( tin_pv4_7_7_  &  (~ n_n4114) ) | ( n_n4114  &  n_n4166 ) ;
 assign pv7_2_2_ = ( n_n3497  &  n_n4105 ) ;
 assign pv3_3_3_ = ( n_n3274  &  n_n4342 ) ;
 assign pv6_4_4_ = ( tin_pv6_4_4_  &  (~ n_n3093) ) | ( n_n3093  &  n_n4065 ) ;
 assign pv2_5_5_ = ( n_n3780  &  n_n4059 ) | ( tin_pv2_5_5_  &  (~ n_n4059) ) ;
 assign pv14_7_7_ = ( n_n3449  &  n_n4241 ) ;
 assign pv9_5_5_ = ( n_n3985  &  n_n4290 ) ;
 assign pv5_6_6_ = ( n_n3567  &  n_n3237 ) ;
 assign pv1_7_7_ = ( tin_pv1_7_7_  &  (~ n_n3544) ) | ( n_n3544  &  n_n4199 ) ;
 assign pv15_7_7_ = ( n_n3079  &  n_n3648 ) ;
 assign pv8_7_7_ = ( n_n3525  &  n_n3529 ) ;
 assign pv4_0_0_ = ( n_n3517  &  n_n3826 ) | ( tin_pv4_0_0_  &  (~ n_n3826) ) ;
 assign pv14_6_6_ = ( n_n3713  &  n_n3262 ) ;
 assign pv12_7_7_ = ( n_n3764  &  n_n3720 ) ;
 assign pv7_3_3_ = ( n_n3411  &  n_n4303 ) ;
 assign pv3_4_4_ = ( n_n3729  &  n_n4162 ) ;
 assign pv15_6_6_ = ( n_n4375  &  n_n3020 ) ;
 assign pv13_7_7_ = ( n_n3372  &  n_n3394 ) ;
 assign pv6_5_5_ = ( n_n4189  &  n_n3348 ) | ( tin_pv6_5_5_  &  (~ n_n3348) ) ;
 assign pv2_6_6_ = ( tin_pv2_6_6_  &  (~ n_n3120) ) | ( n_n3120  &  n_n3385 ) ;
 assign pv14_5_5_ = ( n_n3008  &  n_n3663 ) ;
 assign pv12_6_6_ = ( n_n3782  &  n_n3896 ) ;
 assign pv10_7_7_ = ( n_n3225  &  n_n3521 ) | ( tin_pv10_7_7_  &  (~ n_n3521) ) ;
 assign pv9_6_6_ = ( n_n4243  &  n_n3239 ) ;
 assign pv5_7_7_ = ( n_n3111  &  n_n4005 ) ;
 assign pv1_0_0_ = ( tin_pv1_0_0_  &  (~ n_n3551) ) | ( n_n3551  &  n_n4192 ) ;
 assign pv15_5_5_ = ( n_n3277  &  n_n3674 ) ;
 assign pv13_6_6_ = ( n_n3155  &  n_n3797 ) ;
 assign pv11_7_7_ = ( n_n3376  &  n_n3360 ) | ( tin_pv11_7_7_  &  (~ n_n3360) ) ;
 assign pv8_0_0_ = ( n_n3014  &  n_n4320 ) ;
 assign pv4_1_1_ = ( tin_pv4_1_1_  &  (~ n_n4089) ) | ( n_n4089  &  n_n3722 ) ;
 assign pv14_4_4_ = ( n_n3326  &  n_n3089 ) ;
 assign pv12_5_5_ = ( n_n3619  &  n_n3337 ) ;
 assign pv10_6_6_ = ( tin_pv10_6_6_  &  (~ n_n3570) ) | ( n_n3570  &  n_n3342 ) ;
 assign pv7_4_4_ = ( n_n3073  &  n_n3053 ) ;
 assign pv3_5_5_ = ( n_n3436  &  n_n3142 ) ;
 assign pv15_4_4_ = ( n_n3305  &  n_n3667 ) ;
 assign pv13_5_5_ = ( n_n4139  &  n_n3777 ) ;
 assign pv11_6_6_ = ( n_n4279  &  n_n3504 ) | ( tin_pv11_6_6_  &  (~ n_n3504) ) ;
 assign pv6_6_6_ = ( n_n3429  &  n_n3836 ) | ( tin_pv6_6_6_  &  (~ n_n3836) ) ;
 assign pv2_7_7_ = ( tin_pv2_7_7_  &  (~ n_n4131) ) | ( n_n4131  &  n_n3126 ) ;
 assign pv14_3_3_ = ( n_n3396  &  n_n3316 ) ;
 assign pv12_4_4_ = ( n_n3231  &  n_n3175 ) ;
 assign pv10_5_5_ = ( tin_pv10_5_5_  &  (~ n_n3381) ) | ( n_n3381  &  n_n4247 ) ;
 assign pv9_7_7_ = ( n_n3319  &  n_n3040 ) ;
 assign pv5_0_0_ = ( n_n3195  &  n_n3572 ) ;
 assign pv1_1_1_ = ( tin_pv1_1_1_  &  (~ n_n3215) ) | ( n_n3215  &  n_n3183 ) ;
 assign pv15_3_3_ = ( n_n4172  &  n_n3051 ) ;
 assign pv13_4_4_ = ( n_n3075  &  n_n3758 ) ;
 assign pv11_5_5_ = ( tin_pv11_5_5_  &  (~ n_n3081) ) | ( n_n3081  &  n_n3207 ) ;
 assign pv8_1_1_ = ( n_n3938  &  n_n3883 ) ;
 assign pv4_2_2_ = ( tin_pv4_2_2_  &  (~ n_n4347) ) | ( n_n4347  &  n_n4372 ) ;
 assign n_n4140 = ( wire2275 ) | ( n_n3724  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3935 = ( wire2270 ) | ( pv11_1_1_  &  wire988 ) ;
 assign n_n3444 = ( wire2261 ) | ( wire2262 ) | ( wire2263 ) ;
 assign n_n3007 = ( wire2259 ) | ( n_n3035  &  n_n4157  &  wire894 ) ;
 assign n_n3725 = ( wire2240 ) | ( wire2241 ) | ( wire2242 ) ;
 assign n_n3399 = ( (~ preset)  &  wire1016 ) ;
 assign n_n3143 = ( (~ preset)  &  n_n3144 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3781 = ( (~ preset)  &  n_n3782 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3066 = ( (~ preset)  &  n_n3067 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3507 = ( wire2226 ) | ( pv10_3_3_  &  wire992 ) ;
 assign n_n3224 = ( wire2224 ) | ( n_n4360  &  wire894 ) ;
 assign n_n3179 = ( (~ preset)  &  n_n3180 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3273 = ( (~ preset)  &  n_n3274 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3166 = ( n_n3475  &  wire934 ) | ( n_n3475  &  wire916  &  wire1019 ) | ( (~ n_n3475)  &  wire916  &  (~ wire1019) ) ;
 assign n_n3686 = ( wire2202 ) | ( n_n3458  &  wire894 ) ;
 assign n_n3380 = ( (~ preset)  &  n_n3381 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3096 = ( wire2198 ) | ( n_n3688  &  n_n3624  &  wire894 ) ;
 assign n_n4106 = ( (~ preset)  &  wire1020 ) ;
 assign n_n3496 = ( wire2195 ) | ( n_n3901  &  wire894  &  n_n4367 ) ;
 assign n_n3791 = ( wire2192 ) | ( n_n3916  &  wire894  &  wire1096 ) | ( (~ n_n3916)  &  wire894  &  (~ wire1096) ) ;
 assign n_n3518 = ( wire2166 ) | ( n_n4015  &  wire1004 ) ;
 assign n_n4348 = ( wire2162 ) | ( pv6_0_0_  &  wire990 ) ;
 assign n_n3028 = ( (~ preset)  &  n_n3029 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3618 = ( (~ preset)  &  n_n3619 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3263 = ( (~ preset)  &  n_n3264 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3778 = ( wire2153 ) | ( n_n4288  &  wire894 ) | ( wire894  &  wire6259 ) ;
 assign n_n3227 = ( (~ preset)  &  (~ ngfdn_3)  &  wire1021 ) ;
 assign n_n4113 = ( (~ preset)  &  n_n4114 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3145 = ( (~ preset)  &  n_n3146 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3510 = ( wire2141 ) | ( pv1_5_5_  &  wire994 ) ;
 assign n_n3151 = ( (~ preset)  &  n_n3152 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n129 = ( preset ) | ( n_n3833  &  wire1022 ) | ( (~ n_n3563)  &  (~ wire1022) ) ;
 assign n_n4280 = ( (~ preset)  &  n_n4282 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3304 = ( (~ preset)  &  n_n3305 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3309 = ( wire2126 ) | ( wire1002  &  n_n3363  &  wire1128 ) | ( wire1002  &  (~ n_n3363)  &  (~ wire1128) ) ;
 assign n_n3490 = ( wire2122 ) | ( pv4_5_5_  &  wire997 ) ;
 assign n_n3377 = ( (~ preset)  &  (~ wire1137)  &  wire6290 ) | ( (~ preset)  &  (~ wire1136)  &  wire6290 ) ;
 assign n_n3203 = ( (~ preset)  &  n_n3204 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3023 = ( (~ preset)  &  n_n3024 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4137 = ( (~ preset)  &  n_n4139 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3084 = ( (~ preset)  &  ndn3_15  &  (~ ngfdn_3) ) ;
 assign n_n3131 = ( wire2051 ) | ( n_n3458  &  wire894 ) | ( wire894  &  wire6291 ) ;
 assign n_n4073 = ( wire2029 ) | ( n_n3810  &  n_n4345  &  wire1122 ) | ( n_n3810  &  (~ n_n4345)  &  (~ wire1122) ) ;
 assign n_n3269 = ( wire2027 ) | ( n_n3743  &  wire894 ) ;
 assign n_n3181 = ( wire2023 ) | ( pv1_2_2_  &  wire994 ) ;
 assign n_n3455 = ( (~ preset)  &  n_n3456 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3520 = ( (~ preset)  &  n_n3521 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3080 = ( (~ preset)  &  n_n3081 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3296 = ( wire2007 ) | ( wire1006  &  wire2009 ) | ( wire1006  &  wire6300 ) ;
 assign n_n3668 = ( wire2005 ) | ( n_n3475  &  wire894  &  n_n4367 ) ;
 assign n_n4210 = ( wire2000 ) | ( pv11_2_2_  &  wire988 ) ;
 assign n_n3076 = ( n_n4045  &  n_n4367  &  wire6302 ) | ( n_n4045  &  (~ wire6299)  &  wire6302 ) ;
 assign n_n3148 = ( wire1998 ) | ( n_n4015  &  wire1002 ) ;
 assign n_n3226 = ( wire1996 ) | ( wire1004  &  n_n4345  &  wire1122 ) | ( wire1004  &  (~ n_n4345)  &  (~ wire1122) ) ;
 assign n_n3194 = ( (~ preset)  &  n_n3195 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3523 = ( wire1992 ) | ( n_n3242  &  wire894 ) ;
 assign n_n3727 = ( wire1990 ) | ( n_n3916  &  wire894 ) ;
 assign n_n3875 = ( wire1986 ) | ( pv10_4_4_  &  wire992 ) ;
 assign n_n3614 = ( (~ preset)  &  ndn3_4  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_5  &  (~ ngfdn_3) ) ;
 assign n_n3547 = ( wire1984 ) | ( n_n3946  &  wire894 ) ;
 assign n_n3488 = ( (~ preset)  &  n_n3489 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3762 = ( wire1980 ) | ( n_n3242  &  n_n3170  &  wire894 ) ;
 assign n_n3256 = ( wire1976 ) | ( pv2_3_3_  &  wire999 ) ;
 assign n_n124 = ( preset ) | ( nak3_17 ) | ( wire1971 ) ;
 assign n_n3515 = ( wire1969 ) | ( n_n4159  &  wire894 ) ;
 assign n_n3016 = ( wire1965 ) | ( pv4_1_1_  &  wire997 ) ;
 assign n_n3168 = ( wire1963 ) | ( wire1004  &  n_n3363  &  wire1128 ) | ( wire1004  &  (~ n_n3363)  &  (~ wire1128) ) ;
 assign n_n3011 = ( wire1961 ) | ( n_n3936  &  n_n3099  &  wire894 ) ;
 assign n_n3373 = ( wire1957 ) | ( pv6_5_5_  &  wire990 ) ;
 assign n_n3371 = ( (~ preset)  &  n_n3372 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3343 = ( wire1953 ) | ( n_n4074  &  wire894 ) ;
 assign n_n3018 = ( wire1949 ) | ( n_n3810  &  (~ n_n3975)  &  n_n3974 ) | ( n_n3810  &  n_n3975  &  (~ n_n3974) ) ;
 assign n_n3077 = ( wire1946 ) | ( n_n4233  &  wire894 ) | ( wire894  &  wire6303 ) ;
 assign n_n3312 = ( wire1944 ) | ( n_n3035  &  n_n4157  &  wire894 ) ;
 assign n_n3410 = ( (~ preset)  &  n_n3411 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3230 = ( wire1940 ) | ( n_n4074  &  n_n3578  &  wire894 ) ;
 assign n_n3395 = ( (~ preset)  &  n_n3396 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3431 = ( (~ preset)  &  n_n3432 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3605 = ( (~ preset)  &  n_n3606 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3732 = ( wire1932 ) | ( n_n4224  &  wire894 ) ;
 assign n_n3063 = ( wire1928 ) | ( pv11_6_6_  &  wire988 ) ;
 assign n_n3913 = ( wire1925 ) | ( wire1926 ) | ( wire1927 ) ;
 assign n_n3119 = ( (~ preset)  &  n_n3120 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3220 = ( wire1921 ) | ( n_n4222  &  wire894 ) ;
 assign n_n3172 = ( wire1919 ) | ( n_n3976  &  wire894 ) ;
 assign n_n3070 = ( (~ preset)  &  n_n3851  &  wire936 ) | ( (~ preset)  &  n_n3852  &  (~ wire936) ) ;
 assign n_n3112 = ( wire1914 ) | ( n_n3495  &  wire894 ) | ( wire894  &  wire6310 ) ;
 assign n_n3241 = ( wire1884 ) | ( wire1885 ) ;
 assign n_n3117 = ( wire1882 ) | ( n_n3556  &  n_n4122  &  wire894 ) ;
 assign n_n3375 = ( wire1881 ) | ( n_n3483  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n4088 = ( (~ preset)  &  n_n4089 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3043 = ( wire1876 ) | ( n_n4392  &  wire894 ) ;
 assign n_n3625 = ( wire1874 ) | ( n_n4330  &  wire894 ) ;
 assign n_n3027 = ( wire1870 ) | ( pv11_5_5_  &  wire988 ) ;
 assign n_n3110 = ( wire1868 ) | ( n_n3841  &  wire894  &  wire1078 ) | ( (~ n_n3841)  &  wire894  &  (~ wire1078) ) ;
 assign n_n3320 = ( (~ preset)  &  n_n3321 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3442 = ( (~ preset)  &  n_n3443 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3214 = ( (~ preset)  &  n_n3215 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3751 = ( (~ preset)  &  ndn3_10  &  (~ ngfdn_3) ) | ( (~ preset)  &  nen3_10  &  (~ ngfdn_3) ) ;
 assign n_n4170 = ( wire1859 ) | ( n_n4351  &  wire894 ) | ( wire894  &  wire6322 ) ;
 assign n_n3982 = ( (~ preset)  &  (~ pdn)  &  wire1028 ) ;
 assign n_n3589 = ( (~ preset)  &  n_n3590 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4109 = ( (~ preset)  &  n_n4110 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3941 = ( nlc3_3  &  (~ wire944) ) | ( (~ wire944)  &  nrq3_2  &  wire6324 ) ;
 assign n_n3575 = ( wire1853 ) | ( n_n4211  &  n_n3657  &  wire894 ) ;
 assign n_n4128 = ( (~ preset)  &  n_n4129 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4186 = ( wire1849 ) | ( n_n4071  &  wire894 ) ;
 assign n_n4283 = ( wire1847 ) | ( wire894  &  n_n4116 ) ;
 assign n_n3022 = ( wire1843 ) | ( pv4_2_2_  &  wire997 ) ;
 assign n_n3437 = ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3566 = ( (~ preset)  &  n_n3567 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3032 = ( wire1837 ) | ( pv6_6_6_  &  wire990 ) ;
 assign n_n3074 = ( (~ preset)  &  n_n3075 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3353 = ( wire1833 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3464 = ( wire1830 ) | ( n_n4351  &  wire894 ) | ( wire894  &  wire6322 ) ;
 assign n_n4321 = ( (~ preset)  &  ndn3_5  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_6  &  (~ ngfdn_3) ) ;
 assign n_n3616 = ( (~ preset)  &  n_n3617 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4161 = ( (~ preset)  &  n_n4162 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3206 = ( wire1825 ) | ( n_n4012  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n4119 = ( (~ preset)  &  n_n4120 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3064 = ( (~ preset)  &  n_n3065 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4004 = ( (~ preset)  &  n_n4005 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3265 = ( (~ preset)  &  n_n3266 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3216 = ( wire1812 ) | ( pv6_7_7_  &  wire990 ) ;
 assign n_n3599 = ( (~ preset)  &  n_n3600 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3414 = ( (~ preset)  &  n_n3415 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4242 = ( wire1806 ) | ( n_n4095  &  wire894 ) ;
 assign n_n3871 = ( (~ preset)  &  n_n3872 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3647 = ( (~ preset)  &  n_n3648 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3357 = ( wire1800 ) | ( n_n4211  &  n_n3657  &  wire894 ) ;
 assign n_n3349 = ( (~ preset)  &  n_n3350 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3675 = ( (~ preset)  &  ndn3_6  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_7  &  (~ ngfdn_3) ) ;
 assign n_n3115 = ( (~ preset)  &  n_n3116 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3582 = ( wire1795 ) | ( n_n3766  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3904 = ( wire1792 ) | ( n_n4351  &  wire894 ) ;
 assign n_n4130 = ( (~ preset)  &  n_n4131 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3314 = ( wire1788 ) | ( n_n3085  &  n_n3250  &  wire894 ) ;
 assign n_n3060 = ( wire1786 ) | ( n_n3976  &  wire894 ) ;
 assign n_n3047 = ( wire1784 ) | ( n_n4222  &  wire894 ) ;
 assign n_n3837 = ( wire1780 ) | ( pv1_4_4_  &  wire994 ) ;
 assign n_n3508 = ( wire1776 ) | ( pv1_6_6_  &  wire994 ) ;
 assign n_n3127 = ( wire1774 ) | ( n_n3608  &  wire894 ) ;
 assign n_n3235 = ( wire1771 ) | ( wire1772 ) | ( wire1773 ) ;
 assign n_n4212 = ( (~ preset)  &  n_n4213 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3759 = ( wire1767 ) | ( n_n3688  &  n_n3624  &  wire894 ) ;
 assign n_n4218 = ( (~ preset)  &  ndn3_7  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_8  &  (~ ngfdn_3) ) ;
 assign n_n3251 = ( (~ preset)  &  n_n3252 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3382 = ( n_n4366  &  wire934 ) | ( n_n4366  &  wire916  &  wire1034 ) | ( (~ n_n4366)  &  wire916  &  (~ wire1034) ) ;
 assign n_n3327 = ( wire1755 ) | ( pv2_1_1_  &  wire999 ) ;
 assign n_n3987 = ( wire1752 ) | ( wire1753 ) | ( wire1754 ) ;
 assign n_n3347 = ( (~ preset)  &  n_n3348 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3543 = ( (~ preset)  &  n_n3544 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3100 = ( (~ preset)  &  n_n3101 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4276 = ( wire1745 ) | ( n_n4334  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3895 = ( wire1742 ) | ( n_n3556  &  n_n4122  &  wire894 ) ;
 assign n_n3735 = ( wire1740 ) | ( n_n3495  &  wire894 ) ;
 assign n_n3049 = ( wire1736 ) | ( pv4_6_6_  &  wire997 ) ;
 assign n_n3649 = ( (~ preset)  &  n_n3650 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3306 = ( (~ preset)  &  n_n3307 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4293 = ( wire1728 ) | ( pv1_3_3_  &  wire994 ) ;
 assign n_n3907 = ( (~ n_n4334)  &  wire1014 ) | ( n_n4334  &  wire982 ) | ( n_n4334  &  wire1724 ) ;
 assign n_n3579 = ( wire1716 ) | ( wire1006  &  wire1719 ) | ( wire1006  &  wire6332 ) ;
 assign n_n4163 = ( (~ preset)  &  n_n4164 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3154 = ( wire1711 ) | ( n_n4145  &  wire894 ) ;
 assign n_n3748 = ( (~ preset)  &  n_n3749 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3271 = ( wire1707 ) | ( wire1708 ) ;
 assign n_n4346 = ( (~ preset)  &  n_n4347 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3825 = ( (~ preset)  &  n_n3826 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3359 = ( (~ preset)  &  n_n3360 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3147 = ( wire1699 ) | ( wire1002  &  n_n4345  &  wire1122 ) | ( wire1002  &  (~ n_n4345)  &  (~ wire1122) ) ;
 assign n_n3092 = ( (~ preset)  &  n_n3093 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3156 = ( (~ preset)  &  n_n3157 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3505 = ( wire1693 ) | ( n_n4349  &  wire894 ) ;
 assign n_n3160 = ( (~ preset)  &  n_n3161 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3318 = ( wire1689 ) | ( n_n4233  &  wire894 ) ;
 assign n_n3428 = ( wire1687 ) | ( n_n3892  &  wire894 ) ;
 assign n_n3969 = ( wire1686 ) | ( n_n4125  &  wire894  &  n_n4367 ) ;
 assign n_n3447 = ( wire1683 ) | ( n_n3242  &  n_n3170  &  wire894 ) ;
 assign n_n4081 = ( wire1679 ) | ( pv4_7_7_  &  wire997 ) ;
 assign n_n3302 = ( wire1673 ) | ( wire1002  &  n_n4158 ) ;
 assign n_n3182 = ( wire1671 ) | ( n_n3936  &  n_n3099  &  wire894 ) ;
 assign n_n3129 = ( (~ preset)  &  n_n3130 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3430 = ( (~ preset)  &  nsr4_2  &  (~ wire973) ) ;
 assign n_n4046 = ( wire1659 ) | ( (~ preset)  &  n_n4047  &  (~ n_n4126) ) ;
 assign n_n3123 = ( wire1655 ) | ( pv2_2_2_  &  wire999 ) ;
 assign n_n3238 = ( (~ preset)  &  n_n3239 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3972 = ( wire1647 ) | ( wire1648 ) ;
 assign n_n3889 = ( (~ preset)  &  n_n3890 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4001 = ( wire1642 ) | ( n_n3608  &  wire894 ) | ( wire894  &  wire6272 ) ;
 assign n_n3090 = ( wire1640 ) | ( n_n3085  &  wire894 ) ;
 assign n_n3983 = ( wire1638 ) | ( n_n4288  &  wire894 ) ;
 assign n_n3325 = ( (~ preset)  &  n_n3326 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3540 = ( wire1630 ) | ( wire1006  &  wire1633 ) | ( wire1006  &  wire6337 ) ;
 assign n_n125 = ( preset ) | ( pdn ) | ( nsr4_2  &  wire973 ) ;
 assign n_n3693 = ( wire1621 ) | ( wire1006  &  wire1623 ) | ( wire1006  &  wire6338 ) ;
 assign n_n4373 = ( (~ preset)  &  n_n4375 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3866 = ( (~ preset)  &  (~ nak3_17)  &  wire1041 ) ;
 assign n_n4289 = ( (~ preset)  &  n_n4290 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3459 = ( wire1614 ) | ( wire1004  &  n_n4158 ) ;
 assign n_n4121 = ( wire1612 ) | ( wire1613 ) ;
 assign n_n3773 = ( (~ preset)  &  n_n3774 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3013 = ( (~ preset)  &  n_n3014 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4239 = ( (~ preset)  &  n_n4241 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3950 = ( wire1604 ) | ( n_n4201  &  wire894 ) ;
 assign n_n3236 = ( wire1602 ) | ( n_n4145  &  wire894  &  wire1075 ) | ( (~ n_n4145)  &  wire894  &  (~ wire1075) ) ;
 assign n_n3530 = ( wire1598 ) | ( pv6_2_2_  &  wire990 ) ;
 assign n_n3033 = ( wire1594 ) | ( pv6_4_4_  &  wire990 ) ;
 assign n_n3550 = ( (~ preset)  &  n_n3551 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3378 = ( (~ preset)  &  n_n3379 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3009 = ( wire1580 ) | ( n_n4275  &  wire1042 ) ;
 assign n_n3569 = ( (~ preset)  &  n_n3570 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3853 = ( wire1574 ) | ( pv2_5_5_  &  wire999 ) ;
 assign n_n131 = ( wire1565 ) | ( wire6350 ) ;
 assign n_n3450 = ( wire1561 ) | ( pv2_7_7_  &  wire999 ) ;
 assign n_n4036 = ( (~ preset)  &  n_n4037 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3406 = ( wire1557 ) | ( n_n3898  &  wire894  &  wire1076 ) | ( (~ n_n3898)  &  wire894  &  (~ wire1076) ) ;
 assign n_n4228 = ( wire1551 ) | ( wire1552 ) ;
 assign n_n3701 = ( wire1547 ) | ( pv6_1_1_  &  wire990 ) ;
 assign n_n3338 = ( (~ preset)  &  n_n3339 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4361 = ( wire1541 ) | ( pv10_5_5_  &  wire992 ) ;
 assign n_n3466 = ( wire1538 ) | ( n_n4334  &  (~ n_n3483)  &  wire1014 ) ;
 assign n_n3355 = ( (~ preset)  &  (~ n_n4099)  &  wire1119  &  wire6349 ) | ( (~ preset)  &  n_n4099  &  (~ wire1119)  &  wire6349 ) ;
 assign n_n4184 = ( (~ preset)  &  n_n4185 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3068 = ( wire1534 ) | ( n_n3934  &  wire894  &  n_n4367 ) ;
 assign n_n3642 = ( (~ preset)  &  n_n3643 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3402 = ( wire1529 ) | ( n_n4229  &  wire894 ) ;
 assign n_n3056 = ( wire1527 ) | ( n_n4145  &  wire894 ) ;
 assign n_n3019 = ( wire1524 ) | ( n_n4095  &  wire894 ) | ( wire894  &  wire6321 ) ;
 assign n_n3827 = ( (~ preset)  &  n_n3828 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3629 = ( wire1520 ) | ( n_n3085  &  n_n3250  &  wire894 ) ;
 assign n_n3137 = ( wire1518 ) | ( n_n3968  &  wire894 ) ;
 assign n_n126 = ( preset ) | ( pdn ) | ( (~ ngfdn_3)  &  (~ nrq1_3) ) ;
 assign n_n4063 = ( wire1514 ) | ( n_n3922  &  wire894 ) ;
 assign n_n3677 = ( wire1513 ) | ( n_n4366  &  wire894  &  n_n4367 ) ;
 assign n_n3285 = ( wire1510 ) | ( wire894  &  n_n3741 ) ;
 assign n_n3308 = ( wire1508 ) | ( wire1509 ) ;
 assign n_n4058 = ( (~ preset)  &  n_n4059 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3435 = ( wire1504 ) | ( n_n3898  &  wire894 ) ;
 assign n_n3635 = ( (~ preset)  &  nen3_10  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_9  &  (~ ngfdn_3) ) ;
 assign n_n3460 = ( (~ preset)  &  n_n3461 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4011 = ( wire1500 ) | ( n_n4012  &  wire982 ) ;
 assign n_n3050 = ( (~ preset)  &  n_n3051 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3072 = ( wire1497 ) | ( n_n4047  &  wire894  &  n_n4367 ) ;
 assign n_n3775 = ( wire1494 ) | ( n_n3898  &  wire894 ) ;
 assign n_n3199 = ( wire1492  &  wire6354 ) | ( n_n3832  &  wire6255  &  wire6354 ) ;
 assign n_n3025 = ( wire1488 ) | ( pv10_2_2_  &  wire992 ) ;
 assign n_n3058 = ( wire1486 ) | ( wire1487 ) ;
 assign n_n3258 = ( wire1482 ) | ( pv1_7_7_  &  wire994 ) ;
 assign n_n3503 = ( (~ preset)  &  n_n3504 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n130 = ( wire6357 ) | ( n_n4045  &  wire1477 ) | ( n_n4045  &  wire6356 ) ;
 assign n_n121 = ( (~ wire1006)  &  (~ wire1470) ) | ( (~ wire1470)  &  (~ wire1472)  &  (~ wire6358) ) ;
 assign n_n3134 = ( wire1468 ) | ( n_n4324  &  wire894  &  n_n4367 ) ;
 assign n_n4370 = ( wire1465 ) | ( n_n4383  &  wire894 ) ;
 assign n_n4234 = ( wire1463 ) | ( n_n4229  &  wire894  &  wire1079 ) | ( (~ n_n4229)  &  wire894  &  (~ wire1079) ) ;
 assign n_n3039 = ( (~ preset)  &  n_n3040 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3873 = ( (~ preset)  &  n_n3874 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3998 = ( (~ preset)  &  n_n3999 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3222 = ( wire1455 ) | ( n_n4122  &  wire894 ) ;
 assign n_n3036 = ( (~ preset)  &  (~ pdn)  &  ndn1_34 ) ;
 assign n_n3062 = ( wire1451 ) | ( pv10_1_1_  &  wire992 ) ;
 assign n_n3017 = ( wire1449 ) | ( n_n3810  &  n_n4015 ) ;
 assign n_n3212 = ( wire1447 ) | ( n_n4258  &  wire894 ) ;
 assign n_n3094 = ( (~ preset)  &  n_n3095 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3662 = ( (~ preset)  &  n_n3663 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3217 = ( n_n3724  &  wire947 ) | ( (~ n_n3724)  &  n_n3814  &  wire896 ) ;
 assign n_n3037 = ( (~ preset)  &  n_n3038 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3368 = ( wire1437 ) | ( n_n4337  &  wire894 ) ;
 assign n_n3030 = ( wire1433 ) | ( pv11_0_0_  &  wire988 ) ;
 assign n_n3494 = ( wire1429 ) | ( pv11_4_4_  &  wire988 ) ;
 assign n_n3711 = ( wire1427 ) | ( n_n3556  &  n_n4122  &  wire894 ) ;
 assign n_n3088 = ( wire1425 ) | ( n_n4074  &  n_n3578  &  wire894 ) ;
 assign n_n3210 = ( (~ preset)  &  n_n3211 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3366 = ( (~ preset)  &  n_n3367 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3433 = ( (~ preset)  &  n_n3434 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3125 = ( wire1416 ) | ( n_n4233  &  wire894 ) | ( wire894  &  wire6303 ) ;
 assign n_n4190 = ( wire1414 ) | ( n_n3688  &  n_n3624  &  wire894 ) ;
 assign n_n4134 = ( wire1412 ) | ( n_n3876  &  wire894 ) ;
 assign n_n3052 = ( (~ preset)  &  n_n3053 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3937 = ( (~ preset)  &  n_n3938 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3632 = ( wire1402 ) | ( (~ preset)  &  n_n3769  &  (~ n_n4126) ) ;
 assign n_n4387 = ( wire1400 ) | ( n_n3936  &  n_n3099  &  wire894 ) ;
 assign n_n127 = ( wire944 ) | ( (~ nen3_10)  &  nsr3_17 ) | ( nsr3_17  &  (~ nak3_17) ) ;
 assign n_n3902 = ( (~ preset)  &  n_n3903 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3684 = ( n_n3658  &  wire6361 ) | ( n_n4367  &  wire6268  &  wire6361 ) ;
 assign n_n3046 = ( (~ preset)  &  nrq3_11  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ nsr3_14)  &  (~ ngfdn_3) ) ;
 assign n_n3817 = ( wire1391 ) | ( wire1392 ) | ( wire1393 ) ;
 assign n_n3374 = ( wire1387 ) | ( pv6_3_3_  &  wire990 ) ;
 assign n_n3462 = ( wire1385 ) | ( n_n4316  &  wire894 ) ;
 assign n_n3174 = ( (~ preset)  &  n_n3175 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3054 = ( wire1381 ) | ( n_n3657  &  wire894 ) ;
 assign n_n3200 = ( wire1378 ) | ( n_n3495  &  wire894 ) | ( wire894  &  wire6310 ) ;
 assign n_n3383 = ( wire1375 ) | ( n_n4095  &  wire894 ) | ( wire894  &  wire6321 ) ;
 assign n_n4076 = ( (~ preset)  &  n_n4077 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3141 = ( (~ preset)  &  n_n3142 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3289 = ( wire1365 ) | ( (~ preset)  &  n_n3901  &  (~ n_n4126) ) ;
 assign n_n3552 = ( wire1362 ) | ( (~ n_n3934)  &  n_n3976  &  wire916 ) ;
 assign n_n3821 = ( wire1360 ) | ( n_n4227  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3721 = ( wire1357 ) | ( n_n4160  &  wire894 ) ;
 assign n_n4307 = ( wire1355 ) | ( n_n4182  &  wire894 ) ;
 assign n_n3229 = ( wire1351 ) | ( pv4_0_0_  &  wire997 ) ;
 assign n_n3021 = ( wire1347 ) | ( pv4_4_4_  &  wire997 ) ;
 assign n_n3835 = ( (~ preset)  &  n_n3836 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3469 = ( (~ preset)  &  n_n3470 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3329 = ( wire1341 ) | ( n_n4157  &  wire894 ) ;
 assign n_n3881 = ( wire1339 ) | ( n_n3099  &  wire894 ) ;
 assign n_n3031 = ( wire1335 ) | ( pv10_6_6_  &  wire992 ) ;
 assign n_n4156 = ( wire1333 ) | ( n_n3810  &  n_n4158 ) ;
 assign n_n4086 = ( (~ preset)  &  ndn3_8  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_9  &  (~ ngfdn_3) ) ;
 assign n_n3045 = ( wire1329 ) | ( pv1_1_1_  &  wire994 ) ;
 assign n_n3189 = ( (~ preset)  &  n_n3190 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4028 = ( wire1323 ) | ( wire1006  &  wire1325 ) | ( wire1006  &  wire6366 ) ;
 assign n_n3041 = ( (~ preset)  &  n_n3042 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n133 = ( preset ) | ( pdn ) | ( wire1318 ) ;
 assign n_n122 = ( preset ) | ( wire1315 ) | ( wire1316 ) ;
 assign n_n3187 = ( (~ preset)  &  n_n3188 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4300 = ( wire1312 ) | ( n_n3769  &  wire894  &  n_n4367 ) ;
 assign n_n3249 = ( wire1307 ) | ( pv11_3_3_  &  wire988 ) ;
 assign n_n3169 = ( wire1303 ) | ( pv11_7_7_  &  wire988 ) ;
 assign n_n3757 = ( wire1301 ) | ( n_n3916  &  wire894 ) ;
 assign n_n3908 = ( wire1298 ) | ( n_n3608  &  wire894 ) | ( wire894  &  wire6272 ) ;
 assign n_n3106 = ( wire1295 ) | ( n_n4392  &  wire894 ) | ( wire894  &  wire6306 ) ;
 assign n_n3149 = ( (~ preset)  &  n_n3150 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4317 = ( wire1291 ) | ( n_n3688  &  wire894 ) ;
 assign n_n4359 = ( wire1287 ) | ( pv10_7_7_  &  wire992 ) ;
 assign n_n4245 = ( wire1285 ) | ( n_n4362  &  wire894 ) ;
 assign n_n4196 = ( wire1283 ) | ( n_n3242  &  n_n3170  &  wire894 ) ;
 assign n_n3964 = ( wire1282 ) | ( n_n4275  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3184 = ( wire1280 ) | ( wire896  &  wire6370 ) ;
 assign n_n3010 = ( wire1275 ) | ( pv2_4_4_  &  wire999 ) ;
 assign n_n3122 = ( wire1271 ) | ( pv2_6_6_  &  wire999 ) ;
 assign n_n3512 = ( wire1270 ) | ( n_n3814  &  (~ n_n3830)  &  wire6252 ) ;
 assign n_n3571 = ( wire1267 ) | ( (~ n_n4159)  &  n_n3976  &  wire894 ) | ( n_n4159  &  (~ n_n3976)  &  wire894 ) ;
 assign n_n4165 = ( wire1265 ) | ( n_n4270  &  wire894 ) ;
 assign n_n3519 = ( wire1263 ) | ( wire1004  &  (~ n_n3975)  &  n_n3974 ) | ( wire1004  &  n_n3975  &  (~ n_n3974) ) ;
 assign n_n3392 = ( wire1261 ) | ( n_n3841  &  wire894 ) ;
 assign n_n4094 = ( wire1259 ) | ( wire1260 ) ;
 assign n_n3862 = ( (~ preset)  &  n_n3863 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3719 = ( (~ preset)  &  n_n3720 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3810 = ( (~ preset)  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign n_n3755 = ( wire1251 ) | ( pv10_0_0_  &  wire992 ) ;
 assign n_n3665 = ( wire1248 ) | ( n_n3458  &  wire894 ) | ( wire894  &  wire6291 ) ;
 assign n_n3340 = ( wire1246 ) | ( n_n4299  &  wire894 ) ;
 assign n_n3528 = ( (~ preset)  &  n_n3529 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4207 = ( wire1242 ) | ( n_n3756  &  wire894 ) ;
 assign n_n3585 = ( n_n4324  &  wire934 ) | ( n_n4324  &  wire916  &  wire1062 ) | ( (~ n_n4324)  &  wire916  &  (~ wire1062) ) ;
 assign n_n3336 = ( wire1232 ) | ( n_n3035  &  n_n4157  &  wire894 ) ;
 assign n_n3026 = ( wire1230 ) | ( n_n4227  &  wire947 ) | ( n_n4227  &  wire1586 ) ;
 assign n_n4152 = ( (~ preset)  &  n_n4153 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n128 = ( wire1225 ) | ( wire6376 ) ;
 assign n_n3232 = ( (~ preset)  &  n_n3233 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4262 = ( (~ preset)  &  wire1064 ) ;
 assign n_n3412 = ( wire1218 ) | ( n_n4251  &  wire894 ) ;
 assign n_n3015 = ( wire1214 ) | ( pv4_3_3_  &  wire997 ) ;
 assign n_n3526 = ( wire1212 ) | ( wire1213 ) ;
 assign n_n3440 = ( (~ preset)  &  n_n3441 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3140 = ( (~ preset)  &  n_n4026  &  (~ nak3_17) ) | ( (~ preset)  &  (~ nak3_17)  &  wire1208 ) ;
 assign n_n4339 = ( wire1206 ) | ( n_n4229  &  wire894 ) ;
 assign n_n4100 = ( wire1204 ) | ( n_n3841  &  wire894 ) ;
 assign n_n3275 = ( wire1201 ) | ( n_n4288  &  wire894 ) | ( wire894  &  wire6259 ) ;
 assign n_n4178 = ( wire1199 ) | ( n_n3085  &  n_n3250  &  wire894 ) ;
 assign n_n3877 = ( wire1195 ) | ( pv1_0_0_  &  wire994 ) ;
 assign n_n3538 = ( wire1191 ) | ( pv2_0_0_  &  wire999 ) ;
 assign n_n3680 = ( wire1187 ) | ( wire1006  &  wire1189 ) | ( wire1006  &  wire6379 ) ;
 assign n_n3104 = ( wire1182 ) | ( wire1006  &  wire1184 ) | ( wire1006  &  wire6380 ) ;
 assign n_n3484 = ( wire1179 ) | ( n_n3533  &  wire894 ) ;
 assign n_n3473 = ( (~ preset)  &  n_n4057  &  wire1068 ) ;
 assign n_n3673 = ( (~ preset)  &  n_n3674 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3592 = ( wire1171 ) | ( wire1172 ) | ( n_n3959  &  wire1069 ) ;
 assign n_n3607 = ( wire1168 ) | ( wire1002  &  (~ n_n3975)  &  n_n3974 ) | ( wire1002  &  n_n3975  &  (~ n_n3974) ) ;
 assign n_n3292 = ( wire1165 ) | ( wire1166 ) | ( wire1167 ) ;
 assign n_n4017 = ( (~ preset)  &  n_n4018 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4352 = ( (~ preset)  &  n_n4354 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3796 = ( (~ preset)  &  n_n3797 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3737 = ( wire983 ) | ( n_n4316  &  wire894 ) ;
 assign n_n3644 = ( wire978 ) | ( n_n4392  &  wire894 ) | ( wire894  &  wire6306 ) ;
 assign n_n3059 = ( wire976 ) | ( n_n3810  &  n_n3363  &  wire1128 ) | ( n_n3810  &  (~ n_n3363)  &  (~ wire1128) ) ;
 assign n_n3535 = ( wire974 ) | ( n_n4211  &  n_n3657  &  wire894 ) ;
 assign n_n3804 = ( wire971 ) | ( n_n4074  &  n_n3578  &  wire894 ) ;
 assign n_n3086 = ( (~ preset)  &  n_n3087 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4104 = ( (~ preset)  &  n_n4105 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n3261 = ( (~ preset)  &  n_n3262 ) | ( (~ preset)  &  (~ pdn)  &  nrq1_3 ) ;
 assign n_n4124 = ( n_n4126  &  wire6385 ) | ( (~ preset)  &  n_n4125  &  (~ n_n4126) ) ;
 assign n_n3813 = ( wire946 ) | ( (~ n_n3814)  &  wire896 ) ;
 assign n_n132 = ( (~ wire6389) ) | ( (~ n_n3832)  &  (~ wire921) ) | ( (~ wire921)  &  (~ wire6386) ) ;
 assign n_n123 = ( wire944 ) | ( nsr3_3  &  (~ nrq3_2) ) | ( nsr3_3  &  wire911 ) ;
 assign wire988 = ( (~ preset)  &  ndn3_8  &  (~ ndn3_9) ) ;
 assign wire896 = ( (~ preset)  &  (~ n_n3198)  &  n_n3707  &  n_n3709 ) ;
 assign wire1016 = ( n_n3604  &  n_n3658 ) | ( n_n3604  &  (~ wire6268) ) | ( n_n3604  &  (~ n_n3658)  &  (~ n_n4335) ) | ( (~ n_n3658)  &  n_n4335  &  wire6268 ) ;
 assign wire992 = ( (~ preset)  &  ndn3_7  &  (~ ndn3_8) ) ;
 assign wire894 = ( (~ preset)  &  (~ pdn)  &  (~ nsr1_2)  &  (~ n_n3765) ) ;
 assign wire916 = ( (~ preset)  &  n_n4057  &  (~ n_n3557)  &  n_n4056 ) ;
 assign wire934 = ( (~ preset)  &  (~ n_n4126) ) ;
 assign wire1020 = ( n_n4108 ) | ( pdn  &  (~ ndn1_34) ) | ( (~ pdn)  &  nrq1_3 ) ;
 assign n_n4069 = ( n_n3916  &  wire1096 ) | ( (~ n_n3916)  &  (~ wire1096) ) ;
 assign n_n4015 = ( n_n3363  &  n_n3362  &  wire1129 ) | ( n_n3363  &  (~ wire941)  &  wire1129 ) | ( n_n3362  &  (~ wire941)  &  wire1129 ) | ( (~ n_n3363)  &  (~ n_n3362)  &  (~ wire1129) ) | ( (~ n_n3363)  &  wire941  &  (~ wire1129) ) | ( (~ n_n3362)  &  wire941  &  (~ wire1129) ) ;
 assign wire1004 = ( (~ preset)  &  (~ ndn3_10)  &  nen3_10 ) ;
 assign wire990 = ( (~ preset)  &  ndn3_6  &  (~ ndn3_7) ) ;
 assign wire1021 = ( ndn3_4 ) | ( (~ nsr3_3) ) | ( pready_0_0_  &  nrq3_2 ) ;
 assign wire994 = ( (~ nsr3_3)  &  wire6284 ) | ( pready_0_0_  &  nrq3_2  &  wire6284 ) ;
 assign n_n3563 = ( (~ n_n4360)  &  wire906 ) | ( n_n3653  &  wire906 ) | ( (~ n_n4360)  &  n_n3653  &  wire905 ) ;
 assign wire1022 = ( n_n4067 ) | ( n_n3788 ) | ( (~ wire6254) ) | ( (~ n_n4067)  &  n_n3830 ) ;
 assign wire1002 = ( (~ preset)  &  (~ ndn3_15)  &  ngfdn_3 ) ;
 assign wire997 = ( (~ preset)  &  ndn3_5  &  (~ ndn3_6) ) ;
 assign wire1006 = ( (~ preset)  &  n_n4126 ) | ( (~ preset)  &  n_n3500 ) ;
 assign wire999 = ( (~ preset)  &  ndn3_4  &  (~ ndn3_5) ) ;
 assign nak3_17 = ( (~ n_n4093) ) | ( n_n3788  &  wire1013 ) | ( wire1013  &  wire2264 ) ;
 assign n_n4038 = ( (~ n_n3916)  &  n_n4040  &  n_n4039  &  wire1096 ) | ( n_n3916  &  (~ n_n4040)  &  n_n4039  &  wire1096 ) | ( n_n3916  &  n_n4040  &  (~ n_n4039)  &  wire1096 ) | ( (~ n_n3916)  &  (~ n_n4040)  &  (~ n_n4039)  &  wire1096 ) | ( n_n3916  &  n_n4040  &  n_n4039  &  (~ wire1096) ) | ( (~ n_n3916)  &  (~ n_n4040)  &  n_n4039  &  (~ wire1096) ) | ( (~ n_n3916)  &  n_n4040  &  (~ n_n4039)  &  (~ wire1096) ) | ( n_n3916  &  (~ n_n4040)  &  (~ n_n4039)  &  (~ wire1096) ) ;
 assign n_n3653 = ( n_n3841  &  wire1078 ) | ( (~ n_n3841)  &  (~ wire1078) ) ;
 assign wire944 = ( preset ) | ( pdn ) ;
 assign wire1028 = ( nlc1_2 ) | ( (~ preset_0_0_)  &  (~ nlc1_2)  &  nsr1_2 ) | ( (~ preset_0_0_)  &  nsr1_2  &  n_n4151 ) ;
 assign n_n4116 = ( n_n4316  &  n_n4315  &  n_n4155 ) | ( (~ n_n4316)  &  (~ n_n4315)  &  n_n4155 ) | ( (~ n_n4316)  &  n_n4315  &  (~ n_n4155) ) | ( n_n4316  &  (~ n_n4315)  &  (~ n_n4155) ) ;
 assign n_n3689 = ( (~ n_n3988)  &  n_n3898  &  wire1076  &  n_n3622 ) | ( n_n3988  &  (~ n_n3898)  &  wire1076  &  n_n3622 ) | ( n_n3988  &  n_n3898  &  (~ wire1076)  &  n_n3622 ) | ( (~ n_n3988)  &  (~ n_n3898)  &  (~ wire1076)  &  n_n3622 ) | ( n_n3988  &  n_n3898  &  wire1076  &  (~ n_n3622) ) | ( (~ n_n3988)  &  (~ n_n3898)  &  wire1076  &  (~ n_n3622) ) | ( (~ n_n3988)  &  n_n3898  &  (~ wire1076)  &  (~ n_n3622) ) | ( n_n3988  &  (~ n_n3898)  &  (~ wire1076)  &  (~ n_n3622) ) ;
 assign wire1014 = ( n_n4012  &  wire896  &  wire1012  &  wire6330 ) ;
 assign n_n4158 = ( n_n4345  &  n_n4019  &  wire1086 ) | ( n_n4345  &  n_n3884  &  wire1086 ) | ( n_n4019  &  n_n3884  &  wire1086 ) | ( (~ n_n4345)  &  (~ n_n4019)  &  (~ wire1086) ) | ( (~ n_n4345)  &  (~ n_n3884)  &  (~ wire1086) ) | ( (~ n_n4019)  &  (~ n_n3884)  &  (~ wire1086) ) ;
 assign wire973 = ( pready_0_0_ ) | ( (~ pready_0_0_) ) | ( (~ nsr3_3) ) | ( (~ nrq3_2) ) | ( wire6333 ) ;
 assign wire1041 = ( n_n4067 ) | ( (~ n_n3788)  &  (~ n_n3830)  &  wire6254 ) ;
 assign n_n4079 = ( n_n4145  &  wire1075 ) | ( (~ n_n4145)  &  (~ wire1075) ) ;
 assign wire1012 = ( n_n3724  &  n_n4227  &  n_n3814 ) ;
 assign wire1042 = ( wire947 ) | ( wire1582 ) | ( wire1584 ) | ( wire1586 ) ;
 assign n_n3745 = ( n_n3898  &  wire1076 ) | ( (~ n_n3898)  &  (~ wire1076) ) ;
 assign nrq1_3 = ( (~ nsr1_2) ) | ( preset_0_0_  &  (~ nlc1_2) ) | ( nlc1_2  &  (~ n_n4151) ) ;
 assign n_n3741 = ( (~ n_n4160)  &  n_n4222  &  (~ n_n4159) ) | ( n_n4160  &  (~ n_n4222)  &  (~ n_n4159) ) | ( (~ n_n4160)  &  n_n4222  &  n_n4159  &  n_n3976 ) | ( n_n4160  &  (~ n_n4222)  &  n_n4159  &  n_n3976 ) | ( n_n4160  &  n_n4222  &  n_n4159  &  (~ n_n3976) ) | ( (~ n_n4160)  &  (~ n_n4222)  &  n_n4159  &  (~ n_n3976) ) ;
 assign wire982 = ( wire1726 ) | ( (~ n_n3832)  &  wire6257 ) | ( (~ wire6255)  &  wire6257 ) ;
 assign n_n4256 = ( n_n4229  &  wire1079 ) | ( (~ n_n4229)  &  (~ wire1079) ) ;
 assign wire947 = ( wire1588 ) | ( (~ n_n3832)  &  wire6257 ) | ( (~ wire6255)  &  wire6257 ) ;
 assign n_n4084 = ( (~ n_n4229)  &  n_n3818  &  wire1079  &  n_n3595 ) | ( n_n4229  &  (~ n_n3818)  &  wire1079  &  n_n3595 ) | ( n_n4229  &  n_n3818  &  (~ wire1079)  &  n_n3595 ) | ( (~ n_n4229)  &  (~ n_n3818)  &  (~ wire1079)  &  n_n3595 ) | ( n_n4229  &  n_n3818  &  wire1079  &  (~ n_n3595) ) | ( (~ n_n4229)  &  (~ n_n3818)  &  wire1079  &  (~ n_n3595) ) | ( (~ n_n4229)  &  n_n3818  &  (~ wire1079)  &  (~ n_n3595) ) | ( n_n4229  &  (~ n_n3818)  &  (~ wire1079)  &  (~ n_n3595) ) ;
 assign n_n4133 = ( (~ n_n4159)  &  n_n3976 ) | ( n_n4159  &  (~ n_n3976) ) ;
 assign nrq3_12 = ( nrq3_11  &  (~ ngfdn_3) ) ;
 assign n_n3832 = ( (~ n_n3788)  &  (~ wire2264)  &  wire6254 ) ;
 assign wire1015 = ( n_n3851  &  n_n3831  &  n_n4026 ) | ( n_n3851  &  n_n3831  &  n_n3852 ) | ( n_n3831  &  (~ n_n4026)  &  n_n3852 ) ;
 assign wire1063 = ( (~ n_n3709) ) | ( (~ wire6290) ) | ( wire1137  &  wire1136 ) ;
 assign wire1064 = ( n_n4263 ) | ( (~ nlc3_3)  &  nrq3_2  &  wire6324 ) ;
 assign wire1068 = ( n_n3656 ) | ( n_n4056  &  n_n4098 ) | ( n_n4056  &  (~ wire6349) ) ;
 assign wire923 = ( n_n3959 ) | ( n_n4159  &  n_n3976 ) | ( (~ n_n4159)  &  (~ n_n3976) ) ;
 assign wire1069 = ( wire1173 ) | ( (~ n_n3832)  &  wire6257 ) | ( (~ wire6255)  &  wire6257 ) ;
 assign n_n4297 = ( (~ n_n4145)  &  n_n4080  &  wire1075  &  n_n4078 ) | ( n_n4145  &  (~ n_n4080)  &  wire1075  &  n_n4078 ) | ( n_n4145  &  n_n4080  &  (~ wire1075)  &  n_n4078 ) | ( (~ n_n4145)  &  (~ n_n4080)  &  (~ wire1075)  &  n_n4078 ) | ( n_n4145  &  n_n4080  &  wire1075  &  (~ n_n4078) ) | ( (~ n_n4145)  &  (~ n_n4080)  &  wire1075  &  (~ n_n4078) ) | ( (~ n_n4145)  &  n_n4080  &  (~ wire1075)  &  (~ n_n4078) ) | ( n_n4145  &  (~ n_n4080)  &  (~ wire1075)  &  (~ n_n4078) ) ;
 assign n_n4126 = ( n_n4056  &  wire6270 ) | ( (~ n_n4056)  &  n_n4367  &  wire6268 ) ;
 assign wire1070 = ( (~ n_n4222)  &  (~ n_n3934)  &  n_n4125 ) | ( (~ n_n4222)  &  (~ n_n3976)  &  n_n4125 ) | ( n_n4222  &  (~ n_n3934)  &  (~ n_n4125) ) | ( n_n4222  &  (~ n_n3976)  &  (~ n_n4125) ) | ( n_n4222  &  n_n3934  &  n_n3976  &  n_n4125 ) | ( (~ n_n4222)  &  n_n3934  &  n_n3976  &  (~ n_n4125) ) ;
 assign wire935 = ( n_n4160 ) | ( n_n4383 ) | ( n_n4159 ) ;
 assign n_n3765 = ( preset_0_0_  &  (~ nlc1_2) ) | ( nlc1_2  &  (~ n_n4151) ) ;
 assign n_n4367 = ( n_n3604  &  n_n3658 ) | ( (~ n_n3658)  &  wire6265 ) | ( (~ n_n3658)  &  wire6266 ) ;
 assign wire984 = ( n_n3955 ) | ( (~ n_n3954) ) | ( n_n4029 ) | ( n_n3845 ) ;
 assign n_n4335 = ( wire6265 ) | ( wire6266 ) ;
 assign wire899 = ( n_n4069  &  n_n4082 ) | ( (~ n_n4038)  &  n_n4082 ) | ( n_n4069  &  (~ n_n4038)  &  n_n3986 ) ;
 assign n_n3786 = ( (~ n_n3689)  &  wire899 ) | ( n_n3745  &  wire899 ) | ( (~ n_n3689)  &  n_n3745  &  wire900 ) ;
 assign wire1075 = ( n_n3898  &  n_n4144  &  n_n4223 ) | ( (~ n_n3898)  &  (~ n_n4144)  &  (~ n_n4223) ) | ( n_n3898  &  n_n4144  &  n_n4034 ) | ( n_n4144  &  n_n4223  &  n_n4034 ) | ( (~ n_n3898)  &  (~ n_n4144)  &  (~ n_n4034) ) | ( (~ n_n4144)  &  (~ n_n4223)  &  (~ n_n4034) ) ;
 assign wire1076 = ( n_n3916  &  n_n4223  &  n_n3420 ) | ( (~ n_n3916)  &  (~ n_n4223)  &  (~ n_n3420) ) | ( n_n3916  &  n_n4223  &  n_n4267 ) | ( n_n4223  &  n_n3420  &  n_n4267 ) | ( (~ n_n3916)  &  (~ n_n4223)  &  (~ n_n4267) ) | ( (~ n_n4223)  &  (~ n_n3420)  &  (~ n_n4267) ) ;
 assign n_n3788 = ( (~ n_n3833)  &  n_n4067 ) | ( (~ n_n4067)  &  n_n3563 ) ;
 assign n_n4305 = ( n_n4057  &  (~ n_n3557)  &  n_n4056 ) ;
 assign n_n3656 = ( (~ n_n4056)  &  n_n4367  &  wire6268 ) ;
 assign n_n3500 = ( (~ n_n3493)  &  (~ n_n4045) ) | ( (~ n_n3493)  &  (~ n_n4367)  &  wire6299 ) ;
 assign wire1078 = ( n_n4145  &  n_n4144  &  n_n4268 ) | ( n_n4145  &  n_n4259  &  n_n4268 ) | ( n_n4144  &  n_n4259  &  n_n4268 ) | ( (~ n_n4145)  &  (~ n_n4144)  &  (~ n_n4268) ) | ( (~ n_n4145)  &  (~ n_n4259)  &  (~ n_n4268) ) | ( (~ n_n4144)  &  (~ n_n4259)  &  (~ n_n4268) ) ;
 assign wire1079 = ( n_n4316  &  n_n4181  &  n_n4315 ) | ( (~ n_n4316)  &  (~ n_n4181)  &  (~ n_n4315) ) | ( n_n4316  &  n_n4181  &  n_n4155 ) | ( n_n4181  &  n_n4315  &  n_n4155 ) | ( (~ n_n4316)  &  (~ n_n4181)  &  (~ n_n4155) ) | ( (~ n_n4181)  &  (~ n_n4315)  &  (~ n_n4155) ) ;
 assign wire1013 = ( nen3_10  &  nsr3_17 ) ;
 assign nrq3_15 = ( (~ ndn3_15)  &  ngfdn_3 ) ;
 assign n_n3363 = ( wire2189 ) | ( wire2190 ) | ( wire2191 ) ;
 assign n_n3362 = ( wire6275 ) | ( nrq3_11  &  (~ ngfdn_3)  &  n_n3741 ) ;
 assign n_n4078 = ( n_n3988  &  n_n3622 ) | ( n_n3988  &  (~ n_n3898)  &  wire1076 ) | ( n_n3988  &  n_n3898  &  (~ wire1076) ) | ( (~ n_n3898)  &  wire1076  &  n_n3622 ) | ( n_n3898  &  (~ wire1076)  &  n_n3622 ) ;
 assign n_n3888 = ( n_n4080  &  n_n4078 ) | ( (~ n_n4145)  &  n_n4080  &  wire1075 ) | ( n_n4145  &  n_n4080  &  (~ wire1075) ) | ( (~ n_n4145)  &  wire1075  &  n_n4078 ) | ( n_n4145  &  (~ wire1075)  &  n_n4078 ) ;
 assign n_n4345 = ( n_n4169  &  n_n4168 ) | ( n_n4169  &  wire2049 ) | ( n_n4168  &  wire2049 ) | ( n_n4169  &  wire2050 ) | ( n_n4168  &  wire2050 ) ;
 assign n_n4019 = ( wire6296 ) | ( n_n3916  &  nrq3_12  &  wire1096 ) | ( (~ n_n3916)  &  nrq3_12  &  (~ wire1096) ) ;
 assign n_n3884 = ( wire2035 ) | ( wire2036 ) | ( wire2037 ) ;
 assign wire1086 = ( n_n3334  &  wire1903 ) | ( n_n3334  &  wire1904 ) | ( n_n3334  &  wire1905 ) | ( (~ n_n3334)  &  (~ wire1903)  &  (~ wire1904)  &  (~ wire1905) ) ;
 assign n_n4039 = ( n_n3818  &  n_n3595 ) | ( (~ n_n4229)  &  n_n3818  &  wire1079 ) | ( n_n4229  &  n_n3818  &  (~ wire1079) ) | ( (~ n_n4229)  &  wire1079  &  n_n3595 ) | ( n_n4229  &  (~ wire1079)  &  n_n3595 ) ;
 assign n_n3622 = ( n_n4040  &  n_n4039 ) | ( (~ n_n3916)  &  n_n4040  &  wire1096 ) | ( (~ n_n3916)  &  n_n4039  &  wire1096 ) | ( n_n3916  &  n_n4040  &  (~ wire1096) ) | ( n_n3916  &  n_n4039  &  (~ wire1096) ) ;
 assign n_n3981 = ( wire2175 ) | ( wire2176 ) | ( wire2177 ) ;
 assign wire1088 = ( n_n3981 ) | ( wire2174 ) | ( wire6281 ) ;
 assign n_n3294 = ( n_n3865  &  wire984 ) | ( (~ n_n3865)  &  (~ wire984) ) ;
 assign n_n3334 = ( wire6317 ) | ( n_n3898  &  nrq3_12  &  wire1076 ) | ( (~ n_n3898)  &  nrq3_12  &  (~ wire1076) ) ;
 assign n_n4296 = ( (~ n_n3198)  &  n_n3707  &  n_n3709 ) ;
 assign n_n3324 = ( wire6312 ) | ( n_n3841  &  nrq3_12  &  wire1078 ) | ( (~ n_n3841)  &  nrq3_12  &  (~ wire1078) ) ;
 assign n_n3243 = ( wire1908 ) | ( wire1909 ) | ( wire1910 ) ;
 assign n_n3830 = ( (~ n_n3851)  &  n_n4026 ) | ( (~ n_n4026)  &  (~ n_n3852) ) ;
 assign n_n3869 = ( n_n3916  &  n_n4047 ) | ( n_n3916  &  n_n3870 ) | ( n_n4047  &  n_n3870 ) ;
 assign n_n3205 = ( n_n4366  &  n_n3898 ) | ( n_n4366  &  n_n3869 ) | ( n_n3898  &  n_n3869 ) ;
 assign wire901 = ( (~ n_n3876)  &  n_n4231 ) | ( n_n4069  &  n_n4231 ) | ( (~ n_n3876)  &  n_n4069  &  n_n4254 ) ;
 assign n_n3240 = ( (~ n_n4362)  &  wire901 ) | ( n_n3745  &  wire901 ) | ( (~ n_n4362)  &  n_n3745  &  wire907 ) ;
 assign n_n4181 = ( n_n4160  &  (~ n_n4182) ) | ( n_n4383  &  (~ n_n4182) ) | ( n_n4159  &  (~ n_n4182) ) | ( (~ n_n4160)  &  (~ n_n4383)  &  (~ n_n4159)  &  n_n4182 ) ;
 assign wire1094 = ( n_n4096  &  wire1892 ) | ( n_n4096  &  wire1893 ) | ( n_n4096  &  wire1894 ) | ( (~ n_n4096)  &  (~ wire1892)  &  (~ wire1893)  &  (~ wire1894) ) ;
 assign n_n3870 = ( n_n4229  &  n_n3769 ) | ( n_n4229  &  n_n3899 ) | ( n_n3769  &  n_n3899 ) ;
 assign wire1096 = ( n_n4229  &  n_n4181  &  n_n3420 ) | ( (~ n_n4229)  &  (~ n_n4181)  &  (~ n_n3420) ) | ( n_n4229  &  n_n3420  &  n_n3923 ) | ( n_n4181  &  n_n3420  &  n_n3923 ) | ( (~ n_n4229)  &  (~ n_n3420)  &  (~ n_n3923) ) | ( (~ n_n4181)  &  (~ n_n3420)  &  (~ n_n3923) ) ;
 assign n_n4144 = ( n_n4224  &  (~ n_n4251) ) | ( (~ n_n4251)  &  wire935 ) | ( (~ n_n4251)  &  (~ wire6251) ) | ( (~ n_n4224)  &  n_n4251  &  (~ wire935)  &  wire6251 ) ;
 assign n_n4223 = ( (~ n_n4224)  &  n_n4330 ) | ( (~ n_n4224)  &  n_n4182 ) | ( (~ n_n4224)  &  wire935 ) | ( n_n4224  &  (~ n_n4330)  &  (~ n_n4182)  &  (~ wire935) ) ;
 assign n_n4034 = ( n_n3916  &  n_n4267 ) | ( n_n3916  &  (~ n_n4330)  &  wire1116 ) | ( n_n3916  &  n_n4330  &  (~ wire1116) ) | ( (~ n_n4330)  &  wire1116  &  n_n4267 ) | ( n_n4330  &  (~ wire1116)  &  n_n4267 ) ;
 assign n_n4259 = ( n_n3898  &  n_n4223 ) | ( n_n3898  &  n_n4034 ) | ( n_n4223  &  n_n4034 ) ;
 assign n_n3900 = ( n_n4222  &  n_n4125 ) | ( n_n4222  &  n_n3934  &  n_n3976 ) | ( n_n3934  &  n_n3976  &  n_n4125 ) ;
 assign n_n3124 = ( (~ n_n3959)  &  (~ n_n3741) ) | ( (~ n_n3741)  &  (~ n_n4133) ) | ( n_n3574  &  n_n3959  &  (~ n_n3741) ) | ( (~ n_n3574)  &  n_n3741  &  (~ n_n4133) ) | ( n_n3574  &  (~ n_n3959)  &  n_n3741  &  n_n4133 ) ;
 assign n_n135 = ( (~ n_n3653)  &  wire1137 ) | ( (~ n_n3726)  &  n_n3653  &  n_n3888  &  wire1137 ) | ( n_n3726  &  n_n3653  &  (~ n_n3888)  &  wire1137 ) ;
 assign n_n4315 = ( n_n4160  &  (~ n_n4383) ) | ( (~ n_n4383)  &  n_n4159 ) | ( (~ n_n4160)  &  n_n4383  &  (~ n_n4159) ) ;
 assign wire1104 = ( n_n3334 ) | ( wire1903 ) | ( wire1904 ) | ( wire1905 ) ;
 assign n_n4096 = ( wire6318 ) | ( n_n4145  &  nrq3_12  &  wire1075 ) | ( (~ n_n4145)  &  nrq3_12  &  (~ wire1075) ) ;
 assign wire904 = ( (~ n_n4116)  &  n_n3124 ) | ( (~ n_n3995)  &  n_n4116  &  n_n3124  &  n_n3994 ) | ( n_n3995  &  (~ n_n4116)  &  (~ n_n3124)  &  n_n3994 ) | ( n_n3995  &  n_n4116  &  n_n3124  &  (~ n_n3994) ) | ( (~ n_n3995)  &  (~ n_n4116)  &  (~ n_n3124)  &  (~ n_n3994) ) ;
 assign n_n3986 = ( (~ n_n4256)  &  wire904 ) | ( n_n4084  &  wire904 ) | ( (~ n_n4256)  &  n_n4084  &  wire903 ) ;
 assign n_n3994 = ( n_n3574  &  (~ n_n3741) ) | ( n_n3574  &  wire923 ) | ( (~ n_n3741)  &  wire923 ) ;
 assign n_n3595 = ( n_n3995  &  (~ n_n4116) ) | ( n_n3995  &  n_n3994 ) | ( (~ n_n4116)  &  n_n3994 ) ;
 assign n_n4357 = ( n_n4381  &  n_n4052 ) | ( n_n4381  &  n_n3865 ) | ( n_n4381  &  wire984 ) | ( (~ n_n4381)  &  (~ n_n4052)  &  (~ n_n3865)  &  (~ wire984) ) ;
 assign wire1109 = ( n_n4224 ) | ( n_n4251 ) | ( wire935 ) | ( (~ wire6251) ) ;
 assign n_n4268 = ( (~ n_n4270)  &  wire1109 ) | ( n_n4270  &  (~ wire1109) ) ;
 assign n_n4006 = ( n_n3955  &  n_n4029 ) | ( (~ n_n3954)  &  n_n4029 ) | ( n_n4029  &  n_n3845 ) | ( (~ n_n3955)  &  n_n3954  &  (~ n_n4029)  &  (~ n_n3845) ) ;
 assign n_n3848 = ( n_n3955  &  n_n3845 ) | ( (~ n_n3954)  &  n_n3845 ) | ( (~ n_n3955)  &  n_n3954  &  (~ n_n3845) ) ;
 assign n_n4098 = ( n_n4099  &  wire1119 ) | ( (~ n_n4099)  &  (~ wire1119) ) ;
 assign wire942 = ( (~ n_n4052)  &  n_n3865 ) | ( (~ n_n4052)  &  wire984 ) | ( n_n4052  &  (~ n_n3865)  &  (~ wire984) ) ;
 assign wire1110 = ( n_n4169  &  wire2045 ) | ( n_n4169  &  wire6295 ) | ( (~ n_n4169)  &  (~ wire2045)  &  (~ wire6295) ) ;
 assign n_n3852 = ( n_n4360  &  wire905 ) | ( (~ n_n3653)  &  wire905 ) | ( n_n4360  &  (~ n_n3653)  &  wire906 ) ;
 assign wire903 = ( n_n4116  &  (~ n_n3124) ) | ( n_n3995  &  n_n4116  &  n_n3124  &  n_n3994 ) | ( (~ n_n3995)  &  (~ n_n4116)  &  (~ n_n3124)  &  n_n3994 ) | ( (~ n_n3995)  &  n_n4116  &  n_n3124  &  (~ n_n3994) ) | ( n_n3995  &  (~ n_n4116)  &  (~ n_n3124)  &  (~ n_n3994) ) ;
 assign n_n4082 = ( n_n4256  &  wire903 ) | ( (~ n_n4084)  &  wire903 ) | ( n_n4256  &  (~ n_n4084)  &  wire904 ) ;
 assign nrq3_2 = ( (~ preset_0_0_)  &  (~ nlc1_2)  &  nsr1_2 ) | ( (~ preset_0_0_)  &  nsr1_2  &  n_n4151 ) | ( nlc1_2  &  nsr1_2  &  n_n4151 ) ;
 assign n_n4169 = ( wire2046 ) | ( wire2047 ) | ( wire2048 ) ;
 assign n_n4168 = ( wire6295 ) | ( n_n4229  &  nrq3_12  &  wire1079 ) | ( (~ n_n4229)  &  nrq3_12  &  (~ wire1079) ) ;
 assign n_n4155 = ( (~ n_n4160)  &  n_n4222  &  n_n4159 ) | ( n_n4160  &  n_n4222  &  (~ n_n4159) ) | ( (~ n_n4160)  &  n_n4159  &  n_n3976 ) | ( n_n4222  &  n_n4159  &  n_n3976 ) ;
 assign wire905 = ( n_n4299  &  n_n3253 ) | ( (~ n_n4079)  &  n_n3253 ) | ( n_n4299  &  (~ n_n4079)  &  n_n3240 ) ;
 assign wire1116 = ( n_n4160 ) | ( n_n4383 ) | ( n_n4159 ) | ( n_n4182 ) ;
 assign n_n3420 = ( (~ n_n4330)  &  wire1116 ) | ( n_n4330  &  (~ wire1116) ) ;
 assign wire902 = ( (~ n_n3946)  &  n_n3927 ) | ( n_n4116  &  n_n3927 ) | ( (~ n_n3946)  &  n_n4116  &  (~ n_n3927) ) ;
 assign n_n4231 = ( (~ n_n4258)  &  wire902 ) | ( n_n4256  &  wire902 ) | ( (~ n_n4258)  &  n_n4256  &  wire908 ) ;
 assign wire907 = ( n_n3876  &  n_n4254 ) | ( (~ n_n4069)  &  n_n4254 ) | ( n_n3876  &  (~ n_n4069)  &  n_n4231 ) ;
 assign n_n3253 = ( n_n4362  &  wire907 ) | ( (~ n_n3745)  &  wire907 ) | ( n_n4362  &  (~ n_n3745)  &  wire901 ) ;
 assign wire1119 = ( n_n4381 ) | ( n_n4052 ) | ( n_n3865 ) | ( wire984 ) ;
 assign wire900 = ( (~ n_n4069)  &  n_n3986 ) | ( n_n4038  &  n_n3986 ) | ( (~ n_n4069)  &  n_n4038  &  n_n4082 ) ;
 assign n_n3785 = ( n_n3689  &  wire900 ) | ( (~ n_n3745)  &  wire900 ) | ( n_n3689  &  (~ n_n3745)  &  wire899 ) ;
 assign n_n4097 = ( wire1892 ) | ( wire1893 ) | ( wire1894 ) ;
 assign wire941 = ( (~ n_n3974) ) | ( (~ wire2183)  &  (~ wire2184)  &  (~ wire2185) ) ;
 assign n_n3975 = ( wire2183 ) | ( wire2184 ) | ( wire2185 ) ;
 assign n_n3974 = ( wire6278 ) | ( n_n3934  &  n_n4367  &  nrq3_15 ) ;
 assign wire1122 = ( n_n4019  &  wire2035 ) | ( n_n4019  &  wire2036 ) | ( n_n4019  &  wire2037 ) | ( (~ n_n4019)  &  (~ wire2035)  &  (~ wire2036)  &  (~ wire2037) ) ;
 assign n_n4267 = ( n_n4229  &  n_n4181 ) | ( n_n4229  &  n_n3923 ) | ( n_n4181  &  n_n3923 ) ;
 assign n_n3899 = ( n_n4316  &  n_n3901 ) | ( n_n4316  &  n_n3900 ) | ( n_n3901  &  n_n3900 ) ;
 assign wire906 = ( (~ n_n4299)  &  n_n3240 ) | ( n_n4079  &  n_n3240 ) | ( (~ n_n4299)  &  n_n4079  &  n_n3253 ) ;
 assign wire1128 = ( n_n3975  &  n_n3974  &  wire2188 ) | ( n_n3975  &  n_n3974  &  wire6275 ) | ( (~ n_n3975)  &  (~ wire2188)  &  (~ wire6275) ) | ( (~ n_n3974)  &  (~ wire2188)  &  (~ wire6275) ) ;
 assign wire1129 = ( n_n3981  &  wire2174 ) | ( n_n3981  &  wire6281 ) | ( (~ n_n3981)  &  (~ wire2174)  &  (~ wire6281) ) ;
 assign wire908 = ( n_n3946  &  (~ n_n3927) ) | ( (~ n_n4116)  &  (~ n_n3927) ) | ( n_n3946  &  (~ n_n4116)  &  n_n3927 ) ;
 assign n_n4254 = ( n_n4258  &  wire908 ) | ( (~ n_n4256)  &  wire908 ) | ( n_n4258  &  (~ n_n4256)  &  wire902 ) ;
 assign n_n3923 = ( n_n4316  &  n_n4315 ) | ( n_n4316  &  n_n4155 ) | ( n_n4315  &  n_n4155 ) ;
 assign wire1137 = ( (~ n_n4079)  &  n_n3785 ) | ( n_n4297  &  n_n3785 ) | ( (~ n_n4079)  &  n_n4297  &  n_n3786 ) ;
 assign wire1136 = ( (~ n_n3841)  &  wire1078 ) | ( n_n3841  &  (~ wire1078) ) | ( (~ n_n3726)  &  n_n3841  &  wire1078  &  n_n3888 ) | ( (~ n_n3726)  &  (~ n_n3841)  &  (~ wire1078)  &  n_n3888 ) | ( n_n3726  &  n_n3841  &  wire1078  &  (~ n_n3888) ) | ( n_n3726  &  (~ n_n3841)  &  (~ wire1078)  &  (~ n_n3888) ) ;
 assign n_n3927 = ( (~ n_n3743)  &  n_n3741 ) | ( (~ n_n3743)  &  wire6250 ) | ( n_n3741  &  wire6250 ) ;
 assign wire914 = ( (~ n_n4096)  &  (~ n_n4097) ) | ( (~ n_n4096)  &  (~ wire1898)  &  (~ wire1899) ) | ( (~ n_n4097)  &  (~ wire1898)  &  (~ wire1899) ) ;
 assign wire936 = ( n_n3788 ) | ( wire2264 ) | ( (~ wire6254) ) | ( wire6309 ) ;
 assign wire1155 = ( ndn3_4 ) | ( (~ pready_0_0_)  &  nsr3_3 ) | ( nsr3_3  &  (~ nrq3_2) ) ;
 assign wire1008 = ( (~ n_n3493)  &  (~ n_n4045)  &  n_n4367 ) ;
 assign wire1019 = ( n_n4366  &  n_n4145  &  n_n3898 ) | ( (~ n_n4366)  &  (~ n_n4145)  &  (~ n_n3898) ) | ( n_n4366  &  n_n4145  &  n_n3869 ) | ( n_n4145  &  n_n3898  &  n_n3869 ) | ( (~ n_n4366)  &  (~ n_n4145)  &  (~ n_n3869) ) | ( (~ n_n4145)  &  (~ n_n3898)  &  (~ n_n3869) ) ;
 assign wire1034 = ( n_n3916  &  n_n4047  &  n_n3898 ) | ( (~ n_n3916)  &  (~ n_n4047)  &  (~ n_n3898) ) | ( n_n3916  &  n_n3898  &  n_n3870 ) | ( n_n4047  &  n_n3898  &  n_n3870 ) | ( (~ n_n3916)  &  (~ n_n3898)  &  (~ n_n3870) ) | ( (~ n_n4047)  &  (~ n_n3898)  &  (~ n_n3870) ) ;
 assign wire1038 = ( n_n4047  &  n_n4229  &  n_n3769 ) | ( (~ n_n4047)  &  (~ n_n4229)  &  (~ n_n3769) ) | ( n_n4047  &  n_n4229  &  n_n3899 ) | ( n_n4047  &  n_n3769  &  n_n3899 ) | ( (~ n_n4047)  &  (~ n_n4229)  &  (~ n_n3899) ) | ( (~ n_n4047)  &  (~ n_n3769)  &  (~ n_n3899) ) ;
 assign wire1051 = ( n_n4316  &  n_n3769  &  n_n3901 ) | ( (~ n_n4316)  &  (~ n_n3769)  &  (~ n_n3901) ) | ( n_n4316  &  n_n3769  &  n_n3900 ) | ( n_n3769  &  n_n3901  &  n_n3900 ) | ( (~ n_n4316)  &  (~ n_n3769)  &  (~ n_n3900) ) | ( (~ n_n3769)  &  (~ n_n3901)  &  (~ n_n3900) ) ;
 assign wire1062 = ( n_n3475  &  n_n4145  &  n_n3841 ) | ( (~ n_n3475)  &  (~ n_n4145)  &  (~ n_n3841) ) | ( n_n3475  &  n_n3841  &  n_n3205 ) | ( n_n4145  &  n_n3841  &  n_n3205 ) | ( (~ n_n3475)  &  (~ n_n3841)  &  (~ n_n3205) ) | ( (~ n_n4145)  &  (~ n_n3841)  &  (~ n_n3205) ) ;
 assign wire1082 = ( (~ n_n3707) ) | ( (~ n_n3851)  &  n_n4026 ) | ( (~ n_n4026)  &  (~ n_n3852) ) ;
 assign wire911 = ( (~ tin_pready_0_0_)  &  (~ n_n4108)  &  nsr4_2 ) | ( (~ tin_pready_0_0_)  &  (~ n_n3354)  &  nsr4_2 ) | ( n_n4108  &  (~ n_n3354)  &  nsr4_2 ) ;
 assign wire921 = ( (~ preset)  &  (~ n_n3831) ) | ( (~ preset)  &  wire922 ) | ( (~ preset)  &  wire937 ) ;
 assign wire922 = ( (~ n_n3788)  &  (~ wire2264)  &  wire6254  &  wire6387 ) ;
 assign wire937 = ( (~ n_n3788)  &  wire1082  &  (~ wire2264)  &  wire6254 ) ;
 assign wire946 = ( n_n3814  &  (~ n_n3832)  &  wire6257 ) | ( n_n3814  &  (~ wire6255)  &  wire6257 ) ;
 assign wire971 = ( (~ preset)  &  pdn  &  n_n3806 ) | ( (~ preset)  &  n_n3806  &  (~ nrq1_3) ) ;
 assign wire974 = ( (~ preset)  &  pdn  &  n_n3537 ) | ( (~ preset)  &  n_n3537  &  (~ nrq1_3) ) ;
 assign wire976 = ( (~ preset)  &  (~ nrq3_11)  &  n_n3099 ) | ( (~ preset)  &  ngfdn_3  &  n_n3099 ) ;
 assign wire978 = ( (~ preset)  &  pdn  &  n_n3646 ) | ( (~ preset)  &  n_n3646  &  (~ nrq1_3) ) ;
 assign wire983 = ( (~ preset)  &  pdn  &  n_n3739 ) | ( (~ preset)  &  n_n3739  &  (~ nrq1_3) ) ;
 assign wire1165 = ( (~ preset)  &  n_n4299  &  n_n3832  &  wire6255 ) ;
 assign wire1166 = ( n_n4080  &  (~ n_n3832)  &  wire6257 ) | ( n_n4080  &  (~ wire6255)  &  wire6257 ) ;
 assign wire1167 = ( (~ n_n4080)  &  wire896  &  n_n4079  &  n_n4078 ) | ( n_n4080  &  wire896  &  (~ n_n4079)  &  n_n4078 ) | ( n_n4080  &  wire896  &  n_n4079  &  (~ n_n4078) ) | ( (~ n_n4080)  &  wire896  &  (~ n_n4079)  &  (~ n_n4078) ) ;
 assign wire1168 = ( (~ preset)  &  ndn3_15  &  n_n3608 ) | ( (~ preset)  &  (~ ngfdn_3)  &  n_n3608 ) ;
 assign wire1171 = ( (~ preset)  &  n_n3756  &  n_n3832  &  wire6255 ) ;
 assign wire1172 = ( (~ n_n4159)  &  n_n3976  &  (~ n_n3959)  &  wire896 ) | ( n_n4159  &  (~ n_n3976)  &  (~ n_n3959)  &  wire896 ) ;
 assign wire1173 = ( n_n4159  &  n_n3976  &  wire896 ) | ( (~ n_n4159)  &  (~ n_n3976)  &  wire896 ) ;
 assign wire1179 = ( (~ preset)  &  pdn  &  n_n3486 ) | ( (~ preset)  &  n_n3486  &  (~ nrq1_3) ) ;
 assign wire1182 = ( (~ preset)  &  n_n3865  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1184 = ( n_n3922  &  n_n3656 ) | ( n_n3922  &  wire2011 ) ;
 assign wire1187 = ( (~ preset)  &  n_n3845  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1189 = ( n_n3968  &  n_n3656 ) | ( n_n3968  &  wire2011 ) ;
 assign wire1191 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3931 ) | ( (~ preset)  &  ndn3_5  &  n_n3931 ) ;
 assign wire1195 = ( (~ preset)  &  n_n3878  &  wire1155 ) ;
 assign wire1199 = ( (~ preset)  &  pdn  &  n_n4180 ) | ( (~ preset)  &  n_n4180  &  (~ nrq1_3) ) ;
 assign wire1201 = ( (~ preset)  &  pdn  &  n_n3277 ) | ( (~ preset)  &  n_n3277  &  (~ nrq1_3) ) ;
 assign wire1204 = ( (~ preset)  &  pdn  &  n_n4102 ) | ( (~ preset)  &  n_n4102  &  (~ nrq1_3) ) ;
 assign wire1206 = ( (~ preset)  &  pdn  &  n_n4342 ) | ( (~ preset)  &  n_n4342  &  (~ nrq1_3) ) ;
 assign wire1208 = ( wire1015  &  (~ n_n3788)  &  (~ wire2264)  &  wire6254 ) ;
 assign wire1212 = ( (~ preset)  &  ndn3_10  &  n_n3841 ) | ( (~ preset)  &  (~ nen3_10)  &  n_n3841 ) ;
 assign wire1213 = ( wire1004  &  (~ n_n3324)  &  n_n3243  &  wire914 ) | ( wire1004  &  n_n3324  &  (~ n_n3243)  &  wire914 ) | ( wire1004  &  n_n3324  &  n_n3243  &  (~ wire914) ) | ( wire1004  &  (~ n_n3324)  &  (~ n_n3243)  &  (~ wire914) ) ;
 assign wire1214 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4182 ) | ( (~ preset)  &  ndn3_6  &  n_n4182 ) ;
 assign wire1218 = ( (~ preset)  &  pdn  &  n_n3413 ) | ( (~ preset)  &  n_n3413  &  (~ nrq1_3) ) ;
 assign wire1225 = ( n_n3831  &  n_n3788 ) | ( n_n3831  &  wire2264 ) | ( n_n3831  &  (~ wire6254) ) ;
 assign wire1230 = ( n_n3724  &  (~ n_n4227)  &  n_n3814  &  wire896 ) ;
 assign wire1232 = ( (~ preset)  &  pdn  &  n_n3337 ) | ( (~ preset)  &  n_n3337  &  (~ nrq1_3) ) ;
 assign wire1242 = ( (~ preset)  &  pdn  &  n_n4209 ) | ( (~ preset)  &  n_n4209  &  (~ nrq1_3) ) ;
 assign wire1246 = ( (~ preset)  &  pdn  &  n_n3342 ) | ( (~ preset)  &  n_n3342  &  (~ nrq1_3) ) ;
 assign wire1248 = ( (~ preset)  &  pdn  &  n_n3667 ) | ( (~ preset)  &  n_n3667  &  (~ nrq1_3) ) ;
 assign wire1251 = ( (~ preset)  &  (~ ndn3_7)  &  n_n3756 ) | ( (~ preset)  &  ndn3_8  &  n_n3756 ) ;
 assign wire1259 = ( (~ preset)  &  ndn3_15  &  n_n4095 ) | ( (~ preset)  &  n_n4095  &  (~ ngfdn_3) ) ;
 assign wire1260 = ( wire1002  &  wire1094  &  wire1898 ) | ( wire1002  &  wire1094  &  wire1899 ) | ( wire1002  &  (~ wire1094)  &  (~ wire1898)  &  (~ wire1899) ) ;
 assign wire1261 = ( (~ preset)  &  pdn  &  n_n3394 ) | ( (~ preset)  &  n_n3394  &  (~ nrq1_3) ) ;
 assign wire1263 = ( (~ preset)  &  ndn3_10  &  n_n3976 ) | ( (~ preset)  &  (~ nen3_10)  &  n_n3976 ) ;
 assign wire1265 = ( (~ preset)  &  pdn  &  n_n4166 ) | ( (~ preset)  &  n_n4166  &  (~ nrq1_3) ) ;
 assign wire1267 = ( (~ preset)  &  pdn  &  n_n3572 ) | ( (~ preset)  &  n_n3572  &  (~ nrq1_3) ) ;
 assign wire1270 = ( (~ preset)  &  pdn  &  n_n3514 ) | ( (~ preset)  &  n_n3514  &  (~ nrq1_3) ) ;
 assign wire1271 = ( (~ preset)  &  (~ ndn3_4)  &  n_n4062 ) | ( (~ preset)  &  ndn3_5  &  n_n4062 ) ;
 assign wire1275 = ( (~ preset)  &  (~ ndn3_4)  &  n_n4021 ) | ( (~ preset)  &  ndn3_5  &  n_n4021 ) ;
 assign wire1280 = ( n_n3766  &  wire947 ) | ( n_n3766  &  wire1584 ) | ( n_n3766  &  wire1586 ) ;
 assign wire1282 = ( (~ preset)  &  pdn  &  n_n3966 ) | ( (~ preset)  &  n_n3966  &  (~ nrq1_3) ) ;
 assign wire1283 = ( (~ preset)  &  pdn  &  n_n4199 ) | ( (~ preset)  &  n_n4199  &  (~ nrq1_3) ) ;
 assign wire1285 = ( (~ preset)  &  pdn  &  n_n4247 ) | ( (~ preset)  &  n_n4247  &  (~ nrq1_3) ) ;
 assign wire1287 = ( (~ preset)  &  (~ ndn3_7)  &  n_n4360 ) | ( (~ preset)  &  ndn3_8  &  n_n4360 ) ;
 assign wire1291 = ( (~ preset)  &  pdn  &  n_n4320 ) | ( (~ preset)  &  n_n4320  &  (~ nrq1_3) ) ;
 assign wire1295 = ( (~ preset)  &  pdn  &  n_n3108 ) | ( (~ preset)  &  n_n3108  &  (~ nrq1_3) ) ;
 assign wire1298 = ( (~ preset)  &  pdn  &  n_n3910 ) | ( (~ preset)  &  n_n3910  &  (~ nrq1_3) ) ;
 assign wire1301 = ( (~ preset)  &  pdn  &  n_n3758 ) | ( (~ preset)  &  n_n3758  &  (~ nrq1_3) ) ;
 assign wire1303 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3170 ) | ( (~ preset)  &  ndn3_9  &  n_n3170 ) ;
 assign wire1307 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3250 ) | ( (~ preset)  &  ndn3_9  &  n_n3250 ) ;
 assign wire1312 = ( (~ preset)  &  pdn  &  n_n4303 ) | ( (~ preset)  &  n_n4303  &  (~ nrq1_3) ) ;
 assign wire1315 = ( (~ preset_0_0_)  &  (~ nlc1_2)  &  nsr1_2 ) ;
 assign wire1316 = ( nlc1_2  &  n_n4151 ) | ( (~ nsr1_2)  &  n_n4151 ) | ( preset_0_0_  &  (~ nlc1_2)  &  n_n4151 ) ;
 assign wire1318 = ( nsr3_17  &  nsr3_14 ) | ( n_n4045  &  nsr3_14  &  n_n4367 ) ;
 assign wire1323 = ( (~ preset)  &  n_n4029  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1325 = ( n_n3533  &  n_n3656 ) | ( n_n3533  &  wire2011 ) ;
 assign wire1329 = ( (~ preset)  &  n_n3208  &  wire1155 ) ;
 assign wire1333 = ( (~ preset)  &  (~ nrq3_11)  &  n_n4157 ) | ( (~ preset)  &  n_n4157  &  ngfdn_3 ) ;
 assign wire1335 = ( (~ preset)  &  (~ ndn3_7)  &  n_n4299 ) | ( (~ preset)  &  ndn3_8  &  n_n4299 ) ;
 assign wire1339 = ( (~ preset)  &  pdn  &  n_n3883 ) | ( (~ preset)  &  n_n3883  &  (~ nrq1_3) ) ;
 assign wire1341 = ( (~ preset)  &  pdn  &  n_n3331 ) | ( (~ preset)  &  n_n3331  &  (~ nrq1_3) ) ;
 assign wire1347 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4330 ) | ( (~ preset)  &  ndn3_6  &  n_n4330 ) ;
 assign wire1351 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4159 ) | ( (~ preset)  &  ndn3_6  &  n_n4159 ) ;
 assign wire1355 = ( (~ preset)  &  pdn  &  n_n4309 ) | ( (~ preset)  &  n_n4309  &  (~ nrq1_3) ) ;
 assign wire1357 = ( (~ preset)  &  pdn  &  n_n3722 ) | ( (~ preset)  &  n_n3722  &  (~ nrq1_3) ) ;
 assign wire1360 = ( (~ preset)  &  pdn  &  n_n3823 ) | ( (~ preset)  &  n_n3823  &  (~ nrq1_3) ) ;
 assign wire1362 = ( n_n3934  &  wire1363 ) | ( (~ preset)  &  n_n3934  &  (~ n_n4126) ) ;
 assign wire1363 = ( (~ n_n3976)  &  wire916 ) ;
 assign wire1365 = ( n_n4316  &  n_n3901  &  wire916  &  n_n3900 ) | ( (~ n_n4316)  &  (~ n_n3901)  &  wire916  &  n_n3900 ) | ( (~ n_n4316)  &  n_n3901  &  wire916  &  (~ n_n3900) ) | ( n_n4316  &  (~ n_n3901)  &  wire916  &  (~ n_n3900) ) ;
 assign wire1375 = ( (~ preset)  &  pdn  &  n_n3385 ) | ( (~ preset)  &  n_n3385  &  (~ nrq1_3) ) ;
 assign wire1378 = ( (~ preset)  &  pdn  &  n_n3202 ) | ( (~ preset)  &  n_n3202  &  (~ nrq1_3) ) ;
 assign wire1381 = ( (~ preset)  &  pdn  &  n_n3055 ) | ( (~ preset)  &  n_n3055  &  (~ nrq1_3) ) ;
 assign wire1385 = ( (~ preset)  &  pdn  &  n_n3463 ) | ( (~ preset)  &  n_n3463  &  (~ nrq1_3) ) ;
 assign wire1387 = ( (~ preset)  &  (~ ndn3_6)  &  n_n3533 ) | ( (~ preset)  &  ndn3_7  &  n_n3533 ) ;
 assign wire1391 = ( (~ preset)  &  n_n4258  &  n_n3832  &  wire6255 ) ;
 assign wire1392 = ( n_n3818  &  (~ n_n3832)  &  wire6257 ) | ( n_n3818  &  (~ wire6255)  &  wire6257 ) ;
 assign wire1393 = ( (~ n_n3818)  &  wire896  &  n_n4256  &  n_n3595 ) | ( n_n3818  &  wire896  &  (~ n_n4256)  &  n_n3595 ) | ( n_n3818  &  wire896  &  n_n4256  &  (~ n_n3595) ) | ( (~ n_n3818)  &  wire896  &  (~ n_n4256)  &  (~ n_n3595) ) ;
 assign wire1400 = ( (~ preset)  &  pdn  &  n_n4390 ) | ( (~ preset)  &  n_n4390  &  (~ nrq1_3) ) ;
 assign wire1402 = ( n_n4229  &  wire916  &  wire1051 ) | ( (~ n_n4229)  &  wire916  &  (~ wire1051) ) ;
 assign wire1412 = ( (~ preset)  &  pdn  &  n_n4136 ) | ( (~ preset)  &  n_n4136  &  (~ nrq1_3) ) ;
 assign wire1414 = ( (~ preset)  &  pdn  &  n_n4192 ) | ( (~ preset)  &  n_n4192  &  (~ nrq1_3) ) ;
 assign wire1416 = ( (~ preset)  &  pdn  &  n_n3126 ) | ( (~ preset)  &  n_n3126  &  (~ nrq1_3) ) ;
 assign wire1425 = ( (~ preset)  &  pdn  &  n_n3089 ) | ( (~ preset)  &  n_n3089  &  (~ nrq1_3) ) ;
 assign wire1427 = ( (~ preset)  &  pdn  &  n_n3713 ) | ( (~ preset)  &  n_n3713  &  (~ nrq1_3) ) ;
 assign wire1429 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3578 ) | ( (~ preset)  &  n_n3578  &  ndn3_9 ) ;
 assign wire1433 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3624 ) | ( (~ preset)  &  n_n3624  &  ndn3_9 ) ;
 assign wire1437 = ( (~ preset)  &  pdn  &  n_n3370 ) | ( (~ preset)  &  n_n3370  &  (~ nrq1_3) ) ;
 assign wire1447 = ( (~ preset)  &  pdn  &  n_n3213 ) | ( (~ preset)  &  n_n3213  &  (~ nrq1_3) ) ;
 assign wire1449 = ( (~ preset)  &  n_n3657  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n3657  &  ngfdn_3 ) ;
 assign wire1451 = ( (~ preset)  &  (~ ndn3_7)  &  n_n3743 ) | ( (~ preset)  &  ndn3_8  &  n_n3743 ) ;
 assign wire1455 = ( (~ preset)  &  pdn  &  n_n3223 ) | ( (~ preset)  &  n_n3223  &  (~ nrq1_3) ) ;
 assign wire1463 = ( (~ preset)  &  pdn  &  n_n4236 ) | ( (~ preset)  &  n_n4236  &  (~ nrq1_3) ) ;
 assign wire1465 = ( (~ preset)  &  pdn  &  n_n4372 ) | ( (~ preset)  &  n_n4372  &  (~ nrq1_3) ) ;
 assign wire1468 = ( (~ preset)  &  pdn  &  n_n3136 ) | ( (~ preset)  &  n_n3136  &  (~ nrq1_3) ) ;
 assign wire1470 = ( (~ preset)  &  (~ n_n3954)  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1472 = ( n_n4349  &  n_n3656 ) | ( n_n4349  &  wire2011 ) ;
 assign wire1477 = ( (~ n_n4056)  &  wire6355 ) | ( n_n4098  &  wire6355 ) | ( (~ wire6349)  &  wire6355 ) ;
 assign wire1482 = ( (~ preset)  &  n_n3259  &  wire1155 ) ;
 assign wire1486 = ( (~ preset)  &  n_n3085  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n3085  &  ngfdn_3 ) ;
 assign wire1487 = ( n_n3810  &  wire1110  &  wire2049 ) | ( n_n3810  &  wire1110  &  wire2050 ) | ( n_n3810  &  (~ wire1110)  &  (~ wire2049)  &  (~ wire2050) ) ;
 assign wire1488 = ( (~ preset)  &  (~ ndn3_7)  &  n_n3946 ) | ( (~ preset)  &  ndn3_8  &  n_n3946 ) ;
 assign wire1492 = ( n_n3709  &  (~ wire6290) ) | ( n_n3709  &  wire1137  &  wire1136 ) ;
 assign wire1494 = ( (~ preset)  &  pdn  &  n_n3777 ) | ( (~ preset)  &  n_n3777  &  (~ nrq1_3) ) ;
 assign wire1497 = ( (~ preset)  &  pdn  &  n_n3073 ) | ( (~ preset)  &  n_n3073  &  (~ nrq1_3) ) ;
 assign wire1500 = ( (~ n_n4012)  &  wire896  &  wire1012  &  wire6330 ) ;
 assign wire1504 = ( (~ preset)  &  pdn  &  n_n3436 ) | ( (~ preset)  &  n_n3436  &  (~ nrq1_3) ) ;
 assign wire1508 = ( (~ preset)  &  ndn3_15  &  n_n4351 ) | ( (~ preset)  &  n_n4351  &  (~ ngfdn_3) ) ;
 assign wire1509 = ( wire1002  &  wire1110  &  wire2049 ) | ( wire1002  &  wire1110  &  wire2050 ) | ( wire1002  &  (~ wire1110)  &  (~ wire2049)  &  (~ wire2050) ) ;
 assign wire1510 = ( (~ preset)  &  pdn  &  n_n3287 ) | ( (~ preset)  &  n_n3287  &  (~ nrq1_3) ) ;
 assign wire1513 = ( (~ preset)  &  pdn  &  n_n3679 ) | ( (~ preset)  &  n_n3679  &  (~ nrq1_3) ) ;
 assign wire1514 = ( (~ preset)  &  pdn  &  n_n4065 ) | ( (~ preset)  &  n_n4065  &  (~ nrq1_3) ) ;
 assign wire1518 = ( (~ preset)  &  pdn  &  n_n3138 ) | ( (~ preset)  &  n_n3138  &  (~ nrq1_3) ) ;
 assign wire1520 = ( (~ preset)  &  pdn  &  n_n3631 ) | ( (~ preset)  &  n_n3631  &  (~ nrq1_3) ) ;
 assign wire1524 = ( (~ preset)  &  pdn  &  n_n3020 ) | ( (~ preset)  &  n_n3020  &  (~ nrq1_3) ) ;
 assign wire1527 = ( (~ preset)  &  pdn  &  n_n3057 ) | ( (~ preset)  &  n_n3057  &  (~ nrq1_3) ) ;
 assign wire1529 = ( (~ preset)  &  pdn  &  n_n3404 ) | ( (~ preset)  &  n_n3404  &  (~ nrq1_3) ) ;
 assign wire1534 = ( (~ preset)  &  pdn  &  n_n3069 ) | ( (~ preset)  &  n_n3069  &  (~ nrq1_3) ) ;
 assign wire1538 = ( n_n3483  &  wire982 ) | ( n_n3483  &  wire1539 ) | ( n_n3483  &  wire1724 ) ;
 assign wire1539 = ( (~ n_n4334)  &  wire896 ) ;
 assign wire1541 = ( (~ preset)  &  (~ ndn3_7)  &  n_n4362 ) | ( (~ preset)  &  ndn3_8  &  n_n4362 ) ;
 assign wire1547 = ( (~ preset)  &  (~ ndn3_6)  &  n_n4201 ) | ( (~ preset)  &  ndn3_7  &  n_n4201 ) ;
 assign wire1551 = ( (~ preset)  &  ndn3_10  &  n_n4229 ) | ( (~ preset)  &  n_n4229  &  (~ nen3_10) ) ;
 assign wire1552 = ( wire1004  &  wire1110  &  wire2049 ) | ( wire1004  &  wire1110  &  wire2050 ) | ( wire1004  &  (~ wire1110)  &  (~ wire2049)  &  (~ wire2050) ) ;
 assign wire1557 = ( (~ preset)  &  pdn  &  n_n3408 ) | ( (~ preset)  &  n_n3408  &  (~ nrq1_3) ) ;
 assign wire1561 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3451 ) | ( (~ preset)  &  ndn3_5  &  n_n3451 ) ;
 assign wire1565 = ( n_n4057  &  (~ n_n4056) ) | ( n_n4057  &  n_n4098 ) | ( n_n4057  &  (~ wire6349) ) ;
 assign wire1574 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3854 ) | ( (~ preset)  &  ndn3_5  &  n_n3854 ) ;
 assign wire1580 = ( n_n4296  &  wire6342 ) | ( n_n3832  &  wire6255  &  wire6342 ) ;
 assign wire1582 = ( (~ n_n3766)  &  wire896 ) ;
 assign wire1584 = ( (~ n_n4227)  &  wire896 ) ;
 assign wire1586 = ( (~ n_n3724)  &  wire896 ) ;
 assign wire1588 = ( (~ n_n3814)  &  wire896 ) ;
 assign wire1594 = ( (~ preset)  &  (~ ndn3_6)  &  n_n3922 ) | ( (~ preset)  &  ndn3_7  &  n_n3922 ) ;
 assign wire1598 = ( (~ preset)  &  (~ ndn3_6)  &  n_n3968 ) | ( (~ preset)  &  ndn3_7  &  n_n3968 ) ;
 assign wire1602 = ( (~ preset)  &  pdn  &  n_n3237 ) | ( (~ preset)  &  n_n3237  &  (~ nrq1_3) ) ;
 assign wire1604 = ( (~ preset)  &  pdn  &  n_n3952 ) | ( (~ preset)  &  n_n3952  &  (~ nrq1_3) ) ;
 assign wire1612 = ( (~ preset)  &  n_n4122  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n4122  &  ngfdn_3 ) ;
 assign wire1613 = ( n_n3810  &  wire1094  &  wire1898 ) | ( n_n3810  &  wire1094  &  wire1899 ) | ( n_n3810  &  (~ wire1094)  &  (~ wire1898)  &  (~ wire1899) ) ;
 assign wire1614 = ( (~ preset)  &  ndn3_10  &  n_n3898 ) | ( (~ preset)  &  n_n3898  &  (~ nen3_10) ) ;
 assign wire1621 = ( (~ preset)  &  n_n4099  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1623 = ( n_n4337  &  n_n3656 ) | ( n_n4337  &  wire2011 ) ;
 assign wire1630 = ( (~ preset)  &  n_n4052  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1632 = ( n_n4052  &  n_n3865  &  n_n4305 ) | ( n_n4052  &  wire984  &  n_n4305 ) | ( (~ n_n4052)  &  (~ n_n3865)  &  (~ wire984)  &  n_n4305 ) ;
 assign wire1633 = ( n_n4071  &  n_n3656 ) | ( n_n4071  &  wire2011 ) ;
 assign wire1638 = ( (~ preset)  &  pdn  &  n_n3985 ) | ( (~ preset)  &  n_n3985  &  (~ nrq1_3) ) ;
 assign wire1640 = ( (~ preset)  &  pdn  &  n_n3091 ) | ( (~ preset)  &  n_n3091  &  (~ nrq1_3) ) ;
 assign wire1642 = ( (~ preset)  &  pdn  &  n_n4003 ) | ( (~ preset)  &  n_n4003  &  (~ nrq1_3) ) ;
 assign wire1647 = ( (~ preset)  &  ndn3_10  &  n_n4145 ) | ( (~ preset)  &  n_n4145  &  (~ nen3_10) ) ;
 assign wire1648 = ( wire1004  &  wire1094  &  wire1898 ) | ( wire1004  &  wire1094  &  wire1899 ) | ( wire1004  &  (~ wire1094)  &  (~ wire1898)  &  (~ wire1899) ) ;
 assign wire1655 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3978 ) | ( (~ preset)  &  ndn3_5  &  n_n3978 ) ;
 assign wire1659 = ( n_n3916  &  wire916  &  wire1038 ) | ( (~ n_n3916)  &  wire916  &  (~ wire1038) ) ;
 assign wire1671 = ( (~ preset)  &  pdn  &  n_n3183 ) | ( (~ preset)  &  n_n3183  &  (~ nrq1_3) ) ;
 assign wire1673 = ( (~ preset)  &  ndn3_15  &  n_n4288 ) | ( (~ preset)  &  n_n4288  &  (~ ngfdn_3) ) ;
 assign wire1679 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4270 ) | ( (~ preset)  &  ndn3_6  &  n_n4270 ) ;
 assign wire1683 = ( (~ preset)  &  pdn  &  n_n3449 ) | ( (~ preset)  &  n_n3449  &  (~ nrq1_3) ) ;
 assign wire1686 = ( (~ preset)  &  pdn  &  n_n3971 ) | ( (~ preset)  &  n_n3971  &  (~ nrq1_3) ) ;
 assign wire1687 = ( (~ preset)  &  pdn  &  n_n3429 ) | ( (~ preset)  &  n_n3429  &  (~ nrq1_3) ) ;
 assign wire1689 = ( (~ preset)  &  pdn  &  n_n3319 ) | ( (~ preset)  &  n_n3319  &  (~ nrq1_3) ) ;
 assign wire1693 = ( (~ preset)  &  pdn  &  n_n3506 ) | ( (~ preset)  &  n_n3506  &  (~ nrq1_3) ) ;
 assign wire1699 = ( (~ preset)  &  ndn3_15  &  n_n3458 ) | ( (~ preset)  &  n_n3458  &  (~ ngfdn_3) ) ;
 assign wire1707 = ( (~ preset)  &  ndn3_15  &  n_n4233 ) | ( (~ preset)  &  n_n4233  &  (~ ngfdn_3) ) ;
 assign wire1708 = ( wire1002  &  (~ n_n3324)  &  n_n3243  &  wire914 ) | ( wire1002  &  n_n3324  &  (~ n_n3243)  &  wire914 ) | ( wire1002  &  n_n3324  &  n_n3243  &  (~ wire914) ) | ( wire1002  &  (~ n_n3324)  &  (~ n_n3243)  &  (~ wire914) ) ;
 assign wire1711 = ( (~ preset)  &  pdn  &  n_n3155 ) | ( (~ preset)  &  n_n3155  &  (~ nrq1_3) ) ;
 assign wire1716 = ( (~ preset)  &  n_n3955  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire1719 = ( n_n4201  &  n_n3656 ) | ( n_n4201  &  wire2011 ) ;
 assign wire1724 = ( (~ n_n4012)  &  wire896 ) ;
 assign wire1726 = ( (~ n_n4275)  &  wire896 ) | ( (~ n_n3766)  &  wire896 ) | ( wire896  &  (~ wire1012) ) ;
 assign wire1728 = ( (~ preset)  &  n_n4294  &  wire1155 ) ;
 assign wire1736 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4251 ) | ( (~ preset)  &  ndn3_6  &  n_n4251 ) ;
 assign wire1740 = ( (~ preset)  &  pdn  &  n_n3736 ) | ( (~ preset)  &  n_n3736  &  (~ nrq1_3) ) ;
 assign wire1742 = ( (~ preset)  &  pdn  &  n_n3896 ) | ( (~ preset)  &  n_n3896  &  (~ nrq1_3) ) ;
 assign wire1745 = ( (~ preset)  &  pdn  &  n_n4279 ) | ( (~ preset)  &  n_n4279  &  (~ nrq1_3) ) ;
 assign wire1752 = ( (~ preset)  &  n_n4362  &  n_n3832  &  wire6255 ) ;
 assign wire1753 = ( n_n3988  &  (~ n_n3832)  &  wire6257 ) | ( n_n3988  &  (~ wire6255)  &  wire6257 ) ;
 assign wire1754 = ( (~ n_n3988)  &  wire896  &  n_n3745  &  n_n3622 ) | ( n_n3988  &  wire896  &  (~ n_n3745)  &  n_n3622 ) | ( n_n3988  &  wire896  &  n_n3745  &  (~ n_n3622) ) | ( (~ n_n3988)  &  wire896  &  (~ n_n3745)  &  (~ n_n3622) ) ;
 assign wire1755 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3328 ) | ( (~ preset)  &  ndn3_5  &  n_n3328 ) ;
 assign wire1767 = ( (~ preset)  &  pdn  &  n_n3761 ) | ( (~ preset)  &  n_n3761  &  (~ nrq1_3) ) ;
 assign wire1771 = ( (~ preset)  &  n_n3946  &  n_n3832  &  wire6255 ) ;
 assign wire1772 = ( n_n3995  &  (~ n_n3832)  &  wire6257 ) | ( n_n3995  &  (~ wire6255)  &  wire6257 ) ;
 assign wire1773 = ( (~ n_n3995)  &  wire896  &  n_n4116  &  n_n3994 ) | ( n_n3995  &  wire896  &  (~ n_n4116)  &  n_n3994 ) | ( n_n3995  &  wire896  &  n_n4116  &  (~ n_n3994) ) | ( (~ n_n3995)  &  wire896  &  (~ n_n4116)  &  (~ n_n3994) ) ;
 assign wire1774 = ( (~ preset)  &  pdn  &  n_n3128 ) | ( (~ preset)  &  n_n3128  &  (~ nrq1_3) ) ;
 assign wire1776 = ( (~ preset)  &  n_n3919  &  wire1155 ) ;
 assign wire1780 = ( (~ preset)  &  n_n3886  &  wire1155 ) ;
 assign wire1784 = ( (~ preset)  &  pdn  &  n_n3048 ) | ( (~ preset)  &  n_n3048  &  (~ nrq1_3) ) ;
 assign wire1786 = ( (~ preset)  &  pdn  &  n_n3061 ) | ( (~ preset)  &  n_n3061  &  (~ nrq1_3) ) ;
 assign wire1788 = ( (~ preset)  &  pdn  &  n_n3316 ) | ( (~ preset)  &  n_n3316  &  (~ nrq1_3) ) ;
 assign wire1792 = ( (~ preset)  &  pdn  &  n_n3906 ) | ( (~ preset)  &  n_n3906  &  (~ nrq1_3) ) ;
 assign wire1795 = ( (~ preset)  &  pdn  &  n_n3583 ) | ( (~ preset)  &  n_n3583  &  (~ nrq1_3) ) ;
 assign wire1800 = ( (~ preset)  &  pdn  &  n_n3358 ) | ( (~ preset)  &  n_n3358  &  (~ nrq1_3) ) ;
 assign wire1806 = ( (~ preset)  &  pdn  &  n_n4243 ) | ( (~ preset)  &  n_n4243  &  (~ nrq1_3) ) ;
 assign wire1812 = ( (~ preset)  &  (~ ndn3_6)  &  n_n4337 ) | ( (~ preset)  &  n_n4337  &  ndn3_7 ) ;
 assign wire1825 = ( (~ preset)  &  pdn  &  n_n3207 ) | ( (~ preset)  &  n_n3207  &  (~ nrq1_3) ) ;
 assign wire1830 = ( (~ preset)  &  pdn  &  n_n3465 ) | ( (~ preset)  &  n_n3465  &  (~ nrq1_3) ) ;
 assign wire1833 = ( pdn  &  ndn1_34  &  wire6325 ) | ( (~ pdn)  &  (~ nrq1_3)  &  wire6325 ) | ( ndn1_34  &  (~ nrq1_3)  &  wire6325 ) ;
 assign wire1837 = ( (~ preset)  &  n_n3892  &  (~ ndn3_6) ) | ( (~ preset)  &  n_n3892  &  ndn3_7 ) ;
 assign wire1843 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4383 ) | ( (~ preset)  &  n_n4383  &  ndn3_6 ) ;
 assign wire1847 = ( (~ preset)  &  pdn  &  n_n4286 ) | ( (~ preset)  &  n_n4286  &  (~ nrq1_3) ) ;
 assign wire1849 = ( (~ preset)  &  pdn  &  n_n4189 ) | ( (~ preset)  &  n_n4189  &  (~ nrq1_3) ) ;
 assign wire1853 = ( (~ preset)  &  pdn  &  n_n3576 ) | ( (~ preset)  &  n_n3576  &  (~ nrq1_3) ) ;
 assign wire1859 = ( (~ preset)  &  pdn  &  n_n4172 ) | ( (~ preset)  &  n_n4172  &  (~ nrq1_3) ) ;
 assign wire1868 = ( (~ preset)  &  pdn  &  n_n3111 ) | ( (~ preset)  &  n_n3111  &  (~ nrq1_3) ) ;
 assign wire1870 = ( (~ preset)  &  n_n3035  &  (~ ndn3_8) ) | ( (~ preset)  &  n_n3035  &  ndn3_9 ) ;
 assign wire1874 = ( (~ preset)  &  pdn  &  n_n3627 ) | ( (~ preset)  &  n_n3627  &  (~ nrq1_3) ) ;
 assign wire1876 = ( (~ preset)  &  pdn  &  n_n3044 ) | ( (~ preset)  &  n_n3044  &  (~ nrq1_3) ) ;
 assign wire1881 = ( (~ preset)  &  pdn  &  n_n3376 ) | ( (~ preset)  &  n_n3376  &  (~ nrq1_3) ) ;
 assign wire1882 = ( (~ preset)  &  pdn  &  n_n3118 ) | ( (~ preset)  &  n_n3118  &  (~ nrq1_3) ) ;
 assign wire1884 = ( (~ preset)  &  n_n3242  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n3242  &  ngfdn_3 ) ;
 assign wire1885 = ( n_n3810  &  (~ n_n3324)  &  n_n3243  &  wire914 ) | ( n_n3810  &  n_n3324  &  (~ n_n3243)  &  wire914 ) | ( n_n3810  &  n_n3324  &  n_n3243  &  (~ wire914) ) | ( n_n3810  &  (~ n_n3324)  &  (~ n_n3243)  &  (~ wire914) ) ;
 assign wire1892 = ( (~ ndn3_15)  &  n_n3556  &  n_n4122  &  ngfdn_3 ) ;
 assign wire1893 = ( (~ ndn3_10)  &  n_n3919  &  nen3_10 ) ;
 assign wire1894 = ( n_n4145  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire1896 = ( (~ ndn3_10)  &  nen3_10  &  n_n4062 ) ;
 assign wire1898 = ( n_n4345  &  n_n4019  &  wire1104 ) | ( n_n4345  &  n_n3884  &  wire1104 ) | ( n_n4019  &  n_n3884  &  wire1104 ) ;
 assign wire1899 = ( n_n3334  &  wire1903 ) | ( n_n3334  &  wire1904 ) | ( n_n3334  &  wire1905 ) ;
 assign wire1901 = ( (~ ndn3_10)  &  n_n3854  &  nen3_10 ) ;
 assign wire1903 = ( (~ ndn3_15)  &  n_n3035  &  n_n4157  &  ngfdn_3 ) ;
 assign wire1904 = ( n_n3511  &  (~ ndn3_10)  &  nen3_10 ) ;
 assign wire1905 = ( n_n3898  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire1908 = ( (~ ndn3_15)  &  n_n3242  &  n_n3170  &  ngfdn_3 ) ;
 assign wire1909 = ( (~ ndn3_10)  &  nen3_10  &  n_n3259 ) ;
 assign wire1910 = ( nrq3_11  &  (~ ngfdn_3)  &  n_n3841 ) ;
 assign wire1912 = ( (~ ndn3_10)  &  n_n3451  &  nen3_10 ) ;
 assign wire1914 = ( (~ preset)  &  pdn  &  n_n3113 ) | ( (~ preset)  &  n_n3113  &  (~ nrq1_3) ) ;
 assign wire1919 = ( (~ preset)  &  pdn  &  n_n3173 ) | ( (~ preset)  &  n_n3173  &  (~ nrq1_3) ) ;
 assign wire1921 = ( (~ preset)  &  pdn  &  n_n3221 ) | ( (~ preset)  &  n_n3221  &  (~ nrq1_3) ) ;
 assign wire1925 = ( (~ preset)  &  n_n3876  &  n_n3832  &  wire6255 ) ;
 assign wire1926 = ( n_n4040  &  (~ n_n3832)  &  wire6257 ) | ( n_n4040  &  (~ wire6255)  &  wire6257 ) ;
 assign wire1927 = ( (~ n_n4040)  &  wire896  &  n_n4069  &  n_n4039 ) | ( n_n4040  &  wire896  &  (~ n_n4069)  &  n_n4039 ) | ( n_n4040  &  wire896  &  n_n4069  &  (~ n_n4039) ) | ( (~ n_n4040)  &  wire896  &  (~ n_n4069)  &  (~ n_n4039) ) ;
 assign wire1928 = ( (~ preset)  &  n_n3556  &  (~ ndn3_8) ) | ( (~ preset)  &  n_n3556  &  ndn3_9 ) ;
 assign wire1932 = ( (~ preset)  &  pdn  &  n_n3733 ) | ( (~ preset)  &  n_n3733  &  (~ nrq1_3) ) ;
 assign wire1940 = ( (~ preset)  &  pdn  &  n_n3231 ) | ( (~ preset)  &  n_n3231  &  (~ nrq1_3) ) ;
 assign wire1944 = ( (~ preset)  &  pdn  &  n_n3313 ) | ( (~ preset)  &  n_n3313  &  (~ nrq1_3) ) ;
 assign wire1946 = ( (~ preset)  &  pdn  &  n_n3079 ) | ( (~ preset)  &  n_n3079  &  (~ nrq1_3) ) ;
 assign wire1949 = ( (~ preset)  &  n_n3688  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n3688  &  ngfdn_3 ) ;
 assign wire1953 = ( (~ preset)  &  pdn  &  n_n3344 ) | ( (~ preset)  &  n_n3344  &  (~ nrq1_3) ) ;
 assign wire1957 = ( (~ preset)  &  n_n4071  &  (~ ndn3_6) ) | ( (~ preset)  &  n_n4071  &  ndn3_7 ) ;
 assign wire1961 = ( (~ preset)  &  pdn  &  n_n3012 ) | ( (~ preset)  &  n_n3012  &  (~ nrq1_3) ) ;
 assign wire1963 = ( (~ preset)  &  n_n4222  &  ndn3_10 ) | ( (~ preset)  &  n_n4222  &  (~ nen3_10) ) ;
 assign wire1965 = ( (~ preset)  &  (~ ndn3_5)  &  n_n4160 ) | ( (~ preset)  &  n_n4160  &  ndn3_6 ) ;
 assign wire1969 = ( (~ preset)  &  pdn  &  n_n3517 ) | ( (~ preset)  &  n_n3517  &  (~ nrq1_3) ) ;
 assign wire1971 = ( n_n3707  &  (~ n_n3709) ) | ( n_n3707  &  n_n135 ) | ( n_n3707  &  (~ wire6290) ) ;
 assign wire1976 = ( (~ preset)  &  (~ ndn3_4)  &  n_n3281 ) | ( (~ preset)  &  ndn3_5  &  n_n3281 ) ;
 assign wire1980 = ( (~ preset)  &  pdn  &  n_n3764 ) | ( (~ preset)  &  n_n3764  &  (~ nrq1_3) ) ;
 assign wire1984 = ( (~ preset)  &  pdn  &  n_n3549 ) | ( (~ preset)  &  n_n3549  &  (~ nrq1_3) ) ;
 assign wire1986 = ( (~ preset)  &  n_n3876  &  (~ ndn3_7) ) | ( (~ preset)  &  n_n3876  &  ndn3_8 ) ;
 assign wire1990 = ( (~ preset)  &  pdn  &  n_n3729 ) | ( (~ preset)  &  n_n3729  &  (~ nrq1_3) ) ;
 assign wire1992 = ( (~ preset)  &  pdn  &  n_n3525 ) | ( (~ preset)  &  n_n3525  &  (~ nrq1_3) ) ;
 assign wire1996 = ( (~ preset)  &  n_n3916  &  ndn3_10 ) | ( (~ preset)  &  n_n3916  &  (~ nen3_10) ) ;
 assign wire1998 = ( (~ preset)  &  ndn3_15  &  n_n3495 ) | ( (~ preset)  &  n_n3495  &  (~ ngfdn_3) ) ;
 assign wire2000 = ( (~ preset)  &  n_n4211  &  (~ ndn3_8) ) | ( (~ preset)  &  n_n4211  &  ndn3_9 ) ;
 assign wire2005 = ( (~ preset)  &  pdn  &  n_n3670 ) | ( (~ preset)  &  n_n3670  &  (~ nrq1_3) ) ;
 assign wire2007 = ( (~ preset)  &  n_n4381  &  (~ n_n4126)  &  (~ n_n3500) ) ;
 assign wire2009 = ( n_n3892  &  n_n3656 ) | ( n_n3892  &  wire2011 ) ;
 assign wire2011 = ( (~ n_n3493)  &  (~ n_n4045)  &  (~ n_n4367) ) | ( (~ n_n3493)  &  (~ n_n4367)  &  wire6299 ) ;
 assign wire2023 = ( (~ preset)  &  n_n3858  &  wire1155 ) ;
 assign wire2027 = ( (~ preset)  &  pdn  &  n_n3270 ) | ( (~ preset)  &  n_n3270  &  (~ nrq1_3) ) ;
 assign wire2029 = ( (~ preset)  &  n_n4074  &  (~ nrq3_11) ) | ( (~ preset)  &  n_n4074  &  ngfdn_3 ) ;
 assign wire2035 = ( (~ ndn3_15)  &  n_n4074  &  n_n3578  &  ngfdn_3 ) ;
 assign wire2036 = ( (~ ndn3_10)  &  n_n3886  &  nen3_10 ) ;
 assign wire2037 = ( n_n3916  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire2039 = ( (~ ndn3_10)  &  nen3_10  &  n_n4021 ) ;
 assign wire2044 = ( n_n3281  &  (~ ndn3_10)  &  nen3_10 ) ;
 assign wire2045 = ( n_n4229  &  nrq3_11  &  (~ ngfdn_3)  &  wire1079 ) | ( (~ n_n4229)  &  nrq3_11  &  (~ ngfdn_3)  &  (~ wire1079) ) ;
 assign wire2046 = ( (~ ndn3_15)  &  n_n3085  &  n_n3250  &  ngfdn_3 ) ;
 assign wire2047 = ( (~ ndn3_10)  &  n_n4294  &  nen3_10 ) ;
 assign wire2048 = ( n_n4229  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire2049 = ( n_n3363  &  n_n3362  &  wire1088 ) | ( n_n3363  &  wire1088  &  (~ wire941) ) | ( n_n3362  &  wire1088  &  (~ wire941) ) ;
 assign wire2050 = ( n_n3981  &  wire2174 ) | ( n_n3981  &  wire6281 ) ;
 assign wire2051 = ( (~ preset)  &  pdn  &  n_n3133 ) | ( (~ preset)  &  n_n3133  &  (~ nrq1_3) ) ;
 assign wire2060 = ( (~ n_n3786)  &  (~ n_n3785) ) | ( (~ n_n3786)  &  wire6287 ) ;
 assign wire2061 = ( (~ n_n4145)  &  n_n4080  &  wire1075  &  n_n4078 ) | ( n_n4145  &  n_n4080  &  (~ wire1075)  &  n_n4078 ) | ( (~ n_n4145)  &  (~ n_n4080)  &  wire1075  &  (~ n_n4078) ) | ( n_n4145  &  (~ n_n4080)  &  (~ wire1075)  &  (~ n_n4078) ) ;
 assign wire2122 = ( (~ preset)  &  n_n4224  &  (~ ndn3_5) ) | ( (~ preset)  &  n_n4224  &  ndn3_6 ) ;
 assign wire2126 = ( (~ preset)  &  n_n4392  &  ndn3_15 ) | ( (~ preset)  &  n_n4392  &  (~ ngfdn_3) ) ;
 assign wire2141 = ( (~ preset)  &  n_n3511  &  wire1155 ) ;
 assign wire2153 = ( (~ preset)  &  pdn  &  n_n3780 ) | ( (~ preset)  &  n_n3780  &  (~ nrq1_3) ) ;
 assign wire2162 = ( (~ preset)  &  n_n4349  &  (~ ndn3_6) ) | ( (~ preset)  &  n_n4349  &  ndn3_7 ) ;
 assign wire2166 = ( (~ preset)  &  n_n4316  &  ndn3_10 ) | ( (~ preset)  &  n_n4316  &  (~ nen3_10) ) ;
 assign wire2173 = ( (~ ndn3_10)  &  n_n3978  &  nen3_10 ) ;
 assign wire2174 = ( n_n4316  &  nrq3_12  &  n_n4315  &  n_n4155 ) | ( (~ n_n4316)  &  nrq3_12  &  (~ n_n4315)  &  n_n4155 ) | ( (~ n_n4316)  &  nrq3_12  &  n_n4315  &  (~ n_n4155) ) | ( n_n4316  &  nrq3_12  &  (~ n_n4315)  &  (~ n_n4155) ) ;
 assign wire2175 = ( (~ ndn3_15)  &  n_n4211  &  n_n3657  &  ngfdn_3 ) ;
 assign wire2176 = ( n_n3858  &  (~ ndn3_10)  &  nen3_10 ) ;
 assign wire2177 = ( n_n4316  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire2182 = ( nrq3_11  &  (~ n_n4159)  &  n_n3976  &  (~ ngfdn_3) ) | ( nrq3_11  &  n_n4159  &  (~ n_n3976)  &  (~ ngfdn_3) ) ;
 assign wire2183 = ( (~ ndn3_15)  &  n_n3688  &  n_n3624  &  ngfdn_3 ) ;
 assign wire2184 = ( (~ ndn3_10)  &  nen3_10  &  n_n3878 ) ;
 assign wire2185 = ( nrq3_11  &  n_n3976  &  (~ ngfdn_3) ) ;
 assign wire2187 = ( (~ ndn3_10)  &  n_n3328  &  nen3_10 ) ;
 assign wire2188 = ( nrq3_11  &  (~ ngfdn_3)  &  n_n3741 ) ;
 assign wire2189 = ( n_n3936  &  (~ ndn3_15)  &  ngfdn_3  &  n_n3099 ) ;
 assign wire2190 = ( (~ ndn3_10)  &  nen3_10  &  n_n3208 ) ;
 assign wire2191 = ( n_n4222  &  nrq3_11  &  (~ ngfdn_3) ) ;
 assign wire2192 = ( (~ preset)  &  pdn  &  n_n3793 ) | ( (~ preset)  &  n_n3793  &  (~ nrq1_3) ) ;
 assign wire2195 = ( (~ preset)  &  pdn  &  n_n3497 ) | ( (~ preset)  &  n_n3497  &  (~ nrq1_3) ) ;
 assign wire2198 = ( (~ preset)  &  pdn  &  n_n3098 ) | ( (~ preset)  &  n_n3098  &  (~ nrq1_3) ) ;
 assign wire2202 = ( (~ preset)  &  pdn  &  n_n3687 ) | ( (~ preset)  &  n_n3687  &  (~ nrq1_3) ) ;
 assign wire2224 = ( (~ preset)  &  pdn  &  n_n3225 ) | ( (~ preset)  &  n_n3225  &  (~ nrq1_3) ) ;
 assign wire2226 = ( (~ preset)  &  n_n4258  &  (~ ndn3_7) ) | ( (~ preset)  &  n_n4258  &  ndn3_8 ) ;
 assign wire2240 = ( (~ preset)  &  n_n4360  &  n_n3832  &  wire6255 ) ;
 assign wire2241 = ( n_n3726  &  (~ n_n3832)  &  wire6257 ) | ( n_n3726  &  (~ wire6255)  &  wire6257 ) ;
 assign wire2242 = ( (~ n_n3726)  &  wire896  &  n_n3653  &  n_n3888 ) | ( n_n3726  &  wire896  &  (~ n_n3653)  &  n_n3888 ) | ( n_n3726  &  wire896  &  n_n3653  &  (~ n_n3888) ) | ( (~ n_n3726)  &  wire896  &  (~ n_n3653)  &  (~ n_n3888) ) ;
 assign wire2259 = ( (~ preset)  &  pdn  &  n_n3008 ) | ( (~ preset)  &  n_n3008  &  (~ nrq1_3) ) ;
 assign wire2261 = ( (~ preset)  &  n_n3743  &  n_n3832  &  wire6255 ) ;
 assign wire2262 = ( n_n3574  &  (~ n_n3832)  &  wire6257 ) | ( n_n3574  &  (~ wire6255)  &  wire6257 ) ;
 assign wire2263 = ( (~ n_n3574)  &  wire896  &  n_n3741  &  wire923 ) | ( n_n3574  &  wire896  &  (~ n_n3741)  &  wire923 ) | ( n_n3574  &  wire896  &  n_n3741  &  (~ wire923) ) | ( (~ n_n3574)  &  wire896  &  (~ n_n3741)  &  (~ wire923) ) ;
 assign wire2264 = ( (~ n_n3851)  &  (~ n_n4067)  &  n_n4026 ) | ( (~ n_n4067)  &  (~ n_n4026)  &  (~ n_n3852) ) ;
 assign wire2270 = ( (~ preset)  &  n_n3936  &  (~ ndn3_8) ) | ( (~ preset)  &  n_n3936  &  ndn3_9 ) ;
 assign wire2275 = ( (~ preset)  &  pdn  &  n_n4142 ) | ( (~ preset)  &  n_n4142  &  (~ nrq1_3) ) ;
 assign wire6250 = ( (~ n_n4159)  &  n_n3976  &  (~ n_n3756) ) | ( n_n4159  &  (~ n_n3976)  &  (~ n_n3756) ) ;
 assign wire6251 = ( (~ n_n4182)  &  (~ n_n4330) ) ;
 assign wire6252 = ( n_n3833  &  n_n4067  &  wire894 ) | ( n_n3833  &  wire894  &  (~ n_n3563) ) | ( (~ n_n4067)  &  wire894  &  (~ n_n3563) ) ;
 assign wire6254 = ( nen3_10  &  nsr3_17  &  n_n4093 ) ;
 assign wire6255 = ( wire1015  &  (~ n_n3709) ) ;
 assign wire6257 = ( (~ preset)  &  n_n3198 ) | ( (~ preset)  &  (~ n_n3707) ) | ( (~ preset)  &  (~ n_n3709) ) ;
 assign wire6259 = ( n_n4157  &  n_n3035 ) ;
 assign wire6265 = ( n_n4349 ) | ( n_n4071 ) | ( n_n3892 ) | ( n_n4337 ) ;
 assign wire6266 = ( n_n3968 ) | ( n_n3922 ) | ( n_n4201 ) | ( n_n3533 ) ;
 assign wire6268 = ( n_n4045  &  (~ nsr3_17)  &  nsr3_14 ) ;
 assign wire6270 = ( (~ n_n3557)  &  n_n4057 ) ;
 assign wire6272 = ( n_n3624  &  n_n3688 ) ;
 assign wire6275 = ( wire2187 ) | ( n_n4125  &  n_n4367  &  nrq3_15 ) ;
 assign wire6278 = ( wire2182 ) | ( (~ ndn3_10)  &  nen3_10  &  n_n3931 ) ;
 assign wire6281 = ( wire2173 ) | ( n_n3901  &  n_n4367  &  nrq3_15 ) ;
 assign wire6284 = ( (~ ndn3_4)  &  (~ preset) ) ;
 assign wire6287 = ( (~ n_n4145)  &  wire1075 ) | ( n_n4145  &  (~ wire1075) ) | ( n_n4145  &  (~ n_n4080)  &  wire1075  &  n_n4078 ) | ( (~ n_n4145)  &  (~ n_n4080)  &  (~ wire1075)  &  n_n4078 ) | ( n_n4145  &  n_n4080  &  wire1075  &  (~ n_n4078) ) | ( (~ n_n4145)  &  n_n4080  &  (~ wire1075)  &  (~ n_n4078) ) ;
 assign wire6289 = ( n_n3653 ) | ( wire2061 ) | ( (~ n_n3726)  &  (~ n_n3653)  &  n_n3888 ) | ( n_n3726  &  (~ n_n3653)  &  (~ n_n3888) ) ;
 assign wire6290 = ( n_n4296  &  wire2060 ) | ( n_n4296  &  wire6289 ) ;
 assign wire6291 = ( n_n3578  &  n_n4074 ) ;
 assign wire6295 = ( wire2044 ) | ( n_n3769  &  n_n4367  &  nrq3_15 ) ;
 assign wire6296 = ( wire2039 ) | ( n_n4047  &  n_n4367  &  nrq3_15 ) ;
 assign wire6299 = ( nsr3_14  &  (~ nsr3_17) ) ;
 assign wire6300 = ( n_n4305  &  n_n4357 ) | ( n_n4381  &  wire1008 ) ;
 assign wire6302 = ( n_n3493  &  (~ preset) ) ;
 assign wire6303 = ( n_n3170  &  n_n3242 ) ;
 assign wire6306 = ( n_n3099  &  n_n3936 ) ;
 assign wire6309 = ( (~ n_n3831) ) | ( n_n4026 ) | ( (~ n_n4026)  &  (~ n_n3852) ) ;
 assign wire6310 = ( n_n3657  &  n_n4211 ) ;
 assign wire6312 = ( wire1912 ) | ( n_n4324  &  n_n4367  &  nrq3_15 ) ;
 assign wire6317 = ( wire1901 ) | ( n_n4366  &  n_n4367  &  nrq3_15 ) ;
 assign wire6318 = ( wire1896 ) | ( n_n3475  &  n_n4367  &  nrq3_15 ) ;
 assign wire6321 = ( n_n4122  &  n_n3556 ) ;
 assign wire6322 = ( n_n3250  &  n_n3085 ) ;
 assign wire6324 = ( (~ tin_pready_0_0_)  &  (~ n_n4108)  &  nsr3_3 ) | ( (~ tin_pready_0_0_)  &  (~ n_n3354)  &  nsr3_3 ) | ( n_n4108  &  (~ n_n3354)  &  nsr3_3 ) ;
 assign wire6325 = ( n_n3354  &  (~ preset) ) ;
 assign wire6330 = ( n_n3766  &  n_n4275 ) ;
 assign wire6332 = ( n_n3955  &  wire1008 ) | ( (~ n_n3955)  &  n_n3954  &  n_n4305 ) | ( n_n3955  &  (~ n_n3954)  &  n_n4305 ) ;
 assign wire6333 = ( nlak4_2 ) | ( nlc3_3  &  (~ n_n4263) ) ;
 assign wire6337 = ( wire1632 ) | ( n_n4052  &  wire1008 ) ;
 assign wire6338 = ( n_n4099  &  wire1008 ) | ( n_n4099  &  n_n4305  &  wire1119 ) | ( (~ n_n4099)  &  n_n4305  &  (~ wire1119) ) ;
 assign wire6342 = ( (~ n_n4275)  &  n_n3766  &  wire896  &  wire1012 ) ;
 assign wire6343 = ( (~ n_n3954)  &  (~ n_n3955) ) ;
 assign wire6346 = ( n_n4305  &  (~ n_n4006)  &  (~ n_n3848)  &  wire6343 ) ;
 assign wire6349 = ( (~ n_n3294)  &  (~ n_n4357)  &  wire942  &  wire6346 ) ;
 assign wire6350 = ( preset ) | ( (~ n_n4045) ) | ( (~ n_n4367)  &  wire6299 ) ;
 assign wire6354 = ( n_n3707  &  (~ preset) ) ;
 assign wire6355 = ( n_n4367  &  n_n4057 ) ;
 assign wire6356 = ( (~ nsr3_14) ) | ( nsr3_17 ) ;
 assign wire6357 = ( preset ) | ( (~ n_n4045) ) | ( (~ n_n4367)  &  wire6299 ) ;
 assign wire6358 = ( n_n3954  &  n_n4305 ) | ( (~ n_n3954)  &  wire1008 ) ;
 assign wire6361 = ( (~ preset)  &  n_n4045  &  n_n4367 ) | ( (~ preset)  &  n_n4045  &  (~ wire6299) ) ;
 assign wire6366 = ( n_n4305  &  n_n4006 ) | ( n_n4029  &  wire1008 ) ;
 assign wire6370 = ( n_n3724  &  (~ n_n3766)  &  n_n4227  &  n_n3814 ) ;
 assign wire6374 = ( wire1015  &  n_n3707 ) ;
 assign wire6376 = ( preset ) | ( nak3_17 ) | ( wire1063  &  wire6374 ) ;
 assign wire6379 = ( n_n4305  &  n_n3848 ) | ( n_n3845  &  wire1008 ) ;
 assign wire6380 = ( n_n3865  &  wire1008 ) | ( n_n3865  &  wire984  &  n_n4305 ) | ( (~ n_n3865)  &  (~ wire984)  &  n_n4305 ) ;
 assign wire6385 = ( wire1070  &  wire916 ) ;
 assign wire6386 = ( (~ preset)  &  n_n3709  &  (~ n_n135)  &  wire6290 ) ;
 assign wire6387 = ( n_n3563  &  (~ n_n4067) ) ;
 assign wire6389 = ( n_n4093  &  (~ n_n3788)  &  wire1013  &  (~ wire2264) ) ;


endmodule

