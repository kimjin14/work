module clma (
	pi18, pi106, pi117, pi128, pi139, pi203, pi214, pi225, 
	pi236, pi247, pi258, pi269, pi300, pi311, pi322, pi333, pi344, pi355, 
	pi366, pi377, pi388, pi399, pi17, pi105, pi118, pi127, pi149, pi202, 
	pi215, pi224, pi237, pi246, pi259, pi268, pi312, pi321, pi334, pi343, 
	pi356, pi365, pi378, pi387, pi27, pi108, pi115, pi126, pi159, pi205, 
	pi212, pi223, pi238, pi249, pi256, pi267, pi302, pi320, pi335, pi346, 
	pi353, pi364, pi379, pi397, pi19, pi28, pi107, pi116, pi125, pi169, 
	pi204, pi213, pi222, pi239, pi248, pi257, pi266, pi301, pi310, pi336, 
	pi345, pi354, pi363, pi389, pi398, pi58, pi69, pi135, pi146, pi157, 
	pi168, pi207, pi218, pi229, pi232, pi243, pi254, pi265, pi304, pi315, 
	pi326, pi340, pi351, pi362, pi401, pi412, pi57, pi79, pi109, pi136, 
	pi145, pi158, pi167, pi206, pi219, pi228, pi233, pi242, pi255, pi264, 
	pi303, pi316, pi325, pi330, pi352, pi361, pi400, pi413, pi49, pi67, 
	pi78, pi119, pi137, pi148, pi155, pi166, pi209, pi216, pi227, pi234, 
	pi245, pi252, pi263, pi306, pi313, pi324, pi331, pi342, pi360, pi403, 
	pi410, pi59, pi68, pi77, pi129, pi138, pi147, pi156, pi165, pi208, 
	pi217, pi226, pi235, pi244, pi253, pi262, pi305, pi314, pi323, pi332, 
	pi341, pi350, pi402, pi411, pi87, pi98, pi120, pi131, pi142, pi153, 
	pi164, pi250, pi261, pi88, pi97, pi110, pi132, pi141, pi154, pi163, 
	pi251, pi260, pi89, pi100, pi133, pi144, pi151, pi162, pi230, pi241, 
	pi99, pi134, pi143, pi152, pi161, pi231, pi240, pi102, pi113, pi124, 
	pi160, pi210, pi221, pi101, pi114, pi123, pi150, pi211, pi220, pi104, 
	pi111, pi122, pi140, pi201, pi103, pi112, pi121, pi130, pi200, pi90, 
	pi80, pi190, pclk, pi81, pi92, pi180, pi82, pi91, pi170, pi83, 
	pi94, pi171, pi182, pi193, pi290, pi84, pi93, pi172, pi181, pi194, 
	pi291, pi85, pi96, pi173, pi184, pi191, pi270, pi281, pi86, pi95, 
	pi174, pi183, pi192, pi271, pi280, pi21, pi54, pi65, pi76, pi175, 
	pi186, pi197, pi272, pi283, pi294, pi308, pi319, pi380, pi391, pi405, 
	pi416, pi22, pi53, pi66, pi75, pi176, pi185, pi198, pi273, pi282, 
	pi295, pi307, pi329, pi370, pi392, pi404, pi56, pi63, pi74, pi177, 
	pi188, pi195, pi274, pi285, pi292, pi317, pi328, pi371, pi382, pi407, 
	pi414, pi20, pi55, pi64, pi73, pi178, pi187, pi196, pi275, pi284, 
	pi293, pi309, pi318, pi327, pi372, pi381, pi390, pi406, pi415, pi25, 
	pi50, pi61, pi72, pi179, pi276, pi287, pi298, pi337, pi348, pi359, 
	pi373, pi384, pi395, pi409, pi26, pi62, pi71, pi189, pi277, pi286, 
	pi299, pi338, pi347, pi369, pi374, pi383, pi396, pi408, pi16, pi23, 
	pi52, pi70, pi199, pi278, pi289, pi296, pi339, pi357, pi368, pi375, 
	pi386, pi393, pi15, pi24, pi51, pi60, pi279, pi288, pi297, pi349, 
	pi358, pi367, pi376, pi385, pi394, p__cmx0ad_11, p__cmx0ad_22, p__cmx0ad_33, p__cmx1ad_7, p__cmx0ad_10, 
	p__cmx0ad_23, p__cmx0ad_32, p__cmx1ad_8, p__cmx0ad_24, p__cmx0ad_35, p__cmx1ad_5, p__cmx0ad_25, p__cmx0ad_34, p__cmx1ad_6, p__cmnxcp_0, 
	p__cmx0ad_15, p__cmx1ad_16, p__cmx1ad_27, p__cmxcl_0, p__cmnxcp_1, p__cmx0ad_14, p__cmx1ad_17, p__cmx1ad_26, p__cmxcl_1, p__cmx0ad_13, 
	p__cmx0ad_20, p__cmx0ad_31, p__cmx1ad_9, p__cmx1ad_18, p__cmx1ad_29, p__cmx0ad_12, p__cmx0ad_21, p__cmx0ad_30, p__cmx1ad_19, p__cmx1ad_28, 
	p__cmx0ad_8, p__cmx0ad_9, p__cmx1ad_0, p__cmndst1p0, p__cmx0ad_6, p__cmx0ad_7, p__cmx1ad_3, p__cmndst0p0, p__cmx1ad_4, p__cmx1ad_1, 
	p__cmx1ad_2, p__cmx0ad_0, p__cmx0ad_1, p__cmx0ad_4, p__cmx0ad_5, p__cmxig_0, p__cmx0ad_2, p__cmxig_1, p__cmx0ad_3, p__cmx0ad_19, 
	p__cmx1ad_12, p__cmx1ad_23, p__cmx1ad_34, p__cmxir_0, p__cmx0ad_18, p__cmx1ad_13, p__cmx1ad_22, p__cmx1ad_35, p__cmxir_1, p__cmx0ad_17, 
	p__cmx1ad_14, p__cmx1ad_25, p__cmx1ad_32, p__cmx0ad_16, p__cmx1ad_15, p__cmx1ad_24, p__cmx1ad_33, p__cmx0ad_26, p__cmx1ad_30, p__cmx0ad_27, 
	p__cmx1ad_31, p__cmx0ad_28, p__cmx1ad_10, p__cmx1ad_21, p__cmx0ad_29, p__cmx1ad_11, p__cmx1ad_20);

input pi18;
input pi106;
input pi117;
input pi128;
input pi139;
input pi203;
input pi214;
input pi225;
input pi236;
input pi247;
input pi258;
input pi269;
input pi300;
input pi311;
input pi322;
input pi333;
input pi344;
input pi355;
input pi366;
input pi377;
input pi388;
input pi399;
input pi17;
input pi105;
input pi118;
input pi127;
input pi149;
input pi202;
input pi215;
input pi224;
input pi237;
input pi246;
input pi259;
input pi268;
input pi312;
input pi321;
input pi334;
input pi343;
input pi356;
input pi365;
input pi378;
input pi387;
input pi27;
input pi108;
input pi115;
input pi126;
input pi159;
input pi205;
input pi212;
input pi223;
input pi238;
input pi249;
input pi256;
input pi267;
input pi302;
input pi320;
input pi335;
input pi346;
input pi353;
input pi364;
input pi379;
input pi397;
input pi19;
input pi28;
input pi107;
input pi116;
input pi125;
input pi169;
input pi204;
input pi213;
input pi222;
input pi239;
input pi248;
input pi257;
input pi266;
input pi301;
input pi310;
input pi336;
input pi345;
input pi354;
input pi363;
input pi389;
input pi398;
input pi58;
input pi69;
input pi135;
input pi146;
input pi157;
input pi168;
input pi207;
input pi218;
input pi229;
input pi232;
input pi243;
input pi254;
input pi265;
input pi304;
input pi315;
input pi326;
input pi340;
input pi351;
input pi362;
input pi401;
input pi412;
input pi57;
input pi79;
input pi109;
input pi136;
input pi145;
input pi158;
input pi167;
input pi206;
input pi219;
input pi228;
input pi233;
input pi242;
input pi255;
input pi264;
input pi303;
input pi316;
input pi325;
input pi330;
input pi352;
input pi361;
input pi400;
input pi413;
input pi49;
input pi67;
input pi78;
input pi119;
input pi137;
input pi148;
input pi155;
input pi166;
input pi209;
input pi216;
input pi227;
input pi234;
input pi245;
input pi252;
input pi263;
input pi306;
input pi313;
input pi324;
input pi331;
input pi342;
input pi360;
input pi403;
input pi410;
input pi59;
input pi68;
input pi77;
input pi129;
input pi138;
input pi147;
input pi156;
input pi165;
input pi208;
input pi217;
input pi226;
input pi235;
input pi244;
input pi253;
input pi262;
input pi305;
input pi314;
input pi323;
input pi332;
input pi341;
input pi350;
input pi402;
input pi411;
input pi87;
input pi98;
input pi120;
input pi131;
input pi142;
input pi153;
input pi164;
input pi250;
input pi261;
input pi88;
input pi97;
input pi110;
input pi132;
input pi141;
input pi154;
input pi163;
input pi251;
input pi260;
input pi89;
input pi100;
input pi133;
input pi144;
input pi151;
input pi162;
input pi230;
input pi241;
input pi99;
input pi134;
input pi143;
input pi152;
input pi161;
input pi231;
input pi240;
input pi102;
input pi113;
input pi124;
input pi160;
input pi210;
input pi221;
input pi101;
input pi114;
input pi123;
input pi150;
input pi211;
input pi220;
input pi104;
input pi111;
input pi122;
input pi140;
input pi201;
input pi103;
input pi112;
input pi121;
input pi130;
input pi200;
input pi90;
input pi80;
input pi190;
input pclk;
input pi81;
input pi92;
input pi180;
input pi82;
input pi91;
input pi170;
input pi83;
input pi94;
input pi171;
input pi182;
input pi193;
input pi290;
input pi84;
input pi93;
input pi172;
input pi181;
input pi194;
input pi291;
input pi85;
input pi96;
input pi173;
input pi184;
input pi191;
input pi270;
input pi281;
input pi86;
input pi95;
input pi174;
input pi183;
input pi192;
input pi271;
input pi280;
input pi21;
input pi54;
input pi65;
input pi76;
input pi175;
input pi186;
input pi197;
input pi272;
input pi283;
input pi294;
input pi308;
input pi319;
input pi380;
input pi391;
input pi405;
input pi416;
input pi22;
input pi53;
input pi66;
input pi75;
input pi176;
input pi185;
input pi198;
input pi273;
input pi282;
input pi295;
input pi307;
input pi329;
input pi370;
input pi392;
input pi404;
input pi56;
input pi63;
input pi74;
input pi177;
input pi188;
input pi195;
input pi274;
input pi285;
input pi292;
input pi317;
input pi328;
input pi371;
input pi382;
input pi407;
input pi414;
input pi20;
input pi55;
input pi64;
input pi73;
input pi178;
input pi187;
input pi196;
input pi275;
input pi284;
input pi293;
input pi309;
input pi318;
input pi327;
input pi372;
input pi381;
input pi390;
input pi406;
input pi415;
input pi25;
input pi50;
input pi61;
input pi72;
input pi179;
input pi276;
input pi287;
input pi298;
input pi337;
input pi348;
input pi359;
input pi373;
input pi384;
input pi395;
input pi409;
input pi26;
input pi62;
input pi71;
input pi189;
input pi277;
input pi286;
input pi299;
input pi338;
input pi347;
input pi369;
input pi374;
input pi383;
input pi396;
input pi408;
input pi16;
input pi23;
input pi52;
input pi70;
input pi199;
input pi278;
input pi289;
input pi296;
input pi339;
input pi357;
input pi368;
input pi375;
input pi386;
input pi393;
input pi15;
input pi24;
input pi51;
input pi60;
input pi279;
input pi288;
input pi297;
input pi349;
input pi358;
input pi367;
input pi376;
input pi385;
input pi394;
output p__cmx0ad_11;
output p__cmx0ad_22;
output p__cmx0ad_33;
output p__cmx1ad_7;
output p__cmx0ad_10;
output p__cmx0ad_23;
output p__cmx0ad_32;
output p__cmx1ad_8;
output p__cmx0ad_24;
output p__cmx0ad_35;
output p__cmx1ad_5;
output p__cmx0ad_25;
output p__cmx0ad_34;
output p__cmx1ad_6;
output p__cmnxcp_0;
output p__cmx0ad_15;
output p__cmx1ad_16;
output p__cmx1ad_27;
output p__cmxcl_0;
output p__cmnxcp_1;
output p__cmx0ad_14;
output p__cmx1ad_17;
output p__cmx1ad_26;
output p__cmxcl_1;
output p__cmx0ad_13;
output p__cmx0ad_20;
output p__cmx0ad_31;
output p__cmx1ad_9;
output p__cmx1ad_18;
output p__cmx1ad_29;
output p__cmx0ad_12;
output p__cmx0ad_21;
output p__cmx0ad_30;
output p__cmx1ad_19;
output p__cmx1ad_28;
output p__cmx0ad_8;
output p__cmx0ad_9;
output p__cmx1ad_0;
output p__cmndst1p0;
output p__cmx0ad_6;
output p__cmx0ad_7;
output p__cmx1ad_3;
output p__cmndst0p0;
output p__cmx1ad_4;
output p__cmx1ad_1;
output p__cmx1ad_2;
output p__cmx0ad_0;
output p__cmx0ad_1;
output p__cmx0ad_4;
output p__cmx0ad_5;
output p__cmxig_0;
output p__cmx0ad_2;
output p__cmxig_1;
output p__cmx0ad_3;
output p__cmx0ad_19;
output p__cmx1ad_12;
output p__cmx1ad_23;
output p__cmx1ad_34;
output p__cmxir_0;
output p__cmx0ad_18;
output p__cmx1ad_13;
output p__cmx1ad_22;
output p__cmx1ad_35;
output p__cmxir_1;
output p__cmx0ad_17;
output p__cmx1ad_14;
output p__cmx1ad_25;
output p__cmx1ad_32;
output p__cmx0ad_16;
output p__cmx1ad_15;
output p__cmx1ad_24;
output p__cmx1ad_33;
output p__cmx0ad_26;
output p__cmx1ad_30;
output p__cmx0ad_27;
output p__cmx1ad_31;
output p__cmx0ad_28;
output p__cmx1ad_10;
output p__cmx1ad_21;
output p__cmx0ad_29;
output p__cmx1ad_11;
output p__cmx1ad_20;
wire nv345;
wire n_n13960;
wire n_n13959;
wire nv243;
wire nv294;
wire nv14;
wire nv31;
wire nv43;
wire nv59;
wire nv2;
wire nv349;
wire nv10068;
wire n_n13958;
wire nv437;
wire nv10056;
wire nv499;
wire nv10091;
wire nv10316;
wire nv550;
wire nv10082;
wire n_n13895;
wire nv601;
wire nv10112;
wire nv2153;
wire nv10099;
wire nv3888;
wire nv10135;
wire nv6425;
wire nv10126;
wire nv6437;
wire nv10247;
wire nv8909;
wire nv10143;
wire nv10727;
wire nv8608;
wire n_n424;
wire wire425;
wire wire830;
wire wire856;
wire wire161;
wire wire290;
wire nv10130;
wire wire1289;
wire n_n9245;
wire n_n13643;
wire n_n13271;
wire wire265;
wire wire1323;
wire wire156;
wire wire289;
wire n_n13390;
wire wire711;
wire nv69;
wire nv78;
wire wire326;
wire wire302;
wire wire282;
wire wire514;
wire n_n13789;
wire n_n13786;
wire wire829;
wire wire839;
wire wire911;
wire wire1153;
wire nv251;
wire n_n434;
wire nv6428;
wire wire466;
wire wire594;
wire wire638;
wire wire792;
wire wire988;
wire wire1026;
wire wire1122;
wire wire1299;
wire wire462;
wire wire1002;
wire wire1085;
wire nv10169;
wire wire218;
wire nv354;
wire nv406;
wire nv363;
wire nv401;
wire wire191;
wire wire228;
wire wire260;
wire wire299;
wire wire396;
wire wire412;
wire wire439;
wire wire458;
wire wire1086;
wire n_n1063;
wire wire1343;
wire nv444;
wire wire176;
wire wire262;
wire wire319;
wire wire890;
wire wire177;
wire wire229;
wire wire382;
wire nv10086;
wire n_n450;
wire nv539;
wire wire186;
wire wire630;
wire wire1105;
wire wire1252;
wire wire155;
wire wire190;
wire nv590;
wire n_n11282;
wire nv7447;
wire n_n13096;
wire nv2066;
wire n_n11570;
wire n_n13077;
wire wire175;
wire wire264;
wire wire692;
wire wire708;
wire n_n429;
wire wire510;
wire wire636;
wire nv3311;
wire nv3377;
wire nv3280;
wire nv3369;
wire n_n9587;
wire nv3273;
wire n_n9650;
wire wire158;
wire wire178;
wire wire180;
wire wire294;
wire wire325;
wire wire395;
wire wire399;
wire wire403;
wire wire416;
wire wire438;
wire wire631;
wire wire762;
wire wire1336;
wire n_n8104;
wire wire281;
wire wire509;
wire wire331;
wire wire1165;
wire nv633;
wire wire150;
wire wire172;
wire nv6450;
wire nv10248;
wire n_n13961;
wire wire160;
wire wire202;
wire wire389;
wire wire478;
wire wire725;
wire wire930;
wire wire936;
wire wire1029;
wire nv121;
wire nv158;
wire nv163;
wire n_n13541;
wire n_n13646;
wire n_n13755;
wire n_n13600;
wire wire490;
wire n_n13566;
wire nv116;
wire wire426;
wire wire851;
wire n_n13546;
wire nv212;
wire wire222;
wire wire419;
wire wire318;
wire wire1037;
wire nv222;
wire wire342;
wire wire231;
wire wire768;
wire nv667;
wire wire441;
wire wire269;
wire wire604;
wire wire1032;
wire wire320;
wire wire1097;
wire nv903;
wire nv952;
wire wire157;
wire nv963;
wire nv959;
wire nv758;
wire wire388;
wire wire292;
wire wire357;
wire wire500;
wire n_n12655;
wire nv772;
wire n_n11316;
wire nv699;
wire wire379;
wire wire380;
wire wire1332;
wire nv717;
wire wire184;
wire wire1092;
wire nv1117;
wire nv735;
wire wire1131;
wire nv1138;
wire nv739;
wire nv721;
wire nv1096;
wire nv703;
wire wire459;
wire wire225;
wire wire152;
wire wire272;
wire wire483;
wire wire271;
wire wire211;
wire wire766;
wire wire811;
wire wire816;
wire wire345;
wire wire910;
wire wire1095;
wire nv620;
wire wire317;
wire wire332;
wire nv624;
wire wire1012;
wire nv894;
wire nv890;
wire wire1334;
wire nv923;
wire nv919;
wire n_n12619;
wire wire1039;
wire nv1424;
wire n_n12696;
wire wire436;
wire nv768;
wire wire205;
wire wire1060;
wire nv972;
wire nv968;
wire wire1046;
wire nv1533;
wire nv992;
wire nv988;
wire wire1038;
wire wire224;
wire wire312;
wire nv801;
wire nv797;
wire wire1008;
wire nv914;
wire nv910;
wire wire1312;
wire n_n11076;
wire nv2190;
wire wire1319;
wire nv2176;
wire wire621;
wire nv2186;
wire wire206;
wire wire757;
wire wire924;
wire n_n9294;
wire nv2348;
wire wire365;
wire n_n10860;
wire wire310;
wire wire216;
wire wire314;
wire wire253;
wire wire254;
wire nv2565;
wire wire270;
wire wire347;
wire wire1181;
wire nv2397;
wire wire164;
wire wire240;
wire wire400;
wire wire1194;
wire wire814;
wire wire880;
wire n_n10947;
wire nv2240;
wire wire404;
wire wire847;
wire wire884;
wire n_n10922;
wire n_n10896;
wire wire840;
wire wire881;
wire nv2647;
wire wire321;
wire nv2183;
wire n_n11266;
wire wire907;
wire wire1076;
wire nv2790;
wire n_n9304;
wire n_n10590;
wire n_n10267;
wire wire882;
wire wire1049;
wire wire346;
wire wire1179;
wire n_n10282;
wire nv2622;
wire wire1192;
wire n_n10396;
wire wire1087;
wire nv2946;
wire wire304;
wire wire751;
wire wire866;
wire wire252;
wire wire237;
wire nv2252;
wire nv2235;
wire wire179;
wire wire182;
wire wire166;
wire wire378;
wire nv2340;
wire n_n10835;
wire wire1184;
wire nv2373;
wire wire855;
wire n_n9302;
wire nv3916;
wire wire1281;
wire wire1296;
wire nv3943;
wire n_n8890;
wire nv3918;
wire nv4058;
wire wire870;
wire wire489;
wire wire989;
wire n_n6710;
wire n_n9194;
wire n_n8976;
wire nv3927;
wire wire1180;
wire n_n8862;
wire wire233;
wire wire305;
wire n_n6367;
wire nv3908;
wire nv4045;
wire wire1182;
wire wire632;
wire wire1041;
wire nv4401;
wire wire255;
wire nv3915;
wire n_n7885;
wire wire1065;
wire n_n8085;
wire wire775;
wire nv4932;
wire n_n7095;
wire wire1098;
wire wire834;
wire wire992;
wire wire689;
wire wire1007;
wire n_n8352;
wire wire214;
wire wire374;
wire nv6576;
wire n_n5621;
wire nv669;
wire wire827;
wire wire1047;
wire wire1081;
wire wire721;
wire wire464;
wire n_n2328;
wire n_n4404;
wire nv6462;
wire wire804;
wire n_n4433;
wire wire192;
wire wire196;
wire wire800;
wire n_n4412;
wire n_n5729;
wire n_n4489;
wire wire417;
wire wire193;
wire wire197;
wire wire151;
wire wire173;
wire wire1034;
wire nv7445;
wire n_n3695;
wire nv7647;
wire nv7791;
wire n_n3349;
wire n_n3347;
wire n_n4509;
wire n_n5768;
wire nv10153;
wire n_n4501;
wire n_n5752;
wire n_n5644;
wire n_n3693;
wire n_n5514;
wire nv6589;
wire wire477;
wire wire1074;
wire nv7105;
wire n_n4543;
wire n_n5574;
wire nv6486;
wire nv7050;
wire n_n4473;
wire n_n4611;
wire wire802;
wire nv6472;
wire n_n5580;
wire nv6789;
wire nv8372;
wire n_n3016;
wire nv6859;
wire wire822;
wire wire336;
wire wire1044;
wire wire1063;
wire nv8638;
wire wire405;
wire n_n1241;
wire wire245;
wire wire293;
wire wire316;
wire wire877;
wire wire308;
wire n_n1243;
wire wire1019;
wire wire1075;
wire n_n2176;
wire wire189;
wire wire194;
wire wire295;
wire wire309;
wire wire456;
wire wire700;
wire wire1109;
wire n_n2483;
wire nv839;
wire wire183;
wire wire257;
wire wire476;
wire wire487;
wire wire593;
wire wire626;
wire wire758;
wire wire786;
wire wire1027;
wire wire1322;
wire wire1344;
wire n_n2484;
wire n_n1649;
wire n_n1247;
wire n_n1111;
wire wire361;
wire n_n1119;
wire nv883;
wire n_n1253;
wire n_n1263;
wire n_n1255;
wire wire163;
wire wire171;
wire wire817;
wire n_n1813;
wire wire213;
wire wire506;
wire wire508;
wire wire226;
wire wire154;
wire wire485;
wire nv9492;
wire wire259;
wire nv858;
wire wire853;
wire nv740;
wire n_n1593;
wire nv9031;
wire wire897;
wire n_n2466;
wire wire703;
wire wire999;
wire wire1101;
wire wire278;
wire wire607;
wire wire1082;
wire wire806;
wire n_n2448;
wire wire1304;
wire nv9029;
wire wire341;
wire wire589;
wire n_n2332;
wire wire1146;
wire nv662;
wire nv628;
wire wire418;
wire n_n2327;
wire wire606;
wire n_n1966;
wire wire1302;
wire wire512;
wire nv9129;
wire wire1231;
wire n_n2228;
wire wire461;
wire wire1142;
wire nv9173;
wire n_n2179;
wire n_n2180;
wire wire398;
wire wire770;
wire n_n1566;
wire n_n5610;
wire nv9066;
wire wire951;
wire n_n1574;
wire wire1022;
wire n_n1786;
wire wire952;
wire n_n1756;
wire wire408;
wire wire782;
wire wire860;
wire nv644;
wire n_n13028;
wire wire266;
wire wire348;
wire wire1230;
wire n_n1259;
wire wire327;
wire wire1023;
wire n_n1984;
wire wire701;
wire nv235;
wire wire340;
wire wire381;
wire wire616;
wire n_n12706;
wire nv754;
wire nv942;
wire wire785;
wire nv750;
wire wire1048;
wire nv1162;
wire nv928;
wire wire1036;
wire nv1445;
wire nv873;
wire nv983;
wire nv979;
wire wire1313;
wire wire322;
wire nv2197;
wire wire1111;
wire nv2493;
wire wire238;
wire wire307;
wire wire315;
wire wire706;
wire nv2793;
wire nv3060;
wire nv2534;
wire nv2930;
wire nv2627;
wire nv2330;
wire nv2766;
wire nv2995;
wire nv2314;
wire nv2963;
wire nv2473;
wire nv3109;
wire nv2545;
wire nv3077;
wire nv2857;
wire nv2807;
wire nv2359;
wire wire169;
wire wire763;
wire wire344;
wire wire324;
wire wire1024;
wire wire1061;
wire wire1069;
wire wire1309;
wire wire208;
wire wire1341;
wire n_n9022;
wire nv3961;
wire wire323;
wire wire1185;
wire n_n9141;
wire wire990;
wire n_n8948;
wire wire1103;
wire n_n7845;
wire wire369;
wire wire370;
wire wire613;
wire wire279;
wire wire387;
wire wire473;
wire wire705;
wire wire1028;
wire wire1053;
wire wire1113;
wire wire1203;
wire wire1245;
wire wire1246;
wire wire1288;
wire wire698;
wire wire1031;
wire n_n7837;
wire wire258;
wire n_n9255;
wire wire153;
wire wire437;
wire wire895;
wire wire904;
wire wire1110;
wire n_n7816;
wire n_n7945;
wire n_n7825;
wire wire181;
wire wire227;
wire wire274;
wire wire474;
wire wire765;
wire wire908;
wire wire920;
wire wire1329;
wire wire358;
wire wire1290;
wire wire1292;
wire wire1351;
wire wire201;
wire wire249;
wire wire922;
wire wire1308;
wire n_n7905;
wire wire457;
wire wire1279;
wire n_n7702;
wire n_n6922;
wire wire165;
wire wire268;
wire wire618;
wire wire247;
wire wire818;
wire wire845;
wire wire848;
wire n_n7808;
wire wire311;
wire nv4938;
wire wire991;
wire nv5285;
wire nv4409;
wire wire170;
wire wire484;
wire wire587;
wire wire1118;
wire wire221;
wire wire352;
wire wire263;
wire wire377;
wire wire453;
wire wire699;
wire wire1339;
wire wire788;
wire wire791;
wire nv5843;
wire wire1189;
wire n_n5481;
wire wire801;
wire wire1006;
wire n_n4441;
wire wire826;
wire wire857;
wire wire1064;
wire n_n5520;
wire nv7098;
wire nv7129;
wire wire209;
wire wire199;
wire wire450;
wire wire448;
wire wire251;
wire wire244;
wire wire653;
wire wire203;
wire wire690;
wire wire797;
wire n_n3014;
wire wire335;
wire nv8369;
wire nv10167;
wire wire861;
wire wire501;
wire wire655;
wire wire828;
wire wire1114;
wire wire641;
wire wire673;
wire wire678;
wire wire891;
wire wire1090;
wire wire649;
wire wire652;
wire n_n4481;
wire wire250;
wire wire243;
wire wire898;
wire wire1000;
wire n_n2404;
wire wire820;
wire wire841;
wire wire1248;
wire nv9082;
wire n_n2280;
wire n_n1329;
wire wire1104;
wire n_n2229;
wire wire771;
wire wire934;
wire nv9050;
wire n_n2143;
wire wire1250;
wire wire1196;
wire n_n1891;
wire wire1212;
wire n_n1410;
wire wire835;
wire n_n1394;
wire n_n1858;
wire wire836;
wire wire242;
wire wire974;
wire n_n12782;
wire nv658;
wire wire1310;
wire nv1052;
wire nv764;
wire wire1070;
wire n_n10809;
wire nv2602;
wire nv2694;
wire nv2276;
wire nv2220;
wire nv2641;
wire n_n10412;
wire wire219;
wire wire303;
wire wire313;
wire wire572;
wire wire697;
wire wire953;
wire wire432;
wire wire983;
wire wire1043;
wire wire1080;
wire n_n10795;
wire wire1188;
wire wire794;
wire n_n10796;
wire wire1013;
wire wire1195;
wire wire885;
wire nv2430;
wire wire1186;
wire n_n9177;
wire n_n7913;
wire n_n7877;
wire n_n7893;
wire wire329;
wire wire460;
wire wire1003;
wire wire475;
wire wire611;
wire wire505;
wire nv4389;
wire wire502;
wire wire198;
wire wire449;
wire wire185;
wire wire850;
wire n_n8956;
wire n_n9157;
wire wire187;
wire wire372;
wire wire960;
wire wire442;
wire wire393;
wire nv5283;
wire n_n6749;
wire wire424;
wire wire1284;
wire n_n5908;
wire n_n5604;
wire wire276;
wire wire906;
wire wire963;
wire wire1298;
wire wire1311;
wire wire527;
wire nv7043;
wire wire672;
wire wire832;
wire wire734;
wire wire1306;
wire nv6797;
wire wire1068;
wire wire1123;
wire wire465;
wire wire798;
wire wire468;
wire wire385;
wire wire507;
wire wire1011;
wire wire912;
wire nv8350;
wire n_n2546;
wire wire337;
wire nv6886;
wire wire409;
wire n_n2452;
wire wire1249;
wire n_n5799;
wire n_n2226;
wire n_n1395;
wire nv9297;
wire n_n1859;
wire n_n1558;
wire n_n1229;
wire wire239;
wire nv683;
wire nv1009;
wire nv679;
wire wire1057;
wire nv1073;
wire wire617;
wire wire843;
wire wire1293;
wire wire1014;
wire wire1108;
wire nv821;
wire nv817;
wire wire1318;
wire wire887;
wire wire338;
wire nv6146;
wire nv5862;
wire wire339;
wire wire555;
wire nv6124;
wire n_n7400;
wire wire793;
wire wire833;
wire wire964;
wire wire1316;
wire n_n8112;
wire wire330;
wire wire359;
wire wire401;
wire wire914;
wire wire838;
wire wire1303;
wire nv6104;
wire nv6110;
wire n_n6711;
wire wire684;
wire wire1256;
wire nv6289;
wire wire334;
wire wire574;
wire wire1283;
wire wire1328;
wire wire871;
wire wire928;
wire nv6851;
wire wire204;
wire wire529;
wire wire1096;
wire wire1102;
wire wire446;
wire wire640;
wire wire657;
wire wire1035;
wire wire1340;
wire wire915;
wire wire685;
wire wire447;
wire wire528;
wire n_n1341;
wire n_n1427;
wire n_n1908;
wire n_n1426;
wire wire783;
wire n_n1907;
wire n_n1905;
wire n_n1494;
wire n_n1219;
wire n_n1495;
wire wire975;
wire n_n1491;
wire wire948;
wire wire714;
wire nv1291;
wire nv779;
wire wire1282;
wire nv1183;
wire nv1226;
wire nv1205;
wire nv1270;
wire nv835;
wire nv1249;
wire wire1112;
wire nv783;
wire wire586;
wire wire614;
wire wire1071;
wire wire1210;
wire nv997;
wire wire1058;
wire wire1066;
wire wire1183;
wire wire886;
wire wire883;
wire n_n8968;
wire nv4327;
wire n_n4697;
wire wire1150;
wire n_n4834;
wire n_n4934;
wire wire1091;
wire n_n5328;
wire wire371;
wire wire433;
wire wire585;
wire wire1291;
wire wire899;
wire wire1206;
wire n_n5713;
wire wire273;
wire wire959;
wire wire1285;
wire wire1326;
wire wire422;
wire wire597;
wire wire921;
wire wire837;
wire nv8777;
wire n_n1311;
wire nv9262;
wire n_n2097;
wire n_n2009;
wire n_n2010;
wire n_n2007;
wire n_n1301;
wire nv1556;
wire nv1577;
wire wire1045;
wire wire1073;
wire nv1403;
wire wire248;
wire wire575;
wire wire739;
wire wire1016;
wire wire1093;
wire wire1094;
wire wire1120;
wire wire962;
wire n_n4096;
wire wire918;
wire wire1297;
wire wire1320;
wire n_n1347;
wire n_n1173;
wire n_n1351;
wire wire1275;
wire n_n1335;
wire wire863;
wire wire349;
wire n_n1423;
wire n_n1207;
wire wire878;
wire nv899;
wire wire1033;
wire nv1380;
wire wire943;
wire nv2290;
wire nv2411;
wire wire200;
wire wire916;
wire wire1348;
wire wire486;
wire wire687;
wire wire162;
wire wire968;
wire wire1128;
wire wire492;
wire wire375;
wire nv4630;
wire wire390;
wire wire592;
wire n_n1462;
wire n_n1463;
wire wire972;
wire wire997;
wire wire971;
wire wire1262;
wire n_n1277;
wire n_n1555;
wire n_n1528;
wire wire695;
wire wire970;
wire wire995;
wire wire328;
wire n_n6828;
wire wire306;
wire wire1200;
wire wire230;
wire wire913;
wire wire1324;
wire wire1327;
wire wire691;
wire wire707;
wire wire1198;
wire wire463;
wire wire351;
wire wire727;
wire wire1352;
wire wire1213;
wire n_n1289;
wire n_n1824;
wire n_n1823;
wire n_n1269;
wire n_n1783;
wire wire1264;
wire wire1126;
wire n_n11474;
wire nv1490;
wire nv1359;
wire n_n4541;
wire n_n4542;
wire wire732;
wire wire1337;
wire wire1079;
wire wire1083;
wire wire926;
wire n_n11833;
wire n_n11836;
wire wire368;
wire wire376;
wire wire343;
wire wire812;
wire wire813;
wire n_n12641;
wire wire947;
wire wire1030;
wire nv4575;
wire wire740;
wire wire957;
wire wire722;
wire n_n9515;
wire wire903;
wire n_n9516;
wire wire443;
wire wire754;
wire n_n11295;
wire wire694;
wire nv3202;
wire n_n9647;
wire wire723;
wire wire852;
wire wire933;
wire nv4648;
wire wire1178;
wire n_n8343;
wire n_n7001;
wire n_n6410;
wire wire599;
wire wire391;
wire wire780;
wire wire1211;
wire n_n1992;
wire wire1263;
wire nv10174;
wire nv10178;
wire nv10237;
wire wire980;
wire nv10173;
wire nv10222;
wire nv10162;
wire nv10187;
wire wire493;
wire wire628;
wire wire764;
wire wire868;
wire n_n983;
wire wire480;
wire wire1277;
wire wire499;
wire nv10252;
wire nv4641;
wire wire535;
wire n_n1478;
wire n_n806;
wire wire965;
wire n_n7239;
wire wire188;
wire wire280;
wire wire373;
wire wire440;
wire wire159;
wire wire168;
wire wire283;
wire wire285;
wire wire362;
wire wire367;
wire wire410;
wire wire430;
wire wire445;
wire wire469;
wire wire470;
wire wire479;
wire wire494;
wire wire497;
wire wire511;
wire wire515;
wire wire518;
wire wire520;
wire wire521;
wire wire538;
wire wire539;
wire wire541;
wire wire542;
wire wire544;
wire wire548;
wire wire550;
wire wire551;
wire wire552;
wire wire558;
wire wire559;
wire wire561;
wire wire562;
wire wire563;
wire wire565;
wire wire566;
wire wire568;
wire wire570;
wire wire603;
wire wire609;
wire wire624;
wire wire629;
wire wire651;
wire wire709;
wire wire710;
wire wire724;
wire wire741;
wire wire823;
wire wire825;
wire wire879;
wire wire888;
wire wire894;
wire wire925;
wire wire931;
wire wire932;
wire wire938;
wire wire939;
wire wire944;
wire wire945;
wire wire955;
wire wire956;
wire wire961;
wire wire967;
wire wire969;
wire wire982;
wire wire1001;
wire wire1004;
wire wire1040;
wire wire1042;
wire wire1054;
wire wire1136;
wire wire1137;
wire wire1141;
wire wire1143;
wire wire1145;
wire wire1148;
wire wire1154;
wire wire1155;
wire wire1156;
wire wire1157;
wire wire1159;
wire wire1160;
wire wire1164;
wire wire1166;
wire wire1167;
wire wire1168;
wire wire1169;
wire wire1170;
wire wire1172;
wire wire1174;
wire wire1175;
wire wire1176;
wire wire1191;
wire wire1201;
wire wire1202;
wire wire1207;
wire wire1209;
wire wire1214;
wire wire1215;
wire wire1216;
wire wire1218;
wire wire1221;
wire wire1223;
wire wire1225;
wire wire1228;
wire wire1232;
wire wire1233;
wire wire1235;
wire wire1236;
wire wire1237;
wire wire1238;
wire wire1240;
wire wire1251;
wire wire1254;
wire wire1258;
wire wire1270;
wire wire1273;
wire wire1353;
wire wire1357;
wire wire1358;
wire wire1360;
wire wire1361;
wire wire1362;
wire wire1363;
wire wire1364;
wire wire1365;
wire wire1366;
wire wire1367;
wire wire1371;
wire wire1374;
wire wire1376;
wire wire1380;
wire wire1382;
wire wire1384;
wire wire1385;
wire wire1391;
wire wire1394;
wire wire1395;
wire wire1397;
wire wire1398;
wire wire1400;
wire wire1403;
wire wire1404;
wire wire1406;
wire wire1407;
wire wire1408;
wire wire1416;
wire wire1417;
wire wire1424;
wire wire1426;
wire wire1431;
wire wire1432;
wire wire1433;
wire wire1434;
wire wire1438;
wire wire1439;
wire wire1440;
wire wire1442;
wire wire1444;
wire wire1447;
wire wire1448;
wire wire1454;
wire wire1458;
wire wire1463;
wire wire1465;
wire wire1466;
wire wire1467;
wire wire1471;
wire wire1473;
wire wire1474;
wire wire1479;
wire wire1482;
wire wire1484;
wire wire1485;
wire wire1486;
wire wire1492;
wire wire1493;
wire wire1494;
wire wire1498;
wire wire1501;
wire wire1502;
wire wire1516;
wire wire1517;
wire wire1518;
wire wire1519;
wire wire1535;
wire wire1536;
wire wire1537;
wire wire1538;
wire wire1542;
wire wire1543;
wire wire1547;
wire wire1548;
wire wire1549;
wire wire1550;
wire wire1551;
wire wire1552;
wire wire1553;
wire wire1554;
wire wire1555;
wire wire1556;
wire wire1557;
wire wire1563;
wire wire1566;
wire wire1567;
wire wire1569;
wire wire1571;
wire wire1574;
wire wire1575;
wire wire1578;
wire wire1579;
wire wire1580;
wire wire1585;
wire wire1602;
wire wire1604;
wire wire1606;
wire wire1607;
wire wire1608;
wire wire1610;
wire wire1622;
wire wire1623;
wire wire1625;
wire wire1626;
wire wire1627;
wire wire1628;
wire wire1629;
wire wire1631;
wire wire1634;
wire wire1636;
wire wire1642;
wire wire1643;
wire wire1647;
wire wire1648;
wire wire1649;
wire wire1651;
wire wire1660;
wire wire1662;
wire wire1663;
wire wire1664;
wire wire1665;
wire wire1666;
wire wire1667;
wire wire1668;
wire wire1669;
wire wire1671;
wire wire1672;
wire wire1673;
wire wire1674;
wire wire1676;
wire wire1677;
wire wire1678;
wire wire1680;
wire wire1682;
wire wire1683;
wire wire1684;
wire wire1686;
wire wire1688;
wire wire1689;
wire wire1697;
wire wire1698;
wire wire1699;
wire wire1700;
wire wire1701;
wire wire1705;
wire wire1706;
wire wire1708;
wire wire1710;
wire wire1718;
wire wire1719;
wire wire1720;
wire wire1721;
wire wire1726;
wire wire1732;
wire wire1735;
wire wire1740;
wire wire1742;
wire wire1754;
wire wire1756;
wire wire1763;
wire wire1765;
wire wire1770;
wire wire1772;
wire wire1773;
wire wire1777;
wire wire1783;
wire wire1784;
wire wire1787;
wire wire1791;
wire wire1794;
wire wire1798;
wire wire1803;
wire wire1805;
wire wire1813;
wire wire1827;
wire wire1831;
wire wire1832;
wire wire1833;
wire wire1835;
wire wire1840;
wire wire1845;
wire wire1847;
wire wire1848;
wire wire1849;
wire wire1853;
wire wire1855;
wire wire1860;
wire wire1861;
wire wire1866;
wire wire1872;
wire wire1873;
wire wire1874;
wire wire1875;
wire wire1876;
wire wire1878;
wire wire1879;
wire wire1881;
wire wire1883;
wire wire1886;
wire wire1887;
wire wire1890;
wire wire1892;
wire wire1893;
wire wire1894;
wire wire1895;
wire wire1896;
wire wire1901;
wire wire1903;
wire wire1924;
wire wire1927;
wire wire1928;
wire wire1936;
wire wire1938;
wire wire1941;
wire wire1951;
wire wire1952;
wire wire1953;
wire wire1958;
wire wire1959;
wire wire1970;
wire wire1974;
wire wire1982;
wire wire1983;
wire wire1984;
wire wire1986;
wire wire1987;
wire wire1992;
wire wire1999;
wire wire2001;
wire wire2003;
wire wire2004;
wire wire2005;
wire wire2010;
wire wire2024;
wire wire2025;
wire wire2029;
wire wire2030;
wire wire2035;
wire wire2040;
wire wire2044;
wire wire2045;
wire wire2050;
wire wire2052;
wire wire2054;
wire wire2055;
wire wire2061;
wire wire2062;
wire wire2065;
wire wire2066;
wire wire2067;
wire wire2072;
wire wire2081;
wire wire2083;
wire wire2085;
wire wire2086;
wire wire2087;
wire wire2101;
wire wire2107;
wire wire2108;
wire wire2111;
wire wire2112;
wire wire2115;
wire wire2116;
wire wire2117;
wire wire2118;
wire wire2119;
wire wire2120;
wire wire2121;
wire wire2122;
wire wire2124;
wire wire2126;
wire wire2128;
wire wire2129;
wire wire2130;
wire wire2133;
wire wire2134;
wire wire2137;
wire wire2141;
wire wire2143;
wire wire2145;
wire wire2148;
wire wire2150;
wire wire2151;
wire wire2152;
wire wire2153;
wire wire2154;
wire wire2159;
wire wire2160;
wire wire2165;
wire wire2167;
wire wire2168;
wire wire2169;
wire wire2173;
wire wire2174;
wire wire2175;
wire wire2178;
wire wire2181;
wire wire2182;
wire wire2184;
wire wire2185;
wire wire2187;
wire wire2191;
wire wire2193;
wire wire2197;
wire wire2199;
wire wire2200;
wire wire2201;
wire wire2202;
wire wire2204;
wire wire2207;
wire wire2208;
wire wire2209;
wire wire2210;
wire wire2214;
wire wire2215;
wire wire2216;
wire wire2217;
wire wire2218;
wire wire2220;
wire wire2224;
wire wire2225;
wire wire2227;
wire wire2228;
wire wire2229;
wire wire2230;
wire wire2235;
wire wire2236;
wire wire2237;
wire wire2238;
wire wire2239;
wire wire2240;
wire wire2241;
wire wire2243;
wire wire2244;
wire wire2245;
wire wire2246;
wire wire2250;
wire wire2251;
wire wire2253;
wire wire2254;
wire wire2255;
wire wire2256;
wire wire2257;
wire wire2258;
wire wire2259;
wire wire2260;
wire wire2261;
wire wire2262;
wire wire2263;
wire wire2265;
wire wire2266;
wire wire2267;
wire wire2268;
wire wire2269;
wire wire2270;
wire wire2274;
wire wire2275;
wire wire2277;
wire wire2278;
wire wire2279;
wire wire2285;
wire wire2286;
wire wire2288;
wire wire2289;
wire wire2290;
wire wire2295;
wire wire2298;
wire wire2299;
wire wire2300;
wire wire2301;
wire wire2302;
wire wire2303;
wire wire2304;
wire wire2305;
wire wire2306;
wire wire2308;
wire wire2310;
wire wire2311;
wire wire2313;
wire wire2314;
wire wire2317;
wire wire2318;
wire wire2319;
wire wire2320;
wire wire2321;
wire wire2322;
wire wire2323;
wire wire2324;
wire wire2325;
wire wire2326;
wire wire2327;
wire wire2329;
wire wire2330;
wire wire2331;
wire wire2332;
wire wire2333;
wire wire2334;
wire wire2335;
wire wire2336;
wire wire2341;
wire wire2342;
wire wire2345;
wire wire2346;
wire wire2348;
wire wire2349;
wire wire2350;
wire wire2351;
wire wire2352;
wire wire2353;
wire wire2355;
wire wire2360;
wire wire2364;
wire wire2365;
wire wire2367;
wire wire2368;
wire wire2370;
wire wire2371;
wire wire2374;
wire wire2375;
wire wire2378;
wire wire2379;
wire wire2380;
wire wire2381;
wire wire2382;
wire wire2386;
wire wire2387;
wire wire2389;
wire wire2390;
wire wire2391;
wire wire2398;
wire wire2399;
wire wire2400;
wire wire2402;
wire wire2403;
wire wire2404;
wire wire2406;
wire wire2409;
wire wire2416;
wire wire2418;
wire wire2419;
wire wire2421;
wire wire2422;
wire wire2423;
wire wire2424;
wire wire2426;
wire wire2427;
wire wire2432;
wire wire2433;
wire wire2435;
wire wire2436;
wire wire2437;
wire wire2438;
wire wire2442;
wire wire2446;
wire wire2447;
wire wire2448;
wire wire2456;
wire wire2457;
wire wire2460;
wire wire2469;
wire wire2471;
wire wire2472;
wire wire2474;
wire wire2478;
wire wire2479;
wire wire2482;
wire wire2484;
wire wire2485;
wire wire2486;
wire wire2487;
wire wire2490;
wire wire2491;
wire wire2494;
wire wire2498;
wire wire2499;
wire wire2500;
wire wire2502;
wire wire2508;
wire wire2516;
wire wire2517;
wire wire2519;
wire wire2521;
wire wire2522;
wire wire2524;
wire wire2526;
wire wire2527;
wire wire2529;
wire wire2530;
wire wire2531;
wire wire2532;
wire wire2533;
wire wire2534;
wire wire2538;
wire wire2545;
wire wire2546;
wire wire2547;
wire wire2549;
wire wire2553;
wire wire2554;
wire wire2556;
wire wire2557;
wire wire2558;
wire wire2559;
wire wire2560;
wire wire2562;
wire wire2563;
wire wire2564;
wire wire2566;
wire wire2571;
wire wire2576;
wire wire2585;
wire wire2586;
wire wire2587;
wire wire2591;
wire wire2593;
wire wire2594;
wire wire2595;
wire wire2596;
wire wire2597;
wire wire2600;
wire wire2602;
wire wire2603;
wire wire2604;
wire wire2606;
wire wire2607;
wire wire2608;
wire wire2609;
wire wire2614;
wire wire2615;
wire wire2618;
wire wire2619;
wire wire2620;
wire wire2621;
wire wire2622;
wire wire2624;
wire wire2625;
wire wire2629;
wire wire2631;
wire wire2632;
wire wire2634;
wire wire2635;
wire wire2636;
wire wire2637;
wire wire2639;
wire wire2640;
wire wire2641;
wire wire2642;
wire wire2643;
wire wire2645;
wire wire2646;
wire wire2648;
wire wire2649;
wire wire2652;
wire wire2653;
wire wire2654;
wire wire2655;
wire wire2657;
wire wire2658;
wire wire2659;
wire wire2668;
wire wire2669;
wire wire2671;
wire wire2672;
wire wire2674;
wire wire2675;
wire wire2676;
wire wire2681;
wire wire2684;
wire wire2686;
wire wire2688;
wire wire2691;
wire wire2692;
wire wire2694;
wire wire2695;
wire wire2696;
wire wire2697;
wire wire2698;
wire wire2699;
wire wire2700;
wire wire2701;
wire wire2702;
wire wire2704;
wire wire2705;
wire wire2706;
wire wire2707;
wire wire2708;
wire wire2710;
wire wire2711;
wire wire2713;
wire wire2714;
wire wire2715;
wire wire2717;
wire wire2718;
wire wire2719;
wire wire2720;
wire wire2723;
wire wire2724;
wire wire2729;
wire wire2730;
wire wire2731;
wire wire2732;
wire wire2733;
wire wire2734;
wire wire2735;
wire wire2736;
wire wire2739;
wire wire2741;
wire wire2742;
wire wire2743;
wire wire2744;
wire wire2745;
wire wire2750;
wire wire2752;
wire wire2753;
wire wire2754;
wire wire2755;
wire wire2756;
wire wire2761;
wire wire2762;
wire wire2764;
wire wire2767;
wire wire2770;
wire wire2771;
wire wire2772;
wire wire2775;
wire wire2777;
wire wire2778;
wire wire2780;
wire wire2781;
wire wire2784;
wire wire2785;
wire wire2786;
wire wire2787;
wire wire2788;
wire wire2789;
wire wire2792;
wire wire2794;
wire wire2795;
wire wire2798;
wire wire2800;
wire wire2801;
wire wire2802;
wire wire2803;
wire wire2805;
wire wire2811;
wire wire2812;
wire wire2815;
wire wire2816;
wire wire2817;
wire wire2818;
wire wire2819;
wire wire2820;
wire wire2821;
wire wire2822;
wire wire2826;
wire wire2828;
wire wire2830;
wire wire2831;
wire wire2832;
wire wire2833;
wire wire2834;
wire wire2838;
wire wire2839;
wire wire2840;
wire wire2841;
wire wire2842;
wire wire2845;
wire wire2846;
wire wire2847;
wire wire2850;
wire wire2851;
wire wire2852;
wire wire2855;
wire wire2857;
wire wire2858;
wire wire2860;
wire wire2861;
wire wire2862;
wire wire2863;
wire wire2864;
wire wire2865;
wire wire2866;
wire wire2869;
wire wire2870;
wire wire2871;
wire wire2872;
wire wire2873;
wire wire2875;
wire wire2876;
wire wire2877;
wire wire2878;
wire wire2881;
wire wire2883;
wire wire2884;
wire wire2885;
wire wire2886;
wire wire2889;
wire wire2892;
wire wire2893;
wire wire2894;
wire wire2895;
wire wire2896;
wire wire2897;
wire wire2898;
wire wire2899;
wire wire2900;
wire wire2901;
wire wire2902;
wire wire2906;
wire wire2907;
wire wire2910;
wire wire2911;
wire wire2912;
wire wire2913;
wire wire2915;
wire wire2916;
wire wire2917;
wire wire2918;
wire wire2919;
wire wire2920;
wire wire2926;
wire wire2927;
wire wire2928;
wire wire2932;
wire wire2933;
wire wire2935;
wire wire2936;
wire wire2937;
wire wire2939;
wire wire2946;
wire wire2947;
wire wire2949;
wire wire2950;
wire wire2951;
wire wire2952;
wire wire2954;
wire wire2955;
wire wire2957;
wire wire2958;
wire wire2959;
wire wire2960;
wire wire2961;
wire wire2962;
wire wire2963;
wire wire2964;
wire wire2967;
wire wire2972;
wire wire2980;
wire wire2981;
wire wire2983;
wire wire2984;
wire wire2986;
wire wire2987;
wire wire2990;
wire wire2994;
wire wire2995;
wire wire3000;
wire wire3001;
wire wire3005;
wire wire3006;
wire wire3008;
wire wire3011;
wire wire3015;
wire wire3019;
wire wire3020;
wire wire3023;
wire wire3024;
wire wire3027;
wire wire3030;
wire wire3031;
wire wire3034;
wire wire3036;
wire wire3040;
wire wire3041;
wire wire3042;
wire wire3045;
wire wire3046;
wire wire3047;
wire wire3048;
wire wire3049;
wire wire3050;
wire wire3051;
wire wire3056;
wire wire3057;
wire wire3058;
wire wire3060;
wire wire3064;
wire wire3066;
wire wire3069;
wire wire3074;
wire wire3075;
wire wire3076;
wire wire3083;
wire wire3084;
wire wire3085;
wire wire3086;
wire wire3088;
wire wire3090;
wire wire3091;
wire wire3092;
wire wire3093;
wire wire3096;
wire wire3097;
wire wire3098;
wire wire3099;
wire wire3104;
wire wire3109;
wire wire3110;
wire wire3111;
wire wire3112;
wire wire3114;
wire wire3116;
wire wire3117;
wire wire3118;
wire wire3119;
wire wire3120;
wire wire3121;
wire wire3122;
wire wire3125;
wire wire3126;
wire wire3139;
wire wire3140;
wire wire3141;
wire wire3144;
wire wire3147;
wire wire3149;
wire wire3150;
wire wire3151;
wire wire3153;
wire wire3156;
wire wire3157;
wire wire3158;
wire wire3159;
wire wire3160;
wire wire3161;
wire wire3162;
wire wire3165;
wire wire3166;
wire wire3167;
wire wire3168;
wire wire3169;
wire wire3170;
wire wire3171;
wire wire3173;
wire wire3174;
wire wire3175;
wire wire3176;
wire wire3177;
wire wire3179;
wire wire3182;
wire wire3185;
wire wire3186;
wire wire3187;
wire wire3189;
wire wire3193;
wire wire3195;
wire wire3196;
wire wire3197;
wire wire3199;
wire wire3205;
wire wire3206;
wire wire3214;
wire wire3215;
wire wire3221;
wire wire3222;
wire wire3223;
wire wire3231;
wire wire3233;
wire wire3240;
wire wire3243;
wire wire3246;
wire wire3247;
wire wire3249;
wire wire3251;
wire wire3257;
wire wire3260;
wire wire3266;
wire wire3274;
wire wire3276;
wire wire3277;
wire wire3278;
wire wire3280;
wire wire3292;
wire wire3295;
wire wire3297;
wire wire3301;
wire wire3303;
wire wire3307;
wire wire3308;
wire wire3314;
wire wire3316;
wire wire3318;
wire wire3320;
wire wire3322;
wire wire3326;
wire wire3327;
wire wire3328;
wire wire3337;
wire wire3339;
wire wire3341;
wire wire3349;
wire wire3355;
wire wire3358;
wire wire3375;
wire wire3381;
wire wire3383;
wire wire3387;
wire wire3389;
wire wire3391;
wire wire3393;
wire wire3399;
wire wire3402;
wire wire3405;
wire wire3406;
wire wire3407;
wire wire3410;
wire wire3412;
wire wire3420;
wire wire3426;
wire wire3429;
wire wire3431;
wire wire3435;
wire wire3439;
wire wire3444;
wire wire3448;
wire wire3449;
wire wire3450;
wire wire3453;
wire wire3456;
wire wire3457;
wire wire3458;
wire wire3462;
wire wire3464;
wire wire3466;
wire wire3474;
wire wire3479;
wire wire3482;
wire wire3488;
wire wire3491;
wire wire3493;
wire wire3497;
wire wire3506;
wire wire3512;
wire wire3514;
wire wire3515;
wire wire3516;
wire wire3517;
wire wire3520;
wire wire3521;
wire wire3522;
wire wire3528;
wire wire3529;
wire wire3533;
wire wire3534;
wire wire3537;
wire wire3540;
wire wire3543;
wire wire3544;
wire wire3545;
wire wire3546;
wire wire3547;
wire wire3548;
wire wire3549;
wire wire3551;
wire wire3552;
wire wire3553;
wire wire3554;
wire wire3555;
wire wire3556;
wire wire3557;
wire wire3558;
wire wire3559;
wire wire3561;
wire wire3562;
wire wire3563;
wire wire3564;
wire wire3565;
wire wire3566;
wire wire3567;
wire wire3568;
wire wire3569;
wire wire3571;
wire wire3572;
wire wire3573;
wire wire3576;
wire wire3577;
wire wire3578;
wire wire3580;
wire wire3581;
wire wire3582;
wire wire3584;
wire wire3587;
wire wire3588;
wire wire3589;
wire wire3590;
wire wire3593;
wire wire3594;
wire wire3596;
wire wire3601;
wire wire3602;
wire wire3605;
wire wire3606;
wire wire3607;
wire wire3608;
wire wire3609;
wire wire3610;
wire wire3611;
wire wire3612;
wire wire3615;
wire wire3617;
wire wire3618;
wire wire3623;
wire wire3625;
wire wire3627;
wire wire3628;
wire wire3629;
wire wire3630;
wire wire3631;
wire wire3632;
wire wire3639;
wire wire3641;
wire wire3642;
wire wire3644;
wire wire3645;
wire wire3647;
wire wire3650;
wire wire3651;
wire wire3652;
wire wire3653;
wire wire3655;
wire wire3658;
wire wire3660;
wire wire3661;
wire wire3662;
wire wire3663;
wire wire3664;
wire wire3665;
wire wire3666;
wire wire3667;
wire wire3668;
wire wire3670;
wire wire3676;
wire wire3679;
wire wire3680;
wire wire3681;
wire wire3682;
wire wire3687;
wire wire3690;
wire wire3691;
wire wire3696;
wire wire3698;
wire wire3702;
wire wire3703;
wire wire3704;
wire wire3706;
wire wire3708;
wire wire3709;
wire wire3710;
wire wire3711;
wire wire3712;
wire wire3715;
wire wire3716;
wire wire3717;
wire wire3719;
wire wire3720;
wire wire3721;
wire wire3724;
wire wire3725;
wire wire3727;
wire wire3728;
wire wire3729;
wire wire3730;
wire wire3731;
wire wire3732;
wire wire3735;
wire wire3736;
wire wire3737;
wire wire3739;
wire wire3741;
wire wire3743;
wire wire3744;
wire wire3748;
wire wire3749;
wire wire3750;
wire wire3751;
wire wire3752;
wire wire3755;
wire wire3756;
wire wire3757;
wire wire3759;
wire wire3761;
wire wire3762;
wire wire3763;
wire wire3764;
wire wire3765;
wire wire3768;
wire wire3769;
wire wire3770;
wire wire3773;
wire wire3774;
wire wire3777;
wire wire3778;
wire wire3779;
wire wire3780;
wire wire3782;
wire wire3783;
wire wire3785;
wire wire3786;
wire wire3788;
wire wire3789;
wire wire3792;
wire wire3793;
wire wire3795;
wire wire3796;
wire wire3798;
wire wire3799;
wire wire3801;
wire wire3802;
wire wire3803;
wire wire3804;
wire wire3805;
wire wire3808;
wire wire3809;
wire wire3810;
wire wire3813;
wire wire3814;
wire wire3816;
wire wire3817;
wire wire3818;
wire wire3819;
wire wire3820;
wire wire3821;
wire wire3823;
wire wire3826;
wire wire3827;
wire wire3828;
wire wire3829;
wire wire3830;
wire wire3834;
wire wire3835;
wire wire3838;
wire wire3840;
wire wire3842;
wire wire3843;
wire wire3845;
wire wire3846;
wire wire3849;
wire wire3851;
wire wire3852;
wire wire3855;
wire wire3856;
wire wire3857;
wire wire3858;
wire wire3859;
wire wire3863;
wire wire3864;
wire wire3865;
wire wire3866;
wire wire3867;
wire wire3868;
wire wire3870;
wire wire3874;
wire wire3878;
wire wire3879;
wire wire3880;
wire wire3881;
wire wire3882;
wire wire3883;
wire wire3884;
wire wire3888;
wire wire3889;
wire wire3891;
wire wire3892;
wire wire3893;
wire wire3894;
wire wire3895;
wire wire3896;
wire wire3897;
wire wire3898;
wire wire3899;
wire wire3900;
wire wire3902;
wire wire3903;
wire wire3904;
wire wire3906;
wire wire3907;
wire wire3908;
wire wire3910;
wire wire3912;
wire wire3914;
wire wire3915;
wire wire3916;
wire wire3918;
wire wire3919;
wire wire3920;
wire wire3921;
wire wire3922;
wire wire3923;
wire wire3926;
wire wire3927;
wire wire3929;
wire wire3930;
wire wire3931;
wire wire3934;
wire wire3937;
wire wire3938;
wire wire3939;
wire wire3940;
wire wire3941;
wire wire3942;
wire wire3943;
wire wire3944;
wire wire3945;
wire wire3946;
wire wire3948;
wire wire3950;
wire wire3951;
wire wire3952;
wire wire3955;
wire wire3957;
wire wire3959;
wire wire3961;
wire wire3963;
wire wire3965;
wire wire3969;
wire wire3973;
wire wire3975;
wire wire3977;
wire wire3979;
wire wire3980;
wire wire3981;
wire wire3982;
wire wire3986;
wire wire3987;
wire wire3989;
wire wire3990;
wire wire3991;
wire wire4005;
wire wire4006;
wire wire4017;
wire wire4018;
wire wire4019;
wire wire4020;
wire wire4024;
wire wire4025;
wire wire4027;
wire wire4028;
wire wire4029;
wire wire4037;
wire wire4043;
wire wire4044;
wire wire4046;
wire wire4047;
wire wire4061;
wire wire4062;
wire wire4064;
wire wire4065;
wire wire4066;
wire wire4067;
wire wire4069;
wire wire4070;
wire wire4072;
wire wire4073;
wire wire4077;
wire wire4078;
wire wire4079;
wire wire4082;
wire wire4083;
wire wire4089;
wire wire4090;
wire wire4096;
wire wire4100;
wire wire4101;
wire wire4102;
wire wire4107;
wire wire4108;
wire wire4109;
wire wire4112;
wire wire4113;
wire wire4115;
wire wire4117;
wire wire4118;
wire wire4121;
wire wire4122;
wire wire4123;
wire wire4124;
wire wire4127;
wire wire4128;
wire wire4129;
wire wire4132;
wire wire4134;
wire wire4135;
wire wire4138;
wire wire4139;
wire wire4142;
wire wire4145;
wire wire4147;
wire wire4149;
wire wire4151;
wire wire4158;
wire wire4161;
wire wire4162;
wire wire4163;
wire wire4164;
wire wire4165;
wire wire4167;
wire wire4170;
wire wire4175;
wire wire4176;
wire wire4179;
wire wire4182;
wire wire4183;
wire wire4184;
wire wire4187;
wire wire4189;
wire wire4191;
wire wire4192;
wire wire4193;
wire wire4194;
wire wire4196;
wire wire4197;
wire wire4199;
wire wire4200;
wire wire4201;
wire wire4204;
wire wire4206;
wire wire4208;
wire wire4209;
wire wire4211;
wire wire4213;
wire wire4214;
wire wire4216;
wire wire4217;
wire wire4220;
wire wire4222;
wire wire4226;
wire wire4231;
wire wire4232;
wire wire4235;
wire wire4236;
wire wire4240;
wire wire4241;
wire wire4242;
wire wire4243;
wire wire4244;
wire wire4245;
wire wire4246;
wire wire4247;
wire wire4248;
wire wire4249;
wire wire4250;
wire wire4252;
wire wire4253;
wire wire4254;
wire wire4255;
wire wire4257;
wire wire4258;
wire wire4259;
wire wire4260;
wire wire4263;
wire wire4264;
wire wire4265;
wire wire4266;
wire wire4269;
wire wire4273;
wire wire4276;
wire wire4277;
wire wire4281;
wire wire4282;
wire wire4283;
wire wire4284;
wire wire4286;
wire wire4293;
wire wire4294;
wire wire4295;
wire wire4296;
wire wire4299;
wire wire4300;
wire wire4301;
wire wire4302;
wire wire4303;
wire wire4305;
wire wire4306;
wire wire4307;
wire wire4309;
wire wire4312;
wire wire4313;
wire wire4317;
wire wire4322;
wire wire4323;
wire wire4324;
wire wire4327;
wire wire4331;
wire wire4332;
wire wire4333;
wire wire4334;
wire wire4337;
wire wire4338;
wire wire4341;
wire wire4342;
wire wire4343;
wire wire4344;
wire wire4345;
wire wire4349;
wire wire4350;
wire wire4351;
wire wire4354;
wire wire4357;
wire wire4358;
wire wire4359;
wire wire4361;
wire wire4362;
wire wire4363;
wire wire4365;
wire wire4367;
wire wire4368;
wire wire4369;
wire wire4374;
wire wire4375;
wire wire4376;
wire wire4377;
wire wire4378;
wire wire4383;
wire wire4384;
wire wire4387;
wire wire4392;
wire wire4394;
wire wire4397;
wire wire4400;
wire wire4406;
wire wire4407;
wire wire4409;
wire wire4410;
wire wire4411;
wire wire4415;
wire wire4417;
wire wire4418;
wire wire4419;
wire wire4421;
wire wire4422;
wire wire4423;
wire wire4425;
wire wire4426;
wire wire4428;
wire wire4430;
wire wire4432;
wire wire4433;
wire wire4434;
wire wire4435;
wire wire4436;
wire wire4439;
wire wire4448;
wire wire4449;
wire wire4458;
wire wire4459;
wire wire4462;
wire wire4464;
wire wire4465;
wire wire4466;
wire wire4467;
wire wire4470;
wire wire4471;
wire wire4472;
wire wire4473;
wire wire4474;
wire wire4475;
wire wire4476;
wire wire4478;
wire wire4479;
wire wire4480;
wire wire4481;
wire wire4482;
wire wire4484;
wire wire4491;
wire wire4501;
wire wire4504;
wire wire4505;
wire wire4508;
wire wire4509;
wire wire4510;
wire wire4518;
wire wire4519;
wire wire4520;
wire wire4523;
wire wire4524;
wire wire4525;
wire wire4526;
wire wire4530;
wire wire4531;
wire wire4532;
wire wire4533;
wire wire4536;
wire wire4538;
wire wire4540;
wire wire4544;
wire wire4546;
wire wire4547;
wire wire4548;
wire wire4550;
wire wire4551;
wire wire4553;
wire wire4554;
wire wire4556;
wire wire4558;
wire wire4560;
wire wire4562;
wire wire4564;
wire wire4567;
wire wire4570;
wire wire4574;
wire wire4581;
wire wire4583;
wire wire4585;
wire wire4588;
wire wire4589;
wire wire4590;
wire wire4591;
wire wire4592;
wire wire4596;
wire wire4599;
wire wire4606;
wire wire4607;
wire wire4608;
wire wire4609;
wire wire4613;
wire wire4615;
wire wire4620;
wire wire4624;
wire wire4625;
wire wire4627;
wire wire4632;
wire wire4638;
wire wire4641;
wire wire4642;
wire wire4644;
wire wire4649;
wire wire4651;
wire wire4652;
wire wire4653;
wire wire4655;
wire wire4657;
wire wire4659;
wire wire4660;
wire wire4661;
wire wire4663;
wire wire4667;
wire wire4668;
wire wire4671;
wire wire4674;
wire wire4675;
wire wire4676;
wire wire4678;
wire wire4680;
wire wire4681;
wire wire4685;
wire wire4687;
wire wire4688;
wire wire4690;
wire wire4691;
wire wire4695;
wire wire4697;
wire wire4699;
wire wire4703;
wire wire4704;
wire wire4705;
wire wire4707;
wire wire4709;
wire wire4713;
wire wire4714;
wire wire4717;
wire wire4720;
wire wire4721;
wire wire4722;
wire wire4738;
wire wire4739;
wire wire4743;
wire wire4745;
wire wire4747;
wire wire4751;
wire wire4752;
wire wire4753;
wire wire4757;
wire wire4763;
wire wire4766;
wire wire4767;
wire wire4769;
wire wire4776;
wire wire4778;
wire wire4779;
wire wire4781;
wire wire4782;
wire wire4784;
wire wire4785;
wire wire4787;
wire wire4788;
wire wire4792;
wire wire4793;
wire wire4795;
wire wire4796;
wire wire4797;
wire wire4799;
wire wire4802;
wire wire4803;
wire wire4804;
wire wire4805;
wire wire4807;
wire wire4808;
wire wire4810;
wire wire4811;
wire wire4813;
wire wire4814;
wire wire4817;
wire wire4824;
wire wire4827;
wire wire4833;
wire wire4834;
wire wire4836;
wire wire4837;
wire wire4838;
wire wire4839;
wire wire4843;
wire wire4844;
wire wire4846;
wire wire4847;
wire wire4848;
wire wire4851;
wire wire4853;
wire wire4856;
wire wire4857;
wire wire4861;
wire wire4862;
wire wire4864;
wire wire4865;
wire wire4866;
wire wire4868;
wire wire4875;
wire wire4886;
wire wire4887;
wire wire4889;
wire wire4890;
wire wire4891;
wire wire4892;
wire wire4896;
wire wire4897;
wire wire4899;
wire wire4900;
wire wire4901;
wire wire4904;
wire wire4910;
wire wire4911;
wire wire4912;
wire wire4913;
wire wire4917;
wire wire4921;
wire wire4922;
wire wire4924;
wire wire4925;
wire wire4926;
wire wire4930;
wire wire4931;
wire wire4933;
wire wire4938;
wire wire4942;
wire wire4943;
wire wire4945;
wire wire4950;
wire wire4952;
wire wire4953;
wire wire4957;
wire wire4958;
wire wire4959;
wire wire4967;
wire wire4968;
wire wire4969;
wire wire4970;
wire wire4971;
wire wire4973;
wire wire4981;
wire wire4991;
wire wire4995;
wire wire4997;
wire wire4999;
wire wire5000;
wire wire5002;
wire wire5003;
wire wire5006;
wire wire5009;
wire wire5010;
wire wire5011;
wire wire5012;
wire wire5013;
wire wire5014;
wire wire5015;
wire wire5017;
wire wire5018;
wire wire5019;
wire wire5022;
wire wire5024;
wire wire5025;
wire wire5026;
wire wire5029;
wire wire5030;
wire wire5032;
wire wire5033;
wire wire5034;
wire wire5037;
wire wire5039;
wire wire5040;
wire wire5044;
wire wire5045;
wire wire5046;
wire wire5047;
wire wire5048;
wire wire5049;
wire wire5050;
wire wire5051;
wire wire5052;
wire wire5055;
wire wire5056;
wire wire5058;
wire wire5059;
wire wire5060;
wire wire5063;
wire wire5064;
wire wire5065;
wire wire5066;
wire wire5068;
wire wire5070;
wire wire5071;
wire wire5072;
wire wire5073;
wire wire5075;
wire wire5078;
wire wire5079;
wire wire5080;
wire wire5082;
wire wire5086;
wire wire5087;
wire wire5088;
wire wire5089;
wire wire5090;
wire wire5091;
wire wire5092;
wire wire5094;
wire wire5095;
wire wire5096;
wire wire5097;
wire wire5098;
wire wire5099;
wire wire5101;
wire wire5102;
wire wire5103;
wire wire5107;
wire wire5108;
wire wire5109;
wire wire5110;
wire wire5111;
wire wire5112;
wire wire5113;
wire wire5114;
wire wire5115;
wire wire5116;
wire wire5119;
wire wire5120;
wire wire5125;
wire wire5128;
wire wire5130;
wire wire5131;
wire wire5132;
wire wire5134;
wire wire5135;
wire wire5138;
wire wire5139;
wire wire5140;
wire wire5142;
wire wire5143;
wire wire5144;
wire wire5145;
wire wire5146;
wire wire5148;
wire wire5150;
wire wire5151;
wire wire5152;
wire wire5166;
wire wire5167;
wire wire5168;
wire wire5169;
wire wire5174;
wire wire5178;
wire wire5184;
wire wire5190;
wire wire5196;
wire wire5198;
wire wire5211;
wire wire5215;
wire wire5219;
wire wire5223;
wire wire5239;
wire wire5240;
wire wire5241;
wire wire5242;
wire wire5243;
wire wire5244;
wire wire5245;
wire wire5247;
wire wire5248;
wire wire5249;
wire wire5252;
wire wire5253;
wire wire5254;
wire wire5256;
wire wire5258;
wire wire5261;
wire wire5262;
wire wire5263;
wire wire5264;
wire wire5267;
wire wire5271;
wire wire5273;
wire wire5274;
wire wire5278;
wire wire5279;
wire wire5284;
wire wire5286;
wire wire5287;
wire wire5291;
wire wire5292;
wire wire5300;
wire wire5302;
wire wire5304;
wire wire5305;
wire wire5307;
wire wire5308;
wire wire5309;
wire wire5311;
wire wire5312;
wire wire5315;
wire wire5317;
wire wire5319;
wire wire5325;
wire wire5327;
wire wire5329;
wire wire5334;
wire wire5337;
wire wire5340;
wire wire5344;
wire wire5346;
wire wire5347;
wire wire5348;
wire wire5351;
wire wire5352;
wire wire5353;
wire wire5354;
wire wire5361;
wire wire5362;
wire wire5366;
wire wire5367;
wire wire5368;
wire wire5375;
wire wire5376;
wire wire5377;
wire wire5378;
wire wire5380;
wire wire5381;
wire wire5386;
wire wire5390;
wire wire5391;
wire wire5393;
wire wire5396;
wire wire5397;
wire wire5401;
wire wire5402;
wire wire5404;
wire wire5407;
wire wire5409;
wire wire5414;
wire wire5416;
wire wire5426;
wire wire5429;
wire wire5431;
wire wire5433;
wire wire5435;
wire wire5436;
wire wire5437;
wire wire5439;
wire wire5440;
wire wire5442;
wire wire5443;
wire wire5446;
wire wire5448;
wire wire5450;
wire wire5451;
wire wire5453;
wire wire5454;
wire wire5455;
wire wire5457;
wire wire5463;
wire wire5468;
wire wire5469;
wire wire5470;
wire wire5473;
wire wire5474;
wire wire5475;
wire wire5486;
wire wire5487;
wire wire5494;
wire wire5499;
wire wire5500;
wire wire5501;
wire wire5504;
wire wire5505;
wire wire5507;
wire wire5511;
wire wire5512;
wire wire5513;
wire wire5514;
wire wire5516;
wire wire5517;
wire wire5518;
wire wire5519;
wire wire5520;
wire wire5521;
wire wire5522;
wire wire5523;
wire wire5524;
wire wire5525;
wire wire5528;
wire wire5529;
wire wire5534;
wire wire5535;
wire wire5537;
wire wire5538;
wire wire5539;
wire wire5540;
wire wire5541;
wire wire5542;
wire wire5543;
wire wire5544;
wire wire5545;
wire wire5547;
wire wire5549;
wire wire5553;
wire wire5554;
wire wire5555;
wire wire5557;
wire wire5558;
wire wire5560;
wire wire5561;
wire wire5562;
wire wire5564;
wire wire5565;
wire wire5566;
wire wire5567;
wire wire5576;
wire wire5577;
wire wire5578;
wire wire5579;
wire wire5580;
wire wire5581;
wire wire5583;
wire wire5589;
wire wire5590;
wire wire5591;
wire wire5593;
wire wire5594;
wire wire5598;
wire wire5601;
wire wire5602;
wire wire5603;
wire wire5607;
wire wire5608;
wire wire5610;
wire wire5611;
wire wire5612;
wire wire5613;
wire wire5615;
wire wire5616;
wire wire5618;
wire wire5619;
wire wire5620;
wire wire5621;
wire wire5622;
wire wire5623;
wire wire5624;
wire wire5625;
wire wire5626;
wire wire5627;
wire wire5629;
wire wire5630;
wire wire5632;
wire wire5635;
wire wire5636;
wire wire5637;
wire wire5639;
wire wire5642;
wire wire5643;
wire wire5644;
wire wire5646;
wire wire5647;
wire wire5648;
wire wire5651;
wire wire5653;
wire wire5654;
wire wire5656;
wire wire5657;
wire wire5663;
wire wire5664;
wire wire5665;
wire wire5666;
wire wire5667;
wire wire5668;
wire wire5670;
wire wire5678;
wire wire5682;
wire wire5684;
wire wire5685;
wire wire5687;
wire wire5688;
wire wire5689;
wire wire5693;
wire wire5703;
wire wire5704;
wire wire5705;
wire wire5708;
wire wire5709;
wire wire5710;
wire wire5711;
wire wire5713;
wire wire5714;
wire wire5715;
wire wire5718;
wire wire5723;
wire wire5724;
wire wire5725;
wire wire5728;
wire wire5729;
wire wire5744;
wire wire5745;
wire wire5770;
wire wire5775;
wire wire5778;
wire wire5788;
wire wire5796;
wire wire5797;
wire wire5798;
wire wire5800;
wire wire5801;
wire wire5802;
wire wire5804;
wire wire5808;
wire wire5809;
wire wire5810;
wire wire5812;
wire wire5816;
wire wire5829;
wire wire5837;
wire wire5838;
wire wire5839;
wire wire5841;
wire wire5842;
wire wire5845;
wire wire5847;
wire wire5851;
wire wire5852;
wire wire5855;
wire wire5861;
wire wire5871;
wire wire5873;
wire wire5875;
wire wire5883;
wire wire5884;
wire wire5885;
wire wire5887;
wire wire5889;
wire wire5893;
wire wire5894;
wire wire5895;
wire wire5897;
wire wire5898;
wire wire5902;
wire wire5904;
wire wire5906;
wire wire5914;
wire wire5917;
wire wire5920;
wire wire5921;
wire wire5922;
wire wire5924;
wire wire5926;
wire wire5930;
wire wire5932;
wire wire5935;
wire wire5939;
wire wire5941;
wire wire5945;
wire wire5946;
wire wire5948;
wire wire5960;
wire wire5961;
wire wire5962;
wire wire5963;
wire wire5964;
wire wire5965;
wire wire5966;
wire wire5967;
wire wire5968;
wire wire5975;
wire wire5976;
wire wire5978;
wire wire5979;
wire wire5982;
wire wire5983;
wire wire5984;
wire wire5987;
wire wire5988;
wire wire5989;
wire wire5990;
wire wire5992;
wire wire5999;
wire wire6001;
wire wire6003;
wire wire6004;
wire wire6007;
wire wire6011;
wire wire6012;
wire wire6013;
wire wire6016;
wire wire6017;
wire wire6018;
wire wire6019;
wire wire6025;
wire wire6027;
wire wire6028;
wire wire6030;
wire wire6032;
wire wire6035;
wire wire6038;
wire wire6040;
wire wire6041;
wire wire6042;
wire wire6047;
wire wire6049;
wire wire6050;
wire wire6056;
wire wire6059;
wire wire6062;
wire wire6066;
wire wire6074;
wire wire6077;
wire wire6079;
wire wire6081;
wire wire6087;
wire wire6089;
wire wire6095;
wire wire6103;
wire wire6105;
wire wire6111;
wire wire6114;
wire wire6119;
wire wire6122;
wire wire6123;
wire wire6124;
wire wire6127;
wire wire6132;
wire wire6135;
wire wire6138;
wire wire6140;
wire wire6143;
wire wire6145;
wire wire6152;
wire wire6154;
wire wire6155;
wire wire6156;
wire wire6157;
wire wire6159;
wire wire6161;
wire wire6165;
wire wire6169;
wire wire6170;
wire wire6171;
wire wire6172;
wire wire6174;
wire wire6176;
wire wire6177;
wire wire6179;
wire wire6180;
wire wire6182;
wire wire6184;
wire wire6185;
wire wire6189;
wire wire6190;
wire wire6192;
wire wire6193;
wire wire6196;
wire wire6198;
wire wire6200;
wire wire6202;
wire wire6205;
wire wire6206;
wire wire6207;
wire wire6209;
wire wire6210;
wire wire6217;
wire wire6224;
wire wire6225;
wire wire6226;
wire wire6228;
wire wire6230;
wire wire6231;
wire wire6235;
wire wire6236;
wire wire6239;
wire wire6240;
wire wire6242;
wire wire6243;
wire wire6246;
wire wire6247;
wire wire6249;
wire wire6252;
wire wire6253;
wire wire6255;
wire wire6269;
wire wire6270;
wire wire6271;
wire wire6272;
wire wire6276;
wire wire6281;
wire wire6284;
wire wire6285;
wire wire6287;
wire wire6291;
wire wire6293;
wire wire6295;
wire wire6297;
wire wire6305;
wire wire6308;
wire wire6309;
wire wire6312;
wire wire6314;
wire wire6315;
wire wire6316;
wire wire6318;
wire wire6319;
wire wire6325;
wire wire6326;
wire wire6329;
wire wire6330;
wire wire6332;
wire wire6333;
wire wire6334;
wire wire6337;
wire wire6351;
wire wire6354;
wire wire6355;
wire wire6366;
wire wire6401;
wire wire6402;
wire wire6429;
wire wire6450;
wire wire6453;
wire wire6454;
wire wire6457;
wire wire6475;
wire wire6479;
wire wire6498;
wire wire6499;
wire wire6501;
wire wire6503;
wire wire6505;
wire wire6506;
wire wire6508;
wire wire6509;
wire wire6513;
wire wire6514;
wire wire6515;
wire wire6517;
wire wire6521;
wire wire6524;
wire wire6531;
wire wire6536;
wire wire6537;
wire wire6538;
wire wire6540;
wire wire6541;
wire wire6543;
wire wire6547;
wire wire6549;
wire wire6551;
wire wire6556;
wire wire6557;
wire wire6558;
wire wire6560;
wire wire6561;
wire wire6563;
wire wire6567;
wire wire6569;
wire wire6571;
wire wire6576;
wire wire6577;
wire wire6578;
wire wire6580;
wire wire6581;
wire wire6583;
wire wire6612;
wire wire6613;
wire wire6614;
wire wire6616;
wire wire6617;
wire wire6619;
wire wire6626;
wire wire6628;
wire wire6629;
wire wire6630;
wire wire6633;
wire wire6634;
wire wire6636;
wire wire6640;
wire wire6642;
wire wire6644;
wire wire6647;
wire wire6652;
wire wire6653;
wire wire6655;
wire wire6657;
wire wire6662;
wire wire6663;
wire wire6664;
wire wire6666;
wire wire6667;
wire wire6669;
wire wire6678;
wire wire6679;
wire wire6680;
wire wire6682;
wire wire6683;
wire wire6685;
wire wire6691;
wire wire6692;
wire wire6694;
wire wire6696;
wire wire6701;
wire wire6702;
wire wire6703;
wire wire6705;
wire wire6706;
wire wire6708;
wire wire6714;
wire wire6717;
wire wire6721;
wire wire6722;
wire wire6727;
wire wire6729;
wire wire6731;
wire wire6736;
wire wire6741;
wire wire6742;
wire wire6743;
wire wire6745;
wire wire6746;
wire wire6750;
wire wire6757;
wire wire6758;
wire wire6766;
wire wire6775;
wire wire6780;
wire wire6783;
wire wire6784;
wire wire6785;
wire wire6786;
wire wire6787;
wire wire6788;
wire wire6789;
wire wire6790;
wire wire6795;
wire wire6796;
wire wire6797;
wire wire6799;
wire wire6800;
wire wire6801;
wire wire6802;
wire wire6805;
wire wire6808;
wire wire6809;
wire wire6811;
wire wire6812;
wire wire6814;
wire wire6815;
wire wire6816;
wire wire6818;
wire wire6819;
wire wire6820;
wire wire6821;
wire wire6822;
wire wire6824;
wire wire6826;
wire wire6827;
wire wire6829;
wire wire6831;
wire wire6832;
wire wire6833;
wire wire6834;
wire wire6835;
wire wire6836;
wire wire6838;
wire wire6839;
wire wire6842;
wire wire6844;
wire wire6845;
wire wire6846;
wire wire6847;
wire wire6848;
wire wire6852;
wire wire6854;
wire wire6855;
wire wire6857;
wire wire6858;
wire wire6860;
wire wire6862;
wire wire6864;
wire wire6868;
wire wire6869;
wire wire6870;
wire wire6871;
wire wire6873;
wire wire6874;
wire wire6878;
wire wire6880;
wire wire6883;
wire wire6884;
wire wire6889;
wire wire6890;
wire wire6891;
wire wire6898;
wire wire6899;
wire wire6906;
wire wire6908;
wire wire6909;
wire wire6923;
wire wire6925;
wire wire6926;
wire wire6930;
wire wire6932;
wire wire6935;
wire wire6936;
wire wire6938;
wire wire6940;
wire wire6945;
wire wire6946;
wire wire6949;
wire wire6950;
wire wire6951;
wire wire6952;
wire wire6954;
wire wire6955;
wire wire6956;
wire wire6959;
wire wire6965;
wire wire6966;
wire wire6968;
wire wire6969;
wire wire6973;
wire wire6975;
wire wire6976;
wire wire6978;
wire wire6979;
wire wire6980;
wire wire6986;
wire wire6989;
wire wire6990;
wire wire6991;
wire wire6992;
wire wire6995;
wire wire6996;
wire wire6997;
wire wire6999;
wire wire7000;
wire wire7008;
wire wire7009;
wire wire7010;
wire wire7011;
wire wire7025;
wire wire7027;
wire wire7028;
wire wire7029;
wire wire7030;
wire wire7031;
wire wire7032;
wire wire7035;
wire wire7042;
wire wire7043;
wire wire7044;
wire wire7049;
wire wire7055;
wire wire7056;
wire wire7057;
wire wire7058;
wire wire7059;
wire wire7060;
wire wire7070;
wire wire7072;
wire wire7077;
wire wire7080;
wire wire7087;
wire wire7088;
wire wire7089;
wire wire7090;
wire wire7091;
wire wire7093;
wire wire7095;
wire wire7096;
wire wire7097;
wire wire7099;
wire wire7100;
wire wire7101;
wire wire7107;
wire wire7109;
wire wire7118;
wire wire7119;
wire wire7120;
wire wire7121;
wire wire7122;
wire wire7123;
wire wire7126;
wire wire7129;
wire wire7134;
wire wire7140;
wire wire7144;
wire wire7169;
wire wire7170;
wire wire7172;
wire wire7173;
wire wire7174;
wire wire7175;
wire wire7176;
wire wire7180;
wire wire7181;
wire wire7184;
wire wire7193;
wire wire7194;
wire wire7195;
wire wire28695;
wire wire28698;
wire wire28700;
wire wire28702;
wire wire28705;
wire wire28706;
wire wire28708;
wire wire28710;
wire wire28711;
wire wire28712;
wire wire28713;
wire wire28715;
wire wire28716;
wire wire28718;
wire wire28721;
wire wire28724;
wire wire28729;
wire wire28731;
wire wire28734;
wire wire28735;
wire wire28739;
wire wire28743;
wire wire28746;
wire wire28747;
wire wire28751;
wire wire28755;
wire wire28757;
wire wire28758;
wire wire28760;
wire wire28763;
wire wire28764;
wire wire28765;
wire wire28766;
wire wire28767;
wire wire28770;
wire wire28771;
wire wire28773;
wire wire28775;
wire wire28777;
wire wire28779;
wire wire28781;
wire wire28783;
wire wire28784;
wire wire28786;
wire wire28787;
wire wire28789;
wire wire28790;
wire wire28792;
wire wire28796;
wire wire28798;
wire wire28800;
wire wire28802;
wire wire28805;
wire wire28808;
wire wire28812;
wire wire28815;
wire wire28818;
wire wire28821;
wire wire28822;
wire wire28825;
wire wire28826;
wire wire28829;
wire wire28831;
wire wire28834;
wire wire28838;
wire wire28839;
wire wire28840;
wire wire28842;
wire wire28845;
wire wire28846;
wire wire28848;
wire wire28849;
wire wire28850;
wire wire28851;
wire wire28852;
wire wire28854;
wire wire28855;
wire wire28858;
wire wire28859;
wire wire28863;
wire wire28868;
wire wire28870;
wire wire28873;
wire wire28875;
wire wire28878;
wire wire28882;
wire wire28883;
wire wire28885;
wire wire28886;
wire wire28888;
wire wire28891;
wire wire28892;
wire wire28895;
wire wire28897;
wire wire28898;
wire wire28899;
wire wire28901;
wire wire28902;
wire wire28905;
wire wire28906;
wire wire28910;
wire wire28912;
wire wire28913;
wire wire28914;
wire wire28917;
wire wire28918;
wire wire28919;
wire wire28921;
wire wire28922;
wire wire28923;
wire wire28924;
wire wire28926;
wire wire28927;
wire wire28929;
wire wire28930;
wire wire28931;
wire wire28933;
wire wire28934;
wire wire28935;
wire wire28936;
wire wire28937;
wire wire28938;
wire wire28939;
wire wire28940;
wire wire28944;
wire wire28945;
wire wire28946;
wire wire28949;
wire wire28951;
wire wire28952;
wire wire28954;
wire wire28955;
wire wire28956;
wire wire28959;
wire wire28961;
wire wire28962;
wire wire28963;
wire wire28964;
wire wire28965;
wire wire28966;
wire wire28967;
wire wire28969;
wire wire28971;
wire wire28974;
wire wire28976;
wire wire28977;
wire wire28978;
wire wire28979;
wire wire28980;
wire wire28981;
wire wire28983;
wire wire28986;
wire wire28987;
wire wire28989;
wire wire28990;
wire wire28991;
wire wire28995;
wire wire28999;
wire wire29003;
wire wire29005;
wire wire29006;
wire wire29009;
wire wire29012;
wire wire29015;
wire wire29018;
wire wire29021;
wire wire29022;
wire wire29023;
wire wire29026;
wire wire29027;
wire wire29029;
wire wire29030;
wire wire29033;
wire wire29035;
wire wire29037;
wire wire29038;
wire wire29039;
wire wire29040;
wire wire29041;
wire wire29042;
wire wire29046;
wire wire29050;
wire wire29051;
wire wire29054;
wire wire29057;
wire wire29062;
wire wire29063;
wire wire29067;
wire wire29068;
wire wire29069;
wire wire29070;
wire wire29077;
wire wire29078;
wire wire29079;
wire wire29080;
wire wire29081;
wire wire29082;
wire wire29086;
wire wire29088;
wire wire29089;
wire wire29092;
wire wire29094;
wire wire29095;
wire wire29097;
wire wire29098;
wire wire29099;
wire wire29100;
wire wire29101;
wire wire29102;
wire wire29106;
wire wire29108;
wire wire29111;
wire wire29113;
wire wire29115;
wire wire29117;
wire wire29119;
wire wire29121;
wire wire29122;
wire wire29123;
wire wire29124;
wire wire29125;
wire wire29126;
wire wire29127;
wire wire29128;
wire wire29130;
wire wire29131;
wire wire29136;
wire wire29139;
wire wire29142;
wire wire29144;
wire wire29145;
wire wire29148;
wire wire29149;
wire wire29151;
wire wire29153;
wire wire29155;
wire wire29157;
wire wire29158;
wire wire29159;
wire wire29160;
wire wire29163;
wire wire29165;
wire wire29166;
wire wire29167;
wire wire29168;
wire wire29169;
wire wire29170;
wire wire29171;
wire wire29176;
wire wire29179;
wire wire29181;
wire wire29182;
wire wire29187;
wire wire29188;
wire wire29192;
wire wire29193;
wire wire29194;
wire wire29195;
wire wire29198;
wire wire29203;
wire wire29204;
wire wire29206;
wire wire29207;
wire wire29209;
wire wire29210;
wire wire29211;
wire wire29214;
wire wire29215;
wire wire29217;
wire wire29219;
wire wire29223;
wire wire29225;
wire wire29226;
wire wire29228;
wire wire29231;
wire wire29233;
wire wire29234;
wire wire29236;
wire wire29237;
wire wire29240;
wire wire29241;
wire wire29242;
wire wire29244;
wire wire29247;
wire wire29248;
wire wire29249;
wire wire29252;
wire wire29253;
wire wire29256;
wire wire29259;
wire wire29261;
wire wire29264;
wire wire29268;
wire wire29269;
wire wire29270;
wire wire29271;
wire wire29273;
wire wire29274;
wire wire29276;
wire wire29277;
wire wire29279;
wire wire29280;
wire wire29282;
wire wire29283;
wire wire29286;
wire wire29288;
wire wire29289;
wire wire29291;
wire wire29292;
wire wire29294;
wire wire29296;
wire wire29297;
wire wire29298;
wire wire29299;
wire wire29300;
wire wire29303;
wire wire29306;
wire wire29308;
wire wire29310;
wire wire29311;
wire wire29313;
wire wire29315;
wire wire29316;
wire wire29317;
wire wire29319;
wire wire29320;
wire wire29323;
wire wire29324;
wire wire29325;
wire wire29326;
wire wire29328;
wire wire29331;
wire wire29333;
wire wire29334;
wire wire29335;
wire wire29336;
wire wire29337;
wire wire29338;
wire wire29340;
wire wire29343;
wire wire29344;
wire wire29345;
wire wire29346;
wire wire29347;
wire wire29348;
wire wire29352;
wire wire29353;
wire wire29354;
wire wire29358;
wire wire29360;
wire wire29361;
wire wire29362;
wire wire29366;
wire wire29367;
wire wire29368;
wire wire29371;
wire wire29372;
wire wire29376;
wire wire29377;
wire wire29379;
wire wire29382;
wire wire29385;
wire wire29386;
wire wire29388;
wire wire29393;
wire wire29394;
wire wire29395;
wire wire29397;
wire wire29398;
wire wire29400;
wire wire29403;
wire wire29404;
wire wire29407;
wire wire29408;
wire wire29410;
wire wire29411;
wire wire29413;
wire wire29414;
wire wire29415;
wire wire29417;
wire wire29418;
wire wire29419;
wire wire29420;
wire wire29423;
wire wire29424;
wire wire29425;
wire wire29427;
wire wire29429;
wire wire29430;
wire wire29431;
wire wire29433;
wire wire29437;
wire wire29438;
wire wire29440;
wire wire29441;
wire wire29444;
wire wire29447;
wire wire29449;
wire wire29451;
wire wire29452;
wire wire29454;
wire wire29455;
wire wire29458;
wire wire29460;
wire wire29461;
wire wire29462;
wire wire29465;
wire wire29466;
wire wire29467;
wire wire29468;
wire wire29469;
wire wire29470;
wire wire29471;
wire wire29472;
wire wire29473;
wire wire29474;
wire wire29475;
wire wire29476;
wire wire29479;
wire wire29481;
wire wire29485;
wire wire29486;
wire wire29488;
wire wire29490;
wire wire29491;
wire wire29495;
wire wire29496;
wire wire29497;
wire wire29498;
wire wire29499;
wire wire29501;
wire wire29502;
wire wire29504;
wire wire29505;
wire wire29506;
wire wire29507;
wire wire29508;
wire wire29510;
wire wire29512;
wire wire29513;
wire wire29514;
wire wire29515;
wire wire29517;
wire wire29518;
wire wire29520;
wire wire29521;
wire wire29525;
wire wire29526;
wire wire29527;
wire wire29528;
wire wire29529;
wire wire29530;
wire wire29531;
wire wire29532;
wire wire29533;
wire wire29534;
wire wire29536;
wire wire29537;
wire wire29538;
wire wire29539;
wire wire29540;
wire wire29542;
wire wire29543;
wire wire29544;
wire wire29545;
wire wire29548;
wire wire29550;
wire wire29553;
wire wire29554;
wire wire29555;
wire wire29556;
wire wire29561;
wire wire29562;
wire wire29563;
wire wire29564;
wire wire29565;
wire wire29566;
wire wire29567;
wire wire29568;
wire wire29569;
wire wire29570;
wire wire29571;
wire wire29572;
wire wire29574;
wire wire29575;
wire wire29576;
wire wire29577;
wire wire29578;
wire wire29579;
wire wire29581;
wire wire29582;
wire wire29583;
wire wire29584;
wire wire29586;
wire wire29587;
wire wire29588;
wire wire29589;
wire wire29590;
wire wire29591;
wire wire29592;
wire wire29593;
wire wire29594;
wire wire29595;
wire wire29596;
wire wire29597;
wire wire29598;
wire wire29599;
wire wire29600;
wire wire29601;
wire wire29602;
wire wire29603;
wire wire29604;
wire wire29605;
wire wire29606;
wire wire29609;
wire wire29610;
wire wire29611;
wire wire29612;
wire wire29615;
wire wire29616;
wire wire29617;
wire wire29619;
wire wire29621;
wire wire29622;
wire wire29623;
wire wire29624;
wire wire29625;
wire wire29626;
wire wire29627;
wire wire29628;
wire wire29629;
wire wire29630;
wire wire29631;
wire wire29632;
wire wire29634;
wire wire29635;
wire wire29636;
wire wire29637;
wire wire29639;
wire wire29641;
wire wire29642;
wire wire29644;
wire wire29645;
wire wire29647;
wire wire29648;
wire wire29649;
wire wire29650;
wire wire29651;
wire wire29652;
wire wire29653;
wire wire29655;
wire wire29656;
wire wire29657;
wire wire29658;
wire wire29659;
wire wire29660;
wire wire29662;
wire wire29663;
wire wire29664;
wire wire29665;
wire wire29666;
wire wire29669;
wire wire29670;
wire wire29672;
wire wire29674;
wire wire29675;
wire wire29677;
wire wire29680;
wire wire29681;
wire wire29682;
wire wire29684;
wire wire29685;
wire wire29686;
wire wire29687;
wire wire29690;
wire wire29691;
wire wire29692;
wire wire29693;
wire wire29695;
wire wire29697;
wire wire29699;
wire wire29700;
wire wire29702;
wire wire29703;
wire wire29704;
wire wire29706;
wire wire29707;
wire wire29709;
wire wire29710;
wire wire29711;
wire wire29713;
wire wire29715;
wire wire29716;
wire wire29717;
wire wire29718;
wire wire29719;
wire wire29720;
wire wire29721;
wire wire29723;
wire wire29724;
wire wire29726;
wire wire29727;
wire wire29729;
wire wire29730;
wire wire29733;
wire wire29735;
wire wire29736;
wire wire29739;
wire wire29741;
wire wire29743;
wire wire29745;
wire wire29746;
wire wire29748;
wire wire29749;
wire wire29751;
wire wire29752;
wire wire29753;
wire wire29754;
wire wire29756;
wire wire29757;
wire wire29759;
wire wire29760;
wire wire29761;
wire wire29762;
wire wire29763;
wire wire29764;
wire wire29765;
wire wire29766;
wire wire29767;
wire wire29768;
wire wire29769;
wire wire29770;
wire wire29771;
wire wire29773;
wire wire29774;
wire wire29775;
wire wire29776;
wire wire29779;
wire wire29781;
wire wire29782;
wire wire29784;
wire wire29786;
wire wire29789;
wire wire29790;
wire wire29792;
wire wire29793;
wire wire29794;
wire wire29796;
wire wire29797;
wire wire29798;
wire wire29799;
wire wire29800;
wire wire29802;
wire wire29803;
wire wire29805;
wire wire29806;
wire wire29807;
wire wire29808;
wire wire29809;
wire wire29810;
wire wire29811;
wire wire29812;
wire wire29813;
wire wire29815;
wire wire29816;
wire wire29818;
wire wire29819;
wire wire29821;
wire wire29823;
wire wire29825;
wire wire29827;
wire wire29829;
wire wire29830;
wire wire29831;
wire wire29835;
wire wire29836;
wire wire29838;
wire wire29839;
wire wire29842;
wire wire29843;
wire wire29846;
wire wire29847;
wire wire29848;
wire wire29849;
wire wire29851;
wire wire29852;
wire wire29854;
wire wire29855;
wire wire29856;
wire wire29857;
wire wire29858;
wire wire29859;
wire wire29860;
wire wire29861;
wire wire29862;
wire wire29863;
wire wire29864;
wire wire29865;
wire wire29866;
wire wire29868;
wire wire29869;
wire wire29871;
wire wire29873;
wire wire29876;
wire wire29877;
wire wire29878;
wire wire29880;
wire wire29884;
wire wire29885;
wire wire29886;
wire wire29888;
wire wire29890;
wire wire29892;
wire wire29894;
wire wire29896;
wire wire29898;
wire wire29900;
wire wire29902;
wire wire29905;
wire wire29908;
wire wire29910;
wire wire29912;
wire wire29914;
wire wire29916;
wire wire29918;
wire wire29920;
wire wire29922;
wire wire29924;
wire wire29926;
wire wire29929;
wire wire29932;
wire wire29933;
wire wire29937;
wire wire29940;
wire wire29943;
wire wire29945;
wire wire29946;
wire wire29947;
wire wire29948;
wire wire29949;
wire wire29950;
wire wire29951;
wire wire29952;
wire wire29954;
wire wire29955;
wire wire29958;
wire wire29959;
wire wire29960;
wire wire29961;
wire wire29962;
wire wire29963;
wire wire29964;
wire wire29965;
wire wire29967;
wire wire29968;
wire wire29970;
wire wire29972;
wire wire29973;
wire wire29975;
wire wire29977;
wire wire29979;
wire wire29981;
wire wire29982;
wire wire29985;
wire wire29987;
wire wire29990;
wire wire29992;
wire wire29993;
wire wire29994;
wire wire29995;
wire wire29996;
wire wire29997;
wire wire29998;
wire wire29999;
wire wire30001;
wire wire30003;
wire wire30004;
wire wire30006;
wire wire30007;
wire wire30010;
wire wire30011;
wire wire30013;
wire wire30014;
wire wire30016;
wire wire30018;
wire wire30019;
wire wire30023;
wire wire30025;
wire wire30026;
wire wire30027;
wire wire30028;
wire wire30029;
wire wire30031;
wire wire30032;
wire wire30033;
wire wire30034;
wire wire30035;
wire wire30036;
wire wire30038;
wire wire30040;
wire wire30041;
wire wire30042;
wire wire30043;
wire wire30044;
wire wire30046;
wire wire30047;
wire wire30049;
wire wire30051;
wire wire30052;
wire wire30054;
wire wire30055;
wire wire30057;
wire wire30058;
wire wire30059;
wire wire30060;
wire wire30061;
wire wire30063;
wire wire30064;
wire wire30068;
wire wire30069;
wire wire30071;
wire wire30072;
wire wire30073;
wire wire30074;
wire wire30075;
wire wire30076;
wire wire30078;
wire wire30079;
wire wire30081;
wire wire30084;
wire wire30085;
wire wire30086;
wire wire30090;
wire wire30091;
wire wire30093;
wire wire30094;
wire wire30096;
wire wire30099;
wire wire30100;
wire wire30103;
wire wire30106;
wire wire30108;
wire wire30111;
wire wire30113;
wire wire30114;
wire wire30115;
wire wire30117;
wire wire30118;
wire wire30119;
wire wire30121;
wire wire30123;
wire wire30125;
wire wire30126;
wire wire30128;
wire wire30129;
wire wire30131;
wire wire30133;
wire wire30134;
wire wire30135;
wire wire30138;
wire wire30140;
wire wire30142;
wire wire30146;
wire wire30147;
wire wire30148;
wire wire30149;
wire wire30150;
wire wire30151;
wire wire30152;
wire wire30153;
wire wire30154;
wire wire30156;
wire wire30157;
wire wire30158;
wire wire30160;
wire wire30162;
wire wire30163;
wire wire30164;
wire wire30165;
wire wire30166;
wire wire30168;
wire wire30169;
wire wire30171;
wire wire30173;
wire wire30174;
wire wire30176;
wire wire30177;
wire wire30178;
wire wire30179;
wire wire30181;
wire wire30182;
wire wire30183;
wire wire30185;
wire wire30187;
wire wire30188;
wire wire30189;
wire wire30191;
wire wire30192;
wire wire30194;
wire wire30195;
wire wire30197;
wire wire30198;
wire wire30200;
wire wire30202;
wire wire30204;
wire wire30205;
wire wire30208;
wire wire30209;
wire wire30210;
wire wire30212;
wire wire30213;
wire wire30216;
wire wire30217;
wire wire30218;
wire wire30219;
wire wire30220;
wire wire30223;
wire wire30224;
wire wire30226;
wire wire30227;
wire wire30228;
wire wire30231;
wire wire30232;
wire wire30235;
wire wire30236;
wire wire30238;
wire wire30240;
wire wire30241;
wire wire30243;
wire wire30246;
wire wire30248;
wire wire30250;
wire wire30253;
wire wire30254;
wire wire30257;
wire wire30259;
wire wire30260;
wire wire30263;
wire wire30265;
wire wire30267;
wire wire30268;
wire wire30270;
wire wire30272;
wire wire30273;
wire wire30275;
wire wire30277;
wire wire30279;
wire wire30280;
wire wire30282;
wire wire30283;
wire wire30285;
wire wire30286;
wire wire30287;
wire wire30288;
wire wire30289;
wire wire30290;
wire wire30291;
wire wire30292;
wire wire30293;
wire wire30294;
wire wire30296;
wire wire30297;
wire wire30299;
wire wire30301;
wire wire30302;
wire wire30304;
wire wire30305;
wire wire30306;
wire wire30307;
wire wire30308;
wire wire30309;
wire wire30310;
wire wire30311;
wire wire30313;
wire wire30314;
wire wire30315;
wire wire30316;
wire wire30317;
wire wire30318;
wire wire30321;
wire wire30322;
wire wire30323;
wire wire30326;
wire wire30327;
wire wire30328;
wire wire30329;
wire wire30332;
wire wire30333;
wire wire30336;
wire wire30337;
wire wire30338;
wire wire30340;
wire wire30342;
wire wire30344;
wire wire30346;
wire wire30348;
wire wire30349;
wire wire30351;
wire wire30352;
wire wire30354;
wire wire30356;
wire wire30358;
wire wire30359;
wire wire30360;
wire wire30362;
wire wire30364;
wire wire30367;
wire wire30368;
wire wire30369;
wire wire30370;
wire wire30371;
wire wire30372;
wire wire30374;
wire wire30375;
wire wire30378;
wire wire30379;
wire wire30380;
wire wire30381;
wire wire30382;
wire wire30383;
wire wire30384;
wire wire30385;
wire wire30388;
wire wire30389;
wire wire30390;
wire wire30392;
wire wire30393;
wire wire30397;
wire wire30399;
wire wire30402;
wire wire30404;
wire wire30407;
wire wire30408;
wire wire30409;
wire wire30410;
wire wire30413;
wire wire30414;
wire wire30416;
wire wire30417;
wire wire30419;
wire wire30422;
wire wire30423;
wire wire30424;
wire wire30425;
wire wire30426;
wire wire30427;
wire wire30430;
wire wire30431;
wire wire30432;
wire wire30433;
wire wire30435;
wire wire30436;
wire wire30438;
wire wire30439;
wire wire30441;
wire wire30442;
wire wire30444;
wire wire30445;
wire wire30446;
wire wire30449;
wire wire30450;
wire wire30451;
wire wire30452;
wire wire30455;
wire wire30456;
wire wire30458;
wire wire30461;
wire wire30463;
wire wire30465;
wire wire30467;
wire wire30468;
wire wire30470;
wire wire30472;
wire wire30473;
wire wire30475;
wire wire30477;
wire wire30478;
wire wire30480;
wire wire30482;
wire wire30483;
wire wire30484;
wire wire30485;
wire wire30487;
wire wire30489;
wire wire30491;
wire wire30493;
wire wire30494;
wire wire30496;
wire wire30497;
wire wire30499;
wire wire30501;
wire wire30502;
wire wire30503;
wire wire30505;
wire wire30507;
wire wire30509;
wire wire30510;
wire wire30511;
wire wire30512;
wire wire30515;
wire wire30517;
wire wire30519;
wire wire30521;
wire wire30522;
wire wire30524;
wire wire30525;
wire wire30526;
wire wire30527;
wire wire30528;
wire wire30530;
wire wire30531;
wire wire30532;
wire wire30534;
wire wire30536;
wire wire30537;
wire wire30538;
wire wire30540;
wire wire30541;
wire wire30542;
wire wire30543;
wire wire30544;
wire wire30547;
wire wire30548;
wire wire30549;
wire wire30550;
wire wire30552;
wire wire30553;
wire wire30554;
wire wire30557;
wire wire30558;
wire wire30560;
wire wire30561;
wire wire30562;
wire wire30563;
wire wire30564;
wire wire30566;
wire wire30567;
wire wire30568;
wire wire30569;
wire wire30570;
wire wire30572;
wire wire30573;
wire wire30574;
wire wire30577;
wire wire30578;
wire wire30579;
wire wire30580;
wire wire30581;
wire wire30584;
wire wire30586;
wire wire30588;
wire wire30589;
wire wire30590;
wire wire30592;
wire wire30596;
wire wire30597;
wire wire30598;
wire wire30600;
wire wire30601;
wire wire30602;
wire wire30603;
wire wire30604;
wire wire30605;
wire wire30610;
wire wire30612;
wire wire30613;
wire wire30614;
wire wire30616;
wire wire30620;
wire wire30621;
wire wire30622;
wire wire30624;
wire wire30626;
wire wire30628;
wire wire30629;
wire wire30630;
wire wire30631;
wire wire30634;
wire wire30636;
wire wire30638;
wire wire30639;
wire wire30640;
wire wire30641;
wire wire30644;
wire wire30646;
wire wire30648;
wire wire30649;
wire wire30650;
wire wire30651;
wire wire30652;
wire wire30653;
wire wire30654;
wire wire30655;
wire wire30657;
wire wire30659;
wire wire30661;
wire wire30663;
wire wire30664;
wire wire30665;
wire wire30667;
wire wire30668;
wire wire30669;
wire wire30670;
wire wire30671;
wire wire30673;
wire wire30675;
wire wire30677;
wire wire30679;
wire wire30680;
wire wire30681;
wire wire30683;
wire wire30685;
wire wire30687;
wire wire30689;
wire wire30691;
wire wire30692;
wire wire30696;
wire wire30697;
wire wire30700;
wire wire30701;
wire wire30704;
wire wire30705;
wire wire30707;
wire wire30708;
wire wire30709;
wire wire30711;
wire wire30712;
wire wire30713;
wire wire30714;
wire wire30715;
wire wire30716;
wire wire30717;
wire wire30718;
wire wire30719;
wire wire30720;
wire wire30721;
wire wire30722;
wire wire30723;
wire wire30726;
wire wire30728;
wire wire30729;
wire wire30730;
wire wire30731;
wire wire30732;
wire wire30733;
wire wire30735;
wire wire30737;
wire wire30738;
wire wire30740;
wire wire30742;
wire wire30746;
wire wire30748;
wire wire30749;
wire wire30752;
wire wire30754;
wire wire30755;
wire wire30756;
wire wire30758;
wire wire30759;
wire wire30762;
wire wire30764;
wire wire30765;
wire wire30767;
wire wire30770;
wire wire30772;
wire wire30773;
wire wire30775;
wire wire30776;
wire wire30777;
wire wire30778;
wire wire30779;
wire wire30781;
wire wire30782;
wire wire30784;
wire wire30785;
wire wire30786;
wire wire30788;
wire wire30789;
wire wire30791;
wire wire30793;
wire wire30794;
wire wire30795;
wire wire30797;
wire wire30798;
wire wire30799;
wire wire30800;
wire wire30801;
wire wire30802;
wire wire30803;
wire wire30804;
wire wire30805;
wire wire30806;
wire wire30807;
wire wire30808;
wire wire30813;
wire wire30814;
wire wire30815;
wire wire30817;
wire wire30819;
wire wire30820;
wire wire30823;
wire wire30825;
wire wire30826;
wire wire30827;
wire wire30828;
wire wire30829;
wire wire30832;
wire wire30833;
wire wire30834;
wire wire30835;
wire wire30836;
wire wire30837;
wire wire30838;
wire wire30839;
wire wire30840;
wire wire30841;
wire wire30842;
wire wire30843;
wire wire30844;
wire wire30845;
wire wire30846;
wire wire30847;
wire wire30848;
wire wire30849;
wire wire30850;
wire wire30852;
wire wire30853;
wire wire30854;
wire wire30855;
wire wire30857;
wire wire30858;
wire wire30859;
wire wire30862;
wire wire30863;
wire wire30865;
wire wire30866;
wire wire30869;
wire wire30873;
wire wire30875;
wire wire30876;
wire wire30877;
wire wire30880;
wire wire30882;
wire wire30883;
wire wire30885;
wire wire30887;
wire wire30888;
wire wire30889;
wire wire30890;
wire wire30891;
wire wire30893;
wire wire30894;
wire wire30895;
wire wire30896;
wire wire30897;
wire wire30898;
wire wire30899;
wire wire30900;
wire wire30901;
wire wire30902;
wire wire30903;
wire wire30904;
wire wire30905;
wire wire30906;
wire wire30907;
wire wire30909;
wire wire30910;
wire wire30912;
wire wire30913;
wire wire30914;
wire wire30915;
wire wire30916;
wire wire30917;
wire wire30918;
wire wire30919;
wire wire30920;
wire wire30921;
wire wire30922;
wire wire30923;
wire wire30924;
wire wire30925;
wire wire30927;
wire wire30928;
wire wire30929;
wire wire30930;
wire wire30931;
wire wire30933;
wire wire30935;
wire wire30936;
wire wire30938;
wire wire30940;
wire wire30941;
wire wire30944;
wire wire30947;
wire wire30948;
wire wire30949;
wire wire30950;
wire wire30951;
wire wire30952;
wire wire30953;
wire wire30954;
wire wire30955;
wire wire30956;
wire wire30957;
wire wire30959;
wire wire30960;
wire wire30962;
wire wire30963;
wire wire30964;
wire wire30966;
wire wire30967;
wire wire30968;
wire wire30969;
wire wire30973;
wire wire30974;
wire wire30976;
wire wire30977;
wire wire30980;
wire wire30981;
wire wire30982;
wire wire30983;
wire wire30984;
wire wire30985;
wire wire30986;
wire wire30987;
wire wire30988;
wire wire30989;
wire wire30990;
wire wire30991;
wire wire30993;
wire wire30994;
wire wire30996;
wire wire30999;
wire wire31001;
wire wire31002;
wire wire31005;
wire wire31007;
wire wire31008;
wire wire31009;
wire wire31012;
wire wire31014;
wire wire31015;
wire wire31018;
wire wire31019;
wire wire31022;
wire wire31023;
wire wire31028;
wire wire31032;
wire wire31033;
wire wire31034;
wire wire31037;
wire wire31038;
wire wire31039;
wire wire31040;
wire wire31041;
wire wire31042;
wire wire31043;
wire wire31045;
wire wire31047;
wire wire31049;
wire wire31050;
wire wire31052;
wire wire31055;
wire wire31056;
wire wire31058;
wire wire31059;
wire wire31060;
wire wire31061;
wire wire31062;
wire wire31063;
wire wire31064;
wire wire31065;
wire wire31066;
wire wire31067;
wire wire31068;
wire wire31069;
wire wire31071;
wire wire31072;
wire wire31074;
wire wire31077;
wire wire31079;
wire wire31081;
wire wire31082;
wire wire31085;
wire wire31086;
wire wire31087;
wire wire31088;
wire wire31089;
wire wire31090;
wire wire31092;
wire wire31093;
wire wire31098;
wire wire31099;
wire wire31101;
wire wire31104;
wire wire31105;
wire wire31106;
wire wire31107;
wire wire31108;
wire wire31109;
wire wire31110;
wire wire31112;
wire wire31113;
wire wire31114;
wire wire31115;
wire wire31118;
wire wire31119;
wire wire31121;
wire wire31122;
wire wire31125;
wire wire31130;
wire wire31131;
wire wire31132;
wire wire31136;
wire wire31137;
wire wire31139;
wire wire31140;
wire wire31141;
wire wire31142;
wire wire31144;
wire wire31145;
wire wire31147;
wire wire31148;
wire wire31149;
wire wire31152;
wire wire31155;
wire wire31157;
wire wire31159;
wire wire31160;
wire wire31161;
wire wire31162;
wire wire31163;
wire wire31164;
wire wire31165;
wire wire31166;
wire wire31167;
wire wire31168;
wire wire31169;
wire wire31170;
wire wire31171;
wire wire31172;
wire wire31173;
wire wire31176;
wire wire31177;
wire wire31178;
wire wire31179;
wire wire31180;
wire wire31181;
wire wire31183;
wire wire31184;
wire wire31185;
wire wire31187;
wire wire31188;
wire wire31190;
wire wire31191;
wire wire31192;
wire wire31193;
wire wire31194;
wire wire31195;
wire wire31196;
wire wire31198;
wire wire31199;
wire wire31200;
wire wire31202;
wire wire31203;
wire wire31204;
wire wire31206;
wire wire31207;
wire wire31208;
wire wire31209;
wire wire31211;
wire wire31212;
wire wire31213;
wire wire31214;
wire wire31216;
wire wire31218;
wire wire31220;
wire wire31222;
wire wire31223;
wire wire31227;
wire wire31229;
wire wire31232;
wire wire31233;
wire wire31236;
wire wire31238;
wire wire31240;
wire wire31241;
wire wire31242;
wire wire31244;
wire wire31247;
wire wire31249;
wire wire31250;
wire wire31252;
wire wire31253;
wire wire31254;
wire wire31257;
wire wire31258;
wire wire31260;
wire wire31262;
wire wire31263;
wire wire31264;
wire wire31265;
wire wire31266;
wire wire31267;
wire wire31269;
wire wire31270;
wire wire31271;
wire wire31273;
wire wire31274;
wire wire31276;
wire wire31277;
wire wire31278;
wire wire31279;
wire wire31280;
wire wire31281;
wire wire31282;
wire wire31284;
wire wire31285;
wire wire31286;
wire wire31288;
wire wire31289;
wire wire31290;
wire wire31292;
wire wire31293;
wire wire31294;
wire wire31295;
wire wire31297;
wire wire31298;
wire wire31300;
wire wire31302;
wire wire31303;
wire wire31304;
wire wire31306;
wire wire31308;
wire wire31309;
wire wire31313;
wire wire31315;
wire wire31318;
wire wire31319;
wire wire31322;
wire wire31324;
wire wire31326;
wire wire31327;
wire wire31328;
wire wire31330;
wire wire31333;
wire wire31335;
wire wire31336;
wire wire31338;
wire wire31339;
wire wire31340;
wire wire31343;
wire wire31345;
wire wire31346;
wire wire31347;
wire wire31348;
wire wire31350;
wire wire31352;
wire wire31353;
wire wire31355;
wire wire31356;
wire wire31357;
wire wire31358;
wire wire31360;
wire wire31361;
wire wire31362;
wire wire31364;
wire wire31366;
wire wire31367;
wire wire31368;
wire wire31370;
wire wire31371;
wire wire31372;
wire wire31373;
wire wire31375;
wire wire31376;
wire wire31377;
wire wire31379;
wire wire31380;
wire wire31382;
wire wire31384;
wire wire31385;
wire wire31387;
wire wire31388;
wire wire31390;
wire wire31392;
wire wire31393;
wire wire31396;
wire wire31398;
wire wire31399;
wire wire31401;
wire wire31403;
wire wire31404;
wire wire31406;
wire wire31408;
wire wire31410;
wire wire31412;
wire wire31414;
wire wire31415;
wire wire31417;
wire wire31418;
wire wire31420;
wire wire31425;
wire wire31426;
wire wire31427;
wire wire31428;
wire wire31429;
wire wire31430;
wire wire31434;
wire wire31435;
wire wire31437;
wire wire31438;
wire wire31439;
wire wire31440;
wire wire31442;
wire wire31443;
wire wire31444;
wire wire31446;
wire wire31448;
wire wire31449;
wire wire31450;
wire wire31452;
wire wire31453;
wire wire31454;
wire wire31455;
wire wire31457;
wire wire31458;
wire wire31459;
wire wire31461;
wire wire31462;
wire wire31464;
wire wire31466;
wire wire31467;
wire wire31469;
wire wire31470;
wire wire31471;
wire wire31474;
wire wire31476;
wire wire31478;
wire wire31480;
wire wire31481;
wire wire31483;
wire wire31485;
wire wire31486;
wire wire31488;
wire wire31490;
wire wire31492;
wire wire31494;
wire wire31496;
wire wire31497;
wire wire31499;
wire wire31500;
wire wire31502;
wire wire31507;
wire wire31508;
wire wire31509;
wire wire31510;
wire wire31511;
wire wire31512;
wire wire31516;
wire wire31517;
wire wire31518;
wire wire31519;
wire wire31520;
wire wire31521;
wire wire31523;
wire wire31524;
wire wire31525;
wire wire31527;
wire wire31528;
wire wire31530;
wire wire31531;
wire wire31532;
wire wire31533;
wire wire31534;
wire wire31535;
wire wire31536;
wire wire31538;
wire wire31539;
wire wire31540;
wire wire31542;
wire wire31543;
wire wire31544;
wire wire31546;
wire wire31547;
wire wire31548;
wire wire31549;
wire wire31551;
wire wire31552;
wire wire31554;
wire wire31556;
wire wire31557;
wire wire31558;
wire wire31560;
wire wire31562;
wire wire31563;
wire wire31567;
wire wire31569;
wire wire31572;
wire wire31573;
wire wire31576;
wire wire31578;
wire wire31580;
wire wire31581;
wire wire31582;
wire wire31584;
wire wire31587;
wire wire31589;
wire wire31590;
wire wire31592;
wire wire31593;
wire wire31594;
wire wire31596;
wire wire31598;
wire wire31599;
wire wire31601;
wire wire31602;
wire wire31603;
wire wire31604;
wire wire31606;
wire wire31607;
wire wire31608;
wire wire31610;
wire wire31612;
wire wire31613;
wire wire31614;
wire wire31616;
wire wire31617;
wire wire31618;
wire wire31619;
wire wire31621;
wire wire31622;
wire wire31623;
wire wire31625;
wire wire31626;
wire wire31628;
wire wire31630;
wire wire31631;
wire wire31633;
wire wire31634;
wire wire31635;
wire wire31638;
wire wire31640;
wire wire31642;
wire wire31644;
wire wire31645;
wire wire31647;
wire wire31649;
wire wire31650;
wire wire31652;
wire wire31654;
wire wire31656;
wire wire31658;
wire wire31660;
wire wire31661;
wire wire31663;
wire wire31664;
wire wire31666;
wire wire31671;
wire wire31672;
wire wire31673;
wire wire31674;
wire wire31675;
wire wire31676;
wire wire31680;
wire wire31681;
wire wire31683;
wire wire31684;
wire wire31685;
wire wire31686;
wire wire31688;
wire wire31689;
wire wire31690;
wire wire31692;
wire wire31694;
wire wire31695;
wire wire31696;
wire wire31698;
wire wire31699;
wire wire31700;
wire wire31701;
wire wire31703;
wire wire31704;
wire wire31705;
wire wire31707;
wire wire31708;
wire wire31710;
wire wire31712;
wire wire31713;
wire wire31715;
wire wire31716;
wire wire31718;
wire wire31720;
wire wire31721;
wire wire31724;
wire wire31726;
wire wire31727;
wire wire31729;
wire wire31731;
wire wire31732;
wire wire31734;
wire wire31736;
wire wire31738;
wire wire31740;
wire wire31742;
wire wire31743;
wire wire31745;
wire wire31746;
wire wire31748;
wire wire31753;
wire wire31754;
wire wire31755;
wire wire31756;
wire wire31757;
wire wire31758;
wire wire31762;
wire wire31763;
wire wire31764;
wire wire31765;
wire wire31766;
wire wire31767;
wire wire31769;
wire wire31770;
wire wire31771;
wire wire31773;
wire wire31774;
wire wire31776;
wire wire31777;
wire wire31778;
wire wire31779;
wire wire31780;
wire wire31781;
wire wire31782;
wire wire31784;
wire wire31785;
wire wire31786;
wire wire31788;
wire wire31789;
wire wire31790;
wire wire31792;
wire wire31793;
wire wire31794;
wire wire31795;
wire wire31797;
wire wire31798;
wire wire31799;
wire wire31800;
wire wire31802;
wire wire31804;
wire wire31806;
wire wire31808;
wire wire31809;
wire wire31813;
wire wire31815;
wire wire31818;
wire wire31819;
wire wire31822;
wire wire31824;
wire wire31826;
wire wire31827;
wire wire31828;
wire wire31830;
wire wire31833;
wire wire31835;
wire wire31836;
wire wire31838;
wire wire31839;
wire wire31840;
wire wire31842;
wire wire31844;
wire wire31846;
wire wire31849;
wire wire31851;
wire wire31852;
wire wire31855;
wire wire31858;
wire wire31859;
wire wire31861;
wire wire31864;
wire wire31865;
wire wire31866;
wire wire31869;
wire wire31870;
wire wire31875;
wire wire31876;
wire wire31878;
wire wire31880;
wire wire31882;
wire wire31883;
wire wire31884;
wire wire31885;
wire wire31886;
wire wire31887;
wire wire31888;
wire wire31889;
wire wire31890;
wire wire31891;
wire wire31892;
wire wire31893;
wire wire31894;
wire wire31895;
wire wire31896;
wire wire31897;
wire wire31898;
wire wire31899;
wire wire31900;
wire wire31903;
wire wire31905;
wire wire31906;
wire wire31912;
wire wire31913;
wire wire31914;
wire wire31916;
wire wire31917;
wire wire31918;
wire wire31919;
wire wire31921;
wire wire31922;
wire wire31924;
wire wire31926;
wire wire31928;
wire wire31930;
wire wire31931;
wire wire31932;
wire wire31933;
wire wire31934;
wire wire31935;
wire wire31936;
wire wire31937;
wire wire31939;
wire wire31940;
wire wire31941;
wire wire31943;
wire wire31944;
wire wire31945;
wire wire31946;
wire wire31947;
wire wire31948;
wire wire31949;
wire wire31950;
wire wire31952;
wire wire31954;
wire wire31955;
wire wire31956;
wire wire31957;
wire wire31958;
wire wire31959;
wire wire31960;
wire wire31962;
wire wire31964;
wire wire31967;
wire wire31968;
wire wire31971;
wire wire31972;
wire wire31975;
wire wire31976;
wire wire31979;
wire wire31983;
wire wire31984;
wire wire31985;
wire wire31988;
wire wire31989;
wire wire31990;
wire wire31992;
wire wire31994;
wire wire31995;
wire wire31996;
wire wire31997;
wire wire31998;
wire wire31999;
wire wire32000;
wire wire32001;
wire wire32002;
wire wire32003;
wire wire32004;
wire wire32005;
wire wire32006;
wire wire32009;
wire wire32010;
wire wire32011;
wire wire32012;
wire wire32013;
wire wire32014;
wire wire32016;
wire wire32017;
wire wire32018;
wire wire32019;
wire wire32022;
wire wire32024;
wire wire32025;
wire wire32026;
wire wire32027;
wire wire32029;
wire wire32030;
wire wire32032;
wire wire32033;
wire wire32036;
wire wire32037;
wire wire32040;
wire wire32041;
wire wire32042;
wire wire32043;
wire wire32045;
wire wire32046;
wire wire32047;
wire wire32050;
wire wire32051;
wire wire32053;
wire wire32054;
wire wire32055;
wire wire32056;
wire wire32057;
wire wire32059;
wire wire32061;
wire wire32063;
wire wire32064;
wire wire32065;
wire wire32066;
wire wire32068;
wire wire32069;
wire wire32070;
wire wire32074;
wire wire32076;
wire wire32077;
wire wire32078;
wire wire32079;
wire wire32081;
wire wire32082;
wire wire32083;
wire wire32084;
wire wire32085;
wire wire32086;
wire wire32089;
wire wire32090;
wire wire32091;
wire wire32092;
wire wire32094;
wire wire32095;
wire wire32096;
wire wire32097;
wire wire32099;
wire wire32100;
wire wire32103;
wire wire32104;
wire wire32106;
wire wire32107;
wire wire32109;
wire wire32110;
wire wire32111;
wire wire32112;
wire wire32113;
wire wire32114;
wire wire32116;
wire wire32118;
wire wire32122;
wire wire32124;
wire wire32125;
wire wire32126;
wire wire32130;
wire wire32132;
wire wire32134;
wire wire32137;
wire wire32138;
wire wire32139;
wire wire32141;
wire wire32143;
wire wire32144;
wire wire32145;
wire wire32146;
wire wire32148;
wire wire32149;
wire wire32150;
wire wire32151;
wire wire32152;
wire wire32155;
wire wire32156;
wire wire32157;
wire wire32159;
wire wire32161;
wire wire32162;
wire wire32164;
wire wire32165;
wire wire32168;
wire wire32170;
wire wire32171;
wire wire32173;
wire wire32177;
wire wire32178;
wire wire32181;
wire wire32182;
wire wire32184;
wire wire32186;
wire wire32188;
wire wire32189;
wire wire32191;
wire wire32193;
wire wire32194;
wire wire32196;
wire wire32197;
wire wire32199;
wire wire32200;
wire wire32202;
wire wire32203;
wire wire32206;
wire wire32207;
wire wire32208;
wire wire32210;
wire wire32212;
wire wire32214;
wire wire32216;
wire wire32217;
wire wire32219;
wire wire32221;
wire wire32222;
wire wire32223;
wire wire32224;
wire wire32225;
wire wire32226;
wire wire32227;
wire wire32228;
wire wire32230;
wire wire32231;
wire wire32232;
wire wire32233;
wire wire32235;
wire wire32236;
wire wire32237;
wire wire32238;
wire wire32239;
wire wire32241;
wire wire32243;
wire wire32244;
wire wire32249;
wire wire32250;
wire wire32251;
wire wire32252;
wire wire32253;
wire wire32254;
wire wire32256;
wire wire32257;
wire wire32258;
wire wire32260;
wire wire32261;
wire wire32262;
wire wire32264;
wire wire32267;
wire wire32271;
wire wire32272;
wire wire32273;
wire wire32274;
wire wire32275;
wire wire32277;
wire wire32280;
wire wire32281;
wire wire32282;
wire wire32283;
wire wire32285;
wire wire32288;
wire wire32289;
wire wire32290;
wire wire32291;
wire wire32292;
wire wire32293;
wire wire32294;
wire wire32296;
wire wire32297;
wire wire32299;
wire wire32300;
wire wire32301;
wire wire32303;
wire wire32304;
wire wire32306;
wire wire32308;
wire wire32309;
wire wire32314;
wire wire32315;
wire wire32316;
wire wire32318;
wire wire32319;
wire wire32322;
wire wire32325;
wire wire32330;
wire wire32331;
wire wire32332;
wire wire32334;
wire wire32335;
wire wire32338;
wire wire32340;
wire wire32341;
wire wire32344;
wire wire32349;
wire wire32352;
wire wire32354;
wire wire32355;
wire wire32356;
wire wire32357;
wire wire32358;
wire wire32359;
wire wire32360;
wire wire32361;
wire wire32362;
wire wire32363;
wire wire32364;
wire wire32365;
wire wire32367;
wire wire32368;
wire wire32369;
wire wire32370;
wire wire32371;
wire wire32372;
wire wire32373;
wire wire32375;
wire wire32378;
wire wire32380;
wire wire32382;
wire wire32384;
wire wire32386;
wire wire32387;
wire wire32388;
wire wire32390;
wire wire32391;
wire wire32392;
wire wire32394;
wire wire32395;
wire wire32396;
wire wire32398;
wire wire32401;
wire wire32402;
wire wire32403;
wire wire32406;
wire wire32408;
wire wire32409;
wire wire32410;
wire wire32411;
wire wire32413;
wire wire32415;
wire wire32416;
wire wire32417;
wire wire32418;
wire wire32419;
wire wire32420;
wire wire32421;
wire wire32422;
wire wire32424;
wire wire32425;
wire wire32427;
wire wire32428;
wire wire32430;
wire wire32431;
wire wire32432;
wire wire32433;
wire wire32434;
wire wire32437;
wire wire32438;
wire wire32439;
wire wire32440;
wire wire32442;
wire wire32443;
wire wire32444;
wire wire32446;
wire wire32447;
wire wire32449;
wire wire32450;
wire wire32451;
wire wire32452;
wire wire32453;
wire wire32454;
wire wire32455;
wire wire32456;
wire wire32458;
wire wire32459;
wire wire32463;
wire wire32464;
wire wire32467;
wire wire32468;
wire wire32473;
wire wire32474;
wire wire32476;
wire wire32477;
wire wire32478;
wire wire32481;
wire wire32483;
wire wire32485;
wire wire32486;
wire wire32488;
wire wire32489;
wire wire32490;
wire wire32491;
wire wire32492;
wire wire32493;
wire wire32494;
wire wire32495;
wire wire32496;
wire wire32497;
wire wire32498;
wire wire32499;
wire wire32500;
wire wire32501;
wire wire32502;
wire wire32503;
wire wire32504;
wire wire32505;
wire wire32507;
wire wire32508;
wire wire32509;
wire wire32510;
wire wire32511;
wire wire32513;
wire wire32515;
wire wire32516;
wire wire32518;
wire wire32519;
wire wire32522;
wire wire32523;
wire wire32524;
wire wire32525;
wire wire32527;
wire wire32528;
wire wire32529;
wire wire32531;
wire wire32532;
wire wire32534;
wire wire32535;
wire wire32536;
wire wire32537;
wire wire32538;
wire wire32539;
wire wire32540;
wire wire32542;
wire wire32543;
wire wire32545;
wire wire32546;
wire wire32548;
wire wire32549;
wire wire32550;
wire wire32551;
wire wire32552;
wire wire32553;
wire wire32554;
wire wire32555;
wire wire32556;
wire wire32558;
wire wire32559;
wire wire32563;
wire wire32564;
wire wire32567;
wire wire32568;
wire wire32571;
wire wire32573;
wire wire32576;
wire wire32578;
wire wire32580;
wire wire32581;
wire wire32583;
wire wire32586;
wire wire32587;
wire wire32589;
wire wire32591;
wire wire32592;
wire wire32595;
wire wire32596;
wire wire32599;
wire wire32602;
wire wire32605;
wire wire32606;
wire wire32608;
wire wire32609;
wire wire32611;
wire wire32613;
wire wire32614;
wire wire32616;
wire wire32617;
wire wire32619;
wire wire32621;
wire wire32622;
wire wire32624;
wire wire32627;
wire wire32628;
wire wire32629;
wire wire32630;
wire wire32631;
wire wire32633;
wire wire32634;
wire wire32635;
wire wire32636;
wire wire32638;
wire wire32639;
wire wire32640;
wire wire32641;
wire wire32643;
wire wire32645;
wire wire32647;
wire wire32648;
wire wire32649;
wire wire32651;
wire wire32652;
wire wire32654;
wire wire32655;
wire wire32657;
wire wire32659;
wire wire32660;
wire wire32661;
wire wire32662;
wire wire32663;
wire wire32664;
wire wire32665;
wire wire32666;
wire wire32667;
wire wire32668;
wire wire32669;
wire wire32671;
wire wire32672;
wire wire32673;
wire wire32676;
wire wire32677;
wire wire32678;
wire wire32680;
wire wire32681;
wire wire32682;
wire wire32684;
wire wire32685;
wire wire32687;
wire wire32689;
wire wire32690;
wire wire32691;
wire wire32692;
wire wire32693;
wire wire32694;
wire wire32695;
wire wire32696;
wire wire32697;
wire wire32700;
wire wire32702;
wire wire32703;
wire wire32704;
wire wire32706;
wire wire32709;
wire wire32710;
wire wire32711;
wire wire32712;
wire wire32714;
wire wire32715;
wire wire32717;
wire wire32720;
wire wire32722;
wire wire32724;
wire wire32726;
wire wire32727;
wire wire32728;
wire wire32729;
wire wire32730;
wire wire32731;
wire wire32733;
wire wire32735;
wire wire32736;
wire wire32737;
wire wire32740;
wire wire32741;
wire wire32742;
wire wire32746;
wire wire32748;
wire wire32749;
wire wire32750;
wire wire32751;
wire wire32752;
wire wire32754;
wire wire32756;
wire wire32758;
wire wire32759;
wire wire32761;
wire wire32763;
wire wire32764;
wire wire32765;
wire wire32766;
wire wire32769;
wire wire32771;
wire wire32772;
wire wire32774;
wire wire32776;
wire wire32777;
wire wire32779;
wire wire32780;
wire wire32782;
wire wire32783;
wire wire32784;
wire wire32786;
wire wire32787;
wire wire32789;
wire wire32791;
wire wire32793;
wire wire32794;
wire wire32795;
wire wire32796;
wire wire32798;
wire wire32799;
wire wire32800;
wire wire32801;
wire wire32803;
wire wire32805;
wire wire32806;
wire wire32808;
wire wire32809;
wire wire32810;
wire wire32811;
wire wire32812;
wire wire32814;
wire wire32815;
wire wire32816;
wire wire32817;
wire wire32818;
wire wire32819;
wire wire32820;
wire wire32821;
wire wire32823;
wire wire32825;
wire wire32826;
wire wire32827;
wire wire32828;
wire wire32831;
wire wire32832;
wire wire32836;
wire wire32837;
wire wire32839;
wire wire32841;
wire wire32842;
wire wire32843;
wire wire32844;
wire wire32845;
wire wire32846;
wire wire32847;
wire wire32848;
wire wire32849;
wire wire32850;
wire wire32853;
wire wire32855;
wire wire32857;
wire wire32859;
wire wire32861;
wire wire32862;
wire wire32864;
wire wire32865;
wire wire32867;
wire wire32868;
wire wire32869;
wire wire32870;
wire wire32871;
wire wire32873;
wire wire32874;
wire wire32875;
wire wire32876;
wire wire32879;
wire wire32881;
wire wire32882;
wire wire32883;
wire wire32885;
wire wire32887;
wire wire32888;
wire wire32890;
wire wire32891;
wire wire32893;
wire wire32894;
wire wire32895;
wire wire32898;
wire wire32899;
wire wire32900;
wire wire32902;
wire wire32903;
wire wire32904;
wire wire32905;
wire wire32906;
wire wire32909;
wire wire32910;
wire wire32911;
wire wire32912;
wire wire32914;
wire wire32915;
wire wire32916;
wire wire32919;
wire wire32920;
wire wire32921;
wire wire32922;
wire wire32923;
wire wire32924;
wire wire32925;
wire wire32927;
wire wire32929;
wire wire32930;
wire wire32931;
wire wire32932;
wire wire32933;
wire wire32934;
wire wire32935;
wire wire32936;
wire wire32937;
wire wire32938;
wire wire32939;
wire wire32941;
wire wire32942;
wire wire32943;
wire wire32944;
wire wire32945;
wire wire32946;
wire wire32948;
wire wire32949;
wire wire32950;
wire wire32951;
wire wire32952;
wire wire32953;
wire wire32954;
wire wire32955;
wire wire32956;
wire wire32957;
wire wire32958;
wire wire32959;
wire wire32960;
wire wire32962;
wire wire32963;
wire wire32964;
wire wire32965;
wire wire32966;
wire wire32967;
wire wire32969;
wire wire32970;
wire wire32973;
wire wire32975;
wire wire32976;
wire wire32978;
wire wire32979;
wire wire32982;
wire wire32984;
wire wire32985;
wire wire32986;
wire wire32987;
wire wire32989;
wire wire32990;
wire wire32991;
wire wire32992;
wire wire32994;
wire wire32995;
wire wire32996;
wire wire32997;
wire wire32998;
wire wire33000;
wire wire33001;
wire wire33003;
wire wire33004;
wire wire33007;
wire wire33008;
wire wire33010;
wire wire33011;
wire wire33013;
wire wire33014;
wire wire33015;
wire wire33016;
wire wire33017;
wire wire33018;
wire wire33019;
wire wire33020;
wire wire33021;
wire wire33022;
wire wire33023;
wire wire33024;
wire wire33026;
wire wire33027;
wire wire33028;
wire wire33029;
wire wire33030;
wire wire33032;
wire wire33034;
wire wire33035;
wire wire33036;
wire wire33040;
wire wire33043;
wire wire33044;
wire wire33045;
wire wire33046;
wire wire33047;
wire wire33050;
wire wire33052;
wire wire33055;
wire wire33056;
wire wire33057;
wire wire33058;
wire wire33059;
wire wire33060;
wire wire33062;
wire wire33064;
wire wire33065;
wire wire33066;
wire wire33067;
wire wire33068;
wire wire33069;
wire wire33070;
wire wire33071;
wire wire33072;
wire wire33073;
wire wire33074;
wire wire33075;
wire wire33076;
wire wire33077;
wire wire33078;
wire wire33079;
wire wire33080;
wire wire33081;
wire wire33082;
wire wire33083;
wire wire33085;
wire wire33086;
wire wire33087;
wire wire33091;
wire wire33093;
wire wire33094;
wire wire33095;
wire wire33096;
wire wire33097;
wire wire33098;
wire wire33099;
wire wire33100;
wire wire33101;
wire wire33103;
wire wire33105;
wire wire33106;
wire wire33108;
wire wire33109;
wire wire33111;
wire wire33112;
wire wire33113;
wire wire33114;
wire wire33115;
wire wire33116;
wire wire33117;
wire wire33119;
wire wire33120;
wire wire33121;
wire wire33124;
wire wire33125;
wire wire33127;
wire wire33128;
wire wire33130;
wire wire33131;
wire wire33132;
wire wire33133;
wire wire33134;
wire wire33136;
wire wire33137;
wire wire33138;
wire wire33139;
wire wire33140;
wire wire33143;
wire wire33144;
wire wire33145;
wire wire33146;
wire wire33147;
wire wire33148;
wire wire33149;
wire wire33150;
wire wire33151;
wire wire33152;
wire wire33156;
wire wire33158;
wire wire33159;
wire wire33160;
wire wire33161;
wire wire33162;
wire wire33163;
wire wire33164;
wire wire33166;
wire wire33167;
wire wire33169;
wire wire33170;
wire wire33172;
wire wire33173;
wire wire33174;
wire wire33175;
wire wire33177;
wire wire33178;
wire wire33180;
wire wire33181;
wire wire33183;
wire wire33184;
wire wire33187;
wire wire33188;
wire wire33189;
wire wire33190;
wire wire33191;
wire wire33194;
wire wire33196;
wire wire33197;
wire wire33198;
wire wire33201;
wire wire33202;
wire wire33206;
wire wire33209;
wire wire33210;
wire wire33212;
wire wire33214;
wire wire33215;
wire wire33218;
wire wire33220;
wire wire33223;
wire wire33225;
wire wire33226;
wire wire33227;
wire wire33228;
wire wire33230;
wire wire33234;
wire wire33235;
wire wire33236;
wire wire33238;
wire wire33240;
wire wire33241;
wire wire33242;
wire wire33244;
wire wire33246;
wire wire33249;
wire wire33251;
wire wire33252;
wire wire33254;
wire wire33256;
wire wire33257;
wire wire33258;
wire wire33260;
wire wire33261;
wire wire33262;
wire wire33263;
wire wire33266;
wire wire33267;
wire wire33270;
wire wire33272;
wire wire33274;
wire wire33276;
wire wire33278;
wire wire33279;
wire wire33282;
wire wire33284;
wire wire33288;
wire wire33290;
wire wire33291;
wire wire33293;
wire wire33294;
wire wire33295;
wire wire33296;
wire wire33297;
wire wire33298;
wire wire33299;
wire wire33302;
wire wire33303;
wire wire33304;
wire wire33305;
wire wire33306;
wire wire33307;
wire wire33309;
wire wire33310;
wire wire33319;
wire wire33321;
wire wire33325;
wire wire33327;
wire wire33328;
wire wire33331;
wire wire33333;
wire wire33334;
wire wire33336;
wire wire33339;
wire wire33340;
wire wire33341;
wire wire33342;
wire wire33343;
wire wire33345;
wire wire33346;
wire wire33347;
wire wire33348;
wire wire33349;
wire wire33350;
wire wire33352;
wire wire33355;
wire wire33364;
wire wire33366;
wire wire33370;
wire wire33372;
wire wire33373;
wire wire33376;
wire wire33378;
wire wire33379;
wire wire33381;
wire wire33384;
wire wire33385;
wire wire33386;
wire wire33387;
wire wire33388;
wire wire33390;
wire wire33391;
wire wire33392;
wire wire33393;
wire wire33394;
wire wire33395;
wire wire33398;
wire wire33400;
wire wire33404;
wire wire33406;
wire wire33407;
wire wire33410;
wire wire33412;
wire wire33413;
wire wire33415;
wire wire33417;
wire wire33420;
wire wire33421;
wire wire33426;
wire wire33427;
wire wire33428;
wire wire33429;
wire wire33433;
wire wire33434;
wire wire33438;
wire wire33440;
wire wire33442;
wire wire33444;
wire wire33446;
wire wire33450;
wire wire33452;
wire wire33453;
wire wire33456;
wire wire33458;
wire wire33459;
wire wire33461;
wire wire33462;
wire wire33463;
wire wire33464;
wire wire33465;
wire wire33466;
wire wire33467;
wire wire33470;
wire wire33471;
wire wire33472;
wire wire33473;
wire wire33474;
wire wire33475;
wire wire33476;
wire wire33484;
wire wire33486;
wire wire33487;
wire wire33490;
wire wire33492;
wire wire33496;
wire wire33498;
wire wire33499;
wire wire33501;
wire wire33504;
wire wire33505;
wire wire33506;
wire wire33507;
wire wire33508;
wire wire33510;
wire wire33511;
wire wire33512;
wire wire33513;
wire wire33514;
wire wire33515;
wire wire33518;
wire wire33520;
wire wire33524;
wire wire33526;
wire wire33527;
wire wire33530;
wire wire33532;
wire wire33533;
wire wire33535;
wire wire33537;
wire wire33540;
wire wire33541;
wire wire33544;
wire wire33545;
wire wire33546;
wire wire33547;
wire wire33548;
wire wire33550;
wire wire33551;
wire wire33552;
wire wire33553;
wire wire33554;
wire wire33555;
wire wire33564;
wire wire33566;
wire wire33567;
wire wire33570;
wire wire33572;
wire wire33576;
wire wire33578;
wire wire33579;
wire wire33581;
wire wire33584;
wire wire33585;
wire wire33586;
wire wire33587;
wire wire33588;
wire wire33590;
wire wire33591;
wire wire33592;
wire wire33593;
wire wire33594;
wire wire33595;
wire wire33596;
wire wire33598;
wire wire33599;
wire wire33600;
wire wire33601;
wire wire33603;
wire wire33604;
wire wire33605;
wire wire33608;
wire wire33609;
wire wire33611;
wire wire33612;
wire wire33613;
wire wire33614;
wire wire33616;
wire wire33618;
wire wire33619;
wire wire33621;
wire wire33622;
wire wire33627;
wire wire33628;
wire wire33630;
wire wire33632;
wire wire33634;
wire wire33636;
wire wire33637;
wire wire33638;
wire wire33640;
wire wire33641;
wire wire33642;
wire wire33643;
wire wire33644;
wire wire33645;
wire wire33647;
wire wire33649;
wire wire33651;
wire wire33657;
wire wire33658;
wire wire33660;
wire wire33661;
wire wire33662;
wire wire33663;
wire wire33665;
wire wire33666;
wire wire33668;
wire wire33669;
wire wire33672;
wire wire33674;
wire wire33677;
wire wire33678;
wire wire33679;
wire wire33680;
wire wire33681;
wire wire33682;
wire wire33684;
wire wire33685;
wire wire33686;
wire wire33688;
wire wire33689;
wire wire33691;
wire wire33693;
wire wire33695;
wire wire33696;
wire wire33697;
wire wire33698;
wire wire33699;
wire wire33700;
wire wire33701;
wire wire33702;
wire wire33704;
wire wire33705;
wire wire33706;
wire wire33709;
wire wire33710;
wire wire33713;
wire wire33715;
wire wire33716;
wire wire33721;
wire wire33724;
wire wire33725;
wire wire33727;
wire wire33728;
wire wire33730;
wire wire33732;
wire wire33733;
wire wire33734;
wire wire33735;
wire wire33736;
wire wire33737;
wire wire33738;
wire wire33739;
wire wire33740;
wire wire33741;
wire wire33742;
wire wire33743;
wire wire33744;
wire wire33745;
wire wire33746;
wire wire33748;
wire wire33750;
wire wire33751;
wire wire33753;
wire wire33754;
wire wire33755;
wire wire33756;
wire wire33758;
wire wire33759;
wire wire33760;
wire wire33763;
wire wire33764;
wire wire33765;
wire wire33769;
wire wire33770;
wire wire33773;
wire wire33774;
wire wire33776;
wire wire33777;
wire wire33779;
wire wire33780;
wire wire33782;
wire wire33783;
wire wire33785;
wire wire33786;
wire wire33789;
wire wire33793;
wire wire33795;
wire wire33796;
wire wire33797;
wire wire33799;
wire wire33801;
wire wire33802;
wire wire33803;
wire wire33804;
wire wire33805;
wire wire33806;
wire wire33807;
wire wire33809;
wire wire33812;
wire wire33813;
wire wire33817;
wire wire33818;
wire wire33821;
wire wire33824;
wire wire33825;
wire wire33827;
wire wire33828;
wire wire33830;
wire wire33831;
wire wire33833;
wire wire33834;
wire wire33835;
wire wire33836;
wire wire33837;
wire wire33839;
wire wire33842;
wire wire33844;
wire wire33846;
wire wire33847;
wire wire33848;
wire wire33850;
wire wire33855;
wire wire33856;
wire wire33858;
wire wire33859;
wire wire33860;
wire wire33861;
wire wire33862;
wire wire33863;
wire wire33864;
wire wire33866;
wire wire33868;
wire wire33870;
wire wire33872;
wire wire33875;
wire wire33876;
wire wire33880;
wire wire33881;
wire wire33882;
wire wire33883;
wire wire33885;
wire wire33886;
wire wire33887;
wire wire33889;
wire wire33891;
wire wire33892;
wire wire33893;
wire wire33896;
wire wire33899;
wire wire33900;
wire wire33904;
wire wire33906;
wire wire33907;
wire wire33908;
wire wire33909;
wire wire33910;
wire wire33911;
wire wire33914;
wire wire33915;
wire wire33916;
wire wire33918;
wire wire33919;
wire wire33920;
wire wire33922;
wire wire33923;
wire wire33924;
wire wire33926;
wire wire33927;
wire wire33929;
wire wire33930;
wire wire33931;
wire wire33932;
wire wire33933;
wire wire33935;
wire wire33936;
wire wire33938;
wire wire33939;
wire wire33940;
wire wire33941;
wire wire33943;
wire wire33945;
wire wire33946;
wire wire33947;
wire wire33949;
wire wire33952;
wire wire33954;
wire wire33955;
wire wire33956;
wire wire33958;
wire wire33959;
wire wire33960;
wire wire33961;
wire wire33962;
wire wire33964;
wire wire33965;
wire wire33966;
wire wire33967;
wire wire33968;
wire wire33971;
wire wire33973;
wire wire33976;
wire wire33977;
wire wire33978;
wire wire33979;
wire wire33983;
wire wire33986;
wire wire33987;
wire wire33989;
wire wire33990;
wire wire33992;
wire wire33993;
wire wire33994;
wire wire33996;
wire wire33998;
wire wire34001;
wire wire34002;
wire wire34003;
wire wire34005;
wire wire34007;
wire wire34008;
wire wire34010;
wire wire34011;
wire wire34013;
wire wire34014;
wire wire34015;
wire wire34016;
wire wire34017;
wire wire34019;
wire wire34020;
wire wire34021;
wire wire34022;
wire wire34024;
wire wire34027;
wire wire34028;
wire wire34030;
wire wire34032;
wire wire34033;
wire wire34034;
wire wire34035;
wire wire34036;
wire wire34038;
wire wire34039;
wire wire34040;
wire wire34041;
wire wire34042;
wire wire34043;
wire wire34044;
wire wire34045;
wire wire34046;
wire wire34048;
wire wire34050;
wire wire34053;
wire wire34055;
wire wire34057;
wire wire34059;
wire wire34060;
wire wire34062;
wire wire34063;
wire wire34064;
wire wire34066;
wire wire34067;
wire wire34068;
wire wire34069;
wire wire34070;
wire wire34071;
wire wire34074;
wire wire34075;
wire wire34076;
wire wire34078;
wire wire34080;
wire wire34082;
wire wire34083;
wire wire34084;
wire wire34086;
wire wire34088;
wire wire34089;
wire wire34090;
wire wire34091;
wire wire34092;
wire wire34094;
wire wire34095;
wire wire34096;
wire wire34097;
wire wire34098;
wire wire34099;
wire wire34100;
wire wire34101;
wire wire34102;
wire wire34103;
wire wire34106;
wire wire34108;
wire wire34109;
wire wire34110;
wire wire34111;
wire wire34112;
wire wire34113;
wire wire34115;
wire wire34116;
wire wire34117;
wire wire34119;
wire wire34120;
wire wire34124;
wire wire34125;
wire wire34127;
wire wire34128;
wire wire34129;
wire wire34130;
wire wire34131;
wire wire34132;
wire wire34134;
wire wire34135;
wire wire34136;
wire wire34137;
wire wire34138;
wire wire34139;
wire wire34140;
wire wire34142;
wire wire34143;
wire wire34147;
wire wire34148;
wire wire34150;
wire wire34151;
wire wire34152;
wire wire34153;
wire wire34154;
wire wire34155;
wire wire34156;
wire wire34157;
wire wire34158;
wire wire34159;
wire wire34160;
wire wire34161;
wire wire34162;
wire wire34164;
wire wire34165;
wire wire34167;
wire wire34168;
wire wire34169;
wire wire34170;
wire wire34171;
wire wire34173;
wire wire34174;
wire wire34175;
wire wire34176;
wire wire34177;
wire wire34178;
wire wire34180;
wire wire34182;
wire wire34183;
wire wire34184;
wire wire34185;
wire wire34186;
wire wire34187;
wire wire34188;
wire wire34189;
wire wire34190;
wire wire34191;
wire wire34192;
wire wire34193;
wire wire34194;
wire wire34195;
wire wire34196;
wire wire34197;
wire wire34198;
wire wire34199;
wire wire34201;
wire wire34203;
wire wire34204;
wire wire34206;
wire wire34207;
wire wire34208;
wire wire34209;
wire wire34210;
wire wire34212;
wire wire34213;
wire wire34214;
wire wire34217;
wire wire34220;
wire wire34221;
wire wire34223;
wire wire34224;
wire wire34227;
wire wire34228;
wire wire34230;
wire wire34232;
wire wire34233;
wire wire34234;
wire wire34235;
wire wire34236;
wire wire34238;
wire wire34239;
wire wire34240;
wire wire34241;
wire wire34242;
wire wire34243;
wire wire34244;
wire wire34246;
wire wire34247;
wire wire34248;
wire wire34250;
wire wire34253;
wire wire34255;
wire wire34258;
wire wire34262;
wire wire34263;
wire wire34264;
wire wire34265;
wire wire34266;
wire wire34267;
wire wire34268;
wire wire34271;
wire wire34272;
wire wire34274;
wire wire34275;
wire wire34276;
wire wire34277;
wire wire34278;
wire wire34279;
wire wire34280;
wire wire34281;
wire wire34282;
wire wire34283;
wire wire34284;
wire wire34285;
wire wire34286;
wire wire34287;
wire wire34288;
wire wire34289;
wire wire34291;
wire wire34292;
wire wire34293;
wire wire34295;
wire wire34297;
wire wire34299;
wire wire34301;
wire wire34302;
wire wire34304;
wire wire34305;
wire wire34306;
wire wire34307;
wire wire34308;
wire wire34311;
wire wire34312;
wire wire34313;
wire wire34314;
wire wire34315;
wire wire34316;
wire wire34318;
wire wire34319;
wire wire34320;
wire wire34321;
wire wire34322;
wire wire34323;
wire wire34324;
wire wire34325;
wire wire34326;
wire wire34330;
wire wire34331;
wire wire34333;
wire wire34334;
wire wire34335;
wire wire34337;
wire wire34340;
wire wire34342;
wire wire34344;
wire wire34346;
wire wire34347;
wire wire34348;
wire wire34351;
wire wire34352;
wire wire34353;
wire wire34354;
wire wire34356;
wire wire34357;
wire wire34358;
wire wire34359;
wire wire34360;
wire wire34361;
wire wire34362;
wire wire34363;
wire wire34365;
wire wire34366;
wire wire34369;
wire wire34370;
wire wire34373;
wire wire34374;
wire wire34375;
wire wire34377;
wire wire34378;
wire wire34380;
wire wire34381;
wire wire34383;
wire wire34385;
wire wire34386;
wire wire34387;
wire wire34389;
wire wire34390;
wire wire34391;
wire wire34394;
wire wire34395;
wire wire34397;
wire wire34398;
wire wire34399;
wire wire34400;
wire wire34401;
wire wire34404;
wire wire34406;
wire wire34407;
wire wire34410;
wire wire34412;
wire wire34413;
wire wire34414;
wire wire34415;
wire wire34417;
wire wire34418;
wire wire34419;
wire wire34420;
wire wire34421;
wire wire34423;
wire wire34424;
wire wire34425;
wire wire34426;
wire wire34427;
wire wire34429;
wire wire34430;
wire wire34432;
wire wire34433;
wire wire34434;
wire wire34436;
wire wire34437;
wire wire34438;
wire wire34439;
wire wire34440;
wire wire34441;
wire wire34442;
wire wire34443;
wire wire34444;
wire wire34445;
wire wire34446;
wire wire34447;
wire wire34448;
wire wire34449;
wire wire34450;
wire wire34451;
wire wire34452;
wire wire34454;
wire wire34455;
wire wire34457;
wire wire34458;
wire wire34459;
wire wire34460;
wire wire34461;
wire wire34463;
wire wire34464;
wire wire34465;
wire wire34467;
wire wire34468;
wire wire34470;
wire wire34472;
wire wire34473;
wire wire34474;
wire wire34475;
wire wire34476;
wire wire34477;
wire wire34478;
wire wire34479;
wire wire34480;
wire wire34481;
wire wire34482;
wire wire34483;
wire wire34484;
wire wire34485;
wire wire34486;
wire wire34487;
wire wire34488;
wire wire34489;
wire wire34490;
wire wire34491;
wire wire34492;
wire wire34494;
wire wire34496;
wire wire34498;
wire wire34499;
wire wire34500;
wire wire34501;
wire wire34503;
wire wire34504;
wire wire34505;
wire wire34507;
wire wire34508;
wire wire34509;
wire wire34511;
wire wire34513;
wire wire34518;
wire wire34519;
wire wire34522;
wire wire34523;
wire wire34525;
wire wire34526;
wire wire34527;
wire wire34529;
wire wire34530;
wire wire34532;
wire wire34533;
wire wire34534;
wire wire34536;
wire wire34537;
wire wire34540;
wire wire34542;
wire wire34543;
wire wire34545;
wire wire34547;
wire wire34548;
wire wire34549;
wire wire34550;
wire wire34551;
wire wire34553;
wire wire34555;
wire wire34557;
wire wire34558;
wire wire34560;
wire wire34561;
wire wire34562;
wire wire34563;
wire wire34564;
wire wire34566;
wire wire34567;
wire wire34571;
wire wire34572;
wire wire34573;
wire wire34574;
wire wire34575;
wire wire34579;
wire wire34580;
wire wire34582;
wire wire34584;
wire wire34585;
wire wire34586;
wire wire34588;
wire wire34590;
wire wire34591;
wire wire34593;
wire wire34594;
wire wire34595;
wire wire34596;
wire wire34598;
wire wire34600;
wire wire34602;
wire wire34604;
wire wire34606;
wire wire34608;
wire wire34609;
wire wire34610;
wire wire34612;
wire wire34613;
wire wire34614;
wire wire34615;
wire wire34617;
wire wire34620;
wire wire34621;
wire wire34623;
wire wire34624;
wire wire34626;
wire wire34627;
wire wire34628;
wire wire34629;
wire wire34631;
wire wire34633;
wire wire34636;
wire wire34637;
wire wire34638;
wire wire34640;
wire wire34642;
wire wire34645;
wire wire34647;
wire wire34648;
wire wire34650;
wire wire34651;
wire wire34654;
wire wire34656;
wire wire34659;
wire wire34661;
wire wire34663;
wire wire34664;
wire wire34665;
wire wire34666;
wire wire34670;
wire wire34671;
wire wire34673;
wire wire34675;
wire wire34676;
wire wire34677;
wire wire34678;
wire wire34679;
wire wire34680;
wire wire34681;
wire wire34682;
wire wire34683;
wire wire34684;
wire wire34686;
wire wire34689;
wire wire34690;
wire wire34692;
wire wire34694;
wire wire34695;
wire wire34696;
wire wire34697;
wire wire34699;
wire wire34702;
wire wire34703;
wire wire34705;
wire wire34707;
wire wire34708;
wire wire34709;
wire wire34710;
wire wire34712;
wire wire34714;
wire wire34716;
wire wire34718;
wire wire34719;
wire wire34722;
wire wire34724;
wire wire34725;
wire wire34726;
wire wire34731;
wire wire34733;
wire wire34734;
wire wire34735;
wire wire34739;
wire wire34741;
wire wire34742;
wire wire34744;
wire wire34745;
wire wire34748;
wire wire34749;
wire wire34752;
wire wire34754;
wire wire34755;
wire wire34758;
wire wire34761;
wire wire34763;
wire wire34765;
wire wire34766;
wire wire34767;
wire wire34769;
wire wire34770;
wire wire34771;
wire wire34772;
wire wire34775;
wire wire34776;
wire wire34778;
wire wire34780;
wire wire34782;
wire wire34783;
wire wire34785;
wire wire34790;
wire wire34791;
wire wire34794;
wire wire34795;
wire wire34798;
wire wire34801;
wire wire34803;
wire wire34804;
wire wire34806;
wire wire34810;
wire wire34813;
wire wire34814;
wire wire34815;
wire wire34816;
wire wire34817;
wire wire34819;
wire wire34820;
wire wire34823;
wire wire34825;
wire wire34826;
wire wire34828;
wire wire34830;
wire wire34831;
wire wire34833;
wire wire34834;
wire wire34835;
wire wire34837;
wire wire34838;
wire wire34839;
wire wire34841;
wire wire34843;
wire wire34844;
wire wire34845;
wire wire34846;
wire wire34848;
wire wire34850;
wire wire34851;
wire wire34853;
wire wire34855;
wire wire34857;
wire wire34859;
wire wire34860;
wire wire34861;
wire wire34862;
wire wire34863;
wire wire34865;
wire wire34866;
wire wire34869;
wire wire34871;
wire wire34874;
wire wire34875;
wire wire34876;
wire wire34877;
wire wire34879;
wire wire34880;
wire wire34881;
wire wire34882;
wire wire34883;
wire wire34884;
wire wire34885;
wire wire34886;
wire wire34887;
wire wire34888;
wire wire34890;
wire wire34891;
wire wire34894;
wire wire34895;
wire wire34897;
wire wire34898;
wire wire34899;
wire wire34900;
wire wire34901;
wire wire34902;
wire wire34904;
wire wire34906;
wire wire34907;
wire wire34909;
wire wire34911;
wire wire34912;
wire wire34914;
wire wire34916;
wire wire34917;
wire wire34919;
wire wire34924;
wire wire34925;
wire wire34928;
wire wire34929;
wire wire34931;
wire wire34932;
wire wire34934;
wire wire34935;
wire wire34939;
wire wire34940;
wire wire34942;
wire wire34943;
wire wire34945;
wire wire34947;
wire wire34950;
wire wire34951;
wire wire34954;
wire wire34955;
wire wire34957;
wire wire34958;
wire wire34959;
wire wire34960;
wire wire34962;
wire wire34965;
wire wire34966;
wire wire34967;
wire wire34968;
wire wire34971;
wire wire34973;
wire wire34974;
wire wire34977;
wire wire34981;
wire wire34983;
wire wire34984;
wire wire34987;
wire wire34990;
wire wire34991;
wire wire34992;
wire wire34994;
wire wire34995;
wire wire34996;
wire wire34997;
wire wire34998;
wire wire34999;
wire wire35000;
wire wire35001;
wire wire35003;
wire wire35004;
wire wire35005;
wire wire35006;
wire wire35007;
wire wire35008;
wire wire35009;
wire wire35011;
wire wire35012;
wire wire35014;
wire wire35015;
wire wire35016;
wire wire35017;
wire wire35020;
wire wire35021;
wire wire35023;
wire wire35025;
wire wire35028;
wire wire35030;
wire wire35031;
wire wire35033;
wire wire35034;
wire wire35035;
wire wire35037;
wire wire35038;
wire wire35039;
wire wire35040;
wire wire35041;
wire wire35042;
wire wire35043;
wire wire35044;
wire wire35046;
wire wire35048;
wire wire35051;
wire wire35053;
wire wire35054;
wire wire35055;
wire wire35056;
wire wire35057;
wire wire35058;
wire wire35060;
wire wire35061;
wire wire35062;
wire wire35063;
wire wire35064;
wire wire35065;
wire wire35069;
wire wire35070;
wire wire35071;
wire wire35072;
wire wire35075;
wire wire35076;
wire wire35077;
wire wire35078;
wire wire35079;
wire wire35080;
wire wire35081;
wire wire35082;
wire wire35084;
wire wire35085;
wire wire35088;
wire wire35089;
wire wire35092;
wire wire35093;
wire wire35094;
wire wire35095;
wire wire35096;
wire wire35097;
wire wire35098;
wire wire35099;
wire wire35100;
wire wire35101;
wire wire35102;
wire wire35103;
wire wire35105;
wire wire35106;
wire wire35107;
wire wire35108;
wire wire35109;
wire wire35110;
wire wire35111;
wire wire35112;
wire wire35113;
wire wire35116;
wire wire35117;
wire wire35118;
wire wire35119;
wire wire35120;
wire wire35121;
wire wire35122;
wire wire35123;
wire wire35124;
wire wire35125;
wire wire35129;
wire wire35130;
wire wire35131;
wire wire35133;
wire wire35134;
wire wire35135;
wire wire35136;
wire wire35137;
wire wire35138;
wire wire35139;
wire wire35140;
wire wire35141;
wire wire35142;
wire wire35143;
wire wire35144;
wire wire35145;
wire wire35146;
wire wire35147;
wire wire35148;
wire wire35149;
wire wire35150;
wire wire35151;
wire wire35152;
wire wire35153;
wire wire35156;
wire wire35157;
wire wire35158;
wire wire35159;
wire wire35160;
wire wire35162;
wire wire35163;
wire wire35164;
wire wire35165;
wire wire35166;
wire wire35167;
wire wire35168;
wire wire35169;
wire wire35170;
wire wire35171;
wire wire35172;
wire wire35174;
wire wire35175;
wire wire35176;
wire wire35178;
wire wire35179;
wire wire35181;
wire wire35182;
wire wire35183;
wire wire35184;
wire wire35186;
wire wire35187;
wire wire35188;
wire wire35189;
wire wire35190;
wire wire35191;
wire wire35192;
wire wire35194;
wire wire35196;
wire wire35199;
wire wire35201;
wire wire35202;
wire wire35203;
wire wire35204;
wire wire35206;
wire wire35208;
wire wire35210;
wire wire35211;
wire wire35212;
wire wire35213;
wire wire35214;
wire wire35215;
wire wire35217;
wire wire35218;
wire wire35221;
wire wire35223;
wire wire35224;
wire wire35225;
wire wire35226;
wire wire35227;
wire wire35228;
wire wire35229;
wire wire35231;
wire wire35232;
wire wire35233;
wire wire35234;
wire wire35235;
wire wire35236;
wire wire35237;
wire wire35240;
wire wire35242;
wire wire35243;
wire wire35245;
wire wire35247;
wire wire35248;
wire wire35249;
wire wire35250;
wire wire35251;
wire wire35252;
wire wire35253;
wire wire35254;
wire wire35257;
wire wire35258;
wire wire35261;
wire wire35262;
wire wire35264;
wire wire35265;
wire wire35268;
wire wire35271;
wire wire35272;
wire wire35273;
wire wire35274;
wire wire35275;
wire wire35276;
wire wire35277;
wire wire35278;
wire wire35279;
wire wire35280;
wire wire35281;
wire wire35284;
wire wire35285;
wire wire35286;
wire wire35287;
wire wire35288;
wire wire35289;
wire wire35290;
wire wire35292;
wire wire35294;
wire wire35295;
wire wire35297;
wire wire35298;
wire wire35299;
wire wire35301;
wire wire35303;
wire wire35304;
wire wire35307;
wire wire35308;
wire wire35309;
wire wire35310;
wire wire35311;
wire wire35312;
wire wire35313;
wire wire35314;
wire wire35315;
wire wire35316;
wire wire35317;
wire wire35320;
wire wire35321;
wire wire35322;
wire wire35323;
wire wire35325;
wire wire35326;
wire wire35328;
wire wire35329;
wire wire35330;
wire wire35332;
wire wire35333;
wire wire35336;
wire wire35338;
wire wire35340;
wire wire35342;
wire wire35343;
wire wire35347;
wire wire35348;
wire wire35351;
wire wire35352;
wire wire35353;
wire wire35354;
wire wire35356;
wire wire35359;
wire wire35360;
wire wire35363;
wire wire35365;
wire wire35366;
wire wire35367;
wire wire35368;
wire wire35370;
wire wire35371;
wire wire35372;
wire wire35373;
wire wire35374;
wire wire35375;
wire wire35377;
wire wire35378;
wire wire35379;
wire wire35380;
wire wire35381;
wire wire35382;
wire wire35383;
wire wire35384;
wire wire35386;
wire wire35388;
wire wire35389;
wire wire35390;
wire wire35391;
wire wire35392;
wire wire35393;
wire wire35394;
wire wire35395;
wire wire35396;
wire wire35397;
wire wire35398;
wire wire35399;
wire wire35402;
wire wire35403;
wire wire35406;
wire wire35407;
wire wire35408;
wire wire35411;
wire wire35412;
wire wire35414;
wire wire35416;
wire wire35418;
wire wire35419;
wire wire35421;
wire wire35424;
wire wire35425;
wire wire35426;
wire wire35427;
wire wire35428;
wire wire35429;
wire wire35430;
wire wire35431;
wire wire35433;
wire wire35434;
wire wire35435;
wire wire35437;
wire wire35439;
wire wire35440;
wire wire35443;
wire wire35445;
wire wire35446;
wire wire35448;
wire wire35449;
wire wire35450;
wire wire35452;
wire wire35454;
wire wire35456;
wire wire35458;
wire wire35461;
wire wire35464;
wire wire35466;
wire wire35469;
wire wire35470;
wire wire35471;
wire wire35473;
wire wire35474;
wire wire35475;
wire wire35477;
wire wire35479;
wire wire35481;
wire wire35482;
wire wire35485;
wire wire35487;
wire wire35488;
wire wire35489;
wire wire35490;
wire wire35491;
wire wire35492;
wire wire35493;
wire wire35494;
wire wire35495;
wire wire35496;
wire wire35497;
wire wire35498;
wire wire35500;
wire wire35502;
wire wire35504;
wire wire35505;
wire wire35506;
wire wire35507;
wire wire35510;
wire wire35511;
wire wire35512;
wire wire35514;
wire wire35515;
wire wire35516;
wire wire35518;
wire wire35519;
wire wire35521;
wire wire35522;
wire wire35525;
wire wire35526;
wire wire35527;
wire wire35528;
wire wire35531;
wire wire35532;
wire wire35533;
wire wire35535;
wire wire35536;
wire wire35537;
wire wire35539;
wire wire35540;
wire wire35541;
wire wire35542;
wire wire35544;
wire wire35545;
wire wire35547;
wire wire35549;
wire wire35553;
wire wire35554;
wire wire35557;
wire wire35559;
wire wire35562;
wire wire35563;
wire wire35564;
wire wire35565;
wire wire35566;
wire wire35567;
wire wire35568;
wire wire35569;
wire wire35570;
wire wire35571;
wire wire35572;
wire wire35573;
wire wire35574;
wire wire35575;
wire wire35577;
wire wire35579;
wire wire35581;
wire wire35584;
wire wire35585;
wire wire35587;
wire wire35588;
wire wire35589;
wire wire35590;
wire wire35593;
wire wire35595;
wire wire35597;
wire wire35599;
wire wire35600;
wire wire35602;
wire wire35603;
wire wire35606;
wire wire35608;
wire wire35609;
wire wire35611;
wire wire35613;
wire wire35614;
wire wire35615;
wire wire35616;
wire wire35617;
wire wire35619;
wire wire35620;
wire wire35621;
wire wire35623;
wire wire35626;
wire wire35628;
wire wire35629;
wire wire35631;
wire wire35633;
wire wire35634;
wire wire35636;
wire wire35638;
wire wire35640;
wire wire35641;
wire wire35643;
wire wire35645;
wire wire35648;
wire wire35652;
wire wire35653;
wire wire35655;
wire wire35656;
wire wire35658;
wire wire35659;
wire wire35661;
wire wire35662;
wire wire35663;
wire wire35665;
wire wire35666;
wire wire35667;
wire wire35670;
wire wire35671;
wire wire35673;
wire wire35675;
wire wire35678;
wire wire35679;
wire wire35680;
wire wire35681;
wire wire35682;
wire wire35683;
wire wire35684;
wire wire35685;
wire wire35690;
wire wire35691;
wire wire35694;
wire wire35695;
reg ni39;

reg ni43;

reg ni42;

reg ni41;

reg ni40;

reg ni47;

reg ni46;

reg ni45;

reg ni44;

reg ni48;

reg ni38;

reg ni13;

reg ni2;

reg ni37;

reg ni14;

reg ni36;

reg ni11;

reg ni4;

reg ni35;

reg ni12;

reg ni3;

reg ni34;

reg ni9;

reg ni33;

reg ni10;

reg ni32;

reg ni7;

reg ni31;

reg ni8;

reg ni30;

reg ni5;

reg ni29;

reg ni6;

always  @(posedge pclk)
	ni39<=nv345;

 always  @(posedge pclk)
	ni43<=n_n13960;

 always  @(posedge pclk)
	ni42<=n_n13959;

 always  @(posedge pclk)
	ni41<=nv243;

 always  @(posedge pclk)
	ni40<=nv294;

 always  @(posedge pclk)
	ni47<=nv14;

 always  @(posedge pclk)
	ni46<=nv31;

 always  @(posedge pclk)
	ni45<=nv43;

 always  @(posedge pclk)
	ni44<=nv59;

 always  @(posedge pclk)
	ni48<=nv2;

 always  @(posedge pclk)
	ni38<=nv349;

 always  @(posedge pclk)
	ni13<=nv10068;

 always  @(posedge pclk)
	ni2<=n_n13958;

 always  @(posedge pclk)
	ni37<=nv437;

 always  @(posedge pclk)
	ni14<=nv10056;

 always  @(posedge pclk)
	ni36<=nv499;

 always  @(posedge pclk)
	ni11<=nv10091;

 always  @(posedge pclk)
	ni4<=nv10316;

 always  @(posedge pclk)
	ni35<=nv550;

 always  @(posedge pclk)
	ni12<=nv10082;

 always  @(posedge pclk)
	ni3<=n_n13895;

 always  @(posedge pclk)
	ni34<=nv601;

 always  @(posedge pclk)
	ni9<=nv10112;

 always  @(posedge pclk)
	ni33<=nv2153;

 always  @(posedge pclk)
	ni10<=nv10099;

 always  @(posedge pclk)
	ni32<=nv3888;

 always  @(posedge pclk)
	ni7<=nv10135;

 always  @(posedge pclk)
	ni31<=nv6425;

 always  @(posedge pclk)
	ni8<=nv10126;

 always  @(posedge pclk)
	ni30<=nv6437;

 always  @(posedge pclk)
	ni5<=nv10247;

 always  @(posedge pclk)
	ni29<=nv8909;

 always  @(posedge pclk)
	ni6<=nv10143;

 assign p__cmx0ad_22 = ( pi63  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_7 = ( pi239  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_23 = ( pi64  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_24 = ( pi65  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_5 = ( pi237  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_25 = ( pi66  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_6 = ( pi238  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmnxcp_0 = ( wire35670 ) | ( (~ n_n424)  &  wire35662 ) | ( (~ n_n424)  &  wire35666 ) ;
 assign p__cmx0ad_15 = ( ni9  &  ni10  &  wire1289  &  wire35671 ) ;
 assign p__cmx1ad_16 = ( pi240  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_27 = ( pi251  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmnxcp_1 = ( (~ ni2)  &  (~ wire367)  &  (~ wire35690)  &  (~ wire35691) ) ;
 assign p__cmx0ad_14 = ( (~ pi23)  &  pi24  &  nv10130  &  wire1289 ) | ( pi23  &  (~ pi24)  &  nv10130  &  wire1289 ) ;
 assign p__cmx1ad_17 = ( pi241  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_26 = ( pi250  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_13 = ( pi23  &  nv10130  &  wire1289 ) | ( pi24  &  nv10130  &  wire1289 ) ;
 assign p__cmx0ad_20 = ( pi61  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_31 = ( pi72  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_9 = ( (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_18 = ( pi242  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_29 = ( pi253  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_12 = ( (~ pi24)  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_21 = ( pi62  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_30 = ( pi71  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_19 = ( pi243  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_28 = ( pi252  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_9 = ( ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_0 = ( pi232  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmndst1p0 = ( ni43  &  (~ ni42)  &  (~ ni32) ) | ( ni43  &  (~ ni42)  &  (~ ni30) ) ;
 assign p__cmx0ad_6 = ( pi55  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_7 = ( pi56  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_3 = ( pi235  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmndst0p0 = ( ni38  &  (~ ni37)  &  ni32 ) | ( ni38  &  (~ ni37)  &  (~ ni30) ) ;
 assign p__cmx1ad_4 = ( pi236  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_1 = ( pi233  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_2 = ( pi234  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_0 = ( pi49  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_1 = ( pi50  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_4 = ( pi53  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_5 = ( pi54  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmxig_0 = ( (~ ni33)  &  ni29 ) ;
 assign p__cmx0ad_2 = ( pi51  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmxig_1 = ( ni33  &  ni29 ) ;
 assign p__cmx0ad_3 = ( pi52  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx0ad_19 = ( pi60  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_12 = ( (~ pi27)  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx1ad_23 = ( pi247  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmxir_0 = ( wire168 ) | ( wire1323  &  wire35694 ) ;
 assign p__cmx0ad_18 = ( pi59  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_13 = ( (~ ni2)  &  (~ ni3)  &  (~ wire290)  &  wire156 ) ;
 assign p__cmx1ad_22 = ( pi246  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmxir_1 = ( (~ wire289)  &  wire35695 ) ;
 assign p__cmx0ad_17 = ( pi58  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_14 = ( (~ pi27)  &  pi26  &  n_n13895  &  (~ wire290) ) | ( pi27  &  (~ pi26)  &  n_n13895  &  (~ wire290) ) ;
 assign p__cmx1ad_25 = ( pi249  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_16 = ( pi57  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_15 = ( pi27  &  pi26  &  n_n13895  &  (~ wire290) ) ;
 assign p__cmx1ad_24 = ( pi248  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_26 = ( pi67  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_30 = ( pi254  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_27 = ( pi68  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_31 = ( pi255  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_28 = ( pi69  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_21 = ( pi245  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign p__cmx0ad_29 = ( pi70  &  ni9  &  ni10  &  wire1289 ) ;
 assign p__cmx1ad_20 = ( pi244  &  (~ ni2)  &  (~ ni3)  &  (~ wire290) ) ;
 assign nv345 = ( wire7193 ) | ( wire7194 ) ;
 assign n_n13960 = ( wire28765 ) | ( wire28766 ) | ( wire28770 ) ;
 assign n_n13959 = ( (~ wire7090)  &  (~ wire7095)  &  (~ wire28905)  &  (~ wire28906) ) ;
 assign nv243 = ( wire28944 ) | ( wire28945 ) | ( wire28946 ) ;
 assign nv294 = ( wire7055 ) | ( wire7056 ) | ( wire28986 ) | ( wire28987 ) ;
 assign nv14 = ( wire7042 ) | ( wire7043 ) | ( wire28991 ) ;
 assign nv31 = ( wire7035 ) | ( wire28995 ) | ( wire1002  &  wire1085 ) ;
 assign nv43 = ( wire1002 ) | ( wire7030 ) | ( wire7031 ) | ( wire7032 ) ;
 assign nv59 = ( wire7028 ) | ( wire7029 ) ;
 assign nv2 = ( wire29003 ) | ( pi20  &  (~ ni47)  &  wire7044 ) ;
 assign nv349 = ( wire6997 ) | ( wire29081 ) | ( wire29082 ) | ( wire29086 ) ;
 assign nv10068 = ( wire29102 ) | ( (~ n_n1063)  &  wire1343 ) | ( (~ n_n1063)  &  wire29100 ) ;
 assign n_n13958 = ( (~ ni2)  &  ni3 ) ;
 assign nv437 = ( wire6946 ) | ( wire6951 ) | ( wire29131 ) | ( wire29136 ) ;
 assign nv10056 = ( wire6935 ) | ( wire6936 ) | ( wire29149 ) ;
 assign nv499 = ( wire6923 ) | ( wire6925 ) | ( wire29171 ) | ( wire29176 ) ;
 assign nv10091 = ( wire6973 ) | ( wire6975 ) | ( wire29092 ) | ( wire29094 ) ;
 assign nv10316 = ( ni2  &  ni4 ) | ( (~ ni2)  &  (~ wire29393)  &  (~ wire29394) ) ;
 assign nv550 = ( wire29430 ) | ( wire29431 ) | ( wire29437 ) | ( wire29438 ) ;
 assign nv10082 = ( wire29447 ) | ( n_n450  &  wire29441 ) | ( n_n450  &  wire29444 ) ;
 assign n_n13895 = ( (~ ni2)  &  (~ ni3) ) ;
 assign nv601 = ( wire30336 ) | ( n_n13895  &  (~ wire265)  &  n_n13077 ) ;
 assign nv10112 = ( wire30359 ) | ( wire30360 ) | ( wire30364 ) ;
 assign nv2153 = ( wire31159 ) | ( wire31040  &  wire31042 ) | ( wire31041  &  wire31042 ) ;
 assign nv10099 = ( wire31169 ) | ( wire1323  &  (~ wire31166)  &  (~ wire31167) ) ;
 assign nv3888 = ( wire3516 ) | ( wire3520 ) | ( wire3521 ) | ( wire33246 ) ;
 assign nv10135 = ( wire3512 ) | ( wire3514 ) | ( wire331  &  wire33249 ) ;
 assign nv6425 = ( wire33256 ) | ( nv6428  &  wire33251 ) | ( nv6428  &  wire33252 ) ;
 assign nv10126 = ( wire33262 ) | ( wire33263 ) ;
 assign nv6437 = ( wire34973 ) | ( wire34965  &  wire34967 ) | ( wire34966  &  wire34967 ) ;
 assign nv10247 = ( ni2  &  ni5 ) | ( (~ ni2)  &  (~ nv10248) ) ;
 assign nv8909 = ( wire518 ) | ( wire520 ) | ( wire35621 ) ;
 assign nv10143 = ( ni2  &  ni6 ) | ( (~ ni2)  &  (~ wire515)  &  (~ wire35634) ) ;
 assign nv10727 = ( ni33  &  ni31 ) ;
 assign nv8608 = ( ni31  &  ni30 ) ;
 assign n_n424 = ( wire445 ) | ( wire469 ) | ( wire470 ) | ( wire35648 ) ;
 assign wire425 = ( ni2 ) | ( (~ ni3) ) | ( (~ ni6) ) ;
 assign wire830 = ( (~ ni2)  &  ni4  &  ni3 ) ;
 assign wire856 = ( (~ ni31) ) | ( ni31  &  ni30 ) ;
 assign wire161 = ( pi23 ) | ( pi24 ) ;
 assign wire290 = ( (~ ni13) ) | ( (~ ni14) ) | ( ni11 ) | ( ni12 ) ;
 assign nv10130 = ( ni9  &  ni10 ) ;
 assign wire1289 = ( (~ ni2)  &  (~ ni3)  &  (~ ni7)  &  (~ ni8) ) ;
 assign n_n9245 = ( ni32  &  ni30 ) ;
 assign n_n13643 = ( (~ ni43)  &  (~ ni42) ) ;
 assign n_n13271 = ( ni38  &  (~ ni37) ) ;
 assign wire265 = ( ni9 ) | ( ni7 ) | ( ni8 ) ;
 assign wire1323 = ( (~ ni2)  &  (~ ni3)  &  (~ ni10) ) ;
 assign wire156 = ( pi27 ) | ( pi26 ) ;
 assign wire289 = ( ni13 ) | ( (~ ni14) ) | ( ni11 ) | ( ni12 ) ;
 assign n_n13390 = ( ni33  &  (~ ni32) ) ;
 assign wire711 = ( ni32 ) | ( ni31 ) | ( (~ ni32)  &  (~ ni30) ) ;
 assign nv69 = ( ni43  &  ni42  &  ni41 ) | ( ni43  &  ni42  &  (~ ni41) ) | ( ni43  &  (~ ni42)  &  (~ ni41)  &  ni44 ) ;
 assign nv78 = ( ni43  &  ni42  &  ni41 ) | ( ni43  &  ni42  &  (~ ni41) ) | ( ni43  &  (~ ni41)  &  (~ ni44) ) ;
 assign wire326 = ( (~ pi19)  &  (~ pi20) ) ;
 assign wire302 = ( (~ pi17)  &  (~ pi16) ) ;
 assign wire282 = ( (~ pi19)  &  pi20 ) ;
 assign wire514 = ( (~ ni43) ) | ( (~ ni42)  &  ni41 ) ;
 assign n_n13789 = ( wire7180 ) | ( wire28715 ) | ( wire28716 ) | ( wire28718 ) ;
 assign n_n13786 = ( wire7170 ) | ( wire7173 ) | ( wire28731 ) ;
 assign wire829 = ( (~ ni40)  &  (~ ni32) ) | ( (~ ni40)  &  (~ ni30) ) ;
 assign wire839 = ( ni40  &  (~ ni32) ) | ( ni40  &  (~ ni30) ) ;
 assign wire911 = ( ni32  &  ni31  &  ni30 ) ;
 assign wire1153 = ( (~ ni32) ) | ( (~ ni30) ) | ( ni31  &  ni30 ) ;
 assign nv251 = ( ni41  &  wire290 ) | ( ni41  &  wire638 ) | ( pi27  &  (~ wire290)  &  (~ wire638) ) ;
 assign n_n434 = ( ni41  &  ni33  &  ni32 ) ;
 assign nv6428 = ( ni31 ) | ( (~ ni32)  &  (~ ni30) ) ;
 assign wire466 = ( (~ ni32) ) | ( ni31 ) | ( (~ ni30) ) ;
 assign wire594 = ( ni9  &  ni10  &  (~ wire290) ) ;
 assign wire638 = ( (~ ni33) ) | ( (~ ni32) ) | ( ni31 ) | ( (~ ni30) ) ;
 assign wire792 = ( (~ ni9) ) | ( ni7 ) | ( ni8 ) ;
 assign wire988 = ( (~ ni32) ) | ( ni31 ) | ( (~ ni30) ) | ( ni33  &  ni32 ) ;
 assign wire1026 = ( (~ ni2)  &  (~ ni3)  &  (~ wire281)  &  (~ wire202) ) ;
 assign wire1122 = ( pi27  &  pi24 ) ;
 assign wire1299 = ( pi27  &  (~ pi24) ) ;
 assign wire462 = ( (~ pi26) ) | ( (~ pi23) ) ;
 assign wire1002 = ( (~ pi21)  &  ni32 ) | ( (~ pi21)  &  (~ ni31) ) | ( (~ pi21)  &  ni30 ) ;
 assign wire1085 = ( ni46  &  ni45 ) ;
 assign nv10169 = ( (~ ni30) ) | ( ni31  &  ni30 ) ;
 assign wire218 = ( (~ ni32) ) | ( (~ ni31) ) | ( ni30 ) ;
 assign nv354 = ( ni38  &  ni37 ) | ( ni39  &  ni38  &  (~ ni36) ) ;
 assign nv406 = ( (~ ni39)  &  ni38 ) | ( ni38  &  ni36 ) | ( ni38  &  ni37  &  (~ ni36) ) ;
 assign nv363 = ( (~ ni39)  &  ni38  &  ni37 ) | ( ni38  &  ni37  &  ni36 ) | ( ni38  &  ni37  &  (~ ni36) ) | ( (~ ni39)  &  ni38  &  (~ ni37)  &  (~ ni36) ) ;
 assign nv401 = ( ni39  &  ni38 ) | ( ni38  &  ni37 ) | ( ni38  &  ni36 ) ;
 assign wire191 = ( (~ pi17)  &  pi19 ) ;
 assign wire228 = ( (~ pi17)  &  (~ pi19)  &  pi20 ) ;
 assign wire260 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20) ) ;
 assign wire299 = ( pi17  &  pi19 ) ;
 assign wire396 = ( (~ ni35)  &  ni32 ) | ( (~ ni35)  &  (~ ni31) ) | ( (~ ni35)  &  (~ ni30) ) ;
 assign wire412 = ( ni37  &  ni36  &  ni32 ) | ( ni37  &  ni36  &  (~ ni30) ) ;
 assign wire439 = ( ni35  &  ni32 ) | ( ni35  &  (~ ni31) ) | ( ni35  &  (~ ni30) ) ;
 assign wire458 = ( pi17  &  (~ pi19)  &  pi20 ) ;
 assign wire1086 = ( (~ ni32)  &  (~ ni31)  &  ni30 ) ;
 assign n_n1063 = ( wire6966 ) | ( wire6968 ) | ( wire29098 ) ;
 assign wire1343 = ( ni13  &  (~ ni14) ) ;
 assign nv444 = ( ni39  &  ni43  &  ni44 ) | ( ni39  &  ni42  &  ni44 ) | ( (~ ni39)  &  ni43  &  (~ ni44) ) | ( (~ ni39)  &  ni42  &  (~ ni44) ) ;
 assign wire176 = ( ni36 ) | ( (~ ni35) ) ;
 assign wire262 = ( (~ pi18) ) | ( pi17 ) ;
 assign wire319 = ( ni35  &  ni32 ) | ( ni35  &  (~ ni30) ) ;
 assign wire890 = ( (~ pi18) ) | ( pi17 ) | ( pi20 ) ;
 assign wire177 = ( ni36 ) | ( ni35 ) ;
 assign wire229 = ( ni39 ) | ( ni36 ) ;
 assign wire382 = ( (~ ni38)  &  (~ ni36) ) ;
 assign nv10086 = ( ni13  &  ni14 ) ;
 assign n_n450 = ( wire948 ) | ( wire6940 ) | ( wire29139 ) ;
 assign nv539 = ( ni36  &  ni32 ) ;
 assign wire186 = ( ni11 ) | ( ni12 ) ;
 assign wire630 = ( (~ ni13) ) | ( ni11 ) | ( ni12 ) ;
 assign wire1105 = ( ni9  &  ni10  &  wire1289  &  (~ wire281) ) ;
 assign wire1252 = ( (~ ni33) ) | ( ni32 ) | ( wire290 ) | ( nv6428 ) ;
 assign wire155 = ( pi27 ) | ( (~ pi26) ) ;
 assign wire190 = ( (~ ni11)  &  ni12 ) ;
 assign nv590 = ( ni35  &  ni32 ) ;
 assign n_n11282 = ( ni33  &  ni30 ) ;
 assign nv7447 = ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign n_n13096 = ( wire6789 ) | ( pi26  &  ni35 ) ;
 assign nv2066 = ( wire30327 ) | ( (~ wire289)  &  wire30307 ) | ( (~ wire289)  &  wire30308 ) ;
 assign n_n11570 = ( wire6185 ) | ( wire6190 ) | ( wire29880 ) | ( wire29884 ) ;
 assign n_n13077 = ( wire30236 ) | ( wire6124  &  wire30217 ) | ( wire30216  &  wire30217 ) ;
 assign wire175 = ( ni13 ) | ( (~ ni14) ) | ( ni12 ) ;
 assign wire264 = ( ni11  &  (~ ni9)  &  ni10 ) ;
 assign wire692 = ( pi15  &  (~ wire289) ) ;
 assign wire708 = ( (~ pi15)  &  (~ wire289) ) ;
 assign n_n429 = ( wire5961 ) | ( (~ pi23)  &  ni7 ) | ( pi24  &  ni7 ) ;
 assign wire510 = ( (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire636 = ( (~ ni10) ) | ( ni8 ) | ( ni9  &  ni10 ) ;
 assign nv3311 = ( wire751 ) | ( (~ n_n12619)  &  wire240 ) | ( (~ n_n12619)  &  wire5906 ) ;
 assign nv3377 = ( wire304 ) | ( wire240  &  wire252 ) | ( wire252  &  wire5871 ) ;
 assign nv3280 = ( wire304 ) | ( wire240  &  wire252 ) | ( wire252  &  wire5861 ) ;
 assign nv3369 = ( wire304 ) | ( wire240  &  wire252 ) | ( wire252  &  wire5845 ) ;
 assign n_n9587 = ( wire30426 ) | ( wire252  &  wire5788 ) | ( wire252  &  wire30425 ) ;
 assign nv3273 = ( wire304 ) | ( wire240  &  wire252 ) | ( wire252  &  wire5770 ) ;
 assign n_n9650 = ( wire5079 ) | ( wire30515 ) | ( wire302  &  n_n9647 ) ;
 assign wire158 = ( pi17  &  (~ pi16) ) ;
 assign wire178 = ( (~ pi19)  &  pi21  &  pi22  &  (~ pi20) ) ;
 assign wire180 = ( (~ pi19)  &  pi21  &  pi22  &  pi20 ) ;
 assign wire294 = ( pi20  &  (~ pi16)  &  wire153 ) ;
 assign wire325 = ( (~ pi20)  &  (~ pi16)  &  wire153 ) ;
 assign wire395 = ( (~ pi17)  &  pi16  &  pi15 ) ;
 assign wire399 = ( ni7 ) | ( ni8 ) | ( ni9  &  ni10 ) ;
 assign wire403 = ( pi17  &  pi16  &  pi15 ) ;
 assign wire416 = ( pi17  &  pi16  &  pi15  &  wire152 ) ;
 assign wire438 = ( (~ pi19)  &  pi20  &  wire162 ) | ( (~ pi19)  &  (~ pi20)  &  wire159 ) ;
 assign wire631 = ( ni13 ) | ( ni11 ) | ( ni12 ) ;
 assign wire762 = ( wire30882 ) | ( wire30883 ) | ( pi15  &  wire723 ) ;
 assign wire1336 = ( pi20  &  wire485  &  wire162 ) | ( (~ pi20)  &  wire485  &  wire159 ) ;
 assign n_n8104 = ( wire4478 ) | ( wire4479 ) | ( wire4480 ) | ( wire32134 ) ;
 assign wire281 = ( ni4 ) | ( ni5 ) | ( ni6 ) ;
 assign wire509 = ( (~ ni9)  &  ni10 ) ;
 assign wire331 = ( (~ ni7)  &  ni8 ) ;
 assign wire1165 = ( (~ ni9) ) | ( (~ ni10) ) | ( (~ ni8) ) ;
 assign nv633 = ( ni47 ) | ( ni45 ) | ( (~ ni43)  &  ni42 ) ;
 assign wire150 = ( (~ pi21) ) | ( (~ pi22) ) ;
 assign wire172 = ( ni38 ) | ( (~ ni37) ) ;
 assign nv6450 = ( wire3047 ) | ( wire3049 ) | ( wire33769 ) | ( wire33770 ) ;
 assign nv10248 = ( wire2116 ) | ( wire2117 ) | ( wire2118 ) | ( wire34987 ) ;
 assign n_n13961 =((~ pi18) & pi18);
 assign wire160 = ( (~ pi23) ) | ( pi24 ) ;
 assign wire202 = ( ni7 ) | ( ni8 ) ;
 assign wire389 = ( (~ ni14) ) | ( ni12 ) ;
 assign wire478 = ( (~ ni31) ) | ( (~ ni6) ) ;
 assign wire725 = ( ni4 ) | ( (~ ni5) ) ;
 assign wire930 = ( (~ ni36) ) | ( (~ ni33) ) | ( ni32 ) ;
 assign wire936 = ( (~ ni33) ) | ( (~ ni31) ) | ( ni30 ) ;
 assign wire1029 = ( (~ ni4)  &  (~ ni6) ) ;
 assign nv121 = ( ni43  &  ni42 ) | ( ni43  &  ni41 ) | ( ni43  &  (~ ni44) ) ;
 assign nv158 = ( ni43  &  ni42 ) | ( (~ ni43)  &  (~ ni42) ) | ( (~ ni42)  &  (~ ni41) ) ;
 assign nv163 = ( (~ ni42) ) | ( ni43  &  ni44 ) ;
 assign n_n13541 = ( (~ ni42)  &  ni41 ) | ( ni43  &  ni41  &  ni44 ) ;
 assign n_n13646 = ( (~ ni43)  &  (~ ni42)  &  ni41 ) | ( ni43  &  ni42  &  ni41  &  ni44 ) ;
 assign n_n13755 = ( ni43  &  ni42  &  (~ ni40) ) | ( ni43  &  (~ ni41)  &  (~ ni40) ) ;
 assign n_n13600 = ( (~ ni41)  &  (~ ni40)  &  nv163 ) | ( ni41  &  (~ ni40)  &  nv158  &  nv163 ) ;
 assign wire490 = ( ni39  &  ni44 ) | ( (~ ni39)  &  (~ ni44) ) ;
 assign n_n13566 = ( ni43  &  ni42  &  (~ ni41) ) | ( (~ ni43)  &  (~ ni42)  &  (~ ni41) ) | ( (~ ni42)  &  (~ ni41)  &  ni44 ) ;
 assign nv116 = ( ni43  &  ni41 ) | ( ni43  &  ni42  &  (~ ni41) ) | ( ni43  &  (~ ni42)  &  ni44 ) ;
 assign wire426 = ( ni42 ) | ( (~ ni41) ) ;
 assign wire851 = ( wire7134 ) | ( (~ ni39)  &  (~ ni40)  &  (~ n_n13600) ) ;
 assign n_n13546 = ( ni43  &  ni42  &  (~ ni41) ) | ( (~ ni43)  &  (~ ni42)  &  (~ ni41) ) | ( ni43  &  (~ ni41)  &  (~ ni44) ) ;
 assign nv212 = ( ni39  &  (~ ni43)  &  ni42 ) | ( (~ ni39)  &  (~ ni43)  &  ni42 ) | ( ni39  &  ni42  &  ni44 ) | ( (~ ni39)  &  ni42  &  (~ ni44) ) ;
 assign wire222 = ( ni38 ) | ( ni37 ) ;
 assign wire419 = ( ni43 ) | ( (~ ni42) ) ;
 assign wire318 = ( ni31  &  ni30 ) | ( ni30  &  (~ wire490) ) | ( ni30  &  (~ wire28771) ) ;
 assign wire1037 = ( nv8608  &  n_n9245 ) | ( n_n9245  &  (~ wire490) ) | ( n_n9245  &  (~ wire28771) ) ;
 assign nv222 = ( nv212 ) | ( (~ n_n13755)  &  (~ n_n13566)  &  n_n13546 ) ;
 assign wire342 = ( ni39 ) | ( ni37 ) | ( ni36 ) ;
 assign wire231 = ( (~ ni39) ) | ( ni36 ) ;
 assign wire768 = ( ni33 ) | ( ni32 ) | ( ni31 ) | ( (~ ni32)  &  (~ ni30) ) ;
 assign nv667 = ( ni42 ) | ( nv669 ) | ( (~ ni42)  &  ni41 ) ;
 assign wire441 = ( ni41 ) | ( wire6727 ) | ( ni42  &  (~ ni41) ) | ( (~ ni41)  &  nv669 ) ;
 assign wire269 = ( ni39  &  (~ ni36) ) | ( ni38  &  (~ ni36) ) ;
 assign wire604 = ( wire357 ) | ( (~ ni38)  &  (~ wire229)  &  nv633 ) ;
 assign wire1032 = ( ni38  &  ni36 ) | ( ni38  &  (~ ni35) ) ;
 assign wire320 = ( (~ ni38)  &  ni37 ) | ( (~ ni38)  &  (~ ni37)  &  nv633 ) ;
 assign wire1097 = ( (~ ni38)  &  ni37  &  wire176 ) | ( (~ ni38)  &  (~ ni37)  &  wire176  &  nv633 ) ;
 assign nv903 = ( wire1097 ) | ( wire6682 ) | ( wire6683 ) ;
 assign nv952 = ( n_n12696 ) | ( wire1060 ) | ( wire222  &  wire29518 ) ;
 assign wire157 = ( ni31 ) | ( ni32  &  (~ ni31) ) | ( (~ ni31)  &  ni30 ) ;
 assign nv963 = ( wire1097 ) | ( wire6580 ) | ( wire6581 ) ;
 assign nv959 = ( ni34 ) | ( (~ wire157)  &  (~ wire6581)  &  (~ wire29504) ) ;
 assign nv758 = ( nv669 ) | ( ni42  &  (~ nv669) ) | ( (~ ni41)  &  (~ nv669)  &  wire6766 ) ;
 assign wire388 = ( ni42 ) | ( ni47 ) | ( ni45 ) | ( ni43  &  (~ ni47) ) ;
 assign wire292 = ( (~ ni39)  &  (~ ni36) ) | ( ni38  &  (~ ni36) ) ;
 assign wire357 = ( (~ ni38)  &  ni37  &  (~ ni36) ) ;
 assign wire500 = ( wire357 ) | ( (~ ni38)  &  nv633  &  (~ wire231) ) ;
 assign n_n12655 = ( (~ pi25)  &  ni34 ) ;
 assign nv772 = ( wire6727 ) | ( ni42  &  ni41 ) | ( ni42  &  (~ ni41) ) | ( ni41  &  nv669 ) | ( (~ ni41)  &  nv669 ) ;
 assign n_n11316 = ( (~ pi21)  &  ni34 ) ;
 assign nv699 = ( ni34 ) | ( (~ wire157)  &  (~ wire6742)  &  (~ wire29648) ) ;
 assign wire379 = ( pi21  &  wire224 ) ;
 assign wire380 = ( pi21  &  pi22  &  wire312 ) ;
 assign wire1332 = ( ni34  &  wire6742 ) | ( ni34  &  wire6743 ) | ( ni34  &  wire29647 ) ;
 assign nv717 = ( ni34 ) | ( (~ wire157)  &  (~ wire6703)  &  (~ wire29653) ) ;
 assign wire184 = ( ni34  &  ni31 ) | ( ni34  &  ni33  &  ni29 ) ;
 assign wire1092 = ( ni34  &  wire6701 ) | ( ni34  &  wire6703 ) | ( ni34  &  wire29652 ) ;
 assign nv1117 = ( wire184 ) | ( (~ nv6428)  &  nv717 ) | ( nv717  &  nv721 ) ;
 assign nv735 = ( ni34 ) | ( (~ wire157)  &  (~ wire6691)  &  (~ wire29623) ) ;
 assign wire1131 = ( ni34  &  wire436 ) | ( ni34  &  wire6691 ) | ( ni34  &  wire6692 ) ;
 assign nv1138 = ( wire184 ) | ( (~ nv6428)  &  nv735 ) | ( nv735  &  nv739 ) ;
 assign nv739 = ( wire436 ) | ( wire6691 ) | ( wire6692 ) ;
 assign nv721 = ( wire436 ) | ( wire6701 ) | ( wire6702 ) | ( wire6703 ) ;
 assign nv1096 = ( wire184 ) | ( (~ nv6428)  &  nv699 ) | ( nv699  &  nv703 ) ;
 assign nv703 = ( wire436 ) | ( wire6741 ) | ( wire6742 ) | ( wire6743 ) ;
 assign wire459 = ( (~ ni34) ) | ( pi22  &  pi25 ) ;
 assign wire225 = ( (~ ni34)  &  (~ nv6428) ) | ( pi22  &  pi25  &  (~ ni34) ) | ( pi22  &  pi25  &  (~ nv6428) ) ;
 assign wire152 = ( pi19  &  pi21  &  pi22 ) ;
 assign wire272 = ( pi17  &  pi19  &  pi21  &  pi22 ) ;
 assign wire483 = ( pi22  &  pi25  &  wire184 ) ;
 assign wire271 = ( (~ pi21)  &  ni34 ) | ( (~ pi22)  &  ni34 ) ;
 assign wire211 = ( pi21  &  pi20 ) ;
 assign wire766 = ( (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire811 = ( (~ pi25)  &  wire178 ) ;
 assign wire816 = ( (~ pi19)  &  (~ pi21)  &  ni34 ) | ( (~ pi19)  &  (~ pi22)  &  ni34 ) ;
 assign wire345 = ( pi25  &  wire178 ) ;
 assign wire910 = ( pi25  &  (~ ni34)  &  wire178 ) ;
 assign wire1095 = ( (~ pi19)  &  (~ pi20)  &  pi25 ) ;
 assign nv620 = ( ni34 ) | ( (~ wire157)  &  (~ n_n12782)  &  (~ wire29481) ) ;
 assign wire317 = ( ni34  &  ni31  &  (~ ni29) ) ;
 assign wire332 = ( wire6757 ) | ( (~ ni34)  &  (~ ni29) ) ;
 assign nv624 = ( n_n12782 ) | ( ni36  &  (~ wire172) ) | ( ni36  &  nv628 ) ;
 assign wire1012 = ( ni34  &  n_n12782 ) | ( ni34  &  wire29481 ) ;
 assign nv894 = ( wire1097 ) | ( wire6666 ) | ( wire6667 ) ;
 assign nv890 = ( ni34 ) | ( (~ wire157)  &  (~ wire6667)  &  (~ wire29466) ) ;
 assign wire1334 = ( ni34  &  wire1097 ) | ( ni34  &  wire6666 ) | ( ni34  &  wire6667 ) ;
 assign nv923 = ( wire1075 ) | ( wire6705 ) | ( wire6706 ) ;
 assign nv919 = ( ni34 ) | ( (~ wire157)  &  (~ wire6706)  &  (~ wire29455) ) ;
 assign n_n12619 = ( ni34  &  ni33 ) ;
 assign wire1039 = ( ni34  &  wire1075 ) | ( ni34  &  wire6705 ) | ( ni34  &  wire6706 ) ;
 assign nv1424 = ( wire184 ) | ( (~ nv6428)  &  nv919 ) | ( nv923  &  nv919 ) ;
 assign n_n12696 = ( wire604 ) | ( wire269  &  nv772 ) ;
 assign wire436 = ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign nv768 = ( n_n12696 ) | ( ni36  &  (~ wire172) ) | ( ni36  &  nv772 ) ;
 assign wire205 = ( ni37 ) | ( (~ ni36) ) ;
 assign wire1060 = ( (~ ni38)  &  (~ ni37)  &  ni36  &  nv633 ) ;
 assign nv972 = ( wire1097 ) | ( wire6616 ) | ( wire6617 ) ;
 assign nv968 = ( ni34 ) | ( (~ wire157)  &  (~ wire6617)  &  (~ wire29512) ) ;
 assign wire1046 = ( ni34  &  wire1097 ) | ( ni34  &  wire6616 ) | ( ni34  &  wire6617 ) ;
 assign nv1533 = ( wire184 ) | ( (~ nv6428)  &  nv968 ) | ( nv972  &  nv968 ) ;
 assign nv992 = ( wire1075 ) | ( wire6540 ) | ( wire6541 ) ;
 assign nv988 = ( ni34 ) | ( (~ wire157)  &  (~ wire6541)  &  (~ wire29530) ) ;
 assign wire1038 = ( ni34  &  wire1075 ) | ( ni34  &  wire6540 ) | ( ni34  &  wire6541 ) ;
 assign wire224 = ( (~ pi22)  &  ni34 ) | ( ni34  &  ni31 ) | ( ni34  &  ni30 ) ;
 assign wire312 = ( ni33  &  ni29 ) | ( ni32  &  ni29 ) ;
 assign nv801 = ( wire436 ) | ( wire6612 ) | ( wire6613 ) | ( wire6614 ) ;
 assign nv797 = ( ni34 ) | ( (~ wire157)  &  (~ wire6613)  &  (~ wire29576) ) ;
 assign wire1008 = ( ni34  &  wire6613 ) | ( ni34  &  wire6614 ) | ( ni34  &  wire29575 ) ;
 assign nv914 = ( wire1075 ) | ( wire6745 ) | ( wire6746 ) ;
 assign nv910 = ( ni34 ) | ( (~ wire157)  &  (~ wire6746)  &  (~ wire29449) ) ;
 assign wire1312 = ( ni34  &  wire1075 ) | ( ni34  &  wire6745 ) | ( ni34  &  wire6746 ) ;
 assign n_n11076 = ( wire5946 ) | ( (~ ni43)  &  wire5948 ) | ( (~ ni43)  &  wire30372 ) ;
 assign nv2190 = ( wire30369 ) | ( (~ ni42)  &  nv2186 ) | ( ni43  &  ni42  &  nv2186 ) ;
 assign wire1319 = ( ni41  &  wire5941 ) | ( ni41  &  wire5945 ) | ( ni41  &  wire30369 ) ;
 assign nv2176 = ( ni46  &  ni45 ) | ( ni47  &  (~ ni45)  &  ni48 ) ;
 assign wire621 = ( ni47 ) | ( ni45 ) ;
 assign nv2186 = ( ni46  &  ni45 ) | ( (~ ni47)  &  (~ ni45) ) | ( ni47  &  (~ ni45)  &  ni48 ) ;
 assign wire206 = ( (~ ni31)  &  (~ ni30) ) ;
 assign wire757 = ( ni33  &  ni30 ) | ( ni33  &  ni31  &  (~ ni30) ) | ( ni33  &  ni32  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire924 = ( (~ ni32)  &  (~ ni31)  &  (~ ni30) ) ;
 assign n_n9294 = ( (~ pi22)  &  wire757 ) | ( (~ pi22)  &  nv2186  &  wire924 ) ;
 assign nv2348 = ( n_n11076 ) | ( ni41  &  wire5939 ) | ( ni41  &  wire30370 ) ;
 assign wire365 = ( ni38  &  (~ ni36) ) | ( ni39  &  (~ ni37)  &  (~ ni36) ) ;
 assign n_n10860 = ( wire706 ) | ( wire5926 ) | ( nv2348  &  wire365 ) ;
 assign wire310 = ( ni38  &  ni36 ) | ( (~ ni37)  &  ni36 ) ;
 assign wire216 = ( (~ wire172)  &  nv2176  &  wire926 ) | ( (~ wire172)  &  (~ wire621)  &  wire926 ) | ( (~ wire172)  &  nv2176  &  (~ wire926) ) ;
 assign wire314 = ( ni36  &  wire216 ) ;
 assign wire253 = ( (~ ni40)  &  ni38 ) ;
 assign wire254 = ( ni40  &  ni38 ) ;
 assign nv2565 = ( wire30410 ) | ( (~ ni35)  &  wire5884 ) | ( (~ ni35)  &  wire30409 ) ;
 assign wire270 = ( ni37  &  ni36 ) ;
 assign wire347 = ( (~ ni40)  &  (~ ni37)  &  ni36 ) ;
 assign wire1181 = ( wire314 ) | ( wire346  &  wire5939 ) | ( wire346  &  wire30370 ) ;
 assign nv2397 = ( wire5404 ) | ( wire30470 ) | ( (~ ni36)  &  nv2565 ) ;
 assign wire164 = ( ni33  &  ni31 ) | ( ni33  &  ni32  &  (~ ni31) ) | ( ni33  &  (~ ni31)  &  ni30 ) ;
 assign wire240 = ( ni33  &  ni31 ) | ( ni33  &  (~ ni31)  &  (~ wire7195) ) | ( (~ ni33)  &  (~ ni31)  &  wire866  &  wire7195 ) ;
 assign wire400 = ( ni39  &  ni38  &  (~ ni36) ) | ( ni38  &  ni37  &  (~ ni36) ) | ( (~ ni39)  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire1194 = ( wire5889 ) | ( (~ ni36)  &  wire216 ) ;
 assign wire814 = ( (~ ni39)  &  ni40  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire880 = ( (~ ni40) ) | ( wire216 ) | ( wire5885 ) ;
 assign n_n10947 = ( wire5924 ) | ( wire5926 ) | ( (~ ni36)  &  wire216 ) ;
 assign nv2240 = ( ni41  &  nv2190 ) | ( (~ ni41)  &  wire30370 ) | ( ni43  &  (~ ni41)  &  nv2190 ) ;
 assign wire404 = ( ni39  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire847 = ( ni39  &  (~ ni40)  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire884 = ( ni40 ) | ( wire216 ) | ( wire5810 ) ;
 assign n_n10922 = ( wire5808 ) | ( wire5809 ) | ( n_n10947  &  wire884 ) ;
 assign n_n10896 = ( wire5920 ) | ( wire5921 ) | ( n_n10947  &  wire881 ) ;
 assign wire840 = ( ni39  &  ni40  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire881 = ( (~ ni40) ) | ( wire216 ) | ( wire5922 ) ;
 assign nv2647 = ( n_n11266 ) | ( n_n13643  &  nv2186 ) | ( (~ n_n13643)  &  wire5930 ) ;
 assign wire321 = ( wire216 ) | ( (~ ni37)  &  n_n10282 ) ;
 assign nv2183 = ( n_n11266 ) | ( (~ ni42)  &  nv2176 ) ;
 assign n_n11266 = ( wire5932 ) | ( (~ ni43)  &  wire5945 ) | ( (~ ni43)  &  wire30369 ) ;
 assign wire907 = ( (~ ni41)  &  ni44 ) ;
 assign wire1076 = ( (~ ni41)  &  (~ ni44) ) ;
 assign nv2790 = ( ni41  &  nv2647 ) | ( (~ ni41)  &  (~ ni44)  &  nv2647 ) | ( (~ ni41)  &  ni44  &  nv2183 ) ;
 assign n_n9304 = ( (~ pi21)  &  wire757 ) | ( (~ pi21)  &  wire1085  &  wire924 ) ;
 assign n_n10590 = ( wire30372 ) | ( nv2186  &  wire30371 ) ;
 assign n_n10267 = ( wire1192 ) | ( wire365  &  nv2790 ) ;
 assign wire882 = ( (~ ni40) ) | ( wire216 ) | ( (~ ni39)  &  n_n10282 ) ;
 assign wire1049 = ( wire177  &  wire216 ) | ( (~ ni37)  &  wire177  &  n_n10282 ) ;
 assign wire346 = ( ni40  &  (~ ni37)  &  ni36 ) ;
 assign wire1179 = ( ni36  &  wire216 ) | ( nv2647  &  wire346 ) ;
 assign n_n10282 = ( (~ ni38)  &  wire5941 ) | ( (~ ni38)  &  wire5945 ) | ( (~ ni38)  &  wire30369 ) ;
 assign nv2622 = ( ni41  &  nv2183 ) | ( (~ ni41)  &  (~ ni44)  &  nv2647 ) | ( (~ ni41)  &  ni44  &  nv2183 ) ;
 assign wire1192 = ( (~ ni36)  &  wire216 ) | ( (~ wire342)  &  n_n10282 ) ;
 assign n_n10396 = ( wire1192 ) | ( wire365  &  nv2622 ) ;
 assign wire1087 = ( (~ ni37)  &  ni36  &  n_n10282 ) ;
 assign nv2946 = ( n_n10396 ) | ( wire1087 ) | ( wire222  &  wire30558 ) ;
 assign wire304 = ( wire237 ) | ( ni33  &  ni31 ) ;
 assign wire751 = ( wire237 ) | ( wire5902 ) | ( ni33  &  ni31 ) ;
 assign wire866 = ( wire216 ) | ( wire172  &  n_n11266 ) | ( wire172  &  wire5930 ) ;
 assign wire252 = ( (~ ni34) ) | ( (~ ni33) ) | ( (~ nv6428) ) ;
 assign wire237 = ( ni34  &  ni33  &  wire216 ) | ( ni34  &  ni33  &  wire5904 ) ;
 assign nv2252 = ( wire240 ) | ( ni33  &  wire5470 ) | ( ni33  &  wire30505 ) ;
 assign nv2235 = ( wire5475 ) | ( wire30507 ) | ( (~ ni36)  &  nv2473 ) ;
 assign wire179 = ( pi19  &  pi21  &  pi22  &  (~ pi20) ) ;
 assign wire182 = ( pi19  &  pi21  &  pi22  &  pi20 ) ;
 assign wire166 = ( pi20  &  wire162 ) | ( (~ pi20)  &  wire159 ) ;
 assign wire378 = ( pi19  &  pi20  &  wire162 ) | ( pi19  &  (~ pi20)  &  wire159 ) ;
 assign nv2340 = ( wire240 ) | ( ni33  &  n_n10860 ) | ( ni33  &  wire30439 ) ;
 assign n_n10835 = ( wire5390 ) | ( wire5391 ) | ( n_n10860  &  wire884 ) ;
 assign wire1184 = ( wire314 ) | ( wire347  &  wire5939 ) | ( wire347  &  wire30370 ) ;
 assign nv2373 = ( wire240 ) | ( ni33  &  wire5381 ) | ( ni33  &  wire30480 ) ;
 assign wire855 = ( (~ ni47) ) | ( ni45 ) ;
 assign n_n9302 = ( (~ pi22)  &  wire757 ) | ( (~ pi22)  &  nv2176  &  wire924 ) ;
 assign nv3916 = ( (~ ni42)  &  (~ ni47) ) | ( ni42  &  ni45 ) | ( (~ ni42)  &  ni45 ) | ( ni43  &  ni42  &  (~ ni47) ) ;
 assign wire1281 = ( (~ ni41)  &  ni45 ) | ( ni43  &  (~ ni41)  &  (~ ni47) ) ;
 assign wire1296 = ( ni41  &  nv3916 ) ;
 assign nv3943 = ( wire1296 ) | ( wire4910 ) | ( wire4911 ) | ( wire4912 ) ;
 assign n_n8890 = ( (~ pi25)  &  wire4973 ) | ( (~ pi25)  &  ni32  &  ni30 ) | ( (~ pi25)  &  ni32  &  (~ ni30) ) ;
 assign nv3918 = ( ni45 ) | ( ni43  &  (~ ni47) ) ;
 assign nv4058 = ( wire4853 ) | ( wire4910 ) | ( wire4911 ) | ( wire4912 ) ;
 assign wire870 = ( (~ ni36)  &  (~ wire255) ) | ( nv3915  &  wire31260 ) ;
 assign wire489 = ( (~ wire255) ) | ( (~ ni39)  &  (~ ni38)  &  nv3916 ) ;
 assign wire989 = ( ni40 ) | ( wire489 ) ;
 assign n_n6710 = ( ni32  &  (~ ni30) ) ;
 assign n_n9194 = ( wire4967 ) | ( ni40  &  ni38  &  nv3927 ) ;
 assign n_n8976 = ( wire4957 ) | ( wire4958 ) | ( wire4959 ) ;
 assign nv3927 = ( wire1296 ) | ( wire4968 ) | ( wire4969 ) | ( wire4970 ) ;
 assign wire1180 = ( wire4950 ) | ( ni36  &  (~ wire255) ) ;
 assign n_n8862 = ( ni33  &  (~ wire255) ) | ( ni33  &  wire172  &  nv3916 ) ;
 assign wire233 = ( (~ ni29) ) | ( (~ n_n8862) ) ;
 assign wire305 = ( n_n9245 ) | ( wire4581 ) | ( (~ n_n8862)  &  wire32057 ) ;
 assign n_n6367 = ( ni32  &  (~ ni30) ) | ( (~ ni45)  &  (~ ni31)  &  (~ ni30) ) ;
 assign nv3908 = ( ni32  &  ni30 ) | ( ni32  &  (~ ni30) ) | ( (~ ni45)  &  (~ ni31)  &  (~ ni30) ) ;
 assign nv4045 = ( wire4931 ) | ( wire4968 ) | ( wire4969 ) | ( wire4970 ) ;
 assign wire1182 = ( wire347  &  nv3918 ) | ( ni36  &  (~ wire255) ) ;
 assign wire632 = ( ni38 ) | ( ni37 ) | ( (~ ni36) ) | ( (~ nv3916) ) ;
 assign wire1041 = ( ni38  &  wire31890 ) | ( (~ nv3916)  &  wire31890 ) ;
 assign nv4401 = ( wire305 ) | ( wire233  &  wire4805 ) | ( wire233  &  wire31891 ) ;
 assign wire255 = ( ni38 ) | ( (~ ni37) ) | ( ni47  &  (~ ni45) ) ;
 assign nv3915 = ( (~ wire255) ) | ( ni38  &  nv3916 ) | ( (~ ni37)  &  nv3916 ) ;
 assign n_n7885 = ( n_n6710 ) | ( wire206  &  (~ wire4897)  &  (~ wire31262) ) ;
 assign wire1065 = ( ni32  &  ni31  &  ni30 ) ;
 assign n_n8085 = ( (~ ni33)  &  ni32  &  ni30 ) | ( ni32  &  ni31  &  ni30 ) ;
 assign wire775 = ( ni32  &  (~ ni30) ) | ( (~ ni33)  &  ni32  &  ni30 ) | ( ni32  &  ni31  &  ni30 ) ;
 assign nv4932 = ( pi27  &  ni32 ) | ( pi26  &  ni32 ) | ( (~ pi27)  &  (~ pi26)  &  wire775 ) ;
 assign n_n7095 = ( (~ pi21)  &  ni32  &  wire156 ) | ( (~ pi21)  &  (~ wire156)  &  wire775 ) ;
 assign wire1098 = ( ni36  &  wire323 ) | ( (~ ni35)  &  wire323 ) ;
 assign wire834 = ( (~ ni39)  &  (~ ni40)  &  (~ ni37)  &  (~ ni36) ) ;
 assign wire992 = ( ni40 ) | ( wire492 ) ;
 assign wire689 = ( ni36  &  (~ wire255) ) ;
 assign wire1007 = ( wire4817 ) | ( (~ n_n9022)  &  wire31844 ) ;
 assign n_n8352 = ( (~ ni33)  &  (~ wire255) ) | ( (~ ni33)  &  wire172  &  nv3916 ) ;
 assign wire214 = ( (~ ni29) ) | ( (~ n_n8352) ) ;
 assign wire374 = ( n_n9245 ) | ( wire4061 ) | ( (~ n_n8352)  &  wire31171 ) ;
 assign nv6576 = ( ni47 ) | ( ni45 ) | ( wire6766 ) | ( ni43  &  (~ ni47) ) ;
 assign n_n5621 = ( wire1198 ) | ( nv669  &  wire691 ) | ( wire691  &  wire6766 ) ;
 assign nv669 = ( ni47 ) | ( ni45 ) | ( ni43  &  (~ ni47) ) ;
 assign wire827 = ( (~ ni36)  &  n_n5799  &  (~ wire390) ) | ( n_n5799  &  (~ wire390)  &  wire33267 ) ;
 assign wire1047 = ( ni40  &  (~ ni37)  &  wire3462 ) | ( ni40  &  (~ ni37)  &  wire33267 ) ;
 assign wire1081 = ( (~ ni40)  &  (~ ni37)  &  wire3462 ) | ( (~ ni40)  &  (~ ni37)  &  wire33267 ) ;
 assign wire721 = ( wire33426 ) | ( wire33427 ) | ( wire33428 ) | ( wire33429 ) ;
 assign wire464 = ( n_n2328 ) | ( ni40  &  ni38  &  nv669 ) ;
 assign n_n2328 = ( ni47  &  (~ ni38) ) | ( ni45  &  (~ ni38) ) ;
 assign n_n4404 = ( (~ ni38)  &  (~ wire157)  &  (~ wire621) ) | ( ni38  &  (~ wire157)  &  (~ nv669) ) | ( (~ wire157)  &  (~ wire621)  &  (~ nv669) ) ;
 assign nv6462 = ( wire3474 ) | ( (~ ni42)  &  wire172 ) | ( wire172  &  nv669 ) ;
 assign wire804 = ( n_n2328 ) | ( wire3431 ) | ( wire253  &  nv669 ) ;
 assign n_n4433 = ( wire33510  &  wire33513 ) | ( wire33511  &  wire33513 ) | ( wire33510  &  wire33514 ) | ( wire33511  &  wire33514 ) ;
 assign wire192 = ( ni33 ) | ( (~ ni29) ) | ( (~ nv6462) ) ;
 assign wire196 = ( ni30 ) | ( ni33  &  wire33266 ) | ( (~ nv6462)  &  wire33266 ) ;
 assign wire800 = ( n_n2328 ) | ( wire3493 ) | ( wire254  &  nv669 ) ;
 assign n_n4412 = ( wire33390  &  wire33393 ) | ( wire33391  &  wire33393 ) | ( wire33390  &  wire33394 ) | ( wire33391  &  wire33394 ) ;
 assign n_n5729 = ( wire3301 ) | ( wire3303 ) | ( wire270  &  n_n2328 ) ;
 assign n_n4489 = ( wire33302  &  wire33305 ) | ( wire33303  &  wire33305 ) | ( wire33302  &  wire33306 ) | ( wire33303  &  wire33306 ) ;
 assign wire417 = ( ni36  &  (~ ni32)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire193 = ( (~ ni33) ) | ( (~ ni29) ) | ( (~ nv6462) ) ;
 assign wire197 = ( ni30 ) | ( (~ ni33)  &  wire33776 ) | ( (~ nv6462)  &  wire33776 ) ;
 assign wire151 = ( (~ pi19)  &  pi21  &  pi22 ) ;
 assign wire173 = ( (~ pi21)  &  ni30 ) | ( pi21  &  (~ pi22)  &  ni30 ) ;
 assign wire1034 = ( (~ pi19)  &  (~ pi21)  &  ni30 ) | ( (~ pi19)  &  pi21  &  (~ pi22)  &  ni30 ) ;
 assign nv7445 = ( pi27  &  ni30 ) | ( pi26  &  ni30 ) | ( (~ pi27)  &  (~ pi26)  &  nv7447 ) ;
 assign n_n3695 = ( (~ pi21)  &  ni30  &  wire156 ) | ( (~ pi21)  &  (~ wire156)  &  nv7447 ) ;
 assign nv7647 = ( (~ pi27)  &  ni30 ) | ( pi27  &  (~ ni33)  &  ni30 ) | ( pi27  &  ni31  &  ni30 ) ;
 assign nv7791 = ( pi27  &  ni30 ) | ( (~ pi26)  &  ni30 ) | ( (~ pi27)  &  pi26  &  nv7447 ) ;
 assign n_n3349 = ( (~ pi21)  &  ni30  &  wire155 ) | ( (~ pi21)  &  (~ wire155)  &  nv7447 ) ;
 assign n_n3347 = ( (~ pi22)  &  ni30  &  wire155 ) | ( (~ pi22)  &  (~ wire155)  &  nv7447 ) ;
 assign n_n4509 = ( wire33470  &  wire33473 ) | ( wire33471  &  wire33473 ) | ( wire33470  &  wire33474 ) | ( wire33471  &  wire33474 ) ;
 assign n_n5768 = ( wire3387 ) | ( wire3389 ) | ( wire270  &  n_n2328 ) ;
 assign nv10153 = ( (~ ni30) ) | ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign n_n4501 = ( wire33590  &  wire33593 ) | ( wire33591  &  wire33593 ) | ( wire33590  &  wire33594 ) | ( wire33591  &  wire33594 ) ;
 assign n_n5752 = ( wire707 ) | ( wire3389 ) | ( nv6486  &  wire685 ) ;
 assign n_n5644 = ( wire1200 ) | ( wire3435 ) ;
 assign n_n3693 = ( (~ pi22)  &  ni30  &  wire156 ) | ( (~ pi22)  &  (~ wire156)  &  nv7447 ) ;
 assign n_n5514 = ( wire826 ) | ( wire1064 ) | ( nv6589  &  wire857 ) ;
 assign nv6589 = ( wire6727 ) | ( ni41  &  nv669 ) | ( (~ ni41)  &  nv669 ) ;
 assign wire477 = ( (~ ni36) ) | ( nv9066 ) ;
 assign wire1074 = ( (~ ni37)  &  (~ ni32)  &  (~ ni31)  &  (~ ni30) ) ;
 assign nv7105 = ( wire196 ) | ( wire192  &  wire3214 ) | ( wire192  &  wire3215 ) ;
 assign n_n4543 = ( wire3193 ) | ( (~ ni36)  &  n_n4404 ) | ( n_n4404  &  nv9066 ) ;
 assign n_n5574 = ( wire826 ) | ( wire1064 ) | ( nv6486  &  wire857 ) ;
 assign nv6486 = ( wire6727 ) | ( (~ ni42)  &  ni41 ) | ( ni41  &  nv669 ) | ( (~ ni41)  &  nv669 ) ;
 assign nv7050 = ( wire196 ) | ( wire192  &  wire3307 ) | ( wire192  &  wire3308 ) ;
 assign n_n4473 = ( wire3276 ) | ( (~ ni38)  &  (~ wire157)  &  (~ wire621) ) ;
 assign n_n4611 = ( wire3274 ) | ( wire477  &  wire3276 ) | ( wire477  &  wire3277 ) ;
 assign wire802 = ( wire465 ) | ( ni40  &  ni38  &  nv6486 ) ;
 assign nv6472 = ( nv669 ) | ( wire6766 ) | ( (~ ni42)  &  ni41 ) ;
 assign n_n5580 = ( wire827 ) | ( wire1064 ) | ( nv6472  &  wire861 ) ;
 assign nv6789 = ( wire197 ) | ( wire193  &  wire3326 ) | ( wire193  &  wire3327 ) ;
 assign nv8372 = ( ni33  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign n_n3016 = ( wire3149 ) | ( nv8372  &  wire33939 ) ;
 assign nv6859 = ( wire197 ) | ( wire193  &  wire3214 ) | ( wire193  &  wire3215 ) ;
 assign wire822 = ( pi24  &  ni33  &  ni30 ) | ( pi24  &  ni31  &  ni30 ) ;
 assign wire336 = ( wire3156 ) | ( (~ pi21)  &  wire822 ) | ( (~ pi22)  &  wire822 ) ;
 assign wire1044 = ( pi21  &  pi22  &  pi24 ) ;
 assign wire1063 = ( ni30  &  (~ wire150) ) | ( (~ wire150)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign nv8638 = ( wire336 ) | ( wire3153 ) | ( (~ pi24)  &  wire1063 ) ;
 assign wire405 = ( wire1982 ) | ( (~ pi22)  &  (~ ni29) ) ;
 assign n_n1241 = ( wire405 ) | ( (~ pi22)  &  wire35140 ) | ( (~ pi22)  &  wire35141 ) ;
 assign wire245 = ( ni31  &  (~ ni30)  &  ni29 ) ;
 assign wire293 = ( (~ ni32)  &  ni30  &  ni29 ) ;
 assign wire316 = ( (~ ni31)  &  (~ ni30)  &  ni29 ) ;
 assign wire877 = ( wire1479 ) | ( (~ ni35)  &  wire266  &  wire348 ) ;
 assign wire308 = ( wire35005 ) | ( (~ pi21)  &  ni32 ) | ( (~ pi21)  &  ni30 ) ;
 assign n_n1243 = ( wire308 ) | ( (~ pi21)  &  wire35135 ) | ( (~ pi21)  &  wire35136 ) ;
 assign wire1019 = ( ni38  &  ni36 ) | ( ni38  &  ni35 ) ;
 assign wire1075 = ( (~ ni38)  &  ni37  &  wire177 ) | ( (~ ni38)  &  (~ ni37)  &  wire177  &  nv633 ) ;
 assign n_n2176 = ( wire35325 ) | ( wire316  &  wire6703 ) | ( wire316  &  wire29653 ) ;
 assign wire189 = ( pi21  &  pi22  &  pi20 ) ;
 assign wire194 = ( pi17  &  (~ pi16)  &  wire152 ) ;
 assign wire295 = ( pi17  &  pi19  &  (~ pi16) ) ;
 assign wire309 = ( pi21  &  pi22  &  pi20  &  (~ ni29) ) ;
 assign wire456 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire700 = ( wire309  &  wire259 ) ;
 assign wire1109 = ( (~ ni29)  &  wire259 ) ;
 assign n_n2483 = ( wire35597 ) | ( (~ pi16)  &  wire1148 ) | ( (~ pi16)  &  wire35588 ) ;
 assign nv839 = ( wire436 ) | ( wire6536 ) | ( wire6537 ) | ( wire6538 ) ;
 assign wire183 = ( pi17  &  pi16  &  wire152 ) ;
 assign wire257 = ( pi17  &  pi19  &  pi16 ) ;
 assign wire476 = ( pi17  &  pi25  &  pi16 ) ;
 assign wire487 = ( pi20  &  (~ ni29)  &  wire153 ) ;
 assign wire593 = ( pi17  &  (~ pi19)  &  pi16 ) ;
 assign wire626 = ( wire1567 ) | ( wire35237 ) | ( n_n1824  &  wire35236 ) ;
 assign wire758 = ( wire1623 ) | ( wire1626 ) | ( wire35257 ) | ( wire35258 ) ;
 assign wire786 = ( wire1228 ) | ( wire191  &  wire1952 ) | ( wire191  &  wire35210 ) ;
 assign wire1027 = ( (~ pi17)  &  (~ pi19)  &  pi25 ) ;
 assign wire1322 = ( pi20  &  (~ ni29)  &  wire259  &  wire153 ) ;
 assign wire1344 = ( (~ pi17)  &  pi19  &  pi25 ) ;
 assign n_n2484 = ( wire894 ) | ( wire931 ) | ( wire961 ) | ( wire35559 ) ;
 assign n_n1649 = ( wire35116 ) | ( wire316  &  wire6746 ) | ( wire316  &  wire29449 ) ;
 assign n_n1247 = ( wire308 ) | ( (~ pi21)  &  wire35112 ) | ( (~ pi21)  &  wire35113 ) ;
 assign n_n1111 = ( wire35118 ) | ( wire213  &  wire1535 ) | ( wire213  &  wire35116 ) ;
 assign wire361 = ( (~ pi22) ) | ( ni31 ) | ( ni32  &  (~ ni31) ) | ( (~ ni31)  &  ni30 ) ;
 assign n_n1119 = ( wire35158 ) | ( wire213  &  wire1516 ) | ( wire213  &  wire35156 ) ;
 assign nv883 = ( wire6453 ) | ( wire6454 ) | ( wire29476 ) ;
 assign n_n1253 = ( wire405 ) | ( (~ pi22)  &  wire35102 ) | ( (~ pi22)  &  wire35103 ) ;
 assign n_n1263 = ( wire405 ) | ( (~ pi22)  &  wire860 ) | ( (~ pi22)  &  wire35094 ) ;
 assign n_n1255 = ( wire308 ) | ( (~ pi21)  &  wire35122 ) | ( (~ pi21)  &  wire35123 ) ;
 assign wire163 = ( (~ pi17)  &  (~ pi19) ) ;
 assign wire171 = ( pi20  &  wire153 ) ;
 assign wire817 = ( (~ pi17)  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign n_n1813 = ( wire603 ) | ( wire609 ) | ( wire35506 ) | ( wire35507 ) ;
 assign wire213 = ( pi21  &  pi22  &  (~ pi20) ) ;
 assign wire506 = ( pi21  &  (~ pi22)  &  (~ pi20) ) ;
 assign wire508 = ( wire2065 ) | ( wire218  &  wire34995 ) ;
 assign wire226 = ( pi16  &  pi15 ) ;
 assign wire154 = ( pi17  &  pi16 ) ;
 assign wire485 = ( pi17  &  pi19  &  pi16  &  pi15 ) ;
 assign nv9492 = ( (~ ni38)  &  ni37 ) | ( ni38  &  nv9031 ) | ( (~ ni38)  &  (~ ni37)  &  wire771 ) ;
 assign wire259 = ( (~ pi25) ) | ( ni31 ) | ( ni32  &  (~ ni31) ) | ( (~ ni31)  &  ni30 ) ;
 assign nv858 = ( (~ ni38)  &  ni37 ) | ( ni38  &  wire388 ) | ( (~ ni38)  &  (~ ni37)  &  nv633 ) ;
 assign wire853 = ( wire1391 ) | ( wire1394 ) | ( wire1395 ) | ( wire35017 ) ;
 assign nv740 = ( wire6694 ) | ( (~ ni38)  &  ni37 ) | ( (~ ni38)  &  (~ ni37)  &  nv633 ) ;
 assign n_n1593 = ( wire1196 ) | ( wire1484 ) | ( wire1485 ) | ( wire1486 ) ;
 assign nv9031 = ( ni43 ) | ( ni42 ) | ( ni47 ) ;
 assign wire897 = ( (~ ni39)  &  (~ ni32) ) | ( ni38  &  (~ ni32) ) | ( ni36  &  (~ ni32) ) ;
 assign n_n2466 = ( ni39  &  ni47 ) | ( ni39  &  (~ ni43)  &  ni42 ) ;
 assign wire703 = ( (~ ni38)  &  ni37  &  (~ ni32) ) ;
 assign wire999 = ( wire703 ) | ( n_n2466  &  wire35060 ) ;
 assign wire1101 = ( ni43  &  (~ ni40) ) | ( ni42  &  (~ ni40) ) | ( (~ ni43)  &  (~ ni40)  &  ni45 ) ;
 assign wire278 = ( ni36  &  ni32 ) | ( (~ ni35)  &  ni32 ) ;
 assign wire607 = ( (~ ni38)  &  ni37  &  (~ ni36) ) | ( (~ ni38)  &  (~ ni36)  &  n_n2448 ) ;
 assign wire1082 = ( (~ ni38)  &  ni37  &  wire278 ) | ( (~ ni38)  &  (~ ni37)  &  wire278  &  wire770 ) ;
 assign wire806 = ( ni37  &  ni36  &  ni32 ) | ( ni37  &  (~ ni36)  &  ni35  &  ni32 ) ;
 assign n_n2448 = ( ni39  &  ni45 ) | ( ni39  &  (~ ni43)  &  ni42 ) ;
 assign wire1304 = ( (~ ni38)  &  (~ ni36)  &  n_n2448 ) ;
 assign nv9029 = ( ni41  &  (~ ni40) ) | ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( ni41  &  ni40  &  (~ nv9031) ) | ( ni40  &  (~ ni44)  &  (~ nv9031) ) ;
 assign wire341 = ( ni36  &  (~ ni32) ) ;
 assign wire589 = ( (~ ni38)  &  ni37  &  ni36  &  (~ ni32) ) ;
 assign n_n2332 = ( wire35309 ) | ( (~ ni36)  &  wire35152 ) | ( (~ ni36)  &  wire35153 ) ;
 assign wire1146 = ( ni36  &  ni32 ) | ( (~ ni35)  &  ni32  &  nv9066 ) ;
 assign nv662 = ( wire436 ) | ( wire6662 ) | ( wire6663 ) | ( wire6664 ) ;
 assign nv628 = ( ni42 ) | ( nv669 ) | ( wire6766 ) | ( (~ ni42)  &  ni41 ) ;
 assign wire418 = ( ni30  &  ni29 ) ;
 assign n_n2327 = ( wire1832 ) | ( wire1835 ) | ( wire35311 ) ;
 assign wire606 = ( (~ ni38)  &  ni37  &  (~ ni36) ) | ( (~ ni38)  &  (~ ni36)  &  n_n1966 ) ;
 assign n_n1966 = ( (~ ni39)  &  ni45 ) | ( (~ ni39)  &  (~ ni43)  &  ni42 ) ;
 assign wire1302 = ( (~ ni38)  &  (~ ni36)  &  n_n1966 ) ;
 assign wire512 = ( ni43 ) | ( ni42 ) | ( ni41 ) | ( ni47 ) ;
 assign nv9129 = ( ni41  &  ni40 ) | ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( ni41  &  (~ ni40)  &  (~ nv9031) ) | ( (~ ni40)  &  (~ ni44)  &  (~ nv9031) ) ;
 assign wire1231 = ( wire703 ) | ( (~ ni37)  &  n_n1574  &  wire835 ) ;
 assign n_n2228 = ( wire35289 ) | ( (~ ni36)  &  wire35112 ) | ( (~ ni36)  &  wire35113 ) ;
 assign wire461 = ( (~ ni35)  &  ni32 ) ;
 assign wire1142 = ( ni36  &  ni32 ) | ( ni35  &  ni32  &  nv9066 ) ;
 assign nv9173 = ( ni41  &  ni40 ) | ( ni41  &  (~ ni40) ) | ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( (~ ni41)  &  (~ ni40)  &  ni44 ) ;
 assign n_n2179 = ( wire35321 ) | ( (~ ni36)  &  wire35135 ) | ( (~ ni36)  &  wire35136 ) ;
 assign n_n2180 = ( wire35322 ) | ( (~ nv539)  &  wire35140 ) | ( (~ nv539)  &  wire35141 ) ;
 assign wire398 = ( (~ ni38)  &  ni37 ) | ( (~ ni38)  &  (~ ni37)  &  wire771 ) ;
 assign wire770 = ( ni45 ) | ( (~ ni43)  &  ni42 ) ;
 assign n_n1566 = ( ni45  &  (~ ni38) ) | ( (~ ni43)  &  ni42  &  (~ ni38) ) ;
 assign n_n5610 = ( (~ ni39)  &  ni47 ) | ( (~ ni39)  &  ni45 ) ;
 assign nv9066 = ( ni38 ) | ( ni37 ) | ( ni47  &  (~ ni38) ) | ( ni45  &  (~ ni38) ) ;
 assign wire951 = ( ni37 ) | ( (~ ni36) ) | ( ni39  &  ni38 ) | ( ni38  &  ni36 ) ;
 assign n_n1574 = ( ni47  &  (~ ni38) ) | ( (~ ni43)  &  ni42  &  (~ ni38) ) ;
 assign wire1022 = ( (~ ni37)  &  ni36  &  (~ ni32)  &  n_n1574 ) ;
 assign n_n1786 = ( wire1022 ) | ( wire999  &  wire951 ) | ( wire951  &  wire1883 ) ;
 assign wire952 = ( ni37 ) | ( (~ ni36) ) | ( ni38  &  (~ ni37) ) ;
 assign n_n1756 = ( wire1022 ) | ( wire952  &  wire1000 ) | ( wire952  &  wire1710 ) ;
 assign wire408 = ( ni41 ) | ( (~ ni41)  &  ni44 ) | ( (~ ni41)  &  wire934 ) ;
 assign wire782 = ( ni37 ) | ( (~ ni36) ) | ( (~ ni32) ) ;
 assign wire860 = ( ni32  &  wire35092 ) | ( ni36  &  ni32  &  n_n2404 ) | ( (~ ni36)  &  ni32  &  n_n2404 ) ;
 assign nv644 = ( wire6722 ) | ( wire29474 ) | ( wire29475 ) ;
 assign n_n13028 = ( (~ ni38)  &  ni37 ) | ( ni37  &  wire441 ) ;
 assign wire266 = ( ni32  &  ni30  &  ni29 ) ;
 assign wire348 = ( wire33310 ) | ( (~ ni36)  &  n_n5610 ) | ( ni36  &  nv9066 ) ;
 assign wire1230 = ( wire703 ) | ( (~ ni37)  &  n_n1574  &  wire836 ) ;
 assign n_n1259 = ( wire308 ) | ( (~ pi21)  &  wire35152 ) | ( (~ pi21)  &  wire35153 ) ;
 assign wire327 = ( ni36  &  ni32 ) | ( ni35  &  ni32 ) ;
 assign wire1023 = ( (~ ni38)  &  ni37  &  wire327 ) | ( (~ ni38)  &  (~ ni37)  &  wire770  &  wire327 ) ;
 assign n_n1984 = ( (~ ni39)  &  ni47 ) | ( (~ ni39)  &  (~ ni43)  &  ni42 ) ;
 assign wire701 = ( ni35  &  ni32  &  ni30  &  ni29 ) ;
 assign nv235 = ( nv212 ) | ( nv69  &  (~ nv121)  &  (~ n_n13755) ) ;
 assign wire340 = ( (~ pi17)  &  (~ pi19)  &  pi20 ) | ( (~ pi17)  &  (~ pi19)  &  (~ pi20) ) ;
 assign wire381 = ( (~ pi17)  &  pi19  &  pi20 ) ;
 assign wire616 = ( (~ pi17)  &  pi19  &  (~ pi20) ) ;
 assign n_n12706 = ( wire500 ) | ( nv758  &  wire292 ) ;
 assign nv754 = ( n_n12706 ) | ( ni36  &  (~ wire172) ) | ( ni36  &  nv758 ) ;
 assign nv942 = ( wire1060 ) | ( n_n12706 ) | ( wire222  &  wire29534 ) ;
 assign wire785 = ( wire157 ) | ( wire6722 ) | ( wire29474 ) | ( wire29475 ) ;
 assign nv750 = ( ni34 ) | ( (~ wire157)  &  (~ n_n12706)  &  (~ wire29534) ) ;
 assign wire1048 = ( ni34  &  n_n12706 ) | ( ni34  &  wire29534 ) ;
 assign nv1162 = ( wire184 ) | ( (~ nv6428)  &  nv750 ) | ( nv754  &  nv750 ) ;
 assign nv928 = ( ni34 ) | ( (~ wire320)  &  (~ wire157)  &  (~ wire6694) ) ;
 assign wire1036 = ( ni34  &  wire320 ) | ( ni34  &  wire6694 ) ;
 assign nv1445 = ( wire184 ) | ( (~ nv6428)  &  nv928 ) | ( nv740  &  nv928 ) ;
 assign nv873 = ( wire1060 ) | ( n_n12782 ) | ( wire222  &  wire29481 ) ;
 assign nv983 = ( wire1075 ) | ( wire6560 ) | ( wire6561 ) ;
 assign nv979 = ( ni34 ) | ( (~ wire157)  &  (~ wire6561)  &  (~ wire29526) ) ;
 assign wire1313 = ( ni34  &  wire1075 ) | ( ni34  &  wire6560 ) | ( ni34  &  wire6561 ) ;
 assign wire322 = ( wire216 ) | ( wire5917 ) ;
 assign nv2197 = ( wire314 ) | ( wire1194 ) | ( wire5775 ) | ( wire5839 ) ;
 assign wire1111 = ( (~ ni38)  &  (~ wire205)  &  n_n11266 ) | ( (~ ni38)  &  (~ wire205)  &  wire5930 ) ;
 assign nv2493 = ( wire30384 ) | ( (~ ni35)  &  wire5838 ) | ( (~ ni35)  &  wire30383 ) ;
 assign wire238 = ( ni34  &  (~ ni33)  &  (~ wire157) ) ;
 assign wire307 = ( wire164 ) | ( wire237 ) | ( wire866  &  wire30522 ) ;
 assign wire315 = ( (~ ni34)  &  ni33  &  (~ ni32) ) ;
 assign wire706 = ( (~ ni36)  &  wire216 ) ;
 assign nv2793 = ( wire30603 ) | ( n_n10267  &  wire238 ) | ( wire238  &  wire30528 ) ;
 assign nv3060 = ( n_n10267 ) | ( wire1087 ) | ( wire222  &  wire30528 ) ;
 assign nv2534 = ( n_n10860 ) | ( wire1111 ) | ( wire222  &  wire30439 ) ;
 assign nv2930 = ( wire1087 ) | ( n_n10412 ) | ( wire222  &  wire30538 ) ;
 assign nv2627 = ( wire30667 ) | ( n_n10396  &  wire238 ) | ( wire238  &  wire30558 ) ;
 assign nv2330 = ( wire314 ) | ( wire1194 ) | ( wire5416 ) | ( wire5887 ) ;
 assign nv2766 = ( wire314 ) | ( wire1195 ) | ( wire5549 ) | ( wire5591 ) ;
 assign nv2995 = ( wire30569 ) | ( (~ ni35)  &  wire5705 ) | ( (~ ni35)  &  wire30568 ) ;
 assign nv2314 = ( wire216 ) | ( wire5917 ) | ( ni38  &  nv2240 ) ;
 assign nv2963 = ( wire30549 ) | ( ni35  &  wire5725 ) | ( ni35  &  wire30548 ) ;
 assign nv2473 = ( wire30424 ) | ( ni35  &  wire5797 ) | ( ni35  &  wire30423 ) ;
 assign nv3109 = ( wire30614 ) | ( (~ ni35)  &  wire5590 ) | ( (~ ni35)  &  wire30613 ) ;
 assign nv2545 = ( wire30442 ) | ( ni35  &  wire5376 ) | ( ni35  &  wire30441 ) ;
 assign nv3077 = ( wire30590 ) | ( ni35  &  wire5577 ) | ( ni35  &  wire30589 ) ;
 assign nv2857 = ( wire5583 ) | ( wire30616 ) | ( (~ ni36)  &  nv3109 ) ;
 assign nv2807 = ( wire5567 ) | ( wire30592 ) | ( (~ ni36)  &  nv3077 ) ;
 assign nv2359 = ( wire5368 ) | ( wire30475 ) | ( (~ ni36)  &  nv2545 ) ;
 assign wire169 = ( (~ pi20)  &  wire153 ) ;
 assign wire763 = ( pi20  &  pi16  &  wire153 ) ;
 assign wire344 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire324 = ( pi19  &  pi21  &  pi22  &  pi20 ) | ( pi19  &  pi21  &  pi22  &  (~ pi20) ) ;
 assign wire1024 = ( (~ pi20)  &  pi16  &  wire153 ) ;
 assign wire1061 = ( (~ pi17)  &  pi16 ) ;
 assign wire1069 = ( (~ pi15)  &  ni14 ) ;
 assign wire1309 = ( pi17  &  pi16  &  wire324 ) ;
 assign wire208 = ( pi17  &  pi19  &  pi16 ) | ( (~ pi17)  &  (~ pi19)  &  pi16 ) ;
 assign wire1341 = ( pi20  &  wire208  &  wire162 ) | ( (~ pi20)  &  wire208  &  wire159 ) ;
 assign n_n9022 = ( (~ ni47)  &  (~ ni38) ) | ( ni45  &  (~ ni38) ) ;
 assign nv3961 = ( ni41  &  nv3916 ) | ( (~ ni41)  &  nv3918 ) ;
 assign wire323 = ( (~ ni38)  &  ni37  &  wire855 ) | ( (~ ni38)  &  (~ ni37)  &  nv3916 ) ;
 assign wire1185 = ( wire346  &  nv3918 ) | ( ni36  &  (~ wire255) ) ;
 assign n_n9141 = ( wire4904 ) | ( (~ ni40)  &  ni38  &  nv3943 ) ;
 assign wire990 = ( (~ ni40) ) | ( wire489 ) ;
 assign n_n8948 = ( wire4899 ) | ( wire4900 ) | ( wire4901 ) ;
 assign wire1103 = ( ni36  &  wire323 ) | ( ni35  &  wire323 ) ;
 assign n_n7845 = ( n_n6710 ) | ( wire206  &  (~ wire4922)  &  (~ wire31680) ) ;
 assign wire369 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire370 = ( (~ pi15)  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire613 = ( ni13  &  (~ ni12) ) | ( (~ ni14)  &  (~ ni12) ) ;
 assign wire279 = ( wire170 ) | ( ni32  &  ni30  &  wire181 ) ;
 assign wire387 = ( pi21  &  pi22  &  (~ pi20)  &  pi25 ) ;
 assign wire473 = ( wire32018 ) | ( wire170  &  wire198 ) ;
 assign wire705 = ( pi25  &  (~ pi16) ) ;
 assign wire1028 = ( pi21  &  pi22  &  pi20  &  (~ pi25) ) ;
 assign wire1053 = ( pi21  &  pi22  &  (~ pi20)  &  (~ pi25) ) ;
 assign wire1113 = ( (~ pi25)  &  (~ pi16) ) ;
 assign wire1203 = ( wire908 ) | ( wire476  &  wire4827 ) | ( wire476  &  wire31949 ) ;
 assign wire1245 = ( wire4802 ) | ( wire4803 ) | ( n_n7913  &  wire475 ) ;
 assign wire1246 = ( wire1329 ) | ( wire4776 ) | ( n_n7837  &  wire437 ) ;
 assign wire1288 = ( (~ pi20)  &  wire170 ) | ( (~ pi20)  &  n_n9245  &  wire181 ) ;
 assign wire698 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire1031 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign n_n7837 = ( n_n6710 ) | ( wire206  &  (~ wire4793)  &  (~ wire31598) ) ;
 assign wire258 = ( pi16  &  (~ pi15) ) ;
 assign n_n9255 = ( wire922 ) | ( wire4653 ) | ( wire4678 ) | ( wire32033 ) ;
 assign wire153 = ( (~ pi17)  &  (~ pi19)  &  pi21  &  pi22 ) ;
 assign wire437 = ( (~ pi17)  &  pi25  &  wire182 ) ;
 assign wire895 = ( wire473 ) | ( n_n8890  &  wire153 ) | ( n_n8890  &  wire32019 ) ;
 assign wire904 = ( wire32013 ) | ( (~ pi22)  &  (~ pi16)  &  nv3908 ) ;
 assign wire1110 = ( pi17  &  pi21  &  pi22  &  (~ pi16) ) ;
 assign n_n7816 = ( n_n6710 ) | ( wire206  &  (~ wire4844)  &  (~ wire31352) ) ;
 assign n_n7945 = ( wire4175 ) | ( wire4183 ) | ( wire32831 ) | ( wire32832 ) ;
 assign n_n7825 = ( n_n6710 ) | ( wire206  &  (~ wire4834)  &  (~ wire31434) ) ;
 assign wire181 = ( pi21  &  pi22  &  pi25 ) ;
 assign wire227 = ( (~ pi21)  &  nv4932 ) | ( pi21  &  (~ pi22)  &  nv4938 ) ;
 assign wire274 = ( pi25  &  wire187 ) | ( (~ pi25)  &  wire4448 ) | ( (~ pi25)  &  wire4449 ) ;
 assign wire474 = ( pi25  &  wire182 ) ;
 assign wire765 = ( (~ pi15)  &  (~ ni14) ) ;
 assign wire908 = ( pi25  &  wire152  &  wire154  &  n_n7808 ) ;
 assign wire920 = ( pi15  &  (~ ni14) ) ;
 assign wire1329 = ( n_n6710  &  wire219 ) | ( wire219  &  wire4778 ) | ( wire219  &  wire4779 ) ;
 assign wire358 = ( pi25  &  wire179 ) ;
 assign wire1290 = ( wire474  &  wire31838 ) | ( wire474  &  wire31839 ) | ( wire474  &  wire31840 ) ;
 assign wire1292 = ( wire457  &  wire31338 ) | ( wire457  &  wire31339 ) | ( wire457  &  wire31340 ) ;
 assign wire1351 = ( wire393  &  wire4613 ) | ( wire393  &  wire31347 ) ;
 assign wire201 = ( n_n6922 ) | ( wire4435 ) | ( wire4436 ) ;
 assign wire249 = ( wire32720 ) | ( (~ pi25)  &  wire4433 ) | ( (~ pi25)  &  wire4434 ) ;
 assign wire922 = ( wire311  &  wire928 ) | ( wire311  &  wire4680 ) | ( wire311  &  wire4681 ) ;
 assign wire1308 = ( wire457  &  wire31428 ) | ( wire457  &  wire31429 ) | ( wire457  &  wire31430 ) ;
 assign n_n7905 = ( n_n6710 ) | ( wire206  &  (~ wire4862)  &  (~ wire31762) ) ;
 assign wire457 = ( pi25  &  wire180 ) ;
 assign wire1279 = ( pi25  &  wire158  &  wire152  &  n_n7877 ) ;
 assign n_n7702 = ( wire4112 ) | ( wire4115 ) | ( wire32741 ) | ( wire32742 ) ;
 assign n_n6922 = ( (~ pi27)  &  (~ pi21)  &  ni32 ) | ( pi27  &  (~ pi21)  &  wire775 ) ;
 assign wire165 = ( ni13 ) | ( (~ ni14) ) ;
 assign wire268 = ( (~ ni13)  &  ni14  &  (~ ni11)  &  ni12 ) ;
 assign wire618 = ( ni13  &  (~ ni11)  &  ni12 ) ;
 assign wire247 = ( pi20  &  pi25  &  wire153 ) ;
 assign wire818 = ( (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire845 = ( (~ pi15)  &  wire268 ) ;
 assign wire848 = ( pi15  &  wire268 ) ;
 assign n_n7808 = ( n_n6710 ) | ( wire206  &  (~ wire323)  &  (~ wire4824) ) ;
 assign wire311 = ( pi17  &  pi25  &  pi16  &  wire152 ) ;
 assign nv4938 = ( n_n9245  &  wire156 ) | ( wire156  &  n_n6367 ) | ( (~ wire156)  &  n_n6367 ) | ( (~ wire156)  &  n_n8085 ) ;
 assign wire991 = ( (~ ni40) ) | ( wire492 ) ;
 assign nv5285 = ( n_n9245  &  wire155 ) | ( wire155  &  n_n6367 ) | ( (~ wire155)  &  n_n6367 ) | ( (~ wire155)  &  n_n8085 ) ;
 assign nv4409 = ( wire305 ) | ( wire233  &  wire4811 ) | ( wire233  &  wire31893 ) ;
 assign wire170 = ( (~ pi21)  &  ni32 ) | ( pi21  &  (~ pi22)  &  nv3908 ) ;
 assign wire484 = ( (~ pi17)  &  (~ pi16)  &  wire182 ) ;
 assign wire587 = ( (~ pi17)  &  (~ pi16)  &  wire179 ) ;
 assign wire1118 = ( (~ wire150)  &  wire4973 ) | ( ni32  &  ni30  &  (~ wire150) ) | ( ni32  &  (~ ni30)  &  (~ wire150) ) ;
 assign wire221 = ( (~ pi21)  &  nv5283 ) | ( pi21  &  (~ pi22)  &  nv5285 ) ;
 assign wire352 = ( wire221 ) | ( (~ wire150)  &  wire4458 ) | ( (~ wire150)  &  wire4459 ) ;
 assign wire263 = ( (~ ni13)  &  (~ ni14) ) ;
 assign wire377 = ( (~ ni13)  &  (~ ni14)  &  (~ ni11)  &  ni12 ) ;
 assign wire453 = ( wire227 ) | ( (~ wire150)  &  wire4448 ) | ( (~ wire150)  &  wire4449 ) ;
 assign wire699 = ( (~ ni13)  &  ni14  &  ni11  &  (~ ni12) ) ;
 assign wire1339 = ( ni13  &  ni11 ) | ( (~ ni14)  &  ni11 ) | ( ni11  &  ni12 ) ;
 assign wire788 = ( ni13  &  ni11 ) | ( (~ ni14)  &  ni11 ) | ( ni13  &  ni12 ) | ( ni11  &  ni12 ) ;
 assign wire791 = ( wire201 ) | ( (~ wire150)  &  wire4433 ) | ( (~ wire150)  &  wire4434 ) ;
 assign nv5843 = ( wire32489 ) | ( (~ ni11)  &  wire4419 ) | ( (~ ni11)  &  wire32181 ) ;
 assign wire1189 = ( wire4649 ) | ( ni36  &  (~ wire255) ) ;
 assign n_n5481 = ( (~ pi25)  &  ni30 ) | ( (~ pi25)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire801 = ( wire465 ) | ( wire3383 ) ;
 assign wire1006 = ( (~ ni36)  &  (~ wire157) ) | ( (~ wire157)  &  wire33600 ) ;
 assign n_n4441 = ( wire33550  &  wire33553 ) | ( wire33551  &  wire33553 ) | ( wire33550  &  wire33554 ) | ( wire33551  &  wire33554 ) ;
 assign wire826 = ( (~ ni36)  &  n_n5610  &  (~ wire390) ) | ( n_n5610  &  (~ wire390)  &  wire33310 ) ;
 assign wire857 = ( wire3314 ) | ( (~ ni37)  &  wire3491 ) | ( (~ ni37)  &  wire33310 ) ;
 assign wire1064 = ( ni37  &  (~ ni36)  &  n_n2328 ) ;
 assign n_n5520 = ( wire827 ) | ( wire1064 ) | ( nv6576  &  wire861 ) ;
 assign nv7098 = ( wire196 ) | ( wire192  &  wire3205 ) | ( wire192  &  wire3206 ) ;
 assign nv7129 = ( wire196 ) | ( wire192  &  wire3185 ) | ( wire192  &  wire3186 ) ;
 assign wire209 = ( (~ pi21)  &  nv7647 ) | ( pi21  &  (~ pi22)  &  nv7647 ) ;
 assign wire199 = ( (~ pi17)  &  wire179 ) ;
 assign wire450 = ( wire2563 ) | ( wire196  &  wire171 ) | ( wire171  &  wire2566 ) ;
 assign wire448 = ( pi20  &  wire153 ) | ( (~ pi20)  &  wire153 ) ;
 assign wire251 = ( pi17  &  pi16  &  wire178 ) ;
 assign wire244 = ( pi17  &  pi16  &  wire180 ) ;
 assign wire653 = ( wire34119 ) | ( nv10153  &  wire2545 ) | ( nv10153  &  wire34111 ) ;
 assign wire203 = ( (~ pi17)  &  wire182 ) ;
 assign wire690 = ( (~ pi17)  &  pi27  &  wire182 ) ;
 assign wire797 = ( wire463 ) | ( wire3297 ) ;
 assign n_n3014 = ( wire3147 ) | ( nv8372  &  wire33940 ) ;
 assign wire335 = ( wire3144 ) | ( wire3149 ) | ( nv8372  &  wire33939 ) ;
 assign nv8369 = ( wire335 ) | ( wire3141 ) | ( wire161  &  wire1063 ) ;
 assign nv10167 = ( (~ ni30) ) | ( ni33  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire861 = ( wire3337 ) | ( (~ ni37)  &  wire3462 ) | ( (~ ni37)  &  wire33267 ) ;
 assign wire501 = ( wire385 ) | ( wire197  &  wire199 ) | ( wire199  &  wire3391 ) ;
 assign wire655 = ( wire34465 ) | ( nv10167  &  wire3019 ) | ( nv10167  &  wire34457 ) ;
 assign wire828 = ( (~ pi17)  &  pi24  &  wire182 ) ;
 assign wire1114 = ( (~ pi17)  &  (~ pi24)  &  wire182 ) ;
 assign wire641 = ( wire447 ) | ( wire197  &  wire203 ) | ( wire203  &  wire3316 ) ;
 assign wire673 = ( wire34496 ) | ( nv10167  &  wire2994 ) | ( nv10167  &  wire34488 ) ;
 assign wire678 = ( wire34488 ) | ( wire197  &  wire243 ) | ( wire243  &  wire3249 ) ;
 assign wire891 = ( wire528 ) | ( wire199  &  wire2984 ) | ( wire199  &  wire34484 ) ;
 assign wire1090 = ( (~ pi17)  &  (~ pi24)  &  wire179 ) ;
 assign wire649 = ( wire34395 ) | ( nv10167  &  wire2961 ) | ( nv10167  &  wire33833 ) ;
 assign wire652 = ( wire34436 ) | ( nv10167  &  wire2946 ) | ( nv10167  &  wire34427 ) ;
 assign n_n4481 = ( wire33345  &  wire33348 ) | ( wire33346  &  wire33348 ) | ( wire33345  &  wire33349 ) | ( wire33346  &  wire33349 ) ;
 assign wire250 = ( pi17  &  (~ pi16)  &  wire178 ) ;
 assign wire243 = ( pi17  &  (~ pi16)  &  wire180 ) ;
 assign wire898 = ( ni39  &  (~ ni32) ) | ( ni38  &  (~ ni32) ) | ( ni36  &  (~ ni32) ) ;
 assign wire1000 = ( wire703 ) | ( n_n1984  &  wire35079 ) ;
 assign n_n2404 = ( wire1708 ) | ( (~ ni38)  &  ni37 ) ;
 assign wire820 = ( ni32  &  ni31  &  (~ ni30)  &  ni29 ) ;
 assign wire841 = ( ni36  &  ni32  &  ni30  &  ni29 ) ;
 assign wire1248 = ( ni36  &  wire266 ) | ( wire266  &  wire33310 ) | ( (~ ni36)  &  n_n5610  &  wire266 ) ;
 assign nv9082 = ( ni41  &  ni40 ) | ( ni41  &  (~ ni40) ) | ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( (~ ni41)  &  ni40  &  ni44 ) ;
 assign n_n2280 = ( wire35286 ) | ( (~ ni36)  &  wire35122 ) | ( (~ ni36)  &  wire35123 ) ;
 assign n_n1329 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n2228 ) ;
 assign wire1104 = ( ni43  &  ni40 ) | ( ni42  &  ni40 ) | ( (~ ni43)  &  ni40  &  ni45 ) ;
 assign n_n2229 = ( wire35288 ) | ( (~ nv539)  &  wire35108 ) | ( (~ nv539)  &  wire35109 ) ;
 assign wire771 = ( ni47 ) | ( (~ ni43)  &  ni42 ) ;
 assign wire934 = ( ni43 ) | ( ni42 ) | ( ni45 ) ;
 assign nv9050 = ( ni43 ) | ( ni42 ) | ( (~ ni43)  &  ni45 ) ;
 assign n_n2143 = ( wire35274 ) | ( nv9492  &  wire35273 ) | ( wire1777  &  wire35273 ) ;
 assign wire1250 = ( ni36  &  ni32  &  (~ wire172) ) | ( ni36  &  ni32  &  nv9050 ) ;
 assign wire1196 = ( wire1763 ) | ( nv9066  &  wire266 ) ;
 assign n_n1891 = ( (~ ni40)  &  ni38  &  wire907 ) | ( ni40  &  ni38  &  nv9031 ) | ( (~ ni40)  &  ni38  &  nv9031 ) ;
 assign wire1212 = ( (~ ni38)  &  ni37  &  (~ ni36) ) | ( (~ ni38)  &  (~ ni36)  &  n_n1984 ) ;
 assign n_n1410 = ( wire1212 ) | ( wire1585 ) | ( (~ ni36)  &  n_n1891 ) ;
 assign wire835 = ( ni36  &  (~ ni32) ) | ( ni35  &  (~ ni32) ) ;
 assign n_n1394 = ( wire35031 ) | ( (~ ni35)  &  (~ ni32)  &  n_n1410 ) ;
 assign n_n1858 = ( wire589 ) | ( wire1578 ) | ( wire1579 ) | ( wire1580 ) ;
 assign wire836 = ( ni36  &  (~ ni32) ) | ( (~ ni35)  &  (~ ni32) ) ;
 assign wire242 = ( (~ ni38)  &  ni37 ) | ( (~ ni38)  &  (~ ni37)  &  wire770 ) ;
 assign wire974 = ( wire1992 ) | ( wire348  &  wire701 ) ;
 assign n_n12782 = ( wire500 ) | ( wire292  &  nv628 ) ;
 assign nv658 = ( ni34 ) | ( (~ wire157)  &  (~ wire6663)  &  (~ wire29629) ) ;
 assign wire1310 = ( ni34  &  wire6663 ) | ( ni34  &  wire6664 ) | ( ni34  &  wire29628 ) ;
 assign nv1052 = ( wire184 ) | ( (~ nv6428)  &  nv658 ) | ( nv662  &  nv658 ) ;
 assign nv764 = ( ni34 ) | ( (~ wire157)  &  (~ n_n12696)  &  (~ wire29518) ) ;
 assign wire1070 = ( ni34  &  n_n12696 ) | ( ni34  &  wire29518 ) ;
 assign n_n10809 = ( wire5851 ) | ( wire5852 ) | ( n_n10860  &  wire881 ) ;
 assign nv2602 = ( n_n10590 ) | ( ni41  &  n_n11266 ) | ( ni41  &  wire5930 ) ;
 assign nv2694 = ( wire5648 ) | ( wire30675 ) | ( (~ ni36)  &  nv2995 ) ;
 assign nv2276 = ( wire5507 ) | ( wire30499 ) | ( (~ ni36)  &  nv2493 ) ;
 assign nv2220 = ( wire706 ) | ( wire5924 ) | ( wire5926 ) | ( wire30431 ) ;
 assign nv2641 = ( wire5632 ) | ( wire30659 ) | ( (~ ni36)  &  nv2963 ) ;
 assign n_n10412 = ( wire1195 ) | ( wire400  &  nv2602 ) ;
 assign wire219 = ( (~ pi20)  &  pi25  &  wire153 ) ;
 assign wire303 = ( (~ ni33)  &  (~ ni32)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire313 = ( (~ pi25)  &  wire303 ) ;
 assign wire572 = ( wire5453 ) | ( (~ wire150)  &  wire5454 ) | ( (~ wire150)  &  wire5455 ) ;
 assign wire697 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire953 = ( wire378 ) | ( wire152  &  wire5454 ) | ( wire152  &  wire5455 ) ;
 assign wire432 = ( wire5450 ) | ( wire228  &  n_n9304 ) | ( wire228  &  wire5816 ) ;
 assign wire983 = ( wire5448 ) | ( wire325  &  wire5454 ) | ( wire325  &  wire5455 ) ;
 assign wire1043 = ( pi21  &  pi22  &  (~ pi25)  &  wire303 ) ;
 assign wire1080 = ( pi19  &  pi21  &  pi22  &  pi25 ) ;
 assign n_n10795 = ( wire5439 ) | ( wire5440 ) | ( wire31005 ) ;
 assign wire1188 = ( ni36  &  wire216 ) | ( wire347  &  nv2647 ) ;
 assign wire794 = ( wire432 ) | ( wire169  &  wire5454 ) | ( wire169  &  wire5455 ) ;
 assign n_n10796 = ( wire5348 ) | ( wire5351 ) | ( wire30976 ) | ( wire30977 ) ;
 assign wire1013 = ( wire176  &  wire216 ) | ( (~ ni37)  &  wire176  &  n_n10282 ) ;
 assign wire1195 = ( (~ ni36)  &  wire216 ) | ( wire404  &  n_n10282 ) ;
 assign wire885 = ( ni40 ) | ( wire216 ) | ( ni39  &  n_n10282 ) ;
 assign nv2430 = ( wire240 ) | ( ni33  &  wire5429 ) | ( ni33  &  wire30473 ) ;
 assign wire1186 = ( ni36  &  wire216 ) | ( nv2240  &  wire346 ) ;
 assign n_n9177 = ( wire4868 ) | ( ni40  &  ni38  &  nv3943 ) ;
 assign n_n7913 = ( n_n6710 ) | ( wire206  &  (~ wire4953)  &  (~ wire31516) ) ;
 assign n_n7877 = ( n_n6710 ) | ( wire206  &  (~ wire323)  &  (~ wire4917) ) ;
 assign n_n7893 = ( n_n6710 ) | ( wire206  &  (~ wire4887)  &  (~ wire31176) ) ;
 assign wire329 = ( pi17  &  wire180 ) ;
 assign wire460 = ( pi17  &  wire178 ) ;
 assign wire1003 = ( pi17  &  wire170 ) | ( (~ wire150)  &  wire31935 ) ;
 assign wire475 = ( (~ pi17)  &  pi25  &  wire179 ) ;
 assign wire611 = ( pi21  &  pi22  &  pi20  &  pi25 ) ;
 assign wire505 = ( wire32110 ) | ( wire305  &  wire199 ) | ( wire199  &  wire4562 ) ;
 assign nv4389 = ( wire305 ) | ( wire233  &  wire4681 ) | ( wire233  &  wire31852 ) ;
 assign wire502 = ( wire391 ) | ( wire305  &  wire203 ) | ( wire203  &  wire4533 ) ;
 assign wire198 = ( (~ pi17)  &  (~ pi19) ) | ( (~ pi17)  &  pi20 ) ;
 assign wire449 = ( (~ pi20)  &  nv4401  &  wire153 ) | ( pi20  &  wire153  &  nv4409 ) ;
 assign wire185 = ( (~ pi17)  &  (~ pi19) ) | ( (~ pi17)  &  (~ pi20) ) ;
 assign wire850 = ( (~ pi19)  &  wire170 ) ;
 assign n_n8956 = ( wire4889 ) | ( wire4890 ) | ( wire4891 ) ;
 assign n_n9157 = ( wire4892 ) | ( (~ ni40)  &  ni38  &  nv3927 ) ;
 assign wire187 = ( (~ wire156)  &  n_n8085 ) | ( ni32  &  ni30  &  wire156 ) ;
 assign wire372 = ( n_n7095 ) | ( (~ pi22)  &  nv4938  &  wire204 ) ;
 assign wire960 = ( wire4226 ) | ( wire158  &  wire152  &  wire274 ) ;
 assign wire442 = ( n_n7095 ) | ( (~ pi22)  &  wire211  &  nv4938 ) ;
 assign wire393 = ( pi17  &  pi25  &  (~ pi16)  &  wire152 ) ;
 assign nv5283 = ( pi27  &  ni32 ) | ( (~ pi26)  &  ni32 ) | ( (~ pi27)  &  pi26  &  wire775 ) ;
 assign n_n6749 = ( (~ pi21)  &  ni32  &  wire155 ) | ( (~ pi21)  &  (~ wire155)  &  wire775 ) ;
 assign wire424 = ( ni32  &  (~ ni30) ) | ( ni32  &  ni31  &  ni30 ) | ( ni33  &  ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire1284 = ( (~ pi21)  &  wire424 ) ;
 assign n_n5908 = ( (~ pi21)  &  ni32  &  wire160 ) | ( (~ pi21)  &  (~ wire160)  &  wire424 ) ;
 assign n_n5604 = ( wire1198 ) | ( wire3497 ) ;
 assign wire276 = ( pi25  &  nv7791 ) | ( (~ pi25)  &  wire3157 ) | ( (~ pi25)  &  wire3158 ) ;
 assign wire906 = ( wire311  &  wire3193 ) | ( n_n4404  &  wire477  &  wire311 ) ;
 assign wire963 = ( wire2214 ) | ( wire152  &  wire154  &  wire276 ) ;
 assign wire1298 = ( wire219  &  wire3206 ) | ( (~ n_n5520)  &  wire219  &  wire33611 ) ;
 assign wire1311 = ( wire358  &  wire3393 ) | ( wire358  &  n_n4441  &  wire33555 ) ;
 assign wire527 = ( pi20  &  nv7050  &  wire153 ) | ( (~ pi20)  &  wire153  &  nv7043 ) ;
 assign nv7043 = ( wire196 ) | ( wire192  &  wire3326 ) | ( wire192  &  wire3327 ) ;
 assign wire672 = ( wire34203 ) | ( nv10153  &  wire2498 ) | ( nv10153  &  wire34198 ) ;
 assign wire832 = ( (~ pi17)  &  pi27  &  wire179 ) ;
 assign wire734 = ( (~ pi21)  &  pi20  &  nv7791 ) | ( pi21  &  (~ pi22)  &  pi20  &  nv7791 ) ;
 assign wire1306 = ( (~ pi21)  &  nv7791  &  wire185 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire185 ) ;
 assign nv6797 = ( wire197 ) | ( wire193  &  wire3307 ) | ( wire193  &  wire3308 ) ;
 assign wire1068 = ( (~ ni40)  &  (~ ni37)  &  wire3491 ) | ( (~ ni40)  &  (~ ni37)  &  wire33310 ) ;
 assign wire1123 = ( ni40  &  (~ ni37)  &  wire3491 ) | ( ni40  &  (~ ni37)  &  wire33310 ) ;
 assign wire465 = ( n_n2328 ) | ( (~ wire426)  &  wire253 ) | ( wire253  &  nv669 ) ;
 assign wire798 = ( wire463 ) | ( (~ ni40)  &  ni38  &  nv6486 ) ;
 assign wire468 = ( n_n2328 ) | ( (~ ni40)  &  ni38  &  nv669 ) ;
 assign wire385 = ( pi20  &  nv6859  &  wire153 ) | ( (~ pi20)  &  wire153  &  nv6851 ) ;
 assign wire507 = ( (~ pi17)  &  pi16  &  (~ pi15) ) ;
 assign wire1011 = ( pi19  &  (~ pi21)  &  ni30 ) | ( pi19  &  pi21  &  (~ pi22)  &  ni30 ) ;
 assign wire912 = ( pi21  &  pi22  &  wire268 ) ;
 assign nv8350 = ( wire34814 ) | ( (~ ni11)  &  wire3177 ) | ( (~ ni11)  &  wire33906 ) ;
 assign n_n2546 = ( wire2881 ) | ( nv8372  &  wire34844 ) ;
 assign wire337 = ( wire2878 ) | ( wire2881 ) | ( nv8372  &  wire34844 ) ;
 assign nv6886 = ( wire197 ) | ( wire193  &  wire3185 ) | ( wire193  &  wire3186 ) ;
 assign wire409 = ( ni41 ) | ( (~ ni41)  &  (~ ni44) ) | ( (~ ni41)  &  wire934 ) ;
 assign n_n2452 = ( wire1881 ) | ( (~ ni38)  &  ni37 ) ;
 assign wire1249 = ( ni36  &  wire266 ) | ( wire266  &  wire33267 ) | ( (~ ni36)  &  wire266  &  n_n5799 ) ;
 assign n_n5799 = ( ni39  &  ni47 ) | ( ni39  &  ni45 ) ;
 assign n_n2226 = ( wire35292 ) | ( wire316  &  wire6742 ) | ( wire316  &  wire29648 ) ;
 assign n_n1395 = ( wire35034 ) | ( wire461  &  wire1602 ) | ( wire461  &  wire35033 ) ;
 assign nv9297 = ( wire2005 ) | ( wire4913 ) | ( (~ ni41)  &  ni44 ) ;
 assign n_n1859 = ( wire35243 ) | ( (~ nv539)  &  n_n1395 ) | ( n_n1395  &  wire35242 ) ;
 assign n_n1558 = ( wire1022 ) | ( wire999  &  wire951 ) | ( wire951  &  wire1941 ) ;
 assign n_n1229 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n1558 ) ;
 assign wire239 = ( ni4 ) | ( ni5 ) ;
 assign nv683 = ( wire436 ) | ( wire6678 ) | ( wire6679 ) | ( wire6680 ) ;
 assign nv1009 = ( wire184 ) | ( (~ nv6428)  &  nv620 ) | ( nv620  &  nv624 ) ;
 assign nv679 = ( ni34 ) | ( (~ wire157)  &  (~ wire6680)  &  (~ wire29636) ) ;
 assign wire1057 = ( ni34  &  wire6678 ) | ( ni34  &  wire6680 ) | ( ni34  &  wire29635 ) ;
 assign nv1073 = ( wire184 ) | ( (~ nv6428)  &  nv679 ) | ( nv683  &  nv679 ) ;
 assign wire617 = ( pi19  &  pi21  &  pi20 ) ;
 assign wire843 = ( pi21  &  pi20  &  wire344 ) ;
 assign wire1293 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire1014 = ( pi19  &  (~ pi20)  &  pi25 ) ;
 assign wire1108 = ( pi19  &  (~ pi21)  &  ni34 ) | ( pi19  &  (~ pi22)  &  ni34 ) ;
 assign nv821 = ( wire436 ) | ( wire6556 ) | ( wire6557 ) | ( wire6558 ) ;
 assign nv817 = ( ni34 ) | ( (~ wire157)  &  (~ wire6557)  &  (~ wire29588) ) ;
 assign wire1318 = ( ni34  &  wire6557 ) | ( ni34  &  wire6558 ) | ( ni34  &  wire29587 ) ;
 assign wire887 = ( ni40 ) | ( wire216 ) | ( wire5798 ) ;
 assign wire338 = ( wire4394 ) | ( (~ pi24)  &  wire170 ) | ( pi24  &  wire1284 ) ;
 assign nv6146 = ( wire338 ) | ( wire4392 ) | ( (~ pi24)  &  wire1118 ) ;
 assign nv5862 = ( wire339 ) | ( wire4327 ) | ( wire161  &  wire1118 ) ;
 assign wire339 = ( n_n6410 ) | ( pi21  &  wire4383 ) | ( pi21  &  wire4384 ) ;
 assign wire555 = ( ni13  &  (~ ni11) ) | ( (~ ni14)  &  (~ ni11)  &  (~ ni12) ) ;
 assign nv6124 = ( n_n6367 ) | ( pi27  &  wire1065 ) | ( (~ pi27)  &  wire1065 ) | ( (~ pi27)  &  wire4397 ) ;
 assign n_n7400 = ( wire3719 ) | ( wire3720 ) | ( wire3721 ) | ( wire33052 ) ;
 assign wire793 = ( ni9 ) | ( (~ ni10) ) | ( ni8 ) ;
 assign wire833 = ( ni11  &  (~ ni9)  &  (~ ni10)  &  (~ ni8) ) ;
 assign wire964 = ( wire3706 ) | ( wire158  &  wire152  &  wire280 ) ;
 assign wire1316 = ( (~ ni9)  &  (~ ni10)  &  (~ ni8) ) ;
 assign n_n8112 = ( wire3667 ) | ( wire3668 ) | ( wire3670 ) | ( wire33220 ) ;
 assign wire330 = ( ni11  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire359 = ( (~ ni13)  &  ni14  &  (~ ni11)  &  ni12 ) ;
 assign wire401 = ( ni13 ) | ( ni12 ) | ( (~ ni13)  &  (~ ni14)  &  (~ ni12) ) ;
 assign wire914 = ( pi21  &  (~ pi22) ) ;
 assign wire838 = ( pi26  &  (~ pi24) ) ;
 assign wire1303 = ( ni13  &  (~ ni11) ) ;
 assign nv6104 = ( n_n6710 ) | ( pi27  &  wire1065 ) | ( (~ pi27)  &  wire1065 ) | ( pi27  &  wire4397 ) ;
 assign nv6110 = ( n_n6367 ) | ( pi27  &  wire1065 ) | ( (~ pi27)  &  wire1065 ) | ( pi27  &  wire4397 ) ;
 assign n_n6711 = ( ni32  &  ni31  &  ni30 ) | ( ni33  &  ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire684 = ( wire32184 ) | ( (~ wire150)  &  n_n6710 ) | ( (~ wire150)  &  wire4973 ) ;
 assign wire1256 = ( wire32334 ) | ( (~ pi15)  &  wire32318 ) | ( (~ pi15)  &  wire32319 ) ;
 assign nv6289 = ( wire334 ) | ( wire3596 ) | ( wire160  &  wire1118 ) ;
 assign wire334 = ( n_n5908 ) | ( pi21  &  wire3601 ) | ( pi21  &  wire3602 ) ;
 assign wire574 = ( (~ ni14) ) | ( ni12 ) | ( ni13  &  ni14 ) ;
 assign wire1283 = ( (~ pi17)  &  pi23  &  (~ pi24)  &  wire182 ) ;
 assign wire1328 = ( (~ ni9)  &  ni10  &  (~ ni7)  &  ni8 ) ;
 assign wire871 = ( (~ ni36)  &  (~ wire255) ) | ( nv3915  &  wire31172 ) ;
 assign wire928 = ( n_n6710 ) | ( wire436  &  wire206  &  (~ n_n9022) ) ;
 assign nv6851 = ( wire197 ) | ( wire193  &  wire3205 ) | ( wire193  &  wire3206 ) ;
 assign wire204 = ( pi21  &  (~ pi20) ) ;
 assign wire529 = ( wire34078 ) | ( nv10153  &  wire2402 ) | ( nv10153  &  wire2403 ) ;
 assign wire1096 = ( (~ pi17)  &  pi27  &  wire182 ) | ( (~ pi17)  &  pi26  &  wire182 ) ;
 assign wire1102 = ( (~ pi17)  &  (~ pi27)  &  (~ pi26)  &  wire182 ) ;
 assign wire446 = ( pi20  &  nv7105  &  wire153 ) | ( (~ pi20)  &  wire153  &  nv7098 ) ;
 assign wire640 = ( wire446 ) | ( wire196  &  wire199 ) | ( wire199  &  wire2469 ) ;
 assign wire657 = ( wire34175 ) | ( nv10153  &  wire2446 ) | ( nv10153  &  wire34170 ) ;
 assign wire1035 = ( pi17  &  (~ pi21)  &  ni30 ) | ( pi17  &  pi21  &  (~ pi22)  &  ni30 ) ;
 assign wire1340 = ( (~ pi17)  &  (~ pi19)  &  pi16 ) ;
 assign wire915 = ( pi17  &  pi19  &  pi16  &  pi15 ) | ( (~ pi17)  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire685 = ( ni40  &  ni38  &  ni36 ) | ( ni40  &  (~ ni37)  &  ni36 ) ;
 assign wire447 = ( (~ pi20)  &  nv6789  &  wire153 ) | ( pi20  &  wire153  &  nv6797 ) ;
 assign wire528 = ( wire2980 ) | ( wire34482 ) | ( nv10167  &  wire447 ) ;
 assign n_n1341 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n2332 ) ;
 assign n_n1427 = ( wire34997 ) | ( wire461  &  wire2050 ) | ( wire461  &  wire34996 ) ;
 assign n_n1908 = ( wire35215 ) | ( (~ nv539)  &  n_n1427 ) | ( n_n1427  &  wire35214 ) ;
 assign n_n1426 = ( wire35000 ) | ( wire2040  &  wire34999 ) | ( wire34998  &  wire34999 ) ;
 assign wire783 = ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( (~ ni41)  &  (~ ni40)  &  (~ ni44)  &  (~ nv9031) ) ;
 assign n_n1907 = ( wire35218 ) | ( (~ ni36)  &  n_n1426 ) | ( n_n1426  &  wire35217 ) ;
 assign n_n1905 = ( wire1648 ) | ( wire35221 ) | ( wire245  &  n_n1908 ) ;
 assign n_n1494 = ( wire35043 ) | ( wire2101  &  wire35042 ) | ( wire35041  &  wire35042 ) ;
 assign n_n1219 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n1494 ) ;
 assign n_n1495 = ( wire35040 ) | ( nv590  &  wire2081 ) | ( nv590  &  wire35039 ) ;
 assign wire975 = ( wire2072 ) | ( wire701  &  wire349 ) ;
 assign n_n1491 = ( wire35046 ) | ( wire316  &  wire6581 ) | ( wire316  &  wire29504 ) ;
 assign wire948 = ( (~ ni11)  &  (~ ni12) ) | ( (~ pi27)  &  ni14  &  (~ ni11) ) ;
 assign wire714 = ( (~ nv6428) ) | ( wire29562 ) | ( (~ ni36)  &  nv858 ) ;
 assign nv1291 = ( wire184 ) | ( ni34  &  wire714 ) | ( wire714  &  wire6524 ) ;
 assign nv779 = ( ni34 ) | ( (~ wire157)  &  (~ wire6577)  &  (~ wire29569) ) ;
 assign wire1282 = ( ni34  &  wire6577 ) | ( ni34  &  wire6578 ) | ( ni34  &  wire29568 ) ;
 assign nv1183 = ( wire184 ) | ( (~ nv6428)  &  nv764 ) | ( nv768  &  nv764 ) ;
 assign nv1226 = ( wire184 ) | ( (~ nv6428)  &  nv797 ) | ( nv801  &  nv797 ) ;
 assign nv1205 = ( wire184 ) | ( (~ nv6428)  &  nv779 ) | ( nv779  &  nv783 ) ;
 assign nv1270 = ( wire184 ) | ( (~ nv6428)  &  nv835 ) | ( nv839  &  nv835 ) ;
 assign nv835 = ( ni34 ) | ( (~ wire157)  &  (~ wire6537)  &  (~ wire29593) ) ;
 assign nv1249 = ( wire184 ) | ( (~ nv6428)  &  nv817 ) | ( nv821  &  nv817 ) ;
 assign wire1112 = ( ni34  &  wire6537 ) | ( ni34  &  wire6538 ) | ( ni34  &  wire29592 ) ;
 assign nv783 = ( wire436 ) | ( wire6576 ) | ( wire6577 ) | ( wire6578 ) ;
 assign wire586 = ( pi17  &  pi16  &  (~ pi15)  &  wire152 ) ;
 assign wire614 = ( pi17  &  pi16  &  (~ pi15) ) ;
 assign wire1071 = ( pi17  &  pi19  &  pi16  &  (~ pi15) ) ;
 assign wire1210 = ( wire816 ) | ( pi25  &  wire326  &  wire184 ) ;
 assign nv997 = ( ni34 ) | ( (~ wire157)  &  (~ nv858) ) ;
 assign wire1058 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire1066 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire1183 = ( ni36  &  wire216 ) | ( wire347  &  nv2240 ) ;
 assign wire886 = ( ni40 ) | ( wire216 ) | ( (~ ni39)  &  n_n10282 ) ;
 assign wire883 = ( (~ ni40) ) | ( wire216 ) | ( ni39  &  n_n10282 ) ;
 assign n_n8968 = ( wire4864 ) | ( wire4865 ) | ( wire4866 ) ;
 assign nv4327 = ( wire305 ) | ( wire233  &  wire4613 ) | ( wire233  &  wire31347 ) ;
 assign n_n4697 = ( wire34724 ) | ( (~ ni11)  &  wire33860 ) | ( (~ ni11)  &  wire33861 ) ;
 assign wire1150 = ( wire34032 ) | ( wire34033 ) | ( wire34059 ) | ( wire34060 ) ;
 assign n_n4834 = ( wire3109 ) | ( wire3110 ) | ( wire180  &  n_n4412 ) ;
 assign n_n4934 = ( wire2318 ) | ( wire2323 ) | ( wire33715 ) | ( wire33716 ) ;
 assign wire1091 = ( pi19  &  ni30 ) ;
 assign n_n5328 = ( wire2730 ) | ( wire2731 ) | ( wire2732 ) | ( wire33839 ) ;
 assign wire371 = ( wire3057 ) | ( wire173  &  wire616 ) ;
 assign wire433 = ( wire3084 ) | ( wire3085 ) | ( wire173  &  wire340 ) ;
 assign wire585 = ( wire3069 ) | ( pi17  &  pi16  &  wire443 ) ;
 assign wire1291 = ( pi20  &  wire351 ) ;
 assign wire899 = ( wire3086 ) | ( pi25  &  (~ pi16) ) ;
 assign wire1206 = ( wire906 ) | ( wire476  &  wire3064 ) | ( wire476  &  wire33705 ) ;
 assign n_n5713 = ( wire707 ) | ( wire3303 ) | ( nv6486  &  wire691 ) ;
 assign wire273 = ( pi25  &  nv7445 ) | ( (~ pi25)  &  wire3139 ) | ( (~ pi25)  &  wire3140 ) ;
 assign wire959 = ( wire2798 ) | ( wire158  &  wire152  &  wire273 ) ;
 assign wire1285 = ( pi25  &  wire158  &  wire152  &  n_n4611 ) ;
 assign wire1326 = ( wire345  &  wire3280 ) | ( wire345  &  n_n4489  &  wire33307 ) ;
 assign wire422 = ( (~ pi27)  &  ni33  &  ni30 ) | ( pi27  &  ni31  &  ni30 ) | ( (~ pi27)  &  ni31  &  ni30 ) ;
 assign wire597 = ( (~ pi21)  &  nv7647 ) | ( (~ pi22)  &  nv7647 ) ;
 assign wire921 = ( (~ pi21)  &  (~ ni14) ) | ( (~ pi22)  &  (~ ni14) ) ;
 assign wire837 = ( pi21  &  pi22  &  (~ ni14) ) ;
 assign nv8777 = ( wire337 ) | ( wire2852 ) | ( wire160  &  wire1063 ) ;
 assign n_n1311 = ( wire308 ) | ( (~ pi21)  &  wire999 ) | ( (~ pi21)  &  wire1941 ) ;
 assign nv9262 = ( wire2087 ) | ( wire4971 ) | ( (~ ni41)  &  (~ ni44) ) ;
 assign n_n2097 = ( wire1927 ) | ( wire35228 ) | ( wire35229 ) ;
 assign n_n2009 = ( wire35204 ) | ( (~ ni36)  &  n_n1494 ) | ( n_n1494  &  wire35203 ) ;
 assign n_n2010 = ( wire35202 ) | ( (~ ni36)  &  n_n1495 ) | ( (~ ni32)  &  n_n1495 ) ;
 assign n_n2007 = ( wire35208 ) | ( wire316  &  wire6577 ) | ( wire316  &  wire29569 ) ;
 assign n_n1301 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n2009 ) ;
 assign nv1556 = ( wire184 ) | ( (~ nv6428)  &  nv979 ) | ( nv983  &  nv979 ) ;
 assign nv1577 = ( wire184 ) | ( (~ nv6428)  &  nv988 ) | ( nv992  &  nv988 ) ;
 assign wire1045 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire1073 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign nv1403 = ( wire184 ) | ( (~ nv6428)  &  nv910 ) | ( nv914  &  nv910 ) ;
 assign wire248 = ( pi25  &  nv7647 ) | ( (~ pi25)  &  wire3125 ) | ( (~ pi25)  &  wire3126 ) ;
 assign wire575 = ( wire2688 ) | ( wire153  &  wire248 ) ;
 assign wire739 = ( wire3060 ) | ( wire219  &  wire3205 ) | ( wire219  &  wire3206 ) ;
 assign wire1016 = ( ni11  &  wire369 ) ;
 assign wire1093 = ( (~ pi17)  &  (~ pi27)  &  pi26  &  wire179 ) ;
 assign wire1094 = ( ni11  &  wire370 ) ;
 assign wire1120 = ( (~ pi17)  &  pi27  &  wire179 ) | ( (~ pi17)  &  (~ pi26)  &  wire179 ) ;
 assign wire962 = ( wire2197 ) | ( wire158  &  wire152  &  wire276 ) ;
 assign n_n4096 = ( wire2168 ) | ( wire33977 ) | ( wire33978 ) | ( wire33979 ) ;
 assign wire918 = ( pi25  &  wire152  &  n_n4404  &  wire154 ) ;
 assign wire1297 = ( wire345  &  wire721  &  wire33433 ) | ( wire345  &  wire721  &  wire33434 ) ;
 assign wire1320 = ( wire1006  &  (~ n_n5520)  &  wire219 ) | ( (~ n_n5520)  &  wire219  &  wire33612 ) ;
 assign n_n1347 = ( wire308 ) | ( (~ pi21)  &  wire1000 ) | ( (~ pi21)  &  wire1710 ) ;
 assign n_n1173 = ( wire35314 ) | ( wire213  &  wire1832 ) | ( wire213  &  wire35312 ) ;
 assign n_n1351 = ( wire308 ) | ( (~ pi21)  &  wire999 ) | ( (~ pi21)  &  wire1883 ) ;
 assign wire1275 = ( wire35329 ) | ( wire863  &  wire35328 ) ;
 assign n_n1335 = ( wire405 ) | ( (~ pi22)  &  wire1896 ) | ( (~ pi22)  &  wire35284 ) ;
 assign wire863 = ( ni32  &  wire35162 ) | ( ni36  &  ni32  &  n_n2452 ) | ( (~ ni36)  &  ni32  &  n_n2452 ) ;
 assign wire349 = ( wire33267 ) | ( ni36  &  nv9066 ) | ( (~ ni36)  &  n_n5799 ) ;
 assign n_n1423 = ( wire35003 ) | ( wire316  &  wire6561 ) | ( wire316  &  wire29526 ) ;
 assign n_n1207 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n1426 ) ;
 assign wire878 = ( wire2035 ) | ( (~ ni35)  &  wire266  &  wire349 ) ;
 assign nv899 = ( ni34 ) | ( (~ wire157)  &  (~ wire6683)  &  (~ wire29470) ) ;
 assign wire1033 = ( ni34  &  wire1097 ) | ( ni34  &  wire6682 ) | ( ni34  &  wire6683 ) ;
 assign nv1380 = ( wire184 ) | ( (~ nv6428)  &  nv899 ) | ( nv903  &  nv899 ) ;
 assign wire943 = ( wire157 ) | ( wire6453 ) | ( wire6454 ) | ( wire29476 ) ;
 assign nv2290 = ( wire240 ) | ( ni33  &  wire5501 ) | ( ni33  &  wire30496 ) ;
 assign nv2411 = ( wire240 ) | ( ni33  &  wire5409 ) | ( ni33  &  wire30467 ) ;
 assign wire200 = ( wire164 ) | ( wire5678 ) | ( wire866  &  wire30522 ) ;
 assign wire916 = ( (~ pi20)  &  n_n9304 ) | ( pi21  &  (~ pi20)  &  n_n9302 ) ;
 assign wire1348 = ( pi20  &  wire162 ) ;
 assign wire486 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire213 ) ;
 assign wire687 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire189 ) ;
 assign wire162 = ( n_n9304 ) | ( wire5816 ) | ( pi21  &  n_n9294 ) ;
 assign wire968 = ( wire294  &  wire200 ) | ( wire697  &  wire162 ) ;
 assign wire1128 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire152 ) ;
 assign wire492 = ( (~ wire255) ) | ( ni39  &  (~ ni38)  &  nv3916 ) ;
 assign wire375 = ( n_n8085 ) | ( wire4061 ) | ( (~ n_n8352)  &  wire31171 ) ;
 assign nv4630 = ( wire374 ) | ( wire214  &  wire4681 ) | ( wire214  &  wire31852 ) ;
 assign wire390 = ( ni37 ) | ( ni38  &  (~ ni37) ) ;
 assign wire592 = ( (~ ni37)  &  wire3491 ) | ( (~ ni37)  &  wire33310 ) ;
 assign n_n1462 = ( wire35012 ) | ( ni35  &  (~ ni32)  &  n_n1478 ) ;
 assign n_n1463 = ( wire34991 ) | ( nv590  &  wire1999 ) | ( nv590  &  wire34990 ) ;
 assign wire972 = ( wire1571 ) | ( wire329  &  wire1574 ) | ( wire329  &  wire35247 ) ;
 assign wire997 = ( wire1563 ) | ( wire458  &  wire308 ) | ( wire458  &  wire1569 ) ;
 assign wire971 = ( wire1471 ) | ( wire329  &  wire1473 ) | ( wire329  &  wire35144 ) ;
 assign wire1262 = ( wire35098 ) | ( wire294  &  wire1454 ) | ( wire294  &  wire35097 ) ;
 assign n_n1277 = ( wire1439 ) | ( wire1444 ) | ( wire35407 ) | ( wire35408 ) ;
 assign n_n1555 = ( wire35063 ) | ( wire316  &  nv942 ) ;
 assign n_n1528 = ( wire1022 ) | ( wire952  &  wire1000 ) | ( wire952  &  wire1631 ) ;
 assign wire695 = ( pi17  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire970 = ( wire1382 ) | ( wire329  &  wire1384 ) | ( wire329  &  wire35037 ) ;
 assign wire995 = ( wire1374 ) | ( wire458  &  wire308 ) | ( wire458  &  wire1380 ) ;
 assign wire328 = ( pi17  &  (~ ni29)  &  wire152 ) | ( pi17  &  (~ ni29)  &  wire189 ) ;
 assign n_n6828 = ( wire3756 ) | ( wire3757 ) | ( wire33036 ) | ( wire33040 ) ;
 assign wire306 = ( n_n6711 ) | ( wire4581 ) | ( (~ n_n8862)  &  wire32057 ) ;
 assign wire1200 = ( wire270  &  n_n2328 ) | ( nv669  &  wire691 ) ;
 assign wire230 = ( (~ pi21)  &  ni34 ) | ( pi21  &  (~ pi22)  &  ni34 ) ;
 assign wire913 = ( pi17  &  pi19  &  pi16  &  (~ pi15) ) | ( (~ pi17)  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire1324 = ( pi20  &  pi16  &  (~ pi15)  &  wire153 ) ;
 assign wire1327 = ( (~ pi20)  &  pi16  &  (~ pi15)  &  wire153 ) ;
 assign wire691 = ( (~ ni40)  &  ni38  &  ni36 ) | ( (~ ni40)  &  (~ ni37)  &  ni36 ) ;
 assign wire707 = ( ni37  &  ni36  &  n_n2328 ) ;
 assign wire1198 = ( wire270  &  n_n2328 ) | ( nv669  &  wire685 ) ;
 assign wire463 = ( n_n2328 ) | ( (~ wire426)  &  wire254 ) | ( wire254  &  nv669 ) ;
 assign wire351 = ( (~ pi21)  &  ni30 ) | ( pi21  &  (~ pi22)  &  ni30 ) | ( pi21  &  pi22  &  pi25  &  ni30 ) ;
 assign wire727 = ( wire3090 ) | ( wire173  &  wire381 ) ;
 assign wire1352 = ( wire393  &  wire3276 ) | ( wire393  &  wire3277 ) ;
 assign wire1213 = ( wire388  &  wire293 ) | ( nv9066  &  wire266 ) ;
 assign n_n1289 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n1907 ) ;
 assign n_n1824 = ( wire1250 ) | ( (~ nv539)  &  wire1772 ) | ( (~ nv539)  &  wire1773 ) ;
 assign n_n1823 = ( wire35184 ) | ( (~ ni36)  &  (~ ni32)  &  nv9492 ) ;
 assign n_n1269 = ( wire35004 ) | ( wire35005 ) | ( (~ pi21)  &  n_n1786 ) ;
 assign n_n1783 = ( wire35167 ) | ( wire245  &  wire863 ) | ( wire245  &  wire35164 ) ;
 assign wire1264 = ( wire7099 ) | ( wire28825 ) | ( wire28826 ) | ( wire28829 ) ;
 assign wire1126 = ( (~ ni40)  &  (~ ni38)  &  (~ ni37) ) ;
 assign n_n11474 = ( wire317 ) | ( wire6249 ) | ( nv959  &  wire29508 ) ;
 assign nv1490 = ( wire184 ) | ( ni34  &  (~ nv6428) ) | ( ni34  &  nv952 ) ;
 assign nv1359 = ( wire184 ) | ( (~ nv6428)  &  nv890 ) | ( nv894  &  nv890 ) ;
 assign n_n4541 = ( wire2772 ) | ( wire2777 ) | ( wire34665 ) | ( wire34666 ) ;
 assign n_n4542 = ( wire2753 ) | ( wire2755 ) | ( wire34638 ) | ( wire34640 ) ;
 assign wire732 = ( (~ pi21)  &  pi20  &  nv7445 ) | ( pi21  &  (~ pi22)  &  pi20  &  nv7445 ) ;
 assign wire1337 = ( (~ pi21)  &  nv7445  &  wire185 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire185 ) ;
 assign wire1079 = ( (~ pi15)  &  wire377 ) ;
 assign wire1083 = ( pi15  &  wire377 ) ;
 assign wire926 = ( ni39 ) | ( ni38 ) ;
 assign n_n11833 = ( wire6269 ) | ( wire6271 ) | ( wire29490 ) | ( wire29491 ) ;
 assign n_n11836 = ( wire6226 ) | ( wire6236 ) | ( wire29556 ) | ( wire29561 ) ;
 assign wire368 = ( pi21  &  ni34 ) ;
 assign wire376 = ( pi21  &  pi22  &  ni33  &  (~ ni32) ) ;
 assign wire343 = ( (~ pi21)  &  ni34 ) | ( pi21  &  (~ pi22)  &  ni34 ) | ( pi21  &  pi22  &  (~ pi25)  &  ni34 ) ;
 assign wire812 = ( pi17  &  pi25  &  (~ pi16)  &  wire180 ) ;
 assign wire813 = ( pi17  &  pi25  &  pi16  &  wire180 ) ;
 assign n_n12641 = ( wire30094 ) | ( pi15  &  wire30073 ) | ( pi15  &  wire30074 ) ;
 assign wire947 = ( wire6242 ) | ( wire6243 ) | ( wire29502 ) ;
 assign wire1030 = ( (~ pi20)  &  ni33  &  (~ ni32)  &  wire153 ) ;
 assign nv4575 = ( wire374 ) | ( wire214  &  wire4613 ) | ( wire214  &  wire31347 ) ;
 assign wire740 = ( wire1320 ) | ( wire3104 ) ;
 assign wire957 = ( wire2681 ) | ( wire158  &  wire152  &  wire248 ) ;
 assign wire722 = ( (~ ni43)  &  ni42 ) | ( (~ ni41)  &  ni40 ) ;
 assign n_n9515 = ( wire5616 ) | ( wire5618 ) | ( wire5619 ) | ( wire31101 ) ;
 assign wire903 = ( wire763  &  wire200 ) | ( wire162  &  wire31065 ) ;
 assign n_n9516 = ( wire5535 ) | ( wire5538 ) | ( wire5539 ) | ( wire31082 ) ;
 assign wire443 = ( (~ pi21)  &  ni30 ) | ( (~ pi22)  &  ni30 ) ;
 assign wire754 = ( wire433 ) | ( pi20  &  wire153  &  n_n5481 ) | ( (~ pi20)  &  wire153  &  n_n5481 ) ;
 assign n_n11295 = ( wire31023 ) | ( wire1069  &  n_n10795 ) | ( wire1069  &  n_n10796 ) ;
 assign wire694 = ( wire5247 ) | ( wire5248 ) ;
 assign nv3202 = ( wire304 ) | ( wire240  &  wire252 ) | ( wire252  &  wire5196 ) ;
 assign n_n9647 = ( wire30510 ) | ( wire252  &  wire5184 ) | ( wire252  &  wire30509 ) ;
 assign wire723 = ( wire5145 ) | ( wire5146 ) | ( wire30865 ) | ( wire30866 ) ;
 assign wire852 = ( wire5166 ) | ( wire5168 ) | ( wire5169 ) | ( wire30446 ) ;
 assign wire933 = ( wire5107 ) | ( wire5108 ) | ( wire30819 ) | ( wire30820 ) ;
 assign nv4648 = ( wire374 ) | ( wire214  &  wire4811 ) | ( wire214  &  wire31893 ) ;
 assign wire1178 = ( n_n9245  &  wire151 ) | ( (~ pi19)  &  wire170 ) ;
 assign n_n8343 = ( wire3898 ) | ( wire3904 ) | ( wire31975 ) | ( wire31976 ) ;
 assign n_n7001 = ( wire4024 ) | ( wire4025 ) | ( wire33152 ) | ( wire33156 ) ;
 assign n_n6410 = ( (~ pi21)  &  ni32  &  wire161 ) | ( (~ pi21)  &  (~ wire161)  &  wire424 ) ;
 assign wire599 = ( pi27  &  wire1065 ) | ( (~ pi27)  &  wire1065 ) | ( pi27  &  wire4397 ) ;
 assign wire391 = ( wire4530 ) | ( wire4531 ) | ( wire305  &  wire448 ) ;
 assign wire780 = ( ni40  &  nv9031 ) | ( (~ ni40)  &  nv9031 ) | ( (~ ni41)  &  ni40  &  (~ ni44)  &  (~ nv9031) ) ;
 assign wire1211 = ( (~ ni38)  &  ni37  &  (~ ni36) ) | ( (~ ni38)  &  (~ ni36)  &  n_n2466 ) ;
 assign n_n1992 = ( ni40  &  ni38  &  wire907 ) | ( ni40  &  ni38  &  nv9031 ) | ( (~ ni40)  &  ni38  &  nv9031 ) ;
 assign wire1263 = ( wire1686 ) | ( wire1688 ) | ( wire697  &  n_n1347 ) ;
 assign nv10174 = ( pi27  &  (~ ni30) ) | ( (~ pi27)  &  (~ ni30) ) | ( pi27  &  ni33  &  ni30 ) | ( pi27  &  ni31  &  ni30 ) | ( (~ pi27)  &  ni31  &  ni30 ) ;
 assign nv10178 = ( (~ pi26)  &  (~ ni30) ) | ( pi26  &  nv10173 ) | ( (~ pi26)  &  ni31  &  ni30 ) ;
 assign nv10237 = ( nv10167  &  wire764 ) | ( nv10169  &  wire631  &  (~ wire764) ) ;
 assign wire980 = ( ni13 ) | ( (~ ni14)  &  ni11 ) | ( ni11  &  ni12 ) ;
 assign nv10173 = ( pi27  &  (~ ni30) ) | ( (~ pi27)  &  (~ ni30) ) | ( (~ pi27)  &  ni33  &  ni30 ) | ( pi27  &  ni31  &  ni30 ) | ( (~ pi27)  &  ni31  &  ni30 ) ;
 assign nv10222 = ( (~ ni30)  &  wire160 ) | ( (~ ni30)  &  (~ wire160) ) | ( ni31  &  ni30  &  wire160 ) | ( (~ ni33)  &  ni30  &  (~ wire160) ) | ( ni31  &  ni30  &  (~ wire160) ) ;
 assign nv10162 = ( nv10153 ) | ( (~ pi27)  &  pi26  &  (~ nv10153) ) ;
 assign nv10187 = ( (~ ni30)  &  wire161 ) | ( (~ ni30)  &  (~ wire161) ) | ( ni31  &  ni30  &  wire161 ) | ( (~ ni33)  &  ni30  &  (~ wire161) ) | ( ni31  &  ni30  &  (~ wire161) ) ;
 assign wire493 = ( pi27 ) | ( (~ ni30) ) | ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire628 = ( pi24  &  (~ ni30) ) | ( (~ pi24)  &  (~ ni30) ) | ( pi24  &  (~ ni33)  &  ni30 ) | ( pi24  &  ni31  &  ni30 ) | ( (~ pi24)  &  ni31  &  ni30 ) ;
 assign wire764 = ( (~ ni13)  &  (~ ni11)  &  (~ ni12) ) | ( (~ ni14)  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire868 = ( ni13  &  ni14  &  (~ ni11) ) | ( ni13  &  (~ ni11)  &  ni12 ) ;
 assign n_n983 = ( wire6891 ) | ( wire29352 ) | ( wire29353 ) | ( wire29354 ) ;
 assign wire480 = ( wire764 ) | ( nv10153  &  wire29270 ) | ( (~ wire156)  &  (~ nv10153)  &  wire29270 ) ;
 assign wire1277 = ( ni13  &  nv10167 ) | ( (~ ni12)  &  nv10167 ) | ( nv10167  &  wire29198 ) ;
 assign wire499 = ( pi27 ) | ( (~ pi26) ) | ( wire175 ) | ( nv10153 ) ;
 assign nv10252 = ( wire6822 ) | ( wire6827 ) | ( wire29252 ) | ( wire29253 ) ;
 assign nv4641 = ( wire374 ) | ( wire214  &  wire4805 ) | ( wire214  &  wire31891 ) ;
 assign wire535 = ( pi20  &  wire153  &  nv4648 ) | ( (~ pi20)  &  wire153  &  nv4641 ) ;
 assign n_n1478 = ( wire1212 ) | ( wire2010 ) | ( (~ ni36)  &  n_n1992 ) ;
 assign n_n806 = ( wire6812 ) | ( wire6814 ) | ( nv10237  &  wire29259 ) ;
 assign wire965 = ( wire4082 ) | ( wire152  &  wire154  &  wire280 ) ;
 assign n_n7239 = ( wire3809 ) | ( wire3810 ) | ( wire33087 ) | ( wire33091 ) ;
 assign wire188 = ( (~ wire155)  &  n_n8085 ) | ( ni32  &  ni30  &  wire155 ) ;
 assign wire280 = ( pi25  &  wire188 ) | ( (~ pi25)  &  wire4458 ) | ( (~ pi25)  &  wire4459 ) ;
 assign wire373 = ( n_n6749 ) | ( (~ pi22)  &  wire211  &  nv5285 ) ;
 assign wire440 = ( n_n6749 ) | ( (~ pi22)  &  nv5285  &  wire204 ) ;
 assign wire159 = ( n_n9304 ) | ( pi21  &  n_n9302 ) ;
 assign p__cmx0ad_11 = ( n_n13961 ) ;
 assign p__cmx0ad_33 = ( n_n13961 ) ;
 assign p__cmx0ad_10 = ( n_n13961 ) ;
 assign p__cmx0ad_32 = ( n_n13961 ) ;
 assign p__cmx1ad_8 = ( n_n13961 ) ;
 assign p__cmx0ad_35 = ( n_n13961 ) ;
 assign p__cmx0ad_34 = ( n_n13961 ) ;
 assign p__cmxcl_0 = ( n_n13895 ) ;
 assign p__cmxcl_1 = ( n_n13895 ) ;
 assign p__cmx0ad_8 = ( n_n13961 ) ;
 assign p__cmx1ad_34 = ( n_n13961 ) ;
 assign p__cmx1ad_35 = ( n_n13961 ) ;
 assign p__cmx1ad_32 = ( n_n13961 ) ;
 assign p__cmx1ad_33 = ( n_n13961 ) ;
 assign p__cmx1ad_10 = ( n_n13961 ) ;
 assign p__cmx1ad_11 = ( n_n13961 ) ;
 assign wire168 = ( ni33  &  (~ wire265)  &  wire510 ) | ( (~ ni29)  &  (~ wire265)  &  wire510 ) ;
 assign wire283 = ( (~ ni31)  &  wire35675 ) | ( (~ ni30)  &  wire35675 ) | ( n_n434  &  wire35675 ) ;
 assign wire285 = ( wire830  &  (~ n_n434)  &  wire930 ) ;
 assign wire362 = ( (~ ni2)  &  ni3  &  (~ wire281) ) ;
 assign wire367 = ( n_n13895  &  wire948 ) | ( n_n13895  &  wire6940 ) | ( n_n13895  &  wire29139 ) ;
 assign wire410 = ( ni13  &  (~ ni2)  &  ni14  &  (~ ni3) ) ;
 assign wire430 = ( n_n13895  &  (~ wire494)  &  (~ wire35640)  &  (~ wire35641) ) ;
 assign wire445 = ( (~ ni41)  &  ni4  &  ni32 ) ;
 assign wire469 = ( ni4  &  ni5 ) | ( ni4  &  (~ ni6) ) ;
 assign wire470 = ( ni4  &  (~ ni31) ) | ( ni4  &  (~ ni30) ) | ( ni4  &  n_n434 ) ;
 assign wire479 = ( pi23  &  (~ pi24)  &  (~ ni3)  &  (~ ni7) ) ;
 assign wire494 = ( (~ ni3)  &  wire5961 ) | ( (~ ni3)  &  wire5962 ) ;
 assign wire497 = ( (~ wire725)  &  (~ wire6808)  &  (~ wire6809)  &  wire35623 ) ;
 assign wire511 = ( (~ wire6808)  &  (~ wire6809)  &  wire35628 ) ;
 assign wire515 = ( wire29371  &  wire35629 ) | ( (~ ni7)  &  n_n983  &  wire35629 ) ;
 assign wire518 = ( (~ wire539)  &  (~ wire35616)  &  (~ wire35617)  &  wire35619 ) ;
 assign wire520 = ( wire1289  &  (~ wire539)  &  (~ wire35616)  &  (~ wire35617) ) ;
 assign wire521 = ( ni2  &  ni29 ) | ( ni3  &  ni29 ) ;
 assign wire538 = ( wire35365  &  wire35615 ) | ( wire35366  &  wire35615 ) | ( wire35425  &  wire35615 ) ;
 assign wire539 = ( ni9  &  (~ ni8)  &  wire1201 ) | ( ni9  &  (~ ni8)  &  wire35469 ) ;
 assign wire541 = ( (~ wire793)  &  wire35365 ) | ( (~ wire793)  &  wire35366 ) | ( (~ wire793)  &  wire35425 ) ;
 assign wire542 = ( wire1075  &  wire35471 ) | ( wire6705  &  wire35471 ) | ( wire6706  &  wire35471 ) ;
 assign wire544 = ( wire1473  &  wire35475 ) | ( wire35142  &  wire35475 ) | ( wire35143  &  wire35475 ) ;
 assign wire548 = ( wire565  &  wire35487 ) | ( wire566  &  wire35487 ) | ( wire35485  &  wire35487 ) ;
 assign wire550 = ( n_n1593  &  wire35489 ) | ( wire1482  &  wire35489 ) ;
 assign wire551 = ( wire309  &  wire259  &  wire35490 ) ;
 assign wire552 = ( wire1465  &  wire35491 ) | ( wire1467  &  wire35491 ) | ( wire35131  &  wire35491 ) ;
 assign wire558 = ( wire226  &  wire724 ) | ( wire226  &  wire741 ) | ( wire226  &  wire35522 ) ;
 assign wire559 = ( (~ pi15)  &  n_n2484 ) ;
 assign wire561 = ( wire1075  &  wire309 ) | ( wire309  &  wire6540 ) | ( wire309  &  wire6541 ) ;
 assign wire562 = ( wire211  &  wire405 ) | ( (~ pi22)  &  wire211  &  n_n1395 ) ;
 assign wire563 = ( wire189  &  wire1384 ) | ( wire189  &  wire35037 ) ;
 assign wire565 = ( (~ pi25)  &  wire2024 ) | ( (~ pi25)  &  wire2025 ) | ( (~ pi25)  &  wire35006 ) ;
 assign wire566 = ( pi25  &  wire35373 ) | ( pi25  &  wire35374 ) ;
 assign wire568 = ( wire1097  &  wire35492 ) | ( wire6682  &  wire35492 ) | ( wire6683  &  wire35492 ) ;
 assign wire570 = ( wire1542  &  wire35494 ) | ( wire35159  &  wire35494 ) | ( wire35160  &  wire35494 ) ;
 assign wire603 = ( wire1344  &  wire35393 ) | ( wire1344  &  wire35394 ) ;
 assign wire609 = ( wire1027  &  wire35396 ) | ( wire1027  &  wire35397 ) ;
 assign wire624 = ( wire487  &  wire6453 ) | ( wire487  &  wire6454 ) | ( wire487  &  wire29476 ) ;
 assign wire629 = ( wire228  &  wire308 ) | ( (~ pi21)  &  wire228  &  n_n1756 ) ;
 assign wire651 = ( wire1097  &  wire35511 ) | ( wire6616  &  wire35511 ) | ( wire6617  &  wire35511 ) ;
 assign wire709 = ( wire405  &  wire35512 ) | ( (~ pi22)  &  n_n1463  &  wire35512 ) ;
 assign wire710 = ( wire191  &  wire189  &  wire1986 ) | ( wire191  &  wire189  &  wire35023 ) ;
 assign wire724 = ( wire1344  &  wire35377 ) | ( wire1344  &  wire35378 ) ;
 assign wire741 = ( (~ pi25)  &  wire1207 ) | ( (~ pi25)  &  wire1209 ) ;
 assign wire823 = ( wire6613  &  wire35525 ) | ( wire6614  &  wire35525 ) | ( wire29575  &  wire35525 ) ;
 assign wire825 = ( wire1974  &  wire35527 ) | ( wire1982  &  wire35527 ) | ( wire1983  &  wire35527 ) ;
 assign wire879 = ( wire189  &  wire1663  &  wire35528 ) | ( wire189  &  wire35199  &  wire35528 ) ;
 assign wire888 = ( wire1660  &  wire35531 ) | ( wire35004  &  wire35531 ) | ( wire35005  &  wire35531 ) ;
 assign wire894 = ( wire35211  &  wire35532 ) | ( wire35212  &  wire35532 ) ;
 assign wire925 = ( wire35233  &  wire35533 ) | ( wire35234  &  wire35533 ) ;
 assign wire931 = ( (~ pi25)  &  pi16  &  wire786 ) ;
 assign wire932 = ( wire309  &  wire259  &  wire35535 ) ;
 assign wire938 = ( wire6537  &  wire35536 ) | ( wire6538  &  wire35536 ) | ( wire29592  &  wire35536 ) ;
 assign wire939 = ( wire405  &  wire35537 ) | ( (~ pi22)  &  n_n1859  &  wire35537 ) ;
 assign wire944 = ( wire189  &  wire593  &  wire1574 ) | ( wire189  &  wire593  &  wire35247 ) ;
 assign wire945 = ( wire1642  &  wire35539 ) | ( wire1643  &  wire35539 ) | ( wire35223  &  wire35539 ) ;
 assign wire955 = ( wire1569  &  wire35540 ) | ( wire35004  &  wire35540 ) | ( wire35005  &  wire35540 ) ;
 assign wire956 = ( n_n12696  &  wire35541 ) | ( wire29518  &  wire35541 ) ;
 assign wire961 = ( wire35225  &  wire35542 ) | ( wire35226  &  wire35542 ) ;
 assign wire967 = ( (~ ni29)  &  wire152  &  wire154  &  wire259 ) ;
 assign wire969 = ( wire183  &  wire1608 ) | ( wire183  &  wire35186 ) | ( wire183  &  wire35187 ) ;
 assign wire982 = ( wire309  &  wire593  &  wire259 ) ;
 assign wire1001 = ( wire6701  &  wire35562 ) | ( wire6703  &  wire35562 ) | ( wire29652  &  wire35562 ) ;
 assign wire1004 = ( wire405  &  wire35563 ) | ( (~ pi22)  &  n_n2180  &  wire35563 ) ;
 assign wire1040 = ( wire1783  &  wire35565 ) | ( wire1784  &  wire35565 ) | ( wire35295  &  wire35565 ) ;
 assign wire1042 = ( wire308  &  wire35566 ) | ( (~ pi21)  &  n_n2179  &  wire35566 ) ;
 assign wire1054 = ( wire35294  &  wire35567 ) | ( wire213  &  n_n2226  &  wire35567 ) ;
 assign wire1136 = ( (~ ni29)  &  wire158  &  wire152  &  wire259 ) ;
 assign wire1137 = ( wire194  &  wire1756 ) | ( wire194  &  wire35276 ) | ( wire194  &  wire35277 ) ;
 assign wire1141 = ( wire35329  &  wire35568 ) | ( wire863  &  wire35328  &  wire35568 ) ;
 assign wire1143 = ( wire6678  &  wire35569 ) | ( wire6680  &  wire35569 ) | ( wire29635  &  wire35569 ) ;
 assign wire1145 = ( wire1886  &  wire35571 ) | ( wire35298  &  wire35571 ) | ( wire35299  &  wire35571 ) ;
 assign wire1148 = ( wire35315  &  wire35572 ) | ( wire35316  &  wire35572 ) ;
 assign wire1154 = ( wire308  &  wire35574 ) | ( (~ pi21)  &  n_n2280  &  wire35574 ) ;
 assign wire1155 = ( wire1873  &  wire35575 ) | ( wire1874  &  wire35575 ) | ( wire35336  &  wire35575 ) ;
 assign wire1156 = ( wire1027  &  wire1275 ) | ( wire1027  &  wire1861 ) | ( wire1027  &  wire35338 ) ;
 assign wire1157 = ( wire817  &  wire35262 ) | ( (~ pi22)  &  wire817  &  wire860 ) ;
 assign wire1159 = ( (~ pi25)  &  wire1258 ) | ( (~ pi25)  &  wire260  &  n_n1351 ) ;
 assign wire1160 = ( (~ pi17)  &  pi19  &  wire309  &  wire259 ) ;
 assign wire1164 = ( wire171  &  wire1698 ) | ( wire171  &  wire1700 ) | ( wire171  &  wire35268 ) ;
 assign wire1166 = ( wire405  &  wire34994 ) | ( (~ pi22)  &  n_n1463  &  wire34994 ) ;
 assign wire1167 = ( wire2024  &  wire35009 ) | ( wire2025  &  wire35009 ) | ( wire35006  &  wire35009 ) ;
 assign wire1168 = ( wire1984  &  wire35014 ) | ( wire35004  &  wire35014 ) | ( wire35005  &  wire35014 ) ;
 assign wire1169 = ( wire1394  &  wire35020 ) | ( wire1395  &  wire35020 ) | ( wire35017  &  wire35020 ) ;
 assign wire1170 = ( wire1986  &  wire35025 ) | ( wire35023  &  wire35025 ) ;
 assign wire1172 = ( pi16  &  pi15  &  wire289  &  wire995 ) ;
 assign wire1174 = ( wire289  &  wire226  &  wire1207 ) | ( wire289  &  wire226  &  wire1209 ) ;
 assign wire1175 = ( wire35088  &  wire35089 ) | ( nv952  &  wire35076  &  wire35089 ) ;
 assign wire1176 = ( wire289  &  wire395  &  wire309 ) ;
 assign wire1191 = ( pi15  &  wire289  &  wire35178 ) | ( pi15  &  wire289  &  wire35179 ) ;
 assign wire1201 = ( (~ wire289)  &  wire35365 ) | ( (~ wire289)  &  wire35366 ) | ( (~ wire289)  &  wire35425 ) ;
 assign wire1202 = ( wire289  &  wire1221 ) | ( wire289  &  wire1225 ) | ( wire289  &  wire35456 ) ;
 assign wire1207 = ( (~ pi17)  &  pi19  &  wire2061 ) | ( (~ pi17)  &  pi19  &  wire35048 ) ;
 assign wire1209 = ( (~ pi17)  &  (~ pi19)  &  wire1416 ) | ( (~ pi17)  &  (~ pi19)  &  wire35065 ) ;
 assign wire1214 = ( wire1974  &  wire35427 ) | ( wire1982  &  wire35427 ) | ( wire1983  &  wire35427 ) ;
 assign wire1215 = ( wire1642  &  wire35428 ) | ( wire1643  &  wire35428 ) | ( wire35223  &  wire35428 ) ;
 assign wire1216 = ( wire1660  &  wire35429 ) | ( wire35004  &  wire35429 ) | ( wire35005  &  wire35429 ) ;
 assign wire1218 = ( wire1663  &  wire35431 ) | ( wire35199  &  wire35431 ) ;
 assign wire1221 = ( pi16  &  (~ pi15)  &  wire786 ) ;
 assign wire1223 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire309 ) ;
 assign wire1225 = ( (~ pi15)  &  wire1237 ) | ( (~ pi15)  &  wire35445 ) | ( (~ pi15)  &  wire35446 ) ;
 assign wire1228 = ( (~ pi17)  &  (~ pi19)  &  wire1924 ) | ( (~ pi17)  &  (~ pi19)  &  wire35232 ) ;
 assign wire1232 = ( wire35294  &  wire35433 ) | ( wire213  &  n_n2226  &  wire35433 ) ;
 assign wire1233 = ( wire308  &  wire35434 ) | ( (~ pi21)  &  n_n2280  &  wire35434 ) ;
 assign wire1235 = ( wire344  &  wire35329 ) | ( wire344  &  wire863  &  wire35328 ) ;
 assign wire1236 = ( (~ pi16)  &  wire1718 ) | ( (~ pi16)  &  wire1719 ) ;
 assign wire1237 = ( (~ pi16)  &  wire1726 ) | ( (~ pi16)  &  n_n2176  &  wire329 ) ;
 assign wire1238 = ( (~ pi16)  &  wire1258 ) | ( (~ pi16)  &  wire260  &  n_n1351 ) ;
 assign wire1240 = ( wire484  &  wire1886 ) | ( wire484  &  wire35298 ) | ( wire484  &  wire35299 ) ;
 assign wire1251 = ( wire325  &  wire1873 ) | ( wire325  &  wire1874 ) | ( wire325  &  wire35336 ) ;
 assign wire1254 = ( (~ pi17)  &  (~ pi16)  &  wire309 ) ;
 assign wire1258 = ( (~ ni29)  &  wire153 ) ;
 assign wire1270 = ( (~ pi16)  &  wire1463 ) | ( (~ pi16)  &  wire458  &  n_n1243 ) ;
 assign wire1273 = ( wire484  &  wire1542 ) | ( wire484  &  wire35159 ) | ( wire484  &  wire35160 ) ;
 assign wire1353 = ( wire344  &  wire1492 ) | ( wire344  &  wire1493 ) | ( wire344  &  wire35168 ) ;
 assign wire1357 = ( wire1075  &  wire35367 ) | ( wire6540  &  wire35367 ) | ( wire6541  &  wire35367 ) ;
 assign wire1358 = ( nv952  &  wire35368 ) | ( wire157  &  wire35368 ) ;
 assign wire1360 = ( wire1097  &  wire35370 ) | ( wire6616  &  wire35370 ) | ( wire6617  &  wire35370 ) ;
 assign wire1361 = ( wire405  &  wire35371 ) | ( (~ pi22)  &  n_n1463  &  wire35371 ) ;
 assign wire1362 = ( wire1984  &  wire35372 ) | ( wire35004  &  wire35372 ) | ( wire35005  &  wire35372 ) ;
 assign wire1363 = ( wire35373  &  wire35375 ) | ( wire35374  &  wire35375 ) ;
 assign wire1364 = ( wire395  &  wire182  &  wire1986 ) | ( wire395  &  wire182  &  wire35023 ) ;
 assign wire1365 = ( wire35377  &  wire35379 ) | ( wire35378  &  wire35379 ) ;
 assign wire1366 = ( wire35380  &  wire35382 ) | ( wire35381  &  wire35382 ) ;
 assign wire1367 = ( (~ ni29)  &  wire395  &  wire157  &  wire182 ) ;
 assign wire1371 = ( pi16  &  pi15  &  wire1398 ) | ( pi16  &  pi15  &  wire35088 ) ;
 assign wire1374 = ( pi17  &  pi19  &  wire1376 ) | ( pi17  &  pi19  &  wire35028 ) ;
 assign wire1376 = ( pi21  &  (~ pi22)  &  wire1772 ) | ( pi21  &  (~ pi22)  &  wire1773 ) ;
 assign wire1380 = ( (~ pi21)  &  wire35031 ) | ( (~ pi21)  &  n_n1410  &  wire35030 ) ;
 assign wire1382 = ( wire405  &  wire695 ) | ( (~ pi22)  &  n_n1395  &  wire695 ) ;
 assign wire1384 = ( wire316  &  wire1075 ) | ( wire316  &  wire6540 ) | ( wire316  &  wire6541 ) ;
 assign wire1385 = ( ni40  &  wire388  &  wire293 ) | ( (~ ni40)  &  nv772  &  wire293 ) ;
 assign wire1391 = ( (~ ni29)  &  nv858 ) ;
 assign wire1394 = ( (~ ni31)  &  (~ ni30)  &  ni29  &  nv858 ) ;
 assign wire1395 = ( wire245  &  wire1773 ) | ( wire245  &  nv9050  &  wire35016 ) ;
 assign wire1397 = ( wire1406  &  wire35075 ) | ( wire1407  &  wire35075 ) | ( wire1408  &  wire35075 ) ;
 assign wire1398 = ( pi20  &  nv952  &  wire316  &  wire153 ) ;
 assign wire1400 = ( wire1406  &  wire35078 ) | ( wire1407  &  wire35078 ) | ( wire1408  &  wire35078 ) ;
 assign wire1403 = ( pi20  &  wire266  &  wire348  &  wire153 ) ;
 assign wire1404 = ( wire817  &  wire1982 ) | ( (~ pi22)  &  (~ ni29)  &  wire817 ) ;
 assign wire1406 = ( ni36  &  ni32  &  (~ nv354)  &  n_n1566 ) ;
 assign wire1407 = ( wire390  &  wire1634 ) | ( wire390  &  wire1636 ) | ( wire390  &  wire35072 ) ;
 assign wire1408 = ( (~ nv539)  &  wire35072 ) | ( (~ nv539)  &  nv9297  &  wire35070 ) ;
 assign wire1416 = ( wire213  &  wire35063 ) | ( wire316  &  wire213  &  nv942 ) ;
 assign wire1417 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n1558 ) ;
 assign wire1424 = ( ni36  &  ni32  &  (~ nv354)  &  n_n1566 ) ;
 assign wire1426 = ( nv401  &  wire1936 ) | ( nv401  &  wire1938 ) | ( nv401  &  wire35056 ) ;
 assign wire1431 = ( wire1075  &  wire35383 ) | ( wire6705  &  wire35383 ) | ( wire6706  &  wire35383 ) ;
 assign wire1432 = ( wire943  &  wire35384 ) ;
 assign wire1433 = ( (~ pi16)  &  wire272  &  n_n1593 ) | ( (~ pi16)  &  wire272  &  wire1482 ) ;
 assign wire1434 = ( wire1097  &  wire35386 ) | ( wire6682  &  wire35386 ) | ( wire6683  &  wire35386 ) ;
 assign wire1438 = ( wire1542  &  wire35392 ) | ( wire35159  &  wire35392 ) | ( wire35160  &  wire35392 ) ;
 assign wire1439 = ( wire35393  &  wire35395 ) | ( wire35394  &  wire35395 ) ;
 assign wire1440 = ( (~ ni29)  &  wire302  &  wire157  &  wire182 ) ;
 assign wire1442 = ( (~ pi16)  &  wire1463 ) | ( (~ pi16)  &  wire458  &  n_n1243 ) ;
 assign wire1444 = ( wire344  &  wire35396 ) | ( wire344  &  wire35397 ) ;
 assign wire1447 = ( wire308  &  wire697 ) | ( (~ pi21)  &  n_n1756  &  wire697 ) ;
 assign wire1448 = ( wire294  &  wire1454 ) | ( wire294  &  wire35097 ) ;
 assign wire1454 = ( wire316  &  wire6453 ) | ( wire316  &  wire6454 ) | ( wire316  &  wire29476 ) ;
 assign wire1458 = ( ni41  &  wire35093 ) | ( (~ ni41)  &  ni44  &  wire35093 ) | ( (~ ni41)  &  wire934  &  wire35093 ) ;
 assign wire1463 = ( wire299  &  wire1465 ) | ( wire299  &  wire1467 ) | ( wire299  &  wire35131 ) ;
 assign wire1465 = ( wire1770  &  wire35130 ) | ( wire1772  &  wire35130 ) | ( wire1773  &  wire35130 ) ;
 assign wire1466 = ( pi21  &  wire1982 ) | ( pi21  &  (~ pi22)  &  (~ ni29) ) ;
 assign wire1467 = ( (~ pi21)  &  nv9492 ) | ( (~ pi21)  &  ni41  &  ni38 ) ;
 assign wire1471 = ( n_n1241  &  wire695 ) ;
 assign wire1473 = ( wire316  &  wire1075 ) | ( wire316  &  wire6705 ) | ( wire316  &  wire6706 ) ;
 assign wire1474 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  wire441  &  wire293 ) ;
 assign wire1479 = ( nv9066  &  wire701 ) ;
 assign wire1482 = ( (~ ni29)  &  wire320 ) | ( (~ ni29)  &  wire6694 ) ;
 assign wire1484 = ( nv9492  &  wire35125 ) | ( ni41  &  ni38  &  wire35125 ) ;
 assign wire1485 = ( wire320  &  wire316 ) | ( wire316  &  wire6694 ) ;
 assign wire1486 = ( wire245  &  wire1770 ) | ( wire245  &  wire1772 ) | ( wire245  &  wire1773 ) ;
 assign wire1492 = ( wire506  &  wire863 ) | ( wire506  &  wire1501 ) | ( wire506  &  wire1502 ) ;
 assign wire1493 = ( wire213  &  wire1498 ) | ( wire213  &  wire35167 ) ;
 assign wire1494 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n1786 ) ;
 assign wire1498 = ( wire245  &  wire863 ) | ( wire245  &  wire1501 ) | ( wire245  &  wire1502 ) ;
 assign wire1501 = ( ni41  &  wire35163 ) | ( (~ ni41)  &  (~ ni44)  &  wire35163 ) | ( (~ ni41)  &  wire934  &  wire35163 ) ;
 assign wire1502 = ( (~ ni37)  &  ni36  &  ni32  &  n_n1566 ) ;
 assign wire1516 = ( wire1097  &  wire316 ) | ( wire316  &  wire6666 ) | ( wire316  &  wire6667 ) ;
 assign wire1517 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv667  &  wire293 ) | ( ni40  &  nv6576  &  wire293 ) ;
 assign wire1518 = ( wire245  &  wire1082 ) | ( wire245  &  wire1853 ) | ( wire245  &  wire35149 ) ;
 assign wire1519 = ( wire245  &  wire1230 ) | ( wire245  &  wire1840 ) | ( wire245  &  wire35153 ) ;
 assign wire1535 = ( wire316  &  wire1075 ) | ( wire316  &  wire6745 ) | ( wire316  &  wire6746 ) ;
 assign wire1536 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv6576  &  wire293 ) ;
 assign wire1537 = ( wire245  &  wire1023 ) | ( wire245  &  wire1803 ) | ( wire245  &  wire35109 ) ;
 assign wire1538 = ( wire245  &  wire1231 ) | ( wire245  &  wire1813 ) | ( wire245  &  wire35113 ) ;
 assign wire1542 = ( wire1097  &  wire316 ) | ( wire316  &  wire6682 ) | ( wire316  &  wire6683 ) ;
 assign wire1543 = ( (~ ni40)  &  nv667  &  wire293 ) | ( ni40  &  wire441  &  wire293 ) ;
 assign wire1547 = ( wire6537  &  wire35181 ) | ( wire6538  &  wire35181 ) | ( wire29592  &  wire35181 ) ;
 assign wire1548 = ( wire157  &  wire35182 ) | ( n_n12696  &  wire35182 ) | ( wire29518  &  wire35182 ) ;
 assign wire1549 = ( wire1608  &  wire35188 ) | ( wire35186  &  wire35188 ) | ( wire35187  &  wire35188 ) ;
 assign wire1550 = ( wire6613  &  wire35189 ) | ( wire6614  &  wire35189 ) | ( wire29575  &  wire35189 ) ;
 assign wire1551 = ( wire1974  &  wire35192 ) | ( wire1982  &  wire35192 ) | ( wire1983  &  wire35192 ) ;
 assign wire1552 = ( wire1660  &  wire35196 ) | ( wire35004  &  wire35196 ) | ( wire35005  &  wire35196 ) ;
 assign wire1553 = ( wire182  &  wire507  &  wire1663 ) | ( wire182  &  wire507  &  wire35199 ) ;
 assign wire1554 = ( wire35211  &  wire35213 ) | ( wire35212  &  wire35213 ) ;
 assign wire1555 = ( wire35225  &  wire35227 ) | ( wire35226  &  wire35227 ) ;
 assign wire1556 = ( wire35233  &  wire35235 ) | ( wire35234  &  wire35235 ) ;
 assign wire1557 = ( (~ ni29)  &  wire157  &  wire182  &  wire507 ) ;
 assign wire1563 = ( pi17  &  pi19  &  wire626 ) ;
 assign wire1566 = ( pi21  &  wire1982 ) | ( pi21  &  (~ pi22)  &  (~ ni29) ) ;
 assign wire1567 = ( (~ pi21)  &  wire35184 ) | ( (~ pi21)  &  nv9492  &  wire35183 ) ;
 assign wire1569 = ( (~ pi21)  &  wire1578 ) | ( (~ pi21)  &  wire1580 ) | ( (~ pi21)  &  wire35240 ) ;
 assign wire1571 = ( wire405  &  wire695 ) | ( (~ pi22)  &  n_n1859  &  wire695 ) ;
 assign wire1574 = ( wire316  &  wire6537 ) | ( wire316  &  wire6538 ) | ( wire316  &  wire29592 ) ;
 assign wire1575 = ( ni40  &  wire388  &  wire293 ) | ( (~ ni40)  &  nv772  &  wire293 ) ;
 assign wire1578 = ( (~ ni35)  &  (~ ni32)  &  n_n1410 ) | ( (~ ni35)  &  n_n1410  &  wire35031 ) ;
 assign wire1579 = ( (~ ni40)  &  wire907  &  wire341 ) | ( ni40  &  nv9031  &  wire341 ) | ( (~ ni40)  &  nv9031  &  wire341 ) ;
 assign wire1580 = ( (~ ni36)  &  wire35031 ) | ( (~ ni36)  &  n_n1410  &  wire35030 ) ;
 assign wire1585 = ( (~ ni40)  &  (~ wire231)  &  wire907 ) | ( ni40  &  (~ wire231)  &  nv9031 ) | ( (~ ni40)  &  (~ wire231)  &  nv9031 ) ;
 assign wire1602 = ( (~ ni36)  &  wire1607 ) | ( (~ ni36)  &  wire254  &  nv9050 ) ;
 assign wire1604 = ( (~ ni40)  &  wire907 ) | ( (~ ni40)  &  wire2005 ) | ( (~ ni40)  &  wire4913 ) ;
 assign wire1606 = ( ni40  &  ni38  &  nv9050 ) ;
 assign wire1607 = ( wire253  &  wire907 ) | ( wire253  &  wire2005 ) | ( wire253  &  wire4913 ) ;
 assign wire1608 = ( (~ ni29)  &  wire29562 ) | ( (~ ni36)  &  (~ ni29)  &  nv858 ) ;
 assign wire1610 = ( wire316  &  wire29562 ) | ( (~ ni36)  &  wire316  &  nv858 ) ;
 assign wire1622 = ( wire1634  &  wire35248 ) | ( wire1636  &  wire35248 ) | ( wire35072  &  wire35248 ) ;
 assign wire1623 = ( n_n12696  &  wire35249 ) | ( wire29518  &  wire35249 ) ;
 assign wire1625 = ( wire1000  &  wire35251 ) | ( wire1631  &  wire35251 ) ;
 assign wire1626 = ( wire1634  &  wire35252 ) | ( wire1636  &  wire35252 ) | ( wire35072  &  wire35252 ) ;
 assign wire1627 = ( wire1000  &  wire35253 ) | ( wire1631  &  wire35253 ) ;
 assign wire1628 = ( pi20  &  wire153  &  wire1248 ) ;
 assign wire1629 = ( wire817  &  wire1982 ) | ( (~ pi22)  &  (~ ni29)  &  wire817 ) ;
 assign wire1631 = ( nv9031  &  wire898 ) | ( (~ ni41)  &  ni44  &  wire898 ) ;
 assign wire1634 = ( wire907  &  wire35070 ) | ( wire2005  &  wire35070 ) | ( wire4913  &  wire35070 ) ;
 assign wire1636 = ( nv539  &  wire907 ) | ( nv539  &  wire2005 ) | ( nv539  &  wire4913 ) ;
 assign wire1642 = ( wire213  &  wire1648 ) | ( wire213  &  wire1651 ) | ( wire213  &  wire35221 ) ;
 assign wire1643 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n1907 ) ;
 assign wire1647 = ( ni30  &  ni29  &  wire1142 ) | ( ni30  &  ni29  &  wire1794 ) ;
 assign wire1648 = ( wire316  &  wire6557 ) | ( wire316  &  wire6558 ) | ( wire316  &  wire29587 ) ;
 assign wire1649 = ( (~ ni40)  &  nv758  &  wire293 ) | ( ni40  &  wire388  &  wire293 ) ;
 assign wire1651 = ( ni31  &  (~ ni30)  &  ni29  &  n_n1908 ) ;
 assign wire1660 = ( (~ pi21)  &  wire1667 ) | ( (~ pi21)  &  wire1669 ) | ( (~ pi21)  &  wire35194 ) ;
 assign wire1662 = ( ni30  &  ni29  &  wire1146 ) | ( ni30  &  ni29  &  wire1890 ) ;
 assign wire1663 = ( wire316  &  wire6613 ) | ( wire316  &  wire6614 ) | ( wire316  &  wire29575 ) ;
 assign wire1664 = ( (~ ni40)  &  wire388  &  wire293 ) | ( ni40  &  nv772  &  wire293 ) ;
 assign wire1665 = ( wire245  &  wire1667 ) | ( wire245  &  wire1669 ) | ( wire245  &  wire35194 ) ;
 assign wire1666 = ( wire245  &  wire35191 ) | ( (~ nv539)  &  wire245  &  n_n1463 ) ;
 assign wire1667 = ( ni35  &  (~ ni32)  &  n_n1478 ) | ( ni35  &  n_n1478  &  wire35012 ) ;
 assign wire1668 = ( ni40  &  wire907  &  wire341 ) | ( ni40  &  nv9031  &  wire341 ) | ( (~ ni40)  &  nv9031  &  wire341 ) ;
 assign wire1669 = ( (~ ni36)  &  wire35012 ) | ( (~ ni36)  &  n_n1478  &  wire35011 ) ;
 assign wire1671 = ( wire6701  &  wire35271 ) | ( wire6703  &  wire35271 ) | ( wire29652  &  wire35271 ) ;
 assign wire1672 = ( wire1756  &  wire35278 ) | ( wire35276  &  wire35278 ) | ( wire35277  &  wire35278 ) ;
 assign wire1673 = ( wire785  &  wire35279 ) ;
 assign wire1674 = ( wire6678  &  wire35280 ) | ( wire6680  &  wire35280 ) | ( wire29635  &  wire35280 ) ;
 assign wire1676 = ( wire308  &  wire35287 ) | ( (~ pi21)  &  n_n2280  &  wire35287 ) ;
 assign wire1677 = ( wire1783  &  wire35297 ) | ( wire1784  &  wire35297 ) | ( wire35295  &  wire35297 ) ;
 assign wire1678 = ( wire1886  &  wire35301 ) | ( wire35298  &  wire35301 ) | ( wire35299  &  wire35301 ) ;
 assign wire1680 = ( (~ ni29)  &  wire302  &  wire157  &  wire182 ) ;
 assign wire1682 = ( (~ pi16)  &  wire1718 ) | ( (~ pi16)  &  wire1719 ) ;
 assign wire1683 = ( (~ pi16)  &  wire1726 ) | ( (~ pi16)  &  n_n2176  &  wire329 ) ;
 assign wire1684 = ( wire344  &  wire1275 ) | ( wire344  &  wire1861 ) | ( wire344  &  wire35338 ) ;
 assign wire1686 = ( wire843  &  wire35262 ) | ( (~ pi22)  &  wire860  &  wire843 ) ;
 assign wire1688 = ( wire294  &  wire1698 ) | ( wire294  &  wire1700 ) | ( wire294  &  wire35268 ) ;
 assign wire1689 = ( ni41  &  wire35261 ) | ( (~ ni41)  &  ni44  &  wire35261 ) | ( (~ ni41)  &  wire934  &  wire35261 ) ;
 assign wire1697 = ( wire1708  &  wire35264 ) | ( (~ ni38)  &  ni37  &  wire35264 ) ;
 assign wire1698 = ( wire1302  &  wire820 ) | ( wire820  &  wire1705 ) | ( wire820  &  wire1706 ) ;
 assign wire1699 = ( (~ ni32)  &  ni30  &  ni29  &  wire441 ) ;
 assign wire1700 = ( wire316  &  wire6722 ) | ( wire316  &  wire29474 ) | ( wire316  &  wire29475 ) ;
 assign wire1701 = ( wire245  &  wire1000 ) | ( wire245  &  wire1710 ) ;
 assign wire1705 = ( ni41  &  wire269 ) | ( (~ ni41)  &  ni44  &  wire269 ) | ( (~ ni41)  &  wire269  &  wire934 ) ;
 assign wire1706 = ( (~ ni36)  &  wire1708 ) | ( (~ ni38)  &  ni37  &  (~ ni36) ) ;
 assign wire1708 = ( ni41  &  ni37 ) | ( (~ ni41)  &  ni44  &  ni37 ) | ( (~ ni41)  &  ni37  &  wire934 ) ;
 assign wire1710 = ( ni41  &  wire898 ) | ( nv9031  &  wire898 ) | ( (~ ni41)  &  ni44  &  wire898 ) ;
 assign wire1718 = ( pi17  &  pi19  &  wire1720 ) | ( pi17  &  pi19  &  wire35320 ) ;
 assign wire1719 = ( wire458  &  wire308 ) | ( (~ pi21)  &  wire458  &  n_n2179 ) ;
 assign wire1720 = ( pi21  &  (~ pi22)  &  wire1765 ) | ( pi21  &  (~ pi22)  &  wire35272 ) ;
 assign wire1721 = ( pi21  &  wire1982 ) | ( pi21  &  (~ pi22)  &  (~ ni29) ) ;
 assign wire1726 = ( wire405  &  wire695 ) | ( (~ pi22)  &  n_n2180  &  wire695 ) ;
 assign wire1732 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  wire441  &  wire293 ) ;
 assign wire1735 = ( ni37  &  ni36  &  ni32  &  (~ nv401) ) ;
 assign wire1740 = ( wire357  &  wire461 ) | ( wire382  &  n_n1966  &  wire461 ) ;
 assign wire1742 = ( (~ ni40)  &  wire4913 ) | ( (~ ni41)  &  (~ ni40)  &  ni44 ) ;
 assign wire1754 = ( (~ ni35)  &  ni32  &  wire3491 ) | ( (~ ni35)  &  ni32  &  wire33310 ) ;
 assign wire1756 = ( (~ ni29)  &  wire436 ) | ( (~ ni29)  &  wire6691 ) | ( (~ ni29)  &  wire6692 ) ;
 assign wire1763 = ( ni42  &  wire293 ) | ( nv669  &  wire293 ) | ( (~ ni42)  &  ni41  &  wire293 ) ;
 assign wire1765 = ( (~ nv539)  &  wire1770 ) | ( (~ nv539)  &  wire1772 ) | ( (~ nv539)  &  wire1773 ) ;
 assign wire1770 = ( ni41  &  ni38  &  ni32 ) ;
 assign wire1772 = ( ni38  &  ni32  &  nv9050 ) ;
 assign wire1773 = ( (~ ni38)  &  ni37  &  ni32 ) | ( (~ ni38)  &  (~ ni37)  &  ni32  &  wire770 ) ;
 assign wire1777 = ( ni41  &  ni38 ) ;
 assign wire1783 = ( nv703  &  wire35294 ) | ( nv703  &  wire213  &  n_n2226 ) ;
 assign wire1784 = ( n_n1329  &  wire35294 ) | ( wire213  &  n_n1329  &  n_n2226 ) ;
 assign wire1787 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n2228 ) ;
 assign wire1791 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv6576  &  wire293 ) ;
 assign wire1794 = ( (~ ni35)  &  ni32  &  wire3462 ) | ( (~ ni35)  &  ni32  &  wire33267 ) ;
 assign wire1798 = ( ni37  &  ni36  &  ni32  &  (~ nv401) ) ;
 assign wire1803 = ( wire357  &  wire461 ) | ( wire382  &  n_n2448  &  wire461 ) ;
 assign wire1805 = ( (~ ni40)  &  wire4971 ) | ( (~ ni41)  &  (~ ni40)  &  (~ ni44) ) ;
 assign wire1813 = ( n_n2466  &  wire35110 ) ;
 assign wire1827 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n2332 ) ;
 assign wire1831 = ( ni30  &  ni29  &  wire1146 ) | ( ni30  &  ni29  &  wire1970 ) ;
 assign wire1832 = ( wire316  &  wire6663 ) | ( wire316  &  wire6664 ) | ( wire316  &  wire29628 ) ;
 assign wire1833 = ( ni40  &  nv667  &  wire293 ) | ( (~ ni40)  &  nv667  &  wire293 ) | ( ni40  &  nv6576  &  wire293 ) ;
 assign wire1835 = ( wire245  &  wire1849 ) | ( wire245  &  wire35308 ) ;
 assign wire1840 = ( n_n2466  &  wire35151 ) ;
 assign wire1845 = ( ni41  &  wire35303 ) | ( wire1101  &  wire35303 ) | ( wire1855  &  wire35303 ) ;
 assign wire1847 = ( (~ ni38)  &  (~ ni36)  &  nv590  &  n_n2448 ) ;
 assign wire1848 = ( (~ nv401)  &  wire806 ) ;
 assign wire1849 = ( (~ ni36)  &  wire35148 ) | ( (~ ni32)  &  wire35148 ) | ( (~ ni36)  &  wire35149 ) | ( (~ ni32)  &  wire35149 ) ;
 assign wire1853 = ( nv590  &  wire357 ) | ( wire382  &  nv590  &  n_n2448 ) ;
 assign wire1855 = ( ni40  &  wire4971 ) | ( (~ ni41)  &  ni40  &  (~ ni44) ) ;
 assign wire1860 = ( wire157  &  wire35330 ) | ( n_n12782  &  wire35330 ) | ( wire29481  &  wire35330 ) ;
 assign wire1861 = ( wire213  &  wire1873 ) | ( wire213  &  wire1874 ) | ( wire213  &  wire35336 ) ;
 assign wire1866 = ( pi21  &  (~ pi20)  &  wire1982 ) | ( pi21  &  (~ pi20)  &  wire1983 ) ;
 assign wire1872 = ( wire1881  &  wire35332 ) | ( (~ ni38)  &  ni37  &  wire35332 ) ;
 assign wire1873 = ( wire1304  &  wire820 ) | ( wire820  &  wire1878 ) | ( wire820  &  wire1879 ) ;
 assign wire1874 = ( wire316  &  n_n12782 ) | ( wire316  &  wire29481 ) ;
 assign wire1875 = ( (~ ni32)  &  ni30  &  ni29  &  nv628 ) ;
 assign wire1876 = ( wire245  &  wire999 ) | ( wire245  &  wire1883 ) ;
 assign wire1878 = ( ni41  &  wire292 ) | ( (~ ni41)  &  (~ ni44)  &  wire292 ) | ( (~ ni41)  &  wire292  &  wire934 ) ;
 assign wire1879 = ( (~ ni36)  &  wire1881 ) | ( (~ ni38)  &  ni37  &  (~ ni36) ) ;
 assign wire1881 = ( ni41  &  ni37 ) | ( (~ ni41)  &  (~ ni44)  &  ni37 ) | ( (~ ni41)  &  ni37  &  wire934 ) ;
 assign wire1883 = ( nv9031  &  wire897 ) | ( ni41  &  (~ nv9031)  &  wire897 ) | ( (~ ni44)  &  (~ nv9031)  &  wire897 ) ;
 assign wire1886 = ( wire316  &  wire6678 ) | ( wire316  &  wire6680 ) | ( wire316  &  wire29635 ) ;
 assign wire1887 = ( (~ ni40)  &  nv667  &  wire293 ) | ( ni40  &  wire441  &  wire293 ) ;
 assign wire1890 = ( ni35  &  ni32  &  wire3491 ) | ( ni35  &  ni32  &  wire33310 ) ;
 assign wire1892 = ( ni41  &  wire35281 ) | ( wire1101  &  wire35281 ) | ( wire1903  &  wire35281 ) ;
 assign wire1893 = ( (~ ni38)  &  (~ ni36)  &  nv590  &  n_n1966 ) ;
 assign wire1894 = ( (~ nv401)  &  wire806 ) ;
 assign wire1895 = ( ni36  &  ni32  &  wire1903 ) | ( ni36  &  ni32  &  wire35099 ) ;
 assign wire1896 = ( (~ ni36)  &  wire35102 ) | ( (~ ni32)  &  wire35102 ) | ( (~ ni36)  &  wire35103 ) | ( (~ ni32)  &  wire35103 ) ;
 assign wire1901 = ( nv590  &  wire357 ) | ( wire382  &  nv590  &  n_n1966 ) ;
 assign wire1903 = ( ni40  &  wire4913 ) | ( (~ ni41)  &  ni40  &  ni44 ) ;
 assign wire1924 = ( wire213  &  wire1927 ) | ( wire213  &  wire35228 ) | ( wire213  &  wire35229 ) ;
 assign wire1927 = ( wire316  &  n_n12706 ) | ( wire316  &  wire29534 ) ;
 assign wire1928 = ( (~ ni32)  &  ni30  &  ni29  &  nv758 ) ;
 assign wire1936 = ( wire1076  &  wire35053 ) | ( wire2087  &  wire35053 ) | ( wire4971  &  wire35053 ) ;
 assign wire1938 = ( nv539  &  wire1076 ) | ( nv539  &  wire2087 ) | ( nv539  &  wire4971 ) ;
 assign wire1941 = ( nv9031  &  wire897 ) | ( (~ ni41)  &  (~ ni44)  &  (~ nv9031)  &  wire897 ) ;
 assign wire1951 = ( wire506  &  wire35202 ) | ( (~ nv539)  &  wire506  &  n_n1495 ) ;
 assign wire1952 = ( wire213  &  wire1958 ) | ( wire213  &  wire35208 ) ;
 assign wire1953 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n2009 ) ;
 assign wire1958 = ( wire316  &  wire6577 ) | ( wire316  &  wire6578 ) | ( wire316  &  wire29568 ) ;
 assign wire1959 = ( ni40  &  nv758  &  wire293 ) | ( (~ ni40)  &  wire388  &  wire293 ) ;
 assign wire1970 = ( ni35  &  ni32  &  wire3462 ) | ( ni35  &  ni32  &  wire33267 ) ;
 assign wire1974 = ( (~ pi22)  &  wire35191 ) | ( (~ pi22)  &  (~ nv539)  &  n_n1463 ) ;
 assign wire1982 = ( (~ pi22)  &  (~ ni32) ) | ( (~ pi22)  &  (~ ni31) ) | ( (~ pi22)  &  ni30 ) ;
 assign wire1983 = ( (~ pi22)  &  (~ ni29) ) ;
 assign wire1984 = ( (~ pi21)  &  wire35012 ) | ( (~ pi21)  &  n_n1478  &  wire35011 ) ;
 assign wire1986 = ( wire1097  &  wire316 ) | ( wire316  &  wire6616 ) | ( wire316  &  wire6617 ) ;
 assign wire1987 = ( (~ ni40)  &  wire388  &  wire293 ) | ( ni40  &  nv772  &  wire293 ) ;
 assign wire1992 = ( (~ ni35)  &  nv9066  &  wire266 ) ;
 assign wire1999 = ( (~ ni36)  &  wire2003 ) | ( (~ ni36)  &  wire253  &  nv9050 ) ;
 assign wire2001 = ( ni40  &  wire907 ) | ( ni40  &  wire2005 ) | ( ni40  &  wire4913 ) ;
 assign wire2003 = ( wire254  &  wire907 ) | ( wire254  &  wire2005 ) | ( wire254  &  wire4913 ) ;
 assign wire2004 = ( (~ ni40)  &  ni38  &  nv9050 ) ;
 assign wire2005 = ( ni43  &  ni41 ) | ( ni42  &  ni41 ) | ( (~ ni43)  &  ni41  &  ni45 ) ;
 assign wire2010 = ( ni40  &  (~ wire231)  &  wire907 ) | ( ni40  &  (~ wire231)  &  nv9031 ) | ( (~ ni40)  &  (~ wire231)  &  nv9031 ) ;
 assign wire2024 = ( wire213  &  wire2029 ) | ( wire213  &  wire35003 ) ;
 assign wire2025 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n1426 ) ;
 assign wire2029 = ( wire316  &  wire1075 ) | ( wire316  &  wire6560 ) | ( wire316  &  wire6561 ) ;
 assign wire2030 = ( (~ ni40)  &  nv758  &  wire293 ) | ( ni40  &  wire388  &  wire293 ) ;
 assign wire2035 = ( nv9066  &  wire701 ) ;
 assign wire2040 = ( (~ ni36)  &  wire2045 ) | ( (~ ni36)  &  wire254  &  nv9031 ) ;
 assign wire2044 = ( ni40  &  ni38  &  nv9031 ) ;
 assign wire2045 = ( wire253  &  nv9031 ) | ( (~ ni41)  &  (~ ni44)  &  wire253  &  (~ nv9031) ) ;
 assign wire2050 = ( (~ ni36)  &  wire2055 ) | ( (~ ni36)  &  wire254  &  nv9050 ) ;
 assign wire2052 = ( (~ ni40)  &  wire1076 ) | ( (~ ni40)  &  wire2087 ) | ( (~ ni40)  &  wire4971 ) ;
 assign wire2054 = ( ni40  &  ni38  &  nv9050 ) ;
 assign wire2055 = ( wire253  &  wire1076 ) | ( wire253  &  wire2087 ) | ( wire253  &  wire4971 ) ;
 assign wire2061 = ( wire213  &  wire2066 ) | ( wire213  &  wire35046 ) ;
 assign wire2062 = ( (~ pi20)  &  wire308 ) | ( (~ pi21)  &  (~ pi20)  &  n_n1494 ) ;
 assign wire2065 = ( pi21  &  (~ pi20)  &  (~ ni29) ) ;
 assign wire2066 = ( wire1097  &  wire316 ) | ( wire316  &  wire6580 ) | ( wire316  &  wire6581 ) ;
 assign wire2067 = ( ni40  &  nv758  &  wire293 ) | ( (~ ni40)  &  wire388  &  wire293 ) ;
 assign wire2072 = ( (~ ni35)  &  nv9066  &  wire266 ) ;
 assign wire2081 = ( (~ ni36)  &  wire2085 ) | ( (~ ni36)  &  wire253  &  nv9050 ) ;
 assign wire2083 = ( ni40  &  wire1076 ) | ( ni40  &  wire2087 ) | ( ni40  &  wire4971 ) ;
 assign wire2085 = ( wire254  &  wire1076 ) | ( wire254  &  wire2087 ) | ( wire254  &  wire4971 ) ;
 assign wire2086 = ( (~ ni40)  &  ni38  &  nv9050 ) ;
 assign wire2087 = ( ni43  &  ni41 ) | ( ni42  &  ni41 ) | ( (~ ni43)  &  ni41  &  ni45 ) ;
 assign wire2101 = ( (~ ni36)  &  wire2107 ) | ( (~ ni36)  &  wire253  &  nv9031 ) ;
 assign wire2107 = ( wire254  &  nv9031 ) | ( (~ ni41)  &  (~ ni44)  &  wire254  &  (~ nv9031) ) ;
 assign wire2108 = ( (~ ni40)  &  ni38  &  nv9031 ) ;
 assign wire2111 = ( wire1029  &  (~ wire6808)  &  (~ wire6809)  &  wire34974 ) ;
 assign wire2112 = ( wire6808  &  wire34977 ) | ( wire6809  &  wire34977 ) ;
 assign wire2115 = ( (~ ni4)  &  ni3  &  (~ ni30)  &  (~ ni5) ) ;
 assign wire2116 = ( (~ nv10252)  &  (~ wire6811)  &  wire34981 ) | ( (~ wire6811)  &  (~ wire29256)  &  wire34981 ) ;
 assign wire2117 = ( (~ ni5)  &  (~ ni6) ) ;
 assign wire2118 = ( (~ nv10252)  &  (~ wire6811)  &  wire34983 ) | ( (~ wire6811)  &  (~ wire29256)  &  wire34983 ) ;
 assign wire2119 = ( wire33627  &  wire33662 ) | ( wire33628  &  wire33662 ) | ( wire33660  &  wire33662 ) ;
 assign wire2120 = ( wire2308  &  wire33735 ) | ( wire33733  &  wire33735 ) ;
 assign wire2121 = ( nv6450  &  wire33774 ) ;
 assign wire2122 = ( wire33858  &  wire33863 ) | ( wire33859  &  wire33863 ) | ( wire33861  &  wire33863 ) ;
 assign wire2124 = ( wire3177  &  wire33907 ) | ( wire33906  &  wire33907 ) ;
 assign wire2126 = ( ni2  &  ni30 ) | ( ni3  &  ni30 ) ;
 assign wire2128 = ( wire2892  &  wire33918 ) | ( wire33914  &  wire33918 ) ;
 assign wire2129 = ( wire3150  &  wire33922 ) | ( wire3151  &  wire33922 ) ;
 assign wire2130 = ( wire3157  &  wire33926 ) | ( wire3158  &  wire33926 ) ;
 assign wire2133 = ( (~ pi21)  &  wire33933  &  wire33935 ) | ( (~ pi22)  &  wire33933  &  wire33935 ) ;
 assign wire2134 = ( wire3157  &  wire33938 ) | ( wire3158  &  wire33938 ) ;
 assign wire2137 = ( wire3150  &  wire33949 ) | ( wire3151  &  wire33949 ) ;
 assign wire2141 = ( wire34262  &  wire34347 ) | ( wire34263  &  wire34347 ) | ( wire34346  &  wire34347 ) ;
 assign wire2143 = ( wire2593  &  wire34533 ) | ( wire34532  &  wire34533 ) ;
 assign wire2145 = ( wire2902  &  wire34806 ) | ( wire34803  &  wire34806 ) | ( wire34804  &  wire34806 ) ;
 assign wire2148 = ( ni7  &  wire2828 ) | ( ni7  &  wire2830 ) | ( ni7  &  wire34945 ) ;
 assign wire2150 = ( wire2225  &  wire33986 ) | ( wire33956  &  wire33986 ) ;
 assign wire2151 = ( n_n4412  &  wire181  &  wire33987 ) ;
 assign wire2152 = ( (~ n_n5514)  &  wire1006  &  wire33990 ) | ( (~ n_n5514)  &  wire33609  &  wire33990 ) ;
 assign wire2153 = ( (~ pi17)  &  pi16  &  wire358  &  n_n4441 ) ;
 assign wire2154 = ( wire2218  &  wire33992 ) | ( wire179  &  wire276  &  wire33992 ) ;
 assign wire2159 = ( pi16  &  wire2215 ) | ( pi16  &  wire2216 ) | ( pi16  &  wire2217 ) ;
 assign wire2160 = ( wire154  &  wire2220 ) | ( wire178  &  wire154  &  wire276 ) ;
 assign wire2165 = ( wire2225  &  wire33958 ) | ( wire33956  &  wire33958 ) ;
 assign wire2167 = ( (~ n_n5574)  &  wire1006  &  wire33962 ) | ( (~ n_n5574)  &  wire33604  &  wire33962 ) ;
 assign wire2168 = ( (~ pi17)  &  (~ pi16)  &  n_n4509  &  wire358 ) ;
 assign wire2169 = ( wire2218  &  wire33964 ) | ( wire179  &  wire276  &  wire33964 ) ;
 assign wire2173 = ( (~ n_n5580)  &  wire1006  &  wire33968 ) | ( (~ n_n5580)  &  wire33599  &  wire33968 ) ;
 assign wire2174 = ( (~ pi16)  &  wire2215 ) | ( (~ pi16)  &  wire2216 ) | ( (~ pi16)  &  wire2217 ) ;
 assign wire2175 = ( wire158  &  wire2220 ) | ( wire158  &  wire178  &  wire276 ) ;
 assign wire2178 = ( wire3322  &  wire34035 ) | ( n_n4509  &  wire33475  &  wire34035 ) ;
 assign wire2181 = ( wire3251  &  wire34038 ) | ( n_n4481  &  wire33350  &  wire34038 ) ;
 assign wire2182 = ( wire3327  &  wire34039 ) | ( (~ n_n5580)  &  wire33598  &  wire34039 ) ;
 assign wire2184 = ( wire2225  &  wire34041 ) | ( wire33956  &  wire34041 ) ;
 assign wire2185 = ( wire3308  &  wire34042 ) | ( (~ n_n5574)  &  wire33603  &  wire34042 ) ;
 assign wire2187 = ( wire3318  &  wire34044 ) | ( n_n4501  &  wire33595  &  wire34044 ) ;
 assign wire2191 = ( wire158  &  wire2220 ) | ( wire158  &  wire178  &  wire276 ) ;
 assign wire2193 = ( (~ pi25)  &  wire294  &  wire3157 ) | ( (~ pi25)  &  wire294  &  wire3158 ) ;
 assign wire2197 = ( (~ pi21)  &  nv7791  &  wire295 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire295 ) ;
 assign wire2199 = ( wire3341  &  wire34011 ) | ( n_n4433  &  wire33515  &  wire34011 ) ;
 assign wire2200 = ( wire2225  &  wire34013 ) | ( wire33956  &  wire34013 ) ;
 assign wire2201 = ( wire3189  &  wire34015 ) | ( n_n4412  &  wire33395  &  wire34015 ) ;
 assign wire2202 = ( wire3215  &  wire34017 ) | ( (~ n_n5514)  &  wire33608  &  wire34017 ) ;
 assign wire2204 = ( wire2218  &  wire34019 ) | ( wire179  &  wire276  &  wire34019 ) ;
 assign wire2207 = ( pi16  &  wire219  &  wire3205 ) | ( pi16  &  wire219  &  wire3206 ) ;
 assign wire2208 = ( wire345  &  wire154  &  wire3185 ) | ( wire345  &  wire154  &  wire3186 ) ;
 assign wire2209 = ( pi16  &  wire2215 ) | ( pi16  &  wire2216 ) | ( pi16  &  wire2217 ) ;
 assign wire2210 = ( wire154  &  wire2220 ) | ( wire178  &  wire154  &  wire276 ) ;
 assign wire2214 = ( (~ pi21)  &  nv7791  &  wire257 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire257 ) ;
 assign wire2215 = ( n_n3349  &  wire163 ) | ( n_n3347  &  wire163  &  wire204 ) ;
 assign wire2216 = ( (~ pi20)  &  pi25  &  nv7791  &  wire153 ) ;
 assign wire2217 = ( (~ pi25)  &  wire169  &  wire3157 ) | ( (~ pi25)  &  wire169  &  wire3158 ) ;
 assign wire2218 = ( pi19  &  n_n3349 ) | ( pi19  &  n_n3347  &  wire204 ) ;
 assign wire2220 = ( (~ pi19)  &  n_n3349 ) | ( (~ pi19)  &  n_n3347  &  wire204 ) ;
 assign wire2224 = ( ni30  &  wire155  &  wire181 ) | ( (~ wire155)  &  nv7447  &  wire181 ) ;
 assign wire2225 = ( (~ pi25)  &  (~ wire150)  &  wire3157 ) | ( (~ pi25)  &  (~ wire150)  &  wire3158 ) ;
 assign wire2227 = ( wire196  &  wire34266 ) | ( wire192  &  n_n4501  &  wire34266 ) ;
 assign wire2228 = ( wire1016  &  wire2409  &  wire34268 ) | ( wire1016  &  wire34070  &  wire34268 ) ;
 assign wire2229 = ( wire196  &  wire34271 ) | ( wire192  &  n_n4509  &  wire34271 ) ;
 assign wire2230 = ( wire1093  &  wire2576  &  wire34272 ) | ( wire1093  &  wire34063  &  wire34272 ) ;
 assign wire2235 = ( wire2382  &  wire34281 ) | ( wire2387  &  wire34281 ) | ( wire34089  &  wire34281 ) ;
 assign wire2236 = ( wire2389  &  wire34282 ) | ( wire2390  &  wire34282 ) | ( wire2391  &  wire34282 ) ;
 assign wire2237 = ( (~ pi21)  &  nv7791  &  wire34283 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire34283 ) ;
 assign wire2238 = ( wire1339  &  wire33627 ) | ( wire1339  &  wire33628 ) | ( wire1339  &  wire33660 ) ;
 assign wire2239 = ( ni11  &  wire370  &  wire2435 ) | ( ni11  &  wire370  &  wire34297 ) ;
 assign wire2240 = ( ni11  &  wire370  &  wire2486 ) | ( ni11  &  wire370  &  wire34318 ) ;
 assign wire2241 = ( wire1016  &  wire2533 ) | ( wire1016  &  wire34330 ) | ( wire1016  &  wire34331 ) ;
 assign wire2243 = ( wire832  &  wire2576  &  wire34064 ) | ( wire832  &  wire34063  &  wire34064 ) ;
 assign wire2244 = ( wire196  &  wire34067 ) | ( wire192  &  n_n4509  &  wire34067 ) ;
 assign wire2245 = ( wire196  &  wire34069 ) | ( wire192  &  n_n4501  &  wire34069 ) ;
 assign wire2246 = ( wire690  &  wire2409  &  wire34071 ) | ( wire690  &  wire34070  &  wire34071 ) ;
 assign wire2250 = ( wire2382  &  wire34091 ) | ( wire2387  &  wire34091 ) | ( wire34089  &  wire34091 ) ;
 assign wire2251 = ( wire2389  &  wire34092 ) | ( wire2390  &  wire34092 ) | ( wire2391  &  wire34092 ) ;
 assign wire2253 = ( wire1083  &  wire2269 ) | ( wire1083  &  wire34124 ) | ( wire1083  &  wire34125 ) ;
 assign wire2254 = ( wire1083  &  wire2379 ) | ( wire1083  &  wire34147 ) | ( wire1083  &  wire34148 ) ;
 assign wire2255 = ( (~ pi15)  &  wire377  &  wire2277 ) | ( (~ pi15)  &  wire377  &  wire34182 ) ;
 assign wire2256 = ( (~ pi15)  &  wire377  &  wire2289 ) | ( (~ pi15)  &  wire377  &  wire34212 ) ;
 assign wire2257 = ( wire848  &  wire2427 ) | ( wire848  &  wire34220 ) | ( wire848  &  wire34221 ) ;
 assign wire2258 = ( (~ pi15)  &  wire268  &  wire2367 ) | ( (~ pi15)  &  wire268  &  wire34232 ) ;
 assign wire2259 = ( (~ pi15)  &  wire268  &  wire2418 ) | ( (~ pi15)  &  wire268  &  wire34246 ) ;
 assign wire2260 = ( wire618  &  wire33627 ) | ( wire618  &  wire33628 ) | ( wire618  &  wire33660 ) ;
 assign wire2261 = ( (~ ni11)  &  wire2308 ) | ( (~ ni11)  &  wire33733 ) ;
 assign wire2262 = ( wire196  &  wire34095 ) | ( n_n4433  &  wire192  &  wire34095 ) ;
 assign wire2263 = ( wire2571  &  wire34098 ) | ( wire34096  &  wire34098 ) ;
 assign wire2265 = ( wire2554  &  wire34109 ) | ( wire34108  &  wire34109 ) ;
 assign wire2266 = ( wire2560  &  wire34110 ) | ( wire2562  &  wire34110 ) | ( wire2563  &  wire34110 ) ;
 assign wire2267 = ( pi16  &  wire1337 ) ;
 assign wire2268 = ( pi27  &  wire2545 ) | ( pi26  &  wire2545 ) | ( pi27  &  wire34111 ) | ( pi26  &  wire34111 ) ;
 assign wire2269 = ( (~ pi27)  &  (~ pi26)  &  wire653 ) ;
 assign wire2270 = ( (~ pi21)  &  nv7445  &  wire154 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire154 ) ;
 assign wire2274 = ( wire2456  &  wire34165 ) | ( wire34164  &  wire34165 ) ;
 assign wire2275 = ( pi27  &  pi16  &  wire640 ) | ( pi26  &  pi16  &  wire640 ) ;
 assign wire2277 = ( (~ pi27)  &  (~ pi26)  &  wire657 ) ;
 assign wire2278 = ( pi27  &  wire2446 ) | ( pi26  &  wire2446 ) | ( pi27  &  wire34170 ) | ( pi26  &  wire34170 ) ;
 assign wire2279 = ( (~ pi21)  &  nv7445  &  wire154 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire154 ) ;
 assign wire2285 = ( wire34193  &  wire34194 ) | ( nv10153  &  wire527  &  wire34194 ) ;
 assign wire2286 = ( (~ pi16)  &  wire1337 ) ;
 assign wire2288 = ( (~ pi21)  &  wire158  &  nv7445 ) | ( pi21  &  (~ pi22)  &  wire158  &  nv7445 ) ;
 assign wire2289 = ( (~ pi27)  &  (~ pi26)  &  wire672 ) ;
 assign wire2290 = ( pi27  &  wire2498 ) | ( pi26  &  wire2498 ) | ( pi27  &  wire34198 ) | ( pi26  &  wire34198 ) ;
 assign wire2295 = ( pi19  &  ni30  &  (~ wire175)  &  wire33669 ) ;
 assign wire2298 = ( pi15  &  ni30  &  (~ wire175)  &  wire344 ) ;
 assign wire2299 = ( (~ n_n5580)  &  wire1006  &  wire33678 ) | ( (~ n_n5580)  &  wire33599  &  wire33678 ) ;
 assign wire2300 = ( (~ n_n5574)  &  wire1006  &  wire33680 ) | ( (~ n_n5574)  &  wire33604  &  wire33680 ) ;
 assign wire2301 = ( wire33682  &  wire33684 ) | ( n_n4481  &  wire329  &  wire33684 ) ;
 assign wire2302 = ( wire1006  &  (~ n_n5520)  &  wire33685 ) | ( (~ n_n5520)  &  wire33612  &  wire33685 ) ;
 assign wire2303 = ( (~ n_n5514)  &  wire1006  &  wire33686 ) | ( (~ n_n5514)  &  wire33609  &  wire33686 ) ;
 assign wire2304 = ( pi19  &  ni30  &  (~ wire175)  &  wire395 ) ;
 assign wire2305 = ( wire915  &  wire33688 ) ;
 assign wire2306 = ( n_n4404  &  wire33689 ) ;
 assign wire2308 = ( wire613  &  wire33627 ) | ( wire613  &  wire33628 ) | ( wire613  &  wire33660 ) ;
 assign wire2310 = ( wire3318  &  wire33693 ) | ( n_n4501  &  wire33595  &  wire33693 ) ;
 assign wire2311 = ( wire3322  &  wire33695 ) | ( n_n4509  &  wire33475  &  wire33695 ) ;
 assign wire2313 = ( wire3341  &  wire33697 ) | ( n_n4433  &  wire33515  &  wire33697 ) ;
 assign wire2314 = ( wire3393  &  wire33698 ) | ( n_n4441  &  wire33555  &  wire33698 ) ;
 assign wire2317 = ( wire3308  &  wire33701 ) | ( (~ n_n5574)  &  wire33603  &  wire33701 ) ;
 assign wire2318 = ( wire3098  &  wire33704 ) | ( wire3099  &  wire33704 ) | ( wire33702  &  wire33704 ) ;
 assign wire2319 = ( wire1327  &  wire3206 ) | ( (~ n_n5520)  &  wire1327  &  wire33611 ) ;
 assign wire2320 = ( wire1324  &  wire3215 ) | ( (~ n_n5514)  &  wire1324  &  wire33608 ) ;
 assign wire2321 = ( pi19  &  ni30  &  wire507 ) ;
 assign wire2322 = ( ni30  &  wire913 ) ;
 assign wire2323 = ( wire614  &  wire3064 ) | ( wire614  &  wire33705 ) ;
 assign wire2324 = ( wire586  &  wire3193 ) | ( n_n4404  &  wire477  &  wire586 ) ;
 assign wire2325 = ( wire196  &  wire33630 ) | ( wire192  &  n_n4489  &  wire33630 ) ;
 assign wire2326 = ( wire196  &  wire33632 ) | ( wire192  &  n_n4481  &  wire33632 ) ;
 assign wire2327 = ( wire196  &  wire33634 ) | ( wire192  &  n_n4473  &  wire33634 ) ;
 assign wire2329 = ( wire196  &  wire33636 ) | ( wire192  &  n_n4509  &  wire33636 ) ;
 assign wire2330 = ( wire196  &  wire33637 ) | ( wire192  &  n_n4501  &  wire33637 ) ;
 assign wire2331 = ( wire196  &  wire33638 ) | ( wire192  &  n_n4412  &  wire33638 ) ;
 assign wire2332 = ( wire178  &  wire403  &  wire196 ) | ( wire178  &  wire403  &  wire2549 ) ;
 assign wire2333 = ( wire196  &  wire33640 ) | ( n_n4433  &  wire192  &  wire33640 ) ;
 assign wire2334 = ( wire196  &  wire33641 ) | ( wire192  &  n_n4441  &  wire33641 ) ;
 assign wire2335 = ( wire196  &  wire33642 ) | ( wire2406  &  wire33642 ) ;
 assign wire2336 = ( wire196  &  wire33643 ) | ( wire2404  &  wire33643 ) ;
 assign wire2341 = ( pi16  &  pi15  &  wire2562 ) | ( pi16  &  pi15  &  wire2563 ) ;
 assign wire2342 = ( wire416  &  wire196 ) | ( wire416  &  wire2547 ) ;
 assign wire2345 = ( wire196  &  wire33352 ) | ( wire2500  &  wire33352 ) ;
 assign wire2346 = ( wire196  &  wire33355 ) | ( wire192  &  n_n4611  &  wire33355 ) ;
 assign wire2348 = ( wire180  &  wire196  &  wire614 ) | ( wire180  &  wire614  &  wire2448 ) ;
 assign wire2349 = ( wire178  &  nv7129  &  wire614 ) ;
 assign wire2350 = ( wire196  &  wire33476 ) | ( wire2524  &  wire33476 ) ;
 assign wire2351 = ( wire182  &  wire196  &  wire507 ) | ( wire182  &  wire507  &  wire2474 ) ;
 assign wire2352 = ( wire179  &  wire196  &  wire507 ) | ( wire179  &  wire507  &  wire2469 ) ;
 assign wire2353 = ( wire196  &  wire33596 ) | ( wire2519  &  wire33596 ) ;
 assign wire2355 = ( nv7050  &  wire33605 ) ;
 assign wire2360 = ( wire196  &  wire586 ) | ( wire192  &  n_n4543  &  wire586 ) ;
 assign wire2364 = ( pi27  &  pi16  &  wire2456 ) | ( pi27  &  pi16  &  wire34164 ) ;
 assign wire2365 = ( (~ pi27)  &  pi16  &  wire640 ) ;
 assign wire2367 = ( pi27  &  wire657 ) ;
 assign wire2368 = ( (~ pi27)  &  wire2446 ) | ( (~ pi27)  &  wire34170 ) ;
 assign wire2370 = ( wire196  &  wire34128 ) | ( wire192  &  n_n4509  &  wire34128 ) ;
 assign wire2371 = ( wire2576  &  wire34130 ) | ( wire34063  &  wire34130 ) ;
 assign wire2374 = ( wire2409  &  wire34135 ) | ( wire34070  &  wire34135 ) ;
 assign wire2375 = ( wire196  &  wire34136 ) | ( wire192  &  n_n4501  &  wire34136 ) ;
 assign wire2378 = ( (~ pi21)  &  nv7445  &  wire34139 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire34139 ) ;
 assign wire2379 = ( (~ pi27)  &  (~ pi26)  &  wire2387 ) | ( (~ pi27)  &  (~ pi26)  &  wire34090 ) ;
 assign wire2380 = ( wire156  &  wire2389 ) | ( wire156  &  wire2390 ) | ( wire156  &  wire2391 ) ;
 assign wire2381 = ( (~ pi21)  &  wire158  &  nv7445 ) | ( pi21  &  (~ pi22)  &  wire158  &  nv7445 ) ;
 assign wire2382 = ( n_n4481  &  wire34082 ) ;
 assign wire2386 = ( pi17  &  (~ pi16)  &  nv7447  &  wire178 ) ;
 assign wire2387 = ( nv10153  &  wire2389 ) | ( nv10153  &  wire2390 ) | ( nv10153  &  wire2391 ) ;
 assign wire2389 = ( wire196  &  wire250 ) | ( wire192  &  n_n4489  &  wire250 ) ;
 assign wire2390 = ( wire196  &  wire243 ) | ( wire192  &  n_n4481  &  wire243 ) ;
 assign wire2391 = ( wire196  &  wire194 ) | ( wire192  &  n_n4473  &  wire194 ) ;
 assign wire2398 = ( (~ n_n5580)  &  wire1006  &  wire34075 ) | ( (~ n_n5580)  &  wire33599  &  wire34075 ) ;
 assign wire2399 = ( (~ n_n5574)  &  wire1006  &  wire34076 ) | ( (~ n_n5574)  &  wire33604  &  wire34076 ) ;
 assign wire2400 = ( pi20  &  nv7447  &  wire153 ) | ( (~ pi20)  &  nv7447  &  wire153 ) ;
 assign wire2402 = ( pi20  &  wire196  &  wire153 ) | ( pi20  &  wire153  &  wire2404 ) ;
 assign wire2403 = ( (~ pi20)  &  wire196  &  wire153 ) | ( (~ pi20)  &  wire153  &  wire2406 ) ;
 assign wire2404 = ( wire192  &  (~ n_n5574)  &  wire1006 ) | ( wire192  &  (~ n_n5574)  &  wire33604 ) ;
 assign wire2406 = ( wire192  &  (~ n_n5580)  &  wire1006 ) | ( wire192  &  (~ n_n5580)  &  wire33599 ) ;
 assign wire2409 = ( wire196  &  nv10153 ) | ( wire192  &  nv10153  &  n_n4501 ) ;
 assign wire2416 = ( wire34193  &  wire34238 ) | ( nv10153  &  wire527  &  wire34238 ) ;
 assign wire2418 = ( pi27  &  wire672 ) ;
 assign wire2419 = ( (~ pi27)  &  wire2498 ) | ( (~ pi27)  &  wire34198 ) ;
 assign wire2421 = ( wire196  &  wire34213 ) | ( n_n4433  &  wire192  &  wire34213 ) ;
 assign wire2422 = ( wire2571  &  wire34214 ) | ( wire34096  &  wire34214 ) ;
 assign wire2423 = ( pi27  &  pi16  &  wire2554 ) | ( pi27  &  pi16  &  wire34108 ) ;
 assign wire2424 = ( (~ pi27)  &  pi16  &  wire450 ) | ( (~ pi27)  &  pi16  &  wire2560 ) ;
 assign wire2426 = ( (~ pi27)  &  wire2545 ) | ( (~ pi27)  &  wire34111 ) ;
 assign wire2427 = ( pi27  &  wire653 ) ;
 assign wire2432 = ( wire2456  &  wire34289 ) | ( wire34164  &  wire34289 ) ;
 assign wire2433 = ( pi27  &  pi16  &  wire640 ) | ( (~ pi26)  &  pi16  &  wire640 ) ;
 assign wire2435 = ( (~ pi27)  &  pi26  &  wire657 ) ;
 assign wire2436 = ( pi27  &  wire2446 ) | ( (~ pi26)  &  wire2446 ) | ( pi27  &  wire34170 ) | ( (~ pi26)  &  wire34170 ) ;
 assign wire2437 = ( (~ pi21)  &  nv7791  &  wire154 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire154 ) ;
 assign wire2438 = ( wire3189  &  wire34167 ) | ( n_n4412  &  wire33395  &  wire34167 ) ;
 assign wire2442 = ( pi17  &  pi16  &  nv7447  &  wire178 ) ;
 assign wire2446 = ( wire180  &  wire196  &  wire154 ) | ( wire180  &  wire154  &  wire2448 ) ;
 assign wire2447 = ( wire196  &  wire183 ) | ( wire192  &  n_n4543  &  wire183 ) ;
 assign wire2448 = ( wire192  &  wire3189 ) | ( wire192  &  n_n4412  &  wire33395 ) ;
 assign wire2456 = ( wire196  &  wire34158 ) | ( wire2469  &  wire34158 ) ;
 assign wire2457 = ( wire3393  &  wire34159 ) | ( n_n4441  &  wire33555  &  wire34159 ) ;
 assign wire2460 = ( (~ pi17)  &  nv7447  &  wire179 ) ;
 assign wire2469 = ( wire192  &  wire3393 ) | ( wire192  &  n_n4441  &  wire33555 ) ;
 assign wire2471 = ( wire192  &  wire3341 ) | ( n_n4433  &  wire192  &  wire33515 ) ;
 assign wire2472 = ( wire196  &  nv10153 ) | ( nv10153  &  wire2474 ) ;
 assign wire2474 = ( wire192  &  wire3341 ) | ( n_n4433  &  wire192  &  wire33515 ) ;
 assign wire2478 = ( n_n3349  &  wire34302 ) | ( n_n3347  &  wire204  &  wire34302 ) ;
 assign wire2479 = ( pi21  &  (~ pi20)  &  n_n3347  &  wire698 ) ;
 assign wire2482 = ( (~ pi21)  &  nv7791  &  wire34306 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire34306 ) ;
 assign wire2484 = ( wire34193  &  wire34308 ) | ( nv10153  &  wire527  &  wire34308 ) ;
 assign wire2485 = ( (~ pi21)  &  wire158  &  nv7791 ) | ( pi21  &  (~ pi22)  &  wire158  &  nv7791 ) ;
 assign wire2486 = ( (~ pi27)  &  pi26  &  wire672 ) ;
 assign wire2487 = ( pi27  &  wire2498 ) | ( (~ pi26)  &  wire2498 ) | ( pi27  &  wire34198 ) | ( (~ pi26)  &  wire34198 ) ;
 assign wire2490 = ( wire3251  &  wire34195 ) | ( n_n4481  &  wire33350  &  wire34195 ) ;
 assign wire2491 = ( wire3280  &  wire34196 ) | ( n_n4489  &  wire33307  &  wire34196 ) ;
 assign wire2494 = ( pi17  &  (~ pi16)  &  nv7447  &  wire178 ) ;
 assign wire2498 = ( wire158  &  wire180  &  wire196 ) | ( wire158  &  wire180  &  wire2500 ) ;
 assign wire2499 = ( wire196  &  wire194 ) | ( wire192  &  n_n4611  &  wire194 ) ;
 assign wire2500 = ( wire192  &  wire3251 ) | ( wire192  &  n_n4481  &  wire33350 ) ;
 assign wire2502 = ( wire192  &  wire3280 ) | ( wire192  &  n_n4489  &  wire33307 ) ;
 assign wire2508 = ( pi20  &  nv7447  &  wire153 ) | ( (~ pi20)  &  nv7447  &  wire153 ) ;
 assign wire2516 = ( wire192  &  wire3318 ) | ( wire192  &  n_n4501  &  wire33595 ) ;
 assign wire2517 = ( wire196  &  nv10153 ) | ( nv10153  &  wire2519 ) ;
 assign wire2519 = ( wire192  &  wire3318 ) | ( wire192  &  n_n4501  &  wire33595 ) ;
 assign wire2521 = ( wire192  &  wire3322 ) | ( wire192  &  n_n4509  &  wire33475 ) ;
 assign wire2522 = ( wire196  &  nv10153 ) | ( nv10153  &  wire2524 ) ;
 assign wire2524 = ( wire192  &  wire3322 ) | ( wire192  &  n_n4509  &  wire33475 ) ;
 assign wire2526 = ( wire196  &  wire34320 ) | ( n_n4433  &  wire192  &  wire34320 ) ;
 assign wire2527 = ( wire2571  &  wire34322 ) | ( wire34096  &  wire34322 ) ;
 assign wire2529 = ( wire2554  &  wire34324 ) | ( wire34108  &  wire34324 ) ;
 assign wire2530 = ( wire2560  &  wire34325 ) | ( wire2562  &  wire34325 ) | ( wire2563  &  wire34325 ) ;
 assign wire2531 = ( pi16  &  wire1306 ) ;
 assign wire2532 = ( pi27  &  wire2545 ) | ( (~ pi26)  &  wire2545 ) | ( pi27  &  wire34111 ) | ( (~ pi26)  &  wire34111 ) ;
 assign wire2533 = ( (~ pi27)  &  pi26  &  wire653 ) ;
 assign wire2534 = ( (~ pi21)  &  nv7791  &  wire154 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire154 ) ;
 assign wire2538 = ( wire721  &  wire33433  &  wire34113 ) | ( wire721  &  wire33434  &  wire34113 ) ;
 assign wire2545 = ( wire196  &  wire244 ) | ( wire192  &  n_n4412  &  wire244 ) ;
 assign wire2546 = ( wire152  &  wire196  &  wire154 ) | ( wire152  &  wire154  &  wire2547 ) ;
 assign wire2547 = ( ni33  &  n_n4404 ) | ( (~ ni29)  &  n_n4404 ) | ( n_n4404  &  (~ nv6462) ) ;
 assign wire2549 = ( wire721  &  wire192  &  wire33433 ) | ( wire721  &  wire192  &  wire33434 ) ;
 assign wire2553 = ( wire1006  &  (~ n_n5520)  &  wire34100 ) | ( (~ n_n5520)  &  wire33612  &  wire34100 ) ;
 assign wire2554 = ( wire196  &  wire34101 ) | ( wire192  &  n_n4441  &  wire34101 ) ;
 assign wire2556 = ( (~ n_n5514)  &  wire1006  &  wire34103 ) | ( (~ n_n5514)  &  wire33609  &  wire34103 ) ;
 assign wire2557 = ( pi20  &  nv7447  &  wire153 ) | ( (~ pi20)  &  nv7447  &  wire153 ) ;
 assign wire2558 = ( nv10153  &  wire2562 ) | ( nv10153  &  wire2563 ) ;
 assign wire2559 = ( (~ pi17)  &  nv7447  &  wire179 ) ;
 assign wire2560 = ( wire196  &  wire199 ) | ( wire192  &  n_n4441  &  wire199 ) ;
 assign wire2562 = ( pi20  &  wire196  &  wire153 ) | ( pi20  &  wire153  &  wire2566 ) ;
 assign wire2563 = ( (~ pi20)  &  wire196  &  wire153 ) | ( (~ pi20)  &  wire153  &  wire2564 ) ;
 assign wire2564 = ( wire192  &  wire1006  &  (~ n_n5520) ) | ( wire192  &  (~ n_n5520)  &  wire33612 ) ;
 assign wire2566 = ( wire192  &  (~ n_n5514)  &  wire1006 ) | ( wire192  &  (~ n_n5514)  &  wire33609 ) ;
 assign wire2571 = ( wire196  &  nv10153 ) | ( n_n4433  &  wire192  &  nv10153 ) ;
 assign wire2576 = ( wire196  &  nv10153 ) | ( wire192  &  n_n4509  &  nv10153 ) ;
 assign wire2585 = ( wire268  &  wire422  &  wire34354 ) ;
 assign wire2586 = ( wire837  &  wire3139  &  wire34356 ) | ( wire837  &  wire3140  &  wire34356 ) ;
 assign wire2587 = ( (~ ni14)  &  n_n3695  &  wire34357 ) | ( (~ ni14)  &  n_n3693  &  wire34357 ) ;
 assign wire2591 = ( pi23  &  wire912  &  wire3125 ) | ( pi23  &  wire912  &  wire3126 ) ;
 assign wire2593 = ( (~ ni11)  &  wire2614 ) | ( (~ ni11)  &  wire2615 ) | ( (~ ni11)  &  wire34523 ) ;
 assign wire2594 = ( wire2967  &  wire34369 ) | ( wire34365  &  wire34369 ) ;
 assign wire2595 = ( wire197  &  wire34373 ) | ( wire193  &  n_n4509  &  wire34373 ) ;
 assign wire2596 = ( wire3034  &  wire34377 ) | ( wire34374  &  wire34377 ) ;
 assign wire2597 = ( wire197  &  wire34380 ) | ( n_n4433  &  wire193  &  wire34380 ) ;
 assign wire2600 = ( wire369  &  wire2635  &  wire34387 ) | ( wire369  &  wire2636  &  wire34387 ) ;
 assign wire2602 = ( wire369  &  wire2955  &  wire34407 ) | ( wire369  &  wire34406  &  wire34407 ) ;
 assign wire2603 = ( wire2961  &  wire34410 ) | ( wire2962  &  wire34410 ) | ( wire2963  &  wire34410 ) ;
 assign wire2604 = ( wire2964  &  wire34412 ) | ( wire3195  &  wire34412 ) | ( wire3196  &  wire34412 ) ;
 assign wire2606 = ( n_n3016  &  wire185  &  wire34415 ) | ( wire185  &  wire3144  &  wire34415 ) ;
 assign wire2607 = ( wire2935  &  wire34417 ) | ( wire2936  &  wire34417 ) | ( wire2937  &  wire34417 ) ;
 assign wire2608 = ( wire2928  &  wire34426 ) | ( wire2933  &  wire34426 ) | ( wire34424  &  wire34426 ) ;
 assign wire2609 = ( wire161  &  wire369  &  wire2946 ) | ( wire161  &  wire369  &  wire34427 ) ;
 assign wire2614 = ( wire370  &  wire34472 ) | ( (~ wire161)  &  wire370  &  wire655 ) ;
 assign wire2615 = ( wire370  &  wire34503 ) | ( wire370  &  wire34504 ) ;
 assign wire2618 = ( wire2635  &  wire34445 ) | ( wire2636  &  wire34445 ) ;
 assign wire2619 = ( wire3023  &  wire34455 ) | ( wire34454  &  wire34455 ) ;
 assign wire2620 = ( pi16  &  pi23  &  wire501 ) | ( pi16  &  pi24  &  wire501 ) ;
 assign wire2621 = ( pi16  &  n_n3016  &  wire185 ) | ( pi16  &  wire185  &  wire3144 ) ;
 assign wire2622 = ( pi23  &  wire3019 ) | ( pi24  &  wire3019 ) | ( pi23  &  wire34457 ) | ( pi24  &  wire34457 ) ;
 assign wire2624 = ( pi17  &  pi16  &  n_n3016 ) | ( pi17  &  pi16  &  wire3144 ) ;
 assign wire2625 = ( nv8372  &  wire34475 ) | ( wire3000  &  wire34475 ) | ( wire3001  &  wire34475 ) ;
 assign wire2629 = ( wire2635  &  wire34486 ) | ( wire2636  &  wire34486 ) ;
 assign wire2631 = ( (~ pi16)  &  n_n3016  &  wire185 ) | ( (~ pi16)  &  wire185  &  wire3144 ) ;
 assign wire2632 = ( pi23  &  wire2994 ) | ( pi24  &  wire2994 ) | ( pi23  &  wire34488 ) | ( pi24  &  wire34488 ) ;
 assign wire2634 = ( pi17  &  (~ pi16)  &  n_n3016 ) | ( pi17  &  (~ pi16)  &  wire3144 ) ;
 assign wire2635 = ( wire211  &  wire3147 ) | ( wire211  &  nv8372  &  wire33940 ) ;
 assign wire2636 = ( pi20  &  wire3149 ) | ( pi20  &  nv8372  &  wire33939 ) ;
 assign wire2637 = ( wire3341  &  wire34536 ) | ( n_n4433  &  wire33515  &  wire34536 ) ;
 assign wire2639 = ( wire3189  &  wire34540 ) | ( n_n4412  &  wire33395  &  wire34540 ) ;
 assign wire2640 = ( wire2686  &  wire34542 ) | ( wire152  &  wire248  &  wire34542 ) ;
 assign wire2641 = ( wire345  &  wire3185  &  wire34543 ) | ( wire345  &  wire3186  &  wire34543 ) ;
 assign wire2642 = ( (~ pi15)  &  wire359  &  wire34557 ) | ( (~ pi15)  &  wire359  &  wire34558 ) ;
 assign wire2643 = ( pi15  &  wire359  &  wire34579 ) | ( pi15  &  wire359  &  wire34580 ) ;
 assign wire2645 = ( wire258  &  wire1298  &  wire359 ) | ( wire258  &  wire359  &  wire3060 ) ;
 assign wire2646 = ( wire2684  &  wire34584 ) | ( wire151  &  wire248  &  wire34584 ) ;
 assign wire2648 = ( wire2688  &  wire34586 ) | ( wire153  &  wire248  &  wire34586 ) ;
 assign wire2649 = ( wire818  &  wire2750 ) | ( wire818  &  wire34709 ) | ( wire818  &  wire34710 ) ;
 assign wire2652 = ( wire3318  &  wire34545 ) | ( n_n4501  &  wire33595  &  wire34545 ) ;
 assign wire2653 = ( wire3322  &  wire34547 ) | ( n_n4509  &  wire33475  &  wire34547 ) ;
 assign wire2654 = ( wire2686  &  wire34548 ) | ( wire152  &  wire248  &  wire34548 ) ;
 assign wire2655 = ( wire3251  &  wire34549 ) | ( n_n4481  &  wire33350  &  wire34549 ) ;
 assign wire2657 = ( (~ pi16)  &  wire3096 ) | ( (~ pi16)  &  wire3097 ) ;
 assign wire2658 = ( wire158  &  wire2684 ) | ( wire158  &  wire151  &  wire248 ) ;
 assign wire2659 = ( (~ pi16)  &  wire2688 ) | ( (~ pi16)  &  wire153  &  wire248 ) ;
 assign wire2668 = ( pi16  &  wire1320 ) | ( pi16  &  wire3104 ) ;
 assign wire2669 = ( (~ pi17)  &  pi16  &  wire358  &  n_n4441 ) ;
 assign wire2671 = ( pi17  &  wire2684 ) | ( pi17  &  wire151  &  wire248 ) ;
 assign wire2672 = ( (~ pi17)  &  wire2686 ) | ( (~ pi17)  &  wire152  &  wire248 ) ;
 assign wire2674 = ( (~ pi17)  &  (~ pi16)  &  n_n4509  &  wire358 ) ;
 assign wire2675 = ( (~ pi16)  &  wire3111 ) | ( (~ pi16)  &  wire3112 ) ;
 assign wire2676 = ( (~ pi21)  &  nv7647  &  wire257 ) | ( pi21  &  (~ pi22)  &  nv7647  &  wire257 ) ;
 assign wire2681 = ( (~ pi21)  &  nv7647  &  wire295 ) | ( pi21  &  (~ pi22)  &  nv7647  &  wire295 ) ;
 assign wire2684 = ( (~ pi19)  &  (~ pi21)  &  nv7647 ) | ( (~ pi19)  &  pi21  &  (~ pi22)  &  nv7647 ) ;
 assign wire2686 = ( pi19  &  (~ pi21)  &  nv7647 ) | ( pi19  &  pi21  &  (~ pi22)  &  nv7647 ) ;
 assign wire2688 = ( (~ pi21)  &  nv7647  &  wire163 ) | ( pi21  &  (~ pi22)  &  nv7647  &  wire163 ) ;
 assign wire2691 = ( wire197  &  wire33779 ) | ( wire3320  &  wire33779 ) ;
 assign wire2692 = ( wire197  &  wire33782 ) | ( n_n4433  &  wire193  &  wire33782 ) ;
 assign wire2694 = ( pi20  &  wire369  &  wire351  &  wire33786 ) ;
 assign wire2695 = ( wire3092  &  wire33789 ) | ( (~ pi20)  &  wire351  &  wire33789 ) ;
 assign wire2696 = ( (~ pi25)  &  (~ pi16)  &  wire370  &  wire641 ) ;
 assign wire2697 = ( wire2964  &  wire33793 ) | ( wire3195  &  wire33793 ) | ( wire3196  &  wire33793 ) ;
 assign wire2698 = ( wire197  &  wire33795 ) | ( wire3233  &  wire33795 ) ;
 assign wire2699 = ( wire369  &  wire3439  &  wire33797 ) | ( wire369  &  wire33796  &  wire33797 ) ;
 assign wire2700 = ( wire740  &  wire33799 ) | ( n_n4441  &  wire475  &  wire33799 ) ;
 assign wire2701 = ( (~ pi16)  &  wire370  &  wire727 ) | ( (~ pi16)  &  wire370  &  wire3088 ) ;
 assign wire2702 = ( wire370  &  wire1113  &  wire3246 ) | ( wire370  &  wire1113  &  wire33802 ) ;
 assign wire2704 = ( wire3098  &  wire33805 ) | ( wire3099  &  wire33805 ) | ( wire33702  &  wire33805 ) ;
 assign wire2705 = ( wire3083  &  wire33806 ) | ( wire3084  &  wire33806 ) | ( wire3085  &  wire33806 ) ;
 assign wire2706 = ( wire3083  &  wire33807 ) | ( wire3084  &  wire33807 ) | ( wire3085  &  wire33807 ) ;
 assign wire2707 = ( pi16  &  wire369  &  wire3056 ) | ( pi16  &  wire369  &  wire3057 ) ;
 assign wire2708 = ( wire369  &  wire918 ) | ( wire476  &  wire369  &  n_n4834 ) ;
 assign wire2710 = ( wire369  &  wire3069 ) | ( wire154  &  wire369  &  wire443 ) ;
 assign wire2711 = ( wire370  &  wire2718 ) | ( wire370  &  wire33824 ) | ( wire370  &  wire33825 ) ;
 assign wire2713 = ( wire197  &  wire1028  &  wire33809 ) | ( wire1028  &  wire3339  &  wire33809 ) ;
 assign wire2714 = ( wire3341  &  wire33812 ) | ( n_n4433  &  wire33515  &  wire33812 ) ;
 assign wire2715 = ( pi20  &  wire351  &  wire33813 ) ;
 assign wire2717 = ( pi16  &  wire1298 ) | ( pi16  &  wire3058 ) | ( pi16  &  wire3060 ) ;
 assign wire2718 = ( (~ pi25)  &  wire3179 ) | ( (~ pi25)  &  wire33818 ) ;
 assign wire2719 = ( pi16  &  wire3083 ) | ( pi16  &  wire3084 ) | ( pi16  &  wire3085 ) ;
 assign wire2720 = ( pi16  &  wire3057 ) | ( pi16  &  wire173  &  wire616 ) ;
 assign wire2723 = ( wire351  &  wire33827 ) ;
 assign wire2724 = ( wire197  &  wire33828 ) | ( wire193  &  n_n4509  &  wire33828 ) ;
 assign wire2729 = ( (~ pi16)  &  wire3083 ) | ( (~ pi16)  &  wire3084 ) | ( (~ pi16)  &  wire3085 ) ;
 assign wire2730 = ( pi25  &  (~ pi16)  &  wire3114 ) | ( pi25  &  (~ pi16)  &  wire33682 ) ;
 assign wire2731 = ( wire1113  &  wire3221 ) | ( wire1113  &  wire3222 ) | ( wire1113  &  wire33831 ) ;
 assign wire2732 = ( (~ pi25)  &  (~ pi16)  &  wire2961 ) | ( (~ pi25)  &  (~ pi16)  &  wire33833 ) ;
 assign wire2733 = ( wire3341  &  wire34590 ) | ( n_n4433  &  wire33515  &  wire34590 ) ;
 assign wire2734 = ( wire3189  &  wire34593 ) | ( n_n4412  &  wire33395  &  wire34593 ) ;
 assign wire2735 = ( wire2812  &  wire34595  &  wire34596 ) | ( wire34594  &  wire34595  &  wire34596 ) ;
 assign wire2736 = ( wire3215  &  wire34600 ) | ( (~ n_n5514)  &  wire33608  &  wire34600 ) ;
 assign wire2739 = ( wire2805  &  wire34606 ) | ( wire179  &  wire273  &  wire34606 ) ;
 assign wire2741 = ( wire219  &  wire3205  &  wire34609 ) | ( wire219  &  wire3206  &  wire34609 ) ;
 assign wire2742 = ( wire345  &  wire3185  &  wire34610 ) | ( wire345  &  wire3186  &  wire34610 ) ;
 assign wire2743 = ( wire2800  &  wire34612 ) | ( wire2801  &  wire34612 ) | ( wire2802  &  wire34612 ) ;
 assign wire2744 = ( (~ pi21)  &  nv7445  &  wire34613 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire34613 ) ;
 assign wire2745 = ( wire2803  &  wire34614 ) | ( wire178  &  wire273  &  wire34614 ) ;
 assign wire2750 = ( (~ pi15)  &  (~ ni14)  &  wire34694 ) | ( (~ pi15)  &  (~ ni14)  &  wire34695 ) ;
 assign wire2752 = ( wire2812  &  wire34620 ) | ( wire34594  &  wire34620 ) ;
 assign wire2753 = ( n_n4412  &  wire181  &  wire34621 ) ;
 assign wire2754 = ( (~ n_n5514)  &  wire1006  &  wire34624 ) | ( (~ n_n5514)  &  wire33609  &  wire34624 ) ;
 assign wire2755 = ( (~ pi17)  &  pi16  &  wire358  &  n_n4441 ) ;
 assign wire2756 = ( wire2805  &  wire34626 ) | ( wire179  &  wire273  &  wire34626 ) ;
 assign wire2761 = ( pi16  &  wire2800 ) | ( pi16  &  wire2801 ) | ( pi16  &  wire2802 ) ;
 assign wire2762 = ( wire154  &  wire2803 ) | ( wire178  &  wire154  &  wire273 ) ;
 assign wire2764 = ( (~ pi21)  &  nv7445  &  wire257 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire257 ) ;
 assign wire2767 = ( (~ pi16)  &  n_n3693  &  wire817 ) ;
 assign wire2770 = ( (~ n_n5574)  &  wire1006  &  wire34647 ) | ( (~ n_n5574)  &  wire33604  &  wire34647 ) ;
 assign wire2771 = ( (~ n_n5580)  &  wire1006  &  wire34648 ) | ( (~ n_n5580)  &  wire33599  &  wire34648 ) ;
 assign wire2772 = ( pi25  &  wire158  &  wire180  &  n_n4481 ) ;
 assign wire2775 = ( (~ pi19)  &  (~ pi16)  &  n_n3695 ) ;
 assign wire2777 = ( (~ pi17)  &  (~ pi16)  &  n_n4509  &  wire358 ) ;
 assign wire2778 = ( wire302  &  wire2805 ) | ( wire302  &  wire179  &  wire273 ) ;
 assign wire2780 = ( wire1293  &  wire2812 ) | ( wire1293  &  wire34594 ) ;
 assign wire2781 = ( (~ pi25)  &  wire294  &  wire3139 ) | ( (~ pi25)  &  wire294  &  wire3140 ) ;
 assign wire2784 = ( wire3318  &  wire34671 ) | ( n_n4501  &  wire33595  &  wire34671 ) ;
 assign wire2785 = ( wire2812  &  wire34673 ) | ( wire34594  &  wire34673 ) ;
 assign wire2786 = ( wire3322  &  wire34675 ) | ( n_n4509  &  wire33475  &  wire34675 ) ;
 assign wire2787 = ( wire3251  &  wire34677 ) | ( n_n4481  &  wire33350  &  wire34677 ) ;
 assign wire2788 = ( wire3308  &  wire34679 ) | ( (~ n_n5574)  &  wire33603  &  wire34679 ) ;
 assign wire2789 = ( wire2805  &  wire34680 ) | ( wire179  &  wire273  &  wire34680 ) ;
 assign wire2792 = ( wire3327  &  wire34683 ) | ( (~ n_n5580)  &  wire33598  &  wire34683 ) ;
 assign wire2794 = ( (~ pi16)  &  wire2800 ) | ( (~ pi16)  &  wire2801 ) | ( (~ pi16)  &  wire2802 ) ;
 assign wire2795 = ( wire158  &  wire2803 ) | ( wire158  &  wire178  &  wire273 ) ;
 assign wire2798 = ( (~ pi21)  &  nv7445  &  wire295 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire295 ) ;
 assign wire2800 = ( n_n3695  &  wire163 ) | ( n_n3693  &  wire163  &  wire204 ) ;
 assign wire2801 = ( (~ pi20)  &  pi25  &  nv7445  &  wire153 ) ;
 assign wire2802 = ( (~ pi25)  &  wire169  &  wire3139 ) | ( (~ pi25)  &  wire169  &  wire3140 ) ;
 assign wire2803 = ( (~ pi19)  &  n_n3695 ) | ( (~ pi19)  &  n_n3693  &  wire204 ) ;
 assign wire2805 = ( pi19  &  n_n3695 ) | ( pi19  &  n_n3693  &  wire204 ) ;
 assign wire2811 = ( ni30  &  wire156  &  wire181 ) | ( (~ wire156)  &  nv7447  &  wire181 ) ;
 assign wire2812 = ( (~ pi25)  &  (~ wire150)  &  wire3139 ) | ( (~ pi25)  &  (~ wire150)  &  wire3140 ) ;
 assign wire2815 = ( wire268  &  (~ wire793)  &  wire422  &  wire34820 ) ;
 assign wire2816 = ( wire3157  &  wire34825 ) | ( wire3158  &  wire34825 ) ;
 assign wire2817 = ( wire3150  &  wire34828 ) | ( wire3151  &  wire34828 ) ;
 assign wire2818 = ( wire2892  &  wire34831 ) | ( wire33914  &  wire34831 ) ;
 assign wire2819 = ( wire837  &  wire3139  &  wire34833 ) | ( wire837  &  wire3140  &  wire34833 ) ;
 assign wire2820 = ( (~ ni14)  &  n_n3695  &  wire34835 ) | ( (~ ni14)  &  n_n3693  &  wire34835 ) ;
 assign wire2821 = ( wire2906  &  wire34837 ) | ( wire2907  &  wire34837 ) ;
 assign wire2822 = ( wire2884  &  wire34839 ) | ( wire2885  &  wire34839 ) | ( wire2886  &  wire34839 ) ;
 assign wire2826 = ( wire912  &  wire3125  &  wire34850 ) | ( wire912  &  wire3126  &  wire34850 ) ;
 assign wire2828 = ( wire2850  &  wire34931 ) | ( wire2851  &  wire34931 ) | ( wire34929  &  wire34931 ) ;
 assign wire2830 = ( ni9  &  (~ ni8)  &  nv8350 ) ;
 assign wire2831 = ( wire197  &  wire34853 ) | ( n_n4433  &  wire193  &  wire34853 ) ;
 assign wire2832 = ( wire3034  &  wire34855 ) | ( wire34374  &  wire34855 ) ;
 assign wire2833 = ( wire2967  &  wire34857 ) | ( wire34365  &  wire34857 ) ;
 assign wire2834 = ( wire197  &  wire34859 ) | ( wire193  &  n_n4509  &  wire34859 ) ;
 assign wire2838 = ( wire369  &  wire2955  &  wire34866 ) | ( wire369  &  wire34406  &  wire34866 ) ;
 assign wire2839 = ( wire2961  &  wire34869 ) | ( wire2962  &  wire34869 ) | ( wire2963  &  wire34869 ) ;
 assign wire2840 = ( wire2964  &  wire34871 ) | ( wire3195  &  wire34871 ) | ( wire3196  &  wire34871 ) ;
 assign wire2841 = ( wire369  &  wire1031  &  wire2876 ) | ( wire369  &  wire1031  &  wire2877 ) ;
 assign wire2842 = ( wire369  &  wire698  &  wire2865 ) | ( wire369  &  wire698  &  wire2866 ) ;
 assign wire2845 = ( wire2935  &  wire34876 ) | ( wire2936  &  wire34876 ) | ( wire2937  &  wire34876 ) ;
 assign wire2846 = ( wire2928  &  wire34877 ) | ( wire2933  &  wire34877 ) | ( wire34424  &  wire34877 ) ;
 assign wire2847 = ( wire160  &  wire369  &  wire2946 ) | ( wire160  &  wire369  &  wire34427 ) ;
 assign wire2850 = ( wire370  &  wire2863 ) | ( wire370  &  wire34894 ) | ( wire370  &  wire34895 ) ;
 assign wire2851 = ( wire370  &  wire34911 ) | ( (~ wire160)  &  wire370  &  wire655 ) ;
 assign wire2852 = ( nv8372  &  wire34846 ) | ( (~ wire157)  &  (~ nv6462)  &  wire34846 ) ;
 assign wire2855 = ( nv8372  &  wire34881 ) | ( wire2983  &  wire34881 ) | ( wire2984  &  wire34881 ) ;
 assign wire2857 = ( nv8372  &  wire34884 ) | ( wire3000  &  wire34884 ) | ( wire3001  &  wire34884 ) ;
 assign wire2858 = ( wire2865  &  wire34885 ) | ( wire2866  &  wire34885 ) ;
 assign wire2860 = ( wire34483  &  wire34887 ) | ( nv10167  &  wire447  &  wire34887 ) ;
 assign wire2861 = ( n_n2546  &  wire34888 ) | ( wire2878  &  wire34888 ) ;
 assign wire2862 = ( (~ pi23)  &  wire2994 ) | ( pi24  &  wire2994 ) | ( (~ pi23)  &  wire34488 ) | ( pi24  &  wire34488 ) ;
 assign wire2863 = ( pi23  &  (~ pi24)  &  wire673 ) ;
 assign wire2864 = ( pi17  &  (~ pi16)  &  n_n2546 ) | ( pi17  &  (~ pi16)  &  wire2878 ) ;
 assign wire2865 = ( wire204  &  wire2883 ) | ( nv8372  &  wire204  &  wire34845 ) ;
 assign wire2866 = ( (~ pi20)  &  wire2881 ) | ( (~ pi20)  &  nv8372  &  wire34844 ) ;
 assign wire2869 = ( wire2876  &  wire34901 ) | ( wire2877  &  wire34901 ) ;
 assign wire2870 = ( wire3023  &  wire34902 ) | ( wire34454  &  wire34902 ) ;
 assign wire2871 = ( pi16  &  (~ pi23)  &  wire501 ) | ( pi16  &  pi24  &  wire501 ) ;
 assign wire2872 = ( n_n2546  &  wire34904 ) | ( wire2878  &  wire34904 ) ;
 assign wire2873 = ( (~ pi23)  &  wire3019 ) | ( pi24  &  wire3019 ) | ( (~ pi23)  &  wire34457 ) | ( pi24  &  wire34457 ) ;
 assign wire2875 = ( pi17  &  pi16  &  n_n2546 ) | ( pi17  &  pi16  &  wire2878 ) ;
 assign wire2876 = ( wire211  &  wire2883 ) | ( wire211  &  nv8372  &  wire34845 ) ;
 assign wire2877 = ( pi20  &  wire2881 ) | ( pi20  &  nv8372  &  wire34844 ) ;
 assign wire2878 = ( pi21  &  wire2883 ) | ( pi21  &  nv8372  &  wire34845 ) ;
 assign wire2881 = ( (~ pi21)  &  (~ pi23)  &  ni30 ) | ( (~ pi21)  &  pi24  &  ni30 ) ;
 assign wire2883 = ( (~ pi22)  &  (~ pi23)  &  ni30 ) | ( (~ pi22)  &  pi24  &  ni30 ) ;
 assign wire2884 = ( nv8372  &  wire34361 ) | ( (~ wire157)  &  (~ nv6462)  &  wire34361 ) ;
 assign wire2885 = ( nv8608  &  wire1299 ) | ( wire1299  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire2886 = ( pi24  &  wire3125 ) | ( pi24  &  wire3126 ) ;
 assign wire2889 = ( pi24  &  ni30  &  wire156 ) | ( pi24  &  (~ wire156)  &  nv7447 ) ;
 assign wire2892 = ( pi24  &  ni30  &  wire155 ) | ( pi24  &  (~ wire155)  &  nv7447 ) ;
 assign wire2893 = ( (~ wire156)  &  wire818  &  wire921  &  wire34726 ) ;
 assign wire2894 = ( wire156  &  wire822  &  wire818  &  wire921 ) ;
 assign wire2895 = ( wire359  &  wire3125  &  wire34731 ) | ( wire359  &  wire3126  &  wire34731 ) ;
 assign wire2896 = ( wire837  &  wire3139  &  wire34733 ) | ( wire837  &  wire3140  &  wire34733 ) ;
 assign wire2897 = ( (~ ni14)  &  n_n3695  &  wire34734 ) | ( (~ ni14)  &  n_n3693  &  wire34734 ) ;
 assign wire2898 = ( wire2906  &  wire34735 ) | ( wire2907  &  wire34735 ) ;
 assign wire2899 = ( (~ pi24)  &  wire359  &  wire597 ) ;
 assign wire2900 = ( pi24  &  wire359  &  wire422 ) ;
 assign wire2901 = ( (~ wire157)  &  (~ nv6462)  &  wire1044  &  wire359 ) ;
 assign wire2902 = ( (~ ni11)  &  wire2926 ) | ( (~ ni11)  &  wire2927 ) | ( (~ ni11)  &  wire34795 ) ;
 assign wire2906 = ( nv8608  &  wire34358 ) | ( (~ wire157)  &  (~ nv6462)  &  wire34358 ) ;
 assign wire2907 = ( nv8372  &  wire34359 ) | ( (~ wire157)  &  (~ nv6462)  &  wire34359 ) ;
 assign wire2910 = ( (~ wire1090)  &  wire2967  &  wire34739 ) | ( (~ wire1090)  &  wire34365  &  wire34739 ) ;
 assign wire2911 = ( wire197  &  wire34742 ) | ( wire193  &  n_n4509  &  wire34742 ) ;
 assign wire2912 = ( wire197  &  wire34744 ) | ( n_n4433  &  wire193  &  wire34744 ) ;
 assign wire2913 = ( wire828  &  wire3034  &  wire34745 ) | ( wire828  &  wire34374  &  wire34745 ) ;
 assign wire2915 = ( wire369  &  wire2955  &  wire34749 ) | ( wire369  &  wire34406  &  wire34749 ) ;
 assign wire2916 = ( wire2961  &  wire34752 ) | ( wire2962  &  wire34752 ) | ( wire2963  &  wire34752 ) ;
 assign wire2917 = ( wire2964  &  wire34754 ) | ( wire3195  &  wire34754 ) | ( wire3196  &  wire34754 ) ;
 assign wire2918 = ( wire2935  &  wire34755 ) | ( wire2936  &  wire34755 ) | ( wire2937  &  wire34755 ) ;
 assign wire2919 = ( pi24  &  wire369  &  wire2933 ) | ( pi24  &  wire369  &  wire34425 ) ;
 assign wire2920 = ( (~ pi24)  &  wire369  &  wire2946 ) | ( (~ pi24)  &  wire369  &  wire34427 ) ;
 assign wire2926 = ( wire370  &  wire34769 ) | ( wire370  &  wire34770 ) ;
 assign wire2927 = ( wire370  &  wire34780 ) | ( pi24  &  wire370  &  wire655 ) ;
 assign wire2928 = ( n_n4481  &  wire34418 ) ;
 assign wire2932 = ( pi17  &  (~ pi16)  &  wire178  &  nv8372 ) ;
 assign wire2933 = ( nv10167  &  wire2935 ) | ( nv10167  &  wire2936 ) | ( nv10167  &  wire2937 ) ;
 assign wire2935 = ( wire197  &  wire250 ) | ( n_n4489  &  wire193  &  wire250 ) ;
 assign wire2936 = ( wire197  &  wire243 ) | ( wire193  &  n_n4481  &  wire243 ) ;
 assign wire2937 = ( wire197  &  wire194 ) | ( wire193  &  n_n4473  &  wire194 ) ;
 assign wire2939 = ( wire721  &  wire33433  &  wire34430 ) | ( wire721  &  wire33434  &  wire34430 ) ;
 assign wire2946 = ( wire197  &  wire244 ) | ( n_n4412  &  wire193  &  wire244 ) ;
 assign wire2947 = ( wire152  &  wire197  &  wire154 ) | ( wire152  &  wire154  &  wire3233 ) ;
 assign wire2949 = ( (~ n_n5580)  &  wire1006  &  wire34390 ) | ( (~ n_n5580)  &  wire33599  &  wire34390 ) ;
 assign wire2950 = ( (~ n_n5574)  &  wire1006  &  wire34391 ) | ( (~ n_n5574)  &  wire33604  &  wire34391 ) ;
 assign wire2951 = ( pi20  &  nv8372  &  wire153 ) | ( (~ pi20)  &  nv8372  &  wire153 ) ;
 assign wire2952 = ( (~ pi17)  &  wire182  &  nv8372 ) ;
 assign wire2954 = ( wire1006  &  (~ n_n5520)  &  wire34398 ) | ( (~ n_n5520)  &  wire33612  &  wire34398 ) ;
 assign wire2955 = ( wire197  &  wire34399 ) | ( wire193  &  n_n4441  &  wire34399 ) ;
 assign wire2957 = ( (~ n_n5514)  &  wire1006  &  wire34401 ) | ( (~ n_n5514)  &  wire33609  &  wire34401 ) ;
 assign wire2958 = ( pi20  &  nv8372  &  wire153 ) | ( (~ pi20)  &  nv8372  &  wire153 ) ;
 assign wire2959 = ( nv10167  &  wire3195 ) | ( nv10167  &  wire3196 ) ;
 assign wire2960 = ( (~ pi17)  &  wire179  &  nv8372 ) ;
 assign wire2961 = ( wire197  &  wire203 ) | ( wire193  &  n_n4501  &  wire203 ) ;
 assign wire2962 = ( pi20  &  wire197  &  wire153 ) | ( pi20  &  wire153  &  wire3231 ) ;
 assign wire2963 = ( (~ pi20)  &  wire197  &  wire153 ) | ( (~ pi20)  &  wire153  &  wire3328 ) ;
 assign wire2964 = ( wire197  &  wire199 ) | ( wire193  &  n_n4441  &  wire199 ) ;
 assign wire2967 = ( wire197  &  nv10167 ) | ( wire193  &  n_n4509  &  nv10167 ) ;
 assign wire2972 = ( (~ pi16)  &  (~ pi24)  &  wire641 ) ;
 assign wire2980 = ( wire3308  &  wire34481 ) | ( (~ n_n5574)  &  wire33603  &  wire34481 ) ;
 assign wire2981 = ( pi20  &  nv8372  &  wire153 ) | ( (~ pi20)  &  nv8372  &  wire153 ) ;
 assign wire2983 = ( wire193  &  wire3322 ) | ( wire193  &  n_n4509  &  wire33475 ) ;
 assign wire2984 = ( wire197  &  nv10167 ) | ( nv10167  &  wire3320 ) ;
 assign wire2986 = ( wire3251  &  wire34489 ) | ( n_n4481  &  wire33350  &  wire34489 ) ;
 assign wire2987 = ( wire3280  &  wire34490 ) | ( n_n4489  &  wire33307  &  wire34490 ) ;
 assign wire2990 = ( pi17  &  (~ pi16)  &  wire178  &  nv8372 ) ;
 assign wire2994 = ( wire158  &  wire180  &  wire197 ) | ( wire158  &  wire180  &  wire3249 ) ;
 assign wire2995 = ( wire197  &  wire194 ) | ( wire193  &  n_n4611  &  wire194 ) ;
 assign wire3000 = ( wire193  &  wire3318 ) | ( wire193  &  n_n4501  &  wire33595 ) ;
 assign wire3001 = ( wire197  &  nv10167 ) | ( nv10167  &  wire3316 ) ;
 assign wire3005 = ( pi16  &  pi24  &  wire3023 ) | ( pi16  &  pi24  &  wire34454 ) ;
 assign wire3006 = ( pi16  &  (~ pi24)  &  wire501 ) ;
 assign wire3008 = ( (~ pi24)  &  wire3019 ) | ( (~ pi24)  &  wire34457 ) ;
 assign wire3011 = ( wire3189  &  wire34458 ) | ( n_n4412  &  wire33395  &  wire34458 ) ;
 assign wire3015 = ( pi17  &  pi16  &  wire178  &  nv8372 ) ;
 assign wire3019 = ( wire180  &  wire197  &  wire154 ) | ( wire180  &  wire154  &  wire3187 ) ;
 assign wire3020 = ( wire197  &  wire183 ) | ( wire193  &  n_n4543  &  wire183 ) ;
 assign wire3023 = ( wire197  &  wire34448 ) | ( wire3391  &  wire34448 ) ;
 assign wire3024 = ( wire3393  &  wire34449 ) | ( n_n4441  &  wire33555  &  wire34449 ) ;
 assign wire3027 = ( (~ pi17)  &  wire179  &  nv8372 ) ;
 assign wire3030 = ( wire193  &  wire3341 ) | ( n_n4433  &  wire193  &  wire33515 ) ;
 assign wire3031 = ( wire197  &  nv10167 ) | ( nv10167  &  wire3339 ) ;
 assign wire3034 = ( wire197  &  nv10167 ) | ( n_n4433  &  wire193  &  nv10167 ) ;
 assign wire3036 = ( wire3341  &  wire33738 ) | ( n_n4433  &  wire33515  &  wire33738 ) ;
 assign wire3040 = ( wire33682  &  wire33745 ) | ( n_n4481  &  wire329  &  wire33745 ) ;
 assign wire3041 = ( wire1291  &  wire33746 ) | ( wire189  &  n_n5481  &  wire33746 ) ;
 assign wire3042 = ( (~ pi16)  &  pi15  &  wire3111 ) | ( (~ pi16)  &  pi15  &  wire3112 ) ;
 assign wire3045 = ( pi15  &  wire754 ) | ( pi15  &  wire33750 ) ;
 assign wire3046 = ( pi16  &  (~ pi15)  &  wire739 ) | ( pi16  &  (~ pi15)  &  wire3058 ) ;
 assign wire3047 = ( (~ pi15)  &  wire1206 ) ;
 assign wire3048 = ( wire1031  &  wire1291 ) | ( wire189  &  wire1031  &  n_n5481 ) ;
 assign wire3049 = ( (~ pi15)  &  wire3075 ) | ( (~ pi15)  &  wire3076 ) | ( (~ pi15)  &  wire33756 ) ;
 assign wire3050 = ( wire226  &  wire740 ) | ( wire226  &  n_n4441  &  wire475 ) ;
 assign wire3051 = ( pi15  &  wire918 ) | ( pi15  &  wire476  &  n_n4834 ) ;
 assign wire3056 = ( (~ pi21)  &  ni30  &  wire616 ) | ( pi21  &  (~ pi22)  &  ni30  &  wire616 ) ;
 assign wire3057 = ( (~ pi17)  &  pi25  &  ni30  &  wire179 ) ;
 assign wire3058 = ( wire475  &  wire3393 ) | ( n_n4441  &  wire475  &  wire33555 ) ;
 assign wire3060 = ( wire247  &  wire3215 ) | ( (~ n_n5514)  &  wire247  &  wire33608 ) ;
 assign wire3064 = ( wire180  &  wire3189 ) | ( wire180  &  n_n4412  &  wire33395 ) ;
 assign wire3066 = ( (~ pi19)  &  ni30 ) ;
 assign wire3069 = ( pi17  &  pi25  &  pi16  &  ni30 ) ;
 assign wire3074 = ( (~ pi16)  &  wire433 ) | ( (~ pi16)  &  n_n5481  &  wire448 ) ;
 assign wire3075 = ( wire899  &  wire3098 ) | ( wire899  &  wire3099 ) | ( wire899  &  wire33702 ) ;
 assign wire3076 = ( (~ pi16)  &  wire3088 ) | ( (~ pi16)  &  wire3090 ) | ( (~ pi16)  &  wire3091 ) ;
 assign wire3083 = ( (~ pi21)  &  ni30  &  wire340 ) | ( pi21  &  (~ pi22)  &  ni30  &  wire340 ) ;
 assign wire3084 = ( pi20  &  pi25  &  ni30  &  wire153 ) ;
 assign wire3085 = ( (~ pi20)  &  pi25  &  ni30  &  wire153 ) ;
 assign wire3086 = ( (~ pi21)  &  (~ pi16)  &  ni30 ) | ( (~ pi22)  &  (~ pi16)  &  ni30 ) ;
 assign wire3088 = ( wire437  &  wire3318 ) | ( n_n4501  &  wire437  &  wire33595 ) ;
 assign wire3090 = ( (~ pi17)  &  pi25  &  ni30  &  wire182 ) ;
 assign wire3091 = ( (~ pi21)  &  ni30  &  wire381 ) | ( pi21  &  (~ pi22)  &  ni30  &  wire381 ) ;
 assign wire3092 = ( wire387  &  wire3322 ) | ( n_n4509  &  wire387  &  wire33475 ) ;
 assign wire3093 = ( (~ pi20)  &  wire351 ) ;
 assign wire3096 = ( wire247  &  wire3308 ) | ( (~ n_n5574)  &  wire247  &  wire33603 ) ;
 assign wire3097 = ( wire219  &  wire3327 ) | ( (~ n_n5580)  &  wire219  &  wire33598 ) ;
 assign wire3098 = ( wire460  &  wire3280 ) | ( n_n4489  &  wire460  &  wire33307 ) ;
 assign wire3099 = ( wire329  &  wire3251 ) | ( n_n4481  &  wire329  &  wire33350 ) ;
 assign wire3104 = ( (~ n_n5514)  &  wire247  &  wire1006 ) | ( (~ n_n5514)  &  wire247  &  wire33609 ) ;
 assign wire3109 = ( wire178  &  wire721  &  wire33433 ) | ( wire178  &  wire721  &  wire33434 ) ;
 assign wire3110 = ( (~ pi19)  &  ni30 ) ;
 assign wire3111 = ( (~ n_n5574)  &  wire247  &  wire1006 ) | ( (~ n_n5574)  &  wire247  &  wire33604 ) ;
 assign wire3112 = ( (~ n_n5580)  &  wire1006  &  wire219 ) | ( (~ n_n5580)  &  wire219  &  wire33599 ) ;
 assign wire3114 = ( pi17  &  wire180  &  n_n4481 ) ;
 assign wire3116 = ( pi17  &  ni30 ) ;
 assign wire3117 = ( (~ wire150)  &  wire699  &  wire3157 ) | ( (~ wire150)  &  wire699  &  wire3158 ) ;
 assign wire3118 = ( (~ wire150)  &  wire377  &  wire3139 ) | ( (~ wire150)  &  wire377  &  wire3140 ) ;
 assign wire3119 = ( wire173  &  wire788 ) | ( wire1063  &  wire788 ) ;
 assign wire3120 = ( (~ pi21)  &  nv7791  &  wire699 ) | ( pi21  &  (~ pi22)  &  nv7791  &  wire699 ) ;
 assign wire3121 = ( (~ pi21)  &  nv7445  &  wire377 ) | ( pi21  &  (~ pi22)  &  nv7445  &  wire377 ) ;
 assign wire3122 = ( (~ pi21)  &  nv7647  &  wire268 ) | ( pi21  &  (~ pi22)  &  nv7647  &  wire268 ) ;
 assign wire3125 = ( pi27  &  nv7447 ) | ( pi27  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3126 = ( (~ pi27)  &  ni30 ) | ( (~ pi27)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3139 = ( (~ wire156)  &  nv7447 ) | ( (~ wire156)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3140 = ( ni30  &  wire156 ) | ( wire156  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3141 = ( nv8372  &  wire33941 ) | ( (~ wire157)  &  (~ nv6462)  &  wire33941 ) ;
 assign wire3144 = ( pi21  &  wire3147 ) | ( pi21  &  nv8372  &  wire33940 ) ;
 assign wire3147 = ( (~ pi22)  &  pi23  &  ni30 ) | ( (~ pi22)  &  pi24  &  ni30 ) ;
 assign wire3149 = ( (~ pi21)  &  pi23  &  ni30 ) | ( (~ pi21)  &  pi24  &  ni30 ) ;
 assign wire3150 = ( nv8608  &  (~ wire155) ) | ( (~ wire155)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3151 = ( wire155  &  nv8372 ) | ( wire155  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3153 = ( nv8372  &  wire1044 ) | ( (~ wire157)  &  (~ nv6462)  &  wire1044 ) ;
 assign wire3156 = ( (~ pi21)  &  (~ pi24)  &  ni30 ) | ( pi21  &  (~ pi22)  &  (~ pi24)  &  ni30 ) ;
 assign wire3157 = ( (~ wire155)  &  nv7447 ) | ( (~ wire155)  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3158 = ( ni30  &  wire155 ) | ( wire155  &  (~ wire157)  &  (~ nv6462) ) ;
 assign wire3159 = ( wire197  &  wire33866 ) | ( wire3339  &  wire33866 ) ;
 assign wire3160 = ( wire197  &  wire33868 ) | ( wire3391  &  wire33868 ) ;
 assign wire3161 = ( wire197  &  wire33870 ) | ( wire193  &  n_n4441  &  wire33870 ) ;
 assign wire3162 = ( wire197  &  wire33872 ) | ( n_n4433  &  wire193  &  wire33872 ) ;
 assign wire3165 = ( wire197  &  wire33875 ) | ( wire193  &  n_n4509  &  wire33875 ) ;
 assign wire3166 = ( wire197  &  wire33876 ) | ( wire193  &  n_n4501  &  wire33876 ) ;
 assign wire3167 = ( (~ wire175)  &  wire226  &  wire3195 ) | ( (~ wire175)  &  wire226  &  wire3196 ) ;
 assign wire3168 = ( pi16  &  (~ pi15)  &  (~ wire175)  &  wire385 ) ;
 assign wire3169 = ( (~ wire175)  &  wire173  &  wire208 ) ;
 assign wire3170 = ( wire3221  &  wire33880 ) | ( wire3222  &  wire33880 ) | ( wire33831  &  wire33880 ) ;
 assign wire3171 = ( wire197  &  wire33881 ) | ( wire3231  &  wire33881 ) ;
 assign wire3173 = ( wire197  &  wire33883 ) | ( wire3328  &  wire33883 ) ;
 assign wire3174 = ( (~ wire175)  &  wire403  &  wire3439 ) | ( (~ wire175)  &  wire403  &  wire33796 ) ;
 assign wire3175 = ( (~ pi17)  &  (~ pi16)  &  wire173  &  wire369 ) ;
 assign wire3176 = ( wire370  &  wire3179 ) | ( wire370  &  wire33818 ) ;
 assign wire3177 = ( wire370  &  wire3240 ) | ( wire370  &  wire3243 ) | ( wire370  &  wire33887 ) ;
 assign wire3179 = ( wire180  &  wire197  &  wire154 ) | ( wire180  &  wire154  &  wire3187 ) ;
 assign wire3182 = ( wire197  &  wire183 ) | ( wire193  &  n_n4543  &  wire183 ) ;
 assign wire3185 = ( wire721  &  wire417  &  (~ wire1198)  &  (~ wire3466) ) ;
 assign wire3186 = ( (~ n_n5621)  &  wire721  &  wire33433 ) | ( (~ n_n5621)  &  wire721  &  wire33434 ) ;
 assign wire3187 = ( wire193  &  wire3189 ) | ( n_n4412  &  wire193  &  wire33395 ) ;
 assign wire3189 = ( wire33386  &  wire33392 ) | ( wire33387  &  wire33392 ) | ( wire33391  &  wire33392 ) ;
 assign wire3193 = ( (~ ni37)  &  ni36  &  (~ wire157)  &  (~ nv669) ) ;
 assign wire3195 = ( pi20  &  wire197  &  wire153 ) | ( pi20  &  wire153  &  wire3197 ) ;
 assign wire3196 = ( (~ pi20)  &  wire197  &  wire153 ) | ( (~ pi20)  &  wire153  &  wire3199 ) ;
 assign wire3197 = ( wire193  &  (~ n_n5514)  &  wire1006 ) | ( wire193  &  (~ n_n5514)  &  wire33609 ) ;
 assign wire3199 = ( wire193  &  wire1006  &  (~ n_n5520) ) | ( wire193  &  (~ n_n5520)  &  wire33612 ) ;
 assign wire3205 = ( (~ nv669)  &  wire1074  &  (~ n_n5520)  &  (~ wire6766) ) ;
 assign wire3206 = ( wire477  &  wire1006  &  (~ n_n5520) ) | ( wire477  &  (~ n_n5520)  &  wire33612 ) ;
 assign wire3214 = ( (~ nv669)  &  (~ n_n5514)  &  wire1074  &  (~ wire6727) ) ;
 assign wire3215 = ( (~ n_n5514)  &  wire477  &  wire1006 ) | ( (~ n_n5514)  &  wire477  &  wire33609 ) ;
 assign wire3221 = ( wire197  &  wire460 ) | ( n_n4489  &  wire193  &  wire460 ) ;
 assign wire3222 = ( wire197  &  wire329 ) | ( wire193  &  n_n4481  &  wire329 ) ;
 assign wire3223 = ( wire272  &  wire197 ) | ( wire272  &  wire193  &  n_n4473 ) ;
 assign wire3231 = ( wire193  &  (~ n_n5574)  &  wire1006 ) | ( wire193  &  (~ n_n5574)  &  wire33604 ) ;
 assign wire3233 = ( (~ ni33)  &  n_n4404 ) | ( (~ ni29)  &  n_n4404 ) | ( n_n4404  &  (~ nv6462) ) ;
 assign wire3240 = ( wire197  &  wire484 ) | ( wire484  &  wire3316 ) ;
 assign wire3243 = ( (~ pi16)  &  wire3246 ) | ( (~ pi16)  &  wire33802 ) ;
 assign wire3246 = ( pi17  &  wire180  &  wire197 ) | ( pi17  &  wire180  &  wire3249 ) ;
 assign wire3247 = ( wire272  &  wire197 ) | ( wire272  &  wire193  &  n_n4611 ) ;
 assign wire3249 = ( wire193  &  wire3251 ) | ( wire193  &  n_n4481  &  wire33350 ) ;
 assign wire3251 = ( wire33341  &  wire33347 ) | ( wire33342  &  wire33347 ) | ( wire33346  &  wire33347 ) ;
 assign wire3257 = ( (~ ni37)  &  (~ wire826)  &  (~ wire3491)  &  (~ wire33310) ) ;
 assign wire3260 = ( (~ ni37)  &  (~ nv6486)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire3266 = ( (~ nv6486)  &  (~ wire826)  &  wire33334 ) ;
 assign wire3274 = ( wire426  &  (~ wire157)  &  (~ wire205)  &  (~ nv669) ) ;
 assign wire3276 = ( wire426  &  (~ wire157)  &  (~ nv669)  &  (~ n_n2328) ) ;
 assign wire3277 = ( (~ ni47)  &  (~ ni45)  &  (~ ni38)  &  (~ wire157) ) ;
 assign wire3278 = ( wire193  &  wire3280 ) | ( n_n4489  &  wire193  &  wire33307 ) ;
 assign wire3280 = ( wire33298  &  wire33304 ) | ( wire33299  &  wire33304 ) | ( wire33303  &  wire33304 ) ;
 assign wire3292 = ( (~ ni37)  &  (~ wire827)  &  (~ wire1047)  &  (~ nv6472) ) ;
 assign wire3295 = ( (~ wire827)  &  (~ nv6472)  &  wire33291 ) ;
 assign wire3297 = ( (~ wire426)  &  wire253 ) | ( wire253  &  nv669 ) | ( wire253  &  wire6766 ) ;
 assign wire3301 = ( (~ wire426)  &  wire691 ) | ( nv669  &  wire691 ) | ( wire691  &  wire6766 ) ;
 assign wire3303 = ( nv669  &  wire685 ) | ( (~ ni42)  &  ni41  &  wire685 ) ;
 assign wire3307 = ( wire1074  &  (~ n_n5574)  &  (~ nv6486) ) ;
 assign wire3308 = ( wire477  &  (~ n_n5574)  &  wire1006 ) | ( wire477  &  (~ n_n5574)  &  wire33604 ) ;
 assign wire3314 = ( ni38  &  ni37  &  (~ ni36) ) ;
 assign wire3316 = ( wire193  &  wire3318 ) | ( wire193  &  n_n4501  &  wire33595 ) ;
 assign wire3318 = ( wire33586  &  wire33592 ) | ( wire33587  &  wire33592 ) | ( wire33591  &  wire33592 ) ;
 assign wire3320 = ( wire193  &  wire3322 ) | ( wire193  &  n_n4509  &  wire33475 ) ;
 assign wire3322 = ( wire33466  &  wire33472 ) | ( wire33467  &  wire33472 ) | ( wire33471  &  wire33472 ) ;
 assign wire3326 = ( (~ n_n5580)  &  wire33598 ) ;
 assign wire3327 = ( wire477  &  (~ n_n5580)  &  wire1006 ) | ( wire477  &  (~ n_n5580)  &  wire33599 ) ;
 assign wire3328 = ( wire193  &  (~ n_n5580)  &  wire1006 ) | ( wire193  &  (~ n_n5580)  &  wire33599 ) ;
 assign wire3337 = ( ni38  &  ni37  &  (~ ni36) ) ;
 assign wire3339 = ( wire193  &  wire3341 ) | ( n_n4433  &  wire193  &  wire33515 ) ;
 assign wire3341 = ( wire33506  &  wire33512 ) | ( wire33507  &  wire33512 ) | ( wire33511  &  wire33512 ) ;
 assign wire3349 = ( (~ ni37)  &  (~ wire826)  &  (~ wire3491)  &  (~ wire33310) ) ;
 assign wire3355 = ( (~ ni37)  &  (~ nv6486)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire3358 = ( (~ nv6486)  &  (~ wire826)  &  wire33579 ) ;
 assign wire3375 = ( (~ ni37)  &  (~ wire827)  &  (~ wire1081)  &  (~ nv6472) ) ;
 assign wire3381 = ( (~ wire827)  &  (~ nv6472)  &  wire33459 ) ;
 assign wire3383 = ( (~ wire426)  &  wire254 ) | ( wire254  &  nv669 ) | ( wire254  &  wire6766 ) ;
 assign wire3387 = ( (~ wire426)  &  wire685 ) | ( nv669  &  wire685 ) | ( wire685  &  wire6766 ) ;
 assign wire3389 = ( nv669  &  wire691 ) | ( (~ ni42)  &  ni41  &  wire691 ) ;
 assign wire3391 = ( wire193  &  wire3393 ) | ( wire193  &  n_n4441  &  wire33555 ) ;
 assign wire3393 = ( wire33546  &  wire33552 ) | ( wire33547  &  wire33552 ) | ( wire33551  &  wire33552 ) ;
 assign wire3399 = ( (~ ni37)  &  (~ wire827)  &  (~ wire3462)  &  (~ wire33267) ) ;
 assign wire3402 = ( (~ wire827)  &  (~ wire1081)  &  wire33527 ) ;
 assign wire3405 = ( (~ wire827)  &  (~ wire1047)  &  wire33533 ) ;
 assign wire3406 = ( (~ wire827)  &  (~ wire468)  &  (~ wire3410)  &  wire33535 ) ;
 assign wire3407 = ( (~ wire827)  &  wire1200  &  wire33537 ) | ( (~ wire827)  &  wire3412  &  wire33537 ) ;
 assign wire3410 = ( ni40  &  ni38  &  nv669 ) | ( ni40  &  ni38  &  wire6766 ) ;
 assign wire3412 = ( nv669  &  wire685 ) | ( wire685  &  wire6766 ) ;
 assign wire3420 = ( (~ ni37)  &  (~ wire826)  &  (~ wire3491)  &  (~ wire33310) ) ;
 assign wire3426 = ( (~ ni37)  &  (~ nv6589)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire3429 = ( (~ nv6589)  &  (~ wire826)  &  wire33499 ) ;
 assign wire3431 = ( wire254  &  wire6727 ) | ( ni41  &  wire254  &  nv669 ) | ( (~ ni41)  &  wire254  &  nv669 ) ;
 assign wire3435 = ( wire685  &  wire6727 ) | ( ni41  &  nv669  &  wire685 ) | ( (~ ni41)  &  nv669  &  wire685 ) ;
 assign wire3439 = ( wire180  &  wire197 ) | ( wire180  &  n_n4412  &  wire193 ) ;
 assign wire3444 = ( wire721  &  wire193  &  wire33433 ) | ( wire721  &  wire193  &  wire33434 ) ;
 assign wire3448 = ( (~ wire827)  &  (~ wire464)  &  (~ wire3464)  &  wire33398 ) ;
 assign wire3449 = ( (~ wire827)  &  wire1198  &  wire33400 ) | ( (~ wire827)  &  wire3466  &  wire33400 ) ;
 assign wire3450 = ( (~ ni37)  &  (~ wire827)  &  (~ wire3462)  &  (~ wire33267) ) ;
 assign wire3453 = ( (~ wire827)  &  (~ wire1081)  &  wire33407 ) ;
 assign wire3456 = ( (~ wire827)  &  (~ wire1047)  &  wire33413 ) ;
 assign wire3457 = ( (~ wire827)  &  (~ wire464)  &  (~ wire3464)  &  wire33415 ) ;
 assign wire3458 = ( (~ wire827)  &  wire1198  &  wire33417 ) | ( (~ wire827)  &  wire3466  &  wire33417 ) ;
 assign wire3462 = ( ni39  &  ni47  &  (~ ni36) ) | ( ni39  &  ni45  &  (~ ni36) ) ;
 assign wire3464 = ( (~ ni40)  &  ni38  &  nv669 ) | ( (~ ni40)  &  ni38  &  wire6766 ) ;
 assign wire3466 = ( nv669  &  wire691 ) | ( wire691  &  wire6766 ) ;
 assign wire3474 = ( ni47  &  (~ ni38)  &  ni37 ) | ( ni45  &  (~ ni38)  &  ni37 ) ;
 assign wire3479 = ( (~ ni37)  &  (~ wire826)  &  (~ wire3491)  &  (~ wire33310) ) ;
 assign wire3482 = ( (~ ni37)  &  (~ nv6589)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire3488 = ( (~ nv6589)  &  (~ wire826)  &  wire33379 ) ;
 assign wire3491 = ( (~ ni39)  &  ni47  &  (~ ni36) ) | ( (~ ni39)  &  ni45  &  (~ ni36) ) ;
 assign wire3493 = ( wire253  &  wire6727 ) | ( ni41  &  wire253  &  nv669 ) | ( (~ ni41)  &  wire253  &  nv669 ) ;
 assign wire3497 = ( wire691  &  wire6727 ) | ( ni41  &  nv669  &  wire691 ) | ( (~ ni41)  &  nv669  &  wire691 ) ;
 assign wire3506 = ( ni2  &  ni8 ) | ( ni3  &  ni8 ) ;
 assign wire3512 = ( n_n13895  &  wire1165  &  wire5961 ) | ( n_n13895  &  wire1165  &  wire5962 ) ;
 assign wire3514 = ( ni2  &  ni7 ) | ( ni3  &  ni7 ) ;
 assign wire3515 = ( wire31875  &  wire31918 ) | ( wire31876  &  wire31918 ) | ( wire31916  &  wire31918 ) ;
 assign wire3516 = ( wire3889  &  wire31997 ) | ( wire31995  &  wire31997 ) ;
 assign wire3517 = ( wire32053  &  wire32055 ) | ( (~ pi15)  &  n_n9255  &  wire32055 ) ;
 assign wire3520 = ( wire4419  &  wire32182 ) | ( wire32181  &  wire32182 ) ;
 assign wire3521 = ( wire33240  &  wire33241 ) | ( (~ ni7)  &  n_n8112  &  wire33241 ) ;
 assign wire3522 = ( ni2  &  ni32 ) | ( ni3  &  ni32 ) ;
 assign wire3528 = ( wire818  &  wire453  &  wire1328  &  wire32203 ) ;
 assign wire3529 = ( wire3644  &  wire32216 ) | ( wire3647  &  wire32216 ) | ( wire32212  &  wire32216 ) ;
 assign wire3533 = ( wire4295  &  wire32340 ) | ( wire32338  &  wire32340 ) ;
 assign wire3534 = ( (~ pi24)  &  wire791  &  wire359  &  wire1328 ) ;
 assign wire3537 = ( wire3561  &  wire32485 ) | ( wire3562  &  wire32485 ) | ( wire32483  &  wire32485 ) ;
 assign wire3540 = ( wire4253  &  wire32580 ) | ( wire4254  &  wire32580 ) | ( wire32578  &  wire32580 ) ;
 assign wire3543 = ( wire306  &  wire32357 ) | ( wire233  &  n_n7913  &  wire32357 ) ;
 assign wire3544 = ( wire305  &  wire32360 ) | ( wire233  &  n_n7913  &  wire32360 ) ;
 assign wire3545 = ( wire305  &  wire32363 ) | ( wire233  &  n_n7905  &  wire32363 ) ;
 assign wire3546 = ( (~ wire150)  &  wire4433  &  wire32365 ) | ( (~ wire150)  &  wire4434  &  wire32365 ) ;
 assign wire3547 = ( wire306  &  wire32367 ) | ( wire233  &  n_n7905  &  wire32367 ) ;
 assign wire3548 = ( wire3584  &  wire32369 ) | ( (~ pi20)  &  n_n5908  &  wire32369 ) ;
 assign wire3549 = ( wire4276  &  wire32371 ) | ( wire32228  &  wire32371 ) ;
 assign wire3551 = ( wire3644  &  wire32375 ) | ( wire3647  &  wire32375 ) | ( wire32212  &  wire32375 ) ;
 assign wire3552 = ( (~ pi23)  &  ni11  &  wire352  &  (~ wire574) ) ;
 assign wire3553 = ( (~ wire165)  &  wire4295  &  wire32378 ) | ( (~ wire165)  &  wire32338  &  wire32378 ) ;
 assign wire3554 = ( wire198  &  wire334  &  wire32380 ) ;
 assign wire3555 = ( wire4264  &  wire32408 ) | ( wire4266  &  wire32408 ) | ( wire32406  &  wire32408 ) ;
 assign wire3556 = ( wire4281  &  wire32409 ) | ( wire263  &  wire453  &  wire32409 ) ;
 assign wire3557 = ( wire4282  &  wire32410 ) | ( wire4283  &  wire32410 ) | ( wire4284  &  wire32410 ) ;
 assign wire3558 = ( wire32256  &  wire32411 ) | ( n_n7885  &  wire32251  &  wire32411 ) ;
 assign wire3559 = ( pi15  &  (~ wire289)  &  wire158  &  wire334 ) ;
 assign wire3561 = ( wire708  &  wire3581 ) | ( wire708  &  wire32427 ) | ( wire708  &  wire32428 ) ;
 assign wire3562 = ( wire708  &  wire3594 ) | ( wire708  &  wire32446 ) | ( wire708  &  wire32447 ) ;
 assign wire3563 = ( pi15  &  (~ wire289)  &  wire32463 ) | ( pi15  &  (~ wire289)  &  wire32464 ) ;
 assign wire3564 = ( wire555  &  nv6289 ) ;
 assign wire3565 = ( wire306  &  wire32450 ) | ( wire233  &  n_n7845  &  wire32450 ) ;
 assign wire3566 = ( wire305  &  wire32452 ) | ( wire233  &  n_n7845  &  wire32452 ) ;
 assign wire3567 = ( wire306  &  wire32453 ) | ( wire233  &  n_n7837  &  wire32453 ) ;
 assign wire3568 = ( wire3584  &  wire32454 ) | ( (~ pi20)  &  n_n5908  &  wire32454 ) ;
 assign wire3569 = ( wire4501  &  wire32455 ) | ( wire4504  &  wire32455 ) | ( wire32066  &  wire32455 ) ;
 assign wire3571 = ( pi16  &  wire198  &  wire334 ) ;
 assign wire3572 = ( pi23  &  (~ pi24)  &  wire4317 ) | ( pi23  &  (~ pi24)  &  wire32264 ) ;
 assign wire3573 = ( wire160  &  wire4322 ) | ( wire160  &  wire4323 ) | ( wire160  &  wire4324 ) ;
 assign wire3576 = ( wire305  &  wire32419 ) | ( wire4544  &  wire32419 ) ;
 assign wire3577 = ( wire3584  &  wire32420 ) | ( (~ pi20)  &  n_n5908  &  wire32420 ) ;
 assign wire3578 = ( wire4349  &  wire32421 ) | ( wire32277  &  wire32421 ) ;
 assign wire3580 = ( pi16  &  wire198  &  wire334 ) ;
 assign wire3581 = ( (~ pi23)  &  wire4341 ) | ( pi24  &  wire4341 ) | ( (~ pi23)  &  wire32291 ) | ( pi24  &  wire32291 ) ;
 assign wire3582 = ( (~ wire160)  &  wire4343 ) | ( (~ wire160)  &  wire4344 ) | ( (~ wire160)  &  wire32297 ) ;
 assign wire3584 = ( pi21  &  (~ pi20)  &  wire3601 ) | ( pi21  &  (~ pi20)  &  wire3602 ) ;
 assign wire3587 = ( wire306  &  wire32433 ) | ( wire4387  &  wire32433 ) ;
 assign wire3588 = ( wire211  &  wire3601  &  wire32434 ) | ( wire211  &  wire3602  &  wire32434 ) ;
 assign wire3589 = ( n_n5908  &  wire32437 ) ;
 assign wire3590 = ( wire4378  &  wire32438 ) | ( wire32285  &  wire32438 ) ;
 assign wire3593 = ( (~ wire160)  &  wire4367 ) | ( (~ wire160)  &  wire4368 ) | ( (~ wire160)  &  wire32304 ) ;
 assign wire3594 = ( (~ pi23)  &  wire4374 ) | ( pi24  &  wire4374 ) | ( (~ pi23)  &  wire32306 ) | ( pi24  &  wire32306 ) ;
 assign wire3596 = ( n_n6710  &  wire32413 ) | ( n_n6711  &  wire32413 ) | ( wire4973  &  wire32413 ) ;
 assign wire3601 = ( (~ pi22)  &  (~ wire160)  &  n_n6367 ) | ( (~ pi22)  &  (~ wire160)  &  n_n6711 ) ;
 assign wire3602 = ( (~ pi22)  &  (~ pi23)  &  nv3908 ) | ( (~ pi22)  &  pi24  &  nv3908 ) ;
 assign wire3605 = ( wire305  &  wire32223 ) | ( wire233  &  n_n7905  &  wire32223 ) ;
 assign wire3606 = ( wire305  &  wire32225 ) | ( wire233  &  n_n7845  &  wire32225 ) ;
 assign wire3607 = ( wire4273  &  wire32230 ) | ( wire4276  &  wire32230 ) | ( wire32228  &  wire32230 ) ;
 assign wire3608 = ( wire4309  &  wire32235 ) | ( wire4312  &  wire32235 ) | ( wire32233  &  wire32235 ) ;
 assign wire3609 = ( wire306  &  wire32237 ) | ( wire233  &  n_n7837  &  wire32237 ) ;
 assign wire3610 = ( wire306  &  wire32239 ) | ( wire233  &  n_n7905  &  wire32239 ) ;
 assign wire3611 = ( wire449  &  wire32241 ) | ( wire4491  &  wire32241 ) ;
 assign wire3612 = ( wire4501  &  wire32243 ) | ( wire4504  &  wire32243 ) | ( wire32066  &  wire32243 ) ;
 assign wire3615 = ( wire4282  &  wire32249 ) | ( wire4283  &  wire32249 ) | ( wire4284  &  wire32249 ) ;
 assign wire3617 = ( pi15  &  pi24  &  wire4317 ) | ( pi15  &  pi24  &  wire32264 ) ;
 assign wire3618 = ( wire4322  &  wire32267 ) | ( wire4323  &  wire32267 ) | ( wire4324  &  wire32267 ) ;
 assign wire3623 = ( pi16  &  pi24  &  wire4349 ) | ( pi16  &  pi24  &  wire32277 ) ;
 assign wire3625 = ( (~ pi16)  &  pi24  &  wire4378 ) | ( (~ pi16)  &  pi24  &  wire32285 ) ;
 assign wire3627 = ( wire306  &  wire32288 ) | ( wire4387  &  wire32288 ) ;
 assign wire3628 = ( wire305  &  wire32289 ) | ( wire4564  &  wire32289 ) ;
 assign wire3629 = ( wire305  &  wire32290 ) | ( wire4544  &  wire32290 ) ;
 assign wire3630 = ( (~ pi24)  &  wire4341 ) | ( (~ pi24)  &  wire32291 ) ;
 assign wire3631 = ( pi24  &  wire4343 ) | ( pi24  &  wire4344 ) | ( pi24  &  wire32297 ) ;
 assign wire3632 = ( pi24  &  wire4367 ) | ( pi24  &  wire4368 ) | ( pi24  &  wire32304 ) ;
 assign wire3639 = ( (~ pi21)  &  ni32  &  (~ ni30) ) ;
 assign wire3641 = ( n_n6367  &  wire32206 ) | ( n_n6711  &  wire32206 ) ;
 assign wire3642 = ( n_n6710  &  wire32207 ) | ( n_n6711  &  wire32207 ) | ( wire4973  &  wire32207 ) ;
 assign wire3644 = ( pi26  &  (~ pi24)  &  wire4269 ) | ( pi26  &  (~ pi24)  &  wire32189 ) ;
 assign wire3645 = ( (~ pi21)  &  (~ pi26)  &  (~ pi24)  &  wire424 ) ;
 assign wire3647 = ( wire1044  &  wire4458 ) | ( wire1044  &  wire4459 ) ;
 assign wire3650 = ( wire31592  &  wire32586 ) | ( wire31593  &  wire32586 ) | ( wire31594  &  wire32586 ) ;
 assign wire3651 = ( wire4090  &  wire32591 ) | ( wire32587  &  wire32591 ) ;
 assign wire3652 = ( wire31252  &  wire32595 ) | ( wire31253  &  wire32595 ) | ( wire31254  &  wire32595 ) ;
 assign wire3653 = ( n_n6710  &  wire32599 ) | ( wire4807  &  wire32599 ) | ( wire4808  &  wire32599 ) ;
 assign wire3655 = ( wire4079  &  wire32605 ) | ( wire182  &  wire280  &  wire32605 ) ;
 assign wire3658 = ( n_n6710  &  wire32614 ) | ( wire4813  &  wire32614 ) | ( wire4814  &  wire32614 ) ;
 assign wire3660 = ( wire4078  &  wire32619 ) | ( wire32617  &  wire32619 ) ;
 assign wire3661 = ( wire4083  &  wire32621 ) | ( wire180  &  wire280  &  wire32621 ) ;
 assign wire3662 = ( wire393  &  wire4613  &  wire32622 ) | ( wire393  &  wire31347  &  wire32622 ) ;
 assign wire3663 = ( wire32651  &  wire32681 ) | ( wire32652  &  wire32681 ) | ( wire32680  &  wire32681 ) ;
 assign wire3664 = ( wire3706  &  wire32682 ) | ( wire194  &  wire280  &  wire32682 ) ;
 assign wire3665 = ( wire4064  &  wire32710 ) | ( wire4065  &  wire32710 ) | ( wire32709  &  wire32710 ) ;
 assign wire3666 = ( wire32053  &  wire32711 ) | ( (~ pi15)  &  n_n9255  &  wire32711 ) ;
 assign wire3667 = ( wire1316  &  wire32919 ) | ( (~ ni11)  &  n_n8104  &  wire1316 ) ;
 assign wire3668 = ( ni9  &  (~ ni8)  &  nv5843 ) ;
 assign wire3670 = ( (~ wire793)  &  wire3780 ) | ( (~ wire793)  &  wire33201 ) | ( (~ wire793)  &  wire33202 ) ;
 assign wire3676 = ( wire3704  &  wire32664 ) | ( wire179  &  wire280  &  wire32664 ) ;
 assign wire3679 = ( wire4090  &  wire32667 ) | ( wire32587  &  wire32667 ) ;
 assign wire3680 = ( pi16  &  wire219  &  wire4779 ) | ( pi16  &  wire219  &  wire31895 ) ;
 assign wire3681 = ( pi16  &  wire3703 ) | ( pi16  &  wire32639 ) ;
 assign wire3682 = ( wire154  &  wire4083 ) | ( wire180  &  wire154  &  wire280 ) ;
 assign wire3687 = ( wire4090  &  wire32627 ) | ( wire32587  &  wire32627 ) ;
 assign wire3690 = ( (~ pi17)  &  (~ pi16)  &  wire358  &  n_n7913 ) ;
 assign wire3691 = ( wire3704  &  wire32633 ) | ( wire179  &  wire280  &  wire32633 ) ;
 assign wire3696 = ( n_n6710  &  wire32638 ) | ( wire4804  &  wire32638 ) | ( wire4805  &  wire32638 ) ;
 assign wire3698 = ( (~ pi16)  &  wire3703 ) | ( (~ pi16)  &  wire32639 ) ;
 assign wire3702 = ( (~ pi20)  &  pi25  &  wire153  &  wire188 ) ;
 assign wire3703 = ( (~ pi25)  &  wire169  &  wire4458 ) | ( (~ pi25)  &  wire169  &  wire4459 ) ;
 assign wire3704 = ( pi19  &  wire440 ) ;
 assign wire3706 = ( pi17  &  pi19  &  (~ pi16)  &  wire221 ) ;
 assign wire3708 = ( wire374  &  wire32922 ) | ( wire214  &  n_n7905  &  wire32922 ) ;
 assign wire3709 = ( wire375  &  wire32925 ) | ( wire214  &  n_n7905  &  wire32925 ) ;
 assign wire3710 = ( wire374  &  wire32927 ) | ( wire214  &  n_n7913  &  wire32927 ) ;
 assign wire3711 = ( wire375  &  wire32929 ) | ( wire214  &  n_n7913  &  wire32929 ) ;
 assign wire3712 = ( wire3759  &  wire32931 ) | ( pi20  &  n_n6749  &  wire32931 ) ;
 assign wire3715 = ( wire221  &  wire185  &  wire32939 ) ;
 assign wire3716 = ( wire3989  &  wire32941 ) | ( wire3990  &  wire32941 ) | ( wire3991  &  wire32941 ) ;
 assign wire3717 = ( wire32948  &  wire32949 ) | ( n_n7885  &  wire32943  &  wire32949 ) ;
 assign wire3719 = ( wire1339  &  wire31875 ) | ( wire1339  &  wire31876 ) | ( wire1339  &  wire31916 ) ;
 assign wire3720 = ( wire1094  &  wire3731 ) | ( wire1094  &  wire32978 ) | ( wire1094  &  wire32979 ) ;
 assign wire3721 = ( wire1094  &  wire3743 ) | ( wire1094  &  wire33010 ) | ( wire1094  &  wire33011 ) ;
 assign wire3724 = ( wire375  &  wire32954 ) | ( wire3838  &  wire32954 ) ;
 assign wire3725 = ( wire374  &  wire32955 ) | ( wire3969  &  wire32955 ) ;
 assign wire3727 = ( wire3759  &  wire32957 ) | ( pi20  &  n_n6749  &  wire32957 ) ;
 assign wire3728 = ( wire3834  &  wire32962 ) | ( wire3835  &  wire32962 ) | ( wire32960  &  wire32962 ) ;
 assign wire3729 = ( wire3951  &  wire32963 ) | ( wire3952  &  wire32963 ) | ( wire31859  &  wire32963 ) ;
 assign wire3730 = ( pi16  &  wire221  &  wire185 ) ;
 assign wire3731 = ( pi27  &  wire3826 ) | ( (~ pi26)  &  wire3826 ) | ( pi27  &  wire32964 ) | ( (~ pi26)  &  wire32964 ) ;
 assign wire3732 = ( (~ wire155)  &  wire3828 ) | ( (~ wire155)  &  wire3830 ) | ( (~ wire155)  &  wire32970 ) ;
 assign wire3735 = ( wire375  &  wire32984 ) | ( wire3870  &  wire32984 ) ;
 assign wire3736 = ( wire3863  &  wire32985 ) | ( wire3864  &  wire32985 ) ;
 assign wire3737 = ( wire3865  &  wire32989 ) | ( wire3866  &  wire32989 ) | ( wire3867  &  wire32989 ) ;
 assign wire3739 = ( wire375  &  wire32991 ) | ( wire3868  &  wire32991 ) ;
 assign wire3741 = ( (~ pi22)  &  wire698  &  nv5285  &  wire204 ) ;
 assign wire3743 = ( pi27  &  wire3855 ) | ( (~ pi26)  &  wire3855 ) | ( pi27  &  wire32995 ) | ( (~ pi26)  &  wire32995 ) ;
 assign wire3744 = ( (~ wire155)  &  wire3857 ) | ( (~ wire155)  &  wire3858 ) | ( (~ wire155)  &  wire33001 ) ;
 assign wire3748 = ( wire374  &  wire33014 ) | ( wire214  &  n_n7837  &  wire33014 ) ;
 assign wire3749 = ( wire375  &  wire33016 ) | ( wire214  &  n_n7837  &  wire33016 ) ;
 assign wire3750 = ( wire374  &  wire33017 ) | ( wire214  &  n_n7845  &  wire33017 ) ;
 assign wire3751 = ( wire375  &  wire33018 ) | ( wire214  &  n_n7845  &  wire33018 ) ;
 assign wire3752 = ( wire3759  &  wire33019 ) | ( pi20  &  n_n6749  &  wire33019 ) ;
 assign wire3755 = ( pi16  &  wire221  &  wire185 ) ;
 assign wire3756 = ( wire155  &  wire4027 ) | ( wire155  &  wire4028 ) | ( wire155  &  wire4029 ) ;
 assign wire3757 = ( (~ pi27)  &  pi26  &  wire4037 ) | ( (~ pi27)  &  pi26  &  wire33032 ) ;
 assign wire3759 = ( pi21  &  (~ pi22)  &  pi20  &  nv5285 ) ;
 assign wire3761 = ( wire374  &  wire33057 ) | ( wire214  &  n_n7913  &  wire33057 ) ;
 assign wire3762 = ( wire375  &  wire33060 ) | ( wire214  &  n_n7913  &  wire33060 ) ;
 assign wire3763 = ( wire375  &  wire33062 ) | ( wire214  &  n_n7905  &  wire33062 ) ;
 assign wire3764 = ( wire374  &  wire33064 ) | ( wire214  &  n_n7905  &  wire33064 ) ;
 assign wire3765 = ( wire3823  &  wire33066 ) | ( (~ pi20)  &  n_n7095  &  wire33066 ) ;
 assign wire3768 = ( wire227  &  wire198  &  wire33071 ) ;
 assign wire3769 = ( wire3989  &  wire33072 ) | ( wire3990  &  wire33072 ) | ( wire3991  &  wire33072 ) ;
 assign wire3770 = ( wire32948  &  wire33073 ) | ( n_n7885  &  wire32943  &  wire33073 ) ;
 assign wire3773 = ( wire1079  &  wire3820 ) | ( wire1079  &  wire33108 ) | ( wire1079  &  wire33109 ) ;
 assign wire3774 = ( wire1079  &  wire3851 ) | ( wire1079  &  wire33127 ) | ( wire1079  &  wire33128 ) ;
 assign wire3777 = ( wire845  &  wire3788 ) | ( wire845  &  wire33169 ) | ( wire845  &  wire33170 ) ;
 assign wire3778 = ( wire845  &  wire3798 ) | ( wire845  &  wire33183 ) | ( wire845  &  wire33184 ) ;
 assign wire3779 = ( wire618  &  wire31875 ) | ( wire618  &  wire31876 ) | ( wire618  &  wire31916 ) ;
 assign wire3780 = ( (~ ni11)  &  wire3889 ) | ( (~ ni11)  &  wire31995 ) ;
 assign wire3782 = ( wire374  &  wire33159 ) | ( wire3969  &  wire33159 ) ;
 assign wire3783 = ( wire374  &  wire33160 ) | ( wire3963  &  wire33160 ) ;
 assign wire3785 = ( wire3834  &  wire33162 ) | ( wire3835  &  wire33162 ) | ( wire32960  &  wire33162 ) ;
 assign wire3786 = ( wire3951  &  wire33163 ) | ( wire3952  &  wire33163 ) | ( wire31859  &  wire33163 ) ;
 assign wire3788 = ( (~ pi27)  &  wire3826 ) | ( (~ pi27)  &  wire32964 ) ;
 assign wire3789 = ( pi27  &  wire3828 ) | ( pi27  &  wire3830 ) | ( pi27  &  wire32970 ) ;
 assign wire3792 = ( wire374  &  wire33173 ) | ( wire3955  &  wire33173 ) ;
 assign wire3793 = ( wire374  &  wire33174 ) | ( wire3975  &  wire33174 ) ;
 assign wire3795 = ( (~ pi27)  &  (~ pi16)  &  wire3863 ) | ( (~ pi27)  &  (~ pi16)  &  wire3864 ) ;
 assign wire3796 = ( wire3865  &  wire33177 ) | ( wire3866  &  wire33177 ) | ( wire3867  &  wire33177 ) ;
 assign wire3798 = ( (~ pi27)  &  wire3855 ) | ( (~ pi27)  &  wire32995 ) ;
 assign wire3799 = ( pi27  &  wire3857 ) | ( pi27  &  wire3858 ) | ( pi27  &  wire33001 ) ;
 assign wire3801 = ( wire374  &  wire33076 ) | ( wire214  &  n_n7845  &  wire33076 ) ;
 assign wire3802 = ( wire375  &  wire33078 ) | ( wire214  &  n_n7845  &  wire33078 ) ;
 assign wire3803 = ( wire375  &  wire33079 ) | ( wire214  &  n_n7837  &  wire33079 ) ;
 assign wire3804 = ( wire374  &  wire33080 ) | ( wire214  &  n_n7837  &  wire33080 ) ;
 assign wire3805 = ( wire3823  &  wire33081 ) | ( (~ pi20)  &  n_n7095  &  wire33081 ) ;
 assign wire3808 = ( pi16  &  wire227  &  wire198 ) ;
 assign wire3809 = ( wire156  &  wire4027 ) | ( wire156  &  wire4028 ) | ( wire156  &  wire4029 ) ;
 assign wire3810 = ( (~ pi27)  &  (~ pi26)  &  wire4037 ) | ( (~ pi27)  &  (~ pi26)  &  wire33032 ) ;
 assign wire3813 = ( wire375  &  wire33096 ) | ( wire3840  &  wire33096 ) ;
 assign wire3814 = ( wire375  &  wire33097 ) | ( wire3838  &  wire33097 ) ;
 assign wire3816 = ( wire3823  &  wire33099 ) | ( (~ pi20)  &  n_n7095  &  wire33099 ) ;
 assign wire3817 = ( wire3834  &  wire33100 ) | ( wire3835  &  wire33100 ) | ( wire32960  &  wire33100 ) ;
 assign wire3818 = ( wire3951  &  wire33101 ) | ( wire3952  &  wire33101 ) | ( wire31859  &  wire33101 ) ;
 assign wire3819 = ( pi16  &  wire227  &  wire198 ) ;
 assign wire3820 = ( pi27  &  wire3826 ) | ( pi26  &  wire3826 ) | ( pi27  &  wire32964 ) | ( pi26  &  wire32964 ) ;
 assign wire3821 = ( (~ wire156)  &  wire3828 ) | ( (~ wire156)  &  wire3830 ) | ( (~ wire156)  &  wire32970 ) ;
 assign wire3823 = ( pi21  &  (~ pi22)  &  (~ pi20)  &  nv4938 ) ;
 assign wire3826 = ( wire180  &  wire374  &  wire154 ) | ( wire180  &  wire154  &  wire3961 ) ;
 assign wire3827 = ( pi17  &  pi16  &  wire152  &  nv4630 ) ;
 assign wire3828 = ( wire31510  &  wire32965 ) | ( wire31511  &  wire32965 ) | ( wire31512  &  wire32965 ) ;
 assign wire3829 = ( wire928  &  wire32966 ) | ( wire4680  &  wire32966 ) | ( wire4681  &  wire32966 ) ;
 assign wire3830 = ( wire31428  &  wire32967 ) | ( wire31429  &  wire32967 ) | ( wire31430  &  wire32967 ) ;
 assign wire3834 = ( n_n6710  &  wire32958 ) | ( wire4787  &  wire32958 ) | ( wire4788  &  wire32958 ) ;
 assign wire3835 = ( n_n6710  &  wire32959 ) | ( wire4781  &  wire32959 ) | ( wire4782  &  wire32959 ) ;
 assign wire3838 = ( wire214  &  wire31674 ) | ( wire214  &  wire31675 ) | ( wire214  &  wire31676 ) ;
 assign wire3840 = ( wire214  &  wire31756 ) | ( wire214  &  wire31757 ) | ( wire214  &  wire31758 ) ;
 assign wire3842 = ( wire3863  &  wire33111 ) | ( wire3864  &  wire33111 ) ;
 assign wire3843 = ( wire3865  &  wire33112 ) | ( wire3866  &  wire33112 ) | ( wire3867  &  wire33112 ) ;
 assign wire3845 = ( wire374  &  wire33114 ) | ( wire3955  &  wire33114 ) ;
 assign wire3846 = ( wire374  &  wire33115 ) | ( wire3975  &  wire33115 ) ;
 assign wire3849 = ( (~ pi22)  &  wire211  &  wire698  &  nv4938 ) ;
 assign wire3851 = ( pi27  &  wire3855 ) | ( pi26  &  wire3855 ) | ( pi27  &  wire32995 ) | ( pi26  &  wire32995 ) ;
 assign wire3852 = ( (~ wire156)  &  wire3857 ) | ( (~ wire156)  &  wire3858 ) | ( (~ wire156)  &  wire33001 ) ;
 assign wire3855 = ( wire158  &  wire180  &  wire374 ) | ( wire158  &  wire180  &  wire3957 ) ;
 assign wire3856 = ( pi17  &  (~ pi16)  &  wire152  &  nv4575 ) ;
 assign wire3857 = ( wire31252  &  wire32996 ) | ( wire31253  &  wire32996 ) | ( wire31254  &  wire32996 ) ;
 assign wire3858 = ( wire31338  &  wire32997 ) | ( wire31339  &  wire32997 ) | ( wire31340  &  wire32997 ) ;
 assign wire3859 = ( wire4613  &  wire32998 ) | ( wire31347  &  wire32998 ) ;
 assign wire3863 = ( pi20  &  wire374  &  wire153 ) | ( pi20  &  wire153  &  wire3973 ) ;
 assign wire3864 = ( (~ pi20)  &  wire374  &  wire153 ) | ( (~ pi20)  &  wire153  &  wire3977 ) ;
 assign wire3865 = ( n_n6710  &  wire32986 ) | ( wire4807  &  wire32986 ) | ( wire4808  &  wire32986 ) ;
 assign wire3866 = ( n_n6710  &  wire32987 ) | ( wire4813  &  wire32987 ) | ( wire4814  &  wire32987 ) ;
 assign wire3867 = ( pi20  &  wire153  &  wire375 ) | ( (~ pi20)  &  wire153  &  wire375 ) ;
 assign wire3868 = ( wire214  &  wire31838 ) | ( wire214  &  wire31839 ) | ( wire214  &  wire31840 ) ;
 assign wire3870 = ( wire214  &  wire31592 ) | ( wire214  &  wire31593 ) | ( wire214  &  wire31594 ) ;
 assign wire3874 = ( wire3912  &  wire31926 ) | ( pi19  &  wire170  &  wire31926 ) ;
 assign wire3878 = ( n_n6710  &  wire31934 ) | ( wire4810  &  wire31934 ) | ( wire4811  &  wire31934 ) ;
 assign wire3879 = ( wire31937  &  wire31939 ) | ( n_n7885  &  wire329  &  wire31939 ) ;
 assign wire3880 = ( n_n6710  &  wire31940 ) | ( wire4778  &  wire31940 ) | ( wire4779  &  wire31940 ) ;
 assign wire3881 = ( n_n6710  &  wire31941 ) | ( wire4784  &  wire31941 ) | ( wire4785  &  wire31941 ) ;
 assign wire3882 = ( wire3908  &  wire31943 ) | ( wire344  &  wire170  &  wire31943 ) ;
 assign wire3883 = ( wire3910  &  wire31944 ) | ( wire340  &  wire170  &  wire31944 ) ;
 assign wire3884 = ( wire3912  &  wire31945 ) | ( pi19  &  wire170  &  wire31945 ) ;
 assign wire3888 = ( wire31949  &  wire31950 ) | ( wire178  &  n_n7825  &  wire31950 ) ;
 assign wire3889 = ( wire613  &  wire31875 ) | ( wire613  &  wire31876 ) | ( wire613  &  wire31916 ) ;
 assign wire3891 = ( wire31838  &  wire31952 ) | ( wire31839  &  wire31952 ) | ( wire31840  &  wire31952 ) ;
 assign wire3892 = ( wire31592  &  wire31954 ) | ( wire31593  &  wire31954 ) | ( wire31594  &  wire31954 ) ;
 assign wire3893 = ( wire3912  &  wire31955 ) | ( pi19  &  wire170  &  wire31955 ) ;
 assign wire3894 = ( wire31674  &  wire31956 ) | ( wire31675  &  wire31956 ) | ( wire31676  &  wire31956 ) ;
 assign wire3895 = ( wire31756  &  wire31957 ) | ( wire31757  &  wire31957 ) | ( wire31758  &  wire31957 ) ;
 assign wire3896 = ( n_n6710  &  wire31958 ) | ( wire4807  &  wire31958 ) | ( wire4808  &  wire31958 ) ;
 assign wire3897 = ( n_n6710  &  wire31959 ) | ( wire4813  &  wire31959 ) | ( wire4814  &  wire31959 ) ;
 assign wire3898 = ( wire4608  &  wire31962 ) | ( wire4609  &  wire31962 ) | ( wire31960  &  wire31962 ) ;
 assign wire3899 = ( n_n6710  &  wire1327 ) | ( wire1327  &  wire4781 ) | ( wire1327  &  wire4782 ) ;
 assign wire3900 = ( n_n6710  &  wire1324 ) | ( wire1324  &  wire4787 ) | ( wire1324  &  wire4788 ) ;
 assign wire3902 = ( (~ pi15)  &  wire3908 ) | ( (~ pi15)  &  wire344  &  wire170 ) ;
 assign wire3903 = ( wire258  &  wire3910 ) | ( wire340  &  wire258  &  wire170 ) ;
 assign wire3904 = ( wire614  &  wire1178 ) | ( wire614  &  wire4687 ) | ( wire614  &  wire4688 ) ;
 assign wire3906 = ( (~ pi15)  &  n_n9245  &  wire152  &  wire154 ) ;
 assign wire3907 = ( wire507  &  wire3912 ) | ( pi19  &  wire170  &  wire507 ) ;
 assign wire3908 = ( (~ pi16)  &  ni32  &  ni30  &  wire153 ) ;
 assign wire3910 = ( pi20  &  ni32  &  ni30  &  wire153 ) | ( (~ pi20)  &  ni32  &  ni30  &  wire153 ) ;
 assign wire3912 = ( ni32  &  ni30  &  wire152 ) ;
 assign wire3914 = ( wire374  &  wire31878 ) | ( wire214  &  n_n7893  &  wire31878 ) ;
 assign wire3915 = ( wire374  &  wire31880 ) | ( n_n7885  &  wire214  &  wire31880 ) ;
 assign wire3916 = ( wire374  &  wire31882 ) | ( wire214  &  n_n7877  &  wire31882 ) ;
 assign wire3918 = ( wire374  &  wire31884 ) | ( wire214  &  n_n7913  &  wire31884 ) ;
 assign wire3919 = ( wire374  &  wire31885 ) | ( wire214  &  n_n7905  &  wire31885 ) ;
 assign wire3920 = ( wire374  &  wire31886 ) | ( wire214  &  n_n7816  &  wire31886 ) ;
 assign wire3921 = ( wire374  &  wire31887 ) | ( wire214  &  n_n7825  &  wire31887 ) ;
 assign wire3922 = ( wire374  &  wire31888 ) | ( wire214  &  n_n7837  &  wire31888 ) ;
 assign wire3923 = ( wire374  &  wire31889 ) | ( wire214  &  n_n7845  &  wire31889 ) ;
 assign wire3926 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire170 ) ;
 assign wire3927 = ( pi19  &  wire395  &  wire170 ) ;
 assign wire3929 = ( (~ pi19)  &  wire403  &  wire170 ) ;
 assign wire3930 = ( pi16  &  pi15  &  wire4046 ) | ( pi16  &  pi15  &  wire31899 ) ;
 assign wire3931 = ( wire416  &  wire374 ) | ( wire416  &  wire214  &  n_n7808 ) ;
 assign wire3934 = ( wire374  &  wire31343 ) | ( wire3957  &  wire31343 ) ;
 assign wire3937 = ( wire180  &  wire374  &  wire614 ) | ( wire180  &  wire614  &  wire3961 ) ;
 assign wire3938 = ( wire178  &  wire374  &  wire614 ) | ( wire178  &  wire614  &  wire3965 ) ;
 assign wire3939 = ( wire374  &  wire31596 ) | ( wire3955  &  wire31596 ) ;
 assign wire3940 = ( wire182  &  wire374  &  wire507 ) | ( wire182  &  wire507  &  wire3963 ) ;
 assign wire3941 = ( wire179  &  wire374  &  wire507 ) | ( wire179  &  wire507  &  wire3969 ) ;
 assign wire3942 = ( wire374  &  wire31842 ) | ( wire3975  &  wire31842 ) ;
 assign wire3943 = ( wire374  &  wire31846 ) | ( wire3977  &  wire31846 ) ;
 assign wire3944 = ( wire374  &  wire31849 ) | ( wire3973  &  wire31849 ) ;
 assign wire3945 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire170 ) ;
 assign wire3946 = ( pi19  &  wire170  &  wire507 ) ;
 assign wire3948 = ( (~ pi19)  &  wire170  &  wire614 ) ;
 assign wire3950 = ( wire258  &  wire3951 ) | ( wire258  &  wire3952 ) | ( wire258  &  wire31859 ) ;
 assign wire3951 = ( n_n6710  &  wire31855 ) | ( wire4787  &  wire31855 ) | ( wire4788  &  wire31855 ) ;
 assign wire3952 = ( n_n6710  &  wire31858 ) | ( wire4781  &  wire31858 ) | ( wire4782  &  wire31858 ) ;
 assign wire3955 = ( wire214  &  wire31592 ) | ( wire214  &  wire31593 ) | ( wire214  &  wire31594 ) ;
 assign wire3957 = ( wire214  &  wire31338 ) | ( wire214  &  wire31339 ) | ( wire214  &  wire31340 ) ;
 assign wire3959 = ( wire214  &  wire31252 ) | ( wire214  &  wire31253 ) | ( wire214  &  wire31254 ) ;
 assign wire3961 = ( wire214  &  wire31428 ) | ( wire214  &  wire31429 ) | ( wire214  &  wire31430 ) ;
 assign wire3963 = ( wire214  &  wire31674 ) | ( wire214  &  wire31675 ) | ( wire214  &  wire31676 ) ;
 assign wire3965 = ( wire214  &  wire31510 ) | ( wire214  &  wire31511 ) | ( wire214  &  wire31512 ) ;
 assign wire3969 = ( wire214  &  wire31756 ) | ( wire214  &  wire31757 ) | ( wire214  &  wire31758 ) ;
 assign wire3973 = ( n_n6710  &  wire214 ) | ( wire214  &  wire4813 ) | ( wire214  &  wire4814 ) ;
 assign wire3975 = ( wire214  &  wire31838 ) | ( wire214  &  wire31839 ) | ( wire214  &  wire31840 ) ;
 assign wire3977 = ( n_n6710  &  wire214 ) | ( wire214  &  wire4807 ) | ( wire214  &  wire4808 ) ;
 assign wire3979 = ( wire375  &  wire33130 ) | ( wire214  &  n_n7913  &  wire33130 ) ;
 assign wire3980 = ( wire374  &  wire33131 ) | ( wire214  &  n_n7913  &  wire33131 ) ;
 assign wire3981 = ( wire374  &  wire33132 ) | ( wire214  &  n_n7905  &  wire33132 ) ;
 assign wire3982 = ( wire375  &  wire33133 ) | ( wire214  &  n_n7905  &  wire33133 ) ;
 assign wire3986 = ( (~ pi27)  &  wire3989 ) | ( (~ pi27)  &  wire3990 ) | ( (~ pi27)  &  wire3991 ) ;
 assign wire3987 = ( pi27  &  wire32948 ) | ( pi27  &  n_n7885  &  wire32943 ) ;
 assign wire3989 = ( wire374  &  wire250 ) | ( wire214  &  wire250  &  n_n7893 ) ;
 assign wire3990 = ( wire374  &  wire243 ) | ( n_n7885  &  wire214  &  wire243 ) ;
 assign wire3991 = ( wire374  &  wire194 ) | ( wire214  &  wire194  &  n_n7877 ) ;
 assign wire4005 = ( n_n6710  &  wire32933 ) | ( wire4810  &  wire32933 ) | ( wire4811  &  wire32933 ) ;
 assign wire4006 = ( pi20  &  wire153  &  wire375 ) | ( (~ pi20)  &  wire153  &  wire375 ) ;
 assign wire4017 = ( wire375  &  wire33144 ) | ( wire214  &  n_n7845  &  wire33144 ) ;
 assign wire4018 = ( wire374  &  wire33145 ) | ( wire214  &  n_n7845  &  wire33145 ) ;
 assign wire4019 = ( wire374  &  wire33146 ) | ( wire214  &  n_n7837  &  wire33146 ) ;
 assign wire4020 = ( wire375  &  wire33147 ) | ( wire214  &  n_n7837  &  wire33147 ) ;
 assign wire4024 = ( (~ pi27)  &  wire4027 ) | ( (~ pi27)  &  wire4028 ) | ( (~ pi27)  &  wire4029 ) ;
 assign wire4025 = ( pi27  &  wire33032 ) | ( pi27  &  n_n7825  &  wire33027 ) ;
 assign wire4027 = ( wire374  &  wire251 ) | ( wire214  &  n_n7825  &  wire251 ) ;
 assign wire4028 = ( wire374  &  wire244 ) | ( wire214  &  n_n7816  &  wire244 ) ;
 assign wire4029 = ( wire374  &  wire183 ) | ( wire214  &  wire183  &  n_n7808 ) ;
 assign wire4037 = ( (~ ni29)  &  n_n7825  &  wire251 ) | ( (~ n_n8352)  &  n_n7825  &  wire251 ) ;
 assign wire4043 = ( n_n6710  &  wire33021 ) | ( wire4784  &  wire33021 ) | ( wire4785  &  wire33021 ) ;
 assign wire4044 = ( pi20  &  wire153  &  wire375 ) | ( (~ pi20)  &  wire153  &  wire375 ) ;
 assign wire4046 = ( n_n6710  &  wire31898 ) | ( wire4784  &  wire31898 ) | ( wire4785  &  wire31898 ) ;
 assign wire4047 = ( pi20  &  wire374  &  wire153 ) | ( (~ pi20)  &  wire374  &  wire153 ) ;
 assign wire4061 = ( ni32  &  (~ ni30)  &  ni29 ) ;
 assign wire4062 = ( wire31756  &  wire32685 ) | ( wire31757  &  wire32685 ) | ( wire31758  &  wire32685 ) ;
 assign wire4064 = ( wire31674  &  wire32689 ) | ( wire31675  &  wire32689 ) | ( wire31676  &  wire32689 ) ;
 assign wire4065 = ( wire31510  &  wire32691 ) | ( wire31511  &  wire32691 ) | ( wire31512  &  wire32691 ) ;
 assign wire4066 = ( n_n6710  &  wire32693 ) | ( wire4781  &  wire32693 ) | ( wire4782  &  wire32693 ) ;
 assign wire4067 = ( wire4079  &  wire32694 ) | ( wire182  &  wire280  &  wire32694 ) ;
 assign wire4069 = ( wire4090  &  wire32696 ) | ( wire32587  &  wire32696 ) ;
 assign wire4070 = ( n_n6710  &  wire32697 ) | ( wire4787  &  wire32697 ) | ( wire4788  &  wire32697 ) ;
 assign wire4072 = ( pi16  &  wire4078 ) | ( pi16  &  wire32617 ) ;
 assign wire4073 = ( wire154  &  wire4083 ) | ( wire180  &  wire154  &  wire280 ) ;
 assign wire4077 = ( pi20  &  pi25  &  wire153  &  wire188 ) ;
 assign wire4078 = ( (~ pi25)  &  wire171  &  wire4458 ) | ( (~ pi25)  &  wire171  &  wire4459 ) ;
 assign wire4079 = ( pi19  &  wire373 ) ;
 assign wire4082 = ( pi17  &  pi19  &  pi16  &  wire221 ) ;
 assign wire4083 = ( (~ pi19)  &  wire373 ) ;
 assign wire4089 = ( n_n9245  &  wire155  &  wire181 ) | ( (~ wire155)  &  n_n8085  &  wire181 ) ;
 assign wire4090 = ( (~ pi25)  &  (~ wire150)  &  wire4458 ) | ( (~ pi25)  &  (~ wire150)  &  wire4459 ) ;
 assign wire4096 = ( wire4147  &  wire32722 ) | ( wire152  &  wire249  &  wire32722 ) ;
 assign wire4100 = ( wire4145  &  wire32728 ) | ( wire151  &  wire249  &  wire32728 ) ;
 assign wire4101 = ( wire4149  &  wire32729 ) | ( wire153  &  wire249  &  wire32729 ) ;
 assign wire4102 = ( n_n6922  &  wire32730 ) | ( wire4435  &  wire32730 ) | ( wire4436  &  wire32730 ) ;
 assign wire4107 = ( (~ pi15)  &  wire268  &  wire32771 ) | ( (~ pi15)  &  wire268  &  wire32772 ) ;
 assign wire4108 = ( wire818  &  wire4170 ) | ( wire818  &  wire32904 ) ;
 assign wire4109 = ( wire618  &  wire32053 ) | ( (~ pi15)  &  n_n9255  &  wire618 ) ;
 assign wire4112 = ( (~ pi17)  &  (~ pi16)  &  wire358  &  n_n7913 ) ;
 assign wire4113 = ( wire4147  &  wire32735 ) | ( wire152  &  wire249  &  wire32735 ) ;
 assign wire4115 = ( pi17  &  (~ pi16)  &  wire345  &  n_n7893 ) ;
 assign wire4117 = ( wire158  &  wire4145 ) | ( wire158  &  wire151  &  wire249 ) ;
 assign wire4118 = ( (~ pi16)  &  wire4149 ) | ( (~ pi16)  &  wire153  &  wire249 ) ;
 assign wire4121 = ( wire31674  &  wire32746 ) | ( wire31675  &  wire32746 ) | ( wire31676  &  wire32746 ) ;
 assign wire4122 = ( wire31756  &  wire32748 ) | ( wire31757  &  wire32748 ) | ( wire31758  &  wire32748 ) ;
 assign wire4123 = ( wire4147  &  wire32749 ) | ( wire152  &  wire249  &  wire32749 ) ;
 assign wire4124 = ( wire31510  &  wire32750 ) | ( wire31511  &  wire32750 ) | ( wire31512  &  wire32750 ) ;
 assign wire4127 = ( wire154  &  wire4145 ) | ( wire151  &  wire154  &  wire249 ) ;
 assign wire4128 = ( pi16  &  wire4149 ) | ( pi16  &  wire153  &  wire249 ) ;
 assign wire4129 = ( wire257  &  n_n6922 ) | ( wire257  &  wire4435 ) | ( wire257  &  wire4436 ) ;
 assign wire4132 = ( wire31592  &  wire32761 ) | ( wire31593  &  wire32761 ) | ( wire31594  &  wire32761 ) ;
 assign wire4134 = ( wire4147  &  wire32763 ) | ( wire152  &  wire249  &  wire32763 ) ;
 assign wire4135 = ( wire31252  &  wire32764 ) | ( wire31253  &  wire32764 ) | ( wire31254  &  wire32764 ) ;
 assign wire4138 = ( wire158  &  wire4145 ) | ( wire158  &  wire151  &  wire249 ) ;
 assign wire4139 = ( (~ pi16)  &  wire4149 ) | ( (~ pi16)  &  wire153  &  wire249 ) ;
 assign wire4142 = ( wire295  &  n_n6922 ) | ( wire295  &  wire4435 ) | ( wire295  &  wire4436 ) ;
 assign wire4145 = ( (~ pi19)  &  n_n6922 ) | ( (~ pi19)  &  wire4435 ) | ( (~ pi19)  &  wire4436 ) ;
 assign wire4147 = ( pi19  &  n_n6922 ) | ( pi19  &  wire4435 ) | ( pi19  &  wire4436 ) ;
 assign wire4149 = ( wire163  &  n_n6922 ) | ( wire163  &  wire4435 ) | ( wire163  &  wire4436 ) ;
 assign wire4151 = ( (~ pi27)  &  pi25  &  ni32  &  ni30 ) ;
 assign wire4158 = ( wire4220  &  wire32791 ) | ( wire182  &  wire274  &  wire32791 ) ;
 assign wire4161 = ( wire228  &  wire4236  &  wire32796 ) | ( wire228  &  wire32777  &  wire32796 ) ;
 assign wire4162 = ( wire219  &  wire4779  &  wire32798 ) | ( wire219  &  wire31895  &  wire32798 ) ;
 assign wire4163 = ( wire4187  &  wire32799 ) | ( wire178  &  wire274  &  wire32799 ) ;
 assign wire4164 = ( wire4232  &  wire32801 ) | ( wire32800  &  wire32801 ) ;
 assign wire4165 = ( (~ ni14)  &  wire485  &  wire227 ) ;
 assign wire4167 = ( pi15  &  (~ ni14)  &  n_n7808  &  wire311 ) ;
 assign wire4170 = ( (~ pi15)  &  (~ ni14)  &  wire32887 ) | ( (~ pi15)  &  (~ ni14)  &  wire32888 ) ;
 assign wire4175 = ( (~ pi17)  &  (~ pi16)  &  wire358  &  n_n7913 ) ;
 assign wire4176 = ( wire4204  &  wire32814 ) | ( wire179  &  wire274  &  wire32814 ) ;
 assign wire4179 = ( wire4236  &  wire32817 ) | ( wire32777  &  wire32817 ) ;
 assign wire4182 = ( (~ pi25)  &  wire4448  &  wire32820 ) | ( (~ pi25)  &  wire4449  &  wire32820 ) ;
 assign wire4183 = ( pi17  &  (~ pi16)  &  wire345  &  n_n7893 ) ;
 assign wire4184 = ( wire158  &  wire4187 ) | ( wire158  &  wire178  &  wire274 ) ;
 assign wire4187 = ( (~ pi19)  &  wire372 ) ;
 assign wire4189 = ( wire31674  &  wire32837 ) | ( wire31675  &  wire32837 ) | ( wire31676  &  wire32837 ) ;
 assign wire4191 = ( wire31756  &  wire32841 ) | ( wire31757  &  wire32841 ) | ( wire31758  &  wire32841 ) ;
 assign wire4192 = ( wire31510  &  wire32843 ) | ( wire31511  &  wire32843 ) | ( wire31512  &  wire32843 ) ;
 assign wire4193 = ( n_n6710  &  wire32845 ) | ( wire4787  &  wire32845 ) | ( wire4788  &  wire32845 ) ;
 assign wire4194 = ( wire4204  &  wire32846 ) | ( wire179  &  wire274  &  wire32846 ) ;
 assign wire4196 = ( wire4236  &  wire32848 ) | ( wire32777  &  wire32848 ) ;
 assign wire4197 = ( n_n6710  &  wire32849 ) | ( wire4781  &  wire32849 ) | ( wire4782  &  wire32849 ) ;
 assign wire4199 = ( wire154  &  wire4222 ) | ( wire180  &  wire154  &  wire274 ) ;
 assign wire4200 = ( pi16  &  wire4232 ) | ( pi16  &  wire32800 ) ;
 assign wire4201 = ( pi17  &  pi16  &  wire152  &  wire274 ) ;
 assign wire4204 = ( pi19  &  wire372 ) ;
 assign wire4206 = ( wire31592  &  wire32865 ) | ( wire31593  &  wire32865 ) | ( wire31594  &  wire32865 ) ;
 assign wire4208 = ( wire31252  &  wire32869 ) | ( wire31253  &  wire32869 ) | ( wire31254  &  wire32869 ) ;
 assign wire4209 = ( n_n6710  &  wire32871 ) | ( wire4813  &  wire32871 ) | ( wire4814  &  wire32871 ) ;
 assign wire4211 = ( wire4220  &  wire32873 ) | ( wire182  &  wire274  &  wire32873 ) ;
 assign wire4213 = ( wire4236  &  wire32875 ) | ( wire32777  &  wire32875 ) ;
 assign wire4214 = ( n_n6710  &  wire32876 ) | ( wire4807  &  wire32876 ) | ( wire4808  &  wire32876 ) ;
 assign wire4216 = ( wire158  &  wire4222 ) | ( wire158  &  wire180  &  wire274 ) ;
 assign wire4217 = ( (~ pi16)  &  wire4232 ) | ( (~ pi16)  &  wire32800 ) ;
 assign wire4220 = ( pi19  &  wire442 ) ;
 assign wire4222 = ( (~ pi19)  &  wire442 ) ;
 assign wire4226 = ( pi17  &  pi19  &  (~ pi16)  &  wire227 ) ;
 assign wire4231 = ( (~ pi20)  &  pi25  &  wire153  &  wire187 ) ;
 assign wire4232 = ( (~ pi25)  &  wire169  &  wire4448 ) | ( (~ pi25)  &  wire169  &  wire4449 ) ;
 assign wire4235 = ( n_n9245  &  wire156  &  wire181 ) | ( (~ wire156)  &  n_n8085  &  wire181 ) ;
 assign wire4236 = ( (~ pi25)  &  (~ wire150)  &  wire4448 ) | ( (~ pi25)  &  (~ wire150)  &  wire4449 ) ;
 assign wire4240 = ( wire306  &  wire32493 ) | ( wire233  &  n_n7905  &  wire32493 ) ;
 assign wire4241 = ( wire305  &  wire32496 ) | ( wire233  &  n_n7905  &  wire32496 ) ;
 assign wire4242 = ( (~ wire150)  &  wire4433  &  wire32498 ) | ( (~ wire150)  &  wire4434  &  wire32498 ) ;
 assign wire4243 = ( wire4273  &  wire32500 ) | ( wire4276  &  wire32500 ) | ( wire32228  &  wire32500 ) ;
 assign wire4244 = ( wire4365  &  wire32502 ) | ( pi20  &  n_n6410  &  wire32502 ) ;
 assign wire4245 = ( wire449  &  wire32504 ) | ( wire4491  &  wire32504 ) ;
 assign wire4246 = ( (~ wire165)  &  wire4295  &  wire32505 ) | ( (~ wire165)  &  wire32338  &  wire32505 ) ;
 assign wire4247 = ( wire185  &  wire339  &  wire32507 ) ;
 assign wire4248 = ( wire4264  &  wire32508 ) | ( wire4266  &  wire32508 ) | ( wire32406  &  wire32508 ) ;
 assign wire4249 = ( wire4281  &  wire32509 ) | ( wire263  &  wire453  &  wire32509 ) ;
 assign wire4250 = ( wire4282  &  wire32510 ) | ( wire4283  &  wire32510 ) | ( wire4284  &  wire32510 ) ;
 assign wire4252 = ( pi15  &  (~ wire289)  &  wire158  &  wire339 ) ;
 assign wire4253 = ( wire708  &  wire4337 ) | ( wire708  &  wire32531 ) | ( wire708  &  wire32532 ) ;
 assign wire4254 = ( wire708  &  wire4363 ) | ( wire708  &  wire32545 ) | ( wire708  &  wire32546 ) ;
 assign wire4255 = ( pi15  &  (~ wire289)  &  wire32563 ) | ( pi15  &  (~ wire289)  &  wire32564 ) ;
 assign wire4257 = ( (~ pi27)  &  pi24  &  nv3908  &  wire32382 ) ;
 assign wire4258 = ( n_n6367  &  wire838  &  wire32384 ) | ( wire838  &  n_n6711  &  wire32384 ) ;
 assign wire4259 = ( n_n6710  &  wire32387 ) | ( n_n6711  &  wire32387 ) | ( wire4973  &  wire32387 ) ;
 assign wire4260 = ( n_n6367  &  wire914  &  wire32388 ) | ( n_n8085  &  wire914  &  wire32388 ) ;
 assign wire4263 = ( (~ pi21)  &  wire424  &  wire32394 ) ;
 assign wire4264 = ( wire4269  &  wire32395 ) | ( wire32189  &  wire32395 ) ;
 assign wire4265 = ( wire4439  &  wire32396 ) | ( wire775  &  wire32341  &  wire32396 ) ;
 assign wire4266 = ( wire1044  &  wire263  &  wire4448 ) | ( wire1044  &  wire263  &  wire4449 ) ;
 assign wire4269 = ( (~ wire150)  &  n_n6710 ) | ( (~ wire150)  &  wire599 ) | ( (~ wire150)  &  wire4973 ) ;
 assign wire4273 = ( wire199  &  wire306 ) | ( wire233  &  wire199  &  n_n7913 ) ;
 assign wire4276 = ( n_n6710  &  wire32227 ) | ( wire4810  &  wire32227 ) | ( wire4811  &  wire32227 ) ;
 assign wire4277 = ( pi20  &  wire153  &  wire306 ) | ( (~ pi20)  &  wire153  &  wire306 ) ;
 assign wire4281 = ( n_n6922  &  (~ wire165) ) | ( (~ wire165)  &  wire4435 ) | ( (~ wire165)  &  wire4436 ) ;
 assign wire4282 = ( wire305  &  wire250 ) | ( wire233  &  wire250  &  n_n7893 ) ;
 assign wire4283 = ( wire305  &  wire243 ) | ( wire233  &  n_n7885  &  wire243 ) ;
 assign wire4284 = ( wire305  &  wire194 ) | ( wire233  &  wire194  &  n_n7877 ) ;
 assign wire4286 = ( (~ ni29)  &  n_n7885  &  wire243 ) | ( (~ n_n8862)  &  n_n7885  &  wire243 ) ;
 assign wire4293 = ( pi27  &  (~ wire150)  &  wire1065 ) | ( (~ pi27)  &  (~ wire150)  &  wire1065 ) | ( (~ pi27)  &  (~ wire150)  &  wire4397 ) ;
 assign wire4294 = ( pi27  &  (~ pi21)  &  wire1065 ) | ( (~ pi27)  &  (~ pi21)  &  wire1065 ) | ( (~ pi27)  &  (~ pi21)  &  wire4397 ) ;
 assign wire4295 = ( pi21  &  pi22  &  n_n6710 ) | ( pi21  &  pi22  &  wire4973 ) ;
 assign wire4296 = ( (~ pi21)  &  ni32  &  (~ ni30) ) ;
 assign wire4299 = ( wire306  &  wire32549 ) | ( wire233  &  n_n7837  &  wire32549 ) ;
 assign wire4300 = ( wire305  &  wire32551 ) | ( wire233  &  n_n7837  &  wire32551 ) ;
 assign wire4301 = ( wire305  &  wire32553 ) | ( wire233  &  n_n7845  &  wire32553 ) ;
 assign wire4302 = ( wire4309  &  wire32554 ) | ( wire4312  &  wire32554 ) | ( wire32233  &  wire32554 ) ;
 assign wire4303 = ( wire4365  &  wire32555 ) | ( pi20  &  n_n6410  &  wire32555 ) ;
 assign wire4305 = ( pi16  &  wire185  &  wire339 ) ;
 assign wire4306 = ( (~ pi23)  &  (~ pi24)  &  wire4317 ) | ( (~ pi23)  &  (~ pi24)  &  wire32264 ) ;
 assign wire4307 = ( wire161  &  wire4322 ) | ( wire161  &  wire4323 ) | ( wire161  &  wire4324 ) ;
 assign wire4309 = ( wire199  &  wire306 ) | ( wire233  &  n_n7845  &  wire199 ) ;
 assign wire4312 = ( n_n6710  &  wire32232 ) | ( wire4784  &  wire32232 ) | ( wire4785  &  wire32232 ) ;
 assign wire4313 = ( pi20  &  wire153  &  wire306 ) | ( (~ pi20)  &  wire153  &  wire306 ) ;
 assign wire4317 = ( (~ ni29)  &  n_n7816  &  wire244 ) | ( (~ n_n8862)  &  n_n7816  &  wire244 ) ;
 assign wire4322 = ( wire305  &  wire251 ) | ( wire233  &  n_n7825  &  wire251 ) ;
 assign wire4323 = ( wire305  &  wire244 ) | ( wire233  &  n_n7816  &  wire244 ) ;
 assign wire4324 = ( wire305  &  wire183 ) | ( wire233  &  wire183  &  n_n7808 ) ;
 assign wire4327 = ( n_n6710  &  wire32349 ) | ( n_n6711  &  wire32349 ) | ( wire4973  &  wire32349 ) ;
 assign wire4331 = ( wire305  &  wire32518 ) | ( wire4544  &  wire32518 ) ;
 assign wire4332 = ( wire204  &  wire4383  &  wire32519 ) | ( wire204  &  wire4384  &  wire32519 ) ;
 assign wire4333 = ( n_n6410  &  wire32522 ) ;
 assign wire4334 = ( wire4349  &  wire32523 ) | ( wire32277  &  wire32523 ) ;
 assign wire4337 = ( pi23  &  wire4341 ) | ( pi24  &  wire4341 ) | ( pi23  &  wire32291 ) | ( pi24  &  wire32291 ) ;
 assign wire4338 = ( (~ wire161)  &  wire4343 ) | ( (~ wire161)  &  wire4344 ) | ( (~ wire161)  &  wire32297 ) ;
 assign wire4341 = ( wire180  &  wire305  &  wire154 ) | ( wire180  &  wire154  &  wire4540 ) ;
 assign wire4342 = ( pi17  &  pi16  &  wire152  &  nv4389 ) ;
 assign wire4343 = ( wire31510  &  wire32292 ) | ( wire31511  &  wire32292 ) | ( wire31512  &  wire32292 ) ;
 assign wire4344 = ( wire31428  &  wire32293 ) | ( wire31429  &  wire32293 ) | ( wire31430  &  wire32293 ) ;
 assign wire4345 = ( wire928  &  wire32294 ) | ( wire4680  &  wire32294 ) | ( wire4681  &  wire32294 ) ;
 assign wire4349 = ( wire31674  &  wire32272 ) | ( wire31675  &  wire32272 ) | ( wire31676  &  wire32272 ) ;
 assign wire4350 = ( n_n6710  &  wire32273 ) | ( wire4781  &  wire32273 ) | ( wire4782  &  wire32273 ) ;
 assign wire4351 = ( n_n6710  &  wire32274 ) | ( wire4787  &  wire32274 ) | ( wire4788  &  wire32274 ) ;
 assign wire4354 = ( wire233  &  wire31756 ) | ( wire233  &  wire31757 ) | ( wire233  &  wire31758 ) ;
 assign wire4357 = ( wire305  &  wire32537 ) | ( wire4564  &  wire32537 ) ;
 assign wire4358 = ( wire4365  &  wire32538 ) | ( pi20  &  n_n6410  &  wire32538 ) ;
 assign wire4359 = ( wire4378  &  wire32539 ) | ( wire32285  &  wire32539 ) ;
 assign wire4361 = ( (~ pi16)  &  wire185  &  wire339 ) ;
 assign wire4362 = ( (~ wire161)  &  wire4367 ) | ( (~ wire161)  &  wire4368 ) | ( (~ wire161)  &  wire32304 ) ;
 assign wire4363 = ( pi23  &  wire4374 ) | ( pi24  &  wire4374 ) | ( pi23  &  wire32306 ) | ( pi24  &  wire32306 ) ;
 assign wire4365 = ( pi21  &  pi20  &  wire4383 ) | ( pi21  &  pi20  &  wire4384 ) ;
 assign wire4367 = ( wire31252  &  wire32299 ) | ( wire31253  &  wire32299 ) | ( wire31254  &  wire32299 ) ;
 assign wire4368 = ( wire31338  &  wire32300 ) | ( wire31339  &  wire32300 ) | ( wire31340  &  wire32300 ) ;
 assign wire4369 = ( wire4613  &  wire32301 ) | ( wire31347  &  wire32301 ) ;
 assign wire4374 = ( wire158  &  wire180  &  wire305 ) | ( wire158  &  wire180  &  wire4574 ) ;
 assign wire4375 = ( pi17  &  (~ pi16)  &  wire152  &  nv4327 ) ;
 assign wire4376 = ( n_n6710  &  wire32280 ) | ( wire4807  &  wire32280 ) | ( wire4808  &  wire32280 ) ;
 assign wire4377 = ( n_n6710  &  wire32281 ) | ( wire4813  &  wire32281 ) | ( wire4814  &  wire32281 ) ;
 assign wire4378 = ( wire31592  &  wire32282 ) | ( wire31593  &  wire32282 ) | ( wire31594  &  wire32282 ) ;
 assign wire4383 = ( (~ pi22)  &  (~ wire161)  &  n_n6367 ) | ( (~ pi22)  &  (~ wire161)  &  n_n6711 ) ;
 assign wire4384 = ( (~ pi22)  &  pi23  &  nv3908 ) | ( (~ pi22)  &  pi24  &  nv3908 ) ;
 assign wire4387 = ( wire233  &  wire31838 ) | ( wire233  &  wire31839 ) | ( wire233  &  wire31840 ) ;
 assign wire4392 = ( n_n6710  &  wire1044 ) | ( wire1044  &  n_n6711 ) | ( wire1044  &  wire4973 ) ;
 assign wire4394 = ( (~ pi22)  &  n_n6367  &  wire32244 ) | ( (~ pi22)  &  n_n6711  &  wire32244 ) ;
 assign wire4397 = ( ni33  &  ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire4400 = ( wire170  &  wire788 ) | ( wire1118  &  wire788 ) ;
 assign wire4406 = ( wire305  &  wire32141 ) | ( wire233  &  n_n7837  &  wire32141 ) ;
 assign wire4407 = ( wire305  &  wire32143 ) | ( wire233  &  n_n7845  &  wire32143 ) ;
 assign wire4409 = ( wire305  &  wire32145 ) | ( wire233  &  n_n7913  &  wire32145 ) ;
 assign wire4410 = ( wire305  &  wire32146 ) | ( wire233  &  n_n7905  &  wire32146 ) ;
 assign wire4411 = ( (~ wire175)  &  wire226  &  wire4504 ) | ( (~ wire175)  &  wire226  &  wire32066 ) ;
 assign wire4415 = ( wire4508  &  wire32151 ) | ( wire4509  &  wire32151 ) | ( wire32074  &  wire32151 ) ;
 assign wire4417 = ( wire369  &  wire4481 ) | ( wire369  &  wire4482 ) | ( wire369  &  wire32079 ) ;
 assign wire4418 = ( wire613  &  wire170 ) | ( wire613  &  wire1118 ) ;
 assign wire4419 = ( (~ wire175)  &  wire4426 ) | ( (~ wire175)  &  wire4430 ) | ( (~ wire175)  &  wire32168 ) ;
 assign wire4421 = ( wire182  &  wire305  &  wire507 ) | ( wire182  &  wire507  &  wire4533 ) ;
 assign wire4422 = ( wire179  &  wire305  &  wire507 ) | ( wire179  &  wire507  &  wire4544 ) ;
 assign wire4423 = ( wire305  &  wire32155 ) | ( wire4564  &  wire32155 ) ;
 assign wire4425 = ( wire305  &  wire32157 ) | ( wire4560  &  wire32157 ) ;
 assign wire4426 = ( (~ pi16)  &  (~ pi15)  &  wire4567 ) | ( (~ pi16)  &  (~ pi15)  &  wire32112 ) ;
 assign wire4428 = ( pi19  &  wire170  &  wire507 ) ;
 assign wire4430 = ( wire614  &  wire4536 ) | ( wire614  &  wire32096 ) ;
 assign wire4432 = ( wire258  &  wire4530 ) | ( wire258  &  wire4531 ) | ( wire258  &  wire4532 ) ;
 assign wire4433 = ( pi27  &  n_n6710 ) | ( pi27  &  n_n8085 ) | ( pi27  &  wire4973 ) ;
 assign wire4434 = ( (~ pi27)  &  wire4973 ) | ( (~ pi27)  &  ni32  &  ni30 ) | ( (~ pi27)  &  ni32  &  (~ ni30) ) ;
 assign wire4435 = ( n_n6367  &  wire32344 ) | ( n_n8085  &  wire32344 ) ;
 assign wire4436 = ( (~ pi27)  &  pi21  &  (~ pi22)  &  nv3908 ) ;
 assign wire4439 = ( (~ pi27)  &  (~ pi21)  &  ni32 ) ;
 assign wire4448 = ( (~ wire156)  &  n_n6710 ) | ( (~ wire156)  &  n_n8085 ) | ( (~ wire156)  &  wire4973 ) ;
 assign wire4449 = ( wire156  &  wire4973 ) | ( ni32  &  ni30  &  wire156 ) | ( ni32  &  (~ ni30)  &  wire156 ) ;
 assign wire4458 = ( (~ wire155)  &  n_n6710 ) | ( (~ wire155)  &  n_n8085 ) | ( (~ wire155)  &  wire4973 ) ;
 assign wire4459 = ( wire155  &  wire4973 ) | ( ni32  &  ni30  &  wire155 ) | ( ni32  &  (~ ni30)  &  wire155 ) ;
 assign wire4462 = ( wire305  &  wire32059 ) | ( wire233  &  n_n7845  &  wire32059 ) ;
 assign wire4464 = ( wire305  &  wire32063 ) | ( wire233  &  n_n7905  &  wire32063 ) ;
 assign wire4465 = ( wire4501  &  wire32068 ) | ( wire4504  &  wire32068 ) | ( wire32066  &  wire32068 ) ;
 assign wire4466 = ( (~ pi20)  &  wire170  &  wire32069 ) | ( (~ pi20)  &  wire4857  &  wire32069 ) ;
 assign wire4467 = ( wire4856  &  wire32070 ) | ( n_n7905  &  wire611  &  wire32070 ) ;
 assign wire4470 = ( wire369  &  wire1113  &  wire449 ) | ( wire369  &  wire1113  &  wire4491 ) ;
 assign wire4471 = ( wire4508  &  wire32076 ) | ( wire4509  &  wire32076 ) | ( wire32074  &  wire32076 ) ;
 assign wire4472 = ( wire4481  &  wire32081 ) | ( wire4482  &  wire32081 ) | ( wire32079  &  wire32081 ) ;
 assign wire4473 = ( wire32026  &  wire32082 ) | ( wire170  &  wire185  &  wire32082 ) ;
 assign wire4474 = ( wire31937  &  wire32083 ) | ( n_n7885  &  wire329  &  wire32083 ) ;
 assign wire4475 = ( wire32018  &  wire32084 ) | ( wire170  &  wire198  &  wire32084 ) ;
 assign wire4476 = ( wire170  &  wire32085 ) | ( n_n9245  &  wire181  &  wire32085 ) ;
 assign wire4478 = ( wire370  &  wire4523 ) | ( wire370  &  wire32103 ) | ( wire370  &  wire32104 ) ;
 assign wire4479 = ( wire370  &  wire4550 ) | ( wire370  &  wire4551 ) | ( wire370  &  wire32118 ) ;
 assign wire4480 = ( wire613  &  wire32053 ) | ( (~ pi15)  &  wire613  &  n_n9255 ) ;
 assign wire4481 = ( wire305  &  wire32077 ) | ( wire233  &  n_n7816  &  wire32077 ) ;
 assign wire4482 = ( wire305  &  wire32078 ) | ( wire233  &  n_n7825  &  wire32078 ) ;
 assign wire4484 = ( wire305  &  wire183 ) | ( wire233  &  wire183  &  n_n7808 ) ;
 assign wire4491 = ( wire305  &  wire199 ) | ( wire233  &  wire199  &  n_n7913 ) ;
 assign wire4501 = ( wire305  &  wire203 ) | ( wire233  &  n_n7837  &  wire203 ) ;
 assign wire4504 = ( n_n6710  &  wire32065 ) | ( wire4784  &  wire32065 ) | ( wire4785  &  wire32065 ) ;
 assign wire4505 = ( pi20  &  wire305  &  wire153 ) | ( (~ pi20)  &  wire305  &  wire153 ) ;
 assign wire4508 = ( wire305  &  wire460 ) | ( wire233  &  n_n7893  &  wire460 ) ;
 assign wire4509 = ( wire305  &  wire329 ) | ( wire233  &  n_n7885  &  wire329 ) ;
 assign wire4510 = ( wire272  &  wire305 ) | ( wire272  &  wire233  &  n_n7877 ) ;
 assign wire4518 = ( wire305  &  wire1053  &  wire32086 ) | ( wire1053  &  wire4544  &  wire32086 ) ;
 assign wire4519 = ( wire31756  &  wire32089 ) | ( wire31757  &  wire32089 ) | ( wire31758  &  wire32089 ) ;
 assign wire4520 = ( (~ pi20)  &  wire170  &  wire32090 ) | ( (~ pi20)  &  wire4857  &  wire32090 ) ;
 assign wire4523 = ( wire4536  &  wire32097 ) | ( wire32096  &  wire32097 ) ;
 assign wire4524 = ( pi16  &  wire4657 ) | ( pi16  &  wire4659 ) | ( pi16  &  wire4660 ) ;
 assign wire4525 = ( pi16  &  wire32018 ) | ( pi16  &  wire170  &  wire198 ) ;
 assign wire4526 = ( pi17  &  pi16  &  wire170 ) | ( pi17  &  pi16  &  wire4857 ) ;
 assign wire4530 = ( n_n6710  &  wire32091 ) | ( wire4781  &  wire32091 ) | ( wire4782  &  wire32091 ) ;
 assign wire4531 = ( n_n6710  &  wire32092 ) | ( wire4787  &  wire32092 ) | ( wire4788  &  wire32092 ) ;
 assign wire4532 = ( pi20  &  wire305  &  wire153 ) | ( (~ pi20)  &  wire305  &  wire153 ) ;
 assign wire4533 = ( wire233  &  wire31674 ) | ( wire233  &  wire31675 ) | ( wire233  &  wire31676 ) ;
 assign wire4536 = ( wire178  &  wire305 ) | ( wire178  &  wire4538 ) ;
 assign wire4538 = ( wire233  &  wire31510 ) | ( wire233  &  wire31511 ) | ( wire233  &  wire31512 ) ;
 assign wire4540 = ( wire233  &  wire31428 ) | ( wire233  &  wire31429 ) | ( wire233  &  wire31430 ) ;
 assign wire4544 = ( wire233  &  wire31756 ) | ( wire233  &  wire31757 ) | ( wire233  &  wire31758 ) ;
 assign wire4546 = ( wire31838  &  wire32106 ) | ( wire31839  &  wire32106 ) | ( wire31840  &  wire32106 ) ;
 assign wire4547 = ( wire31592  &  wire32107 ) | ( wire31593  &  wire32107 ) | ( wire31594  &  wire32107 ) ;
 assign wire4548 = ( wire305  &  wire1028  &  wire698 ) | ( wire1028  &  wire698  &  wire4564 ) ;
 assign wire4550 = ( (~ pi25)  &  (~ pi16)  &  wire505 ) ;
 assign wire4551 = ( (~ pi25)  &  (~ pi16)  &  wire4567 ) | ( (~ pi25)  &  (~ pi16)  &  wire32112 ) ;
 assign wire4553 = ( wire705  &  wire4608 ) | ( wire705  &  wire4609 ) | ( wire705  &  wire31960 ) ;
 assign wire4554 = ( (~ pi16)  &  wire32026 ) | ( (~ pi16)  &  wire170  &  wire185 ) ;
 assign wire4556 = ( pi20  &  wire305  &  wire153 ) | ( pi20  &  wire153  &  wire4560 ) ;
 assign wire4558 = ( n_n6710  &  wire233 ) | ( wire233  &  wire4807 ) | ( wire233  &  wire4808 ) ;
 assign wire4560 = ( n_n6710  &  wire233 ) | ( wire233  &  wire4813 ) | ( wire233  &  wire4814 ) ;
 assign wire4562 = ( wire233  &  wire31592 ) | ( wire233  &  wire31593 ) | ( wire233  &  wire31594 ) ;
 assign wire4564 = ( wire233  &  wire31838 ) | ( wire233  &  wire31839 ) | ( wire233  &  wire31840 ) ;
 assign wire4567 = ( pi17  &  wire180  &  wire305 ) | ( pi17  &  wire180  &  wire4574 ) ;
 assign wire4570 = ( wire233  &  wire31252 ) | ( wire233  &  wire31253 ) | ( wire233  &  wire31254 ) ;
 assign wire4574 = ( wire233  &  wire31338 ) | ( wire233  &  wire31339 ) | ( wire233  &  wire31340 ) ;
 assign wire4581 = ( ni32  &  (~ ni30)  &  ni29 ) ;
 assign wire4583 = ( wire31592  &  wire32001 ) | ( wire31593  &  wire32001 ) | ( wire31594  &  wire32001 ) ;
 assign wire4585 = ( wire31838  &  wire32005 ) | ( wire31839  &  wire32005 ) | ( wire31840  &  wire32005 ) ;
 assign wire4588 = ( wire1288  &  wire32010 ) | ( n_n8890  &  wire213  &  wire32010 ) ;
 assign wire4589 = ( wire1288  &  wire32011 ) | ( n_n8890  &  wire213  &  wire32011 ) ;
 assign wire4590 = ( wire4856  &  wire32012 ) | ( n_n7905  &  wire611  &  wire32012 ) ;
 assign wire4591 = ( wire4608  &  wire32014 ) | ( wire4609  &  wire32014 ) | ( wire31960  &  wire32014 ) ;
 assign wire4592 = ( pi15  &  wire904  &  wire4875 ) | ( pi15  &  wire904  &  wire31937 ) ;
 assign wire4596 = ( wire32026  &  wire32027 ) | ( wire170  &  wire185  &  wire32027 ) ;
 assign wire4599 = ( wire403  &  wire279 ) | ( wire403  &  (~ wire150)  &  n_n8890 ) ;
 assign wire4606 = ( n_n6710  &  wire247 ) | ( wire247  &  wire4813 ) | ( wire247  &  wire4814 ) ;
 assign wire4607 = ( n_n6710  &  wire219 ) | ( wire219  &  wire4807 ) | ( wire219  &  wire4808 ) ;
 assign wire4608 = ( wire460  &  wire31252 ) | ( wire460  &  wire31253 ) | ( wire460  &  wire31254 ) ;
 assign wire4609 = ( wire329  &  wire31338 ) | ( wire329  &  wire31339 ) | ( wire329  &  wire31340 ) ;
 assign wire4613 = ( (~ wire323)  &  (~ wire4917)  &  wire31346 ) ;
 assign wire4615 = ( (~ wire1103)  &  (~ wire4896)  &  (~ wire4897)  &  wire31266 ) ;
 assign wire4620 = ( (~ wire4899)  &  (~ wire4900)  &  (~ wire4901)  &  wire31286 ) ;
 assign wire4624 = ( (~ wire4899)  &  (~ wire4900)  &  (~ wire4901)  &  wire31302 ) ;
 assign wire4625 = ( (~ wire1103)  &  (~ wire4896)  &  (~ wire4897)  &  wire31306 ) ;
 assign wire4627 = ( (~ n_n8948)  &  (~ wire1103)  &  (~ wire4896)  &  wire31313 ) ;
 assign wire4632 = ( (~ wire1103)  &  (~ wire4886)  &  (~ wire4887)  &  wire31180 ) ;
 assign wire4638 = ( (~ wire4889)  &  (~ wire4890)  &  (~ wire4891)  &  wire31204 ) ;
 assign wire4641 = ( (~ wire1103)  &  (~ wire4886)  &  (~ wire4887)  &  wire31216 ) ;
 assign wire4642 = ( (~ wire4889)  &  (~ wire4890)  &  (~ wire4891)  &  wire31220 ) ;
 assign wire4644 = ( (~ wire1103)  &  (~ n_n8956)  &  (~ wire4886)  &  wire31227 ) ;
 assign wire4649 = ( ni41  &  wire346  &  nv3916 ) | ( (~ ni41)  &  wire346  &  nv3918 ) ;
 assign wire4651 = ( wire31756  &  wire32029 ) | ( wire31757  &  wire32029 ) | ( wire31758  &  wire32029 ) ;
 assign wire4652 = ( wire1288  &  wire32030 ) | ( n_n8890  &  wire213  &  wire32030 ) ;
 assign wire4653 = ( pi16  &  wire4657 ) | ( pi16  &  wire4659 ) | ( pi16  &  wire4660 ) ;
 assign wire4655 = ( wire154  &  wire279 ) | ( (~ wire150)  &  n_n8890  &  wire154 ) ;
 assign wire4657 = ( wire437  &  wire31674 ) | ( wire437  &  wire31675 ) | ( wire437  &  wire31676 ) ;
 assign wire4659 = ( n_n6710  &  wire247 ) | ( wire247  &  wire4787 ) | ( wire247  &  wire4788 ) ;
 assign wire4660 = ( n_n6710  &  wire219 ) | ( wire219  &  wire4781 ) | ( wire219  &  wire4782 ) ;
 assign wire4661 = ( (~ wire1098)  &  (~ wire4792)  &  (~ wire4793)  &  wire31602 ) ;
 assign wire4663 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31610 ) ;
 assign wire4667 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31626 ) ;
 assign wire4668 = ( (~ wire254)  &  (~ wire4799)  &  wire31630 ) | ( (~ nv4058)  &  (~ wire4799)  &  wire31630 ) ;
 assign wire4671 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31642 ) ;
 assign wire4674 = ( (~ wire1098)  &  (~ wire4792)  &  (~ wire4793)  &  wire31654 ) ;
 assign wire4675 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31658 ) ;
 assign wire4676 = ( (~ wire253)  &  (~ nv4058)  &  wire31661 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31661 ) ;
 assign wire4678 = ( wire476  &  wire1178 ) | ( wire476  &  wire4687 ) | ( wire476  &  wire4688 ) ;
 assign wire4680 = ( (~ wire205)  &  wire206  &  (~ nv3918) ) | ( wire206  &  (~ nv3918)  &  wire4685 ) ;
 assign wire4681 = ( (~ wire323)  &  (~ wire4824)  &  wire31851 ) ;
 assign wire4685 = ( ni38  &  ni36 ) | ( ni47  &  (~ ni45)  &  ni36 ) ;
 assign wire4687 = ( wire180  &  wire31428 ) | ( wire180  &  wire31429 ) | ( wire180  &  wire31430 ) ;
 assign wire4688 = ( wire178  &  wire31510 ) | ( wire178  &  wire31511 ) | ( wire178  &  wire31512 ) ;
 assign wire4690 = ( (~ wire1103)  &  (~ wire4843)  &  (~ wire4844)  &  wire31356 ) ;
 assign wire4691 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31360 ) ;
 assign wire4695 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31376 ) ;
 assign wire4697 = ( (~ wire253)  &  (~ wire4851)  &  wire31384 ) | ( (~ nv4058)  &  (~ wire4851)  &  wire31384 ) ;
 assign wire4699 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31392 ) ;
 assign wire4703 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31408 ) ;
 assign wire4704 = ( (~ wire1103)  &  (~ wire4843)  &  (~ wire4844)  &  wire31412 ) ;
 assign wire4705 = ( (~ wire254)  &  (~ nv4058)  &  wire31415 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31415 ) ;
 assign wire4707 = ( (~ wire1103)  &  (~ wire4833)  &  (~ wire4834)  &  wire31438 ) ;
 assign wire4709 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31446 ) ;
 assign wire4713 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31462 ) ;
 assign wire4714 = ( (~ wire253)  &  (~ wire4839)  &  wire31466 ) | ( (~ nv4045)  &  (~ wire4839)  &  wire31466 ) ;
 assign wire4717 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31478 ) ;
 assign wire4720 = ( (~ wire1103)  &  (~ wire4833)  &  (~ wire4834)  &  wire31490 ) ;
 assign wire4721 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31494 ) ;
 assign wire4722 = ( (~ wire254)  &  (~ nv4045)  &  wire31497 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31497 ) ;
 assign wire4738 = ( (~ wire1098)  &  (~ wire4921)  &  (~ wire4922)  &  wire31684 ) ;
 assign wire4739 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31688 ) ;
 assign wire4743 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31704 ) ;
 assign wire4745 = ( (~ wire254)  &  (~ wire4930)  &  wire31712 ) | ( (~ nv4045)  &  (~ wire4930)  &  wire31712 ) ;
 assign wire4747 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31720 ) ;
 assign wire4751 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31736 ) ;
 assign wire4752 = ( (~ wire1098)  &  (~ wire4921)  &  (~ wire4922)  &  wire31740 ) ;
 assign wire4753 = ( (~ wire253)  &  (~ nv4045)  &  wire31743 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31743 ) ;
 assign wire4757 = ( (~ wire1098)  &  (~ wire4861)  &  (~ wire4862)  &  wire31766 ) ;
 assign wire4763 = ( (~ wire4864)  &  (~ wire4865)  &  (~ wire4866)  &  wire31790 ) ;
 assign wire4766 = ( (~ wire1098)  &  (~ wire4861)  &  (~ wire4862)  &  wire31802 ) ;
 assign wire4767 = ( (~ wire4864)  &  (~ wire4865)  &  (~ wire4866)  &  wire31806 ) ;
 assign wire4769 = ( (~ wire1098)  &  (~ n_n8968)  &  (~ wire4861)  &  wire31813 ) ;
 assign wire4776 = ( n_n6710  &  wire247 ) | ( wire247  &  wire4784 ) | ( wire247  &  wire4785 ) ;
 assign wire4778 = ( (~ wire400)  &  wire1041  &  (~ wire871) ) | ( (~ nv4045)  &  wire1041  &  (~ wire871) ) ;
 assign wire4779 = ( n_n6710  &  wire632 ) | ( wire632  &  wire4781 ) | ( wire632  &  wire4782 ) ;
 assign wire4781 = ( wire206  &  (~ nv4045)  &  wire255  &  (~ wire871) ) ;
 assign wire4782 = ( (~ wire400)  &  wire1007  &  (~ wire871) ) | ( (~ nv4045)  &  wire1007  &  (~ wire871) ) ;
 assign wire4784 = ( (~ wire365)  &  (~ wire870)  &  wire1041 ) | ( (~ nv4058)  &  (~ wire870)  &  wire1041 ) ;
 assign wire4785 = ( n_n6710  &  wire632 ) | ( wire632  &  wire4787 ) | ( wire632  &  wire4788 ) ;
 assign wire4787 = ( wire206  &  (~ nv4058)  &  (~ wire870)  &  wire255 ) ;
 assign wire4788 = ( (~ wire365)  &  (~ wire870)  &  wire1007 ) | ( (~ nv4058)  &  (~ wire870)  &  wire1007 ) ;
 assign wire4792 = ( wire176  &  wire4799 ) | ( wire176  &  wire254  &  nv4058 ) ;
 assign wire4793 = ( ni35  &  wire4795 ) | ( ni35  &  wire4796 ) | ( ni35  &  wire4797 ) ;
 assign wire4795 = ( wire870  &  wire989 ) | ( wire365  &  nv4058  &  wire989 ) ;
 assign wire4796 = ( ni45  &  wire847 ) | ( ni43  &  (~ ni47)  &  wire847 ) ;
 assign wire4797 = ( (~ ni36)  &  wire4799 ) | ( (~ ni36)  &  wire254  &  nv4058 ) ;
 assign wire4799 = ( (~ ni40)  &  ni38  &  nv3918 ) ;
 assign wire4802 = ( n_n6710  &  wire247 ) | ( wire247  &  wire4810 ) | ( wire247  &  wire4811 ) ;
 assign wire4803 = ( n_n6710  &  wire219 ) | ( wire219  &  wire4804 ) | ( wire219  &  wire4805 ) ;
 assign wire4804 = ( (~ wire400)  &  wire1041  &  (~ wire871) ) | ( (~ nv3927)  &  wire1041  &  (~ wire871) ) ;
 assign wire4805 = ( n_n6710  &  wire632 ) | ( wire632  &  wire4807 ) | ( wire632  &  wire4808 ) ;
 assign wire4807 = ( wire206  &  (~ nv3927)  &  wire255  &  (~ wire871) ) ;
 assign wire4808 = ( (~ wire400)  &  wire1007  &  (~ wire871) ) | ( (~ nv3927)  &  wire1007  &  (~ wire871) ) ;
 assign wire4810 = ( (~ wire365)  &  (~ wire870)  &  wire1041 ) | ( (~ nv3943)  &  (~ wire870)  &  wire1041 ) ;
 assign wire4811 = ( n_n6710  &  wire632 ) | ( wire632  &  wire4813 ) | ( wire632  &  wire4814 ) ;
 assign wire4813 = ( wire206  &  (~ nv3943)  &  (~ wire870)  &  wire255 ) ;
 assign wire4814 = ( (~ wire365)  &  (~ wire870)  &  wire1007 ) | ( (~ nv3943)  &  (~ wire870)  &  wire1007 ) ;
 assign wire4817 = ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire4824 = ( ni45  &  ni38 ) | ( ni43  &  (~ ni47)  &  ni38 ) ;
 assign wire4827 = ( wire178  &  n_n7825 ) ;
 assign wire4833 = ( wire177  &  wire4839 ) | ( wire177  &  wire253  &  nv4045 ) ;
 assign wire4834 = ( (~ ni35)  &  wire4836 ) | ( (~ ni35)  &  wire4837 ) | ( (~ ni35)  &  wire4838 ) ;
 assign wire4836 = ( wire991  &  wire871 ) | ( wire400  &  nv4045  &  wire991 ) ;
 assign wire4837 = ( ni45  &  wire814 ) | ( ni43  &  (~ ni47)  &  wire814 ) ;
 assign wire4838 = ( (~ ni36)  &  wire4839 ) | ( (~ ni36)  &  wire253  &  nv4045 ) ;
 assign wire4839 = ( ni40  &  ni38  &  nv3918 ) ;
 assign wire4843 = ( wire177  &  wire4851 ) | ( wire177  &  wire253  &  nv4058 ) ;
 assign wire4844 = ( (~ ni35)  &  wire4846 ) | ( (~ ni35)  &  wire4847 ) | ( (~ ni35)  &  wire4848 ) ;
 assign wire4846 = ( wire870  &  wire990 ) | ( wire365  &  nv4058  &  wire990 ) ;
 assign wire4847 = ( ni45  &  wire840 ) | ( ni43  &  (~ ni47)  &  wire840 ) ;
 assign wire4848 = ( (~ ni36)  &  wire4851 ) | ( (~ ni36)  &  wire253  &  nv4058 ) ;
 assign wire4851 = ( ni40  &  ni38  &  nv3918 ) ;
 assign wire4853 = ( ni41  &  ni45 ) | ( ni43  &  ni41  &  (~ ni47) ) ;
 assign wire4856 = ( pi20  &  wire170 ) | ( pi20  &  n_n9245  &  wire181 ) ;
 assign wire4857 = ( ni32  &  ni30  &  wire181 ) ;
 assign wire4861 = ( wire176  &  wire4868 ) | ( wire176  &  wire254  &  nv3943 ) ;
 assign wire4862 = ( ni35  &  wire4864 ) | ( ni35  &  wire4865 ) | ( ni35  &  wire4866 ) ;
 assign wire4864 = ( wire870  &  wire989 ) | ( wire365  &  nv3943  &  wire989 ) ;
 assign wire4865 = ( ni41  &  wire847  &  nv3916 ) | ( (~ ni41)  &  wire847  &  nv3918 ) ;
 assign wire4866 = ( (~ ni36)  &  wire4868 ) | ( (~ ni36)  &  wire254  &  nv3943 ) ;
 assign wire4868 = ( ni41  &  wire253  &  nv3916 ) | ( (~ ni41)  &  wire253  &  nv3918 ) ;
 assign wire4875 = ( pi17  &  wire180  &  n_n7885 ) ;
 assign wire4886 = ( wire177  &  wire4892 ) | ( wire177  &  wire253  &  nv3927 ) ;
 assign wire4887 = ( (~ ni35)  &  wire4889 ) | ( (~ ni35)  &  wire4890 ) | ( (~ ni35)  &  wire4891 ) ;
 assign wire4889 = ( wire991  &  wire871 ) | ( wire400  &  nv3927  &  wire991 ) ;
 assign wire4890 = ( ni41  &  wire814  &  nv3916 ) | ( (~ ni41)  &  wire814  &  nv3918 ) ;
 assign wire4891 = ( (~ ni36)  &  wire4892 ) | ( (~ ni36)  &  wire253  &  nv3927 ) ;
 assign wire4892 = ( ni41  &  wire254  &  nv3916 ) | ( (~ ni41)  &  wire254  &  nv3918 ) ;
 assign wire4896 = ( wire177  &  wire4904 ) | ( wire177  &  wire253  &  nv3943 ) ;
 assign wire4897 = ( (~ ni35)  &  wire4899 ) | ( (~ ni35)  &  wire4900 ) | ( (~ ni35)  &  wire4901 ) ;
 assign wire4899 = ( wire870  &  wire990 ) | ( wire365  &  nv3943  &  wire990 ) ;
 assign wire4900 = ( ni41  &  wire840  &  nv3916 ) | ( (~ ni41)  &  wire840  &  nv3918 ) ;
 assign wire4901 = ( (~ ni36)  &  wire4904 ) | ( (~ ni36)  &  wire253  &  nv3943 ) ;
 assign wire4904 = ( ni41  &  wire254  &  nv3916 ) | ( (~ ni41)  &  wire254  &  nv3918 ) ;
 assign wire4910 = ( wire4913  &  wire31258 ) | ( (~ ni41)  &  ni44  &  wire31258 ) ;
 assign wire4911 = ( ni42  &  wire1281 ) ;
 assign wire4912 = ( nv3916  &  wire4913 ) | ( (~ ni41)  &  ni44  &  nv3916 ) ;
 assign wire4913 = ( ni43  &  (~ ni41) ) | ( ni42  &  (~ ni41) ) | ( (~ ni41)  &  ni45 ) ;
 assign wire4917 = ( ni41  &  ni38  &  nv3916 ) | ( (~ ni41)  &  ni38  &  nv3918 ) ;
 assign wire4921 = ( wire176  &  wire4930 ) | ( wire176  &  wire254  &  nv4045 ) ;
 assign wire4922 = ( ni35  &  wire4924 ) | ( ni35  &  wire4925 ) | ( ni35  &  wire4926 ) ;
 assign wire4924 = ( wire992  &  wire871 ) | ( wire400  &  nv4045  &  wire992 ) ;
 assign wire4925 = ( ni45  &  wire834 ) | ( ni43  &  (~ ni47)  &  wire834 ) ;
 assign wire4926 = ( (~ ni36)  &  wire4930 ) | ( (~ ni36)  &  wire254  &  nv4045 ) ;
 assign wire4930 = ( (~ ni40)  &  ni38  &  nv3918 ) ;
 assign wire4931 = ( ni41  &  ni45 ) | ( ni43  &  ni41  &  (~ ni47) ) ;
 assign wire4933 = ( (~ wire1098)  &  (~ wire4952)  &  (~ wire4953)  &  wire31520 ) ;
 assign wire4938 = ( (~ wire4957)  &  (~ wire4958)  &  (~ wire4959)  &  wire31540 ) ;
 assign wire4942 = ( (~ wire4957)  &  (~ wire4958)  &  (~ wire4959)  &  wire31556 ) ;
 assign wire4943 = ( (~ wire1098)  &  (~ wire4952)  &  (~ wire4953)  &  wire31560 ) ;
 assign wire4945 = ( (~ n_n8976)  &  (~ wire1098)  &  (~ wire4952)  &  wire31567 ) ;
 assign wire4950 = ( ni41  &  wire347  &  nv3916 ) | ( (~ ni41)  &  wire347  &  nv3918 ) ;
 assign wire4952 = ( wire176  &  wire4967 ) | ( wire176  &  wire254  &  nv3927 ) ;
 assign wire4953 = ( ni35  &  wire4957 ) | ( ni35  &  wire4958 ) | ( ni35  &  wire4959 ) ;
 assign wire4957 = ( wire992  &  wire871 ) | ( wire400  &  nv3927  &  wire992 ) ;
 assign wire4958 = ( ni41  &  nv3916  &  wire834 ) | ( (~ ni41)  &  nv3918  &  wire834 ) ;
 assign wire4959 = ( (~ ni36)  &  wire4967 ) | ( (~ ni36)  &  wire254  &  nv3927 ) ;
 assign wire4967 = ( ni41  &  wire253  &  nv3916 ) | ( (~ ni41)  &  wire253  &  nv3918 ) ;
 assign wire4968 = ( wire4971  &  wire31173 ) | ( (~ ni41)  &  (~ ni44)  &  wire31173 ) ;
 assign wire4969 = ( ni42  &  wire1281 ) ;
 assign wire4970 = ( nv3916  &  wire4971 ) | ( (~ ni41)  &  (~ ni44)  &  nv3916 ) ;
 assign wire4971 = ( ni43  &  (~ ni41) ) | ( ni42  &  (~ ni41) ) | ( (~ ni41)  &  ni45 ) ;
 assign wire4973 = ( (~ wire172)  &  wire206  &  wire255 ) | ( wire206  &  (~ nv3916)  &  wire255 ) ;
 assign wire4981 = ( ni2  &  ni10 ) | ( ni3  &  ni10 ) ;
 assign wire4991 = ( nv10727  &  wire30389 ) | ( wire237  &  wire30389 ) | ( wire5829  &  wire30389 ) ;
 assign wire4995 = ( nv10727  &  wire30414 ) | ( wire237  &  wire30414 ) | ( wire5875  &  wire30414 ) ;
 assign wire4997 = ( n_n9587  &  wire30430 ) ;
 assign wire4999 = ( wire30452  &  wire30455 ) | ( wire252  &  wire852  &  wire30455 ) ;
 assign wire5000 = ( wire5086  &  wire30458 ) | ( wire5087  &  wire30458 ) ;
 assign wire5002 = ( nv3377  &  wire416  &  wire30463 ) ;
 assign wire5003 = ( wire5071  &  wire30493 ) | ( wire5073  &  wire30493 ) | ( wire30489  &  wire30493 ) ;
 assign wire5006 = ( wire5063  &  wire30754 ) | ( wire30704  &  wire30754 ) | ( wire30752  &  wire30754 ) ;
 assign wire5009 = ( wire31139  &  wire31140 ) | ( wire708  &  n_n9515  &  wire31140 ) ;
 assign wire5010 = ( ni2  &  ni33 ) | ( ni3  &  ni33 ) ;
 assign wire5011 = ( wire180  &  wire240  &  wire30705 ) | ( wire180  &  wire5906  &  wire30705 ) ;
 assign wire5012 = ( wire240  &  wire30708 ) | ( ni33  &  nv2493  &  wire30708 ) ;
 assign wire5013 = ( wire180  &  wire240  &  wire30709 ) | ( wire180  &  wire5845  &  wire30709 ) ;
 assign wire5014 = ( wire240  &  wire30712 ) | ( ni33  &  nv2565  &  wire30712 ) ;
 assign wire5015 = ( wire240  &  wire30713 ) | ( ni33  &  nv2314  &  wire30713 ) ;
 assign wire5017 = ( wire240  &  wire30715 ) | ( wire5770  &  wire30715 ) ;
 assign wire5018 = ( wire5788  &  wire30716 ) | ( wire30425  &  wire30716 ) ;
 assign wire5019 = ( wire240  &  wire30717 ) | ( wire5861  &  wire30717 ) ;
 assign wire5022 = ( wire240  &  wire30720 ) | ( wire5871  &  wire30720 ) ;
 assign wire5024 = ( pi15  &  (~ ni14)  &  wire5086 ) | ( pi15  &  (~ ni14)  &  wire5087 ) ;
 assign wire5025 = ( (~ pi15)  &  (~ ni14)  &  wire5033 ) | ( (~ pi15)  &  (~ ni14)  &  wire30728 ) ;
 assign wire5026 = ( (~ pi15)  &  (~ ni14)  &  wire5039 ) | ( (~ pi15)  &  (~ ni14)  &  wire30737 ) ;
 assign wire5029 = ( wire240  &  wire30722 ) | ( ni33  &  nv2276  &  wire30722 ) ;
 assign wire5030 = ( wire158  &  wire240  &  wire324 ) | ( wire158  &  wire324  &  wire5196 ) ;
 assign wire5032 = ( wire325  &  wire240 ) | ( ni33  &  wire325  &  nv2197 ) ;
 assign wire5033 = ( (~ pi17)  &  (~ pi16)  &  wire5184 ) | ( (~ pi17)  &  (~ pi16)  &  wire30509 ) ;
 assign wire5034 = ( wire294  &  wire240 ) | ( ni33  &  wire294  &  nv2220 ) ;
 assign wire5037 = ( wire240  &  wire30730 ) | ( ni33  &  nv2397  &  wire30730 ) ;
 assign wire5039 = ( (~ pi17)  &  pi16  &  wire5125 ) | ( (~ pi17)  &  pi16  &  wire30731 ) ;
 assign wire5040 = ( wire240  &  wire1024 ) | ( ni33  &  nv2330  &  wire1024 ) ;
 assign wire5044 = ( wire5325  &  wire30527 ) | ( wire30525  &  wire30527 ) ;
 assign wire5045 = ( wire30530  &  wire30532 ) | ( wire238  &  nv3060  &  wire30532 ) ;
 assign wire5046 = ( wire307  &  wire30537 ) | ( wire5278  &  wire30537 ) | ( wire5279  &  wire30537 ) ;
 assign wire5047 = ( wire5337  &  wire30542 ) | ( wire30540  &  wire30542 ) ;
 assign wire5048 = ( wire5319  &  wire30557 ) | ( wire30553  &  wire30557 ) | ( wire30554  &  wire30557 ) ;
 assign wire5049 = ( wire30560  &  wire30562 ) | ( nv2946  &  wire238  &  wire30562 ) ;
 assign wire5050 = ( wire5329  &  wire30577 ) | ( wire30573  &  wire30577 ) | ( wire30574  &  wire30577 ) ;
 assign wire5051 = ( wire5426  &  wire30580 ) | ( wire30579  &  wire30580 ) ;
 assign wire5052 = ( wire5361  &  wire30600 ) | ( wire5362  &  wire30600 ) | ( wire30598  &  wire30600 ) ;
 assign wire5055 = ( wire5396  &  wire30624 ) | ( wire5397  &  wire30624 ) | ( wire30622  &  wire30624 ) ;
 assign wire5056 = ( pi15  &  ni14  &  wire5086 ) | ( pi15  &  ni14  &  wire5087 ) ;
 assign wire5058 = ( wire307  &  wire30628 ) | ( wire5291  &  wire30628 ) | ( wire5292  &  wire30628 ) ;
 assign wire5059 = ( wire5286  &  wire30638 ) | ( wire5287  &  wire30638 ) | ( wire30636  &  wire30638 ) ;
 assign wire5060 = ( wire5273  &  wire30648 ) | ( wire5274  &  wire30648 ) | ( wire30646  &  wire30648 ) ;
 assign wire5063 = ( wire1069  &  wire5066 ) | ( wire1069  &  wire5068 ) | ( wire1069  &  wire30685 ) ;
 assign wire5064 = ( wire158  &  wire324  &  wire5487 ) | ( wire158  &  wire324  &  wire30650 ) ;
 assign wire5065 = ( wire325  &  wire30651 ) | ( wire325  &  nv2197  &  wire315 ) ;
 assign wire5066 = ( wire302  &  wire5463 ) | ( wire302  &  wire30664 ) | ( wire302  &  wire30665 ) ;
 assign wire5068 = ( wire158  &  wire5494 ) | ( wire158  &  wire30680 ) | ( wire158  &  wire30681 ) ;
 assign wire5070 = ( wire304  &  wire30468 ) | ( wire252  &  nv2411  &  wire30468 ) ;
 assign wire5071 = ( wire304  &  wire30472 ) | ( wire5223  &  wire30472 ) | ( wire5902  &  wire30472 ) ;
 assign wire5072 = ( wire304  &  wire1309 ) | ( wire252  &  wire1309  &  nv2430 ) ;
 assign wire5073 = ( (~ pi17)  &  pi16  &  wire5198 ) | ( (~ pi17)  &  pi16  &  wire30484 ) ;
 assign wire5075 = ( wire751  &  wire763 ) | ( (~ n_n12619)  &  nv2340  &  wire763 ) ;
 assign wire5078 = ( wire304  &  wire30497 ) | ( wire252  &  nv2290  &  wire30497 ) ;
 assign wire5079 = ( nv10727  &  wire30501 ) | ( wire237  &  wire30501 ) | ( wire5215  &  wire30501 ) ;
 assign wire5080 = ( pi17  &  (~ pi16)  &  wire324  &  nv3202 ) ;
 assign wire5082 = ( nv10727  &  wire325 ) | ( wire325  &  wire237 ) | ( wire325  &  wire5219 ) ;
 assign wire5086 = ( pi20  &  wire344  &  wire162 ) | ( (~ pi20)  &  wire344  &  wire159 ) ;
 assign wire5087 = ( pi20  &  wire295  &  wire162 ) | ( (~ pi20)  &  wire295  &  wire159 ) ;
 assign wire5088 = ( wire5788  &  wire30758 ) | ( wire30425  &  wire30758 ) ;
 assign wire5089 = ( wire240  &  wire30762 ) | ( ni33  &  nv2565  &  wire30762 ) ;
 assign wire5090 = ( wire240  &  wire247  &  wire30765 ) | ( wire247  &  wire5861  &  wire30765 ) ;
 assign wire5091 = ( wire240  &  wire30770 ) | ( ni33  &  nv2493  &  wire30770 ) ;
 assign wire5092 = ( wire240  &  wire219  &  wire30773 ) | ( wire219  &  wire5770  &  wire30773 ) ;
 assign wire5094 = ( wire916  &  wire30781 ) | ( wire5249  &  wire30781 ) ;
 assign wire5095 = ( wire916  &  wire30784 ) | ( wire5249  &  wire30784 ) ;
 assign wire5096 = ( wire240  &  wire813  &  wire30786 ) | ( wire813  &  wire5845  &  wire30786 ) ;
 assign wire5097 = ( wire240  &  wire812  &  wire30789 ) | ( wire812  &  wire5906  &  wire30789 ) ;
 assign wire5098 = ( wire240  &  wire30793 ) | ( ni33  &  nv2314  &  wire30793 ) ;
 assign wire5099 = ( wire240  &  wire311  &  wire30795 ) | ( wire311  &  wire5871  &  wire30795 ) ;
 assign wire5101 = ( wire5239  &  wire30826 ) | ( wire5240  &  wire30826 ) | ( wire5241  &  wire30826 ) ;
 assign wire5102 = ( wire5242  &  wire30828 ) | ( wire5243  &  wire30828 ) | ( wire5244  &  wire30828 ) ;
 assign wire5103 = ( wire263  &  wire5247  &  wire30829 ) | ( wire263  &  wire5248  &  wire30829 ) ;
 assign wire5107 = ( wire5125  &  wire30800 ) | ( wire30731  &  wire30800 ) ;
 assign wire5108 = ( wire5184  &  wire30801 ) | ( wire30509  &  wire30801 ) ;
 assign wire5109 = ( wire240  &  wire30802 ) | ( ni33  &  nv2397  &  wire30802 ) ;
 assign wire5110 = ( wire240  &  wire30803 ) | ( ni33  &  nv2220  &  wire30803 ) ;
 assign wire5111 = ( wire240  &  wire30804 ) | ( ni33  &  nv2330  &  wire30804 ) ;
 assign wire5112 = ( wire240  &  wire30805 ) | ( ni33  &  nv2197  &  wire30805 ) ;
 assign wire5113 = ( nv2340  &  wire30806 ) ;
 assign wire5114 = ( wire240  &  wire30807 ) | ( ni33  &  nv2276  &  wire30807 ) ;
 assign wire5115 = ( wire593  &  wire916 ) | ( wire593  &  wire5249 ) ;
 assign wire5116 = ( wire456  &  wire916 ) | ( wire456  &  wire5249 ) ;
 assign wire5119 = ( wire240  &  wire393 ) | ( wire393  &  wire5196 ) ;
 assign wire5120 = ( pi25  &  wire152  &  wire154  &  nv2430 ) ;
 assign wire5125 = ( wire240  &  wire179 ) | ( ni33  &  wire179  &  nv2359 ) ;
 assign wire5128 = ( nv10727  &  wire30834 ) | ( wire237  &  wire30834 ) | ( wire5211  &  wire30834 ) ;
 assign wire5130 = ( nv10727  &  wire30838 ) | ( wire237  &  wire30838 ) | ( wire5219  &  wire30838 ) ;
 assign wire5131 = ( wire304  &  wire30840 ) | ( wire5223  &  wire30840 ) | ( wire5902  &  wire30840 ) ;
 assign wire5132 = ( nv10727  &  wire30841 ) | ( wire237  &  wire30841 ) | ( wire5190  &  wire30841 ) ;
 assign wire5134 = ( wire5198  &  wire30843 ) | ( wire30484  &  wire30843 ) ;
 assign wire5135 = ( wire304  &  wire30844 ) | ( wire252  &  nv2290  &  wire30844 ) ;
 assign wire5138 = ( wire304  &  wire30847 ) | ( wire252  &  nv2411  &  wire30847 ) ;
 assign wire5139 = ( wire751  &  wire30848 ) | ( (~ n_n12619)  &  nv2340  &  wire30848 ) ;
 assign wire5140 = ( wire304  &  wire30849 ) | ( wire252  &  nv2430  &  wire30849 ) ;
 assign wire5142 = ( (~ pi15)  &  wire5239 ) | ( (~ pi15)  &  wire5240 ) | ( (~ pi15)  &  wire5241 ) ;
 assign wire5143 = ( (~ pi15)  &  wire5242 ) | ( (~ pi15)  &  wire5243 ) | ( (~ pi15)  &  wire5244 ) ;
 assign wire5144 = ( (~ pi15)  &  wire5247 ) | ( (~ pi15)  &  wire5248 ) ;
 assign wire5145 = ( wire30452  &  wire30850 ) | ( wire252  &  wire852  &  wire30850 ) ;
 assign wire5146 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  n_n9587 ) ;
 assign wire5148 = ( nv10727  &  wire30853 ) | ( wire237  &  wire30853 ) | ( wire5875  &  wire30853 ) ;
 assign wire5150 = ( nv3280  &  wire30855 ) ;
 assign wire5151 = ( wire593  &  wire916 ) | ( wire593  &  wire5249 ) ;
 assign wire5152 = ( wire456  &  wire916 ) | ( wire456  &  wire5249 ) ;
 assign wire5166 = ( wire240  &  wire182 ) | ( wire182  &  wire5178 ) ;
 assign wire5167 = ( wire180  &  wire240 ) | ( ni33  &  wire180  &  nv2534 ) ;
 assign wire5168 = ( wire240  &  wire179 ) | ( ni33  &  wire179  &  nv2545 ) ;
 assign wire5169 = ( wire178  &  wire240 ) | ( wire178  &  wire5174 ) ;
 assign wire5174 = ( ni33  &  wire30444 ) | ( ni33  &  wire222  &  nv2330 ) ;
 assign wire5178 = ( ni33  &  wire30438 ) | ( ni35  &  ni33  &  n_n10835 ) ;
 assign wire5184 = ( wire240  &  wire179 ) | ( ni33  &  nv2235  &  wire179 ) ;
 assign wire5190 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2330 ) ;
 assign wire5196 = ( ni33  &  wire30502 ) | ( (~ ni36)  &  ni33  &  nv2314 ) ;
 assign wire5198 = ( wire240  &  wire30477 ) | ( ni33  &  nv2359  &  wire30477 ) ;
 assign wire5211 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2220 ) ;
 assign wire5215 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2276 ) ;
 assign wire5219 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2197 ) ;
 assign wire5223 = ( (~ ni34)  &  wire240 ) | ( (~ ni33)  &  wire240 ) | ( (~ ni34)  &  ni33  &  nv2397 ) ;
 assign wire5239 = ( pi17  &  pi19  &  (~ pi16)  &  wire916 ) ;
 assign wire5240 = ( pi17  &  (~ pi16)  &  wire1348 ) | ( pi17  &  (~ pi16)  &  wire5245 ) ;
 assign wire5241 = ( (~ pi25)  &  wire194  &  wire5745 ) | ( (~ pi25)  &  wire194  &  wire30778 ) ;
 assign wire5242 = ( pi17  &  pi19  &  pi16  &  wire916 ) ;
 assign wire5243 = ( pi17  &  pi16  &  wire1348 ) | ( pi17  &  pi16  &  wire5245 ) ;
 assign wire5244 = ( (~ pi25)  &  wire183  &  wire5745 ) | ( (~ pi25)  &  wire183  &  wire30778 ) ;
 assign wire5245 = ( (~ pi25)  &  wire189  &  wire5745 ) | ( (~ pi25)  &  wire189  &  wire30778 ) ;
 assign wire5247 = ( (~ pi25)  &  wire5745  &  wire30797 ) | ( (~ pi25)  &  wire30778  &  wire30797 ) ;
 assign wire5248 = ( (~ pi17)  &  pi20  &  wire162 ) | ( (~ pi17)  &  (~ pi20)  &  wire159 ) ;
 assign wire5249 = ( (~ pi25)  &  wire213  &  wire5745 ) | ( (~ pi25)  &  wire213  &  wire30778 ) ;
 assign wire5252 = ( wire30534  &  wire30890 ) | ( wire222  &  nv2766  &  wire30890 ) ;
 assign wire5253 = ( wire30530  &  wire30893 ) | ( wire238  &  nv3060  &  wire30893 ) ;
 assign wire5254 = ( wire321  &  wire30895 ) | ( ni38  &  nv2647  &  wire30895 ) ;
 assign wire5256 = ( wire1049  &  wire30899 ) | ( wire5607  &  wire30899 ) | ( wire5608  &  wire30899 ) ;
 assign wire5258 = ( wire307  &  wire30903 ) | ( wire5291  &  wire30903 ) | ( wire5292  &  wire30903 ) ;
 assign wire5261 = ( wire5286  &  wire30913 ) | ( wire5287  &  wire30913 ) | ( wire30636  &  wire30913 ) ;
 assign wire5262 = ( wire5273  &  wire30915 ) | ( wire5274  &  wire30915 ) | ( wire30646  &  wire30915 ) ;
 assign wire5263 = ( wire307  &  wire30917 ) | ( wire5278  &  wire30917 ) | ( wire5279  &  wire30917 ) ;
 assign wire5264 = ( wire151  &  wire5454  &  wire30918 ) | ( wire151  &  wire5455  &  wire30918 ) ;
 assign wire5267 = ( wire152  &  wire5454  &  wire30921 ) | ( wire152  &  wire5455  &  wire30921 ) ;
 assign wire5271 = ( wire30438  &  wire30639 ) | ( ni35  &  n_n10835  &  wire30639 ) ;
 assign wire5273 = ( wire1013  &  wire30641 ) | ( wire5557  &  wire30641 ) | ( wire5558  &  wire30641 ) ;
 assign wire5274 = ( (~ wire157)  &  wire179  &  nv3077  &  wire30524 ) ;
 assign wire5278 = ( wire315  &  wire30444 ) | ( wire222  &  wire315  &  nv2330 ) ;
 assign wire5279 = ( wire238  &  wire30534 ) | ( wire222  &  wire238  &  nv2766 ) ;
 assign wire5284 = ( wire30404  &  wire30629 ) | ( (~ ni35)  &  n_n10809  &  wire30629 ) ;
 assign wire5286 = ( wire1049  &  wire30631 ) | ( wire5607  &  wire30631 ) | ( wire5608  &  wire30631 ) ;
 assign wire5287 = ( wire178  &  (~ wire157)  &  nv3109  &  wire30524 ) ;
 assign wire5291 = ( wire216  &  wire315 ) | ( wire315  &  wire5873 ) | ( wire315  &  wire5917 ) ;
 assign wire5292 = ( wire321  &  wire238 ) | ( ni38  &  nv2647  &  wire238 ) ;
 assign wire5300 = ( wire321  &  wire30922 ) | ( wire5682  &  wire30922 ) ;
 assign wire5302 = ( wire1049  &  wire30924 ) | ( wire5710  &  wire30924 ) | ( wire5711  &  wire30924 ) ;
 assign wire5304 = ( wire158  &  wire1080  &  wire5325 ) | ( wire158  &  wire1080  &  wire30525 ) ;
 assign wire5305 = ( wire1013  &  wire30927 ) | ( wire5684  &  wire30927 ) | ( wire5685  &  wire30927 ) ;
 assign wire5307 = ( wire30560  &  wire30929 ) | ( nv2946  &  wire238  &  wire30929 ) ;
 assign wire5308 = ( wire5319  &  wire30930 ) | ( wire30553  &  wire30930 ) | ( wire30554  &  wire30930 ) ;
 assign wire5309 = ( wire5329  &  wire30931 ) | ( wire30573  &  wire30931 ) | ( wire30574  &  wire30931 ) ;
 assign wire5311 = ( wire5337  &  wire30933 ) | ( wire30540  &  wire30933 ) ;
 assign wire5312 = ( wire158  &  wire151  &  wire5454 ) | ( wire158  &  wire151  &  wire5455 ) ;
 assign wire5315 = ( wire302  &  wire152  &  wire5454 ) | ( wire302  &  wire152  &  wire5455 ) ;
 assign wire5317 = ( wire30422  &  wire30543 ) | ( ni35  &  n_n10922  &  wire30543 ) ;
 assign wire5319 = ( wire1013  &  wire30547 ) | ( wire5684  &  wire30547 ) | ( wire5685  &  wire30547 ) ;
 assign wire5325 = ( (~ wire157)  &  wire321  &  wire30524 ) | ( (~ wire157)  &  wire5682  &  wire30524 ) ;
 assign wire5327 = ( wire30374  &  wire30563 ) | ( (~ ni35)  &  n_n10896  &  wire30563 ) ;
 assign wire5329 = ( wire1049  &  wire30567 ) | ( wire5710  &  wire30567 ) | ( wire5711  &  wire30567 ) ;
 assign wire5334 = ( wire315  &  wire30432 ) | ( wire222  &  wire315  &  nv2220 ) ;
 assign wire5337 = ( wire315  &  wire30416 ) | ( wire222  &  nv2197  &  wire315 ) ;
 assign wire5340 = ( n_n10267  &  wire30951 ) | ( wire30528  &  wire30951 ) ;
 assign wire5344 = ( wire5602  &  wire30956 ) | ( wire5603  &  wire30956 ) | ( wire30610  &  wire30956 ) ;
 assign wire5346 = ( wire154  &  wire1080  &  wire5426 ) | ( wire154  &  wire1080  &  wire30579 ) ;
 assign wire5347 = ( wire5554  &  wire30959 ) | ( wire5555  &  wire30959 ) | ( wire30586  &  wire30959 ) ;
 assign wire5348 = ( wire5361  &  wire30960 ) | ( wire5362  &  wire30960 ) | ( wire30598  &  wire30960 ) ;
 assign wire5351 = ( wire5396  &  wire30963 ) | ( wire5397  &  wire30963 ) | ( wire30622  &  wire30963 ) ;
 assign wire5352 = ( wire30601  &  wire30964 ) | ( wire238  &  nv2766  &  wire30964 ) ;
 assign wire5353 = ( wire151  &  wire154  &  wire5454 ) | ( wire151  &  wire154  &  wire5455 ) ;
 assign wire5354 = ( wire152  &  wire1061  &  wire5454 ) | ( wire152  &  wire1061  &  wire5455 ) ;
 assign wire5361 = ( wire5554  &  wire30588 ) | ( wire5555  &  wire30588 ) | ( wire30586  &  wire30588 ) ;
 assign wire5362 = ( (~ wire157)  &  wire179  &  nv2807  &  wire30524 ) ;
 assign wire5366 = ( wire346  &  wire5895 ) | ( wire346  &  wire5898 ) | ( wire346  &  wire30382 ) ;
 assign wire5367 = ( ni37  &  ni36  &  wire5377 ) | ( ni37  &  ni36  &  wire5378 ) ;
 assign wire5368 = ( ni35  &  wire5376 ) | ( ni35  &  wire30441 ) ;
 assign wire5375 = ( wire834  &  wire5939 ) | ( wire834  &  wire30370 ) ;
 assign wire5376 = ( (~ ni36)  &  wire5377 ) | ( (~ ni36)  &  wire5378 ) ;
 assign wire5377 = ( wire254  &  wire5895 ) | ( wire254  &  wire5898 ) | ( wire254  &  wire30382 ) ;
 assign wire5378 = ( (~ ni40)  &  ni38  &  wire5939 ) | ( (~ ni40)  &  ni38  &  wire30370 ) ;
 assign wire5380 = ( wire270  &  wire5393 ) | ( nv2348  &  wire254  &  wire270 ) ;
 assign wire5381 = ( (~ ni36)  &  wire30438 ) | ( (~ ni36)  &  ni35  &  n_n10835 ) ;
 assign wire5386 = ( wire176  &  wire5393 ) | ( wire176  &  nv2348  &  wire254 ) ;
 assign wire5390 = ( wire847  &  wire5939 ) | ( wire847  &  wire30370 ) ;
 assign wire5391 = ( (~ ni36)  &  wire5393 ) | ( (~ ni36)  &  nv2348  &  wire254 ) ;
 assign wire5393 = ( (~ ni40)  &  ni38  &  wire5939 ) | ( (~ ni40)  &  ni38  &  wire30370 ) ;
 assign wire5396 = ( wire5602  &  wire30612 ) | ( wire5603  &  wire30612 ) | ( wire30610  &  wire30612 ) ;
 assign wire5397 = ( wire178  &  (~ wire157)  &  nv2857  &  wire30524 ) ;
 assign wire5401 = ( wire347  &  wire5895 ) | ( wire347  &  wire5898 ) | ( wire347  &  wire30382 ) ;
 assign wire5402 = ( ni37  &  ni36  &  wire5893 ) | ( ni37  &  ni36  &  wire5894 ) ;
 assign wire5404 = ( (~ ni35)  &  wire5884 ) | ( (~ ni35)  &  wire30409 ) ;
 assign wire5407 = ( wire270  &  wire5855 ) | ( nv2348  &  wire253  &  wire270 ) ;
 assign wire5409 = ( (~ ni36)  &  wire30404 ) | ( (~ ni36)  &  (~ ni35)  &  n_n10809 ) ;
 assign wire5414 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  nv2766 ) ;
 assign wire5416 = ( wire310  &  wire5895 ) | ( wire310  &  wire5898 ) | ( wire310  &  wire30382 ) ;
 assign wire5426 = ( (~ wire157)  &  wire5598  &  wire30524 ) | ( (~ wire157)  &  wire30524  &  wire30578 ) ;
 assign wire5429 = ( (~ ni36)  &  wire216 ) | ( (~ ni36)  &  wire5873 ) | ( (~ ni36)  &  wire5917 ) ;
 assign wire5431 = ( wire314  &  wire30980 ) | ( wire5653  &  wire30980 ) | ( wire5654  &  wire30980 ) ;
 assign wire5433 = ( wire5643  &  wire30982 ) | ( wire5644  &  wire30982 ) | ( wire30671  &  wire30982 ) ;
 assign wire5435 = ( wire307  &  wire30984 ) | ( wire5486  &  wire30984 ) | ( wire5487  &  wire30984 ) ;
 assign wire5436 = ( wire5636  &  wire30985 ) | ( wire5637  &  wire30985 ) | ( wire30655  &  wire30985 ) ;
 assign wire5437 = ( n_n10396  &  wire30986 ) | ( wire30558  &  wire30986 ) ;
 assign wire5439 = ( wire5463  &  wire30988 ) | ( wire30664  &  wire30988 ) | ( wire30665  &  wire30988 ) ;
 assign wire5440 = ( wire5494  &  wire30989 ) | ( wire30680  &  wire30989 ) | ( wire30681  &  wire30989 ) ;
 assign wire5442 = ( wire30651  &  wire30991 ) | ( nv2197  &  wire315  &  wire30991 ) ;
 assign wire5443 = ( wire158  &  wire151  &  wire5454 ) | ( wire158  &  wire151  &  wire5455 ) ;
 assign wire5446 = ( wire302  &  wire152  &  wire5454 ) | ( wire302  &  wire152  &  wire5455 ) ;
 assign wire5448 = ( (~ pi16)  &  wire5450 ) | ( (~ pi16)  &  wire5451 ) ;
 assign wire5450 = ( wire260  &  n_n9304 ) | ( pi21  &  wire260  &  n_n9302 ) ;
 assign wire5451 = ( wire228  &  n_n9304 ) | ( wire228  &  (~ wire157)  &  wire30397 ) ;
 assign wire5453 = ( pi21  &  n_n9294 ) ;
 assign wire5454 = ( ni33  &  wire216  &  wire30906 ) | ( ni33  &  wire5904  &  wire30906 ) ;
 assign wire5455 = ( (~ pi25)  &  wire164 ) ;
 assign wire5457 = ( pi20  &  n_n9304 ) | ( pi20  &  (~ wire157)  &  wire30397 ) ;
 assign wire5463 = ( wire5636  &  wire30657 ) | ( wire5637  &  wire30657 ) | ( wire30655  &  wire30657 ) ;
 assign wire5468 = ( n_n11076  &  wire346 ) | ( wire1319  &  wire346 ) ;
 assign wire5469 = ( wire270  &  wire5812 ) | ( wire253  &  wire270  &  nv2240 ) ;
 assign wire5470 = ( (~ ni36)  &  wire30422 ) | ( (~ ni36)  &  ni35  &  n_n10922 ) ;
 assign wire5473 = ( wire1319  &  wire346 ) | ( wire346  &  wire5898 ) | ( wire346  &  wire30382 ) ;
 assign wire5474 = ( ni37  &  ni36  &  wire5800 ) | ( ni37  &  ni36  &  wire5801 ) ;
 assign wire5475 = ( ni35  &  wire5797 ) | ( ni35  &  wire30423 ) ;
 assign wire5486 = ( wire315  &  wire30502 ) | ( (~ ni36)  &  wire315  &  nv2314 ) ;
 assign wire5487 = ( (~ wire157)  &  wire5654  &  wire30524 ) | ( (~ wire157)  &  wire30524  &  wire30649 ) ;
 assign wire5494 = ( wire5643  &  wire30673 ) | ( wire5644  &  wire30673 ) | ( wire30671  &  wire30673 ) ;
 assign wire5499 = ( n_n11076  &  wire347 ) | ( wire1319  &  wire347 ) ;
 assign wire5500 = ( wire270  &  wire5935 ) | ( wire254  &  wire270  &  nv2240 ) ;
 assign wire5501 = ( (~ ni36)  &  wire30374 ) | ( (~ ni36)  &  (~ ni35)  &  n_n10896 ) ;
 assign wire5504 = ( wire1319  &  wire347 ) | ( wire347  &  wire5898 ) | ( wire347  &  wire30382 ) ;
 assign wire5505 = ( ni37  &  ni36  &  wire5841 ) | ( ni37  &  ni36  &  wire5842 ) ;
 assign wire5507 = ( (~ ni35)  &  wire5838 ) | ( (~ ni35)  &  wire30383 ) ;
 assign wire5511 = ( wire30534  &  wire31045 ) | ( wire222  &  nv2766  &  wire31045 ) ;
 assign wire5512 = ( wire321  &  wire31047 ) | ( ni38  &  nv2647  &  wire31047 ) ;
 assign wire5513 = ( wire1013  &  wire31049 ) | ( wire5557  &  wire31049 ) | ( wire5558  &  wire31049 ) ;
 assign wire5514 = ( nv3077  &  wire486  &  wire31050 ) ;
 assign wire5516 = ( wire1049  &  wire31055 ) | ( wire5607  &  wire31055 ) | ( wire5608  &  wire31055 ) ;
 assign wire5517 = ( nv3109  &  wire486  &  wire31056 ) ;
 assign wire5518 = ( wire916  &  wire31058 ) | ( wire213  &  wire200  &  wire31058 ) ;
 assign wire5519 = ( wire1348  &  wire31059 ) | ( wire189  &  wire200  &  wire31059 ) ;
 assign wire5520 = ( wire916  &  wire31060 ) | ( wire213  &  wire200  &  wire31060 ) ;
 assign wire5521 = ( wire378  &  wire31061 ) | ( wire152  &  wire200  &  wire31061 ) ;
 assign wire5522 = ( wire1348  &  wire31062 ) | ( wire189  &  wire200  &  wire31062 ) ;
 assign wire5523 = ( wire916  &  wire31063 ) | ( wire213  &  wire200  &  wire31063 ) ;
 assign wire5524 = ( wire757  &  wire31064 ) | ( wire5744  &  wire31064 ) | ( wire5745  &  wire31064 ) ;
 assign wire5525 = ( wire692  &  wire5547 ) | ( wire692  &  wire763  &  wire200 ) ;
 assign wire5528 = ( pi15  &  (~ wire289)  &  wire31121 ) | ( pi15  &  (~ wire289)  &  wire31122 ) ;
 assign wire5529 = ( pi20  &  wire289  &  wire162 ) | ( (~ pi20)  &  wire289  &  wire159 ) ;
 assign wire5534 = ( wire5598  &  wire31067 ) | ( wire30578  &  wire31067 ) ;
 assign wire5535 = ( wire5554  &  wire31068 ) | ( wire5555  &  wire31068 ) | ( wire30586  &  wire31068 ) ;
 assign wire5537 = ( n_n10267  &  wire238  &  wire763 ) | ( wire238  &  wire763  &  wire30528 ) ;
 assign wire5538 = ( wire5602  &  wire31071 ) | ( wire5603  &  wire31071 ) | ( wire30610  &  wire31071 ) ;
 assign wire5539 = ( nv2857  &  wire31072 ) ;
 assign wire5540 = ( wire1340  &  wire916 ) | ( wire213  &  wire1340  &  wire200 ) ;
 assign wire5541 = ( wire1031  &  wire1348 ) | ( wire189  &  wire1031  &  wire200 ) ;
 assign wire5542 = ( wire1031  &  wire916 ) | ( wire213  &  wire1031  &  wire200 ) ;
 assign wire5543 = ( wire378  &  wire154 ) | ( wire152  &  wire154  &  wire200 ) ;
 assign wire5544 = ( wire593  &  wire1348 ) | ( wire189  &  wire593  &  wire200 ) ;
 assign wire5545 = ( wire593  &  wire916 ) | ( wire593  &  wire213  &  wire200 ) ;
 assign wire5547 = ( wire162  &  wire31065 ) ;
 assign wire5549 = ( wire310  &  n_n10590 ) | ( ni41  &  wire310  &  nv2647 ) ;
 assign wire5553 = ( wire270  &  wire5564 ) | ( wire254  &  wire270  &  nv2790 ) ;
 assign wire5554 = ( (~ ni36)  &  wire1013 ) | ( (~ ni36)  &  wire5557 ) | ( (~ ni36)  &  wire5558 ) ;
 assign wire5555 = ( ni35  &  wire5560 ) | ( ni35  &  wire5561 ) | ( ni35  &  wire5562 ) ;
 assign wire5557 = ( wire176  &  wire5564 ) | ( wire176  &  wire254  &  nv2790 ) ;
 assign wire5558 = ( ni35  &  wire5560 ) | ( ni35  &  wire5561 ) | ( ni35  &  wire5562 ) ;
 assign wire5560 = ( wire1192  &  wire886 ) | ( wire365  &  nv2790  &  wire886 ) ;
 assign wire5561 = ( wire847  &  nv2647 ) ;
 assign wire5562 = ( (~ ni36)  &  wire5564 ) | ( (~ ni36)  &  wire254  &  nv2790 ) ;
 assign wire5564 = ( (~ ni40)  &  ni38  &  nv2647 ) ;
 assign wire5565 = ( n_n10590  &  wire346 ) | ( ni41  &  nv2647  &  wire346 ) ;
 assign wire5566 = ( ni37  &  ni36  &  wire5578 ) | ( ni37  &  ni36  &  wire5579 ) ;
 assign wire5567 = ( ni35  &  wire5577 ) | ( ni35  &  wire30589 ) ;
 assign wire5576 = ( nv2647  &  wire834 ) ;
 assign wire5577 = ( (~ ni36)  &  wire5578 ) | ( (~ ni36)  &  wire253  &  nv2647 ) ;
 assign wire5578 = ( wire254  &  n_n10590 ) | ( ni41  &  wire254  &  nv2647 ) ;
 assign wire5579 = ( (~ ni40)  &  ni38  &  nv2647 ) ;
 assign wire5580 = ( wire347  &  n_n10590 ) | ( ni41  &  wire347  &  nv2647 ) ;
 assign wire5581 = ( ni37  &  ni36  &  wire5593 ) | ( ni37  &  ni36  &  wire5594 ) ;
 assign wire5583 = ( (~ ni35)  &  wire5590 ) | ( (~ ni35)  &  wire30613 ) ;
 assign wire5589 = ( wire814  &  nv2647 ) ;
 assign wire5590 = ( (~ ni36)  &  wire5594 ) | ( (~ ni36)  &  wire254  &  nv2647 ) ;
 assign wire5591 = ( wire400  &  n_n10590 ) | ( ni41  &  wire400  &  nv2647 ) ;
 assign wire5593 = ( ni40  &  ni38  &  nv2647 ) ;
 assign wire5594 = ( wire253  &  n_n10590 ) | ( ni41  &  wire253  &  nv2647 ) ;
 assign wire5598 = ( (~ ni36)  &  wire321 ) | ( ni38  &  (~ ni36)  &  nv2647 ) ;
 assign wire5601 = ( wire270  &  wire5613 ) | ( wire253  &  wire270  &  nv2790 ) ;
 assign wire5602 = ( (~ ni36)  &  wire1049 ) | ( (~ ni36)  &  wire5607 ) | ( (~ ni36)  &  wire5608 ) ;
 assign wire5603 = ( (~ ni35)  &  wire5610 ) | ( (~ ni35)  &  wire5611 ) | ( (~ ni35)  &  wire5612 ) ;
 assign wire5607 = ( wire177  &  wire5613 ) | ( wire177  &  wire253  &  nv2790 ) ;
 assign wire5608 = ( (~ ni35)  &  wire5610 ) | ( (~ ni35)  &  wire5611 ) | ( (~ ni35)  &  wire5612 ) ;
 assign wire5610 = ( wire882  &  wire1192 ) | ( wire365  &  nv2790  &  wire882 ) ;
 assign wire5611 = ( wire840  &  nv2647 ) ;
 assign wire5612 = ( (~ ni36)  &  wire5613 ) | ( (~ ni36)  &  wire253  &  nv2790 ) ;
 assign wire5613 = ( ni40  &  ni38  &  nv2647 ) ;
 assign wire5615 = ( wire314  &  wire31085 ) | ( wire5653  &  wire31085 ) | ( wire5654  &  wire31085 ) ;
 assign wire5616 = ( wire5636  &  wire31086 ) | ( wire5637  &  wire31086 ) | ( wire30655  &  wire31086 ) ;
 assign wire5618 = ( wire5643  &  wire31088 ) | ( wire5644  &  wire31088 ) | ( wire30671  &  wire31088 ) ;
 assign wire5619 = ( nv2694  &  wire31089 ) ;
 assign wire5620 = ( n_n10412  &  wire31090 ) | ( wire30538  &  wire31090 ) ;
 assign wire5621 = ( wire294  &  n_n10396  &  wire238 ) | ( wire294  &  wire238  &  wire30558 ) ;
 assign wire5622 = ( wire158  &  wire378 ) | ( wire158  &  wire152  &  wire200 ) ;
 assign wire5623 = ( wire698  &  wire1348 ) | ( wire189  &  wire698  &  wire200 ) ;
 assign wire5624 = ( wire698  &  wire916 ) | ( wire213  &  wire698  &  wire200 ) ;
 assign wire5625 = ( wire456  &  wire1348 ) | ( wire189  &  wire456  &  wire200 ) ;
 assign wire5626 = ( wire456  &  wire916 ) | ( wire456  &  wire213  &  wire200 ) ;
 assign wire5627 = ( wire344  &  wire916 ) | ( wire213  &  wire344  &  wire200 ) ;
 assign wire5629 = ( ni40  &  (~ ni37)  &  ni36  &  nv2602 ) ;
 assign wire5630 = ( ni37  &  ni36  &  wire5728 ) | ( ni37  &  ni36  &  wire5729 ) ;
 assign wire5632 = ( ni35  &  wire5723 ) | ( ni35  &  wire5724 ) | ( ni35  &  wire5725 ) ;
 assign wire5635 = ( wire270  &  wire5693 ) | ( wire254  &  wire270  &  nv2622 ) ;
 assign wire5636 = ( ni35  &  wire5687 ) | ( ni35  &  wire5688 ) | ( ni35  &  wire5689 ) ;
 assign wire5637 = ( (~ ni36)  &  wire1013 ) | ( (~ ni36)  &  wire5684 ) | ( (~ ni36)  &  wire5685 ) ;
 assign wire5639 = ( (~ ni41)  &  wire347  &  nv2647 ) | ( ni41  &  wire347  &  nv2183 ) ;
 assign wire5642 = ( wire270  &  wire5718 ) | ( wire253  &  wire270  &  nv2622 ) ;
 assign wire5643 = ( (~ ni35)  &  wire5713 ) | ( (~ ni35)  &  wire5714 ) | ( (~ ni35)  &  wire5715 ) ;
 assign wire5644 = ( (~ ni36)  &  wire1049 ) | ( (~ ni36)  &  wire5710 ) | ( (~ ni36)  &  wire5711 ) ;
 assign wire5646 = ( (~ ni40)  &  (~ ni37)  &  ni36  &  nv2602 ) ;
 assign wire5647 = ( ni37  &  ni36  &  wire5708 ) | ( ni37  &  ni36  &  wire5709 ) ;
 assign wire5648 = ( (~ ni35)  &  wire5703 ) | ( (~ ni35)  &  wire5704 ) | ( (~ ni35)  &  wire5705 ) ;
 assign wire5651 = ( (~ ni41)  &  nv2647  &  wire346 ) | ( ni41  &  nv2183  &  wire346 ) ;
 assign wire5653 = ( (~ ni41)  &  wire310  &  nv2647 ) | ( ni41  &  wire310  &  nv2183 ) ;
 assign wire5654 = ( (~ ni36)  &  wire321 ) | ( (~ ni36)  &  wire5682 ) ;
 assign wire5656 = ( wire321  &  wire31104 ) | ( wire5682  &  wire31104 ) ;
 assign wire5657 = ( wire1013  &  wire31105 ) | ( wire5684  &  wire31105 ) | ( wire5685  &  wire31105 ) ;
 assign wire5663 = ( wire158  &  wire378 ) | ( wire158  &  wire152  &  wire200 ) ;
 assign wire5664 = ( wire698  &  wire1348 ) | ( wire189  &  wire698  &  wire200 ) ;
 assign wire5665 = ( wire698  &  wire916 ) | ( wire213  &  wire698  &  wire200 ) ;
 assign wire5666 = ( wire456  &  wire1348 ) | ( wire189  &  wire456  &  wire200 ) ;
 assign wire5667 = ( wire456  &  wire916 ) | ( wire456  &  wire213  &  wire200 ) ;
 assign wire5668 = ( wire344  &  wire916 ) | ( wire213  &  wire344  &  wire200 ) ;
 assign wire5670 = ( wire697  &  wire162 ) ;
 assign wire5678 = ( ni33  &  (~ wire157)  &  wire216 ) | ( ni33  &  (~ wire157)  &  wire5904 ) ;
 assign wire5682 = ( (~ ni41)  &  ni38  &  nv2647 ) | ( ni41  &  ni38  &  nv2183 ) ;
 assign wire5684 = ( wire176  &  wire5693 ) | ( wire176  &  wire254  &  nv2622 ) ;
 assign wire5685 = ( ni35  &  wire5687 ) | ( ni35  &  wire5688 ) | ( ni35  &  wire5689 ) ;
 assign wire5687 = ( wire1192  &  wire886 ) | ( wire365  &  nv2622  &  wire886 ) ;
 assign wire5688 = ( (~ ni41)  &  wire847  &  nv2647 ) | ( ni41  &  wire847  &  nv2183 ) ;
 assign wire5689 = ( (~ ni36)  &  wire5693 ) | ( (~ ni36)  &  wire254  &  nv2622 ) ;
 assign wire5693 = ( (~ ni41)  &  wire253  &  nv2647 ) | ( ni41  &  wire253  &  nv2183 ) ;
 assign wire5703 = ( wire1195  &  wire883 ) | ( wire400  &  nv2602  &  wire883 ) ;
 assign wire5704 = ( (~ ni41)  &  wire814  &  nv2647 ) | ( ni41  &  wire814  &  nv2183 ) ;
 assign wire5705 = ( (~ ni36)  &  wire5708 ) | ( (~ ni36)  &  wire253  &  nv2602 ) ;
 assign wire5708 = ( (~ ni41)  &  wire254  &  nv2647 ) | ( ni41  &  wire254  &  nv2183 ) ;
 assign wire5709 = ( (~ ni40)  &  ni38  &  nv2602 ) ;
 assign wire5710 = ( wire177  &  wire5718 ) | ( wire177  &  wire253  &  nv2622 ) ;
 assign wire5711 = ( (~ ni35)  &  wire5713 ) | ( (~ ni35)  &  wire5714 ) | ( (~ ni35)  &  wire5715 ) ;
 assign wire5713 = ( wire882  &  wire1192 ) | ( wire365  &  wire882  &  nv2622 ) ;
 assign wire5714 = ( (~ ni41)  &  wire840  &  nv2647 ) | ( ni41  &  wire840  &  nv2183 ) ;
 assign wire5715 = ( (~ ni36)  &  wire5718 ) | ( (~ ni36)  &  wire253  &  nv2622 ) ;
 assign wire5718 = ( (~ ni41)  &  wire254  &  nv2647 ) | ( ni41  &  wire254  &  nv2183 ) ;
 assign wire5723 = ( wire1195  &  wire885 ) | ( wire400  &  nv2602  &  wire885 ) ;
 assign wire5724 = ( (~ ni41)  &  nv2647  &  wire834 ) | ( ni41  &  nv2183  &  wire834 ) ;
 assign wire5725 = ( (~ ni36)  &  wire5729 ) | ( (~ ni36)  &  wire254  &  nv2602 ) ;
 assign wire5728 = ( ni40  &  ni38  &  nv2602 ) ;
 assign wire5729 = ( (~ ni41)  &  wire253  &  nv2647 ) | ( ni41  &  wire253  &  nv2183 ) ;
 assign wire5744 = ( ni33  &  wire924  &  wire216 ) | ( ni33  &  wire924  &  wire5904 ) ;
 assign wire5745 = ( (~ ni33)  &  wire924  &  wire866 ) ;
 assign wire5770 = ( ni33  &  wire30416 ) | ( ni33  &  wire222  &  nv2197 ) ;
 assign wire5775 = ( wire1319  &  wire310 ) | ( wire310  &  wire5898 ) | ( wire310  &  wire30382 ) ;
 assign wire5778 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2314 ) ;
 assign wire5788 = ( wire240  &  wire179 ) | ( ni33  &  wire179  &  nv2473 ) ;
 assign wire5796 = ( nv2240  &  wire834 ) ;
 assign wire5797 = ( (~ ni36)  &  wire5800 ) | ( (~ ni36)  &  wire253  &  nv2240 ) ;
 assign wire5798 = ( ni39  &  (~ ni38)  &  n_n11266 ) | ( ni39  &  (~ ni38)  &  wire5930 ) ;
 assign wire5800 = ( wire1319  &  wire254 ) | ( wire254  &  wire5898 ) | ( wire254  &  wire30382 ) ;
 assign wire5801 = ( (~ ni40)  &  ni38  &  nv2240 ) ;
 assign wire5802 = ( ni33  &  wire30422 ) | ( ni35  &  ni33  &  n_n10922 ) ;
 assign wire5804 = ( wire176  &  wire5812 ) | ( wire176  &  wire253  &  nv2240 ) ;
 assign wire5808 = ( nv2240  &  wire847 ) ;
 assign wire5809 = ( (~ ni36)  &  wire5812 ) | ( (~ ni36)  &  wire253  &  nv2240 ) ;
 assign wire5810 = ( (~ ni39)  &  (~ ni38)  &  n_n11266 ) | ( (~ ni39)  &  (~ ni38)  &  wire5930 ) ;
 assign wire5812 = ( ni40  &  ni38  &  n_n11076 ) | ( ni40  &  ni38  &  wire1319 ) ;
 assign wire5816 = ( (~ pi21)  &  (~ ni45)  &  (~ wire157) ) ;
 assign wire5829 = ( wire240  &  wire252 ) | ( ni33  &  wire252  &  nv2493 ) ;
 assign wire5837 = ( wire814  &  nv2240 ) ;
 assign wire5838 = ( (~ ni36)  &  wire5842 ) | ( (~ ni36)  &  wire254  &  nv2240 ) ;
 assign wire5839 = ( wire1319  &  wire400 ) | ( wire400  &  wire5898 ) | ( wire400  &  wire30382 ) ;
 assign wire5841 = ( ni40  &  ni38  &  nv2240 ) ;
 assign wire5842 = ( wire1319  &  wire253 ) | ( wire253  &  wire5898 ) | ( wire253  &  wire30382 ) ;
 assign wire5845 = ( ni33  &  wire30404 ) | ( (~ ni35)  &  ni33  &  n_n10809 ) ;
 assign wire5847 = ( wire177  &  wire5855 ) | ( wire177  &  nv2348  &  wire253 ) ;
 assign wire5851 = ( wire840  &  wire5939 ) | ( wire840  &  wire30370 ) ;
 assign wire5852 = ( (~ ni36)  &  wire5855 ) | ( (~ ni36)  &  nv2348  &  wire253 ) ;
 assign wire5855 = ( ni40  &  ni38  &  wire5939 ) | ( ni40  &  ni38  &  wire30370 ) ;
 assign wire5861 = ( ni33  &  wire30432 ) | ( ni33  &  wire222  &  nv2220 ) ;
 assign wire5871 = ( ni33  &  wire216 ) | ( ni33  &  wire5873 ) | ( ni33  &  wire5917 ) ;
 assign wire5873 = ( ni38  &  wire5939 ) | ( ni38  &  wire30370 ) ;
 assign wire5875 = ( wire240  &  wire252 ) | ( ni33  &  nv2565  &  wire252 ) ;
 assign wire5883 = ( wire814  &  wire5939 ) | ( wire814  &  wire30370 ) ;
 assign wire5884 = ( (~ ni36)  &  wire5893 ) | ( (~ ni36)  &  wire5894 ) ;
 assign wire5885 = ( ni39  &  (~ ni38)  &  n_n11266 ) | ( ni39  &  (~ ni38)  &  wire5930 ) ;
 assign wire5887 = ( wire400  &  wire5895 ) | ( wire400  &  wire5898 ) | ( wire400  &  wire30382 ) ;
 assign wire5889 = ( (~ ni38)  &  wire404  &  n_n11266 ) | ( (~ ni38)  &  wire404  &  wire5930 ) ;
 assign wire5893 = ( ni40  &  ni38  &  wire5939 ) | ( ni40  &  ni38  &  wire30370 ) ;
 assign wire5894 = ( wire253  &  wire5895 ) | ( wire253  &  wire5898 ) | ( wire253  &  wire30382 ) ;
 assign wire5895 = ( ni41  &  wire5939 ) | ( ni41  &  wire30370 ) ;
 assign wire5897 = ( wire5941  &  wire30380 ) | ( wire5945  &  wire30380 ) | ( wire30369  &  wire30380 ) ;
 assign wire5898 = ( wire5939  &  wire30381 ) | ( wire30370  &  wire30381 ) ;
 assign wire5902 = ( ni34  &  ni33  &  (~ nv6428) ) ;
 assign wire5904 = ( wire172  &  wire5941 ) | ( wire172  &  wire5945 ) | ( wire172  &  wire30369 ) ;
 assign wire5906 = ( ni33  &  wire30374 ) | ( (~ ni35)  &  ni33  &  n_n10896 ) ;
 assign wire5914 = ( wire177  &  wire5935 ) | ( wire177  &  wire254  &  nv2240 ) ;
 assign wire5917 = ( (~ ni38)  &  (~ ni37)  &  n_n11266 ) | ( (~ ni38)  &  (~ ni37)  &  wire5930 ) ;
 assign wire5920 = ( nv2240  &  wire840 ) ;
 assign wire5921 = ( (~ ni36)  &  wire5935 ) | ( (~ ni36)  &  wire254  &  nv2240 ) ;
 assign wire5922 = ( (~ ni39)  &  (~ ni38)  &  n_n11266 ) | ( (~ ni39)  &  (~ ni38)  &  wire5930 ) ;
 assign wire5924 = ( n_n11076  &  wire365 ) | ( wire1319  &  wire365 ) ;
 assign wire5926 = ( (~ ni38)  &  (~ wire342)  &  n_n11266 ) | ( (~ ni38)  &  (~ wire342)  &  wire5930 ) ;
 assign wire5930 = ( (~ ni42)  &  nv2176 ) ;
 assign wire5932 = ( ni43  &  ni42  &  nv2176 ) ;
 assign wire5935 = ( (~ ni40)  &  ni38  &  n_n11076 ) | ( (~ ni40)  &  ni38  &  wire1319 ) ;
 assign wire5939 = ( ni43  &  wire30369 ) | ( ni43  &  ni42  &  nv2186 ) | ( ni43  &  (~ ni42)  &  nv2186 ) ;
 assign wire5941 = ( (~ ni42)  &  nv2186 ) ;
 assign wire5945 = ( ni43  &  ni42  &  nv2186 ) ;
 assign wire5946 = ( ni43  &  (~ ni41)  &  nv2186 ) ;
 assign wire5948 = ( (~ ni43)  &  (~ ni41)  &  ni44  &  nv2186 ) ;
 assign wire5960 = ( ni2  &  ni9 ) | ( ni3  &  ni9 ) ;
 assign wire5961 = ( ni9  &  ni7 ) | ( (~ ni10)  &  ni7 ) | ( ni7  &  ni8 ) ;
 assign wire5962 = ( (~ pi23)  &  ni7 ) | ( pi24  &  ni7 ) ;
 assign wire5963 = ( wire1289  &  wire264  &  wire29692 ) | ( wire1289  &  wire264  &  wire29693 ) ;
 assign wire5964 = ( wire6509  &  wire29743 ) | ( wire6515  &  wire29743 ) | ( wire29741  &  wire29743 ) ;
 assign wire5965 = ( wire6636  &  wire29790 ) | ( wire6642  &  wire29790 ) | ( wire29789  &  wire29790 ) ;
 assign wire5966 = ( wire5990  &  wire29838 ) | ( wire29835  &  wire29838 ) | ( wire29836  &  wire29838 ) ;
 assign wire5967 = ( n_n11570  &  wire29885 ) ;
 assign wire5968 = ( wire29692  &  wire29886 ) | ( wire29693  &  wire29886 ) ;
 assign wire5975 = ( wire29515  &  wire29796 ) | ( (~ ni29)  &  wire1046  &  wire29796 ) ;
 assign wire5976 = ( ni34  &  wire29798 ) | ( (~ nv952)  &  (~ wire157)  &  wire29798 ) ;
 assign wire5978 = ( wire317  &  wire29802 ) | ( wire6252  &  wire29802 ) | ( wire6253  &  wire29802 ) ;
 assign wire5979 = ( ni34  &  wire29803 ) | ( (~ wire157)  &  (~ nv942)  &  wire29803 ) ;
 assign wire5982 = ( wire29532  &  wire29806 ) | ( (~ ni29)  &  wire1038  &  wire29806 ) ;
 assign wire5983 = ( ni34  &  nv942  &  wire29807 ) ;
 assign wire5984 = ( wire29809  &  wire29810 ) | ( (~ wire150)  &  n_n11474  &  wire29810 ) ;
 assign wire5987 = ( ni34  &  wire29813 ) | ( (~ wire157)  &  (~ nv858)  &  wire29813 ) ;
 assign wire5988 = ( ni34  &  wire257  &  nv858 ) ;
 assign wire5989 = ( wire317  &  wire29815 ) | ( wire6246  &  wire29815 ) | ( wire6247  &  wire29815 ) ;
 assign wire5990 = ( wire1073  &  wire6079 ) | ( wire1073  &  wire6081 ) | ( wire1073  &  wire29816 ) ;
 assign wire5992 = ( pi16  &  wire6652 ) | ( pi16  &  wire260  &  wire224 ) ;
 assign wire5999 = ( ni34  &  wire247  &  wire29905 ) | ( wire247  &  (~ wire943)  &  wire29905 ) ;
 assign wire6001 = ( ni34  &  wire29914 ) | ( (~ wire157)  &  (~ nv942)  &  wire29914 ) ;
 assign wire6003 = ( ni34  &  wire29922 ) | ( (~ nv952)  &  (~ wire157)  &  wire29922 ) ;
 assign wire6004 = ( ni34  &  wire29926 ) | ( (~ wire157)  &  (~ nv873)  &  wire29926 ) ;
 assign wire6007 = ( wire289  &  nv928  &  wire393  &  wire29933 ) ;
 assign wire6011 = ( wire6089  &  wire29958 ) | ( wire29954  &  wire29958 ) | ( wire29955  &  wire29958 ) ;
 assign wire6012 = ( wire29967  &  wire29972 ) | ( wire29968  &  wire29972 ) | ( wire29970  &  wire29972 ) ;
 assign wire6013 = ( (~ pi17)  &  wire289  &  wire343  &  wire29973 ) ;
 assign wire6016 = ( ni34  &  wire29977 ) | ( (~ nv952)  &  (~ wire157)  &  wire29977 ) ;
 assign wire6017 = ( ni34  &  (~ nv6428)  &  wire29979 ) | ( ni34  &  nv952  &  wire29979 ) ;
 assign wire6018 = ( ni34  &  wire6617  &  wire29981 ) | ( ni34  &  wire29512  &  wire29981 ) ;
 assign wire6019 = ( ni34  &  wire395  &  nv942  &  wire29982 ) ;
 assign wire6025 = ( wire184  &  wire29995 ) | ( wire6479  &  wire29995 ) ;
 assign wire6027 = ( wire29809  &  wire29997 ) | ( (~ wire150)  &  n_n11474  &  wire29997 ) ;
 assign wire6028 = ( wire6457  &  wire29999 ) | ( wire29998  &  wire29999 ) ;
 assign wire6030 = ( ni34  &  wire30001 ) | ( (~ wire157)  &  (~ nv942)  &  wire30001 ) ;
 assign wire6032 = ( wire184  &  wire30003 ) | ( wire6475  &  wire30003 ) ;
 assign wire6035 = ( wire271  &  wire485 ) | ( pi25  &  wire184  &  wire485 ) ;
 assign wire6038 = ( ni34  &  wire6683  &  wire30016 ) | ( ni34  &  wire29470  &  wire30016 ) ;
 assign wire6040 = ( wire302  &  wire225  &  wire617  &  nv899 ) ;
 assign wire6041 = ( pi25  &  ni34  &  nv873  &  wire1293 ) ;
 assign wire6042 = ( ni34  &  nv883  &  wire30023 ) ;
 assign wire6047 = ( ni34  &  wire225  &  wire843 ) | ( wire225  &  wire843  &  (~ wire943) ) ;
 assign wire6049 = ( ni34  &  wire30032 ) | ( (~ wire157)  &  (~ nv873)  &  wire30032 ) ;
 assign wire6050 = ( wire6366  &  wire30034 ) | ( wire30033  &  wire30034 ) ;
 assign wire6056 = ( wire766  &  nv1424  &  wire30038 ) ;
 assign wire6059 = ( ni34  &  wire320  &  wire30043 ) | ( ni34  &  wire6694  &  wire30043 ) ;
 assign wire6062 = ( pi22  &  pi25  &  wire184  &  wire30047 ) ;
 assign wire6066 = ( wire299  &  wire271 ) | ( pi25  &  wire299  &  wire184 ) ;
 assign wire6074 = ( wire1095  &  wire6079 ) | ( wire1095  &  wire6081 ) | ( wire1095  &  wire29816 ) ;
 assign wire6077 = ( pi22  &  pi25  &  wire184  &  wire766 ) ;
 assign wire6079 = ( pi21  &  ni34  &  wire6561 ) | ( pi21  &  ni34  &  wire29526 ) ;
 assign wire6081 = ( pi21  &  pi22  &  wire6255 ) | ( pi21  &  pi22  &  wire29528 ) ;
 assign wire6087 = ( nv750  &  wire29949 ) ;
 assign wire6089 = ( pi25  &  wire180  &  wire154  &  nv835 ) ;
 assign wire6095 = ( ni34  &  wire29962 ) | ( (~ wire785)  &  wire29962 ) ;
 assign wire6103 = ( ni34  &  wire714  &  wire30096 ) | ( wire714  &  wire6524  &  wire30096 ) ;
 assign wire6105 = ( wire1048  &  wire507  &  wire30100 ) ;
 assign wire6111 = ( ni34  &  wire30115 ) | ( wire6524  &  wire30115 ) ;
 assign wire6114 = ( wire6567  &  wire30119 ) | ( wire6569  &  wire30119 ) | ( wire29713  &  wire30119 ) ;
 assign wire6119 = ( nv1291  &  wire30125 ) ;
 assign wire6122 = ( wire271  &  wire1071 ) | ( pi25  &  wire184  &  wire1071 ) ;
 assign wire6123 = ( wire614  &  wire6132 ) | ( wire614  &  wire30134 ) | ( wire614  &  wire30135 ) ;
 assign wire6124 = ( (~ pi15)  &  wire6152 ) | ( (~ pi15)  &  wire30194 ) | ( (~ pi15)  &  wire30195 ) ;
 assign wire6127 = ( (~ pi19)  &  (~ pi20)  &  (~ nv6428)  &  (~ n_n12655) ) ;
 assign wire6132 = ( wire1095  &  wire6547 ) | ( wire1095  &  wire6549 ) | ( wire1095  &  wire29721 ) ;
 assign wire6135 = ( pi22  &  pi25  &  wire184  &  wire766 ) ;
 assign wire6138 = ( nv1073  &  wire617  &  wire30140 ) ;
 assign wire6140 = ( pi25  &  wire1012  &  wire1293 ) | ( (~ ni34)  &  wire1012  &  wire1293 ) ;
 assign wire6143 = ( ni34  &  nv644  &  wire30148 ) ;
 assign wire6145 = ( wire6429  &  wire30151 ) | ( wire30150  &  wire30151 ) ;
 assign wire6152 = ( (~ pi16)  &  wire30178 ) | ( (~ pi16)  &  wire30179 ) | ( (~ pi16)  &  wire30181 ) ;
 assign wire6154 = ( pi25  &  wire184  &  wire1293 ) ;
 assign wire6155 = ( (~ pi21)  &  ni34  &  wire344 ) | ( (~ pi22)  &  ni34  &  wire344 ) ;
 assign wire6156 = ( pi25  &  (~ nv6428)  &  wire260 ) | ( (~ ni34)  &  (~ nv6428)  &  wire260 ) ;
 assign wire6157 = ( (~ pi20)  &  pi25  &  (~ ni34)  &  wire153 ) ;
 assign wire6159 = ( nv1117  &  wire766  &  wire30160 ) ;
 assign wire6161 = ( ni34  &  wire6691  &  wire30164 ) | ( ni34  &  wire29623  &  wire30164 ) ;
 assign wire6165 = ( pi22  &  pi25  &  wire184  &  wire30169 ) ;
 assign wire6169 = ( wire299  &  wire271 ) | ( pi25  &  wire299  &  wire184 ) ;
 assign wire6170 = ( pi25  &  (~ ni34)  &  wire272 ) ;
 assign wire6171 = ( pi17  &  pi19  &  (~ nv6428)  &  (~ n_n12655) ) ;
 assign wire6172 = ( pi22  &  pi25  &  (~ ni34) ) ;
 assign wire6174 = ( ni34  &  wire228  &  nv883  &  wire29839 ) ;
 assign wire6176 = ( (~ wire150)  &  wire312  &  nv899  &  wire29843 ) ;
 assign wire6177 = ( wire29472  &  wire29846 ) | ( (~ ni29)  &  wire1033  &  wire29846 ) ;
 assign wire6179 = ( wire228  &  wire6281  &  wire29849 ) | ( wire228  &  wire29479  &  wire29849 ) ;
 assign wire6180 = ( ni34  &  wire29851 ) | ( (~ wire157)  &  (~ nv873)  &  wire29851 ) ;
 assign wire6182 = ( (~ wire150)  &  nv919  &  wire312  &  wire1058 ) ;
 assign wire6184 = ( ni34  &  nv873  &  wire29855 ) ;
 assign wire6185 = ( wire6196  &  wire29858 ) | ( wire6198  &  wire29858 ) | ( wire29856  &  wire29858 ) ;
 assign wire6189 = ( wire317  &  wire29862 ) | ( wire6284  &  wire29862 ) | ( wire6285  &  wire29862 ) ;
 assign wire6190 = ( wire1066  &  wire6200 ) | ( wire1066  &  wire6202 ) | ( wire1066  &  wire29863 ) ;
 assign wire6192 = ( pi17  &  pi19  &  (~ pi16)  &  wire1036 ) ;
 assign wire6193 = ( (~ pi16)  &  wire6652 ) | ( (~ pi16)  &  wire260  &  wire224 ) ;
 assign wire6196 = ( pi21  &  ni34  &  wire6667 ) | ( pi21  &  ni34  &  wire29466 ) ;
 assign wire6198 = ( pi21  &  pi22  &  wire6287 ) | ( pi21  &  pi22  &  wire29468 ) ;
 assign wire6200 = ( pi21  &  ni34  &  wire6746 ) | ( pi21  &  ni34  &  wire29449 ) ;
 assign wire6202 = ( pi21  &  pi22  &  wire6334 ) | ( pi21  &  pi22  &  wire29452 ) ;
 assign wire6205 = ( wire29452  &  wire29454 ) | ( (~ ni29)  &  wire1312  &  wire29454 ) ;
 assign wire6206 = ( pi15  &  nv919  &  wire1058  &  wire376 ) ;
 assign wire6207 = ( wire29458  &  wire29460 ) | ( (~ ni29)  &  wire1039  &  wire29460 ) ;
 assign wire6209 = ( pi21  &  pi15  &  ni34  &  wire1066 ) ;
 assign wire6210 = ( pi21  &  pi15  &  ni34  &  wire1058 ) ;
 assign wire6217 = ( ni34  &  wire320  &  wire29495 ) | ( ni34  &  wire6694  &  wire29495 ) ;
 assign wire6224 = ( wire29515  &  wire29517 ) | ( (~ ni29)  &  wire1046  &  wire29517 ) ;
 assign wire6225 = ( ni34  &  wire29521 ) | ( (~ nv952)  &  (~ wire157)  &  wire29521 ) ;
 assign wire6226 = ( wire317  &  wire29525 ) | ( wire6252  &  wire29525 ) | ( wire6253  &  wire29525 ) ;
 assign wire6228 = ( wire29528  &  wire29529 ) | ( (~ ni29)  &  wire1313  &  wire29529 ) ;
 assign wire6230 = ( wire29532  &  wire29533 ) | ( (~ ni29)  &  wire1038  &  wire29533 ) ;
 assign wire6231 = ( ni34  &  wire29536 ) | ( (~ wire157)  &  (~ nv942)  &  wire29536 ) ;
 assign wire6235 = ( ni34  &  wire29540 ) | ( (~ wire157)  &  (~ nv858)  &  wire29540 ) ;
 assign wire6236 = ( wire317  &  wire29542 ) | ( wire6246  &  wire29542 ) | ( wire6247  &  wire29542 ) ;
 assign wire6239 = ( pi16  &  wire6332 ) | ( pi16  &  wire6333 ) ;
 assign wire6240 = ( pi17  &  pi19  &  pi16  &  ni34 ) ;
 assign wire6242 = ( ni34  &  nv858  &  wire29499 ) ;
 assign wire6243 = ( ni34  &  wire29501 ) | ( (~ wire157)  &  (~ nv858)  &  wire29501 ) ;
 assign wire6246 = ( ni34  &  (~ ni29)  &  nv942 ) ;
 assign wire6247 = ( ni34  &  wire332 ) | ( (~ wire157)  &  wire332  &  (~ nv942) ) ;
 assign wire6249 = ( (~ nv6428)  &  wire29507 ) | ( wire6581  &  wire29507 ) | ( wire29504  &  wire29507 ) ;
 assign wire6252 = ( (~ ni34)  &  (~ ni29)  &  (~ nv952)  &  (~ wire157) ) ;
 assign wire6253 = ( ni34  &  (~ ni29)  &  (~ nv6428) ) | ( ni34  &  (~ ni29)  &  nv952 ) ;
 assign wire6255 = ( ni34  &  (~ ni29)  &  wire6561 ) | ( ni34  &  (~ ni29)  &  wire29526 ) ;
 assign wire6269 = ( wire29472  &  wire29473 ) | ( (~ ni29)  &  wire1033  &  wire29473 ) ;
 assign wire6270 = ( ni34  &  wire228  &  wire376 ) | ( wire228  &  (~ wire943)  &  wire376 ) ;
 assign wire6271 = ( wire228  &  (~ wire150)  &  wire6281 ) | ( wire228  &  (~ wire150)  &  wire29479 ) ;
 assign wire6272 = ( ni34  &  wire1030 ) | ( (~ wire157)  &  (~ nv873)  &  wire1030 ) ;
 assign wire6276 = ( wire317  &  wire169 ) | ( wire169  &  wire6284 ) | ( wire169  &  wire6285 ) ;
 assign wire6281 = ( ni34  &  (~ ni29)  &  nv883 ) ;
 assign wire6284 = ( ni34  &  (~ ni29)  &  nv873 ) ;
 assign wire6285 = ( ni34  &  wire332 ) | ( (~ wire157)  &  wire332  &  (~ nv873) ) ;
 assign wire6287 = ( ni34  &  (~ ni29)  &  wire6667 ) | ( ni34  &  (~ ni29)  &  wire29466 ) ;
 assign wire6291 = ( wire29572  &  wire29574 ) | ( (~ ni29)  &  wire1282  &  wire29574 ) ;
 assign wire6293 = ( wire29579  &  wire29581 ) | ( (~ ni29)  &  wire1008  &  wire29581 ) ;
 assign wire6295 = ( wire29584  &  wire29586 ) | ( (~ ni29)  &  wire1070  &  wire29586 ) ;
 assign wire6297 = ( wire29590  &  wire29591 ) | ( (~ ni29)  &  wire1318  &  wire29591 ) ;
 assign wire6305 = ( wire29602  &  wire29603 ) | ( (~ ni29)  &  wire1048  &  wire29603 ) ;
 assign wire6308 = ( pi16  &  wire6332 ) | ( pi16  &  wire6333 ) ;
 assign wire6309 = ( pi17  &  pi19  &  pi16  &  ni34 ) ;
 assign wire6312 = ( wire29632  &  wire29634 ) | ( (~ ni29)  &  wire1310  &  wire29634 ) ;
 assign wire6314 = ( wire29639  &  wire29641 ) | ( (~ ni29)  &  wire1057  &  wire29641 ) ;
 assign wire6315 = ( ni34  &  wire376  &  wire29642 ) | ( (~ wire785)  &  wire376  &  wire29642 ) ;
 assign wire6316 = ( wire228  &  wire6714  &  wire29645 ) | ( wire228  &  wire29644  &  wire29645 ) ;
 assign wire6318 = ( wire29650  &  wire29651 ) | ( (~ ni29)  &  wire1332  &  wire29651 ) ;
 assign wire6319 = ( nv717  &  wire1058  &  wire376 ) ;
 assign wire6325 = ( n_n13390  &  wire158  &  nv735  &  wire152 ) ;
 assign wire6326 = ( wire29662  &  wire29663 ) | ( (~ ni29)  &  wire1012  &  wire29663 ) ;
 assign wire6329 = ( (~ pi16)  &  wire6332 ) | ( (~ pi16)  &  wire6333 ) ;
 assign wire6330 = ( pi17  &  pi19  &  (~ pi16)  &  ni34 ) ;
 assign wire6332 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  ni34 ) ;
 assign wire6333 = ( (~ pi17)  &  (~ pi21)  &  ni34 ) ;
 assign wire6334 = ( ni34  &  (~ ni29)  &  wire6746 ) | ( ni34  &  (~ ni29)  &  wire29449 ) ;
 assign wire6337 = ( ni34  &  (~ ni29)  &  wire6706 ) | ( ni34  &  (~ ni29)  &  wire29455 ) ;
 assign wire6351 = ( wire184  &  wire30265 ) | ( wire6479  &  wire30265 ) ;
 assign wire6354 = ( wire294  &  wire6450  &  wire30270 ) | ( wire294  &  wire30028  &  wire30270 ) ;
 assign wire6355 = ( wire6457  &  wire30272 ) | ( wire29998  &  wire30272 ) ;
 assign wire6366 = ( ni34  &  ni32  &  (~ ni31) ) | ( ni34  &  (~ ni31)  &  ni30 ) ;
 assign wire6401 = ( wire6429  &  wire30291 ) | ( wire30150  &  wire30291 ) ;
 assign wire6402 = ( nv1009  &  wire30292 ) ;
 assign wire6429 = ( ni34  &  (~ nv6428) ) | ( (~ nv6428)  &  (~ wire785) ) ;
 assign wire6450 = ( ni34  &  (~ nv6428) ) | ( (~ nv6428)  &  (~ wire943) ) ;
 assign wire6453 = ( ni36  &  n_n13028 ) | ( (~ ni36)  &  n_n13028 ) | ( n_n13028  &  wire6717 ) | ( n_n13028  &  wire29474 ) ;
 assign wire6454 = ( n_n13271  &  wire6722 ) | ( n_n13271  &  wire29474 ) | ( n_n13271  &  wire29475 ) ;
 assign wire6457 = ( ni34  &  ni32  &  (~ ni31) ) | ( ni34  &  (~ ni31)  &  ni30 ) ;
 assign wire6475 = ( ni34  &  nv858 ) | ( ni34  &  (~ ni31)  &  (~ wire7195) ) ;
 assign wire6479 = ( ni34  &  (~ nv6428) ) | ( ni34  &  wire6581 ) | ( ni34  &  wire29504 ) ;
 assign wire6498 = ( wire228  &  wire1070  &  wire29695 ) ;
 assign wire6499 = ( wire1008  &  wire381  &  wire29697 ) ;
 assign wire6501 = ( wire29579  &  wire29702 ) | ( (~ ni29)  &  wire1008  &  wire29702 ) ;
 assign wire6503 = ( wire29584  &  wire29706 ) | ( (~ ni29)  &  wire1070  &  wire29706 ) ;
 assign wire6505 = ( pi21  &  wire1112  &  wire1045 ) | ( (~ ni34)  &  wire1112  &  wire1045 ) ;
 assign wire6506 = ( ni34  &  n_n12706  &  wire29709 ) | ( ni34  &  wire29534  &  wire29709 ) ;
 assign wire6508 = ( wire29595  &  wire29711 ) | ( (~ ni29)  &  wire1112  &  wire29711 ) ;
 assign wire6509 = ( wire6567  &  wire29715 ) | ( wire6569  &  wire29715 ) | ( wire29713  &  wire29715 ) ;
 assign wire6513 = ( ni34  &  wire29719 ) | ( wire6524  &  wire29719 ) ;
 assign wire6514 = ( wire29602  &  wire29720 ) | ( (~ ni29)  &  wire1048  &  wire29720 ) ;
 assign wire6515 = ( wire1073  &  wire6547 ) | ( wire1073  &  wire6549 ) | ( wire1073  &  wire29721 ) ;
 assign wire6517 = ( pi16  &  wire6652 ) | ( pi16  &  wire260  &  wire224 ) ;
 assign wire6521 = ( ni34  &  wire29565 ) | ( wire6524  &  wire29565 ) ;
 assign wire6524 = ( ni36  &  (~ wire157)  &  (~ wire29562) ) | ( (~ wire157)  &  (~ nv858)  &  (~ wire29562) ) ;
 assign wire6531 = ( ni34  &  (~ ni29)  &  wire6537 ) | ( ni34  &  (~ ni29)  &  wire29593 ) ;
 assign wire6536 = ( ni40  &  ni36  &  wire388 ) | ( (~ ni40)  &  ni36  &  nv772 ) ;
 assign wire6537 = ( (~ ni36)  &  wire1075 ) | ( (~ ni36)  &  wire6540 ) | ( (~ ni36)  &  wire6541 ) ;
 assign wire6538 = ( (~ ni35)  &  wire604 ) | ( (~ ni35)  &  wire6543 ) ;
 assign wire6540 = ( ni40  &  wire388  &  wire1019 ) | ( (~ ni40)  &  nv772  &  wire1019 ) ;
 assign wire6541 = ( (~ ni35)  &  wire604 ) | ( (~ ni35)  &  wire6543 ) ;
 assign wire6543 = ( ni40  &  wire269  &  wire388 ) | ( (~ ni40)  &  wire269  &  nv772 ) ;
 assign wire6547 = ( pi21  &  ni34  &  wire6557 ) | ( pi21  &  ni34  &  wire29588 ) ;
 assign wire6549 = ( pi21  &  pi22  &  wire6551 ) | ( pi21  &  pi22  &  wire29590 ) ;
 assign wire6551 = ( ni34  &  (~ ni29)  &  wire6557 ) | ( ni34  &  (~ ni29)  &  wire29588 ) ;
 assign wire6556 = ( (~ ni40)  &  ni36  &  nv758 ) | ( ni40  &  ni36  &  wire388 ) ;
 assign wire6557 = ( (~ ni36)  &  wire1075 ) | ( (~ ni36)  &  wire6560 ) | ( (~ ni36)  &  wire6561 ) ;
 assign wire6558 = ( (~ ni35)  &  wire500 ) | ( (~ ni35)  &  wire6563 ) ;
 assign wire6560 = ( (~ ni40)  &  nv758  &  wire1019 ) | ( ni40  &  wire388  &  wire1019 ) ;
 assign wire6561 = ( (~ ni35)  &  wire500 ) | ( (~ ni35)  &  wire6563 ) ;
 assign wire6563 = ( (~ ni40)  &  nv758  &  wire292 ) | ( ni40  &  wire388  &  wire292 ) ;
 assign wire6567 = ( pi21  &  ni34  &  wire6577 ) | ( pi21  &  ni34  &  wire29569 ) ;
 assign wire6569 = ( pi21  &  pi22  &  wire6571 ) | ( pi21  &  pi22  &  wire29572 ) ;
 assign wire6571 = ( ni34  &  (~ ni29)  &  wire6577 ) | ( ni34  &  (~ ni29)  &  wire29569 ) ;
 assign wire6576 = ( ni40  &  ni36  &  nv758 ) | ( (~ ni40)  &  ni36  &  wire388 ) ;
 assign wire6577 = ( (~ ni36)  &  wire1097 ) | ( (~ ni36)  &  wire6580 ) | ( (~ ni36)  &  wire6581 ) ;
 assign wire6578 = ( ni35  &  wire500 ) | ( ni35  &  wire6583 ) ;
 assign wire6580 = ( ni40  &  wire1032  &  nv758 ) | ( (~ ni40)  &  wire1032  &  wire388 ) ;
 assign wire6581 = ( ni35  &  wire500 ) | ( ni35  &  wire6583 ) ;
 assign wire6583 = ( ni40  &  nv758  &  wire292 ) | ( (~ ni40)  &  wire388  &  wire292 ) ;
 assign wire6612 = ( (~ ni40)  &  ni36  &  wire388 ) | ( ni40  &  ni36  &  nv772 ) ;
 assign wire6613 = ( (~ ni36)  &  wire1097 ) | ( (~ ni36)  &  wire6616 ) | ( (~ ni36)  &  wire6617 ) ;
 assign wire6614 = ( ni35  &  wire604 ) | ( ni35  &  wire6619 ) ;
 assign wire6616 = ( (~ ni40)  &  wire1032  &  wire388 ) | ( ni40  &  wire1032  &  nv772 ) ;
 assign wire6617 = ( ni35  &  wire604 ) | ( ni35  &  wire6619 ) ;
 assign wire6619 = ( (~ ni40)  &  wire269  &  wire388 ) | ( ni40  &  wire269  &  nv772 ) ;
 assign wire6626 = ( ni34  &  wire228  &  nv644  &  wire29746 ) ;
 assign wire6628 = ( wire29639  &  wire29751 ) | ( (~ ni29)  &  wire1057  &  wire29751 ) ;
 assign wire6629 = ( ni34  &  wire29753 ) | ( (~ wire785)  &  wire29753 ) ;
 assign wire6630 = ( wire228  &  wire6714  &  wire29754 ) | ( wire228  &  wire29644  &  wire29754 ) ;
 assign wire6633 = ( (~ wire150)  &  nv717  &  wire312  &  wire1058 ) ;
 assign wire6634 = ( wire29655  &  wire29759 ) | ( (~ ni29)  &  wire1092  &  wire29759 ) ;
 assign wire6636 = ( wire6653  &  wire29763 ) | ( wire6655  &  wire29763 ) | ( wire29761  &  wire29763 ) ;
 assign wire6640 = ( wire29662  &  wire29767 ) | ( (~ ni29)  &  wire1012  &  wire29767 ) ;
 assign wire6642 = ( wire1066  &  wire6729 ) | ( wire1066  &  wire6731 ) | ( wire1066  &  wire29768 ) ;
 assign wire6644 = ( (~ pi16)  &  wire6652 ) | ( (~ pi16)  &  wire260  &  wire224 ) ;
 assign wire6647 = ( ni34  &  wire6691  &  wire29624 ) | ( ni34  &  wire29623  &  wire29624 ) ;
 assign wire6652 = ( (~ pi17)  &  (~ pi21)  &  ni34 ) ;
 assign wire6653 = ( pi21  &  ni34  &  wire6663 ) | ( pi21  &  ni34  &  wire29629 ) ;
 assign wire6655 = ( pi21  &  pi22  &  wire6657 ) | ( pi21  &  pi22  &  wire29632 ) ;
 assign wire6657 = ( ni34  &  (~ ni29)  &  wire6663 ) | ( ni34  &  (~ ni29)  &  wire29629 ) ;
 assign wire6662 = ( ni40  &  ni36  &  nv667 ) | ( (~ ni40)  &  ni36  &  nv667 ) | ( ni40  &  ni36  &  nv6576 ) ;
 assign wire6663 = ( (~ ni36)  &  wire1097 ) | ( (~ ni36)  &  wire6666 ) | ( (~ ni36)  &  wire6667 ) ;
 assign wire6664 = ( ni35  &  wire500 ) | ( ni35  &  wire6669 ) ;
 assign wire6666 = ( ni40  &  nv667  &  wire1032 ) | ( (~ ni40)  &  nv667  &  wire1032 ) | ( ni40  &  wire1032  &  nv6576 ) ;
 assign wire6667 = ( ni35  &  wire500 ) | ( ni35  &  wire6669 ) ;
 assign wire6669 = ( ni40  &  nv667  &  wire292 ) | ( (~ ni40)  &  nv667  &  wire292 ) | ( ni40  &  wire292  &  nv6576 ) ;
 assign wire6678 = ( ni35  &  wire604 ) | ( ni35  &  wire6685 ) ;
 assign wire6679 = ( (~ ni40)  &  ni36  &  nv667 ) | ( ni40  &  ni36  &  wire441 ) ;
 assign wire6680 = ( (~ ni36)  &  wire1097 ) | ( (~ ni36)  &  wire6682 ) | ( (~ ni36)  &  wire6683 ) ;
 assign wire6682 = ( (~ ni40)  &  nv667  &  wire1032 ) | ( ni40  &  wire441  &  wire1032 ) ;
 assign wire6683 = ( ni35  &  wire604 ) | ( ni35  &  wire6685 ) ;
 assign wire6685 = ( (~ ni40)  &  nv667  &  wire269 ) | ( ni40  &  wire441  &  wire269 ) ;
 assign wire6691 = ( (~ ni36)  &  wire320 ) | ( (~ ni36)  &  wire6694 ) ;
 assign wire6692 = ( ni42  &  ni36 ) | ( ni36  &  nv669 ) | ( (~ ni42)  &  ni41  &  ni36 ) ;
 assign wire6694 = ( ni42  &  ni38 ) | ( ni38  &  nv669 ) | ( (~ ni42)  &  ni41  &  ni38 ) ;
 assign wire6696 = ( ni34  &  (~ ni29)  &  wire6703 ) | ( ni34  &  (~ ni29)  &  wire29653 ) ;
 assign wire6701 = ( (~ ni35)  &  wire604 ) | ( (~ ni35)  &  wire6708 ) ;
 assign wire6702 = ( ni40  &  ni36  &  nv667 ) | ( (~ ni40)  &  ni36  &  wire441 ) ;
 assign wire6703 = ( (~ ni36)  &  wire1075 ) | ( (~ ni36)  &  wire6705 ) | ( (~ ni36)  &  wire6706 ) ;
 assign wire6705 = ( ni40  &  nv667  &  wire1019 ) | ( (~ ni40)  &  wire441  &  wire1019 ) ;
 assign wire6706 = ( (~ ni35)  &  wire604 ) | ( (~ ni35)  &  wire6708 ) ;
 assign wire6708 = ( ni40  &  nv667  &  wire269 ) | ( (~ ni40)  &  wire441  &  wire269 ) ;
 assign wire6714 = ( ni34  &  (~ ni29)  &  nv644 ) ;
 assign wire6717 = ( (~ ni37)  &  ni36  &  wire441 ) ;
 assign wire6721 = ( (~ ni39)  &  (~ ni38)  &  (~ ni36)  &  nv633 ) ;
 assign wire6722 = ( (~ ni38)  &  ni37  &  (~ ni36) ) | ( ni37  &  (~ ni36)  &  wire441 ) ;
 assign wire6727 = ( (~ ni43)  &  (~ ni42)  &  (~ ni41)  &  ni44 ) ;
 assign wire6729 = ( pi21  &  ni34  &  wire6742 ) | ( pi21  &  ni34  &  wire29648 ) ;
 assign wire6731 = ( pi21  &  pi22  &  wire6736 ) | ( pi21  &  pi22  &  wire29650 ) ;
 assign wire6736 = ( ni34  &  (~ ni29)  &  wire6742 ) | ( ni34  &  (~ ni29)  &  wire29648 ) ;
 assign wire6741 = ( ni40  &  ni36  &  nv667 ) | ( (~ ni40)  &  ni36  &  nv667 ) | ( (~ ni40)  &  ni36  &  nv6576 ) ;
 assign wire6742 = ( (~ ni36)  &  wire1075 ) | ( (~ ni36)  &  wire6745 ) | ( (~ ni36)  &  wire6746 ) ;
 assign wire6743 = ( (~ ni35)  &  wire500 ) | ( (~ ni35)  &  wire6750 ) ;
 assign wire6745 = ( ni40  &  nv667  &  wire1019 ) | ( (~ ni40)  &  nv667  &  wire1019 ) | ( (~ ni40)  &  nv6576  &  wire1019 ) ;
 assign wire6746 = ( (~ ni35)  &  wire500 ) | ( (~ ni35)  &  wire6750 ) ;
 assign wire6750 = ( ni40  &  nv667  &  wire292 ) | ( (~ ni40)  &  nv667  &  wire292 ) | ( (~ ni40)  &  wire292  &  nv6576 ) ;
 assign wire6757 = ( ni32  &  (~ ni31)  &  (~ ni29) ) | ( (~ ni31)  &  ni30  &  (~ ni29) ) ;
 assign wire6758 = ( (~ ni34)  &  (~ ni29) ) ;
 assign wire6766 = ( (~ ni43)  &  (~ ni42)  &  (~ ni41)  &  (~ ni44) ) ;
 assign wire6775 = ( (~ wire290)  &  n_n11282  &  wire29397  &  wire29398 ) ;
 assign wire6780 = ( (~ wire6789)  &  (~ wire6790)  &  wire29414  &  wire29415 ) ;
 assign wire6783 = ( pi23  &  (~ wire290)  &  wire1105  &  n_n13096 ) ;
 assign wire6784 = ( ni35  &  wire768  &  wire29424 ) | ( pi23  &  (~ wire768)  &  wire29424 ) ;
 assign wire6785 = ( ni35  &  wire768  &  wire29425 ) | ( pi23  &  (~ wire768)  &  wire29425 ) ;
 assign wire6786 = ( ni35  &  wire290  &  (~ nv10130) ) | ( ni35  &  wire290  &  (~ wire1289) ) ;
 assign wire6787 = ( (~ ni9)  &  wire29427 ) | ( (~ ni10)  &  wire29427 ) | ( (~ wire1289)  &  wire29427 ) ;
 assign wire6788 = ( ni2  &  ni35 ) | ( ni35  &  ni3 ) | ( ni35  &  wire281 ) ;
 assign wire6789 = ( pi26  &  (~ ni32)  &  (~ ni31)  &  ni30 ) ;
 assign wire6790 = ( pi26  &  ni35 ) ;
 assign wire6795 = ( wire6808  &  wire29179 ) | ( wire6809  &  wire29179 ) ;
 assign wire6796 = ( (~ ni5)  &  (~ nv10252)  &  wire29261 ) | ( (~ nv10252)  &  (~ n_n806)  &  wire29261 ) ;
 assign wire6797 = ( (~ nv10252)  &  (~ wire6811)  &  wire29264 ) | ( (~ wire6811)  &  (~ wire29256)  &  wire29264 ) ;
 assign wire6799 = ( (~ ni5)  &  (~ nv10252)  &  wire29372 ) | ( (~ nv10252)  &  (~ n_n806)  &  wire29372 ) ;
 assign wire6800 = ( (~ ni3)  &  (~ ni6)  &  (~ nv10252)  &  (~ wire6811) ) ;
 assign wire6801 = ( (~ nv10252)  &  (~ wire6811)  &  wire29377 ) | ( (~ wire6811)  &  (~ wire29256)  &  wire29377 ) ;
 assign wire6802 = ( (~ nv10252)  &  (~ wire6811)  &  wire29379 ) | ( (~ wire6811)  &  (~ wire29256)  &  wire29379 ) ;
 assign wire6805 = ( wire29371  &  wire29382 ) | ( (~ ni7)  &  n_n983  &  wire29382 ) ;
 assign wire6808 = ( ni36  &  (~ ni32)  &  ni31  &  ni30 ) ;
 assign wire6809 = ( ni41  &  ni32  &  ni31  &  ni30 ) ;
 assign wire6811 = ( ni5  &  n_n806 ) ;
 assign wire6812 = ( ni6  &  (~ wire399)  &  wire764 ) ;
 assign wire6814 = ( ni6  &  (~ wire399)  &  nv10153 ) ;
 assign wire6815 = ( wire699  &  nv10174  &  wire29181  &  wire29182 ) ;
 assign wire6816 = ( nv10167  &  wire29187  &  wire29188 ) ;
 assign wire6818 = ( wire175  &  nv10167  &  wire29194  &  wire29195 ) ;
 assign wire6819 = ( wire6846  &  wire29204 ) | ( wire6847  &  wire29204 ) | ( wire6848  &  wire29204 ) ;
 assign wire6820 = ( wire6854  &  wire29207 ) | ( wire359  &  nv10173  &  wire29207 ) ;
 assign wire6821 = ( wire6846  &  wire29210 ) | ( wire6847  &  wire29210 ) | ( wire6848  &  wire29210 ) ;
 assign wire6822 = ( wire6842  &  wire29215 ) | ( wire6845  &  wire29215 ) | ( wire29211  &  wire29215 ) ;
 assign wire6824 = ( wire175  &  wire264  &  nv10167  &  wire29219 ) ;
 assign wire6826 = ( wire6838  &  wire29231 ) | ( wire6839  &  wire29231 ) | ( wire29228  &  wire29231 ) ;
 assign wire6827 = ( wire6842  &  wire29233 ) | ( wire6845  &  wire29233 ) | ( wire29211  &  wire29233 ) ;
 assign wire6829 = ( wire175  &  wire264  &  wire331  &  nv10167 ) ;
 assign wire6831 = ( wire6838  &  wire29237 ) | ( wire6839  &  wire29237 ) | ( wire29228  &  wire29237 ) ;
 assign wire6832 = ( wire1328  &  wire6846 ) | ( wire1328  &  wire6847 ) | ( wire1328  &  wire6848 ) ;
 assign wire6833 = ( (~ wire202)  &  wire6838 ) | ( (~ wire202)  &  wire6839 ) | ( (~ wire202)  &  wire29228 ) ;
 assign wire6834 = ( ni9  &  wire6838 ) | ( ni9  &  wire6839 ) | ( ni9  &  wire29228 ) ;
 assign wire6835 = ( pi26  &  (~ wire175)  &  wire264  &  nv10174 ) ;
 assign wire6836 = ( (~ ni30)  &  wire29223 ) | ( ni33  &  ni30  &  wire29223 ) | ( ni31  &  ni30  &  wire29223 ) ;
 assign wire6838 = ( pi27  &  (~ ni14) ) | ( pi26  &  (~ ni14) ) | ( (~ ni14)  &  nv10153 ) ;
 assign wire6839 = ( pi27  &  ni11 ) | ( (~ pi26)  &  ni11 ) | ( ni11  &  nv10153 ) ;
 assign wire6842 = ( n_n450  &  wire1277 ) | ( wire1277  &  wire6847 ) | ( wire1277  &  wire6848 ) ;
 assign wire6844 = ( (~ pi23)  &  (~ pi24)  &  wire6854 ) | ( (~ pi23)  &  (~ pi24)  &  wire6855 ) ;
 assign wire6845 = ( (~ wire160)  &  wire6846 ) | ( (~ wire160)  &  wire6847 ) | ( (~ wire160)  &  wire6848 ) ;
 assign wire6846 = ( wire948  &  wire1277 ) | ( wire1277  &  wire6940 ) | ( wire1277  &  wire29139 ) ;
 assign wire6847 = ( (~ pi24)  &  n_n450 ) | ( (~ pi24)  &  wire6852 ) ;
 assign wire6848 = ( pi24  &  wire6854 ) | ( pi24  &  wire359  &  nv10173 ) ;
 assign wire6852 = ( (~ ni11)  &  nv10153 ) | ( (~ pi27)  &  pi26  &  (~ ni11)  &  (~ nv10153) ) ;
 assign wire6854 = ( (~ pi26)  &  wire377  &  nv10174 ) ;
 assign wire6855 = ( wire359  &  nv10173 ) ;
 assign wire6857 = ( wire480  &  wire29274 ) | ( wire493  &  wire29271  &  wire29274 ) ;
 assign wire6858 = ( wire6898  &  wire29277 ) | ( wire268  &  nv10174  &  wire29277 ) ;
 assign wire6860 = ( (~ pi26)  &  nv10169  &  wire29283 ) | ( pi26  &  nv10173  &  wire29283 ) ;
 assign wire6862 = ( nv10167  &  wire764  &  wire29288 ) ;
 assign wire6864 = ( (~ wire399)  &  wire29296 ) ;
 assign wire6868 = ( wire6906  &  wire29300 ) | ( wire6908  &  wire29300 ) | ( wire29291  &  wire29300 ) ;
 assign wire6869 = ( (~ wire399)  &  nv10153  &  (~ wire574) ) | ( (~ wire155)  &  (~ wire399)  &  (~ nv10153)  &  (~ wire574) ) ;
 assign wire6870 = ( ni13  &  (~ wire399)  &  nv10153 ) ;
 assign wire6871 = ( (~ wire399)  &  wire480 ) ;
 assign wire6873 = ( wire268  &  wire493  &  wire29303 ) ;
 assign wire6874 = ( nv10153  &  wire377  &  wire29306 ) | ( (~ wire156)  &  (~ nv10153)  &  wire377  &  wire29306 ) ;
 assign wire6878 = ( wire480  &  wire29317 ) | ( wire493  &  wire29271  &  wire29317 ) ;
 assign wire6880 = ( wire264  &  wire628  &  wire29320 ) ;
 assign wire6883 = ( ni13  &  (~ wire290)  &  wire628  &  wire29326 ) ;
 assign wire6884 = ( ni13  &  wire509  &  wire628  &  wire29328 ) ;
 assign wire6889 = ( nv10167  &  wire764  &  wire29337 ) ;
 assign wire6890 = ( ni13  &  wire628  &  wire29338 ) ;
 assign wire6891 = ( ni9  &  ni8  &  wire29291 ) | ( ni9  &  ni8  &  wire29292 ) ;
 assign wire6898 = ( pi26  &  nv10169  &  wire377 ) | ( (~ pi26)  &  wire377  &  nv10173 ) ;
 assign wire6899 = ( wire268  &  nv10174 ) ;
 assign wire6906 = ( (~ pi26)  &  nv10169  &  wire29289 ) | ( pi26  &  nv10173  &  wire29289 ) ;
 assign wire6908 = ( pi26  &  nv10169  &  wire377 ) | ( (~ pi26)  &  wire377  &  nv10173 ) ;
 assign wire6909 = ( wire359  &  nv10174 ) ;
 assign wire6923 = ( (~ wire290)  &  (~ wire1122)  &  wire1105  &  wire29153 ) ;
 assign wire6925 = ( ni36  &  wire768  &  wire29159 ) | ( pi24  &  (~ wire768)  &  wire29159 ) ;
 assign wire6926 = ( n_n13895  &  (~ wire1252)  &  (~ wire281)  &  wire29160 ) ;
 assign wire6930 = ( ni36  &  wire768  &  wire29167 ) | ( pi24  &  (~ wire768)  &  wire29167 ) ;
 assign wire6932 = ( ni2  &  ni36 ) | ( ni36  &  ni3 ) | ( ni36  &  wire281 ) ;
 assign wire6935 = ( n_n450  &  wire29097  &  wire29142 ) | ( n_n450  &  wire29098  &  wire29142 ) ;
 assign wire6936 = ( n_n450  &  wire29097  &  wire29145 ) | ( n_n450  &  wire29098  &  wire29145 ) ;
 assign wire6938 = ( ni2  &  ni14 ) | ( ni14  &  ni3 ) ;
 assign wire6940 = ( (~ pi27)  &  pi26  &  (~ ni11) ) ;
 assign wire6945 = ( p__cmndst0p0  &  nv354  &  wire177  &  wire29106 ) ;
 assign wire6946 = ( nv354  &  wire29111 ) ;
 assign wire6949 = ( p__cmndst0p0  &  (~ wire890)  &  wire29117 ) ;
 assign wire6950 = ( (~ ni31)  &  ni30  &  nv444  &  wire29119 ) ;
 assign wire6951 = ( wire29124  &  wire29125 ) | ( nv444  &  wire29122  &  wire29125 ) ;
 assign wire6952 = ( wire6956  &  wire29126 ) | ( wire6959  &  wire29126 ) | ( wire29124  &  wire29126 ) ;
 assign wire6954 = ( (~ wire890)  &  wire6956 ) | ( (~ wire890)  &  wire6959 ) | ( (~ wire890)  &  wire29124 ) ;
 assign wire6955 = ( (~ pi18)  &  wire6959 ) | ( pi17  &  wire6959 ) | ( (~ pi18)  &  wire29124 ) | ( pi17  &  wire29124 ) ;
 assign wire6956 = ( (~ ni32)  &  (~ ni31)  &  ni30  &  nv444 ) ;
 assign wire6959 = ( ni37  &  (~ ni30)  &  nv444 ) ;
 assign wire6965 = ( ni13  &  ni2 ) | ( ni13  &  ni3 ) ;
 assign wire6966 = ( pi27  &  ni14  &  (~ ni11)  &  ni12 ) ;
 assign wire6968 = ( (~ ni13)  &  (~ ni14)  &  (~ ni11) ) ;
 assign wire6969 = ( ni13  &  ni14  &  (~ ni11) ) ;
 assign wire6973 = ( ni13  &  ni11  &  (~ ni12) ) ;
 assign wire6975 = ( ni2  &  ni11 ) | ( ni11  &  ni3 ) ;
 assign wire6976 = ( nv354  &  wire29005  &  wire29006 ) ;
 assign wire6978 = ( nv401  &  wire439  &  wire29012 ) ;
 assign wire6979 = ( nv406  &  wire439  &  wire29015 ) ;
 assign wire6980 = ( nv401  &  wire396  &  wire29018 ) ;
 assign wire6986 = ( wire396  &  wire29037 ) ;
 assign wire6989 = ( nv401  &  wire260  &  wire29042 ) ;
 assign wire6990 = ( pi15  &  ni32  &  nv401  &  wire260 ) ;
 assign wire6991 = ( nv406  &  wire228  &  wire29046 ) ;
 assign wire6992 = ( pi15  &  ni32  &  nv406  &  wire228 ) ;
 assign wire6995 = ( (~ pi17)  &  pi15  &  (~ wire711) ) ;
 assign wire6996 = ( pi17  &  pi15  &  (~ wire711) ) ;
 assign wire6997 = ( (~ pi15)  &  wire7010 ) | ( (~ pi15)  &  wire7011 ) | ( (~ pi15)  &  wire29067 ) ;
 assign wire6999 = ( ni38  &  (~ ni36)  &  ni35  &  (~ ni30) ) ;
 assign wire7000 = ( ni38  &  (~ ni36)  &  ni35  &  ni32 ) ;
 assign wire7008 = ( nv354  &  wire319  &  wire616 ) ;
 assign wire7009 = ( nv363  &  wire319  &  wire381 ) ;
 assign wire7010 = ( ni32  &  nv354  &  wire260 ) | ( (~ ni30)  &  nv354  &  wire260 ) ;
 assign wire7011 = ( ni32  &  nv363  &  wire228 ) | ( (~ ni30)  &  nv363  &  wire228 ) ;
 assign wire7025 = ( ni48  &  ni32  &  ni31  &  (~ ni30) ) ;
 assign wire7027 = ( pi22  &  ni48 ) ;
 assign wire7028 = ( ni44  &  (~ ni32) ) | ( ni44  &  (~ ni30) ) | ( ni44  &  ni31  &  ni30 ) ;
 assign wire7029 = ( ni33  &  ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire7030 = ( ni45  &  wire425 ) | ( wire425  &  wire1002 ) | ( ni45  &  wire239 ) | ( wire1002  &  wire239 ) ;
 assign wire7031 = ( ni45  &  (~ ni31) ) | ( ni45  &  ni31  &  ni30 ) ;
 assign wire7032 = ( ni45  &  ni32 ) ;
 assign wire7035 = ( pi20  &  (~ ni45)  &  wire1002 ) ;
 assign wire7042 = ( (~ pi22)  &  ni30  &  (~ wire425)  &  (~ wire239) ) ;
 assign wire7043 = ( ni47  &  wire425 ) | ( ni47  &  wire239 ) | ( wire425  &  wire7044 ) | ( wire239  &  wire7044 ) ;
 assign wire7044 = ( (~ pi22)  &  (~ ni32) ) | ( (~ pi22)  &  (~ ni31) ) | ( (~ pi22)  &  ni30 ) ;
 assign wire7049 = ( (~ wire290)  &  nv10130  &  wire1026  &  wire28959 ) ;
 assign wire7055 = ( wire7058  &  wire28977 ) | ( wire7059  &  wire28977 ) | ( wire28974  &  wire28977 ) ;
 assign wire7056 = ( wire7058  &  wire28978 ) | ( wire7059  &  wire28978 ) | ( wire28974  &  wire28978 ) ;
 assign wire7057 = ( ni40  &  ni2 ) | ( ni40  &  ni3 ) | ( ni40  &  wire281 ) ;
 assign wire7058 = ( (~ wire290)  &  (~ nv10153)  &  wire28971 ) ;
 assign wire7059 = ( ni40  &  wire290 ) | ( ni40  &  nv6428 ) ;
 assign wire7060 = ( ni40  &  (~ ni33) ) | ( ni40  &  (~ ni30) ) ;
 assign wire7070 = ( (~ wire290)  &  nv10130  &  wire1026  &  wire28924 ) ;
 assign wire7072 = ( pi24  &  (~ wire290)  &  nv10130  &  wire28929 ) ;
 assign wire7077 = ( ni41  &  ni2 ) | ( ni41  &  ni3 ) | ( ni41  &  wire281 ) ;
 assign wire7080 = ( wire318  &  wire28775 ) | ( wire7144  &  wire28775 ) ;
 assign wire7087 = ( (~ pi18)  &  (~ pi16)  &  nv158  &  wire28798 ) ;
 assign wire7088 = ( n_n13646  &  wire318  &  wire28800 ) | ( n_n13646  &  wire7144  &  wire28800 ) ;
 assign wire7089 = ( (~ ni38)  &  (~ ni37)  &  nv158  &  wire28802 ) ;
 assign wire7090 = ( pi18  &  (~ pi17)  &  pi16  &  wire1264 ) ;
 assign wire7091 = ( wire7109  &  wire28849 ) | ( wire28846  &  wire28849 ) | ( wire28848  &  wire28849 ) ;
 assign wire7093 = ( (~ pi18)  &  pi16  &  wire7140 ) | ( (~ pi18)  &  pi16  &  wire28852 ) ;
 assign wire7095 = ( wire302  &  wire7122 ) | ( wire302  &  wire7123 ) | ( wire302  &  wire28892 ) ;
 assign wire7096 = ( pi17  &  pi16  &  wire7140 ) | ( pi17  &  pi16  &  wire28852 ) ;
 assign wire7097 = ( (~ wire1126)  &  (~ wire722)  &  wire28805 ) ;
 assign wire7099 = ( (~ nv235)  &  (~ wire1126)  &  wire28812 ) ;
 assign wire7100 = ( pi20  &  (~ ni30)  &  (~ wire722)  &  wire28815 ) ;
 assign wire7101 = ( pi20  &  (~ ni30)  &  n_n13546  &  wire28818 ) ;
 assign wire7107 = ( (~ wire1126)  &  (~ wire722)  &  wire28831 ) ;
 assign wire7109 = ( ni38  &  (~ ni30)  &  (~ nv222) ) | ( ni37  &  (~ ni30)  &  (~ nv222) ) ;
 assign wire7118 = ( n_n13546  &  (~ wire1126)  &  wire28854  &  wire28855 ) ;
 assign wire7119 = ( n_n13566  &  (~ wire1126)  &  wire28858  &  wire28859 ) ;
 assign wire7120 = ( pi18  &  ni41  &  nv158  &  wire28863 ) ;
 assign wire7121 = ( pi18  &  (~ ni30)  &  nv158  &  wire1126 ) ;
 assign wire7122 = ( (~ wire851)  &  (~ wire7126)  &  (~ wire28875)  &  wire28878 ) ;
 assign wire7123 = ( (~ wire28885)  &  (~ wire28886)  &  wire28888 ) ;
 assign wire7126 = ( ni39  &  (~ nv78)  &  (~ n_n13755)  &  nv116 ) ;
 assign wire7129 = ( ni39  &  (~ nv69)  &  nv121  &  (~ n_n13755) ) ;
 assign wire7134 = ( ni39  &  (~ ni43)  &  ni42 ) | ( ni39  &  ni42  &  ni44 ) ;
 assign wire7140 = ( (~ nv212)  &  wire318 ) | ( (~ nv212)  &  wire7144 ) ;
 assign wire7144 = ( ni38  &  (~ ni30) ) | ( ni37  &  (~ ni30) ) ;
 assign wire7169 = ( (~ nv69)  &  (~ n_n13755)  &  wire28721 ) ;
 assign wire7170 = ( (~ nv78)  &  (~ n_n13755)  &  wire28724 ) ;
 assign wire7172 = ( (~ ni32)  &  (~ nv69)  &  wire260 ) | ( (~ ni30)  &  (~ nv69)  &  wire260 ) ;
 assign wire7173 = ( (~ ni32)  &  (~ nv78)  &  wire228 ) | ( (~ ni30)  &  (~ nv78)  &  wire228 ) ;
 assign wire7174 = ( (~ pi17)  &  ni32  &  ni31  &  ni30 ) ;
 assign wire7175 = ( wire839  &  (~ nv116)  &  wire28695 ) ;
 assign wire7176 = ( wire839  &  (~ nv121)  &  wire28698 ) ;
 assign wire7180 = ( wire260  &  (~ nv116)  &  wire28706 ) ;
 assign wire7181 = ( wire228  &  (~ nv121)  &  wire28708 ) ;
 assign wire7184 = ( pi16  &  ni32  &  ni31  &  ni30 ) ;
 assign wire7193 = ( ni39  &  ni32 ) | ( ni39  &  ni31 ) | ( ni39  &  (~ ni32)  &  (~ ni30) ) ;
 assign wire7194 = ( ni33  &  (~ ni32)  &  (~ ni31)  &  ni30 ) ;
 assign wire7195 = ( (~ ni32)  &  (~ ni30) ) ;
 assign wire28695 = ( (~ pi17)  &  (~ pi20)  &  pi16 ) ;
 assign wire28698 = ( (~ pi17)  &  pi20  &  pi16 ) ;
 assign wire28700 = ( (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire28702 = ( (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire28705 = ( (~ pi17)  &  pi19  &  pi16  &  (~ ni43) ) ;
 assign wire28706 = ( pi16  &  (~ ni32) ) | ( pi16  &  (~ ni30) ) ;
 assign wire28708 = ( pi16  &  (~ ni32) ) | ( pi16  &  (~ ni30) ) ;
 assign wire28710 = ( pi17  &  pi16  &  (~ ni43) ) ;
 assign wire28711 = ( (~ ni43)  &  (~ ni32) ) | ( (~ ni43)  &  (~ ni30) ) ;
 assign wire28712 = ( (~ ni40)  &  (~ n_n9245)  &  wire28705 ) | ( ni40  &  (~ n_n9245)  &  wire28710 ) ;
 assign wire28713 = ( wire7184 ) | ( wire257  &  wire28711 ) ;
 assign wire28715 = ( wire7176 ) | ( wire829  &  (~ nv121)  &  wire28702 ) ;
 assign wire28716 = ( wire7181 ) | ( wire28712 ) | ( wire28713 ) ;
 assign wire28718 = ( wire7175 ) | ( wire829  &  (~ nv116)  &  wire28700 ) ;
 assign wire28721 = ( (~ pi17)  &  (~ pi20)  &  (~ ni32) ) | ( (~ pi17)  &  (~ pi20)  &  (~ ni30) ) ;
 assign wire28724 = ( (~ pi17)  &  pi20  &  (~ ni32) ) | ( (~ pi17)  &  pi20  &  (~ ni30) ) ;
 assign wire28729 = ( wire7174 ) | ( wire829  &  wire191  &  (~ n_n13755) ) ;
 assign wire28731 = ( wire7169 ) | ( wire7172 ) | ( wire28729 ) ;
 assign wire28734 = ( (~ ni40)  &  (~ ni32) ) | ( (~ ni40)  &  (~ ni31) ) | ( (~ ni40)  &  (~ ni30) ) | ( ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire28735 = ( pi17  &  (~ pi19)  &  (~ wire829)  &  wire28734 ) ;
 assign wire28739 = ( nv78  &  wire282  &  (~ wire839)  &  (~ wire911) ) ;
 assign wire28743 = ( nv69  &  wire326  &  (~ wire839)  &  (~ wire911) ) ;
 assign wire28746 = ( ni40  &  (~ ni32) ) | ( ni40  &  (~ ni31) ) | ( ni40  &  (~ ni30) ) | ( ni32  &  (~ ni31)  &  ni30 ) ;
 assign wire28747 = ( pi17  &  (~ pi19)  &  (~ wire514)  &  wire28746 ) ;
 assign wire28751 = ( nv78  &  wire282  &  (~ wire514)  &  (~ wire911) ) ;
 assign wire28755 = ( nv69  &  wire326  &  (~ wire514)  &  (~ wire911) ) ;
 assign wire28757 = ( (~ pi17)  &  (~ ni32) ) | ( pi19  &  (~ ni32) ) | ( (~ pi17)  &  (~ ni30) ) | ( pi19  &  (~ ni30) ) ;
 assign wire28758 = ( ni43  &  ni42  &  wire28757 ) | ( ni43  &  (~ ni41)  &  wire28757 ) ;
 assign wire28760 = ( (~ pi17)  &  (~ wire1153) ) | ( pi19  &  (~ wire1153) ) ;
 assign wire28763 = ( pi16  &  (~ n_n13789) ) | ( (~ n_n13789)  &  (~ n_n13786)  &  wire28735 ) ;
 assign wire28764 = ( (~ n_n13789)  &  (~ n_n13786)  &  wire28739 ) | ( (~ n_n13789)  &  (~ n_n13786)  &  wire28743 ) ;
 assign wire28765 = ( (~ n_n13789)  &  (~ n_n13786)  &  wire28747 ) | ( (~ n_n13789)  &  (~ n_n13786)  &  wire28751 ) ;
 assign wire28766 = ( (~ n_n13789)  &  (~ n_n13786)  &  wire28755 ) | ( (~ n_n13789)  &  (~ n_n13786)  &  wire28758 ) ;
 assign wire28767 = ( wire302  &  (~ n_n13789)  &  (~ n_n13786) ) | ( (~ n_n13789)  &  (~ n_n13786)  &  wire28760 ) ;
 assign wire28770 = ( wire28763 ) | ( wire28764 ) | ( wire28767 ) ;
 assign wire28771 = ( ni38  &  ni32 ) | ( ni37  &  ni32 ) ;
 assign wire28773 = ( ni39  &  ni42 ) | ( ni39  &  (~ ni41) ) ;
 assign wire28775 = ( (~ pi18)  &  (~ pi16)  &  (~ nv212)  &  wire28773 ) ;
 assign wire28777 = ( ni39  &  (~ ni43)  &  (~ ni42) ) ;
 assign wire28779 = ( (~ pi18)  &  (~ pi16)  &  (~ nv212)  &  wire28777 ) ;
 assign wire28781 = ( (~ pi18)  &  (~ pi16)  &  (~ ni39) ) ;
 assign wire28783 = ( (~ n_n13541)  &  (~ nv212)  &  wire28781 ) ;
 assign wire28784 = ( pi17  &  (~ pi16)  &  ni39 ) ;
 assign wire28786 = ( ni42  &  (~ nv212)  &  wire28784 ) | ( (~ ni41)  &  (~ nv212)  &  wire28784 ) ;
 assign wire28787 = ( ni39  &  (~ ni43)  &  (~ ni42) ) ;
 assign wire28789 = ( pi17  &  (~ pi16)  &  (~ nv212)  &  wire28787 ) ;
 assign wire28790 = ( pi17  &  (~ pi16)  &  (~ ni39) ) ;
 assign wire28792 = ( (~ n_n13541)  &  (~ nv212)  &  wire28790 ) ;
 assign wire28796 = ( (~ pi18)  &  (~ pi16)  &  (~ ni39)  &  n_n13646 ) ;
 assign wire28798 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28800 = ( pi17  &  (~ pi16)  &  (~ ni39) ) ;
 assign wire28802 = ( pi17  &  (~ pi16)  &  (~ ni30) ) ;
 assign wire28805 = ( pi20  &  (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28808 = ( pi20  &  (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28812 = ( pi20  &  ni38  &  (~ ni30) ) | ( pi20  &  ni37  &  (~ ni30) ) ;
 assign wire28815 = ( ni43  &  (~ ni38)  &  (~ ni37) ) | ( (~ ni42)  &  (~ ni38)  &  (~ ni37) ) ;
 assign wire28818 = ( ni43  &  (~ ni38)  &  (~ ni37) ) | ( (~ ni42)  &  (~ ni38)  &  (~ ni37) ) ;
 assign wire28821 = ( ni43  &  ni38 ) | ( (~ ni42)  &  ni38 ) | ( ni43  &  ni37 ) | ( (~ ni42)  &  ni37 ) ;
 assign wire28822 = ( pi20  &  (~ ni30)  &  wire28821 ) ;
 assign wire28825 = ( wire1037 ) | ( n_n13546  &  (~ wire1126)  &  wire28808 ) ;
 assign wire28826 = ( wire7097 ) | ( wire7100 ) | ( wire7101 ) ;
 assign wire28829 = ( (~ nv235)  &  wire28822 ) | ( pi20  &  wire318  &  (~ nv235) ) ;
 assign wire28831 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28834 = ( ni40  &  (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28838 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28839 = ( ni43  &  ni41 ) | ( (~ ni42)  &  ni41 ) | ( ni43  &  (~ ni40) ) | ( (~ ni42)  &  (~ ni40) ) ;
 assign wire28840 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28842 = ( ni38  &  (~ ni30) ) | ( ni37  &  (~ ni30) ) ;
 assign wire28845 = ( n_n13566  &  wire28834 ) | ( n_n13566  &  wire419  &  wire28840 ) ;
 assign wire28846 = ( wire7107 ) | ( wire28845 ) | ( wire28838  &  wire28839 ) ;
 assign wire28848 = ( wire318  &  (~ nv222) ) | ( wire419  &  (~ nv222)  &  wire28842 ) ;
 assign wire28849 = ( pi18  &  (~ pi17)  &  (~ pi20)  &  pi16 ) ;
 assign wire28850 = ( (~ pi16)  &  (~ pi18) ) ;
 assign wire28851 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28852 = ( wire1037 ) | ( ni43  &  wire28851 ) | ( (~ ni42)  &  wire28851 ) ;
 assign wire28854 = ( pi20  &  pi18 ) ;
 assign wire28855 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28858 = ( (~ pi20)  &  pi18 ) ;
 assign wire28859 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28863 = ( (~ ni38)  &  (~ ni37)  &  (~ ni30) ) ;
 assign wire28868 = ( (~ ni40)  &  (~ ni39) ) ;
 assign wire28870 = ( (~ ni39)  &  (~ n_n13646)  &  (~ n_n13546) ) ;
 assign wire28873 = ( (~ ni39)  &  (~ ni43)  &  ni42 ) | ( (~ ni39)  &  ni42  &  (~ ni44) ) ;
 assign wire28875 = ( (~ n_n13600)  &  wire28870 ) | ( (~ n_n13646)  &  (~ n_n13600)  &  wire28873 ) ;
 assign wire28878 = ( pi18  &  pi20  &  wire318 ) | ( pi18  &  pi20  &  wire7144 ) ;
 assign wire28882 = ( (~ ni39)  &  (~ n_n13646)  &  (~ n_n13566) ) ;
 assign wire28883 = ( (~ ni39)  &  ni42  &  (~ ni44) ) | ( ni39  &  (~ ni43)  &  ni42  &  ni44 ) ;
 assign wire28885 = ( (~ n_n13600)  &  wire28882 ) | ( (~ n_n13646)  &  (~ n_n13600)  &  wire28883 ) ;
 assign wire28886 = ( wire7129 ) | ( wire7134 ) | ( (~ n_n13600)  &  wire28868 ) ;
 assign wire28888 = ( pi18  &  (~ pi20)  &  wire318 ) | ( pi18  &  (~ pi20)  &  wire7144 ) ;
 assign wire28891 = ( wire7120 ) | ( wire7121 ) | ( pi18  &  wire1037 ) ;
 assign wire28892 = ( wire7118 ) | ( wire7119 ) | ( wire28891 ) ;
 assign wire28895 = ( wire7087 ) | ( wire7089 ) | ( wire1037  &  wire28850 ) ;
 assign wire28897 = ( wire318  &  wire28779 ) | ( wire7144  &  wire28779 ) | ( wire318  &  wire28783 ) | ( wire7144  &  wire28783 ) ;
 assign wire28898 = ( wire318  &  wire28786 ) | ( wire7144  &  wire28786 ) | ( wire318  &  wire28789 ) | ( wire7144  &  wire28789 ) ;
 assign wire28899 = ( wire318  &  wire28792 ) | ( wire7144  &  wire28792 ) | ( wire318  &  wire28796 ) | ( wire7144  &  wire28796 ) ;
 assign wire28901 = ( wire7080 ) | ( wire28897 ) | ( wire158  &  wire1037 ) ;
 assign wire28902 = ( wire28899 ) | ( wire28898 ) ;
 assign wire28905 = ( wire7088 ) | ( wire7093 ) | ( wire28895 ) | ( wire28902 ) ;
 assign wire28906 = ( wire7091 ) | ( wire7096 ) | ( wire28901 ) ;
 assign wire28910 = ( pi24  &  ni9  &  (~ ni33)  &  ni10 ) ;
 assign wire28912 = ( wire290  &  (~ wire466)  &  wire28910 ) ;
 assign wire28913 = ( ni41  &  pi24 ) ;
 assign wire28914 = ( ni9  &  ni10  &  (~ wire290)  &  wire28913 ) ;
 assign wire28917 = ( (~ pi24)  &  ni41  &  (~ ni32) ) | ( (~ pi24)  &  ni41  &  (~ ni30) ) ;
 assign wire28918 = ( ni9  &  ni10  &  (~ wire290)  &  wire28917 ) ;
 assign wire28919 = ( ni41  &  ni9  &  ni10 ) ;
 assign wire28921 = ( wire290  &  wire466  &  wire28919 ) ;
 assign wire28922 = ( ni9  &  ni10  &  (~ wire290)  &  wire1299 ) ;
 assign wire28923 = ( n_n13895  &  (~ wire638)  &  (~ wire281)  &  (~ wire202) ) ;
 assign wire28924 = ( pi27  &  pi24  &  (~ wire466) ) ;
 assign wire28926 = ( pi27  &  pi24  &  ni41 ) ;
 assign wire28927 = ( ni9  &  ni10  &  (~ wire290)  &  wire28926 ) ;
 assign wire28929 = ( n_n13895  &  (~ wire988)  &  (~ wire281)  &  (~ wire202) ) ;
 assign wire28930 = ( ni41  &  ni31 ) | ( ni41  &  (~ ni32)  &  (~ ni30) ) ;
 assign wire28931 = ( ni9  &  ni10  &  (~ wire290)  &  wire28930 ) ;
 assign wire28933 = ( ni9  &  ni10  &  wire290  &  n_n434 ) ;
 assign wire28934 = ( ni9  &  (~ ni10) ) ;
 assign wire28935 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire28934 ) ;
 assign wire28936 = ( (~ ni2)  &  (~ ni3)  &  wire792  &  (~ wire281) ) ;
 assign wire28937 = ( wire7077 ) | ( wire1026  &  wire28912 ) ;
 assign wire28938 = ( wire1026  &  wire28918 ) | ( wire1026  &  wire28921 ) ;
 assign wire28939 = ( wire1026  &  wire28927 ) | ( wire1026  &  wire28931 ) ;
 assign wire28940 = ( wire1026  &  wire28933 ) | ( wire638  &  wire1026  &  wire28914 ) ;
 assign wire28944 = ( wire7070 ) | ( wire28940 ) | ( wire28922  &  wire28923 ) ;
 assign wire28945 = ( wire7072 ) | ( wire28937 ) | ( wire28938 ) | ( wire28939 ) ;
 assign wire28946 = ( nv251  &  wire28935 ) | ( nv251  &  wire28936 ) ;
 assign wire28949 = ( pi23  &  ni9  &  (~ ni33)  &  ni10 ) ;
 assign wire28951 = ( wire290  &  (~ wire466)  &  wire28949 ) ;
 assign wire28952 = ( ni40  &  ni9  &  ni10 ) ;
 assign wire28954 = ( wire290  &  wire988  &  wire28952 ) ;
 assign wire28955 = ( (~ pi23)  &  pi26 ) ;
 assign wire28956 = ( ni9  &  ni10  &  (~ wire290)  &  wire28955 ) ;
 assign wire28959 = ( (~ pi23)  &  ni40  &  wire466 ) ;
 assign wire28961 = ( pi23  &  ni9  &  ni10  &  (~ wire290) ) ;
 assign wire28962 = ( n_n13895  &  (~ wire988)  &  (~ wire281)  &  (~ wire202) ) ;
 assign wire28963 = ( ni40  &  (~ ni32) ) | ( ni40  &  (~ ni33)  &  (~ ni30) ) ;
 assign wire28964 = ( ni9  &  ni10  &  (~ wire290)  &  wire28963 ) ;
 assign wire28965 = ( pi26  &  ni40  &  (~ ni32) ) | ( pi26  &  ni40  &  (~ ni30) ) ;
 assign wire28966 = ( ni9  &  ni10  &  (~ wire290)  &  wire28965 ) ;
 assign wire28967 = ( pi26  &  pi23  &  (~ wire466) ) ;
 assign wire28969 = ( ni40  &  ni31 ) | ( ni40  &  (~ ni30) ) ;
 assign wire28971 = ( pi26  &  ni32  &  ni30 ) ;
 assign wire28974 = ( wire7060 ) | ( pi26  &  ni40 ) | ( ni40  &  (~ ni32) ) ;
 assign wire28976 = ( ni9  &  (~ ni10) ) ;
 assign wire28977 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire28976 ) ;
 assign wire28978 = ( (~ ni2)  &  (~ ni3)  &  wire792  &  (~ wire281) ) ;
 assign wire28979 = ( wire7057 ) | ( wire1026  &  wire28951 ) ;
 assign wire28980 = ( wire1026  &  wire28964 ) | ( wire1026  &  wire28966 ) ;
 assign wire28981 = ( wire1026  &  wire28954 ) | ( (~ wire638)  &  wire1026  &  wire28956 ) ;
 assign wire28983 = ( wire594  &  wire1026  &  wire28967 ) | ( wire594  &  wire1026  &  wire28969 ) ;
 assign wire28986 = ( wire7049 ) | ( wire28981 ) | ( wire28961  &  wire28962 ) ;
 assign wire28987 = ( wire28979 ) | ( wire28980 ) | ( wire28983 ) ;
 assign wire28989 = ( ni47  &  (~ ni32) ) | ( ni47  &  (~ ni31) ) | ( ni47  &  ni30 ) ;
 assign wire28990 = ( (~ pi22)  &  (~ ni32) ) | ( (~ pi22)  &  (~ ni31) ) ;
 assign wire28991 = ( (~ wire425)  &  (~ wire239)  &  wire28989 ) | ( (~ wire425)  &  (~ wire239)  &  wire28990 ) ;
 assign wire28995 = ( pi21  &  ni46 ) | ( ni46  &  (~ ni32)  &  (~ wire856) ) ;
 assign wire28999 = ( ni48  &  ni47 ) ;
 assign wire29003 = ( wire7025 ) | ( wire7027 ) | ( wire218  &  wire28999 ) ;
 assign wire29005 = ( (~ ni35)  &  ni32 ) | ( (~ ni35)  &  (~ ni30) ) ;
 assign wire29006 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi15) ) ;
 assign wire29009 = ( (~ pi15)  &  (~ ni35)  &  ni32 ) | ( (~ pi15)  &  (~ ni35)  &  (~ ni30) ) ;
 assign wire29012 = ( (~ pi17)  &  (~ pi20)  &  pi15 ) ;
 assign wire29015 = ( (~ pi17)  &  pi20  &  pi15 ) ;
 assign wire29018 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi15 ) ;
 assign wire29021 = ( (~ ni36)  &  ni32 ) | ( (~ ni36)  &  (~ ni30) ) ;
 assign wire29022 = ( pi17  &  pi19  &  (~ pi15)  &  ni38 ) ;
 assign wire29023 = ( ni38  &  ni37  &  ni36 ) ;
 assign wire29026 = ( wire6999 ) | ( (~ ni32)  &  (~ ni31)  &  ni30 ) ;
 assign wire29027 = ( wire7000 ) | ( wire319  &  wire29023 ) ;
 assign wire29029 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi15) ) ;
 assign wire29030 = ( pi17  &  (~ pi19)  &  pi20  &  pi15 ) ;
 assign wire29033 = ( pi17  &  pi15  &  ni38 ) ;
 assign wire29035 = ( pi17  &  pi19  &  (~ pi15)  &  ni38 ) ;
 assign wire29037 = ( (~ pi17)  &  pi19  &  pi15  &  ni38 ) ;
 assign wire29038 = ( ni38  &  pi15 ) ;
 assign wire29039 = ( pi17  &  pi19  &  (~ ni31) ) | ( pi17  &  pi19  &  (~ ni30) ) ;
 assign wire29040 = ( ni38  &  pi15 ) ;
 assign wire29041 = ( pi17  &  pi19  &  ni32 ) ;
 assign wire29042 = ( pi15  &  (~ ni31) ) | ( pi15  &  (~ ni30) ) ;
 assign wire29046 = ( pi15  &  (~ ni31) ) | ( pi15  &  (~ ni30) ) ;
 assign wire29050 = ( pi17  &  pi19  &  (~ pi15) ) ;
 assign wire29051 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi15) ) ;
 assign wire29054 = ( ni38  &  ni32 ) | ( ni38  &  (~ ni30) ) ;
 assign wire29057 = ( (~ pi17)  &  pi19  &  ni38  &  (~ ni35) ) ;
 assign wire29062 = ( wire191  &  wire1086 ) | ( wire191  &  (~ wire1019)  &  wire29054 ) ;
 assign wire29063 = ( wire1086  &  wire340 ) | ( wire412  &  wire29057 ) ;
 assign wire29067 = ( wire7008 ) | ( wire7009 ) | ( wire29062 ) | ( wire29063 ) ;
 assign wire29068 = ( wire29021  &  wire29022 ) | ( wire29038  &  wire29039 ) ;
 assign wire29069 = ( wire29040  &  wire29041 ) | ( wire1086  &  wire29050 ) ;
 assign wire29070 = ( wire439  &  wire29033 ) | ( wire412  &  wire29035 ) ;
 assign wire29077 = ( wire29070 ) | ( nv406  &  wire396  &  wire29030 ) ;
 assign wire29078 = ( wire6986 ) | ( wire6989 ) | ( wire6990 ) | ( wire6991 ) ;
 assign wire29079 = ( wire6992 ) | ( wire6995 ) | ( wire6996 ) | ( wire29068 ) ;
 assign wire29080 = ( wire6976 ) | ( nv363  &  wire458  &  wire29009 ) ;
 assign wire29081 = ( wire29026  &  wire29029 ) | ( wire29027  &  wire29029 ) | ( wire29026  &  wire29051 ) | ( wire29027  &  wire29051 ) ;
 assign wire29082 = ( wire6978 ) | ( wire6979 ) | ( wire6980 ) | ( wire29069 ) ;
 assign wire29086 = ( wire29077 ) | ( wire29078 ) | ( wire29079 ) | ( wire29080 ) ;
 assign wire29088 = ( ni13  &  (~ ni2)  &  ni14  &  (~ ni3) ) ;
 assign wire29089 = ( (~ ni13)  &  ni11 ) | ( (~ ni14)  &  ni11 ) ;
 assign wire29092 = ( (~ ni14)  &  ni11 ) | ( (~ ni13)  &  ni11  &  ni12 ) ;
 assign wire29094 = ( wire190  &  wire29088 ) | ( wire155  &  wire29089 ) ;
 assign wire29095 = ( wire6973 ) | ( wire6975 ) | ( wire29092 ) ;
 assign wire29097 = ( wire6966 ) | ( (~ ni13)  &  (~ ni14)  &  (~ ni11) ) ;
 assign wire29098 = ( wire6969 ) | ( (~ ni33)  &  (~ wire631) ) | ( (~ ni29)  &  (~ wire631) ) ;
 assign wire29099 = ( (~ ni13)  &  (~ ni2)  &  ni14  &  (~ ni3) ) ;
 assign wire29100 = ( wire29094  &  wire29099 ) | ( wire29095  &  wire29099 ) ;
 assign wire29101 = ( (~ ni2)  &  (~ ni11)  &  (~ ni3) ) ;
 assign wire29102 = ( wire6965 ) | ( (~ wire29097)  &  (~ wire29098)  &  wire29101 ) ;
 assign wire29106 = ( pi18  &  (~ pi17)  &  pi20  &  (~ pi15) ) ;
 assign wire29108 = ( pi15  &  ni38  &  (~ ni37) ) ;
 assign wire29111 = ( pi20  &  (~ wire262)  &  wire319  &  wire29108 ) ;
 assign wire29113 = ( pi15  &  (~ ni32)  &  (~ ni31)  &  ni30 ) ;
 assign wire29115 = ( (~ ni38)  &  (~ ni36)  &  ni35 ) ;
 assign wire29117 = ( (~ ni39)  &  (~ ni36)  &  ni35 ) ;
 assign wire29119 = ( (~ pi18)  &  (~ ni32) ) | ( pi17  &  (~ ni32) ) ;
 assign wire29121 = ( ni37  &  ni32  &  ni30 ) ;
 assign wire29122 = ( (~ ni30)  &  ni37 ) ;
 assign wire29123 = ( (~ ni38)  &  ni37  &  (~ ni30) ) | ( (~ ni38)  &  ni37  &  ni32  &  ni30 ) ;
 assign wire29124 = ( wire29123 ) | ( ni39  &  ni44  &  wire29121 ) | ( (~ ni39)  &  (~ ni44)  &  wire29121 ) ;
 assign wire29125 = ( (~ pi18)  &  pi15 ) | ( pi17  &  pi15 ) | ( pi20  &  pi15 ) ;
 assign wire29126 = ( pi18  &  (~ pi17)  &  (~ pi15) ) ;
 assign wire29127 = ( ni36  &  (~ pi15) ) ;
 assign wire29128 = ( p__cmndst0p0  &  wire29127 ) | ( p__cmndst0p0  &  (~ wire890)  &  wire29115 ) ;
 assign wire29130 = ( wire29128 ) | ( nv444  &  wire890  &  wire29113 ) ;
 assign wire29131 = ( wire6945 ) | ( wire6949 ) | ( wire6950 ) ;
 assign wire29136 = ( wire6952 ) | ( wire6954 ) | ( wire6955 ) | ( wire29130 ) ;
 assign wire29139 = ( ni13  &  (~ ni11) ) | ( pi27  &  (~ ni14)  &  (~ ni11) ) ;
 assign wire29142 = ( (~ ni13)  &  (~ ni2)  &  ni14  &  (~ ni3) ) ;
 assign wire29144 = ( (~ ni2)  &  ni12  &  (~ ni3) ) ;
 assign wire29145 = ( (~ ni13)  &  wire29144 ) | ( (~ ni14)  &  wire29144 ) ;
 assign wire29148 = ( (~ ni2)  &  (~ ni14)  &  (~ ni3) ) ;
 assign wire29149 = ( wire6938 ) | ( (~ wire29097)  &  (~ wire29098)  &  wire29148 ) ;
 assign wire29151 = ( pi24  &  (~ ni33)  &  (~ ni32) ) ;
 assign wire29153 = ( (~ ni31)  &  ni30  &  wire29151 ) ;
 assign wire29155 = ( pi27  &  (~ pi24)  &  ni33  &  (~ ni32) ) ;
 assign wire29157 = ( (~ ni31)  &  ni30  &  (~ wire290)  &  wire29155 ) ;
 assign wire29158 = ( ni13  &  (~ ni14)  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire29159 = ( nv10130  &  wire1289  &  (~ wire281)  &  wire29158 ) ;
 assign wire29160 = ( pi27  &  (~ ni9) ) | ( pi27  &  (~ ni10) ) | ( pi27  &  (~ wire1289) ) ;
 assign wire29163 = ( pi27  &  pi24  &  (~ wire290)  &  (~ wire711) ) ;
 assign wire29165 = ( ni36  &  (~ wire290)  &  nv6428 ) ;
 assign wire29166 = ( ni36  &  (~ ni9) ) | ( ni36  &  (~ ni10) ) | ( ni36  &  (~ wire1289) ) ;
 assign wire29167 = ( nv10130  &  wire1289  &  wire630  &  (~ wire281) ) ;
 assign wire29168 = ( ni36  &  ni32  &  (~ wire290) ) ;
 assign wire29169 = ( wire6932 ) | ( wire1105  &  wire29157 ) ;
 assign wire29170 = ( wire1105  &  wire29163 ) | ( wire1105  &  wire29165 ) ;
 assign wire29171 = ( wire1252  &  wire29166 ) | ( wire1105  &  wire29168 ) ;
 assign wire29176 = ( wire6926 ) | ( wire6930 ) | ( wire29169 ) | ( wire29170 ) ;
 assign wire29179 = ( ni4  &  ni3  &  (~ ni5)  &  ni6 ) ;
 assign wire29181 = ( (~ pi23)  &  (~ pi24)  &  (~ ni10) ) ;
 assign wire29182 = ( pi26  &  (~ ni9)  &  (~ ni7)  &  ni8 ) ;
 assign wire29187 = ( (~ pi23)  &  (~ pi24)  &  (~ ni7)  &  ni8 ) ;
 assign wire29188 = ( (~ pi26)  &  ni11  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire29192 = ( ni11  &  (~ ni9)  &  (~ ni7)  &  ni8 ) ;
 assign wire29193 = ( pi23  &  (~ ni10)  &  wire29192 ) | ( pi24  &  (~ ni10)  &  wire29192 ) ;
 assign wire29194 = ( (~ ni9)  &  ni11 ) ;
 assign wire29195 = ( (~ ni10)  &  (~ ni7)  &  ni8 ) ;
 assign wire29198 = ( (~ ni14)  &  pi26 ) ;
 assign wire29203 = ( (~ ni9)  &  ni10  &  ni7  &  (~ ni8) ) ;
 assign wire29204 = ( wire1277  &  wire29203 ) ;
 assign wire29206 = ( pi23  &  (~ pi24)  &  (~ ni9)  &  ni10 ) ;
 assign wire29207 = ( ni7  &  (~ ni8)  &  wire29206 ) ;
 assign wire29209 = ( (~ pi23)  &  (~ pi24)  &  (~ ni9)  &  ni10 ) ;
 assign wire29210 = ( ni7  &  (~ ni8)  &  wire29209 ) ;
 assign wire29211 = ( wire6844 ) | ( pi24  &  n_n450 ) | ( pi24  &  wire6852 ) ;
 assign wire29214 = ( (~ ni9)  &  ni10  &  (~ ni8) ) ;
 assign wire29215 = ( pi24  &  ni7  &  wire29214 ) ;
 assign wire29217 = ( (~ pi23)  &  ni7  &  (~ ni8) ) | ( pi24  &  ni7  &  (~ ni8) ) ;
 assign wire29219 = ( (~ ni8)  &  ni7 ) ;
 assign wire29223 = ( (~ pi26)  &  ni11  &  (~ ni9)  &  ni10 ) ;
 assign wire29225 = ( pi23  &  (~ pi24)  &  ni7  &  (~ ni8) ) ;
 assign wire29226 = ( (~ ni11)  &  ni14 ) ;
 assign wire29228 = ( wire948 ) | ( wire980 ) | ( nv10153  &  wire29226 ) ;
 assign wire29231 = ( (~ ni9)  &  (~ ni10)  &  ni7  &  (~ ni8) ) ;
 assign wire29233 = ( (~ ni9)  &  (~ ni10)  &  (~ ni7)  &  ni8 ) ;
 assign wire29234 = ( (~ pi24)  &  (~ ni7)  &  ni8  &  wire264 ) ;
 assign wire29236 = ( pi24  &  (~ ni7)  &  ni8 ) ;
 assign wire29237 = ( ni8  &  ni7 ) ;
 assign wire29240 = ( wire6815 ) | ( wire6816 ) | ( wire6818 ) ;
 assign wire29241 = ( wire6824 ) | ( wire6829 ) | ( wire499  &  wire29193 ) ;
 assign wire29242 = ( wire499  &  wire29234 ) | ( wire264  &  wire499  &  wire29217 ) ;
 assign wire29244 = ( wire6835  &  wire29225 ) | ( wire6836  &  wire29225 ) | ( wire6835  &  wire29236 ) | ( wire6836  &  wire29236 ) ;
 assign wire29247 = ( wire6834 ) | ( wire6833 ) ;
 assign wire29248 = ( wire6820 ) | ( wire29240 ) | ( wire29244 ) ;
 assign wire29249 = ( wire6826 ) | ( wire6831 ) | ( wire29241 ) | ( wire29242 ) ;
 assign wire29252 = ( wire29249 ) | ( wire6832 ) ;
 assign wire29253 = ( wire6819 ) | ( wire6821 ) | ( wire29247 ) | ( wire29248 ) ;
 assign wire29256 = ( (~ ni6)  &  ni5 ) ;
 assign wire29259 = ( wire399  &  ni6 ) ;
 assign wire29261 = ( ni4  &  (~ ni3) ) | ( (~ ni3)  &  (~ ni5) ) ;
 assign wire29264 = ( ni4  &  (~ ni3)  &  ni5 ) ;
 assign wire29268 = ( (~ ni9)  &  ni10  &  ni7  &  (~ ni8) ) ;
 assign wire29269 = ( wire868  &  wire29268 ) ;
 assign wire29270 = ( (~ ni13)  &  (~ ni14)  &  (~ ni11) ) ;
 assign wire29271 = ( (~ ni13)  &  ni14  &  (~ ni11) ) ;
 assign wire29273 = ( pi23  &  (~ pi24)  &  (~ ni9)  &  ni10 ) ;
 assign wire29274 = ( ni7  &  (~ ni8)  &  wire29273 ) ;
 assign wire29276 = ( (~ pi23)  &  (~ ni9)  &  ni10 ) | ( pi24  &  (~ ni9)  &  ni10 ) ;
 assign wire29277 = ( ni7  &  (~ ni8)  &  wire29276 ) ;
 assign wire29279 = ( pi23  &  (~ pi24)  &  ni7  &  (~ ni8) ) ;
 assign wire29280 = ( (~ wire175)  &  wire264  &  wire29279 ) ;
 assign wire29282 = ( (~ pi23)  &  ni7  &  (~ ni8) ) | ( pi24  &  ni7  &  (~ ni8) ) ;
 assign wire29283 = ( (~ wire175)  &  wire264  &  wire29282 ) ;
 assign wire29286 = ( ni7  &  (~ ni8)  &  wire175  &  wire264 ) ;
 assign wire29288 = ( (~ ni9)  &  ni10  &  ni7  &  (~ ni8) ) ;
 assign wire29289 = ( (~ ni13)  &  ni14  &  ni11  &  (~ ni12) ) ;
 assign wire29291 = ( wire6909 ) | ( (~ wire186)  &  nv10237 ) | ( nv10237  &  wire980 ) ;
 assign wire29292 = ( wire6908 ) | ( wire6906 ) ;
 assign wire29294 = ( (~ ni9)  &  (~ ni10)  &  ni7  &  (~ ni8) ) ;
 assign wire29296 = ( pi27  &  (~ ni13)  &  ni14  &  (~ ni11) ) ;
 assign wire29297 = ( ni9  &  ni10  &  (~ ni8) ) ;
 assign wire29298 = ( ni11  &  (~ ni14) ) ;
 assign wire29299 = ( ni12  &  ni14 ) ;
 assign wire29300 = ( ni9  &  ni7 ) | ( ni7  &  ni8 ) ;
 assign wire29303 = ( pi24  &  (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29306 = ( pi24  &  (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29308 = ( (~ pi23)  &  (~ pi24)  &  ni8 ) ;
 assign wire29310 = ( (~ wire175)  &  wire330  &  wire29308 ) ;
 assign wire29311 = ( pi23  &  ni8 ) | ( pi24  &  ni8 ) ;
 assign wire29313 = ( (~ wire175)  &  wire330  &  wire29311 ) ;
 assign wire29315 = ( (~ ni9)  &  (~ ni10)  &  ni8  &  wire868 ) ;
 assign wire29316 = ( (~ pi23)  &  (~ pi24)  &  ni8 ) ;
 assign wire29317 = ( (~ ni9)  &  (~ ni10)  &  wire29316 ) ;
 assign wire29319 = ( pi24  &  (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29320 = ( (~ ni14)  &  ni8 ) | ( ni12  &  ni8 ) ;
 assign wire29323 = ( (~ pi24)  &  (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29324 = ( pi23  &  ni8 ) | ( pi24  &  ni8 ) ;
 assign wire29325 = ( (~ ni9)  &  (~ ni10)  &  wire29324 ) ;
 assign wire29326 = ( (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29328 = ( (~ ni11)  &  ni12  &  ni8 ) ;
 assign wire29331 = ( pi24  &  ni8  &  (~ wire175)  &  wire264 ) ;
 assign wire29333 = ( (~ pi24)  &  ni8  &  (~ wire175)  &  wire264 ) ;
 assign wire29334 = ( ni13  &  ni8 ) | ( (~ ni14)  &  ni8 ) | ( ni12  &  ni8 ) ;
 assign wire29335 = ( ni11  &  (~ ni9)  &  (~ ni10)  &  wire29334 ) ;
 assign wire29336 = ( (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29337 = ( (~ ni9)  &  (~ ni10)  &  ni8 ) ;
 assign wire29338 = ( ni11  &  (~ ni9)  &  ni10  &  ni8 ) ;
 assign wire29340 = ( wire764  &  wire29319 ) | ( nv10167  &  wire764  &  wire29336 ) ;
 assign wire29343 = ( nv10162  &  wire29310 ) | ( nv10187  &  wire29315 ) ;
 assign wire29344 = ( wire6880 ) | ( nv10153  &  wire29331 ) | ( (~ wire155)  &  (~ nv10153)  &  wire29331 ) ;
 assign wire29345 = ( wire6873 ) | ( wire6889 ) | ( nv10187  &  wire29335 ) ;
 assign wire29346 = ( wire6883 ) | ( nv10178  &  wire29313 ) ;
 assign wire29347 = ( wire6884 ) | ( nv10178  &  wire29333 ) ;
 assign wire29348 = ( wire6874 ) | ( wire6890 ) | ( wire29340 ) ;
 assign wire29352 = ( wire6878 ) | ( wire29343 ) | ( wire29344 ) ;
 assign wire29353 = ( wire6898  &  wire29323 ) | ( wire6899  &  wire29323 ) | ( wire6898  &  wire29325 ) | ( wire6899  &  wire29325 ) ;
 assign wire29354 = ( wire29345 ) | ( wire29346 ) | ( wire29347 ) | ( wire29348 ) ;
 assign wire29358 = ( (~ wire399)  &  nv10153  &  wire29298 ) | ( (~ wire399)  &  nv10153  &  wire29299 ) ;
 assign wire29360 = ( nv10222  &  wire29269 ) | ( nv10162  &  wire29280 ) ;
 assign wire29361 = ( wire6869 ) | ( nv10222  &  wire29286 ) ;
 assign wire29362 = ( wire6862 ) | ( wire6864 ) | ( wire6870 ) | ( wire29358 ) ;
 assign wire29366 = ( wire6857 ) | ( wire29361 ) | ( wire29362 ) ;
 assign wire29367 = ( wire6858 ) | ( wire6860 ) | ( wire6871 ) | ( wire29360 ) ;
 assign wire29368 = ( wire29291  &  wire29294 ) | ( wire29292  &  wire29294 ) | ( wire29291  &  wire29297 ) | ( wire29292  &  wire29297 ) ;
 assign wire29371 = ( wire6868 ) | ( wire29366 ) | ( wire29367 ) | ( wire29368 ) ;
 assign wire29372 = ( (~ ni3)  &  wire29371 ) | ( (~ ni3)  &  (~ ni7)  &  n_n983 ) ;
 assign wire29376 = ( ni5  &  (~ ni3) ) ;
 assign wire29377 = ( wire29371  &  wire29376 ) | ( (~ ni7)  &  n_n983  &  wire29376 ) ;
 assign wire29379 = ( (~ ni3)  &  ni5  &  (~ ni6) ) ;
 assign wire29382 = ( (~ ni3)  &  (~ ni4) ) ;
 assign wire29385 = ( (~ ni4)  &  ni3  &  (~ ni5) ) | ( (~ ni4)  &  (~ ni3)  &  (~ ni6) ) ;
 assign wire29386 = ( (~ ni4)  &  (~ ni3)  &  (~ ni5) ) | ( (~ ni4)  &  ni3  &  wire478 ) | ( ni4  &  ni3  &  ni5  &  (~ wire478) ) ;
 assign wire29388 = ( wire6795 ) | ( wire29385 ) | ( wire29386 ) ;
 assign wire29393 = ( wire6796 ) | ( wire6802 ) | ( wire6805 ) | ( wire29388 ) ;
 assign wire29394 = ( wire6797 ) | ( wire6799 ) | ( wire6800 ) | ( wire6801 ) ;
 assign wire29395 = ( pi26  &  ni33  &  (~ ni32) ) ;
 assign wire29397 = ( (~ ni9)  &  wire29395 ) | ( (~ ni10)  &  wire29395 ) | ( (~ wire1289)  &  wire29395 ) ;
 assign wire29398 = ( (~ ni2)  &  (~ ni3)  &  (~ nv7447)  &  (~ wire281) ) ;
 assign wire29400 = ( pi26  &  ni33  &  (~ ni32) ) ;
 assign wire29403 = ( (~ wire290)  &  wire462  &  (~ nv10169)  &  wire29400 ) ;
 assign wire29404 = ( pi23  &  (~ ni33)  &  (~ ni32) ) ;
 assign wire29407 = ( (~ wire290)  &  wire462  &  (~ nv10169)  &  wire29404 ) ;
 assign wire29408 = ( (~ pi26)  &  ni35 ) | ( (~ pi23)  &  ni35 ) ;
 assign wire29410 = ( ni31  &  (~ wire290)  &  wire29408 ) | ( (~ ni30)  &  (~ wire290)  &  wire29408 ) ;
 assign wire29411 = ( (~ pi26)  &  ni35  &  ni32 ) | ( (~ pi23)  &  ni35  &  ni32 ) ;
 assign wire29413 = ( (~ ni31)  &  ni30  &  (~ wire290)  &  wire29411 ) ;
 assign wire29414 = ( ni35  &  ni32  &  (~ wire290) ) ;
 assign wire29415 = ( n_n13895  &  (~ nv10130)  &  (~ wire281) ) | ( n_n13895  &  (~ wire281)  &  wire202 ) ;
 assign wire29417 = ( ni35  &  (~ ni33) ) | ( ni35  &  (~ ni30) ) ;
 assign wire29418 = ( (~ ni9)  &  wire29417 ) | ( (~ ni10)  &  wire29417 ) | ( (~ wire1289)  &  wire29417 ) ;
 assign wire29419 = ( ni31  &  ni35 ) ;
 assign wire29420 = ( (~ ni9)  &  wire29419 ) | ( (~ ni10)  &  wire29419 ) | ( (~ wire1289)  &  wire29419 ) ;
 assign wire29423 = ( ni13  &  (~ ni14)  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire29424 = ( nv10130  &  wire1289  &  (~ wire281)  &  wire29423 ) ;
 assign wire29425 = ( nv10130  &  wire1289  &  wire630  &  (~ wire281) ) ;
 assign wire29427 = ( ni35  &  pi26 ) ;
 assign wire29429 = ( wire6788 ) | ( wire1105  &  wire29403 ) ;
 assign wire29430 = ( wire1105  &  wire29407 ) | ( wire1105  &  wire29410 ) ;
 assign wire29431 = ( wire6786 ) | ( wire6787 ) | ( wire1105  &  wire29413 ) ;
 assign wire29433 = ( (~ wire6789)  &  (~ wire6790)  &  wire29418 ) | ( (~ wire6789)  &  (~ wire6790)  &  wire29420 ) ;
 assign wire29437 = ( wire6775 ) | ( wire6780 ) | ( wire29433 ) ;
 assign wire29438 = ( wire6783 ) | ( wire6784 ) | ( wire6785 ) | ( wire29429 ) ;
 assign wire29440 = ( (~ ni2)  &  (~ ni12)  &  (~ ni3) ) ;
 assign wire29441 = ( ni13  &  ni14  &  wire29440 ) ;
 assign wire29444 = ( (~ ni13)  &  ni12 ) | ( (~ ni14)  &  ni12 ) ;
 assign wire29447 = ( ni12  &  (~ n_n13895) ) | ( ni11  &  ni12  &  (~ nv10086) ) | ( ni11  &  (~ ni12)  &  n_n13895  &  nv10086 ) ;
 assign wire29449 = ( wire6745 ) | ( wire1075 ) ;
 assign wire29451 = ( pi15  &  wire1066  &  wire376 ) ;
 assign wire29452 = ( wire317 ) | ( nv910  &  wire6757 ) | ( nv910  &  wire6758 ) ;
 assign wire29454 = ( pi21  &  pi22  &  pi15  &  wire1066 ) ;
 assign wire29455 = ( wire6705 ) | ( wire1075 ) ;
 assign wire29458 = ( wire317 ) | ( nv919  &  wire6757 ) | ( nv919  &  wire6758 ) ;
 assign wire29460 = ( pi21  &  pi22  &  pi15  &  wire1058 ) ;
 assign wire29461 = ( pi15  &  ni33  &  (~ ni32) ) ;
 assign wire29462 = ( pi17  &  (~ pi16)  &  wire152  &  wire29461 ) ;
 assign wire29465 = ( ni34  &  pi15 ) ;
 assign wire29466 = ( wire6666 ) | ( wire1097 ) ;
 assign wire29467 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  wire376 ) ;
 assign wire29468 = ( wire317 ) | ( nv890  &  wire6757 ) | ( nv890  &  wire6758 ) ;
 assign wire29469 = ( pi21  &  pi22  &  wire616 ) ;
 assign wire29470 = ( wire6682 ) | ( wire1097 ) ;
 assign wire29471 = ( (~ pi17)  &  pi19  &  pi20  &  wire376 ) ;
 assign wire29472 = ( wire317 ) | ( nv899  &  wire6757 ) | ( nv899  &  wire6758 ) ;
 assign wire29473 = ( pi21  &  pi22  &  wire381 ) ;
 assign wire29474 = ( wire6721 ) | ( wire441  &  wire269 ) ;
 assign wire29475 = ( (~ ni38)  &  ni37  &  ni36 ) | ( ni37  &  ni36  &  wire441 ) | ( (~ ni37)  &  ni36  &  wire441 ) ;
 assign wire29476 = ( wire1060 ) | ( wire6722 ) | ( wire29474 ) ;
 assign wire29479 = ( wire317 ) | ( ni34  &  wire332 ) | ( wire332  &  (~ wire943) ) ;
 assign wire29481 = ( ni36  &  nv628 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29485 = ( wire6332 ) | ( wire6333 ) | ( wire228  &  wire368 ) ;
 assign wire29486 = ( wire29485 ) | ( pi20  &  wire191  &  wire368 ) | ( (~ pi20)  &  wire191  &  wire368 ) ;
 assign wire29488 = ( wire6272 ) | ( wire29486 ) | ( nv890  &  wire29467 ) ;
 assign wire29490 = ( wire6276 ) | ( wire6287  &  wire29469 ) | ( wire29468  &  wire29469 ) ;
 assign wire29491 = ( wire6270 ) | ( wire29488 ) | ( nv899  &  wire29471 ) ;
 assign wire29495 = ( pi17  &  (~ pi16)  &  (~ ni29)  &  wire152 ) ;
 assign wire29496 = ( wire158  &  wire152  &  wire6757 ) | ( wire158  &  wire152  &  wire6758 ) ;
 assign wire29497 = ( wire158  &  n_n11316 ) | ( wire158  &  wire152  &  wire317 ) ;
 assign wire29498 = ( wire29497 ) | ( nv928  &  wire29496 ) ;
 assign wire29499 = ( pi17  &  pi16  &  (~ ni29)  &  wire152 ) ;
 assign wire29501 = ( wire152  &  wire154  &  wire6757 ) | ( wire152  &  wire154  &  wire6758 ) ;
 assign wire29502 = ( n_n11316  &  wire154 ) | ( wire152  &  wire317  &  wire154 ) ;
 assign wire29504 = ( wire6580 ) | ( wire1097 ) ;
 assign wire29505 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29506 = ( wire29505  &  wire376 ) ;
 assign wire29507 = ( (~ ni29)  &  ni34 ) ;
 assign wire29508 = ( (~ ni29)  &  (~ ni34) ) ;
 assign wire29510 = ( pi21  &  pi22  &  pi16 ) ;
 assign wire29512 = ( wire6616 ) | ( wire1097 ) ;
 assign wire29513 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29514 = ( wire29513  &  wire376 ) ;
 assign wire29515 = ( wire317 ) | ( nv968  &  wire6757 ) | ( nv968  &  wire6758 ) ;
 assign wire29517 = ( pi21  &  pi22  &  pi16  &  wire381 ) ;
 assign wire29518 = ( ni36  &  nv772 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29520 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29521 = ( wire29520  &  wire376 ) ;
 assign wire29525 = ( pi21  &  pi22  &  pi16  &  wire228 ) ;
 assign wire29526 = ( wire6560 ) | ( wire1075 ) ;
 assign wire29527 = ( wire376  &  wire1073 ) ;
 assign wire29528 = ( wire317 ) | ( nv979  &  wire6757 ) | ( nv979  &  wire6758 ) ;
 assign wire29529 = ( pi21  &  pi22  &  wire1073 ) ;
 assign wire29530 = ( wire6540 ) | ( wire1075 ) ;
 assign wire29531 = ( wire376  &  wire1045 ) ;
 assign wire29532 = ( wire317 ) | ( nv988  &  wire6757 ) | ( nv988  &  wire6758 ) ;
 assign wire29533 = ( pi21  &  pi22  &  wire1045 ) ;
 assign wire29534 = ( ni36  &  nv758 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29536 = ( (~ pi20)  &  pi16  &  n_n13390  &  wire153 ) ;
 assign wire29537 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29538 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29539 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29540 = ( ni33  &  (~ ni32)  &  wire152  &  wire154 ) ;
 assign wire29542 = ( (~ pi20)  &  pi16  &  wire153 ) ;
 assign wire29543 = ( pi21  &  ni34  &  wire1045 ) | ( pi21  &  ni34  &  wire1073 ) ;
 assign wire29544 = ( wire6240 ) | ( pi21  &  ni34  &  wire29537 ) ;
 assign wire29545 = ( pi21  &  ni34  &  wire29538 ) | ( pi21  &  ni34  &  wire29539 ) ;
 assign wire29548 = ( wire6239 ) | ( wire29543 ) | ( wire29544 ) | ( wire29545 ) ;
 assign wire29550 = ( wire947 ) | ( wire6235 ) | ( wire29548 ) ;
 assign wire29553 = ( nv968  &  wire29514 ) | ( nv979  &  wire29527 ) ;
 assign wire29554 = ( wire6225 ) | ( wire29550 ) | ( nv988  &  wire29531 ) ;
 assign wire29555 = ( wire6231 ) | ( wire29553 ) | ( nv959  &  wire29506 ) ;
 assign wire29556 = ( wire29554 ) | ( wire616  &  n_n11474  &  wire29510 ) ;
 assign wire29561 = ( wire6224 ) | ( wire6228 ) | ( wire6230 ) | ( wire29555 ) ;
 assign wire29562 = ( ni36  &  wire388 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29563 = ( pi17  &  pi16  &  (~ ni29)  &  wire152 ) ;
 assign wire29564 = ( wire29562  &  wire29563 ) | ( (~ ni36)  &  nv858  &  wire29563 ) ;
 assign wire29565 = ( wire152  &  wire154  &  wire6757 ) | ( wire152  &  wire154  &  wire6758 ) ;
 assign wire29566 = ( n_n11316  &  wire154 ) | ( wire152  &  wire317  &  wire154 ) ;
 assign wire29567 = ( wire29566 ) | ( ni34  &  wire29564 ) | ( wire6524  &  wire29564 ) ;
 assign wire29568 = ( wire6576 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29569 = ( wire436 ) | ( wire6576 ) | ( wire6578 ) ;
 assign wire29570 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29571 = ( wire29570  &  wire376 ) ;
 assign wire29572 = ( wire317 ) | ( nv779  &  wire6757 ) | ( nv779  &  wire6758 ) ;
 assign wire29574 = ( pi21  &  pi22  &  pi16  &  wire616 ) ;
 assign wire29575 = ( wire6612 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29576 = ( wire436 ) | ( wire6612 ) | ( wire6614 ) ;
 assign wire29577 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29578 = ( wire29577  &  wire376 ) ;
 assign wire29579 = ( wire317 ) | ( nv797  &  wire6757 ) | ( nv797  &  wire6758 ) ;
 assign wire29581 = ( pi21  &  pi22  &  pi16  &  wire381 ) ;
 assign wire29582 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29583 = ( wire29582  &  wire376 ) ;
 assign wire29584 = ( wire317 ) | ( nv764  &  wire6757 ) | ( nv764  &  wire6758 ) ;
 assign wire29586 = ( pi21  &  pi22  &  pi16  &  wire228 ) ;
 assign wire29587 = ( wire6556 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29588 = ( wire436 ) | ( wire6556 ) | ( wire6558 ) ;
 assign wire29589 = ( wire376  &  wire1073 ) ;
 assign wire29590 = ( wire317 ) | ( nv817  &  wire6757 ) | ( nv817  &  wire6758 ) ;
 assign wire29591 = ( pi21  &  pi22  &  wire1073 ) ;
 assign wire29592 = ( wire6536 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29593 = ( wire436 ) | ( wire6536 ) | ( wire6538 ) ;
 assign wire29594 = ( wire376  &  wire1045 ) ;
 assign wire29595 = ( wire317 ) | ( nv835  &  wire6757 ) | ( nv835  &  wire6758 ) ;
 assign wire29596 = ( pi21  &  pi22  &  wire1045 ) ;
 assign wire29597 = ( (~ pi20)  &  pi16  &  n_n13390  &  wire153 ) ;
 assign wire29598 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29599 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29600 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29601 = ( ni33  &  (~ ni32)  &  wire152  &  wire154 ) ;
 assign wire29602 = ( wire317 ) | ( nv750  &  wire6757 ) | ( nv750  &  wire6758 ) ;
 assign wire29603 = ( (~ pi20)  &  pi16  &  wire153 ) ;
 assign wire29604 = ( pi21  &  ni34  &  wire1045 ) | ( pi21  &  ni34  &  wire1073 ) ;
 assign wire29605 = ( wire6309 ) | ( pi21  &  ni34  &  wire29598 ) ;
 assign wire29606 = ( pi21  &  ni34  &  wire29599 ) | ( pi21  &  ni34  &  wire29600 ) ;
 assign wire29609 = ( wire6308 ) | ( wire29604 ) | ( wire29605 ) | ( wire29606 ) ;
 assign wire29610 = ( wire29609 ) | ( ni34  &  wire29601 ) | ( wire6524  &  wire29601 ) ;
 assign wire29611 = ( wire6521 ) | ( wire29567 ) | ( wire29610 ) ;
 assign wire29612 = ( nv764  &  wire29583 ) | ( nv750  &  wire29597 ) ;
 assign wire29615 = ( wire6295 ) | ( wire6305 ) | ( wire29611 ) | ( wire29612 ) ;
 assign wire29616 = ( nv779  &  wire29571 ) | ( nv797  &  wire29578 ) ;
 assign wire29617 = ( nv817  &  wire29589 ) | ( nv835  &  wire29594 ) ;
 assign wire29619 = ( wire29615 ) | ( wire29616 ) | ( wire29617 ) ;
 assign wire29621 = ( wire6297 ) | ( wire6531  &  wire29596 ) | ( wire29595  &  wire29596 ) ;
 assign wire29622 = ( wire6291 ) | ( wire6293 ) | ( wire29619 ) ;
 assign wire29623 = ( wire6692 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29624 = ( pi17  &  (~ pi16)  &  (~ ni29)  &  wire152 ) ;
 assign wire29625 = ( wire158  &  wire152  &  wire6757 ) | ( wire158  &  wire152  &  wire6758 ) ;
 assign wire29626 = ( wire158  &  n_n11316 ) | ( wire158  &  wire152  &  wire317 ) ;
 assign wire29627 = ( wire29626 ) | ( nv735  &  wire29625 ) ;
 assign wire29628 = ( wire6662 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29629 = ( wire436 ) | ( wire6662 ) | ( wire6664 ) ;
 assign wire29630 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29631 = ( wire29630  &  wire376 ) ;
 assign wire29632 = ( wire317 ) | ( nv658  &  wire6757 ) | ( nv658  &  wire6758 ) ;
 assign wire29634 = ( pi21  &  pi22  &  (~ pi16)  &  wire616 ) ;
 assign wire29635 = ( wire6679 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29636 = ( wire436 ) | ( wire6678 ) | ( wire6679 ) ;
 assign wire29637 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29639 = ( wire317 ) | ( nv679  &  wire6757 ) | ( nv679  &  wire6758 ) ;
 assign wire29641 = ( pi21  &  pi22  &  (~ pi16)  &  wire381 ) ;
 assign wire29642 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29644 = ( wire317 ) | ( ni34  &  wire332 ) | ( wire332  &  (~ wire785) ) ;
 assign wire29645 = ( pi21  &  pi22  &  (~ pi16) ) ;
 assign wire29647 = ( wire6741 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29648 = ( wire436 ) | ( wire6741 ) | ( wire6743 ) ;
 assign wire29649 = ( wire376  &  wire1066 ) ;
 assign wire29650 = ( wire317 ) | ( nv699  &  wire6757 ) | ( nv699  &  wire6758 ) ;
 assign wire29651 = ( pi21  &  pi22  &  wire1066 ) ;
 assign wire29652 = ( wire6702 ) | ( (~ ni38)  &  ni37  &  ni36 ) ;
 assign wire29653 = ( wire436 ) | ( wire6701 ) | ( wire6702 ) ;
 assign wire29655 = ( wire317 ) | ( nv717  &  wire6757 ) | ( nv717  &  wire6758 ) ;
 assign wire29656 = ( pi21  &  pi22  &  wire1058 ) ;
 assign wire29657 = ( (~ pi20)  &  (~ pi16)  &  n_n13390  &  wire153 ) ;
 assign wire29658 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29659 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29660 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29662 = ( wire317 ) | ( nv620  &  wire6757 ) | ( nv620  &  wire6758 ) ;
 assign wire29663 = ( (~ pi20)  &  (~ pi16)  &  wire153 ) ;
 assign wire29664 = ( pi21  &  ni34  &  wire1058 ) | ( pi21  &  ni34  &  wire1066 ) ;
 assign wire29665 = ( wire6330 ) | ( pi21  &  ni34  &  wire29658 ) ;
 assign wire29666 = ( pi21  &  ni34  &  wire29659 ) | ( pi21  &  ni34  &  wire29660 ) ;
 assign wire29669 = ( wire6329 ) | ( wire29664 ) | ( wire29665 ) | ( wire29666 ) ;
 assign wire29670 = ( wire29669 ) | ( nv620  &  wire29657 ) ;
 assign wire29672 = ( wire6325 ) | ( wire6647 ) | ( wire29627 ) | ( wire29670 ) ;
 assign wire29674 = ( wire6315 ) | ( wire6326 ) | ( wire29672 ) ;
 assign wire29675 = ( nv658  &  wire29631 ) | ( nv699  &  wire29649 ) ;
 assign wire29677 = ( wire6316 ) | ( nv679  &  wire376  &  wire29637 ) ;
 assign wire29680 = ( wire6319 ) | ( wire29674 ) | ( wire29675 ) | ( wire29677 ) ;
 assign wire29681 = ( wire6312 ) | ( wire6318 ) | ( wire29680 ) ;
 assign wire29682 = ( wire6314 ) | ( wire6696  &  wire29656 ) | ( wire29655  &  wire29656 ) ;
 assign wire29684 = ( wire6209 ) | ( wire6210 ) | ( wire295  &  wire29465 ) ;
 assign wire29685 = ( wire29684 ) | ( nv928  &  wire29462 ) ;
 assign wire29686 = ( wire29685 ) | ( pi15  &  wire6217 ) | ( pi15  &  wire29498 ) ;
 assign wire29687 = ( wire29686 ) | ( nv910  &  wire29451 ) ;
 assign wire29690 = ( wire6205 ) | ( wire6206 ) | ( wire6207 ) | ( wire29687 ) ;
 assign wire29691 = ( wire29690 ) | ( (~ pi16)  &  pi15  &  n_n11833 ) ;
 assign wire29692 = ( pi15  &  n_n11836 ) | ( (~ pi15)  &  wire29681 ) | ( (~ pi15)  &  wire29682 ) ;
 assign wire29693 = ( wire29691 ) | ( (~ pi15)  &  wire29621 ) | ( (~ pi15)  &  wire29622 ) ;
 assign wire29695 = ( pi21  &  pi16 ) | ( pi16  &  (~ ni34) ) ;
 assign wire29697 = ( pi21  &  pi16 ) | ( pi16  &  (~ ni34) ) ;
 assign wire29699 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29700 = ( pi21  &  pi22  &  wire312  &  wire29699 ) ;
 assign wire29702 = ( pi21  &  pi22  &  pi16  &  wire381 ) ;
 assign wire29703 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29704 = ( pi21  &  pi22  &  wire312  &  wire29703 ) ;
 assign wire29706 = ( pi21  &  pi22  &  pi16  &  wire228 ) ;
 assign wire29707 = ( (~ pi20)  &  pi16  &  wire312  &  wire153 ) ;
 assign wire29709 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire29710 = ( pi21  &  pi22  &  wire312  &  wire1045 ) ;
 assign wire29711 = ( pi21  &  pi22  &  wire1045 ) ;
 assign wire29713 = ( pi21  &  wire224 ) | ( wire380  &  nv779 ) ;
 assign wire29715 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29716 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29717 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29718 = ( pi17  &  pi16  &  wire152  &  wire312 ) ;
 assign wire29719 = ( wire257  &  wire29562 ) | ( (~ ni36)  &  wire257  &  nv858 ) ;
 assign wire29720 = ( (~ pi20)  &  pi16  &  wire153 ) ;
 assign wire29721 = ( pi21  &  wire224 ) | ( wire380  &  nv817 ) ;
 assign wire29723 = ( wire224  &  wire257 ) | ( pi21  &  wire224  &  wire29716 ) ;
 assign wire29724 = ( pi21  &  wire224  &  wire1045 ) | ( pi21  &  wire224  &  wire29717 ) ;
 assign wire29726 = ( wire6517 ) | ( wire29723 ) | ( wire29724 ) ;
 assign wire29727 = ( wire29726 ) | ( ni34  &  wire29718 ) | ( wire6524  &  wire29718 ) ;
 assign wire29729 = ( wire6513 ) | ( wire6521 ) | ( wire29567 ) | ( wire29727 ) ;
 assign wire29730 = ( nv764  &  wire29704 ) | ( nv750  &  wire29707 ) ;
 assign wire29733 = ( wire6498 ) | ( wire6506 ) | ( wire29729 ) | ( wire29730 ) ;
 assign wire29735 = ( wire6503 ) | ( wire6514 ) | ( wire29733 ) ;
 assign wire29736 = ( nv797  &  wire29700 ) | ( nv835  &  wire29710 ) ;
 assign wire29739 = ( wire6499 ) | ( wire6505 ) | ( wire29735 ) | ( wire29736 ) ;
 assign wire29741 = ( wire6501 ) | ( wire6508 ) | ( wire29739 ) ;
 assign wire29743 = ( (~ pi15)  &  (~ wire265)  &  (~ wire289)  &  wire510 ) ;
 assign wire29745 = ( pi21  &  (~ pi16)  &  wire381 ) | ( (~ pi16)  &  (~ ni34)  &  wire381 ) ;
 assign wire29746 = ( pi21  &  (~ pi16) ) | ( (~ pi16)  &  (~ ni34) ) ;
 assign wire29748 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29749 = ( pi21  &  pi22  &  wire312  &  wire29748 ) ;
 assign wire29751 = ( pi21  &  pi22  &  (~ pi16)  &  wire381 ) ;
 assign wire29752 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29753 = ( pi21  &  pi22  &  wire312  &  wire29752 ) ;
 assign wire29754 = ( pi21  &  pi22  &  (~ pi16) ) ;
 assign wire29756 = ( (~ pi20)  &  (~ pi16)  &  wire312  &  wire153 ) ;
 assign wire29757 = ( pi21  &  wire1058 ) | ( (~ ni34)  &  wire1058 ) ;
 assign wire29759 = ( pi21  &  pi22  &  wire1058 ) ;
 assign wire29760 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29761 = ( pi21  &  wire224 ) | ( wire380  &  nv658 ) ;
 assign wire29762 = ( wire29761 ) | ( pi21  &  wire1310 ) | ( (~ ni34)  &  wire1310 ) ;
 assign wire29763 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29764 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29765 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29766 = ( pi17  &  (~ pi16)  &  wire152  &  wire312 ) ;
 assign wire29767 = ( (~ pi20)  &  (~ pi16)  &  wire153 ) ;
 assign wire29768 = ( nv699  &  wire380 ) | ( pi21  &  wire224 ) ;
 assign wire29769 = ( wire29768 ) | ( pi21  &  wire1332 ) | ( (~ ni34)  &  wire1332 ) ;
 assign wire29770 = ( wire224  &  wire295 ) | ( pi21  &  wire224  &  wire29764 ) ;
 assign wire29771 = ( pi21  &  wire224  &  wire1058 ) | ( pi21  &  wire224  &  wire29765 ) ;
 assign wire29773 = ( wire6644 ) | ( wire29770 ) | ( wire29771 ) ;
 assign wire29774 = ( wire29773 ) | ( nv620  &  wire29756 ) ;
 assign wire29775 = ( wire1012  &  wire29760 ) | ( nv735  &  wire29766 ) ;
 assign wire29776 = ( wire29774 ) | ( wire1131  &  wire295 ) ;
 assign wire29779 = ( wire6629 ) | ( wire6647 ) | ( wire29627 ) | ( wire29775 ) ;
 assign wire29781 = ( wire6626 ) | ( wire6640 ) | ( wire29776 ) | ( wire29779 ) ;
 assign wire29782 = ( wire6630 ) | ( nv679  &  wire29749 ) ;
 assign wire29784 = ( wire1057  &  wire29745 ) | ( wire1092  &  wire29757 ) ;
 assign wire29786 = ( wire6633 ) | ( wire29781 ) | ( wire29782 ) | ( wire29784 ) ;
 assign wire29789 = ( wire6628 ) | ( wire6634 ) | ( wire29786 ) ;
 assign wire29790 = ( (~ pi15)  &  (~ wire265)  &  (~ wire289)  &  wire510 ) ;
 assign wire29792 = ( pi21  &  pi16  &  wire381 ) | ( pi16  &  (~ ni34)  &  wire381 ) ;
 assign wire29793 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29794 = ( pi21  &  pi22  &  wire312  &  wire29793 ) ;
 assign wire29796 = ( pi21  &  pi22  &  pi16  &  wire381 ) ;
 assign wire29797 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29798 = ( pi21  &  pi22  &  wire312  &  wire29797 ) ;
 assign wire29799 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29800 = ( pi21  &  ni34  &  wire29799 ) ;
 assign wire29802 = ( pi21  &  pi22  &  pi16  &  wire228 ) ;
 assign wire29803 = ( (~ pi20)  &  pi16  &  wire312  &  wire153 ) ;
 assign wire29805 = ( pi21  &  pi22  &  wire312  &  wire1045 ) ;
 assign wire29806 = ( pi21  &  pi22  &  wire1045 ) ;
 assign wire29807 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire29808 = ( wire379 ) | ( wire368  &  wire6581 ) | ( wire368  &  wire29504 ) ;
 assign wire29809 = ( wire29808 ) | ( (~ wire150)  &  nv959  &  wire312 ) ;
 assign wire29810 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire29811 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire29812 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire29813 = ( pi17  &  pi16  &  wire152  &  wire312 ) ;
 assign wire29815 = ( (~ pi20)  &  pi16  &  wire153 ) ;
 assign wire29816 = ( pi21  &  wire224 ) | ( wire380  &  nv979 ) ;
 assign wire29818 = ( wire224  &  wire257 ) | ( pi21  &  wire224  &  wire29811 ) ;
 assign wire29819 = ( pi21  &  wire224  &  wire1045 ) | ( pi21  &  wire224  &  wire29812 ) ;
 assign wire29821 = ( wire5992 ) | ( wire29818 ) | ( wire29819 ) ;
 assign wire29823 = ( wire5987 ) | ( wire5988 ) | ( wire29821 ) ;
 assign wire29825 = ( wire947 ) | ( wire29823 ) | ( nv952  &  wire29800 ) ;
 assign wire29827 = ( wire5979 ) | ( nv968  &  wire29794 ) ;
 assign wire29829 = ( wire5976 ) | ( wire29825 ) | ( wire1046  &  wire29792 ) ;
 assign wire29830 = ( wire29827 ) | ( (~ n_n11316)  &  wire1038  &  wire1045 ) ;
 assign wire29831 = ( wire5978 ) | ( wire5983 ) | ( nv988  &  wire29805 ) ;
 assign wire29835 = ( wire5984 ) | ( wire5989 ) | ( wire29829 ) ;
 assign wire29836 = ( wire5975 ) | ( wire5982 ) | ( wire29830 ) | ( wire29831 ) ;
 assign wire29838 = ( pi15  &  (~ wire265)  &  (~ wire289)  &  wire510 ) ;
 assign wire29839 = ( pi21  &  (~ pi16) ) | ( (~ pi16)  &  (~ ni34) ) ;
 assign wire29842 = ( pi21  &  (~ pi16)  &  wire381 ) | ( (~ pi16)  &  (~ ni34)  &  wire381 ) ;
 assign wire29843 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29846 = ( pi21  &  pi22  &  (~ pi16)  &  wire381 ) ;
 assign wire29847 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29848 = ( pi21  &  pi22  &  wire312  &  wire29847 ) ;
 assign wire29849 = ( pi21  &  pi22  &  (~ pi16) ) ;
 assign wire29851 = ( (~ pi20)  &  (~ pi16)  &  wire312  &  wire153 ) ;
 assign wire29852 = ( pi21  &  wire1058 ) | ( (~ ni34)  &  wire1058 ) ;
 assign wire29854 = ( pi21  &  pi22  &  wire1058 ) ;
 assign wire29855 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29856 = ( wire380  &  nv890 ) | ( pi21  &  wire224 ) ;
 assign wire29857 = ( wire29856 ) | ( pi21  &  wire1334 ) | ( (~ ni34)  &  wire1334 ) ;
 assign wire29858 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire29859 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire29860 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire29861 = ( pi17  &  (~ pi16)  &  wire152  &  wire312 ) ;
 assign wire29862 = ( (~ pi20)  &  (~ pi16)  &  wire153 ) ;
 assign wire29863 = ( pi21  &  wire224 ) | ( wire380  &  nv910 ) ;
 assign wire29864 = ( wire29863 ) | ( pi21  &  wire1312 ) | ( (~ ni34)  &  wire1312 ) ;
 assign wire29865 = ( wire224  &  wire295 ) | ( pi21  &  wire224  &  wire29859 ) ;
 assign wire29866 = ( pi21  &  wire224  &  wire1058 ) | ( pi21  &  wire224  &  wire29860 ) ;
 assign wire29868 = ( wire6193 ) | ( wire29865 ) | ( wire29866 ) ;
 assign wire29869 = ( wire29868 ) | ( nv928  &  wire29861 ) ;
 assign wire29871 = ( wire6192 ) | ( wire6217 ) | ( wire29498 ) | ( wire29869 ) ;
 assign wire29873 = ( wire6180 ) | ( wire6184 ) | ( wire29871 ) ;
 assign wire29876 = ( wire1033  &  wire29842 ) | ( wire1039  &  wire29852 ) ;
 assign wire29877 = ( wire6176 ) | ( wire6182 ) | ( wire6189 ) | ( wire29873 ) ;
 assign wire29878 = ( wire29876 ) | ( ni34  &  wire29848 ) | ( (~ wire943)  &  wire29848 ) ;
 assign wire29880 = ( wire6177 ) | ( wire6337  &  wire29854 ) | ( wire29458  &  wire29854 ) ;
 assign wire29884 = ( wire6174 ) | ( wire6179 ) | ( wire29877 ) | ( wire29878 ) ;
 assign wire29885 = ( pi15  &  (~ wire265)  &  (~ wire289)  &  wire510 ) ;
 assign wire29886 = ( (~ wire265)  &  wire175  &  wire510 ) ;
 assign wire29888 = ( pi25  &  pi15  &  (~ ni10) ) ;
 assign wire29890 = ( wire289  &  wire178  &  wire154  &  wire29888 ) ;
 assign wire29892 = ( (~ pi16)  &  pi15  &  (~ ni10) ) ;
 assign wire29894 = ( wire289  &  wire475  &  wire29892 ) ;
 assign wire29896 = ( pi16  &  pi15  &  (~ ni10) ) ;
 assign wire29898 = ( wire289  &  wire475  &  wire29896 ) ;
 assign wire29900 = ( pi25  &  pi15  &  (~ ni10) ) ;
 assign wire29902 = ( wire289  &  wire158  &  wire178  &  wire29900 ) ;
 assign wire29905 = ( (~ pi16)  &  pi15  &  (~ ni10)  &  wire289 ) ;
 assign wire29908 = ( (~ pi16)  &  pi15  &  (~ ni10) ) ;
 assign wire29910 = ( wire289  &  wire437  &  wire29908 ) ;
 assign wire29912 = ( pi16  &  pi15  &  (~ ni10) ) ;
 assign wire29914 = ( wire289  &  wire219  &  wire29912 ) ;
 assign wire29916 = ( pi16  &  pi15  &  (~ ni10) ) ;
 assign wire29918 = ( wire289  &  wire437  &  wire29916 ) ;
 assign wire29920 = ( pi16  &  pi15  &  (~ ni10) ) ;
 assign wire29922 = ( wire289  &  wire247  &  wire29920 ) ;
 assign wire29924 = ( (~ pi16)  &  pi15  &  (~ ni10) ) ;
 assign wire29926 = ( wire289  &  wire219  &  wire29924 ) ;
 assign wire29929 = ( pi15  &  (~ ni10)  &  wire289  &  wire813 ) ;
 assign wire29932 = ( pi15  &  (~ ni10)  &  wire289  &  wire812 ) ;
 assign wire29933 = ( (~ ni10)  &  pi15 ) ;
 assign wire29937 = ( pi17  &  (~ pi16)  &  pi15  &  (~ ni10) ) ;
 assign wire29940 = ( pi17  &  pi16  &  pi15  &  (~ ni10) ) ;
 assign wire29943 = ( pi15  &  (~ ni10)  &  wire289 ) ;
 assign wire29945 = ( (~ pi17)  &  pi25  &  pi16  &  wire179 ) ;
 assign wire29946 = ( (~ pi17)  &  pi25  &  pi16  &  wire182 ) ;
 assign wire29947 = ( pi17  &  pi25  &  pi16  &  wire178 ) ;
 assign wire29948 = ( pi20  &  pi25  &  pi16  &  wire153 ) ;
 assign wire29949 = ( (~ pi20)  &  pi25  &  pi16  &  wire153 ) ;
 assign wire29950 = ( pi17  &  pi16  &  wire343 ) | ( (~ pi17)  &  pi16  &  wire343 ) ;
 assign wire29951 = ( wire29950 ) | ( ni34  &  wire311 ) | ( wire311  &  wire6524 ) ;
 assign wire29952 = ( wire29951 ) | ( nv764  &  wire29948 ) ;
 assign wire29954 = ( wire6087 ) | ( wire29952 ) | ( nv779  &  wire29945 ) ;
 assign wire29955 = ( nv797  &  wire29946 ) | ( nv817  &  wire29947 ) ;
 assign wire29958 = ( (~ pi15)  &  (~ ni10)  &  wire289 ) ;
 assign wire29959 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire179 ) ;
 assign wire29960 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire29961 = ( pi17  &  pi25  &  (~ pi16)  &  wire178 ) ;
 assign wire29962 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire29963 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire29964 = ( pi17  &  (~ pi16)  &  wire343 ) | ( (~ pi17)  &  (~ pi16)  &  wire343 ) ;
 assign wire29965 = ( wire29964 ) | ( nv620  &  wire29963 ) ;
 assign wire29967 = ( wire6095 ) | ( wire29965 ) | ( nv735  &  wire393 ) ;
 assign wire29968 = ( nv658  &  wire29959 ) | ( nv699  &  wire29961 ) ;
 assign wire29970 = ( nv717  &  wire812 ) | ( nv679  &  wire29960 ) ;
 assign wire29972 = ( (~ pi15)  &  (~ ni10)  &  wire289 ) ;
 assign wire29973 = ( (~ ni10)  &  pi15 ) ;
 assign wire29975 = ( pi22  &  pi25  &  (~ ni34) ) ;
 assign wire29977 = ( wire395  &  wire766  &  wire29975 ) ;
 assign wire29979 = ( wire395  &  wire459  &  wire766 ) ;
 assign wire29981 = ( wire395  &  wire459  &  wire617 ) ;
 assign wire29982 = ( (~ pi19)  &  (~ pi20)  &  pi25 ) | ( (~ pi19)  &  (~ pi20)  &  (~ ni34) ) ;
 assign wire29985 = ( (~ nv6428)  &  (~ n_n12655)  &  wire485 ) | ( (~ n_n12655)  &  wire485  &  nv858 ) ;
 assign wire29987 = ( pi22  &  (~ pi25)  &  wire395  &  wire766 ) ;
 assign wire29990 = ( pi22  &  (~ pi25)  &  wire395  &  wire617 ) ;
 assign wire29992 = ( wire395  &  wire225  &  wire617 ) ;
 assign wire29993 = ( (~ ni34)  &  pi15 ) ;
 assign wire29994 = ( pi25  &  wire152  &  wire154  &  wire29993 ) ;
 assign wire29995 = ( (~ pi25)  &  wire395  &  wire179 ) ;
 assign wire29996 = ( pi25  &  (~ ni34)  &  wire395  &  wire179 ) ;
 assign wire29997 = ( pi19  &  (~ pi20)  &  pi25  &  wire395 ) ;
 assign wire29998 = ( wire184 ) | ( ni34  &  nv942 ) ;
 assign wire29999 = ( (~ pi25)  &  wire178  &  wire395 ) ;
 assign wire30001 = ( wire395  &  wire910 ) | ( wire395  &  wire6127 ) ;
 assign wire30003 = ( (~ pi25)  &  pi15  &  wire152  &  wire154 ) ;
 assign wire30004 = ( (~ pi19)  &  pi21  &  pi20  &  wire459 ) ;
 assign wire30006 = ( pi22  &  (~ pi25)  &  wire766 ) ;
 assign wire30007 = ( wire766  &  wire6172 ) | ( (~ nv6428)  &  wire459  &  wire766 ) ;
 assign wire30010 = ( wire816 ) | ( wire6077 ) | ( nv988  &  wire30007 ) ;
 assign wire30011 = ( wire910  &  nv979 ) | ( wire1038  &  wire30004 ) ;
 assign wire30013 = ( wire811  &  nv1556 ) | ( nv1577  &  wire30006 ) ;
 assign wire30014 = ( wire30010 ) | ( wire30011 ) | ( wire30013 ) ;
 assign wire30016 = ( (~ pi17)  &  (~ pi16)  &  wire459  &  wire617 ) ;
 assign wire30018 = ( (~ pi17)  &  pi22  &  (~ pi25)  &  (~ pi16) ) ;
 assign wire30019 = ( pi19  &  pi21  &  pi20  &  wire30018 ) ;
 assign wire30023 = ( pi21  &  pi20  &  wire459  &  wire344 ) ;
 assign wire30025 = ( (~ pi17)  &  (~ pi25)  &  (~ pi16)  &  wire179 ) ;
 assign wire30026 = ( pi25  &  (~ ni34)  &  wire302  &  wire179 ) ;
 assign wire30027 = ( (~ pi17)  &  (~ pi16)  &  wire1014 ) ;
 assign wire30028 = ( wire184 ) | ( ni34  &  nv883 ) ;
 assign wire30029 = ( pi22  &  (~ pi25)  &  wire211  &  wire344 ) ;
 assign wire30031 = ( (~ pi17)  &  (~ pi16)  &  wire617 ) ;
 assign wire30032 = ( (~ pi16)  &  wire6156 ) | ( (~ pi16)  &  wire6157 ) ;
 assign wire30033 = ( wire184 ) | ( ni34  &  nv873 ) ;
 assign wire30034 = ( (~ pi20)  &  (~ pi25)  &  (~ pi16)  &  wire153 ) ;
 assign wire30035 = ( pi17  &  (~ ni34) ) | ( pi17  &  pi22  &  pi25 ) ;
 assign wire30036 = ( (~ pi19)  &  pi21  &  pi20  &  wire30035 ) ;
 assign wire30038 = ( pi17  &  pi22  &  (~ pi25) ) ;
 assign wire30040 = ( pi17  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire30041 = ( wire6172  &  wire30040 ) | ( (~ nv6428)  &  wire459  &  wire30040 ) ;
 assign wire30042 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi25 ) ;
 assign wire30043 = ( pi17  &  pi19  &  pi25 ) | ( pi17  &  pi19  &  (~ ni34) ) ;
 assign wire30044 = ( pi17  &  pi25  &  (~ ni34)  &  wire178 ) ;
 assign wire30046 = ( pi17  &  (~ pi25)  &  wire178 ) ;
 assign wire30047 = ( pi17  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire30049 = ( wire272  &  (~ pi25) ) ;
 assign wire30051 = ( wire6062 ) | ( wire6066 ) | ( pi17  &  wire816 ) ;
 assign wire30052 = ( wire30051 ) | ( nv928  &  wire6170 ) | ( nv928  &  wire6171 ) ;
 assign wire30054 = ( wire6059 ) | ( wire30052 ) | ( nv1445  &  wire30049 ) ;
 assign wire30055 = ( wire30054 ) | ( nv910  &  wire30044 ) ;
 assign wire30057 = ( wire1039  &  wire30036 ) | ( nv1403  &  wire30046 ) ;
 assign wire30058 = ( wire30055 ) | ( wire30057 ) | ( nv919  &  wire30041 ) ;
 assign wire30059 = ( wire6056 ) | ( wire6202  &  wire30042 ) | ( wire29864  &  wire30042 ) ;
 assign wire30060 = ( wire6154 ) | ( wire6155 ) | ( wire302  &  wire1108 ) ;
 assign wire30061 = ( wire483  &  wire30031 ) | ( wire483  &  wire211  &  wire344 ) ;
 assign wire30063 = ( wire6049 ) | ( wire30060 ) | ( wire30061 ) ;
 assign wire30064 = ( wire6041 ) | ( nv890  &  wire30026 ) ;
 assign wire30068 = ( wire6040 ) | ( wire6050 ) | ( nv1359  &  wire30025 ) ;
 assign wire30069 = ( wire6038 ) | ( wire6047 ) | ( wire30063 ) | ( wire30064 ) ;
 assign wire30071 = ( wire6042 ) | ( wire6198  &  wire30027 ) | ( wire29857  &  wire30027 ) ;
 assign wire30072 = ( wire30068 ) | ( wire30069 ) | ( nv1380  &  wire30019 ) ;
 assign wire30073 = ( wire30071 ) | ( wire6450  &  wire30029 ) | ( wire30028  &  wire30029 ) ;
 assign wire30074 = ( wire30072 ) | ( (~ pi16)  &  wire30058 ) | ( (~ pi16)  &  wire30059 ) ;
 assign wire30075 = ( wire395  &  wire1108 ) | ( wire395  &  wire483  &  wire766 ) ;
 assign wire30076 = ( wire6035 ) | ( wire395  &  wire483  &  wire617 ) ;
 assign wire30078 = ( wire30075 ) | ( wire30076 ) | ( wire395  &  wire1210 ) ;
 assign wire30079 = ( nv997  &  wire29985 ) | ( nv997  &  wire29994 ) ;
 assign wire30081 = ( wire6032 ) | ( wire30078 ) | ( wire30079 ) ;
 assign wire30084 = ( wire6019 ) | ( nv1490  &  wire29987 ) ;
 assign wire30085 = ( nv968  &  wire29992 ) | ( nv959  &  wire29996 ) ;
 assign wire30086 = ( wire6016 ) | ( wire6017 ) | ( wire6030 ) | ( wire30081 ) ;
 assign wire30090 = ( wire6018 ) | ( wire6025 ) | ( wire30084 ) | ( wire30085 ) ;
 assign wire30091 = ( wire6028 ) | ( wire30086 ) | ( nv1533  &  wire29990 ) ;
 assign wire30093 = ( wire6027 ) | ( wire30090 ) | ( wire30091 ) ;
 assign wire30094 = ( wire30093 ) | ( wire403  &  wire6074 ) | ( wire403  &  wire30014 ) ;
 assign wire30096 = ( pi25  &  wire1071 ) | ( (~ ni34)  &  wire1071 ) ;
 assign wire30099 = ( wire459  &  wire766  &  wire507 ) ;
 assign wire30100 = ( (~ pi19)  &  (~ pi20)  &  pi25 ) | ( (~ pi19)  &  (~ pi20)  &  (~ ni34) ) ;
 assign wire30103 = ( wire459  &  wire507  &  wire617 ) ;
 assign wire30106 = ( pi22  &  (~ pi25)  &  wire766  &  wire507 ) ;
 assign wire30108 = ( wire225  &  wire766  &  wire507 ) ;
 assign wire30111 = ( pi22  &  (~ pi25)  &  wire507  &  wire617 ) ;
 assign wire30113 = ( wire225  &  wire507  &  wire617 ) ;
 assign wire30114 = ( (~ ni34)  &  (~ pi15) ) ;
 assign wire30115 = ( pi25  &  wire152  &  wire154  &  wire30114 ) ;
 assign wire30117 = ( (~ pi25)  &  wire179  &  wire507 ) ;
 assign wire30118 = ( pi25  &  (~ ni34)  &  wire179  &  wire507 ) ;
 assign wire30119 = ( pi19  &  (~ pi20)  &  pi25  &  wire507 ) ;
 assign wire30121 = ( (~ pi25)  &  wire178  &  wire507 ) ;
 assign wire30123 = ( wire910  &  wire507 ) | ( wire507  &  wire6127 ) ;
 assign wire30125 = ( (~ pi25)  &  (~ pi15)  &  wire152  &  wire154 ) ;
 assign wire30126 = ( (~ pi19)  &  pi21  &  pi20  &  wire459 ) ;
 assign wire30128 = ( pi22  &  (~ pi25)  &  wire766 ) ;
 assign wire30129 = ( wire766  &  wire6172 ) | ( (~ nv6428)  &  wire459  &  wire766 ) ;
 assign wire30131 = ( wire6135 ) | ( wire816 ) ;
 assign wire30133 = ( wire910  &  nv817 ) | ( wire1112  &  wire30126 ) ;
 assign wire30134 = ( wire30131 ) | ( wire30133 ) | ( nv835  &  wire30129 ) ;
 assign wire30135 = ( wire811  &  nv1249 ) | ( nv1270  &  wire30128 ) ;
 assign wire30138 = ( (~ pi17)  &  (~ pi16)  &  wire459  &  wire617 ) ;
 assign wire30140 = ( (~ pi17)  &  pi22  &  (~ pi25)  &  (~ pi16) ) ;
 assign wire30142 = ( (~ pi17)  &  (~ pi16)  &  wire617 ) ;
 assign wire30146 = ( (~ pi17)  &  (~ pi25)  &  (~ pi16)  &  wire179 ) ;
 assign wire30147 = ( pi25  &  (~ ni34)  &  wire302  &  wire179 ) ;
 assign wire30148 = ( pi21  &  pi20  &  wire459  &  wire344 ) ;
 assign wire30149 = ( (~ pi17)  &  (~ pi16)  &  wire1014 ) ;
 assign wire30150 = ( wire184 ) | ( ni34  &  nv644 ) ;
 assign wire30151 = ( pi22  &  (~ pi25)  &  wire211  &  wire344 ) ;
 assign wire30152 = ( pi21  &  pi20  &  wire225  &  wire344 ) ;
 assign wire30153 = ( (~ pi17)  &  (~ pi16)  &  wire617 ) ;
 assign wire30154 = ( (~ pi16)  &  wire6156 ) | ( (~ pi16)  &  wire6157 ) ;
 assign wire30156 = ( (~ pi20)  &  (~ pi25)  &  (~ pi16)  &  wire153 ) ;
 assign wire30157 = ( pi17  &  (~ ni34) ) | ( pi17  &  pi22  &  pi25 ) ;
 assign wire30158 = ( (~ pi19)  &  pi21  &  pi20  &  wire30157 ) ;
 assign wire30160 = ( pi17  &  pi22  &  (~ pi25) ) ;
 assign wire30162 = ( pi17  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire30163 = ( wire6172  &  wire30162 ) | ( (~ nv6428)  &  wire459  &  wire30162 ) ;
 assign wire30164 = ( pi17  &  pi19  &  pi25 ) | ( pi17  &  pi19  &  (~ ni34) ) ;
 assign wire30165 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi25 ) ;
 assign wire30166 = ( pi17  &  pi25  &  (~ ni34)  &  wire178 ) ;
 assign wire30168 = ( pi17  &  (~ pi25)  &  wire178 ) ;
 assign wire30169 = ( pi17  &  (~ pi19)  &  pi21  &  pi20 ) ;
 assign wire30171 = ( wire272  &  (~ pi25) ) ;
 assign wire30173 = ( wire6165 ) | ( wire6169 ) | ( pi17  &  wire816 ) ;
 assign wire30174 = ( wire30173 ) | ( nv735  &  wire6170 ) | ( nv735  &  wire6171 ) ;
 assign wire30176 = ( wire6161 ) | ( wire30174 ) | ( nv1138  &  wire30171 ) ;
 assign wire30177 = ( wire30176 ) | ( nv699  &  wire30166 ) ;
 assign wire30178 = ( wire30177 ) | ( nv717  &  wire30163 ) ;
 assign wire30179 = ( wire1092  &  wire30158 ) | ( nv1096  &  wire30168 ) ;
 assign wire30181 = ( wire6159 ) | ( wire6731  &  wire30165 ) | ( wire29769  &  wire30165 ) ;
 assign wire30182 = ( wire6154 ) | ( wire6155 ) | ( wire302  &  wire1108 ) ;
 assign wire30183 = ( wire483  &  wire30153 ) | ( wire483  &  wire211  &  wire344 ) ;
 assign wire30185 = ( wire30182 ) | ( wire30183 ) | ( nv620  &  wire30154 ) ;
 assign wire30187 = ( wire6140 ) | ( wire30185 ) | ( nv1009  &  wire30156 ) ;
 assign wire30188 = ( wire30187 ) | ( ni34  &  wire30152 ) | ( (~ wire785)  &  wire30152 ) ;
 assign wire30189 = ( wire6143 ) | ( nv658  &  wire30147 ) ;
 assign wire30191 = ( wire6145 ) | ( wire225  &  nv679  &  wire30142 ) ;
 assign wire30192 = ( wire30188 ) | ( wire30189 ) | ( wire1057  &  wire30138 ) ;
 assign wire30194 = ( wire30191 ) | ( wire30192 ) | ( nv1052  &  wire30146 ) ;
 assign wire30195 = ( wire6138 ) | ( wire6655  &  wire30149 ) | ( wire29762  &  wire30149 ) ;
 assign wire30197 = ( wire507  &  wire1108 ) | ( wire483  &  wire766  &  wire507 ) ;
 assign wire30198 = ( wire6122 ) | ( wire483  &  wire507  &  wire617 ) ;
 assign wire30200 = ( wire30197 ) | ( wire30198 ) | ( wire507  &  wire1210 ) ;
 assign wire30202 = ( wire6103 ) | ( wire6111 ) | ( wire30200 ) ;
 assign wire30204 = ( nv764  &  wire30108 ) | ( nv750  &  wire30123 ) ;
 assign wire30205 = ( wire6119 ) | ( wire30202 ) | ( wire1070  &  wire30099 ) ;
 assign wire30208 = ( nv1183  &  wire30106 ) | ( nv1162  &  wire30121 ) ;
 assign wire30209 = ( wire6105 ) | ( wire30204 ) | ( wire30205 ) | ( wire30208 ) ;
 assign wire30210 = ( nv797  &  wire30113 ) | ( nv779  &  wire30118 ) ;
 assign wire30212 = ( wire30209 ) | ( wire30210 ) | ( wire1008  &  wire30103 ) ;
 assign wire30213 = ( nv1226  &  wire30111 ) | ( nv1205  &  wire30117 ) ;
 assign wire30216 = ( wire6114 ) | ( wire6123 ) | ( wire30212 ) | ( wire30213 ) ;
 assign wire30217 = ( (~ wire289)  &  (~ ni10) ) ;
 assign wire30218 = ( wire289  &  wire343  &  wire29937 ) | ( wire289  &  wire343  &  wire29940 ) ;
 assign wire30219 = ( wire30218 ) | ( wire6013 ) ;
 assign wire30220 = ( wire30219 ) | ( wire311  &  nv997  &  wire29943 ) ;
 assign wire30223 = ( nv890  &  wire29894 ) | ( nv910  &  wire29902 ) ;
 assign wire30224 = ( wire6001 ) | ( wire6004 ) | ( wire6007 ) | ( wire30220 ) ;
 assign wire30226 = ( nv979  &  wire29890 ) | ( nv959  &  wire29898 ) ;
 assign wire30227 = ( nv899  &  wire29910 ) | ( nv968  &  wire29918 ) ;
 assign wire30228 = ( nv988  &  wire29929 ) | ( nv919  &  wire29932 ) ;
 assign wire30231 = ( wire6003 ) | ( wire30223 ) | ( wire30224 ) | ( wire30228 ) ;
 assign wire30232 = ( wire5999 ) | ( wire30226 ) | ( wire30227 ) ;
 assign wire30235 = ( wire6011 ) | ( wire6012 ) | ( wire30231 ) | ( wire30232 ) ;
 assign wire30236 = ( wire30235 ) | ( (~ ni10)  &  (~ wire289)  &  n_n12641 ) ;
 assign wire30238 = ( pi15  &  (~ pi16) ) ;
 assign wire30240 = ( pi17  &  (~ wire289)  &  wire178  &  wire30238 ) ;
 assign wire30241 = ( pi15  &  (~ pi16) ) ;
 assign wire30243 = ( pi17  &  (~ wire289)  &  wire180  &  wire30241 ) ;
 assign wire30246 = ( (~ pi16)  &  pi15  &  (~ wire289)  &  wire272 ) ;
 assign wire30248 = ( pi17  &  (~ pi16)  &  pi15 ) ;
 assign wire30250 = ( (~ wire289)  &  pi15 ) ;
 assign wire30253 = ( pi15  &  (~ wire289)  &  wire484 ) ;
 assign wire30254 = ( pi17  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire30257 = ( (~ wire289)  &  wire180  &  wire403 ) ;
 assign wire30259 = ( (~ wire289)  &  wire178  &  wire403 ) ;
 assign wire30260 = ( (~ pi17)  &  pi19  &  pi16  &  pi15 ) ;
 assign wire30263 = ( (~ wire289)  &  wire395  &  wire182 ) ;
 assign wire30265 = ( (~ wire289)  &  wire395  &  wire179 ) ;
 assign wire30267 = ( pi15  &  (~ wire289)  &  wire325 ) ;
 assign wire30268 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire30270 = ( (~ wire289)  &  pi15 ) ;
 assign wire30272 = ( (~ pi20)  &  (~ wire289)  &  wire226  &  wire153 ) ;
 assign wire30273 = ( pi20  &  (~ wire289)  &  wire226  &  wire153 ) ;
 assign wire30275 = ( pi15  &  (~ wire289)  &  wire152  &  wire154 ) ;
 assign wire30277 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire178 ) ;
 assign wire30279 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire180 ) ;
 assign wire30280 = ( (~ pi15)  &  (~ pi16) ) ;
 assign wire30282 = ( pi17  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire30283 = ( (~ pi17)  &  pi19  &  pi16  &  (~ pi15) ) ;
 assign wire30285 = ( pi17  &  pi16  &  (~ pi15)  &  wire178 ) ;
 assign wire30286 = ( pi17  &  pi16  &  (~ pi15)  &  wire180 ) ;
 assign wire30287 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire179 ) ;
 assign wire30288 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire182 ) ;
 assign wire30289 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire30290 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire30291 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire30292 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire30293 = ( wire230  &  wire30282 ) | ( wire230  &  wire30283 ) ;
 assign wire30294 = ( wire230  &  wire913 ) | ( (~ pi16)  &  (~ pi15)  &  wire230 ) ;
 assign wire30296 = ( wire30293 ) | ( wire30294 ) | ( nv1291  &  wire586 ) ;
 assign wire30297 = ( wire30296 ) | ( nv1138  &  wire272  &  wire30280 ) ;
 assign wire30299 = ( nv1183  &  wire1324 ) | ( nv1162  &  wire1327 ) ;
 assign wire30301 = ( wire6401 ) | ( wire6402 ) | ( wire30297 ) | ( wire30299 ) ;
 assign wire30302 = ( nv1096  &  wire30277 ) | ( nv1052  &  wire30289 ) ;
 assign wire30304 = ( nv1117  &  wire30279 ) | ( nv1249  &  wire30285 ) ;
 assign wire30305 = ( nv1270  &  wire30286 ) | ( nv1205  &  wire30287 ) ;
 assign wire30306 = ( nv1226  &  wire30288 ) | ( nv1073  &  wire30290 ) ;
 assign wire30307 = ( wire30301 ) | ( wire30302 ) | ( wire30304 ) ;
 assign wire30308 = ( wire30306 ) | ( wire30305 ) ;
 assign wire30309 = ( ni34  &  wire289 ) | ( (~ wire289)  &  wire230  &  wire30248 ) ;
 assign wire30310 = ( (~ wire289)  &  wire230  &  wire30254 ) | ( (~ wire289)  &  wire230  &  wire30260 ) ;
 assign wire30311 = ( (~ wire289)  &  wire915  &  wire230 ) | ( (~ wire289)  &  wire230  &  wire30268 ) ;
 assign wire30313 = ( wire30309 ) | ( wire30310 ) | ( wire30311 ) ;
 assign wire30314 = ( wire30313 ) | ( wire184  &  wire30275 ) | ( wire6475  &  wire30275 ) ;
 assign wire30315 = ( wire30314 ) | ( nv1445  &  wire30246 ) ;
 assign wire30316 = ( wire30315 ) | ( wire6366  &  wire30267 ) | ( wire30033  &  wire30267 ) ;
 assign wire30317 = ( nv1403  &  wire30240 ) | ( nv1490  &  wire30273 ) ;
 assign wire30318 = ( wire6351 ) | ( wire587  &  nv1359  &  wire30250 ) ;
 assign wire30321 = ( nv1424  &  wire30243 ) | ( nv1380  &  wire30253 ) ;
 assign wire30322 = ( nv1577  &  wire30257 ) | ( nv1556  &  wire30259 ) ;
 assign wire30323 = ( wire6355 ) | ( wire30316 ) | ( nv1533  &  wire30263 ) ;
 assign wire30326 = ( wire6354 ) | ( wire30317 ) | ( wire30318 ) | ( wire30321 ) ;
 assign wire30327 = ( wire30322 ) | ( wire30323 ) | ( wire30326 ) ;
 assign wire30328 = ( (~ ni2)  &  (~ ni3)  &  wire265 ) ;
 assign wire30329 = ( ni2  &  ni34 ) | ( (~ ni2)  &  ni3  &  ni34 ) ;
 assign wire30332 = ( wire5964 ) | ( wire5966 ) | ( wire30329 ) ;
 assign wire30333 = ( wire5965 ) | ( wire5967 ) | ( nv2066  &  wire30328 ) ;
 assign wire30336 = ( wire5963 ) | ( wire5968 ) | ( wire30332 ) | ( wire30333 ) ;
 assign wire30337 = ( (~ ni2)  &  (~ ni3)  &  (~ ni9) ) | ( (~ ni2)  &  (~ ni3)  &  (~ ni10) ) ;
 assign wire30338 = ( ni9  &  (~ ni33)  &  ni29 ) | ( (~ ni33)  &  ni10  &  ni29 ) ;
 assign wire30340 = ( (~ wire636)  &  wire30337  &  wire30338 ) ;
 assign wire30342 = ( (~ ni9)  &  ni10 ) | ( ni9  &  (~ ni10) ) ;
 assign wire30344 = ( (~ pi24)  &  ni8  &  wire510  &  wire30342 ) ;
 assign wire30346 = ( (~ ni9)  &  ni8 ) | ( (~ ni10)  &  ni8 ) ;
 assign wire30348 = ( (~ pi24)  &  (~ ni7)  &  wire510  &  wire30346 ) ;
 assign wire30349 = ( (~ ni2)  &  (~ ni3)  &  (~ ni7) ) ;
 assign wire30351 = ( (~ ni33)  &  ni29  &  (~ wire636)  &  wire30349 ) ;
 assign wire30352 = ( (~ ni2)  &  (~ ni3)  &  ni7 ) ;
 assign wire30354 = ( (~ ni9)  &  ni10  &  wire30352 ) | ( ni9  &  (~ ni10)  &  wire30352 ) ;
 assign wire30356 = ( ni9  &  (~ ni10) ) ;
 assign wire30358 = ( ni9  &  (~ ni10)  &  (~ ni7) ) ;
 assign wire30359 = ( wire5960 ) | ( wire5961  &  wire30340 ) | ( wire5962  &  wire30340 ) ;
 assign wire30360 = ( wire5961  &  wire30344 ) | ( wire5962  &  wire30344 ) | ( (~ wire5961)  &  (~ wire5962)  &  wire30348 ) ;
 assign wire30362 = ( wire5961  &  wire30356 ) | ( wire5962  &  wire30356 ) | ( (~ wire5961)  &  (~ wire5962)  &  wire30358 ) ;
 assign wire30364 = ( wire30362 ) | ( (~ n_n429)  &  wire30351 ) | ( n_n429  &  wire30354 ) ;
 assign wire30367 = ( ni44  &  ni42 ) ;
 assign wire30368 = ( (~ ni43)  &  ni42  &  (~ ni44) ) ;
 assign wire30369 = ( nv2176  &  wire30367 ) | ( (~ wire621)  &  wire30367 ) | ( nv2176  &  wire30368 ) ;
 assign wire30370 = ( wire5945 ) | ( wire30369 ) | ( n_n13643  &  nv2176 ) ;
 assign wire30371 = ( (~ ni43)  &  (~ ni41)  &  ni44 ) ;
 assign wire30372 = ( ni43  &  (~ ni41)  &  nv2176 ) | ( (~ ni41)  &  (~ ni44)  &  nv2176 ) ;
 assign wire30374 = ( wire5914 ) | ( wire177  &  wire216 ) | ( wire177  &  wire5917 ) ;
 assign wire30375 = ( pi17  &  (~ pi16)  &  pi15 ) ;
 assign wire30378 = ( wire510  &  wire180  &  (~ wire399) ) ;
 assign wire30379 = ( wire631  &  wire30375  &  wire30378 ) ;
 assign wire30380 = ( ni43  &  (~ ni41)  &  (~ ni44) ) | ( (~ ni43)  &  (~ ni42)  &  (~ ni41)  &  (~ ni44) ) ;
 assign wire30381 = ( ni43  &  ni42  &  (~ ni41)  &  ni44 ) | ( (~ ni43)  &  (~ ni42)  &  (~ ni41)  &  ni44 ) ;
 assign wire30382 = ( wire5897 ) | ( ni43  &  n_n11076 ) | ( ni42  &  n_n11076 ) ;
 assign wire30383 = ( wire5837 ) | ( wire1194  &  wire880 ) | ( wire880  &  wire5839 ) ;
 assign wire30384 = ( wire177  &  wire322 ) | ( wire177  &  wire5841 ) | ( wire177  &  wire5842 ) ;
 assign wire30385 = ( pi17  &  (~ pi16)  &  pi15 ) ;
 assign wire30388 = ( wire510  &  wire178  &  (~ wire399) ) ;
 assign wire30389 = ( wire631  &  wire30385  &  wire30388 ) ;
 assign wire30390 = ( pi15  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30392 = ( (~ wire399)  &  wire631  &  wire30390 ) ;
 assign wire30393 = ( pi17  &  (~ pi16)  &  wire324  &  wire30392 ) ;
 assign wire30397 = ( (~ ni45)  &  (~ pi21) ) ;
 assign wire30399 = ( pi17  &  (~ pi16)  &  pi15 ) ;
 assign wire30402 = ( wire510  &  (~ wire399)  &  wire631  &  wire30399 ) ;
 assign wire30404 = ( wire5847 ) | ( wire177  &  wire216 ) | ( wire177  &  wire5917 ) ;
 assign wire30407 = ( wire510  &  wire180  &  (~ wire399) ) ;
 assign wire30408 = ( wire403  &  wire631  &  wire30407 ) ;
 assign wire30409 = ( wire5883 ) | ( wire1194  &  wire880 ) | ( wire880  &  wire5887 ) ;
 assign wire30410 = ( wire177  &  wire322 ) | ( wire177  &  wire5893 ) | ( wire177  &  wire5894 ) ;
 assign wire30413 = ( wire510  &  wire178  &  (~ wire399) ) ;
 assign wire30414 = ( wire403  &  wire631  &  wire30413 ) ;
 assign wire30416 = ( wire1111 ) | ( wire706 ) | ( wire5839 ) | ( wire5889 ) ;
 assign wire30417 = ( pi15  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30419 = ( (~ wire399)  &  wire631  &  wire30417 ) ;
 assign wire30422 = ( wire5804 ) | ( wire176  &  wire216 ) | ( wire176  &  wire5917 ) ;
 assign wire30423 = ( wire5796 ) | ( wire1194  &  wire887 ) | ( wire887  &  wire5839 ) ;
 assign wire30424 = ( wire176  &  wire322 ) | ( wire176  &  wire5800 ) | ( wire176  &  wire5801 ) ;
 assign wire30425 = ( wire378 ) | ( wire240  &  wire182 ) | ( wire182  &  wire5802 ) ;
 assign wire30426 = ( wire378 ) | ( nv10727  &  wire324 ) | ( wire237  &  wire324 ) ;
 assign wire30427 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire30430 = ( wire510  &  (~ wire399)  &  wire631  &  wire30427 ) ;
 assign wire30431 = ( wire314 ) | ( n_n11076  &  wire310 ) | ( wire1319  &  wire310 ) ;
 assign wire30432 = ( wire1111 ) | ( wire706 ) | ( wire5924 ) | ( wire5926 ) ;
 assign wire30433 = ( pi15  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30435 = ( (~ wire399)  &  wire631  &  wire30433 ) ;
 assign wire30436 = ( pi20  &  (~ pi16)  &  wire153  &  wire30435 ) ;
 assign wire30438 = ( wire5386 ) | ( wire176  &  wire216 ) | ( wire176  &  wire5917 ) ;
 assign wire30439 = ( nv2348  &  wire310 ) | ( ni36  &  wire216 ) ;
 assign wire30441 = ( wire5375 ) | ( wire1194  &  wire887 ) | ( wire887  &  wire5887 ) ;
 assign wire30442 = ( wire176  &  wire322 ) | ( wire176  &  wire5377 ) | ( wire176  &  wire5378 ) ;
 assign wire30444 = ( wire1111 ) | ( wire706 ) | ( wire5887 ) | ( wire5889 ) ;
 assign wire30445 = ( pi19  &  pi20  &  wire162 ) | ( (~ pi19)  &  pi20  &  wire162 ) | ( pi19  &  (~ pi20)  &  wire159 ) | ( (~ pi19)  &  (~ pi20)  &  wire159 ) ;
 assign wire30446 = ( wire5167 ) | ( wire30445 ) ;
 assign wire30449 = ( pi19  &  pi20  &  wire162 ) | ( (~ pi19)  &  pi20  &  wire162 ) | ( pi19  &  (~ pi20)  &  wire159 ) | ( (~ pi19)  &  (~ pi20)  &  wire159 ) ;
 assign wire30450 = ( wire30449 ) | ( nv10727  &  wire324 ) | ( wire237  &  wire324 ) ;
 assign wire30451 = ( pi20  &  nv10727  &  wire151 ) | ( (~ pi20)  &  nv10727  &  wire151 ) | ( pi20  &  wire237  &  wire151 ) | ( (~ pi20)  &  wire237  &  wire151 ) ;
 assign wire30452 = ( wire30451 ) | ( wire30450 ) ;
 assign wire30455 = ( wire510  &  wire395  &  (~ wire399)  &  wire631 ) ;
 assign wire30456 = ( pi15  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30458 = ( (~ wire399)  &  wire631  &  wire30456 ) ;
 assign wire30461 = ( wire510  &  (~ wire399)  &  wire403  &  wire631 ) ;
 assign wire30463 = ( wire510  &  (~ wire399)  &  wire631 ) ;
 assign wire30465 = ( wire1181 ) | ( nv2348  &  wire347 ) ;
 assign wire30467 = ( wire5407 ) | ( wire30465 ) | ( (~ ni35)  &  n_n10809 ) ;
 assign wire30468 = ( pi17  &  pi16  &  wire180 ) ;
 assign wire30470 = ( wire1181 ) | ( wire5401 ) | ( wire5402 ) ;
 assign wire30472 = ( pi17  &  pi16  &  wire178 ) ;
 assign wire30473 = ( wire314 ) | ( wire310  &  wire5939 ) | ( wire310  &  wire30370 ) ;
 assign wire30475 = ( wire1184 ) | ( wire5366 ) | ( wire5367 ) ;
 assign wire30477 = ( (~ ni34)  &  wire179 ) | ( (~ ni33)  &  wire179 ) | ( (~ nv6428)  &  wire179 ) ;
 assign wire30478 = ( wire1184 ) | ( nv2348  &  wire346 ) ;
 assign wire30480 = ( wire5380 ) | ( wire30478 ) | ( ni35  &  n_n10835 ) ;
 assign wire30482 = ( wire378 ) | ( nv10727  &  wire179 ) | ( wire237  &  wire179 ) ;
 assign wire30483 = ( wire30482 ) | ( wire304  &  wire182 ) | ( wire182  &  wire5902 ) ;
 assign wire30484 = ( wire30483 ) | ( (~ n_n12619)  &  wire182  &  nv2373 ) ;
 assign wire30485 = ( wire1341 ) | ( pi17  &  pi16  &  wire438 ) ;
 assign wire30487 = ( wire5072 ) | ( wire304  &  wire1024 ) | ( wire1024  &  wire5190 ) ;
 assign wire30489 = ( wire5070 ) | ( wire5075 ) | ( wire30485 ) | ( wire30487 ) ;
 assign wire30491 = ( (~ pi15)  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30493 = ( (~ wire399)  &  wire631  &  wire30491 ) ;
 assign wire30494 = ( wire314 ) | ( wire5499 ) | ( nv2240  &  wire346 ) ;
 assign wire30496 = ( wire5500 ) | ( wire30494 ) | ( (~ ni35)  &  n_n10896 ) ;
 assign wire30497 = ( pi17  &  (~ pi16)  &  wire180 ) ;
 assign wire30499 = ( wire1186 ) | ( wire5504 ) | ( wire5505 ) ;
 assign wire30501 = ( pi17  &  (~ pi16)  &  wire178 ) ;
 assign wire30502 = ( ni36  &  wire216 ) | ( wire310  &  nv2240 ) ;
 assign wire30503 = ( wire314 ) | ( wire5468 ) | ( wire347  &  nv2240 ) ;
 assign wire30505 = ( wire5469 ) | ( wire30503 ) | ( ni35  &  n_n10922 ) ;
 assign wire30507 = ( wire1183 ) | ( wire5473 ) | ( wire5474 ) ;
 assign wire30509 = ( wire378 ) | ( nv2252  &  wire182 ) ;
 assign wire30510 = ( wire378 ) | ( nv10727  &  wire324 ) | ( wire237  &  wire324 ) ;
 assign wire30511 = ( pi17  &  pi19  &  (~ pi16)  &  wire166 ) | ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire166 ) | ( (~ pi17)  &  (~ pi19)  &  (~ pi16)  &  wire166 ) ;
 assign wire30512 = ( wire30511 ) | ( wire294  &  wire304 ) | ( wire294  &  wire5211 ) ;
 assign wire30515 = ( wire5078 ) | ( wire5080 ) | ( wire5082 ) | ( wire30512 ) ;
 assign wire30517 = ( (~ pi15)  &  (~ ni2)  &  (~ ni3)  &  ni10 ) ;
 assign wire30519 = ( (~ wire399)  &  wire631  &  wire30517 ) ;
 assign wire30521 = ( wire510  &  (~ wire399)  &  wire631 ) ;
 assign wire30522 = ( wire303  &  (~ ni34) ) ;
 assign wire30524 = ( (~ ni33)  &  ni34 ) ;
 assign wire30525 = ( wire307 ) | ( wire315  &  nv2314 ) ;
 assign wire30526 = ( ni14  &  pi15 ) ;
 assign wire30527 = ( pi17  &  (~ pi16)  &  wire324  &  wire30526 ) ;
 assign wire30528 = ( ni36  &  wire216 ) | ( wire310  &  nv2790 ) ;
 assign wire30530 = ( wire307 ) | ( wire315  &  nv2534 ) ;
 assign wire30531 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30532 = ( wire30531  &  wire180 ) ;
 assign wire30534 = ( wire1195 ) | ( wire5591 ) | ( (~ wire205)  &  n_n10282 ) ;
 assign wire30536 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30537 = ( wire30536  &  wire178 ) ;
 assign wire30538 = ( ni36  &  wire216 ) | ( wire310  &  nv2602 ) ;
 assign wire30540 = ( wire307 ) | ( (~ wire157)  &  nv2930  &  wire30524 ) ;
 assign wire30541 = ( ni14  &  pi15 ) ;
 assign wire30542 = ( (~ pi20)  &  (~ pi16)  &  wire153  &  wire30541 ) ;
 assign wire30543 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire182 ) ;
 assign wire30544 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire179 ) ;
 assign wire30547 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire182 ) ;
 assign wire30548 = ( wire5724 ) | ( wire5723 ) ;
 assign wire30549 = ( wire176  &  wire321 ) | ( wire176  &  wire5728 ) | ( wire176  &  wire5729 ) ;
 assign wire30550 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire179 ) ;
 assign wire30552 = ( wire378 ) | ( pi20  &  wire152  &  wire307 ) | ( (~ pi20)  &  wire152  &  wire307 ) ;
 assign wire30553 = ( wire5317 ) | ( wire30552 ) ;
 assign wire30554 = ( nv2473  &  wire30544 ) | ( nv2963  &  wire30550 ) ;
 assign wire30557 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  ni14 ) ;
 assign wire30558 = ( ni36  &  wire216 ) | ( wire310  &  nv2622 ) ;
 assign wire30560 = ( wire5334 ) | ( wire307 ) ;
 assign wire30561 = ( ni14  &  pi15 ) ;
 assign wire30562 = ( pi20  &  (~ pi16)  &  wire153  &  wire30561 ) ;
 assign wire30563 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire180 ) ;
 assign wire30564 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire178 ) ;
 assign wire30566 = ( wire5710 ) | ( wire1049 ) ;
 assign wire30567 = ( ni34  &  (~ ni33)  &  wire180  &  (~ wire157) ) ;
 assign wire30568 = ( wire5704 ) | ( wire5703 ) ;
 assign wire30569 = ( wire177  &  wire321 ) | ( wire177  &  wire5708 ) | ( wire177  &  wire5709 ) ;
 assign wire30570 = ( ni34  &  (~ ni33)  &  wire178  &  (~ wire157) ) ;
 assign wire30572 = ( wire438 ) | ( pi20  &  wire151  &  wire307 ) | ( (~ pi20)  &  wire151  &  wire307 ) ;
 assign wire30573 = ( wire5327 ) | ( wire30572 ) ;
 assign wire30574 = ( nv2493  &  wire30564 ) | ( nv2995  &  wire30570 ) ;
 assign wire30577 = ( pi17  &  (~ pi16)  &  pi15  &  ni14 ) ;
 assign wire30578 = ( ni36  &  wire216 ) | ( wire310  &  nv2647 ) ;
 assign wire30579 = ( wire307 ) | ( wire315  &  wire5429 ) | ( wire315  &  wire30473 ) ;
 assign wire30580 = ( pi17  &  pi16  &  wire324  &  wire1069 ) ;
 assign wire30581 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire182 ) ;
 assign wire30584 = ( wire5557 ) | ( wire1013 ) ;
 assign wire30586 = ( wire1188 ) | ( wire5553 ) | ( nv2790  &  wire346 ) ;
 assign wire30588 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire182 ) ;
 assign wire30589 = ( wire5576 ) | ( wire1195  &  wire885 ) | ( wire885  &  wire5591 ) ;
 assign wire30590 = ( wire176  &  wire321 ) | ( wire176  &  wire5578 ) | ( wire176  &  wire5579 ) ;
 assign wire30592 = ( wire1188 ) | ( wire5565 ) | ( wire5566 ) ;
 assign wire30596 = ( wire378 ) | ( pi20  &  wire152  &  wire307 ) | ( (~ pi20)  &  wire152  &  wire307 ) ;
 assign wire30597 = ( wire30596 ) | ( wire5381  &  wire30581 ) | ( wire30480  &  wire30581 ) ;
 assign wire30598 = ( wire30597 ) | ( wire179  &  wire315  &  nv2359 ) ;
 assign wire30600 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  ni14 ) ;
 assign wire30601 = ( wire307 ) | ( wire315  &  nv2330 ) ;
 assign wire30602 = ( (~ pi20)  &  pi16  &  wire1069  &  wire153 ) ;
 assign wire30603 = ( wire307 ) | ( n_n10860  &  wire315 ) | ( wire315  &  wire30439 ) ;
 assign wire30604 = ( pi20  &  pi16  &  wire1069  &  wire153 ) ;
 assign wire30605 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire180 ) ;
 assign wire30610 = ( wire1179 ) | ( wire5601 ) | ( wire347  &  nv2790 ) ;
 assign wire30612 = ( ni34  &  (~ ni33)  &  wire180  &  (~ wire157) ) ;
 assign wire30613 = ( wire5589 ) | ( wire1195  &  wire883 ) | ( wire883  &  wire5591 ) ;
 assign wire30614 = ( wire177  &  wire321 ) | ( wire177  &  wire5593 ) | ( wire177  &  wire5594 ) ;
 assign wire30616 = ( wire1179 ) | ( wire5580 ) | ( wire5581 ) ;
 assign wire30620 = ( wire438 ) | ( pi20  &  wire151  &  wire307 ) | ( (~ pi20)  &  wire151  &  wire307 ) ;
 assign wire30621 = ( wire30620 ) | ( wire5409  &  wire30605 ) | ( wire30467  &  wire30605 ) ;
 assign wire30622 = ( wire30621 ) | ( wire178  &  nv2397  &  wire315 ) ;
 assign wire30624 = ( pi17  &  pi16  &  (~ pi15)  &  ni14 ) ;
 assign wire30626 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30628 = ( pi15  &  ni14  &  wire152  &  wire154 ) ;
 assign wire30629 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire180 ) ;
 assign wire30630 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire178 ) ;
 assign wire30631 = ( ni34  &  (~ ni33)  &  wire180  &  (~ wire157) ) ;
 assign wire30634 = ( wire438 ) | ( pi20  &  wire151  &  wire307 ) | ( (~ pi20)  &  wire151  &  wire307 ) ;
 assign wire30636 = ( wire5284 ) | ( wire30634 ) | ( nv2565  &  wire30630 ) ;
 assign wire30638 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30639 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire182 ) ;
 assign wire30640 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire179 ) ;
 assign wire30641 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire182 ) ;
 assign wire30644 = ( wire378 ) | ( pi20  &  wire152  &  wire307 ) | ( (~ pi20)  &  wire152  &  wire307 ) ;
 assign wire30646 = ( wire5271 ) | ( wire30644 ) | ( nv2545  &  wire30640 ) ;
 assign wire30648 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30649 = ( wire5653 ) | ( ni36  &  wire216 ) ;
 assign wire30650 = ( wire5486 ) | ( wire307 ) ;
 assign wire30651 = ( wire307 ) | ( wire238  &  n_n10412 ) | ( wire238  &  wire30538 ) ;
 assign wire30652 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire182 ) ;
 assign wire30653 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire179 ) ;
 assign wire30654 = ( wire314 ) | ( wire5639 ) | ( wire346  &  nv2622 ) ;
 assign wire30655 = ( wire5635 ) | ( wire30654 ) ;
 assign wire30657 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire182 ) ;
 assign wire30659 = ( wire314 ) | ( wire5629 ) | ( wire5630 ) | ( wire5639 ) ;
 assign wire30661 = ( ni34  &  (~ ni33)  &  (~ wire157)  &  wire179 ) ;
 assign wire30663 = ( wire378 ) | ( pi20  &  wire152  &  wire307 ) | ( (~ pi20)  &  wire152  &  wire307 ) ;
 assign wire30664 = ( wire30663 ) | ( wire5470  &  wire30652 ) | ( wire30505  &  wire30652 ) ;
 assign wire30665 = ( nv2235  &  wire30653 ) | ( nv2641  &  wire30661 ) ;
 assign wire30667 = ( wire307 ) | ( wire315  &  nv2220 ) ;
 assign wire30668 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire180 ) ;
 assign wire30669 = ( (~ ni34)  &  ni33  &  (~ ni32)  &  wire178 ) ;
 assign wire30670 = ( wire314 ) | ( wire5651 ) | ( wire347  &  nv2622 ) ;
 assign wire30671 = ( wire5642 ) | ( wire30670 ) ;
 assign wire30673 = ( ni34  &  (~ ni33)  &  wire180  &  (~ wire157) ) ;
 assign wire30675 = ( wire314 ) | ( wire5646 ) | ( wire5647 ) | ( wire5651 ) ;
 assign wire30677 = ( ni34  &  (~ ni33)  &  wire178  &  (~ wire157) ) ;
 assign wire30679 = ( wire438 ) | ( pi20  &  wire151  &  wire307 ) | ( (~ pi20)  &  wire151  &  wire307 ) ;
 assign wire30680 = ( wire30679 ) | ( wire5501  &  wire30668 ) | ( wire30496  &  wire30668 ) ;
 assign wire30681 = ( nv2276  &  wire30669 ) | ( nv2694  &  wire30677 ) ;
 assign wire30683 = ( wire5065 ) | ( wire5086 ) | ( wire5087 ) ;
 assign wire30685 = ( wire5064 ) | ( wire30683 ) | ( wire294  &  nv2627 ) ;
 assign wire30687 = ( wire1069  &  wire1341 ) | ( wire438  &  wire30626 ) ;
 assign wire30689 = ( wire5056 ) | ( wire30687 ) | ( ni14  &  wire1336 ) ;
 assign wire30691 = ( wire5044 ) | ( wire5058 ) | ( wire30689 ) ;
 assign wire30692 = ( wire5051 ) | ( wire5414  &  wire30602 ) | ( wire30601  &  wire30602 ) ;
 assign wire30696 = ( wire5045 ) | ( wire30692 ) | ( nv2793  &  wire30604 ) ;
 assign wire30697 = ( wire5046 ) | ( wire5047 ) | ( wire5049 ) | ( wire30691 ) ;
 assign wire30700 = ( wire5060 ) | ( wire5059 ) ;
 assign wire30701 = ( wire5048 ) | ( wire5050 ) | ( wire30696 ) | ( wire30697 ) ;
 assign wire30704 = ( wire5052 ) | ( wire5055 ) | ( wire30700 ) | ( wire30701 ) ;
 assign wire30705 = ( pi17  &  (~ pi16)  &  pi15  &  (~ ni14) ) ;
 assign wire30707 = ( pi17  &  (~ pi16)  &  pi15  &  (~ ni14) ) ;
 assign wire30708 = ( wire178  &  wire30707 ) ;
 assign wire30709 = ( pi17  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire30711 = ( pi17  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire30712 = ( wire30711  &  wire178 ) ;
 assign wire30713 = ( pi17  &  (~ pi16)  &  wire324  &  wire920 ) ;
 assign wire30714 = ( pi17  &  (~ pi16)  &  pi15  &  (~ ni14) ) ;
 assign wire30715 = ( (~ pi20)  &  (~ pi16)  &  wire153  &  wire920 ) ;
 assign wire30716 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  (~ ni14) ) ;
 assign wire30717 = ( pi20  &  (~ pi16)  &  wire153  &  wire920 ) ;
 assign wire30718 = ( (~ pi17)  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire30719 = ( pi17  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire30720 = ( pi15  &  (~ ni14)  &  wire152  &  wire154 ) ;
 assign wire30721 = ( pi17  &  (~ pi16)  &  wire180 ) ;
 assign wire30722 = ( pi17  &  (~ pi16)  &  wire178 ) ;
 assign wire30723 = ( pi17  &  pi19  &  (~ pi16)  &  wire166 ) | ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire166 ) | ( (~ pi17)  &  (~ pi19)  &  (~ pi16)  &  wire166 ) ;
 assign wire30726 = ( wire5030 ) | ( wire5032 ) | ( wire5034 ) | ( wire30723 ) ;
 assign wire30728 = ( wire5029 ) | ( wire30726 ) | ( nv2290  &  wire30721 ) ;
 assign wire30729 = ( pi17  &  pi16  &  wire180 ) ;
 assign wire30730 = ( pi17  &  pi16  &  wire178 ) ;
 assign wire30731 = ( wire378 ) | ( wire182  &  nv2373 ) ;
 assign wire30732 = ( wire1341 ) | ( pi17  &  pi16  &  wire438 ) ;
 assign wire30733 = ( wire30732 ) | ( nv2340  &  wire763 ) ;
 assign wire30735 = ( wire5040 ) | ( wire30733 ) | ( wire1309  &  nv2430 ) ;
 assign wire30737 = ( wire5037 ) | ( wire30735 ) | ( nv2411  &  wire30729 ) ;
 assign wire30738 = ( wire438  &  wire30714 ) | ( wire438  &  wire30719 ) ;
 assign wire30740 = ( wire5024 ) | ( wire30738 ) | ( (~ ni14)  &  wire1336 ) ;
 assign wire30742 = ( wire5015 ) | ( wire5022 ) | ( wire30740 ) ;
 assign wire30746 = ( wire5012 ) | ( wire5017 ) | ( wire5019 ) | ( wire30742 ) ;
 assign wire30748 = ( wire5011 ) | ( wire5013 ) | ( wire5014 ) | ( wire30746 ) ;
 assign wire30749 = ( wire5018 ) | ( wire852  &  wire30718 ) ;
 assign wire30752 = ( wire5025 ) | ( wire5026 ) | ( wire30748 ) | ( wire30749 ) ;
 assign wire30754 = ( wire510  &  (~ wire399)  &  (~ wire631) ) ;
 assign wire30755 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30756 = ( (~ pi16)  &  (~ ni13)  &  (~ ni14) ) | ( (~ pi15)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire30758 = ( (~ pi17)  &  pi25  &  wire30755  &  wire30756 ) ;
 assign wire30759 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30762 = ( wire593  &  wire387  &  wire263  &  wire30759 ) ;
 assign wire30764 = ( (~ pi16)  &  (~ ni13)  &  (~ ni14) ) | ( (~ pi15)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire30765 = ( pi15  &  (~ ni11)  &  (~ ni12)  &  wire30764 ) ;
 assign wire30767 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30770 = ( wire456  &  wire387  &  wire263  &  wire30767 ) ;
 assign wire30772 = ( (~ pi16)  &  (~ ni13)  &  (~ ni14) ) | ( (~ pi15)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire30773 = ( pi15  &  (~ ni11)  &  (~ ni12)  &  wire30772 ) ;
 assign wire30775 = ( pi16  &  pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30776 = ( (~ pi17)  &  pi25  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire30777 = ( wire30776  &  wire30775 ) ;
 assign wire30778 = ( wire5744 ) | ( wire757 ) ;
 assign wire30779 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30781 = ( (~ ni13)  &  (~ ni14)  &  wire593  &  wire30779 ) ;
 assign wire30782 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30784 = ( (~ ni13)  &  (~ ni14)  &  wire456  &  wire30782 ) ;
 assign wire30785 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30786 = ( (~ ni13)  &  (~ ni14)  &  wire30785 ) ;
 assign wire30788 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30789 = ( (~ ni13)  &  (~ ni14)  &  wire30788 ) ;
 assign wire30791 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30793 = ( (~ ni13)  &  (~ ni14)  &  wire393  &  wire30791 ) ;
 assign wire30794 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30795 = ( (~ ni13)  &  (~ ni14)  &  wire30794 ) ;
 assign wire30797 = ( (~ pi17)  &  pi21  &  pi22 ) ;
 assign wire30798 = ( wire5244 ) | ( wire257  &  wire916 ) ;
 assign wire30799 = ( wire5241 ) | ( wire295  &  wire916 ) ;
 assign wire30800 = ( (~ pi17)  &  pi25  &  pi16 ) ;
 assign wire30801 = ( (~ pi17)  &  pi25  &  (~ pi16) ) ;
 assign wire30802 = ( pi17  &  (~ pi19)  &  pi16  &  wire387 ) ;
 assign wire30803 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30804 = ( (~ pi20)  &  pi25  &  pi16  &  wire153 ) ;
 assign wire30805 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30806 = ( pi20  &  pi25  &  pi16  &  wire153 ) ;
 assign wire30807 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire387 ) ;
 assign wire30808 = ( wire5110 ) | ( wire5247 ) | ( wire5248 ) ;
 assign wire30813 = ( wire5240 ) | ( wire5243 ) | ( wire30798 ) | ( wire30799 ) ;
 assign wire30814 = ( wire5111 ) | ( wire5112 ) | ( wire5113 ) | ( wire5115 ) ;
 assign wire30815 = ( wire5116 ) | ( wire5119 ) | ( wire5120 ) | ( wire30808 ) ;
 assign wire30817 = ( wire30813 ) | ( wire30814 ) | ( wire30815 ) ;
 assign wire30819 = ( wire5109 ) | ( nv2290  &  wire812 ) ;
 assign wire30820 = ( wire5114 ) | ( wire30817 ) | ( nv2411  &  wire813 ) ;
 assign wire30823 = ( (~ pi15)  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30825 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30826 = ( (~ ni13)  &  (~ ni14)  &  wire30825 ) ;
 assign wire30827 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30828 = ( (~ ni13)  &  (~ ni14)  &  wire30827 ) ;
 assign wire30829 = ( pi15  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire30832 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire30833 = ( (~ pi16)  &  (~ pi15) ) ;
 assign wire30834 = ( pi20  &  pi25  &  wire153  &  wire30833 ) ;
 assign wire30835 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire30836 = ( wire30835  &  wire387 ) ;
 assign wire30837 = ( (~ pi16)  &  (~ pi15) ) ;
 assign wire30838 = ( (~ pi20)  &  pi25  &  wire153  &  wire30837 ) ;
 assign wire30839 = ( pi17  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire30840 = ( wire30839  &  wire387 ) ;
 assign wire30841 = ( (~ pi20)  &  pi25  &  wire258  &  wire153 ) ;
 assign wire30842 = ( pi25  &  (~ pi15)  &  wire158  &  wire152 ) ;
 assign wire30843 = ( (~ pi17)  &  pi25  &  pi16  &  (~ pi15) ) ;
 assign wire30844 = ( pi25  &  (~ pi15)  &  wire158  &  wire180 ) ;
 assign wire30845 = ( pi17  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire30846 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire30847 = ( pi25  &  (~ pi15)  &  wire180  &  wire154 ) ;
 assign wire30848 = ( pi20  &  pi25  &  wire258  &  wire153 ) ;
 assign wire30849 = ( pi25  &  (~ pi15)  &  wire152  &  wire154 ) ;
 assign wire30850 = ( (~ pi17)  &  pi25  &  pi16 ) ;
 assign wire30852 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30853 = ( pi17  &  (~ pi19)  &  pi16  &  wire387 ) ;
 assign wire30854 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire387 ) ;
 assign wire30855 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30857 = ( wire5152 ) | ( wire304  &  wire393 ) | ( wire393  &  wire5778 ) ;
 assign wire30858 = ( wire5243 ) | ( wire30798 ) | ( nv3377  &  wire311 ) ;
 assign wire30859 = ( wire694 ) | ( wire5151 ) | ( wire5240 ) | ( wire30799 ) ;
 assign wire30862 = ( wire30857 ) | ( wire30858 ) | ( nv3273  &  wire30852 ) ;
 assign wire30863 = ( wire5150 ) | ( wire30859 ) | ( nv3369  &  wire813 ) ;
 assign wire30865 = ( wire5148 ) | ( wire304  &  wire30854 ) | ( wire5829  &  wire30854 ) ;
 assign wire30866 = ( wire30862 ) | ( wire30863 ) | ( nv3311  &  wire812 ) ;
 assign wire30869 = ( wire916  &  wire30845 ) | ( wire5249  &  wire30845 ) | ( wire916  &  wire30846 ) | ( wire5249  &  wire30846 ) ;
 assign wire30873 = ( wire5140 ) | ( nv3202  &  wire30842 ) ;
 assign wire30875 = ( wire5128 ) | ( wire5139 ) | ( wire5144 ) | ( wire30869 ) ;
 assign wire30876 = ( wire5130 ) | ( wire5132 ) | ( wire30873 ) ;
 assign wire30877 = ( wire5142 ) | ( wire5143 ) | ( wire30875 ) ;
 assign wire30880 = ( wire5138 ) | ( wire304  &  wire30836 ) | ( wire5215  &  wire30836 ) ;
 assign wire30882 = ( wire5135 ) | ( wire30876 ) | ( wire30877 ) | ( wire30880 ) ;
 assign wire30883 = ( wire5131 ) | ( wire5134 ) | ( n_n9647  &  wire30832 ) ;
 assign wire30885 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30887 = ( wire228  &  wire1043  &  wire30885 ) ;
 assign wire30888 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30889 = ( (~ pi20)  &  wire153  &  wire30888 ) ;
 assign wire30890 = ( (~ pi25)  &  wire303  &  wire30889 ) ;
 assign wire30891 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30893 = ( wire228  &  wire181  &  wire30891 ) ;
 assign wire30894 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30895 = ( (~ pi25)  &  wire152  &  wire303  &  wire30894 ) ;
 assign wire30896 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30897 = ( (~ pi25)  &  wire178  &  wire303  &  wire30896 ) ;
 assign wire30898 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30899 = ( (~ pi25)  &  wire180  &  wire303  &  wire30898 ) ;
 assign wire30900 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30901 = ( (~ pi25)  &  wire179  &  wire303  &  wire30900 ) ;
 assign wire30902 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30903 = ( wire30902  &  wire1080 ) ;
 assign wire30904 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30905 = ( (~ pi25)  &  wire182  &  wire303  &  wire30904 ) ;
 assign wire30906 = ( (~ pi25)  &  (~ ni32)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire30907 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30909 = ( pi25 ) | ( (~ pi20)  &  n_n9302 ) ;
 assign wire30910 = ( pi20  &  n_n9294 ) | ( (~ pi20)  &  n_n9304 ) ;
 assign wire30912 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30913 = ( wire5457  &  wire30912 ) | ( wire30909  &  wire30912 ) | ( wire30910  &  wire30912 ) ;
 assign wire30914 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30915 = ( wire5457  &  wire30914 ) | ( wire30909  &  wire30914 ) | ( wire30910  &  wire30914 ) ;
 assign wire30916 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30917 = ( (~ pi20)  &  pi25  &  wire153  &  wire30916 ) ;
 assign wire30918 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30919 = ( pi17  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30920 = ( pi16  &  pi15  &  ni14 ) ;
 assign wire30921 = ( (~ pi17)  &  pi16  &  pi15  &  ni14 ) ;
 assign wire30922 = ( (~ pi25)  &  wire158  &  wire152  &  wire303 ) ;
 assign wire30923 = ( (~ pi25)  &  wire158  &  wire178  &  wire303 ) ;
 assign wire30924 = ( (~ pi25)  &  wire158  &  wire180  &  wire303 ) ;
 assign wire30925 = ( (~ pi25)  &  wire302  &  wire179  &  wire303 ) ;
 assign wire30927 = ( (~ pi25)  &  wire302  &  wire182  &  wire303 ) ;
 assign wire30928 = ( (~ pi25)  &  (~ wire150)  &  wire303  &  wire697 ) ;
 assign wire30929 = ( pi21  &  pi22  &  pi25  &  wire697 ) ;
 assign wire30930 = ( wire302  &  wire5457 ) | ( wire302  &  wire30909 ) | ( wire302  &  wire30910 ) ;
 assign wire30931 = ( wire158  &  wire5457 ) | ( wire158  &  wire30909 ) | ( wire158  &  wire30910 ) ;
 assign wire30933 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30935 = ( wire5315 ) | ( pi17  &  (~ pi16)  &  wire953 ) ;
 assign wire30936 = ( wire983 ) | ( wire5312 ) | ( wire572  &  wire697 ) ;
 assign wire30938 = ( wire30936 ) | ( wire325  &  nv2930  &  wire313 ) ;
 assign wire30940 = ( wire5300 ) | ( wire5304 ) | ( wire30935 ) | ( wire30938 ) ;
 assign wire30941 = ( nv2995  &  wire30923 ) | ( nv2963  &  wire30925 ) ;
 assign wire30944 = ( wire5302 ) | ( wire5311 ) | ( nv2946  &  wire30928 ) ;
 assign wire30947 = ( wire5305 ) | ( wire5307 ) | ( wire5308 ) ;
 assign wire30948 = ( wire5309 ) | ( wire30940 ) | ( wire30941 ) | ( wire30944 ) ;
 assign wire30949 = ( ni14  &  pi15 ) ;
 assign wire30950 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire30951 = ( (~ pi25)  &  (~ wire150)  &  wire303  &  wire30950 ) ;
 assign wire30952 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire30953 = ( pi21  &  pi22  &  pi25  &  wire30952 ) ;
 assign wire30954 = ( (~ pi25)  &  wire152  &  wire154  &  wire303 ) ;
 assign wire30955 = ( (~ pi25)  &  wire178  &  wire154  &  wire303 ) ;
 assign wire30956 = ( (~ pi25)  &  wire180  &  wire154  &  wire303 ) ;
 assign wire30957 = ( (~ pi25)  &  wire179  &  wire1061  &  wire303 ) ;
 assign wire30959 = ( (~ pi25)  &  wire182  &  wire1061  &  wire303 ) ;
 assign wire30960 = ( wire1061  &  wire5457 ) | ( wire1061  &  wire30909 ) | ( wire1061  &  wire30910 ) ;
 assign wire30962 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire30963 = ( wire154  &  wire5457 ) | ( wire154  &  wire30909 ) | ( wire154  &  wire30910 ) ;
 assign wire30964 = ( (~ pi20)  &  pi25  &  pi16  &  wire153 ) ;
 assign wire30966 = ( wire154  &  wire953 ) | ( wire572  &  wire30962 ) ;
 assign wire30967 = ( wire5353 ) | ( wire5354 ) | ( pi16  &  wire794 ) ;
 assign wire30968 = ( wire30966 ) | ( wire5598  &  wire30954 ) | ( wire30578  &  wire30954 ) ;
 assign wire30969 = ( wire30967 ) | ( nv2766  &  wire1024  &  wire313 ) ;
 assign wire30973 = ( wire5346 ) | ( wire30969 ) | ( nv2793  &  wire30953 ) ;
 assign wire30974 = ( wire5340 ) | ( wire5352 ) | ( wire30968 ) | ( wire30973 ) ;
 assign wire30976 = ( wire5344 ) | ( nv2807  &  wire30957 ) ;
 assign wire30977 = ( wire5347 ) | ( wire30974 ) | ( nv2857  &  wire30955 ) ;
 assign wire30980 = ( (~ pi25)  &  wire158  &  wire152  &  wire303 ) ;
 assign wire30981 = ( (~ pi25)  &  wire158  &  wire178  &  wire303 ) ;
 assign wire30982 = ( (~ pi25)  &  wire158  &  wire180  &  wire303 ) ;
 assign wire30983 = ( (~ pi25)  &  wire302  &  wire179  &  wire303 ) ;
 assign wire30984 = ( pi17  &  (~ pi16)  &  wire1080 ) ;
 assign wire30985 = ( (~ pi25)  &  wire302  &  wire182  &  wire303 ) ;
 assign wire30986 = ( (~ pi25)  &  (~ wire150)  &  wire303  &  wire697 ) ;
 assign wire30987 = ( pi21  &  pi22  &  pi25  &  wire697 ) ;
 assign wire30988 = ( wire302  &  wire5457 ) | ( wire302  &  wire30909 ) | ( wire302  &  wire30910 ) ;
 assign wire30989 = ( wire158  &  wire5457 ) | ( wire158  &  wire30909 ) | ( wire158  &  wire30910 ) ;
 assign wire30990 = ( (~ pi25)  &  wire325  &  wire303 ) ;
 assign wire30991 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire30993 = ( wire5446 ) | ( n_n10412  &  wire30990 ) | ( wire30538  &  wire30990 ) ;
 assign wire30994 = ( wire572  &  wire697 ) | ( wire158  &  wire953 ) ;
 assign wire30996 = ( wire983 ) | ( wire5443 ) | ( wire30993 ) | ( wire30994 ) ;
 assign wire30999 = ( wire5431 ) | ( wire5437 ) | ( wire5442 ) | ( wire30996 ) ;
 assign wire31001 = ( wire5435 ) | ( wire30999 ) | ( nv2627  &  wire30987 ) ;
 assign wire31002 = ( nv2694  &  wire30981 ) | ( nv2641  &  wire30983 ) ;
 assign wire31005 = ( wire5433 ) | ( wire5436 ) | ( wire31001 ) | ( wire31002 ) ;
 assign wire31007 = ( wire5264 ) | ( wire5254 ) ;
 assign wire31008 = ( wire5267 ) | ( wire228  &  wire572  &  wire30907 ) ;
 assign wire31009 = ( wire953  &  wire30919 ) | ( wire794  &  wire30920 ) ;
 assign wire31012 = ( wire5258 ) | ( wire31007 ) | ( wire31008 ) | ( wire31009 ) ;
 assign wire31014 = ( wire5252 ) | ( wire31012 ) | ( nv3060  &  wire30887 ) ;
 assign wire31015 = ( nv3109  &  wire30897 ) | ( nv3077  &  wire30901 ) ;
 assign wire31018 = ( wire31015 ) | ( wire5558  &  wire30905 ) | ( wire30584  &  wire30905 ) ;
 assign wire31019 = ( wire5253 ) | ( wire5256 ) | ( wire5263 ) | ( wire31014 ) ;
 assign wire31022 = ( wire5261 ) | ( wire5262 ) | ( wire31018 ) | ( wire31019 ) ;
 assign wire31023 = ( wire31022 ) | ( wire30947  &  wire30949 ) | ( wire30948  &  wire30949 ) ;
 assign wire31028 = ( wire5090 ) | ( wire5094 ) | ( wire5098 ) | ( wire5099 ) ;
 assign wire31032 = ( wire5092 ) | ( wire5095 ) | ( wire5097 ) | ( wire5103 ) ;
 assign wire31033 = ( wire5089 ) | ( wire5101 ) | ( wire5102 ) ;
 assign wire31034 = ( wire5091 ) | ( wire5096 ) | ( wire31028 ) ;
 assign wire31037 = ( wire31032 ) | ( wire31033 ) | ( wire852  &  wire30777 ) ;
 assign wire31038 = ( wire5088 ) | ( wire31034 ) | ( wire31037 ) ;
 assign wire31039 = ( wire31038 ) | ( wire263  &  wire933  &  wire30823 ) ;
 assign wire31040 = ( wire31039 ) | ( (~ ni11)  &  ni12  &  wire762 ) ;
 assign wire31041 = ( wire762  &  wire1303 ) | ( (~ wire631)  &  n_n11295 ) ;
 assign wire31042 = ( (~ ni2)  &  (~ ni3)  &  (~ ni10)  &  (~ wire265) ) ;
 assign wire31043 = ( (~ ni2)  &  (~ ni3)  &  (~ wire202)  &  wire330 ) ;
 assign wire31045 = ( pi15  &  (~ wire289)  &  wire1340  &  wire486 ) ;
 assign wire31047 = ( pi15  &  (~ wire289)  &  wire154  &  wire1128 ) ;
 assign wire31049 = ( pi15  &  (~ wire289)  &  wire1031  &  wire687 ) ;
 assign wire31050 = ( pi15  &  (~ wire289)  &  wire1031 ) ;
 assign wire31052 = ( pi15  &  (~ wire289)  &  (~ wire157)  &  wire30524 ) ;
 assign wire31055 = ( pi15  &  (~ wire289)  &  wire593  &  wire687 ) ;
 assign wire31056 = ( pi15  &  (~ wire289)  &  wire593 ) ;
 assign wire31058 = ( pi15  &  (~ wire289)  &  wire1340 ) ;
 assign wire31059 = ( pi15  &  (~ wire289)  &  wire1031 ) ;
 assign wire31060 = ( pi15  &  (~ wire289)  &  wire1031 ) ;
 assign wire31061 = ( pi17  &  pi16  &  pi15  &  (~ wire289) ) ;
 assign wire31062 = ( pi15  &  (~ wire289)  &  wire593 ) ;
 assign wire31063 = ( pi15  &  (~ wire289)  &  wire593 ) ;
 assign wire31064 = ( pi21  &  pi22  &  wire289 ) ;
 assign wire31065 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire31066 = ( (~ wire157)  &  wire213  &  wire1340  &  wire30524 ) ;
 assign wire31067 = ( (~ wire157)  &  wire152  &  wire154  &  wire30524 ) ;
 assign wire31068 = ( (~ wire157)  &  wire189  &  wire1031  &  wire30524 ) ;
 assign wire31069 = ( (~ wire157)  &  wire213  &  wire1031  &  wire30524 ) ;
 assign wire31071 = ( (~ wire157)  &  wire189  &  wire593  &  wire30524 ) ;
 assign wire31072 = ( (~ wire157)  &  wire593  &  wire213  &  wire30524 ) ;
 assign wire31074 = ( wire5540 ) | ( nv2766  &  wire31066 ) ;
 assign wire31077 = ( wire903 ) | ( wire5534 ) | ( wire5545 ) ;
 assign wire31079 = ( wire5541 ) | ( wire5542 ) | ( wire5543 ) | ( wire5544 ) ;
 assign wire31081 = ( wire5537 ) | ( wire31074 ) | ( wire31077 ) | ( wire31079 ) ;
 assign wire31082 = ( wire31081 ) | ( nv2807  &  wire31069 ) ;
 assign wire31085 = ( wire158  &  (~ wire157)  &  wire152  &  wire30524 ) ;
 assign wire31086 = ( (~ wire157)  &  wire189  &  wire698  &  wire30524 ) ;
 assign wire31087 = ( (~ wire157)  &  wire213  &  wire698  &  wire30524 ) ;
 assign wire31088 = ( (~ wire157)  &  wire189  &  wire456  &  wire30524 ) ;
 assign wire31089 = ( (~ wire157)  &  wire456  &  wire213  &  wire30524 ) ;
 assign wire31090 = ( (~ wire157)  &  wire213  &  wire344  &  wire30524 ) ;
 assign wire31092 = ( wire5620 ) | ( wire5670 ) | ( wire294  &  wire200 ) ;
 assign wire31093 = ( wire5623 ) | ( wire5622 ) ;
 assign wire31098 = ( wire5624 ) | ( wire5625 ) | ( wire5626 ) | ( wire5627 ) ;
 assign wire31099 = ( wire5615 ) | ( wire5621 ) | ( wire31092 ) | ( wire31093 ) ;
 assign wire31101 = ( wire31098 ) | ( wire31099 ) | ( nv2641  &  wire31087 ) ;
 assign wire31104 = ( wire158  &  (~ wire157)  &  wire152  &  wire30524 ) ;
 assign wire31105 = ( (~ wire157)  &  wire189  &  wire698  &  wire30524 ) ;
 assign wire31106 = ( (~ wire157)  &  wire213  &  wire698  &  wire30524 ) ;
 assign wire31107 = ( (~ wire157)  &  wire189  &  wire456  &  wire30524 ) ;
 assign wire31108 = ( (~ wire157)  &  wire456  &  wire213  &  wire30524 ) ;
 assign wire31109 = ( (~ wire157)  &  wire213  &  wire344  &  wire30524 ) ;
 assign wire31110 = ( ni34  &  (~ ni33)  &  wire294  &  (~ wire157) ) ;
 assign wire31112 = ( wire5663 ) | ( nv2930  &  wire31109 ) ;
 assign wire31113 = ( wire5665 ) | ( wire5664 ) ;
 assign wire31114 = ( wire5667 ) | ( wire5666 ) ;
 assign wire31115 = ( wire968 ) | ( wire5656 ) | ( wire5668 ) ;
 assign wire31118 = ( wire31112 ) | ( wire31113 ) | ( wire31114 ) | ( wire31115 ) ;
 assign wire31119 = ( nv2963  &  wire31106 ) | ( nv2995  &  wire31108 ) ;
 assign wire31121 = ( wire31118 ) | ( wire31119 ) | ( nv2946  &  wire31110 ) ;
 assign wire31122 = ( wire5657 ) | ( wire5711  &  wire31107 ) | ( wire30566  &  wire31107 ) ;
 assign wire31125 = ( wire5512 ) | ( wire5518 ) | ( wire5524 ) | ( wire5529 ) ;
 assign wire31130 = ( wire5521 ) | ( wire5522 ) | ( wire5523 ) | ( wire5525 ) ;
 assign wire31131 = ( wire5511 ) | ( wire5519 ) | ( wire5520 ) | ( wire31125 ) ;
 assign wire31132 = ( wire31130 ) | ( nv3060  &  wire763  &  wire31052 ) ;
 assign wire31136 = ( wire5514 ) | ( wire5517 ) | ( wire31131 ) | ( wire31132 ) ;
 assign wire31137 = ( wire5513 ) | ( wire5516 ) | ( wire31136 ) ;
 assign wire31139 = ( wire5528 ) | ( wire31137 ) | ( wire708  &  n_n9516 ) ;
 assign wire31140 = ( (~ ni2)  &  (~ ni3)  &  wire265 ) ;
 assign wire31141 = ( wire5010 ) | ( wire438  &  wire30402 ) ;
 assign wire31142 = ( wire438  &  wire30461 ) | ( wire1336  &  wire30521 ) ;
 assign wire31144 = ( wire5000 ) | ( wire31141 ) | ( wire31142 ) ;
 assign wire31145 = ( wire31144 ) | ( wire304  &  wire30393 ) | ( wire5778  &  wire30393 ) ;
 assign wire31147 = ( wire5002 ) | ( wire31145 ) | ( nv3280  &  wire30436 ) ;
 assign wire31148 = ( wire31147 ) | ( nv3273  &  wire325  &  wire30419 ) ;
 assign wire31149 = ( nv3311  &  wire30379 ) | ( nv3369  &  wire30408 ) ;
 assign wire31152 = ( wire4991 ) | ( wire4995 ) | ( wire31148 ) | ( wire31149 ) ;
 assign wire31155 = ( wire4997 ) | ( wire4999 ) | ( wire5003 ) | ( wire31152 ) ;
 assign wire31157 = ( wire5009 ) | ( wire31155 ) | ( n_n9650  &  wire30519 ) ;
 assign wire31159 = ( wire5006 ) | ( wire31157 ) | ( wire762  &  wire31043 ) ;
 assign wire31160 = ( (~ pi23)  &  (~ pi24)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire31161 = ( (~ ni9)  &  (~ ni7)  &  (~ ni8) ) | ( (~ ni10)  &  (~ ni7)  &  (~ ni8) ) | ( ni9  &  ni10  &  (~ ni7)  &  ni8 ) ;
 assign wire31162 = ( wire331  &  wire31160 ) | ( pi24  &  wire509  &  wire331 ) ;
 assign wire31163 = ( (~ pi25)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire31164 = ( (~ ni7)  &  ni10 ) ;
 assign wire31165 = ( (~ ni33)  &  ni10  &  ni29 ) ;
 assign wire31166 = ( wire31161  &  wire31163 ) | ( wire31162  &  wire31163 ) | ( (~ wire31161)  &  (~ wire31162)  &  wire31164 ) ;
 assign wire31167 = ( ni8  &  wire31161 ) | ( ni8  &  wire31162 ) | ( wire31161  &  wire31165 ) | ( wire31162  &  wire31165 ) ;
 assign wire31168 = ( (~ ni7)  &  ni10 ) ;
 assign wire31169 = ( wire4981 ) | ( (~ wire31166)  &  (~ wire31167)  &  wire31168 ) ;
 assign wire31170 = ( (~ ni33)  &  (~ ni32)  &  ni29 ) ;
 assign wire31171 = ( (~ ni31)  &  (~ ni30)  &  wire31170 ) ;
 assign wire31172 = ( ni39  &  (~ ni38)  &  (~ ni36)  &  nv3916 ) ;
 assign wire31173 = ( (~ ni43)  &  (~ ni42)  &  ni44 ) ;
 assign wire31176 = ( wire4886 ) | ( ni36  &  wire323 ) | ( ni35  &  wire323 ) ;
 assign wire31177 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31178 = ( ni40  &  wire31177 ) | ( ni37  &  wire31177 ) | ( (~ ni36)  &  wire31177 ) ;
 assign wire31179 = ( (~ ni36)  &  (~ wire4649)  &  wire31178 ) | ( wire255  &  (~ wire4649)  &  wire31178 ) ;
 assign wire31180 = ( (~ wire4889)  &  (~ wire4890)  &  (~ wire4891)  &  wire31179 ) ;
 assign wire31181 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31183 = ( (~ ni36)  &  wire31181 ) | ( ni40  &  (~ ni37)  &  wire31181 ) ;
 assign wire31184 = ( (~ ni36)  &  (~ wire4649)  &  wire31183 ) | ( wire255  &  (~ wire4649)  &  wire31183 ) ;
 assign wire31185 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31187 = ( (~ ni36)  &  wire31185 ) | ( ni40  &  (~ ni37)  &  wire31185 ) ;
 assign wire31188 = ( (~ ni36)  &  (~ wire4649)  &  wire31187 ) | ( wire255  &  (~ wire4649)  &  wire31187 ) ;
 assign wire31190 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31191 = ( ni40  &  ni36  &  ni35 ) | ( ni37  &  ni36  &  ni35 ) ;
 assign wire31192 = ( wire31191  &  wire31190 ) ;
 assign wire31193 = ( (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31194 = ( (~ ni36)  &  (~ wire4649)  &  wire31193 ) | ( wire255  &  (~ wire4649)  &  wire31193 ) ;
 assign wire31195 = ( (~ wire253)  &  (~ wire4892)  &  wire31194 ) | ( (~ nv3927)  &  (~ wire4892)  &  wire31194 ) ;
 assign wire31196 = ( (~ wire4889)  &  (~ wire4890)  &  (~ wire4891)  &  wire31195 ) ;
 assign wire31198 = ( ni35  &  (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31199 = ( (~ ni36)  &  (~ wire4649)  &  wire31198 ) | ( wire255  &  (~ wire4649)  &  wire31198 ) ;
 assign wire31200 = ( (~ wire253)  &  (~ wire4892)  &  wire31199 ) | ( (~ nv3927)  &  (~ wire4892)  &  wire31199 ) ;
 assign wire31202 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31203 = ( (~ ni36)  &  (~ wire4649)  &  wire31202 ) | ( wire255  &  (~ wire4649)  &  wire31202 ) ;
 assign wire31204 = ( (~ wire253)  &  (~ wire4892)  &  wire31203 ) | ( (~ nv3927)  &  (~ wire4892)  &  wire31203 ) ;
 assign wire31206 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31207 = ( ni40  &  wire31206 ) | ( ni37  &  wire31206 ) | ( (~ ni36)  &  wire31206 ) ;
 assign wire31208 = ( (~ ni36)  &  (~ wire4649)  &  wire31207 ) | ( wire255  &  (~ wire4649)  &  wire31207 ) ;
 assign wire31209 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31211 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4649)  &  wire31209 ) ;
 assign wire31212 = ( (~ wire4889)  &  (~ wire4890)  &  (~ wire4891)  &  wire31211 ) ;
 assign wire31213 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31214 = ( (~ ni37)  &  wire31213 ) | ( (~ ni36)  &  wire31213 ) ;
 assign wire31216 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4649)  &  wire31214 ) ;
 assign wire31218 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31220 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4649)  &  wire31218 ) ;
 assign wire31222 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31223 = ( ni36  &  ni35  &  wire31222 ) ;
 assign wire31227 = ( wire206  &  (~ nv3927)  &  (~ wire1189)  &  (~ n_n9157) ) ;
 assign wire31229 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31232 = ( (~ nv3927)  &  (~ wire1189)  &  (~ n_n9157)  &  wire31229 ) ;
 assign wire31233 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31236 = ( (~ nv3927)  &  (~ wire1189)  &  (~ n_n9157)  &  wire31233 ) ;
 assign wire31238 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31240 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4649)  &  wire31238 ) ;
 assign wire31241 = ( n_n6710 ) | ( (~ wire689)  &  (~ wire4649)  &  wire31192 ) ;
 assign wire31242 = ( wire31241 ) | ( (~ nv3927)  &  (~ wire1189)  &  wire31223 ) ;
 assign wire31244 = ( wire31242 ) | ( (~ n_n9157)  &  wire31208 ) | ( (~ n_n9157)  &  wire31240 ) ;
 assign wire31247 = ( wire31244 ) | ( (~ n_n8956)  &  wire31188 ) | ( (~ n_n8956)  &  wire31236 ) ;
 assign wire31249 = ( (~ wire4887)  &  (~ wire31176)  &  wire31184 ) | ( (~ wire4887)  &  (~ wire31176)  &  wire31196 ) ;
 assign wire31250 = ( (~ wire4887)  &  (~ wire31176)  &  wire31200 ) | ( (~ wire4887)  &  (~ wire31176)  &  wire31212 ) ;
 assign wire31252 = ( wire31247 ) | ( (~ wire4887)  &  (~ wire31176)  &  wire31232 ) ;
 assign wire31253 = ( wire4632 ) | ( wire4638 ) | ( wire4642 ) | ( wire31249 ) ;
 assign wire31254 = ( wire4641 ) | ( wire4644 ) | ( wire31250 ) ;
 assign wire31257 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire178 ) ;
 assign wire31258 = ( (~ ni43)  &  (~ ni42)  &  (~ ni44) ) ;
 assign wire31260 = ( (~ ni39)  &  (~ ni38)  &  (~ ni36)  &  nv3916 ) ;
 assign wire31262 = ( wire4896 ) | ( ni36  &  wire323 ) | ( ni35  &  wire323 ) ;
 assign wire31263 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31264 = ( ni40  &  wire31263 ) | ( ni37  &  wire31263 ) | ( (~ ni36)  &  wire31263 ) ;
 assign wire31265 = ( (~ ni36)  &  (~ wire4649)  &  wire31264 ) | ( wire255  &  (~ wire4649)  &  wire31264 ) ;
 assign wire31266 = ( (~ wire4899)  &  (~ wire4900)  &  (~ wire4901)  &  wire31265 ) ;
 assign wire31267 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31269 = ( (~ ni36)  &  wire31267 ) | ( ni40  &  (~ ni37)  &  wire31267 ) ;
 assign wire31270 = ( (~ ni36)  &  (~ wire4649)  &  wire31269 ) | ( wire255  &  (~ wire4649)  &  wire31269 ) ;
 assign wire31271 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31273 = ( (~ ni36)  &  wire31271 ) | ( ni40  &  (~ ni37)  &  wire31271 ) ;
 assign wire31274 = ( (~ ni36)  &  (~ wire4649)  &  wire31273 ) | ( wire255  &  (~ wire4649)  &  wire31273 ) ;
 assign wire31276 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31277 = ( ni40  &  ni36  &  ni35 ) | ( ni37  &  ni36  &  ni35 ) ;
 assign wire31278 = ( wire31277  &  wire31276 ) ;
 assign wire31279 = ( (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31280 = ( (~ ni36)  &  (~ wire4649)  &  wire31279 ) | ( wire255  &  (~ wire4649)  &  wire31279 ) ;
 assign wire31281 = ( (~ wire253)  &  (~ wire4904)  &  wire31280 ) | ( (~ nv3943)  &  (~ wire4904)  &  wire31280 ) ;
 assign wire31282 = ( (~ wire4899)  &  (~ wire4900)  &  (~ wire4901)  &  wire31281 ) ;
 assign wire31284 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31285 = ( (~ ni36)  &  (~ wire4649)  &  wire31284 ) | ( wire255  &  (~ wire4649)  &  wire31284 ) ;
 assign wire31286 = ( (~ wire253)  &  (~ wire4904)  &  wire31285 ) | ( (~ nv3943)  &  (~ wire4904)  &  wire31285 ) ;
 assign wire31288 = ( ni35  &  (~ ni31)  &  (~ ni30)  &  (~ wire347) ) ;
 assign wire31289 = ( (~ ni36)  &  (~ wire4649)  &  wire31288 ) | ( wire255  &  (~ wire4649)  &  wire31288 ) ;
 assign wire31290 = ( (~ wire253)  &  (~ wire4904)  &  wire31289 ) | ( (~ nv3943)  &  (~ wire4904)  &  wire31289 ) ;
 assign wire31292 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31293 = ( ni40  &  wire31292 ) | ( ni37  &  wire31292 ) | ( (~ ni36)  &  wire31292 ) ;
 assign wire31294 = ( (~ ni36)  &  (~ wire4649)  &  wire31293 ) | ( wire255  &  (~ wire4649)  &  wire31293 ) ;
 assign wire31295 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31297 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4649)  &  wire31295 ) ;
 assign wire31298 = ( (~ wire4899)  &  (~ wire4900)  &  (~ wire4901)  &  wire31297 ) ;
 assign wire31300 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31302 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4649)  &  wire31300 ) ;
 assign wire31303 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31304 = ( (~ ni37)  &  wire31303 ) | ( (~ ni36)  &  wire31303 ) ;
 assign wire31306 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4649)  &  wire31304 ) ;
 assign wire31308 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31309 = ( ni36  &  ni35  &  wire31308 ) ;
 assign wire31313 = ( wire206  &  (~ nv3943)  &  (~ n_n9141)  &  (~ wire1189) ) ;
 assign wire31315 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31318 = ( (~ nv3943)  &  (~ n_n9141)  &  (~ wire1189)  &  wire31315 ) ;
 assign wire31319 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31322 = ( (~ nv3943)  &  (~ n_n9141)  &  (~ wire1189)  &  wire31319 ) ;
 assign wire31324 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31326 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4649)  &  wire31324 ) ;
 assign wire31327 = ( n_n6710 ) | ( (~ wire689)  &  (~ wire4649)  &  wire31278 ) ;
 assign wire31328 = ( wire31327 ) | ( (~ nv3943)  &  (~ wire1189)  &  wire31309 ) ;
 assign wire31330 = ( wire31328 ) | ( (~ n_n9141)  &  wire31294 ) | ( (~ n_n9141)  &  wire31326 ) ;
 assign wire31333 = ( wire31330 ) | ( (~ n_n8948)  &  wire31270 ) | ( (~ n_n8948)  &  wire31318 ) ;
 assign wire31335 = ( (~ wire4897)  &  (~ wire31262)  &  wire31274 ) | ( (~ wire4897)  &  (~ wire31262)  &  wire31282 ) ;
 assign wire31336 = ( (~ wire4897)  &  (~ wire31262)  &  wire31290 ) | ( (~ wire4897)  &  (~ wire31262)  &  wire31298 ) ;
 assign wire31338 = ( wire31333 ) | ( (~ wire4897)  &  (~ wire31262)  &  wire31322 ) ;
 assign wire31339 = ( wire4615 ) | ( wire4620 ) | ( wire4624 ) | ( wire31335 ) ;
 assign wire31340 = ( wire4625 ) | ( wire4627 ) | ( wire31336 ) ;
 assign wire31343 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire180 ) ;
 assign wire31345 = ( wire206  &  wire4685 ) | ( (~ ni37)  &  ni36  &  wire206 ) ;
 assign wire31346 = ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31347 = ( wire928 ) | ( (~ nv3961)  &  wire31345 ) ;
 assign wire31348 = ( (~ pi15)  &  (~ pi16) ) ;
 assign wire31350 = ( (~ pi15)  &  (~ pi16) ) ;
 assign wire31352 = ( wire4843 ) | ( ni36  &  wire323 ) | ( ni35  &  wire323 ) ;
 assign wire31353 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31355 = ( (~ wire347)  &  (~ wire1185)  &  wire31353 ) ;
 assign wire31356 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31355 ) ;
 assign wire31357 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31358 = ( (~ ni36) ) | ( ni40  &  (~ ni37) ) ;
 assign wire31360 = ( (~ wire1185)  &  wire31357  &  wire31358 ) ;
 assign wire31361 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31362 = ( (~ ni36) ) | ( ni40  &  (~ ni37) ) ;
 assign wire31364 = ( (~ wire1185)  &  wire31361  &  wire31362 ) ;
 assign wire31366 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31367 = ( ni40  &  ni36  &  ni35 ) | ( ni37  &  ni36  &  ni35 ) ;
 assign wire31368 = ( wire31367  &  wire31366 ) ;
 assign wire31370 = ( (~ ni31)  &  (~ ni30)  &  (~ wire347)  &  (~ wire1185) ) ;
 assign wire31371 = ( (~ wire253)  &  (~ wire4851)  &  wire31370 ) | ( (~ nv4058)  &  (~ wire4851)  &  wire31370 ) ;
 assign wire31372 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31371 ) ;
 assign wire31373 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31375 = ( (~ wire347)  &  (~ wire1185)  &  wire31373 ) ;
 assign wire31376 = ( (~ wire253)  &  (~ wire4851)  &  wire31375 ) | ( (~ nv4058)  &  (~ wire4851)  &  wire31375 ) ;
 assign wire31377 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31379 = ( (~ wire347)  &  (~ wire1185)  &  wire31377 ) ;
 assign wire31380 = ( (~ wire253)  &  (~ wire4851)  &  wire31379 ) | ( (~ nv4058)  &  (~ wire4851)  &  wire31379 ) ;
 assign wire31382 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31384 = ( (~ wire347)  &  (~ wire1185)  &  wire31382 ) ;
 assign wire31385 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31387 = ( (~ nv4058)  &  (~ wire1185)  &  wire31385 ) ;
 assign wire31388 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31387 ) ;
 assign wire31390 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31392 = ( (~ nv4058)  &  (~ wire1185)  &  wire31390 ) ;
 assign wire31393 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31396 = ( (~ wire270)  &  (~ nv4058)  &  (~ wire1185)  &  wire31393 ) ;
 assign wire31398 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31399 = ( ni36  &  ni35  &  wire31398 ) ;
 assign wire31401 = ( (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31403 = ( (~ wire254)  &  (~ nv4058)  &  wire31401 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31401 ) ;
 assign wire31404 = ( (~ wire4846)  &  (~ wire4847)  &  (~ wire4848)  &  wire31403 ) ;
 assign wire31406 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31408 = ( (~ wire254)  &  (~ nv4058)  &  wire31406 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31406 ) ;
 assign wire31410 = ( ni35  &  (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31412 = ( (~ wire254)  &  (~ nv4058)  &  wire31410 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31410 ) ;
 assign wire31414 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31415 = ( (~ wire1185)  &  wire31414 ) ;
 assign wire31417 = ( ni32  &  (~ ni30) ) | ( (~ wire1185)  &  wire31368 ) ;
 assign wire31418 = ( wire31417 ) | ( (~ nv4058)  &  (~ wire1185)  &  wire31399 ) ;
 assign wire31420 = ( wire4697 ) | ( wire4705 ) | ( wire31418 ) ;
 assign wire31425 = ( (~ wire4844)  &  (~ wire31352)  &  wire31364 ) | ( (~ wire4844)  &  (~ wire31352)  &  wire31372 ) ;
 assign wire31426 = ( (~ wire4844)  &  (~ wire31352)  &  wire31380 ) | ( (~ wire4844)  &  (~ wire31352)  &  wire31388 ) ;
 assign wire31427 = ( (~ wire4844)  &  (~ wire31352)  &  wire31396 ) | ( (~ wire4844)  &  (~ wire31352)  &  wire31404 ) ;
 assign wire31428 = ( wire4691 ) | ( wire4703 ) | ( wire4704 ) | ( wire31420 ) ;
 assign wire31429 = ( wire4690 ) | ( wire4695 ) | ( wire4699 ) | ( wire31425 ) ;
 assign wire31430 = ( wire31427 ) | ( wire31426 ) ;
 assign wire31434 = ( wire4833 ) | ( ni36  &  wire323 ) | ( ni35  &  wire323 ) ;
 assign wire31435 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31437 = ( (~ wire347)  &  (~ wire1185)  &  wire31435 ) ;
 assign wire31438 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31437 ) ;
 assign wire31439 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31440 = ( (~ ni36) ) | ( ni40  &  (~ ni37) ) ;
 assign wire31442 = ( (~ wire1185)  &  wire31439  &  wire31440 ) ;
 assign wire31443 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31444 = ( (~ ni36) ) | ( ni40  &  (~ ni37) ) ;
 assign wire31446 = ( (~ wire1185)  &  wire31443  &  wire31444 ) ;
 assign wire31448 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31449 = ( ni40  &  ni36  &  ni35 ) | ( ni37  &  ni36  &  ni35 ) ;
 assign wire31450 = ( wire31449  &  wire31448 ) ;
 assign wire31452 = ( (~ ni31)  &  (~ ni30)  &  (~ wire347)  &  (~ wire1185) ) ;
 assign wire31453 = ( (~ wire253)  &  (~ wire4839)  &  wire31452 ) | ( (~ nv4045)  &  (~ wire4839)  &  wire31452 ) ;
 assign wire31454 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31453 ) ;
 assign wire31455 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31457 = ( (~ wire347)  &  (~ wire1185)  &  wire31455 ) ;
 assign wire31458 = ( (~ wire253)  &  (~ wire4839)  &  wire31457 ) | ( (~ nv4045)  &  (~ wire4839)  &  wire31457 ) ;
 assign wire31459 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31461 = ( (~ wire347)  &  (~ wire1185)  &  wire31459 ) ;
 assign wire31462 = ( (~ wire253)  &  (~ wire4839)  &  wire31461 ) | ( (~ nv4045)  &  (~ wire4839)  &  wire31461 ) ;
 assign wire31464 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31466 = ( (~ wire347)  &  (~ wire1185)  &  wire31464 ) ;
 assign wire31467 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31469 = ( (~ nv4045)  &  (~ wire1185)  &  wire31467 ) ;
 assign wire31470 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31469 ) ;
 assign wire31471 = ( ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31474 = ( (~ wire270)  &  (~ nv4045)  &  (~ wire1185)  &  wire31471 ) ;
 assign wire31476 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31478 = ( (~ nv4045)  &  (~ wire1185)  &  wire31476 ) ;
 assign wire31480 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31481 = ( ni36  &  ni35  &  wire31480 ) ;
 assign wire31483 = ( (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31485 = ( (~ wire254)  &  (~ nv4045)  &  wire31483 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31483 ) ;
 assign wire31486 = ( (~ wire4836)  &  (~ wire4837)  &  (~ wire4838)  &  wire31485 ) ;
 assign wire31488 = ( ni35  &  (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31490 = ( (~ wire254)  &  (~ nv4045)  &  wire31488 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31488 ) ;
 assign wire31492 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire1185) ) ;
 assign wire31494 = ( (~ wire254)  &  (~ nv4045)  &  wire31492 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31492 ) ;
 assign wire31496 = ( ni36  &  ni35  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31497 = ( (~ wire1185)  &  wire31496 ) ;
 assign wire31499 = ( ni32  &  (~ ni30) ) | ( (~ wire1185)  &  wire31450 ) ;
 assign wire31500 = ( wire31499 ) | ( (~ nv4045)  &  (~ wire1185)  &  wire31481 ) ;
 assign wire31502 = ( wire4714 ) | ( wire4722 ) | ( wire31500 ) ;
 assign wire31507 = ( (~ wire4834)  &  (~ wire31434)  &  wire31442 ) | ( (~ wire4834)  &  (~ wire31434)  &  wire31454 ) ;
 assign wire31508 = ( (~ wire4834)  &  (~ wire31434)  &  wire31458 ) | ( (~ wire4834)  &  (~ wire31434)  &  wire31470 ) ;
 assign wire31509 = ( (~ wire4834)  &  (~ wire31434)  &  wire31474 ) | ( (~ wire4834)  &  (~ wire31434)  &  wire31486 ) ;
 assign wire31510 = ( wire4709 ) | ( wire4720 ) | ( wire4721 ) | ( wire31502 ) ;
 assign wire31511 = ( wire4707 ) | ( wire4713 ) | ( wire4717 ) | ( wire31507 ) ;
 assign wire31512 = ( wire31509 ) | ( wire31508 ) ;
 assign wire31516 = ( wire4952 ) | ( ni36  &  wire323 ) | ( (~ ni35)  &  wire323 ) ;
 assign wire31517 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31518 = ( (~ ni40)  &  wire31517 ) | ( ni37  &  wire31517 ) | ( (~ ni36)  &  wire31517 ) ;
 assign wire31519 = ( (~ ni36)  &  (~ wire4950)  &  wire31518 ) | ( wire255  &  (~ wire4950)  &  wire31518 ) ;
 assign wire31520 = ( (~ wire4957)  &  (~ wire4958)  &  (~ wire4959)  &  wire31519 ) ;
 assign wire31521 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31523 = ( (~ ni36)  &  wire31521 ) | ( (~ ni40)  &  (~ ni37)  &  wire31521 ) ;
 assign wire31524 = ( (~ ni36)  &  (~ wire4950)  &  wire31523 ) | ( wire255  &  (~ wire4950)  &  wire31523 ) ;
 assign wire31525 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31527 = ( (~ ni36)  &  wire31525 ) | ( (~ ni40)  &  (~ ni37)  &  wire31525 ) ;
 assign wire31528 = ( (~ ni36)  &  (~ wire4950)  &  wire31527 ) | ( wire255  &  (~ wire4950)  &  wire31527 ) ;
 assign wire31530 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31531 = ( (~ ni40)  &  ni36  &  (~ ni35) ) | ( ni37  &  ni36  &  (~ ni35) ) ;
 assign wire31532 = ( wire31531  &  wire31530 ) ;
 assign wire31533 = ( (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31534 = ( (~ ni36)  &  (~ wire4950)  &  wire31533 ) | ( wire255  &  (~ wire4950)  &  wire31533 ) ;
 assign wire31535 = ( (~ wire254)  &  (~ wire4967)  &  wire31534 ) | ( (~ nv3927)  &  (~ wire4967)  &  wire31534 ) ;
 assign wire31536 = ( (~ wire4957)  &  (~ wire4958)  &  (~ wire4959)  &  wire31535 ) ;
 assign wire31538 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31539 = ( (~ ni36)  &  (~ wire4950)  &  wire31538 ) | ( wire255  &  (~ wire4950)  &  wire31538 ) ;
 assign wire31540 = ( (~ wire254)  &  (~ wire4967)  &  wire31539 ) | ( (~ nv3927)  &  (~ wire4967)  &  wire31539 ) ;
 assign wire31542 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31543 = ( (~ ni36)  &  (~ wire4950)  &  wire31542 ) | ( wire255  &  (~ wire4950)  &  wire31542 ) ;
 assign wire31544 = ( (~ wire254)  &  (~ wire4967)  &  wire31543 ) | ( (~ nv3927)  &  (~ wire4967)  &  wire31543 ) ;
 assign wire31546 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31547 = ( (~ ni40)  &  wire31546 ) | ( ni37  &  wire31546 ) | ( (~ ni36)  &  wire31546 ) ;
 assign wire31548 = ( (~ ni36)  &  (~ wire4950)  &  wire31547 ) | ( wire255  &  (~ wire4950)  &  wire31547 ) ;
 assign wire31549 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31551 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4950)  &  wire31549 ) ;
 assign wire31552 = ( (~ wire4957)  &  (~ wire4958)  &  (~ wire4959)  &  wire31551 ) ;
 assign wire31554 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31556 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4950)  &  wire31554 ) ;
 assign wire31557 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31558 = ( (~ ni37)  &  wire31557 ) | ( (~ ni36)  &  wire31557 ) ;
 assign wire31560 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4950)  &  wire31558 ) ;
 assign wire31562 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31563 = ( ni36  &  (~ ni35)  &  wire31562 ) ;
 assign wire31567 = ( wire206  &  (~ n_n9194)  &  (~ nv3927)  &  (~ wire1180) ) ;
 assign wire31569 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31572 = ( (~ n_n9194)  &  (~ nv3927)  &  (~ wire1180)  &  wire31569 ) ;
 assign wire31573 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31576 = ( (~ n_n9194)  &  (~ nv3927)  &  (~ wire1180)  &  wire31573 ) ;
 assign wire31578 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31580 = ( (~ nv3927)  &  (~ wire689)  &  (~ wire4950)  &  wire31578 ) ;
 assign wire31581 = ( n_n6710 ) | ( (~ wire689)  &  (~ wire4950)  &  wire31532 ) ;
 assign wire31582 = ( wire31581 ) | ( (~ nv3927)  &  (~ wire1180)  &  wire31563 ) ;
 assign wire31584 = ( wire31582 ) | ( (~ n_n9194)  &  wire31548 ) | ( (~ n_n9194)  &  wire31580 ) ;
 assign wire31587 = ( wire31584 ) | ( (~ n_n8976)  &  wire31524 ) | ( (~ n_n8976)  &  wire31572 ) ;
 assign wire31589 = ( (~ wire4953)  &  (~ wire31516)  &  wire31528 ) | ( (~ wire4953)  &  (~ wire31516)  &  wire31536 ) ;
 assign wire31590 = ( (~ wire4953)  &  (~ wire31516)  &  wire31544 ) | ( (~ wire4953)  &  (~ wire31516)  &  wire31552 ) ;
 assign wire31592 = ( wire31587 ) | ( (~ wire4953)  &  (~ wire31516)  &  wire31576 ) ;
 assign wire31593 = ( wire4933 ) | ( wire4938 ) | ( wire4942 ) | ( wire31589 ) ;
 assign wire31594 = ( wire4943 ) | ( wire4945 ) | ( wire31590 ) ;
 assign wire31596 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire31598 = ( wire4792 ) | ( ni36  &  wire323 ) | ( (~ ni35)  &  wire323 ) ;
 assign wire31599 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31601 = ( (~ wire346)  &  (~ wire1182)  &  wire31599 ) ;
 assign wire31602 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31601 ) ;
 assign wire31603 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31604 = ( (~ ni36) ) | ( (~ ni40)  &  (~ ni37) ) ;
 assign wire31606 = ( (~ wire1182)  &  wire31603  &  wire31604 ) ;
 assign wire31607 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31608 = ( (~ ni36) ) | ( (~ ni40)  &  (~ ni37) ) ;
 assign wire31610 = ( (~ wire1182)  &  wire31607  &  wire31608 ) ;
 assign wire31612 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31613 = ( (~ ni40)  &  ni36  &  (~ ni35) ) | ( ni37  &  ni36  &  (~ ni35) ) ;
 assign wire31614 = ( wire31613  &  wire31612 ) ;
 assign wire31616 = ( (~ ni31)  &  (~ ni30)  &  (~ wire346)  &  (~ wire1182) ) ;
 assign wire31617 = ( (~ wire254)  &  (~ wire4799)  &  wire31616 ) | ( (~ nv4058)  &  (~ wire4799)  &  wire31616 ) ;
 assign wire31618 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31617 ) ;
 assign wire31619 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31621 = ( (~ wire346)  &  (~ wire1182)  &  wire31619 ) ;
 assign wire31622 = ( (~ wire254)  &  (~ wire4799)  &  wire31621 ) | ( (~ nv4058)  &  (~ wire4799)  &  wire31621 ) ;
 assign wire31623 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31625 = ( (~ wire346)  &  (~ wire1182)  &  wire31623 ) ;
 assign wire31626 = ( (~ wire254)  &  (~ wire4799)  &  wire31625 ) | ( (~ nv4058)  &  (~ wire4799)  &  wire31625 ) ;
 assign wire31628 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31630 = ( (~ wire346)  &  (~ wire1182)  &  wire31628 ) ;
 assign wire31631 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31633 = ( (~ nv4058)  &  (~ wire1182)  &  wire31631 ) ;
 assign wire31634 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31633 ) ;
 assign wire31635 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31638 = ( (~ wire270)  &  (~ nv4058)  &  (~ wire1182)  &  wire31635 ) ;
 assign wire31640 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31642 = ( (~ nv4058)  &  (~ wire1182)  &  wire31640 ) ;
 assign wire31644 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31645 = ( ni36  &  (~ ni35)  &  wire31644 ) ;
 assign wire31647 = ( (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31649 = ( (~ wire253)  &  (~ nv4058)  &  wire31647 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31647 ) ;
 assign wire31650 = ( (~ wire4795)  &  (~ wire4796)  &  (~ wire4797)  &  wire31649 ) ;
 assign wire31652 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31654 = ( (~ wire253)  &  (~ nv4058)  &  wire31652 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31652 ) ;
 assign wire31656 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31658 = ( (~ wire253)  &  (~ nv4058)  &  wire31656 ) | ( (~ nv3918)  &  (~ nv4058)  &  wire31656 ) ;
 assign wire31660 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31661 = ( (~ wire1182)  &  wire31660 ) ;
 assign wire31663 = ( ni32  &  (~ ni30) ) | ( (~ wire1182)  &  wire31614 ) ;
 assign wire31664 = ( wire31663 ) | ( (~ nv4058)  &  (~ wire1182)  &  wire31645 ) ;
 assign wire31666 = ( wire4668 ) | ( wire4676 ) | ( wire31664 ) ;
 assign wire31671 = ( (~ wire4793)  &  (~ wire31598)  &  wire31606 ) | ( (~ wire4793)  &  (~ wire31598)  &  wire31618 ) ;
 assign wire31672 = ( (~ wire4793)  &  (~ wire31598)  &  wire31622 ) | ( (~ wire4793)  &  (~ wire31598)  &  wire31634 ) ;
 assign wire31673 = ( (~ wire4793)  &  (~ wire31598)  &  wire31638 ) | ( (~ wire4793)  &  (~ wire31598)  &  wire31650 ) ;
 assign wire31674 = ( wire4663 ) | ( wire4674 ) | ( wire4675 ) | ( wire31666 ) ;
 assign wire31675 = ( wire4661 ) | ( wire4667 ) | ( wire4671 ) | ( wire31671 ) ;
 assign wire31676 = ( wire31673 ) | ( wire31672 ) ;
 assign wire31680 = ( wire4921 ) | ( ni36  &  wire323 ) | ( (~ ni35)  &  wire323 ) ;
 assign wire31681 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31683 = ( (~ wire346)  &  (~ wire1182)  &  wire31681 ) ;
 assign wire31684 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31683 ) ;
 assign wire31685 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31686 = ( (~ ni36) ) | ( (~ ni40)  &  (~ ni37) ) ;
 assign wire31688 = ( (~ wire1182)  &  wire31685  &  wire31686 ) ;
 assign wire31689 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31690 = ( (~ ni36) ) | ( (~ ni40)  &  (~ ni37) ) ;
 assign wire31692 = ( (~ wire1182)  &  wire31689  &  wire31690 ) ;
 assign wire31694 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31695 = ( (~ ni40)  &  ni36  &  (~ ni35) ) | ( ni37  &  ni36  &  (~ ni35) ) ;
 assign wire31696 = ( wire31695  &  wire31694 ) ;
 assign wire31698 = ( (~ ni31)  &  (~ ni30)  &  (~ wire346)  &  (~ wire1182) ) ;
 assign wire31699 = ( (~ wire254)  &  (~ wire4930)  &  wire31698 ) | ( (~ nv4045)  &  (~ wire4930)  &  wire31698 ) ;
 assign wire31700 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31699 ) ;
 assign wire31701 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31703 = ( (~ wire346)  &  (~ wire1182)  &  wire31701 ) ;
 assign wire31704 = ( (~ wire254)  &  (~ wire4930)  &  wire31703 ) | ( (~ nv4045)  &  (~ wire4930)  &  wire31703 ) ;
 assign wire31705 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31707 = ( (~ wire346)  &  (~ wire1182)  &  wire31705 ) ;
 assign wire31708 = ( (~ wire254)  &  (~ wire4930)  &  wire31707 ) | ( (~ nv4045)  &  (~ wire4930)  &  wire31707 ) ;
 assign wire31710 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31712 = ( (~ wire346)  &  (~ wire1182)  &  wire31710 ) ;
 assign wire31713 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31715 = ( (~ nv4045)  &  (~ wire1182)  &  wire31713 ) ;
 assign wire31716 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31715 ) ;
 assign wire31718 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31720 = ( (~ nv4045)  &  (~ wire1182)  &  wire31718 ) ;
 assign wire31721 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31724 = ( (~ wire270)  &  (~ nv4045)  &  (~ wire1182)  &  wire31721 ) ;
 assign wire31726 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31727 = ( ni36  &  (~ ni35)  &  wire31726 ) ;
 assign wire31729 = ( (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31731 = ( (~ wire253)  &  (~ nv4045)  &  wire31729 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31729 ) ;
 assign wire31732 = ( (~ wire4924)  &  (~ wire4925)  &  (~ wire4926)  &  wire31731 ) ;
 assign wire31734 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31736 = ( (~ wire253)  &  (~ nv4045)  &  wire31734 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31734 ) ;
 assign wire31738 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30)  &  (~ wire1182) ) ;
 assign wire31740 = ( (~ wire253)  &  (~ nv4045)  &  wire31738 ) | ( (~ nv3918)  &  (~ nv4045)  &  wire31738 ) ;
 assign wire31742 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31743 = ( (~ wire1182)  &  wire31742 ) ;
 assign wire31745 = ( ni32  &  (~ ni30) ) | ( (~ wire1182)  &  wire31696 ) ;
 assign wire31746 = ( wire31745 ) | ( (~ nv4045)  &  (~ wire1182)  &  wire31727 ) ;
 assign wire31748 = ( wire4745 ) | ( wire4753 ) | ( wire31746 ) ;
 assign wire31753 = ( (~ wire4922)  &  (~ wire31680)  &  wire31692 ) | ( (~ wire4922)  &  (~ wire31680)  &  wire31700 ) ;
 assign wire31754 = ( (~ wire4922)  &  (~ wire31680)  &  wire31708 ) | ( (~ wire4922)  &  (~ wire31680)  &  wire31716 ) ;
 assign wire31755 = ( (~ wire4922)  &  (~ wire31680)  &  wire31724 ) | ( (~ wire4922)  &  (~ wire31680)  &  wire31732 ) ;
 assign wire31756 = ( wire4739 ) | ( wire4751 ) | ( wire4752 ) | ( wire31748 ) ;
 assign wire31757 = ( wire4738 ) | ( wire4743 ) | ( wire4747 ) | ( wire31753 ) ;
 assign wire31758 = ( wire31755 ) | ( wire31754 ) ;
 assign wire31762 = ( wire4861 ) | ( ni36  &  wire323 ) | ( (~ ni35)  &  wire323 ) ;
 assign wire31763 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31764 = ( (~ ni40)  &  wire31763 ) | ( ni37  &  wire31763 ) | ( (~ ni36)  &  wire31763 ) ;
 assign wire31765 = ( (~ ni36)  &  (~ wire4950)  &  wire31764 ) | ( wire255  &  (~ wire4950)  &  wire31764 ) ;
 assign wire31766 = ( (~ wire4864)  &  (~ wire4865)  &  (~ wire4866)  &  wire31765 ) ;
 assign wire31767 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31769 = ( (~ ni36)  &  wire31767 ) | ( (~ ni40)  &  (~ ni37)  &  wire31767 ) ;
 assign wire31770 = ( (~ ni36)  &  (~ wire4950)  &  wire31769 ) | ( wire255  &  (~ wire4950)  &  wire31769 ) ;
 assign wire31771 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31773 = ( (~ ni36)  &  wire31771 ) | ( (~ ni40)  &  (~ ni37)  &  wire31771 ) ;
 assign wire31774 = ( (~ ni36)  &  (~ wire4950)  &  wire31773 ) | ( wire255  &  (~ wire4950)  &  wire31773 ) ;
 assign wire31776 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31777 = ( (~ ni40)  &  ni36  &  (~ ni35) ) | ( ni37  &  ni36  &  (~ ni35) ) ;
 assign wire31778 = ( wire31777  &  wire31776 ) ;
 assign wire31779 = ( (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31780 = ( (~ ni36)  &  (~ wire4950)  &  wire31779 ) | ( wire255  &  (~ wire4950)  &  wire31779 ) ;
 assign wire31781 = ( (~ wire254)  &  (~ wire4868)  &  wire31780 ) | ( (~ nv3943)  &  (~ wire4868)  &  wire31780 ) ;
 assign wire31782 = ( (~ wire4864)  &  (~ wire4865)  &  (~ wire4866)  &  wire31781 ) ;
 assign wire31784 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31785 = ( (~ ni36)  &  (~ wire4950)  &  wire31784 ) | ( wire255  &  (~ wire4950)  &  wire31784 ) ;
 assign wire31786 = ( (~ wire254)  &  (~ wire4868)  &  wire31785 ) | ( (~ nv3943)  &  (~ wire4868)  &  wire31785 ) ;
 assign wire31788 = ( ni36  &  (~ ni31)  &  (~ ni30)  &  (~ wire346) ) ;
 assign wire31789 = ( (~ ni36)  &  (~ wire4950)  &  wire31788 ) | ( wire255  &  (~ wire4950)  &  wire31788 ) ;
 assign wire31790 = ( (~ wire254)  &  (~ wire4868)  &  wire31789 ) | ( (~ nv3943)  &  (~ wire4868)  &  wire31789 ) ;
 assign wire31792 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31793 = ( (~ ni40)  &  wire31792 ) | ( ni37  &  wire31792 ) | ( (~ ni36)  &  wire31792 ) ;
 assign wire31794 = ( (~ ni36)  &  (~ wire4950)  &  wire31793 ) | ( wire255  &  (~ wire4950)  &  wire31793 ) ;
 assign wire31795 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31797 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4950)  &  wire31795 ) ;
 assign wire31798 = ( (~ wire4864)  &  (~ wire4865)  &  (~ wire4866)  &  wire31797 ) ;
 assign wire31799 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31800 = ( (~ ni37)  &  wire31799 ) | ( (~ ni36)  &  wire31799 ) ;
 assign wire31802 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4950)  &  wire31800 ) ;
 assign wire31804 = ( (~ ni37)  &  ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31806 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4950)  &  wire31804 ) ;
 assign wire31808 = ( (~ ni37)  &  (~ ni31)  &  (~ ni30) ) | ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31809 = ( ni36  &  (~ ni35)  &  wire31808 ) ;
 assign wire31813 = ( wire206  &  (~ nv3943)  &  (~ wire1180)  &  (~ n_n9177) ) ;
 assign wire31815 = ( (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31818 = ( (~ nv3943)  &  (~ wire1180)  &  (~ n_n9177)  &  wire31815 ) ;
 assign wire31819 = ( ni36  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31822 = ( (~ nv3943)  &  (~ wire1180)  &  (~ n_n9177)  &  wire31819 ) ;
 assign wire31824 = ( ni36  &  (~ ni35)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31826 = ( (~ nv3943)  &  (~ wire689)  &  (~ wire4950)  &  wire31824 ) ;
 assign wire31827 = ( n_n6710 ) | ( (~ wire689)  &  (~ wire4950)  &  wire31778 ) ;
 assign wire31828 = ( wire31827 ) | ( (~ nv3943)  &  (~ wire1180)  &  wire31809 ) ;
 assign wire31830 = ( wire31828 ) | ( (~ n_n9177)  &  wire31794 ) | ( (~ n_n9177)  &  wire31826 ) ;
 assign wire31833 = ( wire31830 ) | ( (~ n_n8968)  &  wire31774 ) | ( (~ n_n8968)  &  wire31822 ) ;
 assign wire31835 = ( (~ wire4862)  &  (~ wire31762)  &  wire31770 ) | ( (~ wire4862)  &  (~ wire31762)  &  wire31782 ) ;
 assign wire31836 = ( (~ wire4862)  &  (~ wire31762)  &  wire31786 ) | ( (~ wire4862)  &  (~ wire31762)  &  wire31798 ) ;
 assign wire31838 = ( wire31833 ) | ( (~ wire4862)  &  (~ wire31762)  &  wire31818 ) ;
 assign wire31839 = ( wire4757 ) | ( wire4763 ) | ( wire4767 ) | ( wire31835 ) ;
 assign wire31840 = ( wire4766 ) | ( wire4769 ) | ( wire31836 ) ;
 assign wire31842 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire31844 = ( (~ ni38)  &  ni37  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31846 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire31849 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire31851 = ( (~ ni36)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31852 = ( wire4680 ) | ( wire928 ) ;
 assign wire31855 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire31858 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire31859 = ( pi20  &  wire374  &  wire153 ) | ( (~ pi20)  &  wire374  &  wire153 ) ;
 assign wire31861 = ( wire170  &  wire913 ) | ( pi17  &  wire170  &  wire31350 ) ;
 assign wire31864 = ( wire3945 ) | ( wire3946 ) | ( wire3948 ) | ( wire31861 ) ;
 assign wire31865 = ( wire31864 ) | ( wire272  &  nv4575  &  wire31348 ) ;
 assign wire31866 = ( wire31865 ) | ( wire586  &  nv4630 ) ;
 assign wire31869 = ( wire3943 ) | ( wire3944 ) | ( wire3950 ) | ( wire31866 ) ;
 assign wire31870 = ( wire31869 ) | ( wire374  &  wire31257 ) | ( wire3959  &  wire31257 ) ;
 assign wire31875 = ( wire3934 ) | ( wire3937 ) | ( wire3938 ) | ( wire3939 ) ;
 assign wire31876 = ( wire3940 ) | ( wire3941 ) | ( wire3942 ) | ( wire31870 ) ;
 assign wire31878 = ( pi17  &  (~ pi16)  &  pi15  &  wire178 ) ;
 assign wire31880 = ( pi17  &  (~ pi16)  &  pi15  &  wire180 ) ;
 assign wire31882 = ( (~ pi16)  &  pi15  &  wire272 ) ;
 assign wire31883 = ( pi15  &  (~ pi16) ) ;
 assign wire31884 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire179 ) ;
 assign wire31885 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire182 ) ;
 assign wire31886 = ( pi17  &  pi16  &  pi15  &  wire180 ) ;
 assign wire31887 = ( pi17  &  pi16  &  pi15  &  wire178 ) ;
 assign wire31888 = ( (~ pi17)  &  pi16  &  pi15  &  wire182 ) ;
 assign wire31889 = ( (~ pi17)  &  pi16  &  pi15  &  wire179 ) ;
 assign wire31890 = ( (~ ni38)  &  (~ ni37)  &  (~ ni31)  &  (~ ni30) ) ;
 assign wire31891 = ( wire4804 ) | ( ni32  &  (~ ni30) ) ;
 assign wire31892 = ( (~ pi20)  &  (~ pi16)  &  pi15  &  wire153 ) ;
 assign wire31893 = ( wire4810 ) | ( ni32  &  (~ ni30) ) ;
 assign wire31894 = ( pi20  &  (~ pi16)  &  pi15  &  wire153 ) ;
 assign wire31895 = ( wire4778 ) | ( ni32  &  (~ ni30) ) ;
 assign wire31896 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire31897 = ( wire4784 ) | ( ni32  &  (~ ni30) ) ;
 assign wire31898 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire31899 = ( wire4047 ) | ( wire4779  &  wire31896 ) | ( wire31895  &  wire31896 ) ;
 assign wire31900 = ( wire170  &  wire915 ) | ( pi17  &  wire170  &  wire31883 ) ;
 assign wire31903 = ( wire3926 ) | ( wire3927 ) | ( wire3929 ) | ( wire31900 ) ;
 assign wire31905 = ( wire3916 ) | ( wire3931 ) | ( wire31903 ) ;
 assign wire31906 = ( wire31905 ) | ( nv4641  &  wire31892 ) ;
 assign wire31912 = ( wire3923 ) | ( wire3930 ) | ( nv4648  &  wire31894 ) ;
 assign wire31913 = ( wire3914 ) | ( wire3915 ) | ( wire3918 ) | ( wire31906 ) ;
 assign wire31914 = ( wire3919 ) | ( wire3920 ) | ( wire3921 ) | ( wire3922 ) ;
 assign wire31916 = ( wire31912 ) | ( wire31913 ) | ( wire31914 ) ;
 assign wire31917 = ( ni11  &  (~ ni9)  &  ni10 ) | ( ni12  &  (~ ni9)  &  ni10 ) ;
 assign wire31918 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire31917 ) ;
 assign wire31919 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire31921 = ( (~ wire175)  &  wire182  &  wire31919 ) ;
 assign wire31922 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire31924 = ( (~ wire175)  &  wire179  &  wire31922 ) ;
 assign wire31926 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  (~ wire175) ) ;
 assign wire31928 = ( (~ wire175)  &  wire395  &  wire182 ) ;
 assign wire31930 = ( (~ wire175)  &  wire395  &  wire179 ) ;
 assign wire31931 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire31932 = ( (~ pi20)  &  (~ pi16)  &  wire153  &  wire31931 ) ;
 assign wire31933 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire31934 = ( pi20  &  (~ pi16)  &  wire153  &  wire31933 ) ;
 assign wire31935 = ( pi17  &  ni32  &  ni30 ) ;
 assign wire31936 = ( wire1003 ) | ( wire272  &  n_n7877 ) ;
 assign wire31937 = ( wire31936 ) | ( pi17  &  wire178  &  n_n7893 ) ;
 assign wire31939 = ( (~ pi16)  &  pi15  &  (~ wire175) ) ;
 assign wire31940 = ( (~ pi20)  &  (~ wire175)  &  wire226  &  wire153 ) ;
 assign wire31941 = ( pi20  &  (~ wire175)  &  wire226  &  wire153 ) ;
 assign wire31943 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire31944 = ( pi16  &  pi15  &  (~ wire175) ) ;
 assign wire31945 = ( (~ pi17)  &  pi16  &  pi15  &  (~ wire175) ) ;
 assign wire31946 = ( (~ ni13)  &  ni14  &  (~ ni12)  &  wire485 ) ;
 assign wire31947 = ( pi15  &  (~ wire175)  &  wire152  &  wire154 ) ;
 assign wire31948 = ( ni32  &  ni30  &  (~ wire175) ) ;
 assign wire31949 = ( wire1178 ) | ( wire180  &  n_n7816 ) ;
 assign wire31950 = ( pi17  &  pi16  &  pi15  &  (~ wire175) ) ;
 assign wire31952 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire31954 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire31955 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire31956 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire182 ) ;
 assign wire31957 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire179 ) ;
 assign wire31958 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire31959 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire31960 = ( wire1003 ) | ( wire272  &  wire4613 ) | ( wire272  &  wire31347 ) ;
 assign wire31962 = ( (~ pi15)  &  (~ pi16) ) ;
 assign wire31964 = ( wire3906 ) | ( wire170  &  wire1071 ) ;
 assign wire31967 = ( wire3907 ) | ( wire586  &  wire4681 ) | ( wire586  &  wire31852 ) ;
 assign wire31968 = ( wire3893 ) | ( wire3902 ) | ( wire3903 ) | ( wire31964 ) ;
 assign wire31971 = ( wire3899 ) | ( wire3897 ) ;
 assign wire31972 = ( wire3896 ) | ( wire3900 ) | ( wire31967 ) | ( wire31968 ) ;
 assign wire31975 = ( wire3894 ) | ( wire3892 ) ;
 assign wire31976 = ( wire3891 ) | ( wire3895 ) | ( wire31971 ) | ( wire31972 ) ;
 assign wire31979 = ( wire170  &  wire31946 ) | ( wire416  &  wire31948 ) ;
 assign wire31983 = ( wire3874 ) | ( wire3882 ) | ( wire3883 ) | ( wire31979 ) ;
 assign wire31984 = ( wire3884 ) | ( wire31983 ) | ( n_n7808  &  wire31947 ) ;
 assign wire31985 = ( wire31984 ) | ( wire4805  &  wire31932 ) | ( wire31891  &  wire31932 ) ;
 assign wire31988 = ( wire3878 ) | ( wire3880 ) | ( n_n7905  &  wire31921 ) ;
 assign wire31989 = ( n_n7913  &  wire31924 ) | ( n_n7837  &  wire31928 ) ;
 assign wire31990 = ( wire3881 ) | ( wire31985 ) | ( n_n7845  &  wire31930 ) ;
 assign wire31992 = ( wire31988 ) | ( wire31989 ) | ( wire31990 ) ;
 assign wire31994 = ( wire3879 ) | ( wire3888 ) | ( wire31992 ) ;
 assign wire31995 = ( wire31994 ) | ( (~ wire175)  &  n_n8343 ) ;
 assign wire31996 = ( (~ ni11)  &  (~ ni9)  &  ni10 ) ;
 assign wire31997 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire31996 ) ;
 assign wire31998 = ( (~ pi17)  &  pi19  &  pi16  &  pi15 ) ;
 assign wire31999 = ( wire31998  &  wire387 ) ;
 assign wire32000 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire32001 = ( wire32000  &  wire387 ) ;
 assign wire32002 = ( pi21  &  pi22  &  pi20  &  pi15 ) ;
 assign wire32003 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire32002 ) ;
 assign wire32004 = ( (~ pi16)  &  (~ pi15) ) ;
 assign wire32005 = ( (~ pi17)  &  pi25  &  wire182  &  wire32004 ) ;
 assign wire32006 = ( (~ pi16)  &  pi15 ) ;
 assign wire32009 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire213 ) ;
 assign wire32010 = ( (~ pi17)  &  pi19  &  pi16  &  pi15 ) ;
 assign wire32011 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire32012 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  pi15 ) ;
 assign wire32013 = ( pi25  &  (~ pi16) ) | ( (~ pi21)  &  (~ pi16)  &  ni32 ) ;
 assign wire32014 = ( wire904  &  (~ pi15) ) ;
 assign wire32016 = ( (~ pi17)  &  ni32  &  ni30 ) ;
 assign wire32017 = ( pi25  &  ni32  &  ni30 ) ;
 assign wire32018 = ( wire611  &  wire32016 ) | ( wire153  &  wire32017 ) ;
 assign wire32019 = ( (~ pi17)  &  pi21  &  pi22  &  pi20 ) ;
 assign wire32022 = ( (~ pi16)  &  (~ pi15) ) ;
 assign wire32024 = ( (~ pi17)  &  ni32  &  ni30 ) ;
 assign wire32025 = ( pi25  &  ni32  &  ni30 ) ;
 assign wire32026 = ( wire387  &  wire32024 ) | ( wire153  &  wire32025 ) ;
 assign wire32027 = ( (~ pi16)  &  pi15 ) ;
 assign wire32029 = ( (~ pi17)  &  pi19  &  pi16  &  wire387 ) ;
 assign wire32030 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32032 = ( wire4652 ) | ( wire4655 ) | ( pi16  &  wire895 ) ;
 assign wire32033 = ( wire4651 ) | ( wire32032 ) ;
 assign wire32036 = ( n_n8890  &  wire32009 ) | ( n_n8890  &  wire153  &  wire32006 ) ;
 assign wire32037 = ( wire4596 ) | ( n_n8890  &  wire1110 ) | ( n_n8890  &  wire32003 ) ;
 assign wire32040 = ( wire32037 ) | ( (~ pi16)  &  (~ pi15)  &  wire895 ) ;
 assign wire32041 = ( wire4588 ) | ( wire32036 ) | ( wire226  &  wire895 ) ;
 assign wire32042 = ( wire4589 ) | ( wire4599 ) | ( wire32040 ) ;
 assign wire32043 = ( wire32041 ) | ( wire4606  &  wire32022 ) | ( wire4607  &  wire32022 ) ;
 assign wire32045 = ( wire32042 ) | ( wire32043 ) | ( n_n7845  &  wire31999 ) ;
 assign wire32046 = ( wire4590 ) | ( wire32045 ) ;
 assign wire32047 = ( (~ pi16)  &  pi15  &  wire1245 ) | ( pi16  &  pi15  &  wire1246 ) ;
 assign wire32050 = ( wire4583 ) | ( wire4585 ) | ( wire32047 ) ;
 assign wire32051 = ( wire4592 ) | ( wire32046 ) | ( pi15  &  wire1203 ) ;
 assign wire32053 = ( wire4591 ) | ( wire32050 ) | ( wire32051 ) ;
 assign wire32054 = ( ni11  &  (~ ni9)  &  (~ ni10) ) | ( ni12  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire32055 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire32054 ) ;
 assign wire32056 = ( ni33  &  (~ ni32)  &  ni29 ) ;
 assign wire32057 = ( (~ ni31)  &  (~ ni30)  &  wire32056 ) ;
 assign wire32059 = ( wire369  &  wire1053  &  wire1031 ) ;
 assign wire32061 = ( wire369  &  wire387  &  wire1031 ) ;
 assign wire32063 = ( wire369  &  wire1028  &  wire698 ) ;
 assign wire32064 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32065 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32066 = ( wire4505 ) | ( wire4779  &  wire32064 ) | ( wire31895  &  wire32064 ) ;
 assign wire32068 = ( (~ pi25)  &  pi16  &  wire369 ) ;
 assign wire32069 = ( (~ pi17)  &  pi19  &  pi16  &  wire369 ) ;
 assign wire32070 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire369 ) ;
 assign wire32074 = ( wire4510 ) | ( pi17  &  wire170 ) ;
 assign wire32076 = ( (~ pi25)  &  (~ pi16)  &  wire369 ) ;
 assign wire32077 = ( pi17  &  pi16  &  wire180 ) ;
 assign wire32078 = ( pi17  &  pi16  &  wire178 ) ;
 assign wire32079 = ( wire4484 ) | ( (~ pi19)  &  wire154  &  wire170 ) ;
 assign wire32081 = ( wire369  &  (~ pi25) ) ;
 assign wire32082 = ( wire369  &  (~ pi16) ) ;
 assign wire32083 = ( pi25  &  (~ pi16)  &  wire369 ) ;
 assign wire32084 = ( wire369  &  pi16 ) ;
 assign wire32085 = ( pi17  &  pi16  &  wire369 ) ;
 assign wire32086 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32089 = ( (~ pi17)  &  pi19  &  pi16  &  wire387 ) ;
 assign wire32090 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32091 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32092 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32094 = ( pi16  &  (~ pi25) ) ;
 assign wire32095 = ( pi17  &  (~ pi25)  &  pi16  &  wire152 ) ;
 assign wire32096 = ( wire850 ) | ( wire180  &  wire305 ) | ( wire180  &  wire4540 ) ;
 assign wire32097 = ( pi17  &  (~ pi25)  &  pi16 ) ;
 assign wire32099 = ( wire4520 ) | ( wire4525 ) | ( wire4526 ) ;
 assign wire32100 = ( wire32099 ) | ( nv4389  &  wire32095 ) ;
 assign wire32103 = ( wire4518 ) | ( wire4519 ) | ( wire4524 ) | ( wire32100 ) ;
 assign wire32104 = ( wire922 ) | ( wire4678 ) | ( wire502  &  wire32094 ) ;
 assign wire32106 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire611 ) ;
 assign wire32107 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire179 ) ;
 assign wire32109 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32110 = ( wire4556 ) | ( wire305  &  wire169 ) | ( wire169  &  wire4558 ) ;
 assign wire32111 = ( pi17  &  wire170 ) | ( wire272  &  nv4327 ) ;
 assign wire32112 = ( wire32111 ) | ( wire305  &  wire460 ) | ( wire460  &  wire4570 ) ;
 assign wire32113 = ( wire4554 ) | ( wire170  &  wire32109 ) | ( wire4857  &  wire32109 ) ;
 assign wire32114 = ( wire32113 ) | ( (~ pi16)  &  wire4606 ) | ( (~ pi16)  &  wire4607 ) ;
 assign wire32116 = ( wire4546 ) | ( wire4547 ) | ( wire32114 ) ;
 assign wire32118 = ( wire4548 ) | ( wire4553 ) | ( wire32116 ) ;
 assign wire32122 = ( wire4466 ) | ( wire4473 ) | ( wire4475 ) | ( wire4476 ) ;
 assign wire32124 = ( wire4462 ) | ( wire32122 ) | ( n_n7845  &  wire32061 ) ;
 assign wire32125 = ( wire4467 ) | ( wire4464 ) ;
 assign wire32126 = ( (~ pi16)  &  wire369  &  wire1245 ) | ( pi16  &  wire369  &  wire1246 ) ;
 assign wire32130 = ( wire4474 ) | ( wire32124 ) | ( wire32125 ) | ( wire32126 ) ;
 assign wire32132 = ( wire4465 ) | ( wire4470 ) | ( wire369  &  wire1203 ) ;
 assign wire32134 = ( wire4471 ) | ( wire4472 ) | ( wire32130 ) | ( wire32132 ) ;
 assign wire32137 = ( (~ ni11)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire32138 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire32137 ) ;
 assign wire32139 = ( n_n13895  &  wire265  &  wire186  &  (~ wire281) ) ;
 assign wire32141 = ( (~ wire175)  &  wire395  &  wire182 ) ;
 assign wire32143 = ( (~ wire175)  &  wire395  &  wire179 ) ;
 assign wire32144 = ( (~ pi17)  &  pi16  &  pi15  &  (~ wire175) ) ;
 assign wire32145 = ( (~ pi17)  &  (~ pi16)  &  wire179  &  wire369 ) ;
 assign wire32146 = ( (~ pi17)  &  (~ pi16)  &  wire182  &  wire369 ) ;
 assign wire32148 = ( (~ pi20)  &  (~ pi16)  &  wire369  &  wire153 ) ;
 assign wire32149 = ( pi20  &  (~ pi16)  &  wire369  &  wire153 ) ;
 assign wire32150 = ( pi17  &  pi19  &  pi16  &  wire369 ) | ( (~ pi17)  &  (~ pi19)  &  pi16  &  wire369 ) ;
 assign wire32151 = ( wire369  &  (~ pi16) ) ;
 assign wire32152 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire32155 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire32156 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire32157 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire32159 = ( (~ pi15)  &  wire302  &  wire170 ) | ( (~ pi15)  &  wire208  &  wire170 ) ;
 assign wire32161 = ( wire4428 ) | ( wire32159 ) | ( nv4389  &  wire586 ) ;
 assign wire32162 = ( wire32161 ) | ( wire305  &  wire32156 ) | ( wire4558  &  wire32156 ) ;
 assign wire32164 = ( wire4425 ) | ( wire4432 ) | ( wire32162 ) ;
 assign wire32165 = ( wire32164 ) | ( wire305  &  wire32152 ) | ( wire4562  &  wire32152 ) ;
 assign wire32168 = ( wire4421 ) | ( wire4422 ) | ( wire4423 ) | ( wire32165 ) ;
 assign wire32170 = ( wire170  &  wire32150 ) | ( pi19  &  wire170  &  wire32144 ) ;
 assign wire32171 = ( wire32170 ) | ( wire302  &  wire369  &  wire170 ) ;
 assign wire32173 = ( wire4418 ) | ( wire32171 ) | ( nv4401  &  wire32148 ) ;
 assign wire32177 = ( wire4410 ) | ( wire4411 ) | ( nv4409  &  wire32149 ) ;
 assign wire32178 = ( wire4406 ) | ( wire4407 ) | ( wire4409 ) | ( wire32173 ) ;
 assign wire32181 = ( wire4415 ) | ( wire4417 ) | ( wire32177 ) | ( wire32178 ) ;
 assign wire32182 = ( (~ ni11)  &  n_n13895  &  wire265  &  (~ wire281) ) ;
 assign wire32184 = ( n_n6711 ) | ( wire3639 ) | ( n_n6367  &  wire914 ) ;
 assign wire32186 = ( pi26  &  pi24  &  (~ ni14) ) ;
 assign wire32188 = ( wire818  &  wire1328  &  wire32186 ) ;
 assign wire32189 = ( (~ pi21)  &  nv6104 ) | ( pi21  &  (~ pi22)  &  nv6110 ) ;
 assign wire32191 = ( (~ pi26)  &  pi24  &  (~ ni14) ) ;
 assign wire32193 = ( wire818  &  wire1328  &  wire32191 ) ;
 assign wire32194 = ( pi26  &  pi24 ) ;
 assign wire32196 = ( wire264  &  wire331  &  (~ wire574)  &  wire32194 ) ;
 assign wire32197 = ( (~ pi26)  &  pi24 ) ;
 assign wire32199 = ( wire264  &  wire331  &  (~ wire574)  &  wire32197 ) ;
 assign wire32200 = ( pi21  &  (~ pi22)  &  pi24 ) ;
 assign wire32202 = ( wire359  &  wire1328  &  wire32200 ) ;
 assign wire32203 = ( (~ ni14)  &  (~ pi24) ) ;
 assign wire32206 = ( pi21  &  (~ pi22)  &  (~ pi26)  &  (~ pi24) ) ;
 assign wire32207 = ( pi21  &  pi22  &  (~ pi26)  &  (~ pi24) ) ;
 assign wire32208 = ( pi21  &  (~ pi22)  &  pi24 ) ;
 assign wire32210 = ( wire3641 ) | ( wire3645 ) | ( nv5285  &  wire32208 ) ;
 assign wire32212 = ( wire3642 ) | ( wire32210 ) | ( pi24  &  n_n6749 ) ;
 assign wire32214 = ( (~ pi23)  &  (~ ni7)  &  ni8 ) ;
 assign wire32216 = ( (~ wire175)  &  wire330  &  wire32214 ) ;
 assign wire32217 = ( pi23  &  (~ ni7)  &  ni8 ) ;
 assign wire32219 = ( (~ wire175)  &  wire330  &  wire32217 ) ;
 assign wire32221 = ( (~ pi24)  &  wire264  &  wire331  &  (~ wire574) ) ;
 assign wire32222 = ( pi15  &  (~ pi16) ) ;
 assign wire32223 = ( (~ pi17)  &  (~ pi24)  &  wire182  &  wire32222 ) ;
 assign wire32224 = ( pi15  &  pi16 ) ;
 assign wire32225 = ( (~ pi17)  &  (~ pi24)  &  wire179  &  wire32224 ) ;
 assign wire32226 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32227 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32228 = ( wire4277 ) | ( wire4805  &  wire32226 ) | ( wire31891  &  wire32226 ) ;
 assign wire32230 = ( (~ pi16)  &  pi15  &  pi24 ) ;
 assign wire32231 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32232 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32233 = ( wire4313 ) | ( wire4779  &  wire32231 ) | ( wire31895  &  wire32231 ) ;
 assign wire32235 = ( pi16  &  pi15  &  pi24 ) ;
 assign wire32236 = ( pi15  &  pi16 ) ;
 assign wire32237 = ( (~ pi17)  &  pi24  &  wire182  &  wire32236 ) ;
 assign wire32238 = ( pi15  &  (~ pi16) ) ;
 assign wire32239 = ( (~ pi17)  &  pi24  &  wire182  &  wire32238 ) ;
 assign wire32241 = ( (~ pi16)  &  pi15  &  (~ pi24) ) ;
 assign wire32243 = ( pi16  &  pi15  &  (~ pi24) ) ;
 assign wire32244 = ( pi24  &  pi21 ) ;
 assign wire32249 = ( (~ pi24)  &  pi15 ) ;
 assign wire32250 = ( (~ ni29)  &  wire158  &  wire178 ) | ( wire158  &  wire178  &  (~ n_n8862) ) ;
 assign wire32251 = ( (~ ni29)  &  wire158  &  wire180 ) | ( wire158  &  wire180  &  (~ n_n8862) ) ;
 assign wire32252 = ( (~ ni29)  &  wire158  &  wire152 ) | ( wire158  &  wire152  &  (~ n_n8862) ) ;
 assign wire32253 = ( wire250  &  wire306 ) | ( n_n7877  &  wire32252 ) ;
 assign wire32254 = ( wire158  &  wire180  &  wire306 ) | ( wire158  &  wire152  &  wire306 ) ;
 assign wire32256 = ( wire32253 ) | ( wire32254 ) | ( n_n7893  &  wire32250 ) ;
 assign wire32257 = ( pi24  &  pi15 ) ;
 assign wire32258 = ( (~ ni29)  &  wire178  &  wire154 ) | ( wire178  &  (~ n_n8862)  &  wire154 ) ;
 assign wire32260 = ( (~ ni29)  &  wire152  &  wire154 ) | ( wire152  &  (~ n_n8862)  &  wire154 ) ;
 assign wire32261 = ( wire251  &  wire306 ) | ( n_n7808  &  wire32260 ) ;
 assign wire32262 = ( wire180  &  wire154  &  wire306 ) | ( wire152  &  wire154  &  wire306 ) ;
 assign wire32264 = ( wire32261 ) | ( wire32262 ) | ( n_n7825  &  wire32258 ) ;
 assign wire32267 = ( (~ pi24)  &  pi15 ) ;
 assign wire32271 = ( (~ pi17)  &  pi16  &  pi24  &  wire179 ) ;
 assign wire32272 = ( (~ pi17)  &  (~ ni29)  &  wire182 ) | ( (~ pi17)  &  wire182  &  (~ n_n8862) ) ;
 assign wire32273 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32274 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32275 = ( wire203  &  wire306 ) | ( pi20  &  wire153  &  wire306 ) | ( (~ pi20)  &  wire153  &  wire306 ) ;
 assign wire32277 = ( wire4350 ) | ( wire4351 ) | ( wire32275 ) ;
 assign wire32280 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32281 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8862)  &  wire153 ) ;
 assign wire32282 = ( (~ pi17)  &  (~ ni29)  &  wire179 ) | ( (~ pi17)  &  wire179  &  (~ n_n8862) ) ;
 assign wire32283 = ( wire448  &  wire306 ) | ( (~ pi17)  &  wire179  &  wire306 ) ;
 assign wire32285 = ( wire4376 ) | ( wire4377 ) | ( wire32283 ) ;
 assign wire32288 = ( (~ pi17)  &  (~ pi16)  &  pi24  &  wire182 ) ;
 assign wire32289 = ( (~ pi17)  &  (~ pi16)  &  (~ pi24)  &  wire182 ) ;
 assign wire32290 = ( (~ pi17)  &  pi16  &  (~ pi24)  &  wire179 ) ;
 assign wire32291 = ( wire4342 ) | ( wire305  &  wire251 ) | ( wire251  &  wire4538 ) ;
 assign wire32292 = ( (~ ni29)  &  wire178  &  wire154 ) | ( wire178  &  (~ n_n8862)  &  wire154 ) ;
 assign wire32293 = ( (~ ni29)  &  wire180  &  wire154 ) | ( wire180  &  (~ n_n8862)  &  wire154 ) ;
 assign wire32294 = ( (~ ni29)  &  wire152  &  wire154 ) | ( wire152  &  (~ n_n8862)  &  wire154 ) ;
 assign wire32296 = ( wire180  &  wire154  &  wire306 ) | ( wire152  &  wire154  &  wire306 ) ;
 assign wire32297 = ( wire4345 ) | ( wire32296 ) | ( wire251  &  wire306 ) ;
 assign wire32299 = ( (~ ni29)  &  wire158  &  wire178 ) | ( wire158  &  wire178  &  (~ n_n8862) ) ;
 assign wire32300 = ( (~ ni29)  &  wire158  &  wire180 ) | ( wire158  &  wire180  &  (~ n_n8862) ) ;
 assign wire32301 = ( (~ ni29)  &  wire158  &  wire152 ) | ( wire158  &  wire152  &  (~ n_n8862) ) ;
 assign wire32303 = ( wire158  &  wire180  &  wire306 ) | ( wire158  &  wire152  &  wire306 ) ;
 assign wire32304 = ( wire4369 ) | ( wire32303 ) | ( wire250  &  wire306 ) ;
 assign wire32306 = ( wire4375 ) | ( wire305  &  wire250 ) | ( wire250  &  wire4570 ) ;
 assign wire32308 = ( (~ pi17)  &  wire338 ) | ( pi17  &  pi16  &  wire338 ) | ( pi17  &  (~ pi16)  &  wire338 ) ;
 assign wire32309 = ( wire32308 ) | ( wire306  &  wire32271 ) | ( wire4354  &  wire32271 ) ;
 assign wire32314 = ( wire3623 ) | ( wire3625 ) | ( wire3627 ) | ( wire3628 ) ;
 assign wire32315 = ( (~ pi16)  &  (~ pi24)  &  wire505 ) | ( pi16  &  (~ pi24)  &  wire502 ) ;
 assign wire32316 = ( wire3629 ) | ( wire3631 ) | ( wire3632 ) | ( wire32309 ) ;
 assign wire32318 = ( wire32315 ) | ( (~ pi24)  &  wire4374 ) | ( (~ pi24)  &  wire32306 ) ;
 assign wire32319 = ( wire3630 ) | ( wire32314 ) | ( wire32316 ) ;
 assign wire32322 = ( pi17  &  pi16  &  pi15  &  wire338 ) | ( (~ pi17)  &  pi16  &  pi15  &  wire338 ) | ( pi17  &  (~ pi16)  &  pi15  &  wire338 ) | ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire338 ) ;
 assign wire32325 = ( wire3610 ) | ( wire4286  &  wire32257 ) | ( wire32256  &  wire32257 ) ;
 assign wire32330 = ( wire3605 ) | ( wire3615 ) | ( wire3617 ) | ( wire32322 ) ;
 assign wire32331 = ( wire3606 ) | ( wire3607 ) | ( wire3609 ) | ( wire3618 ) ;
 assign wire32332 = ( wire3608 ) | ( wire3611 ) | ( wire3612 ) | ( wire32325 ) ;
 assign wire32334 = ( wire32330 ) | ( wire32331 ) | ( wire32332 ) ;
 assign wire32335 = ( (~ ni13)  &  ni14  &  (~ ni11)  &  (~ ni12) ) ;
 assign wire32338 = ( wire4293 ) | ( wire4294 ) | ( wire4296 ) ;
 assign wire32340 = ( pi24  &  wire359  &  wire1328 ) ;
 assign wire32341 = ( (~ pi21)  &  pi27 ) ;
 assign wire32344 = ( pi27  &  pi21  &  (~ pi22) ) ;
 assign wire32349 = ( pi21  &  pi22  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32352 = ( (~ ni7)  &  ni8  &  wire330  &  wire401 ) ;
 assign wire32354 = ( wire555  &  wire1328 ) ;
 assign wire32355 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32356 = ( pi23  &  (~ pi24)  &  wire213  &  wire32355 ) ;
 assign wire32357 = ( pi15  &  (~ wire289)  &  wire32356 ) ;
 assign wire32358 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32359 = ( (~ pi23)  &  wire213  &  wire32358 ) | ( pi24  &  wire213  &  wire32358 ) ;
 assign wire32360 = ( pi15  &  (~ wire289)  &  wire32359 ) ;
 assign wire32361 = ( (~ pi16)  &  (~ pi23) ) | ( (~ pi16)  &  pi24 ) ;
 assign wire32362 = ( pi15  &  (~ wire289)  &  wire32361 ) ;
 assign wire32363 = ( (~ pi17)  &  wire182  &  wire32362 ) ;
 assign wire32364 = ( (~ pi23)  &  (~ ni11)  &  ni12 ) | ( pi24  &  (~ ni11)  &  ni12 ) ;
 assign wire32365 = ( (~ ni13)  &  ni14  &  wire32364 ) ;
 assign wire32367 = ( (~ pi16)  &  pi15  &  (~ wire289)  &  wire1283 ) ;
 assign wire32368 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32369 = ( pi15  &  (~ wire289)  &  wire32368 ) ;
 assign wire32370 = ( (~ pi16)  &  pi23  &  (~ pi24) ) ;
 assign wire32371 = ( pi15  &  (~ wire289)  &  wire32370 ) ;
 assign wire32372 = ( (~ pi16)  &  (~ pi23) ) | ( (~ pi16)  &  pi24 ) ;
 assign wire32373 = ( pi15  &  (~ wire289)  &  wire32372 ) ;
 assign wire32375 = ( pi23  &  ni11  &  (~ wire574) ) ;
 assign wire32378 = ( pi23  &  (~ pi24)  &  (~ ni11)  &  ni12 ) ;
 assign wire32380 = ( (~ pi16)  &  pi15  &  (~ wire289) ) ;
 assign wire32382 = ( pi21  &  (~ pi22)  &  (~ ni13)  &  ni14 ) ;
 assign wire32384 = ( pi21  &  (~ pi22)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32386 = ( pi21  &  pi22  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32387 = ( pi26  &  (~ pi24)  &  wire32386 ) ;
 assign wire32388 = ( pi27  &  pi24  &  (~ ni13)  &  ni14 ) ;
 assign wire32390 = ( (~ pi24)  &  (~ ni13)  &  ni14 ) ;
 assign wire32391 = ( pi21  &  (~ pi22)  &  wire32390 ) ;
 assign wire32392 = ( pi24  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32394 = ( pi26  &  (~ pi24)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32395 = ( (~ pi26)  &  (~ pi24)  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32396 = ( pi24  &  (~ ni13)  &  ni14 ) ;
 assign wire32398 = ( pi24  &  (~ ni13)  &  (~ ni14) ) ;
 assign wire32401 = ( wire4257 ) | ( wire4258 ) | ( nv6124  &  wire32391 ) ;
 assign wire32402 = ( wire4265 ) | ( nv4938  &  wire914  &  wire32392 ) ;
 assign wire32403 = ( wire4260 ) | ( wire4263 ) | ( n_n7095  &  wire32398 ) ;
 assign wire32406 = ( wire4259 ) | ( wire32401 ) | ( wire32402 ) | ( wire32403 ) ;
 assign wire32408 = ( pi23  &  (~ ni11)  &  ni12 ) ;
 assign wire32409 = ( (~ pi23)  &  (~ ni11)  &  ni12 ) ;
 assign wire32410 = ( (~ pi23)  &  pi15  &  (~ wire289) ) | ( pi15  &  pi24  &  (~ wire289) ) ;
 assign wire32411 = ( pi23  &  pi15  &  (~ pi24)  &  (~ wire289) ) ;
 assign wire32413 = ( pi21  &  pi22  &  pi23  &  (~ pi24) ) ;
 assign wire32415 = ( (~ ni14)  &  ni11 ) | ( ni11  &  ni12 ) | ( ni13  &  ni14  &  ni11 ) ;
 assign wire32416 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32417 = ( pi23  &  (~ pi24)  &  wire213  &  wire32416 ) ;
 assign wire32418 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32419 = ( (~ pi23)  &  wire213  &  wire32418 ) | ( pi24  &  wire213  &  wire32418 ) ;
 assign wire32420 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32421 = ( pi16  &  pi23  &  (~ pi24) ) ;
 assign wire32422 = ( pi16  &  (~ pi23) ) | ( pi16  &  pi24 ) ;
 assign wire32424 = ( wire3577 ) | ( wire3580 ) | ( wire154  &  wire334 ) ;
 assign wire32425 = ( wire32424 ) | ( wire306  &  wire32417 ) | ( wire4354  &  wire32417 ) ;
 assign wire32427 = ( wire32425 ) | ( wire3582 ) ;
 assign wire32428 = ( wire3576 ) | ( wire3578 ) | ( wire502  &  wire32422 ) ;
 assign wire32430 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32431 = ( (~ pi23)  &  wire189  &  wire32430 ) | ( pi24  &  wire189  &  wire32430 ) ;
 assign wire32432 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32433 = ( pi23  &  (~ pi24)  &  wire189  &  wire32432 ) ;
 assign wire32434 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32437 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32438 = ( (~ pi16)  &  pi23  &  (~ pi24) ) ;
 assign wire32439 = ( (~ pi16)  &  (~ pi23) ) | ( (~ pi16)  &  pi24 ) ;
 assign wire32440 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32442 = ( wire3588 ) | ( wire3589 ) | ( wire334  &  wire32440 ) ;
 assign wire32443 = ( wire32442 ) | ( pi17  &  (~ pi16)  &  wire334 ) ;
 assign wire32444 = ( wire32443 ) | ( wire305  &  wire32431 ) | ( wire4564  &  wire32431 ) ;
 assign wire32446 = ( wire32444 ) | ( wire3593 ) ;
 assign wire32447 = ( wire3587 ) | ( wire3590 ) | ( wire505  &  wire32439 ) ;
 assign wire32449 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32450 = ( pi23  &  (~ pi24)  &  wire213  &  wire32449 ) ;
 assign wire32451 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32452 = ( (~ pi23)  &  wire213  &  wire32451 ) | ( pi24  &  wire213  &  wire32451 ) ;
 assign wire32453 = ( (~ pi17)  &  pi16  &  (~ wire160)  &  wire182 ) ;
 assign wire32454 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32455 = ( pi16  &  (~ pi23) ) | ( pi16  &  pi24 ) ;
 assign wire32456 = ( pi16  &  pi23  &  (~ pi24) ) ;
 assign wire32458 = ( wire3568 ) | ( wire3571 ) | ( wire154  &  wire334 ) ;
 assign wire32459 = ( wire32458 ) | ( wire4312  &  wire32456 ) | ( wire32233  &  wire32456 ) ;
 assign wire32463 = ( wire3567 ) | ( wire3569 ) | ( wire32459 ) ;
 assign wire32464 = ( wire3565 ) | ( wire3566 ) | ( wire3572 ) | ( wire3573 ) ;
 assign wire32467 = ( wire3548 ) | ( wire3553 ) | ( wire3554 ) | ( wire3559 ) ;
 assign wire32468 = ( wire3546 ) | ( nv6289  &  wire32415 ) ;
 assign wire32473 = ( wire3551 ) | ( wire3556 ) | ( wire3564 ) | ( wire32467 ) ;
 assign wire32474 = ( wire3552 ) | ( wire3555 ) | ( wire32468 ) | ( wire32473 ) ;
 assign wire32476 = ( wire3544 ) | ( wire3543 ) ;
 assign wire32477 = ( wire3547 ) | ( wire3545 ) ;
 assign wire32478 = ( wire3549 ) | ( wire32474 ) | ( wire449  &  wire32373 ) ;
 assign wire32481 = ( wire3558 ) | ( wire32476 ) | ( wire32477 ) | ( wire32478 ) ;
 assign wire32483 = ( wire3557 ) | ( wire3563 ) | ( wire32481 ) ;
 assign wire32485 = ( (~ ni9)  &  ni10  &  ni7  &  (~ ni8) ) ;
 assign wire32486 = ( (~ ni7)  &  ni8  &  wire264  &  wire401 ) ;
 assign wire32488 = ( wire377  &  wire453 ) | ( wire352  &  wire699 ) ;
 assign wire32489 = ( wire4400 ) | ( wire32488 ) | ( wire268  &  wire791 ) ;
 assign wire32490 = ( (~ ni10)  &  ni7 ) | ( ni7  &  ni8 ) | ( ni9  &  ni10  &  ni7 ) ;
 assign wire32491 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32492 = ( (~ pi23)  &  (~ pi24)  &  wire189  &  wire32491 ) ;
 assign wire32493 = ( pi15  &  (~ wire289)  &  wire32492 ) ;
 assign wire32494 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32495 = ( pi23  &  wire189  &  wire32494 ) | ( pi24  &  wire189  &  wire32494 ) ;
 assign wire32496 = ( pi15  &  (~ wire289)  &  wire32495 ) ;
 assign wire32497 = ( pi23  &  (~ ni11)  &  ni12 ) | ( pi24  &  (~ ni11)  &  ni12 ) ;
 assign wire32498 = ( (~ ni13)  &  ni14  &  wire32497 ) ;
 assign wire32499 = ( (~ pi16)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32500 = ( pi15  &  (~ wire289)  &  wire32499 ) ;
 assign wire32501 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32502 = ( pi15  &  (~ wire289)  &  wire32501 ) ;
 assign wire32503 = ( (~ pi16)  &  pi23 ) | ( (~ pi16)  &  pi24 ) ;
 assign wire32504 = ( pi15  &  (~ wire289)  &  wire32503 ) ;
 assign wire32505 = ( (~ pi23)  &  (~ pi24)  &  (~ ni11)  &  ni12 ) ;
 assign wire32507 = ( (~ pi16)  &  pi15  &  (~ wire289) ) ;
 assign wire32508 = ( (~ pi23)  &  (~ ni11)  &  ni12 ) ;
 assign wire32509 = ( pi23  &  (~ ni11)  &  ni12 ) ;
 assign wire32510 = ( pi23  &  pi15  &  (~ wire289) ) | ( pi15  &  pi24  &  (~ wire289) ) ;
 assign wire32511 = ( (~ pi23)  &  pi15  &  (~ pi24)  &  (~ wire289) ) ;
 assign wire32513 = ( pi16  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32515 = ( (~ pi17)  &  pi19  &  wire213  &  wire32513 ) ;
 assign wire32516 = ( pi16  &  pi23 ) | ( pi16  &  pi24 ) ;
 assign wire32518 = ( (~ pi17)  &  pi19  &  wire213  &  wire32516 ) ;
 assign wire32519 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32522 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire32523 = ( pi16  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32524 = ( pi16  &  pi23 ) | ( pi16  &  pi24 ) ;
 assign wire32525 = ( (~ pi17)  &  (~ pi19)  &  pi16 ) | ( (~ pi17)  &  pi20  &  pi16 ) ;
 assign wire32527 = ( wire4332 ) | ( wire4333 ) | ( wire339  &  wire32525 ) ;
 assign wire32528 = ( wire32527 ) | ( pi17  &  pi16  &  wire339 ) ;
 assign wire32529 = ( wire32528 ) | ( wire306  &  wire32515 ) | ( wire4354  &  wire32515 ) ;
 assign wire32531 = ( wire32529 ) | ( wire4338 ) ;
 assign wire32532 = ( wire4331 ) | ( wire4334 ) | ( wire502  &  wire32524 ) ;
 assign wire32534 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32535 = ( (~ pi23)  &  (~ pi24)  &  wire189  &  wire32534 ) ;
 assign wire32536 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32537 = ( pi23  &  wire189  &  wire32536 ) | ( pi24  &  wire189  &  wire32536 ) ;
 assign wire32538 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32539 = ( (~ pi16)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32540 = ( (~ pi16)  &  pi23 ) | ( (~ pi16)  &  pi24 ) ;
 assign wire32542 = ( wire4358 ) | ( wire4361 ) | ( wire158  &  wire339 ) ;
 assign wire32543 = ( wire32542 ) | ( wire306  &  wire32535 ) | ( wire4387  &  wire32535 ) ;
 assign wire32545 = ( wire32543 ) | ( wire4362 ) ;
 assign wire32546 = ( wire4357 ) | ( wire4359 ) | ( wire505  &  wire32540 ) ;
 assign wire32548 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32549 = ( (~ pi23)  &  (~ pi24)  &  wire189  &  wire32548 ) ;
 assign wire32550 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32551 = ( pi23  &  wire189  &  wire32550 ) | ( pi24  &  wire189  &  wire32550 ) ;
 assign wire32552 = ( pi16  &  pi23 ) | ( pi16  &  pi24 ) ;
 assign wire32553 = ( (~ pi17)  &  wire179  &  wire32552 ) ;
 assign wire32554 = ( pi16  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire32555 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32556 = ( pi16  &  pi23 ) | ( pi16  &  pi24 ) ;
 assign wire32558 = ( wire4303 ) | ( wire4305 ) | ( wire154  &  wire339 ) ;
 assign wire32559 = ( wire32558 ) | ( wire4504  &  wire32556 ) | ( wire32066  &  wire32556 ) ;
 assign wire32563 = ( wire4301 ) | ( wire4302 ) | ( wire32559 ) ;
 assign wire32564 = ( wire4299 ) | ( wire4300 ) | ( wire4306 ) | ( wire4307 ) ;
 assign wire32567 = ( wire4244 ) | ( wire4246 ) | ( wire4247 ) | ( wire4252 ) ;
 assign wire32568 = ( wire4242 ) | ( nv5862  &  wire555 ) ;
 assign wire32571 = ( wire4248 ) | ( wire4249 ) | ( wire32567 ) | ( wire32568 ) ;
 assign wire32573 = ( wire4241 ) | ( wire4286  &  wire32511 ) | ( wire32256  &  wire32511 ) ;
 assign wire32576 = ( wire4240 ) | ( wire4243 ) | ( wire4250 ) | ( wire32571 ) ;
 assign wire32578 = ( wire4245 ) | ( wire4255 ) | ( wire32573 ) | ( wire32576 ) ;
 assign wire32580 = ( (~ ni9)  &  (~ ni10)  &  (~ ni7)  &  ni8 ) ;
 assign wire32581 = ( ni9  &  (~ ni7)  &  ni8 ) ;
 assign wire32583 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32586 = ( wire370  &  wire181  &  wire833  &  wire32583 ) ;
 assign wire32587 = ( wire4089 ) | ( pi21  &  (~ pi22)  &  nv5285 ) ;
 assign wire32589 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32591 = ( wire370  &  wire833  &  wire32589 ) ;
 assign wire32592 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32595 = ( wire370  &  wire181  &  wire833  &  wire32592 ) ;
 assign wire32596 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32599 = ( wire370  &  wire181  &  wire833  &  wire32596 ) ;
 assign wire32602 = ( (~ pi17)  &  (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32605 = ( (~ pi17)  &  (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32606 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32608 = ( wire370  &  wire833  &  wire32606 ) ;
 assign wire32609 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32611 = ( wire370  &  wire833  &  wire32609 ) ;
 assign wire32613 = ( (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32614 = ( pi20  &  pi25  &  wire153  &  wire32613 ) ;
 assign wire32616 = ( pi17  &  (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32617 = ( wire4077 ) | ( (~ pi17)  &  (~ pi19)  &  wire373 ) ;
 assign wire32619 = ( (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32621 = ( pi17  &  (~ pi16)  &  wire370  &  wire833 ) ;
 assign wire32622 = ( wire833  &  wire370 ) ;
 assign wire32624 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32627 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32628 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32629 = ( pi21  &  pi22  &  pi25  &  wire32628 ) ;
 assign wire32630 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32631 = ( pi21  &  pi22  &  pi25  &  wire32630 ) ;
 assign wire32633 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire32634 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire32635 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32636 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32638 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire32639 = ( wire3702 ) | ( (~ pi17)  &  (~ pi19)  &  wire440 ) ;
 assign wire32640 = ( n_n7877  &  wire393 ) | ( wire440  &  wire32634 ) ;
 assign wire32641 = ( wire32640 ) | ( wire158  &  wire178  &  wire280 ) ;
 assign wire32643 = ( wire4090  &  wire32635 ) | ( wire32587  &  wire32635 ) | ( wire4090  &  wire32636 ) | ( wire32587  &  wire32636 ) ;
 assign wire32645 = ( wire3691 ) | ( wire4811  &  wire32631 ) | ( wire31893  &  wire32631 ) ;
 assign wire32647 = ( wire3698 ) | ( wire32641 ) | ( wire32643 ) ;
 assign wire32648 = ( wire964 ) | ( wire3687 ) | ( wire3696 ) | ( wire32645 ) ;
 assign wire32649 = ( wire32647 ) | ( wire181  &  n_n7905  &  wire32624 ) ;
 assign wire32651 = ( wire3690 ) | ( wire158  &  wire345  &  n_n7893 ) ;
 assign wire32652 = ( wire32648 ) | ( wire32649 ) | ( n_n7885  &  wire32629 ) ;
 assign wire32654 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire32655 = ( pi21  &  pi22  &  pi25  &  wire32654 ) ;
 assign wire32657 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire32659 = ( (~ pi17)  &  pi25  &  pi16  &  wire179 ) ;
 assign wire32660 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32661 = ( pi21  &  pi22  &  pi25  &  wire32660 ) ;
 assign wire32662 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire32663 = ( pi21  &  pi22  &  pi25  &  wire32662 ) ;
 assign wire32664 = ( pi16  &  (~ pi17) ) ;
 assign wire32665 = ( pi17  &  pi25  &  pi16  &  wire180 ) ;
 assign wire32666 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32667 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire32668 = ( wire908 ) | ( wire4082 ) | ( wire183  &  wire280 ) ;
 assign wire32669 = ( wire4090  &  wire32657 ) | ( wire32587  &  wire32657 ) | ( wire4090  &  wire32666 ) | ( wire32587  &  wire32666 ) ;
 assign wire32671 = ( wire3676 ) | ( wire4785  &  wire32663 ) | ( wire31897  &  wire32663 ) ;
 assign wire32672 = ( wire32668 ) | ( wire3682 ) ;
 assign wire32673 = ( wire3679 ) | ( wire3681 ) | ( wire32669 ) ;
 assign wire32676 = ( n_n7837  &  wire32655 ) | ( n_n7845  &  wire32659 ) ;
 assign wire32677 = ( n_n7825  &  wire32661 ) | ( n_n7816  &  wire32665 ) ;
 assign wire32678 = ( wire3680 ) | ( wire32671 ) | ( wire32672 ) | ( wire32673 ) ;
 assign wire32680 = ( wire32676 ) | ( wire32677 ) | ( wire32678 ) ;
 assign wire32681 = ( wire833  &  wire369 ) ;
 assign wire32682 = ( wire833  &  wire370 ) ;
 assign wire32684 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire32685 = ( pi21  &  pi22  &  pi25  &  wire32684 ) ;
 assign wire32687 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  pi16 ) ;
 assign wire32689 = ( (~ pi17)  &  pi25  &  pi16  &  wire182 ) ;
 assign wire32690 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32691 = ( pi21  &  pi22  &  pi25  &  wire32690 ) ;
 assign wire32692 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32693 = ( pi21  &  pi22  &  pi25  &  wire32692 ) ;
 assign wire32694 = ( pi16  &  (~ pi17) ) ;
 assign wire32695 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32696 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32697 = ( pi20  &  pi25  &  pi16  &  wire153 ) ;
 assign wire32700 = ( wire4090  &  wire32687 ) | ( wire32587  &  wire32687 ) | ( wire4090  &  wire32695 ) | ( wire32587  &  wire32695 ) ;
 assign wire32702 = ( wire922 ) | ( wire4066 ) | ( wire4067 ) ;
 assign wire32703 = ( wire965 ) | ( wire4070 ) | ( wire4073 ) ;
 assign wire32704 = ( wire4069 ) | ( wire4072 ) | ( wire32700 ) ;
 assign wire32706 = ( wire32702 ) | ( wire32703 ) | ( wire32704 ) ;
 assign wire32709 = ( wire4062 ) | ( wire32706 ) | ( wire154  &  wire1308 ) ;
 assign wire32710 = ( wire833  &  wire370 ) ;
 assign wire32711 = ( ni13  &  wire833 ) | ( (~ ni14)  &  wire833 ) | ( ni12  &  wire833 ) ;
 assign wire32712 = ( (~ pi17)  &  pi16  &  pi15 ) ;
 assign wire32714 = ( pi25  &  wire182  &  wire268  &  wire32712 ) ;
 assign wire32715 = ( (~ pi17)  &  pi16  &  pi15 ) ;
 assign wire32717 = ( pi25  &  wire179  &  wire268  &  wire32715 ) ;
 assign wire32720 = ( wire4151 ) | ( pi27  &  pi25  &  n_n8085 ) ;
 assign wire32722 = ( (~ pi17)  &  pi16  &  pi15  &  wire268 ) ;
 assign wire32724 = ( pi25  &  wire180  &  wire403  &  wire268 ) ;
 assign wire32726 = ( pi25  &  wire178  &  wire403  &  wire268 ) ;
 assign wire32727 = ( pi16  &  pi15  &  wire268 ) ;
 assign wire32728 = ( pi17  &  pi16  &  pi15  &  wire268 ) ;
 assign wire32729 = ( pi16  &  pi15  &  wire268 ) ;
 assign wire32730 = ( wire485  &  wire268 ) ;
 assign wire32731 = ( pi15  &  wire152  &  wire154  &  wire268 ) ;
 assign wire32733 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire32735 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire32736 = ( pi17  &  pi25  &  (~ pi16)  &  wire180 ) ;
 assign wire32737 = ( wire1279 ) | ( wire4142 ) | ( wire194  &  wire249 ) ;
 assign wire32740 = ( wire4113 ) | ( wire4117 ) | ( wire4118 ) | ( wire32737 ) ;
 assign wire32741 = ( n_n7905  &  wire32733 ) | ( n_n7885  &  wire32736 ) ;
 assign wire32742 = ( wire32740 ) | ( (~ pi16)  &  wire4802 ) | ( (~ pi16)  &  wire4803 ) ;
 assign wire32746 = ( (~ pi17)  &  pi25  &  pi16  &  wire182 ) ;
 assign wire32748 = ( (~ pi17)  &  pi25  &  pi16  &  wire179 ) ;
 assign wire32749 = ( pi16  &  (~ pi17) ) ;
 assign wire32750 = ( pi17  &  pi25  &  pi16  &  wire178 ) ;
 assign wire32751 = ( wire4129 ) | ( wire311  &  wire4681 ) | ( wire311  &  wire31852 ) ;
 assign wire32752 = ( wire32751 ) | ( wire152  &  wire154  &  wire249 ) ;
 assign wire32754 = ( wire4127 ) | ( pi16  &  wire4659 ) | ( pi16  &  wire4660 ) ;
 assign wire32756 = ( wire4123 ) | ( wire4128 ) | ( wire32752 ) | ( wire32754 ) ;
 assign wire32758 = ( wire4124 ) | ( wire4122 ) ;
 assign wire32759 = ( wire4121 ) | ( wire32756 ) | ( wire154  &  wire1308 ) ;
 assign wire32761 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire179 ) ;
 assign wire32763 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire32764 = ( pi17  &  pi25  &  (~ pi16)  &  wire178 ) ;
 assign wire32765 = ( wire1351 ) | ( wire4142 ) | ( wire194  &  wire249 ) ;
 assign wire32766 = ( wire4134 ) | ( (~ pi16)  &  wire4606 ) | ( (~ pi16)  &  wire4607 ) ;
 assign wire32769 = ( wire4138 ) | ( wire4139 ) | ( wire32765 ) | ( wire32766 ) ;
 assign wire32771 = ( wire4135 ) | ( (~ pi17)  &  (~ pi16)  &  wire1290 ) ;
 assign wire32772 = ( wire4132 ) | ( wire32769 ) | ( wire158  &  wire1292 ) ;
 assign wire32774 = ( pi19  &  (~ pi20)  &  pi16  &  pi15 ) ;
 assign wire32776 = ( (~ pi17)  &  (~ ni14)  &  wire181  &  wire32774 ) ;
 assign wire32777 = ( wire4235 ) | ( pi21  &  (~ pi22)  &  nv4938 ) ;
 assign wire32779 = ( pi19  &  (~ pi20)  &  pi16  &  pi15 ) ;
 assign wire32780 = ( (~ pi17)  &  (~ ni14)  &  wire32779 ) ;
 assign wire32782 = ( (~ pi17)  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32783 = ( pi25  &  wire182  &  wire32782 ) ;
 assign wire32784 = ( (~ pi19)  &  pi20  &  (~ ni14) ) ;
 assign wire32786 = ( wire403  &  wire181  &  wire32784 ) ;
 assign wire32787 = ( pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32789 = ( wire228  &  wire181  &  wire32787 ) ;
 assign wire32791 = ( (~ pi17)  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32793 = ( (~ pi19)  &  pi20  &  (~ ni14)  &  wire403 ) ;
 assign wire32794 = ( pi17  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32795 = ( pi25  &  wire178  &  wire32794 ) ;
 assign wire32796 = ( pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32798 = ( pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32799 = ( pi17  &  pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32800 = ( wire4231 ) | ( (~ pi17)  &  (~ pi19)  &  wire372 ) ;
 assign wire32801 = ( pi16  &  pi15  &  (~ ni14) ) ;
 assign wire32803 = ( pi15  &  (~ ni14)  &  wire152  &  wire154 ) ;
 assign wire32805 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32806 = ( pi21  &  pi22  &  pi25  &  wire32805 ) ;
 assign wire32808 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire32809 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32810 = ( pi21  &  pi22  &  pi25  &  wire32809 ) ;
 assign wire32811 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32812 = ( pi21  &  pi22  &  pi25  &  wire32811 ) ;
 assign wire32814 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire32815 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire32816 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32817 = ( (~ pi17)  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32818 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire32819 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire32820 = ( pi20  &  (~ pi16)  &  wire153 ) ;
 assign wire32821 = ( wire442  &  wire32815 ) | ( wire187  &  wire32818 ) ;
 assign wire32823 = ( wire4182 ) | ( wire32821 ) | ( n_n7877  &  wire393 ) ;
 assign wire32825 = ( wire4236  &  wire32808 ) | ( wire32777  &  wire32808 ) | ( wire4236  &  wire32816 ) | ( wire32777  &  wire32816 ) ;
 assign wire32826 = ( wire4179 ) | ( wire4805  &  wire32812 ) | ( wire31891  &  wire32812 ) ;
 assign wire32827 = ( wire4176 ) | ( wire4811  &  wire32819 ) | ( wire31893  &  wire32819 ) ;
 assign wire32828 = ( wire960 ) | ( wire4184 ) | ( wire32823 ) ;
 assign wire32831 = ( n_n7905  &  wire32806 ) | ( n_n7885  &  wire32810 ) ;
 assign wire32832 = ( wire32825 ) | ( wire32826 ) | ( wire32827 ) | ( wire32828 ) ;
 assign wire32836 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire32837 = ( pi21  &  pi22  &  pi25  &  wire32836 ) ;
 assign wire32839 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire32841 = ( (~ pi17)  &  pi25  &  pi16  &  wire179 ) ;
 assign wire32842 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32843 = ( pi21  &  pi22  &  pi25  &  wire32842 ) ;
 assign wire32844 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire32845 = ( pi21  &  pi22  &  pi25  &  wire32844 ) ;
 assign wire32846 = ( pi16  &  (~ pi17) ) ;
 assign wire32847 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  pi16 ) ;
 assign wire32848 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire32849 = ( (~ pi20)  &  pi25  &  pi16  &  wire153 ) ;
 assign wire32850 = ( wire922 ) | ( wire257  &  wire227 ) ;
 assign wire32853 = ( wire4236  &  wire32839 ) | ( wire32777  &  wire32839 ) | ( wire4236  &  wire32847 ) | ( wire32777  &  wire32847 ) ;
 assign wire32855 = ( wire4193 ) | ( wire4197 ) | ( wire4201 ) | ( wire32850 ) ;
 assign wire32857 = ( wire4196 ) | ( wire4200 ) | ( wire32853 ) ;
 assign wire32859 = ( wire4194 ) | ( wire4199 ) | ( wire32855 ) | ( wire32857 ) ;
 assign wire32861 = ( wire4192 ) | ( wire4191 ) ;
 assign wire32862 = ( wire4189 ) | ( wire32859 ) | ( wire154  &  wire1308 ) ;
 assign wire32864 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32865 = ( pi21  &  pi22  &  pi25  &  wire32864 ) ;
 assign wire32867 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32868 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32869 = ( pi21  &  pi22  &  pi25  &  wire32868 ) ;
 assign wire32870 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32871 = ( pi21  &  pi22  &  pi25  &  wire32870 ) ;
 assign wire32873 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire32874 = ( pi17  &  (~ pi19)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32875 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire32876 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire32879 = ( wire4236  &  wire32867 ) | ( wire32777  &  wire32867 ) | ( wire4236  &  wire32874 ) | ( wire32777  &  wire32874 ) ;
 assign wire32881 = ( wire1351 ) | ( wire4209 ) | ( wire4211 ) ;
 assign wire32882 = ( wire960 ) | ( wire4214 ) | ( wire4216 ) ;
 assign wire32883 = ( wire4213 ) | ( wire4217 ) | ( wire32879 ) ;
 assign wire32885 = ( wire32881 ) | ( wire32882 ) | ( wire32883 ) ;
 assign wire32887 = ( wire4208 ) | ( (~ pi17)  &  (~ pi16)  &  wire1290 ) ;
 assign wire32888 = ( wire4206 ) | ( wire32885 ) | ( wire158  &  wire1292 ) ;
 assign wire32890 = ( wire4165 ) | ( wire4167 ) | ( wire274  &  wire32803 ) ;
 assign wire32891 = ( wire4236  &  wire32780 ) | ( wire32777  &  wire32780 ) | ( wire4236  &  wire32793 ) | ( wire32777  &  wire32793 ) ;
 assign wire32893 = ( wire32890 ) | ( wire4785  &  wire32789 ) | ( wire31897  &  wire32789 ) ;
 assign wire32894 = ( wire4163 ) | ( wire4158 ) ;
 assign wire32895 = ( wire4161 ) | ( wire4164 ) | ( wire32891 ) ;
 assign wire32898 = ( n_n7845  &  wire32776 ) | ( n_n7837  &  wire32783 ) ;
 assign wire32899 = ( n_n7816  &  wire32786 ) | ( n_n7825  &  wire32795 ) ;
 assign wire32900 = ( wire4162 ) | ( wire32893 ) | ( wire32894 ) | ( wire32895 ) ;
 assign wire32902 = ( wire32898 ) | ( wire32899 ) | ( wire32900 ) ;
 assign wire32903 = ( wire32902 ) | ( pi15  &  (~ ni14)  &  n_n7945 ) ;
 assign wire32904 = ( wire32903 ) | ( wire765  &  wire32861 ) | ( wire765  &  wire32862 ) ;
 assign wire32905 = ( wire4102 ) | ( wire848  &  n_n7808  &  wire311 ) ;
 assign wire32906 = ( wire32905 ) | ( wire249  &  wire32731 ) ;
 assign wire32909 = ( wire4096 ) | ( wire4100 ) | ( wire4101 ) | ( wire32906 ) ;
 assign wire32910 = ( n_n7837  &  wire32714 ) | ( n_n7845  &  wire32717 ) ;
 assign wire32911 = ( n_n7816  &  wire32724 ) | ( n_n7825  &  wire32726 ) ;
 assign wire32912 = ( wire32909 ) | ( wire1329  &  wire32727 ) | ( wire4776  &  wire32727 ) ;
 assign wire32914 = ( wire32910 ) | ( wire32911 ) | ( wire32912 ) ;
 assign wire32915 = ( wire32914 ) | ( pi15  &  n_n7702  &  wire268 ) ;
 assign wire32916 = ( wire32915 ) | ( wire845  &  wire32758 ) | ( wire845  &  wire32759 ) ;
 assign wire32919 = ( wire4107 ) | ( wire4108 ) | ( wire4109 ) | ( wire32916 ) ;
 assign wire32920 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32921 = ( pi27  &  wire189  &  wire32920 ) | ( (~ pi26)  &  wire189  &  wire32920 ) ;
 assign wire32922 = ( ni11  &  wire369  &  wire32921 ) ;
 assign wire32923 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32924 = ( (~ pi27)  &  pi26  &  wire189  &  wire32923 ) ;
 assign wire32925 = ( ni11  &  wire369  &  wire32924 ) ;
 assign wire32927 = ( (~ pi16)  &  ni11  &  wire369  &  wire1120 ) ;
 assign wire32929 = ( (~ pi16)  &  ni11  &  wire369  &  wire1093 ) ;
 assign wire32930 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire32931 = ( ni11  &  wire369  &  wire32930 ) ;
 assign wire32932 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32933 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32934 = ( wire4006 ) | ( wire4805  &  wire32932 ) | ( wire31891  &  wire32932 ) ;
 assign wire32935 = ( (~ pi27)  &  pi26  &  (~ pi16) ) ;
 assign wire32936 = ( ni11  &  wire369  &  wire32935 ) ;
 assign wire32937 = ( pi27  &  (~ pi16) ) | ( (~ pi26)  &  (~ pi16) ) ;
 assign wire32938 = ( ni11  &  wire369  &  wire32937 ) ;
 assign wire32939 = ( (~ pi16)  &  ni11  &  wire369 ) ;
 assign wire32941 = ( pi27  &  ni11  &  wire369 ) | ( (~ pi26)  &  ni11  &  wire369 ) ;
 assign wire32942 = ( (~ ni29)  &  wire158  &  wire178 ) | ( wire158  &  wire178  &  (~ n_n8352) ) ;
 assign wire32943 = ( (~ ni29)  &  wire158  &  wire180 ) | ( wire158  &  wire180  &  (~ n_n8352) ) ;
 assign wire32944 = ( (~ ni29)  &  wire158  &  wire152 ) | ( wire158  &  wire152  &  (~ n_n8352) ) ;
 assign wire32945 = ( wire250  &  wire375 ) | ( n_n7877  &  wire32944 ) ;
 assign wire32946 = ( wire158  &  wire180  &  wire375 ) | ( wire158  &  wire152  &  wire375 ) ;
 assign wire32948 = ( wire32945 ) | ( wire32946 ) | ( n_n7893  &  wire32942 ) ;
 assign wire32949 = ( (~ pi27)  &  pi26  &  ni11  &  wire369 ) ;
 assign wire32950 = ( pi17  &  (~ pi16)  &  ni11  &  wire369 ) ;
 assign wire32951 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32952 = ( pi27  &  wire189  &  wire32951 ) | ( (~ pi26)  &  wire189  &  wire32951 ) ;
 assign wire32953 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32954 = ( (~ pi27)  &  pi26  &  wire189  &  wire32953 ) ;
 assign wire32955 = ( (~ pi17)  &  pi16  &  wire155  &  wire179 ) ;
 assign wire32956 = ( (~ pi17)  &  pi16  &  (~ wire155)  &  wire179 ) ;
 assign wire32957 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire32958 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32959 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32960 = ( pi20  &  wire153  &  wire375 ) | ( (~ pi20)  &  wire153  &  wire375 ) ;
 assign wire32962 = ( (~ pi27)  &  pi26  &  pi16 ) ;
 assign wire32963 = ( pi27  &  pi16 ) | ( (~ pi26)  &  pi16 ) ;
 assign wire32964 = ( wire3827 ) | ( wire374  &  wire251 ) | ( wire251  &  wire3965 ) ;
 assign wire32965 = ( (~ ni29)  &  wire178  &  wire154 ) | ( wire178  &  (~ n_n8352)  &  wire154 ) ;
 assign wire32966 = ( (~ ni29)  &  wire152  &  wire154 ) | ( wire152  &  (~ n_n8352)  &  wire154 ) ;
 assign wire32967 = ( (~ ni29)  &  wire180  &  wire154 ) | ( wire180  &  (~ n_n8352)  &  wire154 ) ;
 assign wire32969 = ( wire180  &  wire154  &  wire375 ) | ( wire152  &  wire154  &  wire375 ) ;
 assign wire32970 = ( wire3829 ) | ( wire32969 ) | ( wire251  &  wire375 ) ;
 assign wire32973 = ( wire3727 ) | ( wire3730 ) | ( wire154  &  wire221 ) ;
 assign wire32975 = ( wire3728 ) | ( wire3729 ) | ( wire32973 ) ;
 assign wire32976 = ( wire32975 ) | ( wire374  &  wire32952 ) | ( wire3963  &  wire32952 ) ;
 assign wire32978 = ( wire3732 ) | ( wire375  &  wire32956 ) | ( wire3840  &  wire32956 ) ;
 assign wire32979 = ( wire3724 ) | ( wire3725 ) | ( wire32976 ) ;
 assign wire32982 = ( pi27  &  wire213  &  wire698 ) | ( (~ pi26)  &  wire213  &  wire698 ) ;
 assign wire32984 = ( (~ pi27)  &  pi26  &  wire213  &  wire698 ) ;
 assign wire32985 = ( pi27  &  (~ pi16) ) | ( (~ pi26)  &  (~ pi16) ) ;
 assign wire32986 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32987 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire32989 = ( (~ pi27)  &  pi26  &  (~ pi16) ) ;
 assign wire32990 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire32991 = ( (~ pi17)  &  (~ pi16)  &  (~ wire155)  &  wire182 ) ;
 assign wire32992 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire32994 = ( (~ pi17)  &  (~ pi16)  &  wire155  &  wire182 ) ;
 assign wire32995 = ( wire3856 ) | ( wire374  &  wire250 ) | ( wire250  &  wire3959 ) ;
 assign wire32996 = ( (~ ni29)  &  wire158  &  wire178 ) | ( wire158  &  wire178  &  (~ n_n8352) ) ;
 assign wire32997 = ( (~ ni29)  &  wire158  &  wire180 ) | ( wire158  &  wire180  &  (~ n_n8352) ) ;
 assign wire32998 = ( (~ ni29)  &  wire158  &  wire152 ) | ( wire158  &  wire152  &  (~ n_n8352) ) ;
 assign wire33000 = ( wire158  &  wire180  &  wire375 ) | ( wire158  &  wire152  &  wire375 ) ;
 assign wire33001 = ( wire3859 ) | ( wire33000 ) | ( wire250  &  wire375 ) ;
 assign wire33003 = ( wire3741 ) | ( wire440  &  wire32990 ) ;
 assign wire33004 = ( wire221  &  wire32992 ) | ( pi17  &  (~ pi16)  &  wire221 ) ;
 assign wire33007 = ( wire3736 ) | ( wire3737 ) | ( wire33003 ) | ( wire33004 ) ;
 assign wire33008 = ( wire33007 ) | ( wire374  &  wire32982 ) | ( wire3955  &  wire32982 ) ;
 assign wire33010 = ( wire3744 ) | ( wire374  &  wire32994 ) | ( wire3975  &  wire32994 ) ;
 assign wire33011 = ( wire3735 ) | ( wire3739 ) | ( wire33008 ) ;
 assign wire33013 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33014 = ( pi27  &  wire189  &  wire33013 ) | ( (~ pi26)  &  wire189  &  wire33013 ) ;
 assign wire33015 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33016 = ( (~ pi27)  &  pi26  &  wire189  &  wire33015 ) ;
 assign wire33017 = ( (~ pi17)  &  pi16  &  wire155  &  wire179 ) ;
 assign wire33018 = ( (~ pi17)  &  pi16  &  (~ wire155)  &  wire179 ) ;
 assign wire33019 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33020 = ( (~ pi20)  &  (~ ni29)  &  wire153 ) | ( (~ pi20)  &  (~ n_n8352)  &  wire153 ) ;
 assign wire33021 = ( pi20  &  (~ ni29)  &  wire153 ) | ( pi20  &  (~ n_n8352)  &  wire153 ) ;
 assign wire33022 = ( wire4044 ) | ( wire4779  &  wire33020 ) | ( wire31895  &  wire33020 ) ;
 assign wire33023 = ( (~ pi27)  &  pi26  &  pi16 ) ;
 assign wire33024 = ( pi27  &  pi16 ) | ( (~ pi26)  &  pi16 ) ;
 assign wire33026 = ( (~ ni29)  &  wire180  &  wire154 ) | ( wire180  &  (~ n_n8352)  &  wire154 ) ;
 assign wire33027 = ( (~ ni29)  &  wire178  &  wire154 ) | ( wire178  &  (~ n_n8352)  &  wire154 ) ;
 assign wire33028 = ( (~ ni29)  &  wire152  &  wire154 ) | ( wire152  &  (~ n_n8352)  &  wire154 ) ;
 assign wire33029 = ( wire244  &  wire375 ) | ( n_n7808  &  wire33028 ) ;
 assign wire33030 = ( wire178  &  wire154  &  wire375 ) | ( wire152  &  wire154  &  wire375 ) ;
 assign wire33032 = ( wire33029 ) | ( wire33030 ) | ( n_n7816  &  wire33026 ) ;
 assign wire33034 = ( wire3752 ) | ( wire3755 ) | ( wire154  &  wire221 ) ;
 assign wire33035 = ( wire33034 ) | ( wire4043  &  wire33023 ) | ( wire33022  &  wire33023 ) ;
 assign wire33036 = ( wire3748 ) | ( wire4046  &  wire33024 ) | ( wire31899  &  wire33024 ) ;
 assign wire33040 = ( wire3749 ) | ( wire3750 ) | ( wire3751 ) | ( wire33035 ) ;
 assign wire33043 = ( wire3712 ) | ( wire3715 ) | ( wire221  &  wire32950 ) ;
 assign wire33044 = ( wire33043 ) | ( wire4005  &  wire32936 ) | ( wire32934  &  wire32936 ) ;
 assign wire33045 = ( wire3709 ) | ( wire3708 ) ;
 assign wire33046 = ( wire3711 ) | ( wire3710 ) ;
 assign wire33047 = ( wire33044 ) | ( wire535  &  wire32938 ) ;
 assign wire33050 = ( wire3717 ) | ( wire33045 ) | ( wire33046 ) | ( wire33047 ) ;
 assign wire33052 = ( wire3716 ) | ( wire33050 ) | ( wire1016  &  n_n6828 ) ;
 assign wire33055 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire33056 = ( pi27  &  wire213  &  wire33055 ) | ( pi26  &  wire213  &  wire33055 ) ;
 assign wire33057 = ( pi15  &  wire377  &  wire33056 ) ;
 assign wire33058 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire33059 = ( (~ pi27)  &  (~ pi26)  &  wire213  &  wire33058 ) ;
 assign wire33060 = ( pi15  &  wire377  &  wire33059 ) ;
 assign wire33062 = ( (~ pi16)  &  pi15  &  wire377  &  wire1102 ) ;
 assign wire33064 = ( (~ pi16)  &  pi15  &  wire377  &  wire1096 ) ;
 assign wire33065 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire33066 = ( pi15  &  wire377  &  wire33065 ) ;
 assign wire33067 = ( (~ pi27)  &  (~ pi26)  &  (~ pi16) ) ;
 assign wire33068 = ( pi15  &  wire377  &  wire33067 ) ;
 assign wire33069 = ( pi27  &  (~ pi16) ) | ( pi26  &  (~ pi16) ) ;
 assign wire33070 = ( pi15  &  wire377  &  wire33069 ) ;
 assign wire33071 = ( (~ pi16)  &  pi15  &  wire377 ) ;
 assign wire33072 = ( pi27  &  pi15  &  wire377 ) | ( pi26  &  pi15  &  wire377 ) ;
 assign wire33073 = ( (~ pi27)  &  (~ pi26)  &  pi15  &  wire377 ) ;
 assign wire33074 = ( pi17  &  (~ pi16)  &  pi15  &  wire377 ) ;
 assign wire33075 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33076 = ( pi27  &  wire213  &  wire33075 ) | ( pi26  &  wire213  &  wire33075 ) ;
 assign wire33077 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33078 = ( (~ pi27)  &  (~ pi26)  &  wire213  &  wire33077 ) ;
 assign wire33079 = ( (~ pi17)  &  pi16  &  (~ wire156)  &  wire182 ) ;
 assign wire33080 = ( (~ pi17)  &  pi16  &  wire156  &  wire182 ) ;
 assign wire33081 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33082 = ( (~ pi27)  &  (~ pi26)  &  pi16 ) ;
 assign wire33083 = ( pi27  &  pi16 ) | ( pi26  &  pi16 ) ;
 assign wire33085 = ( wire3805 ) | ( wire3808 ) | ( wire154  &  wire227 ) ;
 assign wire33086 = ( wire33085 ) | ( wire4043  &  wire33082 ) | ( wire33022  &  wire33082 ) ;
 assign wire33087 = ( wire3801 ) | ( wire4046  &  wire33083 ) | ( wire31899  &  wire33083 ) ;
 assign wire33091 = ( wire3802 ) | ( wire3803 ) | ( wire3804 ) | ( wire33086 ) ;
 assign wire33093 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33094 = ( pi27  &  wire213  &  wire33093 ) | ( pi26  &  wire213  &  wire33093 ) ;
 assign wire33095 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33096 = ( (~ pi27)  &  (~ pi26)  &  wire213  &  wire33095 ) ;
 assign wire33097 = ( (~ pi17)  &  pi16  &  (~ wire156)  &  wire182 ) ;
 assign wire33098 = ( (~ pi17)  &  pi16  &  wire156  &  wire182 ) ;
 assign wire33099 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33100 = ( (~ pi27)  &  (~ pi26)  &  pi16 ) ;
 assign wire33101 = ( pi27  &  pi16 ) | ( pi26  &  pi16 ) ;
 assign wire33103 = ( wire3816 ) | ( wire3819 ) | ( wire154  &  wire227 ) ;
 assign wire33105 = ( wire3817 ) | ( wire3818 ) | ( wire33103 ) ;
 assign wire33106 = ( wire33105 ) | ( wire374  &  wire33094 ) | ( wire3969  &  wire33094 ) ;
 assign wire33108 = ( wire3821 ) | ( wire374  &  wire33098 ) | ( wire3963  &  wire33098 ) ;
 assign wire33109 = ( wire3813 ) | ( wire3814 ) | ( wire33106 ) ;
 assign wire33111 = ( pi27  &  (~ pi16) ) | ( pi26  &  (~ pi16) ) ;
 assign wire33112 = ( (~ pi27)  &  (~ pi26)  &  (~ pi16) ) ;
 assign wire33113 = ( (~ pi27)  &  (~ pi26)  &  wire189  &  wire698 ) ;
 assign wire33114 = ( (~ pi17)  &  (~ pi16)  &  wire156  &  wire179 ) ;
 assign wire33115 = ( pi27  &  wire189  &  wire698 ) | ( pi26  &  wire189  &  wire698 ) ;
 assign wire33116 = ( (~ pi17)  &  (~ pi16)  &  (~ wire156)  &  wire179 ) ;
 assign wire33117 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire33119 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire33120 = ( wire3849 ) | ( wire442  &  wire33117 ) ;
 assign wire33121 = ( wire227  &  wire33119 ) | ( pi17  &  (~ pi16)  &  wire227 ) ;
 assign wire33124 = ( wire3842 ) | ( wire3843 ) | ( wire33120 ) | ( wire33121 ) ;
 assign wire33125 = ( wire33124 ) | ( wire375  &  wire33113 ) | ( wire3868  &  wire33113 ) ;
 assign wire33127 = ( wire3852 ) | ( wire375  &  wire33116 ) | ( wire3870  &  wire33116 ) ;
 assign wire33128 = ( wire3845 ) | ( wire3846 ) | ( wire33125 ) ;
 assign wire33130 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire179 ) ;
 assign wire33131 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire179 ) ;
 assign wire33132 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire182 ) ;
 assign wire33133 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire182 ) ;
 assign wire33134 = ( (~ pi16)  &  pi27 ) ;
 assign wire33136 = ( pi17  &  (~ pi16)  &  wire201 ) | ( (~ pi17)  &  (~ pi16)  &  wire201 ) ;
 assign wire33137 = ( wire33136 ) | ( wire4005  &  wire33134 ) | ( wire32934  &  wire33134 ) ;
 assign wire33138 = ( wire3980 ) | ( wire3979 ) ;
 assign wire33139 = ( wire3982 ) | ( wire3981 ) ;
 assign wire33140 = ( wire33137 ) | ( (~ pi27)  &  (~ pi16)  &  wire535 ) ;
 assign wire33143 = ( wire3987 ) | ( wire33138 ) | ( wire33139 ) | ( wire33140 ) ;
 assign wire33144 = ( (~ pi17)  &  pi27  &  pi16  &  wire179 ) ;
 assign wire33145 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire179 ) ;
 assign wire33146 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire182 ) ;
 assign wire33147 = ( (~ pi17)  &  pi27  &  pi16  &  wire182 ) ;
 assign wire33148 = ( pi16  &  pi27 ) ;
 assign wire33149 = ( pi16  &  (~ pi27) ) ;
 assign wire33150 = ( pi17  &  pi16  &  wire201 ) | ( (~ pi17)  &  pi16  &  wire201 ) ;
 assign wire33151 = ( wire33150 ) | ( wire4043  &  wire33148 ) | ( wire33022  &  wire33148 ) ;
 assign wire33152 = ( wire4017 ) | ( wire4046  &  wire33149 ) | ( wire31899  &  wire33149 ) ;
 assign wire33156 = ( wire4018 ) | ( wire4019 ) | ( wire4020 ) | ( wire33151 ) ;
 assign wire33158 = ( (~ pi17)  &  pi27  &  pi16  &  wire179 ) ;
 assign wire33159 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire179 ) ;
 assign wire33160 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire182 ) ;
 assign wire33161 = ( (~ pi17)  &  pi27  &  pi16  &  wire182 ) ;
 assign wire33162 = ( pi16  &  pi27 ) ;
 assign wire33163 = ( pi16  &  (~ pi27) ) ;
 assign wire33164 = ( pi17  &  pi16  &  wire201 ) | ( (~ pi17)  &  pi16  &  wire201 ) ;
 assign wire33166 = ( wire3785 ) | ( wire3786 ) | ( wire33164 ) ;
 assign wire33167 = ( wire33166 ) | ( wire375  &  wire33158 ) | ( wire3840  &  wire33158 ) ;
 assign wire33169 = ( wire3789 ) | ( wire375  &  wire33161 ) | ( wire3838  &  wire33161 ) ;
 assign wire33170 = ( wire3782 ) | ( wire3783 ) | ( wire33167 ) ;
 assign wire33172 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire179 ) ;
 assign wire33173 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire179 ) ;
 assign wire33174 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire182 ) ;
 assign wire33175 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire182 ) ;
 assign wire33177 = ( (~ pi16)  &  pi27 ) ;
 assign wire33178 = ( pi17  &  (~ pi16)  &  wire201 ) | ( (~ pi17)  &  (~ pi16)  &  wire201 ) ;
 assign wire33180 = ( wire3795 ) | ( wire3796 ) | ( wire33178 ) ;
 assign wire33181 = ( wire33180 ) | ( wire375  &  wire33172 ) | ( wire3870  &  wire33172 ) ;
 assign wire33183 = ( wire3799 ) | ( wire375  &  wire33175 ) | ( wire3868  &  wire33175 ) ;
 assign wire33184 = ( wire3792 ) | ( wire3793 ) | ( wire33181 ) ;
 assign wire33187 = ( wire3765 ) | ( wire3768 ) | ( wire227  &  wire33074 ) ;
 assign wire33188 = ( wire33187 ) | ( wire4005  &  wire33068 ) | ( wire32934  &  wire33068 ) ;
 assign wire33189 = ( wire3762 ) | ( wire3761 ) ;
 assign wire33190 = ( wire3764 ) | ( wire3763 ) ;
 assign wire33191 = ( wire33188 ) | ( wire535  &  wire33070 ) ;
 assign wire33194 = ( wire3770 ) | ( wire33189 ) | ( wire33190 ) | ( wire33191 ) ;
 assign wire33196 = ( wire3769 ) | ( wire33194 ) | ( wire1083  &  n_n7239 ) ;
 assign wire33197 = ( wire848  &  n_n7001 ) | ( wire848  &  wire3986 ) | ( wire848  &  wire33143 ) ;
 assign wire33198 = ( wire33197 ) | ( wire33196 ) ;
 assign wire33201 = ( wire3779 ) | ( wire3778 ) ;
 assign wire33202 = ( wire3773 ) | ( wire3774 ) | ( wire3777 ) | ( wire33198 ) ;
 assign wire33206 = ( wire4090  &  wire32608 ) | ( wire32587  &  wire32608 ) | ( wire4090  &  wire32611 ) | ( wire32587  &  wire32611 ) ;
 assign wire33209 = ( wire3651 ) | ( wire3658 ) | ( wire3664 ) ;
 assign wire33210 = ( wire3653 ) | ( wire3660 ) | ( wire3662 ) | ( wire33206 ) ;
 assign wire33212 = ( wire3655 ) | ( wire3661 ) | ( wire33209 ) | ( wire33210 ) ;
 assign wire33214 = ( wire3652 ) | ( wire1290  &  wire32602 ) ;
 assign wire33215 = ( wire3650 ) | ( wire33212 ) | ( wire1292  &  wire32616 ) ;
 assign wire33218 = ( wire3663 ) | ( wire3665 ) | ( wire33214 ) | ( wire33215 ) ;
 assign wire33220 = ( wire3666 ) | ( wire33218 ) | ( n_n7400  &  (~ wire793) ) ;
 assign wire33223 = ( wire684  &  wire32188 ) | ( nv6124  &  wire32202 ) ;
 assign wire33225 = ( wire4269  &  wire32193 ) | ( wire32189  &  wire32193 ) | ( wire4269  &  wire32196 ) | ( wire32189  &  wire32196 ) ;
 assign wire33226 = ( wire3533 ) | ( wire33223 ) | ( wire684  &  wire32199 ) ;
 assign wire33227 = ( nv5862  &  wire32352 ) | ( nv6146  &  wire32354 ) ;
 assign wire33228 = ( wire33225 ) | ( nv6146  &  wire32486 ) ;
 assign wire33230 = ( wire352  &  wire32219 ) | ( wire352  &  wire32221 ) ;
 assign wire33234 = ( wire3529 ) | ( wire3534 ) | ( wire33227 ) | ( wire33228 ) ;
 assign wire33235 = ( wire3528 ) | ( wire33226 ) | ( wire33230 ) | ( wire33234 ) ;
 assign wire33236 = ( wire33235 ) | ( wire1256  &  wire1328  &  wire32335 ) ;
 assign wire33238 = ( nv5843  &  wire32490 ) | ( nv5843  &  wire32581 ) ;
 assign wire33240 = ( wire3537 ) | ( wire3540 ) | ( wire33236 ) | ( wire33238 ) ;
 assign wire33241 = ( (~ ni2)  &  (~ ni3)  &  wire281 ) ;
 assign wire33242 = ( wire3522 ) | ( wire170  &  wire32139 ) | ( wire1118  &  wire32139 ) ;
 assign wire33244 = ( wire3515 ) | ( wire3517 ) | ( wire33242 ) ;
 assign wire33246 = ( wire33244 ) | ( n_n8104  &  wire32138 ) ;
 assign wire33249 = ( (~ ni2)  &  (~ ni3)  &  ni9  &  ni10 ) ;
 assign wire33251 = ( (~ ni38)  &  (~ ni2)  &  ni37  &  (~ ni3) ) ;
 assign wire33252 = ( (~ pi21)  &  (~ ni2)  &  (~ ni3) ) | ( (~ pi22)  &  (~ ni2)  &  (~ ni3) ) ;
 assign wire33254 = ( pi21  &  ni31 ) | ( ni2  &  ni31 ) | ( ni3  &  ni31 ) ;
 assign wire33256 = ( wire33254 ) | ( n_n13895  &  nv6428  &  nv633 ) ;
 assign wire33257 = ( (~ ni2)  &  (~ ni3)  &  ni9  &  ni10 ) ;
 assign wire33258 = ( (~ ni9)  &  wire33257 ) | ( (~ ni10)  &  wire33257 ) | ( (~ ni8)  &  wire33257 ) ;
 assign wire33260 = ( (~ ni2)  &  (~ ni3)  &  ni8  &  wire1165 ) ;
 assign wire33261 = ( (~ ni2)  &  (~ ni3)  &  (~ ni7) ) ;
 assign wire33262 = ( wire3506 ) | ( (~ wire31161)  &  (~ wire31162)  &  wire33258 ) ;
 assign wire33263 = ( (~ wire31161)  &  (~ wire31162)  &  wire33260 ) | ( (~ wire31161)  &  (~ wire31162)  &  wire33261 ) ;
 assign wire33266 = ( (~ ni33)  &  (~ ni32)  &  (~ ni31)  &  ni29 ) ;
 assign wire33267 = ( (~ ni39)  &  (~ ni36) ) | ( ni38  &  (~ ni36) ) | ( ni37  &  (~ ni36) ) ;
 assign wire33270 = ( (~ wire1081)  &  (~ wire463)  &  (~ wire3297) ) ;
 assign wire33272 = ( (~ wire1081)  &  wire707 ) | ( (~ wire1081)  &  wire3301 ) | ( (~ wire1081)  &  wire3303 ) ;
 assign wire33274 = ( ni37 ) | ( (~ wire3462)  &  (~ wire33267) ) ;
 assign wire33276 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire1081) ) ;
 assign wire33278 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire1081) ) ;
 assign wire33279 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33282 = ( (~ wire827)  &  (~ wire1047)  &  (~ nv6472) ) ;
 assign wire33284 = ( (~ wire827)  &  (~ wire1047)  &  (~ nv6472) ) ;
 assign wire33288 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire6766) ) ;
 assign wire33290 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire6766) ) ;
 assign wire33291 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33293 = ( ni35 ) | ( (~ wire827)  &  (~ wire1081)  &  wire33279 ) ;
 assign wire33294 = ( wire3295 ) | ( (~ ni37)  &  (~ wire827)  &  wire33274 ) ;
 assign wire33295 = ( (~ wire797)  &  wire33276 ) | ( n_n5729  &  wire33278 ) ;
 assign wire33296 = ( (~ wire797)  &  wire33282 ) | ( n_n5729  &  wire33284 ) ;
 assign wire33297 = ( wire3292 ) | ( (~ wire463)  &  (~ wire3297)  &  wire33288 ) ;
 assign wire33298 = ( wire33293 ) | ( n_n5729  &  wire33290 ) ;
 assign wire33299 = ( (~ wire827)  &  (~ wire1047)  &  wire33270 ) | ( (~ wire827)  &  (~ wire1047)  &  wire33272 ) ;
 assign wire33302 = ( wire33293 ) | ( wire33299 ) | ( n_n5729  &  wire33290 ) ;
 assign wire33303 = ( wire33294 ) | ( wire33295 ) | ( wire33296 ) | ( wire33297 ) ;
 assign wire33304 = ( wire417  &  (~ wire707)  &  (~ wire3301)  &  (~ wire3303) ) ;
 assign wire33305 = ( (~ wire157)  &  (~ wire463)  &  (~ wire3297) ) ;
 assign wire33306 = ( (~ ni36)  &  (~ ni35)  &  (~ wire157) ) ;
 assign wire33307 = ( (~ n_n5729)  &  wire33298 ) | ( (~ n_n5729)  &  wire33299 ) | ( (~ n_n5729)  &  wire33303 ) ;
 assign wire33309 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire178 ) ;
 assign wire33310 = ( ni39  &  (~ ni36) ) | ( ni38  &  (~ ni36) ) | ( ni37  &  (~ ni36) ) ;
 assign wire33319 = ( (~ nv6486)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33321 = ( (~ nv6486)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33325 = ( wire426  &  (~ nv669)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33327 = ( wire426  &  (~ nv669)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33328 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33331 = ( wire426  &  (~ nv669)  &  (~ nv6486)  &  (~ wire826) ) ;
 assign wire33333 = ( wire426  &  (~ nv669)  &  (~ nv6486)  &  (~ wire826) ) ;
 assign wire33334 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33336 = ( ni35 ) | ( (~ wire826)  &  (~ wire1068)  &  wire33328 ) ;
 assign wire33339 = ( (~ wire826)  &  (~ wire798)  &  (~ wire592) ) | ( (~ wire826)  &  n_n5713  &  (~ wire592) ) ;
 assign wire33340 = ( (~ wire798)  &  wire33319 ) | ( n_n5713  &  wire33321 ) ;
 assign wire33341 = ( (~ wire798)  &  wire33325 ) | ( n_n5713  &  wire33327 ) ;
 assign wire33342 = ( (~ wire798)  &  wire33331 ) | ( n_n5713  &  wire33333 ) ;
 assign wire33343 = ( wire3257 ) | ( wire3260 ) | ( wire3266 ) | ( wire33336 ) ;
 assign wire33345 = ( wire33342 ) | ( wire33341 ) ;
 assign wire33346 = ( wire33339 ) | ( wire33340 ) | ( wire33343 ) ;
 assign wire33347 = ( (~ n_n5713)  &  wire417 ) ;
 assign wire33348 = ( (~ wire157)  &  (~ wire253)  &  (~ wire463) ) | ( (~ wire157)  &  (~ nv6486)  &  (~ wire463) ) ;
 assign wire33349 = ( (~ ni36)  &  (~ ni35)  &  (~ wire157) ) ;
 assign wire33350 = ( (~ n_n5713)  &  wire33341 ) | ( (~ n_n5713)  &  wire33342 ) | ( (~ n_n5713)  &  wire33346 ) ;
 assign wire33352 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire180 ) ;
 assign wire33355 = ( (~ pi16)  &  (~ pi15)  &  wire272 ) ;
 assign wire33364 = ( (~ nv6589)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33366 = ( (~ nv6589)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33370 = ( (~ nv669)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33372 = ( (~ nv669)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33373 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33376 = ( (~ nv669)  &  (~ wire826)  &  (~ wire6727) ) ;
 assign wire33378 = ( (~ nv669)  &  (~ wire826)  &  (~ wire6727) ) ;
 assign wire33379 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33381 = ( ni35 ) | ( (~ wire826)  &  (~ wire1068)  &  wire33373 ) ;
 assign wire33384 = ( (~ wire800)  &  (~ wire826)  &  (~ wire592) ) | ( (~ wire826)  &  n_n5604  &  (~ wire592) ) ;
 assign wire33385 = ( (~ wire800)  &  wire33364 ) | ( n_n5604  &  wire33366 ) ;
 assign wire33386 = ( (~ wire800)  &  wire33370 ) | ( n_n5604  &  wire33372 ) ;
 assign wire33387 = ( (~ wire800)  &  wire33376 ) | ( n_n5604  &  wire33378 ) ;
 assign wire33388 = ( wire3479 ) | ( wire3482 ) | ( wire3488 ) | ( wire33381 ) ;
 assign wire33390 = ( wire33387 ) | ( wire33386 ) ;
 assign wire33391 = ( wire33384 ) | ( wire33385 ) | ( wire33388 ) ;
 assign wire33392 = ( wire417  &  (~ wire1198)  &  (~ wire3497) ) ;
 assign wire33393 = ( (~ wire157)  &  (~ wire464)  &  (~ wire3493) ) ;
 assign wire33394 = ( (~ ni36)  &  (~ ni35)  &  (~ wire157) ) ;
 assign wire33395 = ( (~ wire1198)  &  (~ wire3497)  &  wire33390 ) | ( (~ wire1198)  &  (~ wire3497)  &  wire33391 ) ;
 assign wire33398 = ( ni37 ) | ( (~ wire3462)  &  (~ wire33267) ) ;
 assign wire33400 = ( ni37 ) | ( (~ wire3462)  &  (~ wire33267) ) ;
 assign wire33404 = ( (~ wire1081)  &  (~ wire464)  &  (~ wire3464) ) ;
 assign wire33406 = ( (~ wire1081)  &  wire1198 ) | ( (~ wire1081)  &  wire3466 ) ;
 assign wire33407 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33410 = ( (~ wire1047)  &  (~ wire464)  &  (~ wire3464) ) ;
 assign wire33412 = ( (~ wire1047)  &  wire1198 ) | ( (~ wire1047)  &  wire3466 ) ;
 assign wire33413 = ( (~ ni37)  &  (~ nv669)  &  (~ wire6766) ) ;
 assign wire33415 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ wire6766) ) ;
 assign wire33417 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ wire6766) ) ;
 assign wire33420 = ( (~ ni37)  &  (~ nv669)  &  (~ wire6766) ) ;
 assign wire33421 = ( ni35 ) | ( (~ wire827)  &  wire33420 ) ;
 assign wire33426 = ( (~ nv669)  &  (~ wire827)  &  wire33404 ) | ( (~ nv669)  &  (~ wire827)  &  wire33406 ) ;
 assign wire33427 = ( (~ nv6576)  &  (~ wire827)  &  wire33410 ) | ( (~ nv6576)  &  (~ wire827)  &  wire33412 ) ;
 assign wire33428 = ( wire3453 ) | ( wire3456 ) | ( wire3457 ) | ( wire3458 ) ;
 assign wire33429 = ( wire3448 ) | ( wire3449 ) | ( wire3450 ) | ( wire33421 ) ;
 assign wire33433 = ( (~ wire157)  &  (~ wire464)  &  (~ wire3464) ) ;
 assign wire33434 = ( (~ ni36)  &  (~ ni35)  &  (~ wire157) ) ;
 assign wire33438 = ( (~ wire1081)  &  (~ wire465)  &  (~ wire3383) ) ;
 assign wire33440 = ( (~ wire1081)  &  wire707 ) | ( (~ wire1081)  &  wire3387 ) | ( (~ wire1081)  &  wire3389 ) ;
 assign wire33442 = ( ni37 ) | ( (~ wire3462)  &  (~ wire33267) ) ;
 assign wire33444 = ( (~ wire827)  &  (~ wire1081)  &  (~ nv6472) ) ;
 assign wire33446 = ( (~ wire827)  &  (~ wire1081)  &  (~ nv6472) ) ;
 assign wire33450 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire1047) ) ;
 assign wire33452 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire1047) ) ;
 assign wire33453 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33456 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire6766) ) ;
 assign wire33458 = ( wire426  &  (~ nv669)  &  (~ wire827)  &  (~ wire6766) ) ;
 assign wire33459 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33461 = ( (~ ni35) ) | ( (~ wire827)  &  (~ wire1047)  &  wire33453 ) ;
 assign wire33462 = ( wire3381 ) | ( (~ ni37)  &  (~ wire827)  &  wire33442 ) ;
 assign wire33463 = ( (~ wire801)  &  wire33444 ) | ( n_n5768  &  wire33446 ) ;
 assign wire33464 = ( wire3375 ) | ( (~ wire465)  &  (~ wire3383)  &  wire33450 ) ;
 assign wire33465 = ( n_n5768  &  wire33452 ) | ( (~ wire801)  &  wire33456 ) ;
 assign wire33466 = ( wire33461 ) | ( n_n5768  &  wire33458 ) ;
 assign wire33467 = ( (~ wire827)  &  (~ wire1047)  &  wire33438 ) | ( (~ wire827)  &  (~ wire1047)  &  wire33440 ) ;
 assign wire33470 = ( wire33461 ) | ( wire33467 ) | ( n_n5768  &  wire33458 ) ;
 assign wire33471 = ( wire33462 ) | ( wire33463 ) | ( wire33464 ) | ( wire33465 ) ;
 assign wire33472 = ( wire417  &  (~ wire707)  &  (~ wire3387)  &  (~ wire3389) ) ;
 assign wire33473 = ( (~ wire157)  &  (~ wire465)  &  (~ wire3383) ) ;
 assign wire33474 = ( (~ ni36)  &  ni35  &  (~ wire157) ) ;
 assign wire33475 = ( (~ n_n5768)  &  wire33466 ) | ( (~ n_n5768)  &  wire33467 ) | ( (~ n_n5768)  &  wire33471 ) ;
 assign wire33476 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire33484 = ( (~ nv669)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33486 = ( (~ nv669)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33487 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33490 = ( (~ nv6589)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33492 = ( (~ nv6589)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33496 = ( (~ nv669)  &  (~ wire826)  &  (~ wire6727) ) ;
 assign wire33498 = ( (~ nv669)  &  (~ wire826)  &  (~ wire6727) ) ;
 assign wire33499 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33501 = ( (~ ni35) ) | ( (~ wire826)  &  (~ wire1123)  &  wire33487 ) ;
 assign wire33504 = ( (~ wire804)  &  (~ wire826)  &  (~ wire592) ) | ( n_n5644  &  (~ wire826)  &  (~ wire592) ) ;
 assign wire33505 = ( (~ wire804)  &  wire33484 ) | ( n_n5644  &  wire33486 ) ;
 assign wire33506 = ( (~ wire804)  &  wire33490 ) | ( n_n5644  &  wire33492 ) ;
 assign wire33507 = ( (~ wire804)  &  wire33496 ) | ( n_n5644  &  wire33498 ) ;
 assign wire33508 = ( wire3420 ) | ( wire3426 ) | ( wire3429 ) | ( wire33501 ) ;
 assign wire33510 = ( wire33507 ) | ( wire33506 ) ;
 assign wire33511 = ( wire33504 ) | ( wire33505 ) | ( wire33508 ) ;
 assign wire33512 = ( wire417  &  (~ wire1200)  &  (~ wire3435) ) ;
 assign wire33513 = ( (~ wire157)  &  (~ wire468)  &  (~ wire3431) ) ;
 assign wire33514 = ( (~ ni36)  &  ni35  &  (~ wire157) ) ;
 assign wire33515 = ( (~ wire1200)  &  (~ wire3435)  &  wire33510 ) | ( (~ wire1200)  &  (~ wire3435)  &  wire33511 ) ;
 assign wire33518 = ( (~ wire1081)  &  (~ wire468)  &  (~ wire3410) ) ;
 assign wire33520 = ( (~ wire1081)  &  wire1200 ) | ( (~ wire1081)  &  wire3412 ) ;
 assign wire33524 = ( (~ wire1081)  &  (~ wire468)  &  (~ wire3410) ) ;
 assign wire33526 = ( (~ wire1081)  &  wire1200 ) | ( (~ wire1081)  &  wire3412 ) ;
 assign wire33527 = ( (~ ni37)  &  (~ nv669)  &  (~ wire6766) ) ;
 assign wire33530 = ( (~ wire1047)  &  (~ wire468)  &  (~ wire3410) ) ;
 assign wire33532 = ( (~ wire1047)  &  wire1200 ) | ( (~ wire1047)  &  wire3412 ) ;
 assign wire33533 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ ni37) ) ;
 assign wire33535 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ wire6766) ) ;
 assign wire33537 = ( (~ ni43)  &  (~ ni47)  &  (~ ni45)  &  (~ wire6766) ) ;
 assign wire33540 = ( (~ ni37)  &  (~ nv669)  &  (~ wire6766) ) ;
 assign wire33541 = ( (~ ni35) ) | ( (~ wire827)  &  wire33540 ) ;
 assign wire33544 = ( wire33541 ) | ( (~ wire827)  &  (~ wire1047)  &  wire33518 ) ;
 assign wire33545 = ( wire3399 ) | ( (~ wire827)  &  (~ wire1047)  &  wire33520 ) ;
 assign wire33546 = ( (~ nv6576)  &  (~ wire827)  &  wire33524 ) | ( (~ nv6576)  &  (~ wire827)  &  wire33526 ) ;
 assign wire33547 = ( (~ nv669)  &  (~ wire827)  &  wire33530 ) | ( (~ nv669)  &  (~ wire827)  &  wire33532 ) ;
 assign wire33548 = ( wire3402 ) | ( wire3405 ) | ( wire3406 ) | ( wire3407 ) ;
 assign wire33550 = ( wire33547 ) | ( wire33546 ) ;
 assign wire33551 = ( wire33544 ) | ( wire33545 ) | ( wire33548 ) ;
 assign wire33552 = ( wire417  &  (~ wire1200)  &  (~ wire3412) ) ;
 assign wire33553 = ( (~ wire157)  &  (~ wire468)  &  (~ wire3410) ) ;
 assign wire33554 = ( (~ ni36)  &  ni35  &  (~ wire157) ) ;
 assign wire33555 = ( (~ wire1200)  &  (~ wire3412)  &  wire33550 ) | ( (~ wire1200)  &  (~ wire3412)  &  wire33551 ) ;
 assign wire33564 = ( wire426  &  (~ nv669)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33566 = ( wire426  &  (~ nv669)  &  (~ wire826)  &  (~ wire1123) ) ;
 assign wire33567 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33570 = ( (~ nv6486)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33572 = ( (~ nv6486)  &  (~ wire826)  &  (~ wire1068) ) ;
 assign wire33576 = ( wire426  &  (~ nv669)  &  (~ nv6486)  &  (~ wire826) ) ;
 assign wire33578 = ( wire426  &  (~ nv669)  &  (~ nv6486)  &  (~ wire826) ) ;
 assign wire33579 = ( ni42  &  (~ ni37)  &  (~ nv669) ) | ( (~ ni41)  &  (~ ni37)  &  (~ nv669) ) ;
 assign wire33581 = ( (~ ni35) ) | ( (~ wire826)  &  (~ wire1123)  &  wire33567 ) ;
 assign wire33584 = ( n_n5752  &  (~ wire826)  &  (~ wire592) ) | ( (~ wire802)  &  (~ wire826)  &  (~ wire592) ) ;
 assign wire33585 = ( (~ wire802)  &  wire33564 ) | ( n_n5752  &  wire33566 ) ;
 assign wire33586 = ( (~ wire802)  &  wire33570 ) | ( n_n5752  &  wire33572 ) ;
 assign wire33587 = ( (~ wire802)  &  wire33576 ) | ( n_n5752  &  wire33578 ) ;
 assign wire33588 = ( wire3349 ) | ( wire3355 ) | ( wire3358 ) | ( wire33581 ) ;
 assign wire33590 = ( wire33587 ) | ( wire33586 ) ;
 assign wire33591 = ( wire33584 ) | ( wire33585 ) | ( wire33588 ) ;
 assign wire33592 = ( (~ n_n5752)  &  wire417 ) ;
 assign wire33593 = ( (~ wire157)  &  (~ wire254)  &  (~ wire465) ) | ( (~ wire157)  &  (~ nv6486)  &  (~ wire465) ) ;
 assign wire33594 = ( (~ ni36)  &  ni35  &  (~ wire157) ) ;
 assign wire33595 = ( (~ n_n5752)  &  wire33586 ) | ( (~ n_n5752)  &  wire33587 ) | ( (~ n_n5752)  &  wire33591 ) ;
 assign wire33596 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire33598 = ( wire426  &  (~ nv669)  &  wire1074  &  (~ wire6766) ) ;
 assign wire33599 = ( (~ wire157)  &  (~ n_n2328)  &  (~ nv6472) ) ;
 assign wire33600 = ( (~ ni47)  &  (~ ni45)  &  (~ ni38) ) ;
 assign wire33601 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire33603 = ( (~ nv6486)  &  wire1074 ) ;
 assign wire33604 = ( (~ wire157)  &  (~ n_n2328)  &  (~ nv6486) ) ;
 assign wire33605 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire33608 = ( (~ nv669)  &  wire1074  &  (~ wire6727) ) ;
 assign wire33609 = ( (~ wire157)  &  (~ n_n2328)  &  (~ nv6589) ) ;
 assign wire33611 = ( (~ nv669)  &  wire1074  &  (~ wire6766) ) ;
 assign wire33612 = ( (~ wire157)  &  (~ nv669)  &  (~ n_n2328)  &  (~ wire6766) ) ;
 assign wire33613 = ( pi17  &  (~ pi16)  &  (~ pi15)  &  wire173 ) | ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire173 ) ;
 assign wire33614 = ( pi19  &  wire173  &  wire507 ) | ( (~ pi19)  &  wire173  &  wire614 ) ;
 assign wire33616 = ( wire33613 ) | ( wire33614 ) | ( wire173  &  wire913 ) ;
 assign wire33618 = ( wire2346 ) | ( wire2360 ) | ( wire33616 ) ;
 assign wire33619 = ( wire33618 ) | ( nv7043  &  wire33601 ) ;
 assign wire33621 = ( wire2355 ) | ( wire33619 ) | ( wire258  &  wire446 ) ;
 assign wire33622 = ( wire33621 ) | ( wire196  &  wire33309 ) | ( wire2502  &  wire33309 ) ;
 assign wire33627 = ( wire2345 ) | ( wire2349 ) | ( wire2350 ) | ( wire2352 ) ;
 assign wire33628 = ( wire2348 ) | ( wire2351 ) | ( wire2353 ) | ( wire33622 ) ;
 assign wire33630 = ( pi17  &  (~ pi16)  &  pi15  &  wire178 ) ;
 assign wire33632 = ( pi17  &  (~ pi16)  &  pi15  &  wire180 ) ;
 assign wire33634 = ( (~ pi16)  &  pi15  &  wire272 ) ;
 assign wire33636 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire179 ) ;
 assign wire33637 = ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire182 ) ;
 assign wire33638 = ( pi17  &  pi16  &  pi15  &  wire180 ) ;
 assign wire33640 = ( (~ pi17)  &  pi16  &  pi15  &  wire182 ) ;
 assign wire33641 = ( (~ pi17)  &  pi16  &  pi15  &  wire179 ) ;
 assign wire33642 = ( (~ pi20)  &  (~ pi16)  &  pi15  &  wire153 ) ;
 assign wire33643 = ( pi20  &  (~ pi16)  &  pi15  &  wire153 ) ;
 assign wire33644 = ( pi17  &  (~ pi16)  &  pi15  &  wire173 ) | ( (~ pi17)  &  (~ pi16)  &  pi15  &  wire173 ) ;
 assign wire33645 = ( pi19  &  wire395  &  wire173 ) | ( (~ pi19)  &  wire403  &  wire173 ) ;
 assign wire33647 = ( wire33644 ) | ( wire33645 ) | ( wire173  &  wire915 ) ;
 assign wire33649 = ( wire2327 ) | ( wire2342 ) | ( wire33647 ) ;
 assign wire33651 = ( wire2335 ) | ( wire2336 ) | ( wire33649 ) ;
 assign wire33657 = ( wire2325 ) | ( wire2333 ) | ( wire2341 ) | ( wire33651 ) ;
 assign wire33658 = ( wire2326 ) | ( wire2329 ) | ( wire2332 ) | ( wire2334 ) ;
 assign wire33660 = ( wire2330 ) | ( wire2331 ) | ( wire33657 ) | ( wire33658 ) ;
 assign wire33661 = ( ni11  &  (~ ni9)  &  ni10 ) | ( ni12  &  (~ ni9)  &  ni10 ) ;
 assign wire33662 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire33661 ) ;
 assign wire33663 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire33665 = ( (~ wire175)  &  wire182  &  wire33663 ) ;
 assign wire33666 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire33668 = ( (~ wire175)  &  wire179  &  wire33666 ) ;
 assign wire33669 = ( (~ pi17)  &  (~ pi16)  &  pi15 ) ;
 assign wire33672 = ( (~ wire175)  &  wire395  &  wire182 ) ;
 assign wire33674 = ( (~ wire175)  &  wire395  &  wire179 ) ;
 assign wire33677 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire33678 = ( (~ pi20)  &  (~ pi16)  &  wire153  &  wire33677 ) ;
 assign wire33679 = ( pi15  &  (~ ni13)  &  ni14  &  (~ ni12) ) ;
 assign wire33680 = ( pi20  &  (~ pi16)  &  wire153  &  wire33679 ) ;
 assign wire33681 = ( wire3116 ) | ( wire272  &  wire3276 ) | ( wire272  &  wire3277 ) ;
 assign wire33682 = ( wire33681 ) | ( pi17  &  wire178  &  n_n4489 ) ;
 assign wire33684 = ( (~ pi16)  &  pi15  &  (~ wire175) ) ;
 assign wire33685 = ( (~ pi20)  &  (~ wire175)  &  wire226  &  wire153 ) ;
 assign wire33686 = ( pi20  &  (~ wire175)  &  wire226  &  wire153 ) ;
 assign wire33688 = ( (~ ni13)  &  ni14  &  (~ ni12)  &  ni30 ) ;
 assign wire33689 = ( pi15  &  (~ wire175)  &  wire152  &  wire154 ) ;
 assign wire33691 = ( pi17  &  pi16  &  pi15  &  (~ wire175) ) ;
 assign wire33693 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire182 ) ;
 assign wire33695 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15)  &  wire179 ) ;
 assign wire33696 = ( (~ pi17)  &  (~ pi16)  &  (~ pi15) ) ;
 assign wire33697 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire182 ) ;
 assign wire33698 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire179 ) ;
 assign wire33699 = ( ni30  &  (~ pi15) ) ;
 assign wire33700 = ( (~ pi20)  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire33701 = ( pi20  &  (~ pi16)  &  (~ pi15)  &  wire153 ) ;
 assign wire33702 = ( pi17  &  ni30 ) | ( wire272  &  n_n4611 ) ;
 assign wire33704 = ( (~ pi15)  &  (~ pi16) ) ;
 assign wire33705 = ( wire3066 ) | ( wire178  &  wire3185 ) | ( wire178  &  wire3186 ) ;
 assign wire33706 = ( wire1091  &  wire33696 ) | ( wire344  &  wire33699 ) ;
 assign wire33709 = ( wire2321 ) | ( wire2322 ) | ( wire2324 ) | ( wire33706 ) ;
 assign wire33710 = ( wire33709 ) | ( wire3326  &  wire33700 ) | ( wire3327  &  wire33700 ) ;
 assign wire33713 = ( wire2317 ) | ( wire2319 ) | ( wire2320 ) | ( wire33710 ) ;
 assign wire33715 = ( wire2310 ) | ( wire2314 ) ;
 assign wire33716 = ( wire2311 ) | ( wire2313 ) | ( wire33713 ) ;
 assign wire33721 = ( wire2295 ) | ( wire2298 ) | ( wire2304 ) | ( wire2305 ) ;
 assign wire33724 = ( wire2302 ) | ( wire2300 ) ;
 assign wire33725 = ( wire2299 ) | ( wire2303 ) | ( wire2306 ) | ( wire33721 ) ;
 assign wire33727 = ( wire33724 ) | ( wire33725 ) | ( n_n4509  &  wire33668 ) ;
 assign wire33728 = ( n_n4501  &  wire33665 ) | ( n_n4441  &  wire33674 ) ;
 assign wire33730 = ( wire33727 ) | ( wire33728 ) | ( n_n4433  &  wire33672 ) ;
 assign wire33732 = ( wire2301 ) | ( wire33730 ) | ( n_n4834  &  wire33691 ) ;
 assign wire33733 = ( wire33732 ) | ( (~ wire175)  &  n_n4934 ) ;
 assign wire33734 = ( (~ ni11)  &  (~ ni9)  &  ni10 ) ;
 assign wire33735 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire33734 ) ;
 assign wire33736 = ( pi17  &  pi21  &  pi22  &  pi16 ) ;
 assign wire33737 = ( (~ pi17)  &  pi19  &  pi16  &  (~ pi15) ) ;
 assign wire33738 = ( wire33737  &  wire611 ) ;
 assign wire33739 = ( (~ pi17)  &  pi19  &  pi16  &  pi15 ) ;
 assign wire33740 = ( wire33739  &  wire611 ) ;
 assign wire33741 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  pi15 ) ;
 assign wire33742 = ( wire33741  &  wire611 ) ;
 assign wire33743 = ( (~ pi16)  &  pi15 ) ;
 assign wire33744 = ( (~ pi17)  &  pi25  &  wire179  &  wire33743 ) ;
 assign wire33745 = ( pi15  &  wire3086 ) | ( pi25  &  (~ pi16)  &  pi15 ) ;
 assign wire33746 = ( (~ pi17)  &  pi19  &  pi15 ) ;
 assign wire33748 = ( wire1110  &  pi15 ) ;
 assign wire33750 = ( wire371 ) | ( (~ pi17)  &  wire179  &  n_n5481 ) ;
 assign wire33751 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire213 ) ;
 assign wire33753 = ( wire1110  &  n_n5481 ) | ( wire484  &  n_n5481 ) | ( n_n5481  &  wire33751 ) ;
 assign wire33754 = ( wire33753 ) | ( wire3074 ) ;
 assign wire33755 = ( wire33754 ) | ( (~ pi16)  &  wire3096 ) | ( (~ pi16)  &  wire3097 ) ;
 assign wire33756 = ( wire33755 ) | ( wire698  &  wire3092 ) | ( wire698  &  wire3093 ) ;
 assign wire33758 = ( wire585 ) | ( n_n5481  &  wire33736 ) | ( n_n5481  &  wire33748 ) ;
 assign wire33759 = ( wire3048 ) | ( wire3041 ) ;
 assign wire33760 = ( wire33758 ) | ( wire258  &  wire754 ) | ( wire258  &  wire33750 ) ;
 assign wire33763 = ( wire3042 ) | ( wire3045 ) | ( wire33759 ) | ( wire33760 ) ;
 assign wire33764 = ( wire33763 ) | ( n_n4509  &  wire33744 ) ;
 assign wire33765 = ( n_n4433  &  wire33740 ) | ( n_n4501  &  wire33742 ) ;
 assign wire33769 = ( wire3036 ) | ( wire3046 ) | ( wire33765 ) ;
 assign wire33770 = ( wire3040 ) | ( wire3050 ) | ( wire3051 ) | ( wire33764 ) ;
 assign wire33773 = ( ni11  &  (~ ni9)  &  (~ ni10) ) | ( ni12  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33774 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire33773 ) ;
 assign wire33776 = ( ni33  &  (~ ni32)  &  (~ ni31)  &  ni29 ) ;
 assign wire33777 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire33779 = ( wire370  &  wire1053  &  wire33777 ) ;
 assign wire33780 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33782 = ( wire369  &  wire1028  &  wire33780 ) ;
 assign wire33783 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33785 = ( wire369  &  wire611  &  wire33783 ) ;
 assign wire33786 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33789 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire370 ) ;
 assign wire33793 = ( (~ pi25)  &  pi16  &  wire369 ) ;
 assign wire33795 = ( (~ pi25)  &  wire152  &  wire154  &  wire369 ) ;
 assign wire33796 = ( wire1034 ) | ( wire178  &  wire197 ) | ( wire178  &  wire3444 ) ;
 assign wire33797 = ( pi17  &  (~ pi25)  &  pi16 ) ;
 assign wire33799 = ( wire369  &  pi16 ) ;
 assign wire33801 = ( wire3247 ) | ( wire1035 ) ;
 assign wire33802 = ( wire33801 ) | ( wire197  &  wire460 ) | ( wire460  &  wire3278 ) ;
 assign wire33803 = ( (~ pi25)  &  (~ pi16)  &  wire370 ) ;
 assign wire33804 = ( wire370  &  (~ pi16) ) ;
 assign wire33805 = ( pi25  &  (~ pi16)  &  wire370 ) ;
 assign wire33806 = ( wire370  &  (~ pi16) ) ;
 assign wire33807 = ( wire369  &  pi16 ) ;
 assign wire33809 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33812 = ( (~ pi17)  &  pi19  &  pi16  &  wire611 ) ;
 assign wire33813 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire33817 = ( wire3182 ) | ( pi17  &  pi16  &  wire1034 ) ;
 assign wire33818 = ( wire33817 ) | ( wire178  &  wire154  &  nv6886 ) ;
 assign wire33821 = ( wire585 ) | ( wire2715 ) | ( wire2719 ) | ( wire2720 ) ;
 assign wire33824 = ( wire2713 ) | ( wire2714 ) | ( wire2717 ) | ( wire33821 ) ;
 assign wire33825 = ( wire1206 ) | ( (~ pi25)  &  pi16  &  wire501 ) ;
 assign wire33827 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire33828 = ( (~ pi17)  &  pi19  &  (~ pi16)  &  wire1053 ) ;
 assign wire33830 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire33831 = ( wire3223 ) | ( wire1035 ) ;
 assign wire33833 = ( wire2962 ) | ( wire197  &  wire169 ) | ( wire169  &  wire3328 ) ;
 assign wire33834 = ( wire2723 ) | ( (~ pi16)  &  wire3090 ) | ( (~ pi16)  &  wire3091 ) ;
 assign wire33835 = ( wire33834 ) | ( wire2729 ) ;
 assign wire33836 = ( wire33835 ) | ( (~ pi16)  &  wire3111 ) | ( (~ pi16)  &  wire3112 ) ;
 assign wire33837 = ( wire33836 ) | ( n_n4509  &  wire387  &  wire698 ) ;
 assign wire33839 = ( wire2724 ) | ( wire33837 ) | ( n_n4501  &  wire33830 ) ;
 assign wire33842 = ( wire2694 ) | ( wire2710 ) ;
 assign wire33844 = ( wire2706 ) | ( wire2705 ) ;
 assign wire33846 = ( wire2698 ) | ( wire2707 ) | ( wire33842 ) | ( wire33844 ) ;
 assign wire33847 = ( wire33846 ) | ( wire3096  &  wire33804 ) | ( wire3097  &  wire33804 ) ;
 assign wire33848 = ( wire33847 ) | ( n_n4433  &  wire33785 ) ;
 assign wire33850 = ( wire2692 ) | ( wire2700 ) | ( wire33848 ) ;
 assign wire33855 = ( wire2691 ) | ( wire2695 ) | ( wire2697 ) | ( wire33850 ) ;
 assign wire33856 = ( wire2699 ) | ( wire2701 ) | ( wire2704 ) | ( wire2708 ) ;
 assign wire33858 = ( wire33856 ) | ( wire3246  &  wire33803 ) | ( wire33802  &  wire33803 ) ;
 assign wire33859 = ( wire2696 ) | ( wire33855 ) | ( wire369  &  n_n5328 ) ;
 assign wire33860 = ( wire2702 ) | ( wire33856 ) | ( wire33859 ) ;
 assign wire33861 = ( wire2711 ) | ( nv6450  &  wire613 ) ;
 assign wire33862 = ( (~ ni11)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33863 = ( n_n13895  &  (~ wire281)  &  (~ wire202)  &  wire33862 ) ;
 assign wire33864 = ( n_n13895  &  wire265  &  wire186  &  (~ wire281) ) ;
 assign wire33866 = ( (~ wire175)  &  wire182  &  wire507 ) ;
 assign wire33868 = ( (~ wire175)  &  wire179  &  wire507 ) ;
 assign wire33870 = ( (~ wire175)  &  wire395  &  wire179 ) ;
 assign wire33872 = ( (~ wire175)  &  wire395  &  wire182 ) ;
 assign wire33875 = ( (~ pi17)  &  (~ pi16)  &  wire179  &  wire369 ) ;
 assign wire33876 = ( (~ pi17)  &  (~ pi16)  &  wire182  &  wire369 ) ;
 assign wire33880 = ( (~ pi16)  &  wire369 ) | ( (~ pi15)  &  wire369 ) ;
 assign wire33881 = ( pi20  &  (~ pi16)  &  wire369  &  wire153 ) ;
 assign wire33882 = ( pi15  &  (~ wire175)  &  wire152  &  wire154 ) ;
 assign wire33883 = ( (~ pi20)  &  (~ pi16)  &  wire369  &  wire153 ) ;
 assign wire33885 = ( wire302  &  wire173 ) | ( wire325  &  nv6789 ) ;
 assign wire33886 = ( wire33885 ) | ( wire294  &  nv6797 ) ;
 assign wire33887 = ( wire33886 ) | ( wire197  &  wire587 ) | ( wire587  &  wire3320 ) ;
 assign wire33889 = ( (~ wire175)  &  wire395  &  wire1011 ) | ( (~ wire175)  &  wire507  &  wire1011 ) ;
 assign wire33891 = ( wire3169 ) | ( wire3175 ) | ( wire33889 ) ;
 assign wire33892 = ( wire33891 ) | ( wire197  &  wire33882 ) | ( wire3233  &  wire33882 ) ;
 assign wire33893 = ( wire33892 ) | ( wire173  &  wire613 ) | ( wire1063  &  wire613 ) ;
 assign wire33896 = ( wire3167 ) | ( wire3171 ) | ( wire3173 ) | ( wire33893 ) ;
 assign wire33899 = ( wire3166 ) | ( wire3162 ) ;
 assign wire33900 = ( wire3161 ) | ( wire3165 ) | ( wire3168 ) | ( wire33896 ) ;
 assign wire33904 = ( wire3159 ) | ( wire3160 ) | ( wire33899 ) | ( wire33900 ) ;
 assign wire33906 = ( wire3170 ) | ( wire3174 ) | ( wire3176 ) | ( wire33904 ) ;
 assign wire33907 = ( (~ ni11)  &  n_n13895  &  wire265  &  (~ wire281) ) ;
 assign wire33908 = ( pi24  &  ni31  &  ni30 ) ;
 assign wire33909 = ( (~ pi27)  &  pi26  &  (~ ni7)  &  ni8 ) ;
 assign wire33910 = ( (~ pi21)  &  wire33908 ) | ( (~ pi22)  &  wire33908 ) ;
 assign wire33911 = ( (~ wire175)  &  wire264  &  wire33909 ) ;
 assign wire33914 = ( (~ pi24)  &  nv8608  &  wire155 ) | ( (~ pi24)  &  nv8608  &  (~ wire155) ) | ( (~ pi24)  &  wire155  &  n_n11282 ) ;
 assign wire33915 = ( (~ pi23)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33916 = ( (~ pi21)  &  (~ ni7)  &  ni8 ) | ( (~ pi22)  &  (~ ni7)  &  ni8 ) ;
 assign wire33918 = ( wire699  &  wire33915  &  wire33916 ) ;
 assign wire33919 = ( (~ pi23)  &  (~ pi24)  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33920 = ( pi21  &  pi22  &  (~ ni7)  &  ni8 ) ;
 assign wire33922 = ( wire699  &  wire33919  &  wire33920 ) ;
 assign wire33923 = ( pi23  &  (~ ni9)  &  (~ ni10) ) | ( pi24  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33924 = ( pi21  &  pi22  &  (~ ni7)  &  ni8 ) ;
 assign wire33926 = ( wire699  &  wire33923  &  wire33924 ) ;
 assign wire33927 = ( pi23  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33929 = ( (~ ni7)  &  ni8  &  wire699  &  wire33927 ) ;
 assign wire33930 = ( (~ pi26)  &  (~ ni7)  &  ni8 ) ;
 assign wire33931 = ( (~ pi21)  &  wire33930 ) | ( (~ pi22)  &  wire33930 ) ;
 assign wire33932 = ( (~ wire175)  &  wire264  &  wire822 ) ;
 assign wire33933 = ( pi27  &  (~ ni7)  &  ni8 ) ;
 assign wire33935 = ( (~ wire175)  &  wire264  &  wire822 ) ;
 assign wire33936 = ( (~ pi24)  &  (~ ni7)  &  ni8 ) ;
 assign wire33938 = ( (~ wire175)  &  wire264  &  (~ wire150)  &  wire33936 ) ;
 assign wire33939 = ( (~ pi21)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire33940 = ( (~ pi22)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire33941 = ( pi21  &  pi22  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire33943 = ( ni11  &  (~ ni9)  &  (~ ni10) ) ;
 assign wire33945 = ( (~ ni7)  &  ni8  &  wire401  &  wire33943 ) ;
 assign wire33946 = ( (~ pi24)  &  (~ ni7)  &  ni8 ) ;
 assign wire33947 = ( (~ wire175)  &  wire264  &  wire33946 ) ;
 assign wire33949 = ( (~ wire175)  &  wire264  &  wire331  &  wire1044 ) ;
 assign wire33952 = ( (~ ni7)  &  ni8  &  wire264  &  wire401 ) ;
 assign wire33954 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire33955 = ( pi21  &  pi22  &  pi25  &  wire33954 ) ;
 assign wire33956 = ( wire2224 ) | ( pi21  &  n_n3347 ) ;
 assign wire33958 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire33959 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire33960 = ( pi21  &  pi22  &  pi25  &  wire33959 ) ;
 assign wire33961 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire33962 = ( pi21  &  pi22  &  pi25  &  wire33961 ) ;
 assign wire33964 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire33965 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire33966 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire33967 = ( pi17  &  pi25  &  (~ pi16)  &  wire178 ) ;
 assign wire33968 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire33971 = ( wire1352 ) | ( wire2167 ) | ( wire2173 ) ;
 assign wire33973 = ( wire2225  &  wire33965 ) | ( wire33956  &  wire33965 ) | ( wire2225  &  wire33966 ) | ( wire33956  &  wire33966 ) ;
 assign wire33976 = ( wire962 ) | ( wire2165 ) | ( wire33973 ) ;
 assign wire33977 = ( wire2174 ) | ( wire33971 ) | ( n_n4489  &  wire33967 ) ;
 assign wire33978 = ( wire2169 ) | ( wire2175 ) | ( wire33976 ) ;
 assign wire33979 = ( n_n4501  &  wire33955 ) | ( n_n4481  &  wire33960 ) ;
 assign wire33983 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire33986 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire33987 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire33989 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire33990 = ( pi21  &  pi22  &  pi25  &  wire33989 ) ;
 assign wire33992 = ( pi16  &  (~ pi17) ) ;
 assign wire33993 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire33994 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire33996 = ( wire918 ) | ( wire2152 ) | ( pi16  &  wire1320 ) ;
 assign wire33998 = ( wire2225  &  wire33993 ) | ( wire33956  &  wire33993 ) | ( wire2225  &  wire33994 ) | ( wire33956  &  wire33994 ) ;
 assign wire34001 = ( wire963 ) | ( wire2150 ) | ( wire33998 ) ;
 assign wire34002 = ( wire2154 ) | ( wire2159 ) | ( wire2160 ) | ( wire33996 ) ;
 assign wire34003 = ( wire34001 ) | ( n_n4433  &  wire181  &  wire33983 ) ;
 assign wire34005 = ( wire34002 ) | ( pi17  &  pi16  &  wire1297 ) ;
 assign wire34007 = ( wire2151 ) | ( wire2153 ) | ( wire34003 ) | ( wire34005 ) ;
 assign wire34008 = ( (~ ni7)  &  (~ ni8)  &  wire369  &  wire330 ) ;
 assign wire34010 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire34011 = ( pi21  &  pi22  &  pi25  &  wire34010 ) ;
 assign wire34013 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire34014 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34015 = ( pi21  &  pi22  &  pi25  &  wire34014 ) ;
 assign wire34016 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34017 = ( pi21  &  pi22  &  pi25  &  wire34016 ) ;
 assign wire34019 = ( pi16  &  (~ pi17) ) ;
 assign wire34020 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34021 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34022 = ( wire906 ) | ( wire2214 ) | ( wire183  &  wire276 ) ;
 assign wire34024 = ( wire2225  &  wire34020 ) | ( wire33956  &  wire34020 ) | ( wire2225  &  wire34021 ) | ( wire33956  &  wire34021 ) ;
 assign wire34027 = ( wire2200 ) | ( wire2202 ) | ( wire34022 ) ;
 assign wire34028 = ( wire2204 ) | ( wire2209 ) | ( wire34024 ) ;
 assign wire34030 = ( wire2207 ) | ( wire2210 ) | ( wire34027 ) | ( wire34028 ) ;
 assign wire34032 = ( wire2201 ) | ( (~ pi17)  &  pi16  &  wire1311 ) ;
 assign wire34033 = ( wire2199 ) | ( wire2208 ) | ( wire34030 ) ;
 assign wire34034 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire34035 = ( pi21  &  pi22  &  pi25  &  wire34034 ) ;
 assign wire34036 = ( (~ pi17)  &  (~ pi16)  &  wire182 ) ;
 assign wire34038 = ( pi21  &  pi22  &  pi25  &  wire1058 ) ;
 assign wire34039 = ( pi21  &  pi22  &  pi25  &  wire1293 ) ;
 assign wire34040 = ( (~ pi17)  &  (~ pi16)  &  wire617 ) ;
 assign wire34041 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire34042 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire34043 = ( (~ pi16)  &  ni30  &  wire155 ) | ( (~ pi16)  &  (~ wire155)  &  nv7447 ) ;
 assign wire34044 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire34045 = ( n_n3347  &  wire34040 ) | ( (~ pi16)  &  n_n3347  &  wire817 ) ;
 assign wire34046 = ( wire302  &  n_n3349 ) | ( wire247  &  wire34043 ) ;
 assign wire34048 = ( wire34045 ) | ( wire34046 ) | ( n_n4611  &  wire393 ) ;
 assign wire34050 = ( wire2193 ) | ( wire34048 ) | ( wire276  &  wire34036 ) ;
 assign wire34053 = ( wire1293  &  wire2225 ) | ( wire1058  &  wire2225 ) | ( wire1293  &  wire33956 ) | ( wire1058  &  wire33956 ) ;
 assign wire34055 = ( wire962 ) | ( wire2182 ) | ( wire2184 ) | ( wire2185 ) ;
 assign wire34057 = ( wire2191 ) | ( wire34050 ) | ( wire34053 ) | ( wire34055 ) ;
 assign wire34059 = ( wire2187 ) | ( wire2181 ) ;
 assign wire34060 = ( wire2178 ) | ( wire34057 ) | ( wire158  &  wire1326 ) ;
 assign wire34062 = ( (~ ni7)  &  (~ ni8)  &  wire370  &  wire330 ) ;
 assign wire34063 = ( nv7447 ) | ( wire192  &  n_n4509 ) ;
 assign wire34064 = ( (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34066 = ( (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34067 = ( (~ pi17)  &  (~ pi27)  &  wire179  &  wire34066 ) ;
 assign wire34068 = ( (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34069 = ( (~ pi17)  &  (~ pi27)  &  wire182  &  wire34068 ) ;
 assign wire34070 = ( nv7447 ) | ( wire192  &  n_n4501 ) ;
 assign wire34071 = ( (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34074 = ( (~ pi27)  &  (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34075 = ( ni33  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34076 = ( ni33  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34078 = ( wire2398 ) | ( wire2399 ) | ( wire2400 ) ;
 assign wire34080 = ( pi27  &  (~ pi16)  &  pi15  &  wire268 ) ;
 assign wire34082 = ( ni33  &  wire243 ) | ( (~ ni29)  &  wire243 ) | ( (~ nv6462)  &  wire243 ) ;
 assign wire34083 = ( ni33  &  wire250 ) | ( (~ ni29)  &  wire250 ) | ( (~ nv6462)  &  wire250 ) ;
 assign wire34084 = ( wire158  &  wire152  &  wire3276 ) | ( wire158  &  wire152  &  wire3277 ) ;
 assign wire34086 = ( nv7447  &  wire158  &  wire180 ) | ( nv7447  &  wire158  &  wire152 ) ;
 assign wire34088 = ( wire2386 ) | ( wire34086 ) | ( wire192  &  wire34084 ) ;
 assign wire34089 = ( wire34088 ) | ( n_n4489  &  wire34083 ) ;
 assign wire34090 = ( wire34089 ) | ( n_n4481  &  wire34082 ) ;
 assign wire34091 = ( pi27  &  pi15  &  wire268 ) ;
 assign wire34092 = ( (~ pi27)  &  pi15  &  wire268 ) ;
 assign wire34094 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34095 = ( pi27  &  wire189  &  wire34094 ) | ( pi26  &  wire189  &  wire34094 ) ;
 assign wire34096 = ( nv7447 ) | ( n_n4433  &  wire192 ) ;
 assign wire34097 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34098 = ( (~ pi27)  &  (~ pi26)  &  wire189  &  wire34097 ) ;
 assign wire34099 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34100 = ( ni33  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34101 = ( (~ pi17)  &  wire179  &  nv10153 ) ;
 assign wire34102 = ( ni33  &  wire199 ) | ( (~ ni29)  &  wire199 ) | ( (~ nv6462)  &  wire199 ) ;
 assign wire34103 = ( ni33  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34106 = ( wire2553 ) | ( wire2556 ) | ( wire2557 ) | ( wire2559 ) ;
 assign wire34108 = ( wire2558 ) | ( wire34106 ) | ( n_n4441  &  wire34102 ) ;
 assign wire34109 = ( (~ pi27)  &  (~ pi26)  &  pi16 ) ;
 assign wire34110 = ( pi27  &  pi16 ) | ( pi26  &  pi16 ) ;
 assign wire34111 = ( wire2546 ) | ( wire196  &  wire251 ) | ( wire251  &  wire2549 ) ;
 assign wire34112 = ( ni33  &  wire244 ) | ( (~ ni29)  &  wire244 ) | ( (~ nv6462)  &  wire244 ) ;
 assign wire34113 = ( ni33  &  wire251 ) | ( (~ ni29)  &  wire251 ) | ( (~ nv6462)  &  wire251 ) ;
 assign wire34115 = ( nv7447  &  wire180  &  wire154 ) | ( nv7447  &  wire152  &  wire154 ) ;
 assign wire34116 = ( wire34115 ) | ( nv7447  &  wire178  &  wire154 ) ;
 assign wire34117 = ( wire34116 ) | ( n_n4404  &  wire192  &  wire183 ) ;
 assign wire34119 = ( wire2538 ) | ( wire34117 ) | ( n_n4412  &  wire34112 ) ;
 assign wire34120 = ( wire2270 ) | ( wire732  &  wire34099 ) ;
 assign wire34124 = ( wire2262 ) | ( wire2263 ) | ( wire2267 ) | ( wire34120 ) ;
 assign wire34125 = ( wire2265 ) | ( wire2266 ) | ( wire2268 ) ;
 assign wire34127 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34128 = ( pi27  &  wire213  &  wire34127 ) | ( pi26  &  wire213  &  wire34127 ) ;
 assign wire34129 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34130 = ( (~ pi27)  &  (~ pi26)  &  wire213  &  wire34129 ) ;
 assign wire34131 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34132 = ( pi21  &  (~ pi20)  &  wire34131 ) ;
 assign wire34134 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire34135 = ( (~ pi17)  &  (~ pi16)  &  (~ wire156)  &  wire182 ) ;
 assign wire34136 = ( (~ pi17)  &  (~ pi16)  &  wire156  &  wire182 ) ;
 assign wire34137 = ( pi27  &  (~ pi16) ) | ( pi26  &  (~ pi16) ) ;
 assign wire34138 = ( (~ pi27)  &  (~ pi26)  &  (~ pi16) ) ;
 assign wire34139 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire34140 = ( n_n3693  &  wire34132 ) | ( n_n3695  &  wire34134 ) ;
 assign wire34142 = ( wire2378 ) | ( wire2381 ) | ( wire34140 ) ;
 assign wire34143 = ( wire34142 ) | ( wire2402  &  wire34137 ) | ( wire2403  &  wire34137 ) ;
 assign wire34147 = ( wire2374 ) | ( wire2375 ) | ( wire529  &  wire34138 ) ;
 assign wire34148 = ( wire2370 ) | ( wire2371 ) | ( wire2380 ) | ( wire34143 ) ;
 assign wire34150 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34151 = ( pi27  &  wire189  &  wire34150 ) | ( pi26  &  wire189  &  wire34150 ) ;
 assign wire34152 = ( wire2471 ) | ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34153 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34154 = ( (~ pi27)  &  (~ pi26)  &  wire189  &  wire34153 ) ;
 assign wire34155 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34156 = ( ni33  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34157 = ( ni33  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34158 = ( (~ pi17)  &  wire179  &  nv10153 ) ;
 assign wire34159 = ( ni33  &  wire199 ) | ( (~ ni29)  &  wire199 ) | ( (~ nv6462)  &  wire199 ) ;
 assign wire34160 = ( wire2460 ) | ( pi20  &  nv7447  &  wire153 ) | ( (~ pi20)  &  nv7447  &  wire153 ) ;
 assign wire34161 = ( wire34160 ) | ( wire3205  &  wire34156 ) | ( wire3206  &  wire34156 ) ;
 assign wire34162 = ( wire34161 ) | ( wire3214  &  wire34157 ) | ( wire3215  &  wire34157 ) ;
 assign wire34164 = ( wire2457 ) | ( wire34162 ) | ( nv10153  &  wire446 ) ;
 assign wire34165 = ( (~ pi27)  &  (~ pi26)  &  pi16 ) ;
 assign wire34167 = ( ni33  &  wire244 ) | ( (~ ni29)  &  wire244 ) | ( (~ nv6462)  &  wire244 ) ;
 assign wire34168 = ( ni33  &  wire251 ) | ( (~ ni29)  &  wire251 ) | ( (~ nv6462)  &  wire251 ) ;
 assign wire34169 = ( ni33  &  wire183 ) | ( (~ ni29)  &  wire183 ) | ( (~ nv6462)  &  wire183 ) ;
 assign wire34170 = ( wire2447 ) | ( wire178  &  wire154  &  nv7129 ) ;
 assign wire34171 = ( nv7447  &  wire180  &  wire154 ) | ( nv7447  &  wire152  &  wire154 ) ;
 assign wire34173 = ( wire2442 ) | ( wire34171 ) | ( n_n4543  &  wire34169 ) ;
 assign wire34174 = ( wire34173 ) | ( wire3185  &  wire34168 ) | ( wire3186  &  wire34168 ) ;
 assign wire34175 = ( wire34174 ) | ( wire2438 ) ;
 assign wire34176 = ( wire2279 ) | ( wire732  &  wire34155 ) ;
 assign wire34177 = ( wire34176 ) | ( pi16  &  wire1337 ) ;
 assign wire34178 = ( wire34177 ) | ( wire196  &  wire34151 ) | ( wire2474  &  wire34151 ) ;
 assign wire34180 = ( wire34178 ) | ( wire2472  &  wire34154 ) | ( wire34152  &  wire34154 ) ;
 assign wire34182 = ( wire2274 ) | ( wire2275 ) | ( wire2278 ) | ( wire34180 ) ;
 assign wire34183 = ( pi27  &  wire189  &  wire698 ) | ( pi26  &  wire189  &  wire698 ) ;
 assign wire34184 = ( wire2516 ) | ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34185 = ( (~ pi27)  &  (~ pi26)  &  wire189  &  wire698 ) ;
 assign wire34186 = ( wire2521 ) | ( (~ ni33)  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34187 = ( (~ pi17)  &  (~ pi16)  &  (~ wire156)  &  wire179 ) ;
 assign wire34188 = ( (~ pi17)  &  (~ pi16)  &  wire156  &  wire179 ) ;
 assign wire34189 = ( pi27  &  (~ pi16) ) | ( pi26  &  (~ pi16) ) ;
 assign wire34190 = ( ni33  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34191 = ( ni33  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34192 = ( wire2508 ) | ( wire3326  &  wire34190 ) | ( wire3327  &  wire34190 ) ;
 assign wire34193 = ( wire34192 ) | ( wire3307  &  wire34191 ) | ( wire3308  &  wire34191 ) ;
 assign wire34194 = ( (~ pi27)  &  (~ pi26)  &  (~ pi16) ) ;
 assign wire34195 = ( ni33  &  wire243 ) | ( (~ ni29)  &  wire243 ) | ( (~ nv6462)  &  wire243 ) ;
 assign wire34196 = ( ni33  &  wire250 ) | ( (~ ni29)  &  wire250 ) | ( (~ nv6462)  &  wire250 ) ;
 assign wire34197 = ( ni33  &  wire194 ) | ( (~ ni29)  &  wire194 ) | ( (~ nv6462)  &  wire194 ) ;
 assign wire34198 = ( wire2499 ) | ( wire196  &  wire250 ) | ( wire250  &  wire2502 ) ;
 assign wire34199 = ( nv7447  &  wire158  &  wire180 ) | ( nv7447  &  wire158  &  wire152 ) ;
 assign wire34201 = ( wire2494 ) | ( wire34199 ) | ( n_n4611  &  wire34197 ) ;
 assign wire34203 = ( wire2490 ) | ( wire2491 ) | ( wire34201 ) ;
 assign wire34204 = ( wire2288 ) | ( wire698  &  wire732 ) ;
 assign wire34206 = ( wire2286 ) | ( wire34204 ) | ( wire527  &  wire34189 ) ;
 assign wire34207 = ( wire34206 ) | ( wire196  &  wire34188 ) | ( wire2524  &  wire34188 ) ;
 assign wire34208 = ( wire2285 ) | ( wire196  &  wire34183 ) | ( wire2519  &  wire34183 ) ;
 assign wire34209 = ( wire34207 ) | ( wire2522  &  wire34187 ) | ( wire34186  &  wire34187 ) ;
 assign wire34210 = ( wire34208 ) | ( wire2517  &  wire34185 ) | ( wire34184  &  wire34185 ) ;
 assign wire34212 = ( wire2290 ) | ( wire34209 ) | ( wire34210 ) ;
 assign wire34213 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire182 ) ;
 assign wire34214 = ( (~ pi17)  &  pi27  &  pi16  &  wire182 ) ;
 assign wire34217 = ( pi17  &  pi16  &  wire209 ) | ( (~ pi17)  &  pi16  &  wire209 ) ;
 assign wire34220 = ( wire2421 ) | ( wire2422 ) | ( wire34217 ) ;
 assign wire34221 = ( wire2423 ) | ( wire2424 ) | ( wire2426 ) ;
 assign wire34223 = ( (~ pi17)  &  (~ pi27)  &  pi16  &  wire182 ) ;
 assign wire34224 = ( (~ pi17)  &  pi27  &  pi16  &  wire182 ) ;
 assign wire34227 = ( pi17  &  pi16  &  wire209 ) | ( (~ pi17)  &  pi16  &  wire209 ) ;
 assign wire34228 = ( wire34227 ) | ( wire196  &  wire34223 ) | ( wire2474  &  wire34223 ) ;
 assign wire34230 = ( wire34228 ) | ( wire2472  &  wire34224 ) | ( wire34152  &  wire34224 ) ;
 assign wire34232 = ( wire2364 ) | ( wire2365 ) | ( wire2368 ) | ( wire34230 ) ;
 assign wire34233 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire179 ) ;
 assign wire34234 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire179 ) ;
 assign wire34235 = ( (~ pi17)  &  (~ pi27)  &  (~ pi16)  &  wire182 ) ;
 assign wire34236 = ( (~ pi17)  &  pi27  &  (~ pi16)  &  wire182 ) ;
 assign wire34238 = ( (~ pi16)  &  pi27 ) ;
 assign wire34239 = ( pi17  &  (~ pi16)  &  wire209 ) | ( (~ pi17)  &  (~ pi16)  &  wire209 ) ;
 assign wire34240 = ( wire34239 ) | ( (~ pi27)  &  (~ pi16)  &  wire527 ) ;
 assign wire34241 = ( wire34240 ) | ( wire196  &  wire34234 ) | ( wire2524  &  wire34234 ) ;
 assign wire34242 = ( wire2416 ) | ( wire196  &  wire34235 ) | ( wire2519  &  wire34235 ) ;
 assign wire34243 = ( wire34241 ) | ( wire2522  &  wire34233 ) | ( wire34186  &  wire34233 ) ;
 assign wire34244 = ( wire34242 ) | ( wire2517  &  wire34236 ) | ( wire34184  &  wire34236 ) ;
 assign wire34246 = ( wire2419 ) | ( wire34243 ) | ( wire34244 ) ;
 assign wire34247 = ( pi17  &  (~ pi16)  &  wire848  &  wire209 ) | ( (~ pi17)  &  (~ pi16)  &  wire848  &  wire209 ) ;
 assign wire34248 = ( wire34247 ) | ( wire2402  &  wire34074 ) | ( wire2403  &  wire34074 ) ;
 assign wire34250 = ( wire2245 ) | ( wire529  &  wire34080 ) ;
 assign wire34253 = ( wire2243 ) | ( wire2244 ) | ( wire2251 ) | ( wire34248 ) ;
 assign wire34255 = ( wire2246 ) | ( wire2250 ) | ( wire34250 ) | ( wire34253 ) ;
 assign wire34258 = ( wire2253 ) | ( wire2260 ) | ( wire34255 ) ;
 assign wire34262 = ( wire2254 ) | ( wire2255 ) | ( wire2257 ) | ( wire2261 ) ;
 assign wire34263 = ( wire2256 ) | ( wire2258 ) | ( wire2259 ) | ( wire34258 ) ;
 assign wire34264 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34265 = ( pi27  &  wire189  &  wire34264 ) | ( (~ pi26)  &  wire189  &  wire34264 ) ;
 assign wire34266 = ( ni11  &  wire369  &  wire34265 ) ;
 assign wire34267 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34268 = ( (~ pi27)  &  pi26  &  wire189  &  wire34267 ) ;
 assign wire34271 = ( (~ pi16)  &  ni11  &  wire369  &  wire1120 ) ;
 assign wire34272 = ( (~ pi16)  &  ni11  &  wire369 ) ;
 assign wire34274 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34275 = ( ni11  &  wire369  &  wire34274 ) ;
 assign wire34276 = ( pi27  &  (~ pi16) ) | ( (~ pi26)  &  (~ pi16) ) ;
 assign wire34277 = ( ni11  &  wire369  &  wire34276 ) ;
 assign wire34278 = ( (~ pi27)  &  pi26  &  (~ pi16) ) ;
 assign wire34279 = ( ni11  &  wire369  &  wire34278 ) ;
 assign wire34280 = ( (~ pi16)  &  ni11  &  wire369 ) ;
 assign wire34281 = ( (~ pi27)  &  pi26  &  ni11  &  wire369 ) ;
 assign wire34282 = ( pi27  &  ni11  &  wire369 ) | ( (~ pi26)  &  ni11  &  wire369 ) ;
 assign wire34283 = ( pi17  &  (~ pi16)  &  ni11  &  wire369 ) ;
 assign wire34284 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34285 = ( pi27  &  wire189  &  wire34284 ) | ( (~ pi26)  &  wire189  &  wire34284 ) ;
 assign wire34286 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34287 = ( (~ pi27)  &  pi26  &  wire189  &  wire34286 ) ;
 assign wire34288 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34289 = ( (~ pi27)  &  pi26  &  pi16 ) ;
 assign wire34291 = ( wire2437 ) | ( wire734  &  wire34288 ) ;
 assign wire34292 = ( wire34291 ) | ( pi16  &  wire1306 ) ;
 assign wire34293 = ( wire34292 ) | ( wire196  &  wire34285 ) | ( wire2474  &  wire34285 ) ;
 assign wire34295 = ( wire34293 ) | ( wire2472  &  wire34287 ) | ( wire34152  &  wire34287 ) ;
 assign wire34297 = ( wire2432 ) | ( wire2433 ) | ( wire2436 ) | ( wire34295 ) ;
 assign wire34299 = ( (~ pi27)  &  pi26  &  wire213  &  wire698 ) ;
 assign wire34301 = ( pi27  &  wire213  &  wire698 ) | ( (~ pi26)  &  wire213  &  wire698 ) ;
 assign wire34302 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire34304 = ( (~ pi17)  &  (~ pi16)  &  (~ wire155)  &  wire182 ) ;
 assign wire34305 = ( (~ pi17)  &  (~ pi16)  &  wire155  &  wire182 ) ;
 assign wire34306 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire34307 = ( pi27  &  (~ pi16) ) | ( (~ pi26)  &  (~ pi16) ) ;
 assign wire34308 = ( (~ pi27)  &  pi26  &  (~ pi16) ) ;
 assign wire34311 = ( wire2478 ) | ( wire2479 ) | ( wire2482 ) | ( wire2485 ) ;
 assign wire34312 = ( wire34311 ) | ( wire527  &  wire34307 ) ;
 assign wire34313 = ( wire34312 ) | ( wire196  &  wire34301 ) | ( wire2524  &  wire34301 ) ;
 assign wire34314 = ( wire2484 ) | ( wire196  &  wire34305 ) | ( wire2519  &  wire34305 ) ;
 assign wire34315 = ( wire34313 ) | ( wire2522  &  wire34299 ) | ( wire34186  &  wire34299 ) ;
 assign wire34316 = ( wire34314 ) | ( wire2517  &  wire34304 ) | ( wire34184  &  wire34304 ) ;
 assign wire34318 = ( wire2487 ) | ( wire34315 ) | ( wire34316 ) ;
 assign wire34319 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34320 = ( pi27  &  wire189  &  wire34319 ) | ( (~ pi26)  &  wire189  &  wire34319 ) ;
 assign wire34321 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34322 = ( (~ pi27)  &  pi26  &  wire189  &  wire34321 ) ;
 assign wire34323 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34324 = ( (~ pi27)  &  pi26  &  pi16 ) ;
 assign wire34325 = ( pi27  &  pi16 ) | ( (~ pi26)  &  pi16 ) ;
 assign wire34326 = ( wire2534 ) | ( wire734  &  wire34323 ) ;
 assign wire34330 = ( wire2526 ) | ( wire2527 ) | ( wire2531 ) | ( wire34326 ) ;
 assign wire34331 = ( wire2529 ) | ( wire2530 ) | ( wire2532 ) ;
 assign wire34333 = ( wire2237 ) | ( wire734  &  wire34275 ) ;
 assign wire34334 = ( wire34333 ) | ( wire1306  &  wire34280 ) ;
 assign wire34335 = ( wire34334 ) | ( wire2402  &  wire34277 ) | ( wire2403  &  wire34277 ) ;
 assign wire34337 = ( wire2227 ) | ( wire529  &  wire34279 ) ;
 assign wire34340 = ( wire2229 ) | ( wire2230 ) | ( wire2236 ) | ( wire34335 ) ;
 assign wire34342 = ( wire2228 ) | ( wire2235 ) | ( wire34337 ) | ( wire34340 ) ;
 assign wire34344 = ( wire2238 ) | ( wire2241 ) | ( wire34342 ) ;
 assign wire34346 = ( wire2239 ) | ( wire2240 ) | ( wire34344 ) ;
 assign wire34347 = ( (~ ni9)  &  ni10  &  (~ ni7)  &  (~ ni8) ) ;
 assign wire34348 = ( (~ ni7)  &  (~ ni8)  &  wire175  &  wire330 ) ;
 assign wire34351 = ( (~ pi24)  &  nv8608  &  wire156 ) | ( (~ pi24)  &  nv8608  &  (~ wire156) ) | ( (~ pi24)  &  wire156  &  n_n11282 ) ;
 assign wire34352 = ( (~ pi23)  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34353 = ( (~ pi21)  &  (~ ni14)  &  wire34352 ) | ( (~ pi22)  &  (~ ni14)  &  wire34352 ) ;
 assign wire34354 = ( (~ pi21)  &  (~ pi23)  &  (~ pi24) ) | ( (~ pi22)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire34356 = ( pi23  &  wire818 ) | ( pi24  &  wire818 ) ;
 assign wire34357 = ( pi23  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34358 = ( (~ pi27)  &  (~ pi26)  &  wire837 ) ;
 assign wire34359 = ( pi27  &  wire837 ) | ( pi26  &  wire837 ) ;
 assign wire34360 = ( (~ pi23)  &  (~ pi24)  &  wire818 ) ;
 assign wire34361 = ( (~ pi24)  &  (~ pi27) ) ;
 assign wire34362 = ( wire2885 ) | ( wire2884 ) ;
 assign wire34363 = ( pi21  &  pi22  &  (~ pi23)  &  wire268 ) ;
 assign wire34365 = ( nv8372 ) | ( wire193  &  n_n4509 ) ;
 assign wire34366 = ( (~ pi16)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire34369 = ( wire191  &  wire213  &  wire369  &  wire34366 ) ;
 assign wire34370 = ( (~ pi16)  &  pi23 ) | ( (~ pi16)  &  pi24 ) ;
 assign wire34373 = ( wire191  &  wire213  &  wire369  &  wire34370 ) ;
 assign wire34374 = ( nv8372 ) | ( n_n4433  &  wire193 ) ;
 assign wire34375 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34377 = ( (~ wire161)  &  wire189  &  wire369  &  wire34375 ) ;
 assign wire34378 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34380 = ( wire161  &  wire189  &  wire369  &  wire34378 ) ;
 assign wire34381 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34383 = ( pi21  &  (~ pi20)  &  wire369  &  wire34381 ) ;
 assign wire34385 = ( (~ pi17)  &  pi19  &  (~ pi20)  &  (~ pi16) ) ;
 assign wire34386 = ( wire369  &  wire34385 ) ;
 assign wire34387 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34389 = ( (~ ni33)  &  wire203 ) | ( (~ ni29)  &  wire203 ) | ( (~ nv6462)  &  wire203 ) ;
 assign wire34390 = ( (~ ni33)  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34391 = ( (~ ni33)  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34394 = ( wire2949 ) | ( wire2950 ) | ( wire2951 ) | ( wire2952 ) ;
 assign wire34395 = ( wire34394 ) | ( n_n4501  &  wire34389 ) ;
 assign wire34397 = ( (~ pi16)  &  (~ pi23)  &  (~ pi24)  &  wire369 ) ;
 assign wire34398 = ( (~ ni33)  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34399 = ( (~ pi17)  &  wire179  &  nv10167 ) ;
 assign wire34400 = ( (~ ni33)  &  wire199 ) | ( (~ ni29)  &  wire199 ) | ( (~ nv6462)  &  wire199 ) ;
 assign wire34401 = ( (~ ni33)  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34404 = ( wire2954 ) | ( wire2957 ) | ( wire2958 ) | ( wire2960 ) ;
 assign wire34406 = ( wire2959 ) | ( wire34404 ) | ( n_n4441  &  wire34400 ) ;
 assign wire34407 = ( pi16  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire34410 = ( (~ pi16)  &  pi23  &  wire369 ) | ( (~ pi16)  &  pi24  &  wire369 ) ;
 assign wire34412 = ( pi16  &  pi23  &  wire369 ) | ( pi16  &  pi24  &  wire369 ) ;
 assign wire34413 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire34414 = ( wire34413  &  wire369 ) ;
 assign wire34415 = ( wire369  &  pi16 ) ;
 assign wire34417 = ( pi23  &  wire369 ) | ( pi24  &  wire369 ) ;
 assign wire34418 = ( (~ ni33)  &  wire243 ) | ( (~ ni29)  &  wire243 ) | ( (~ nv6462)  &  wire243 ) ;
 assign wire34419 = ( (~ ni33)  &  wire250 ) | ( (~ ni29)  &  wire250 ) | ( (~ nv6462)  &  wire250 ) ;
 assign wire34420 = ( wire158  &  wire152  &  wire3276 ) | ( wire158  &  wire152  &  wire3277 ) ;
 assign wire34421 = ( wire158  &  wire180  &  nv8372 ) | ( wire158  &  wire152  &  nv8372 ) ;
 assign wire34423 = ( wire2932 ) | ( wire34421 ) | ( wire193  &  wire34420 ) ;
 assign wire34424 = ( wire34423 ) | ( n_n4489  &  wire34419 ) ;
 assign wire34425 = ( wire34424 ) | ( n_n4481  &  wire34418 ) ;
 assign wire34426 = ( (~ pi23)  &  (~ pi24)  &  wire369 ) ;
 assign wire34427 = ( wire2947 ) | ( wire197  &  wire251 ) | ( wire251  &  wire3444 ) ;
 assign wire34429 = ( (~ ni33)  &  wire244 ) | ( (~ ni29)  &  wire244 ) | ( (~ nv6462)  &  wire244 ) ;
 assign wire34430 = ( (~ ni33)  &  wire251 ) | ( (~ ni29)  &  wire251 ) | ( (~ nv6462)  &  wire251 ) ;
 assign wire34432 = ( wire180  &  nv8372  &  wire154 ) | ( wire152  &  nv8372  &  wire154 ) ;
 assign wire34433 = ( wire34432 ) | ( wire178  &  nv8372  &  wire154 ) ;
 assign wire34434 = ( wire34433 ) | ( n_n4404  &  wire193  &  wire183 ) ;
 assign wire34436 = ( wire2939 ) | ( wire34434 ) | ( n_n4412  &  wire34429 ) ;
 assign wire34437 = ( (~ pi23)  &  (~ pi24)  &  wire369 ) ;
 assign wire34438 = ( pi17  &  (~ pi16)  &  wire369 ) ;
 assign wire34439 = ( pi17  &  pi16  &  wire369 ) ;
 assign wire34440 = ( wire3030 ) | ( ni33  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34441 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34442 = ( (~ pi23)  &  (~ pi24)  &  wire189  &  wire34441 ) ;
 assign wire34443 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34444 = ( pi23  &  wire189  &  wire34443 ) | ( pi24  &  wire189  &  wire34443 ) ;
 assign wire34445 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34446 = ( (~ ni33)  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34447 = ( (~ ni33)  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34448 = ( (~ pi17)  &  wire179  &  nv10167 ) ;
 assign wire34449 = ( (~ ni33)  &  wire199 ) | ( (~ ni29)  &  wire199 ) | ( (~ nv6462)  &  wire199 ) ;
 assign wire34450 = ( wire3027 ) | ( pi20  &  nv8372  &  wire153 ) | ( (~ pi20)  &  nv8372  &  wire153 ) ;
 assign wire34451 = ( wire34450 ) | ( wire3205  &  wire34446 ) | ( wire3206  &  wire34446 ) ;
 assign wire34452 = ( wire34451 ) | ( wire3214  &  wire34447 ) | ( wire3215  &  wire34447 ) ;
 assign wire34454 = ( wire3024 ) | ( wire34452 ) | ( nv10167  &  wire385 ) ;
 assign wire34455 = ( pi16  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire34457 = ( wire3020 ) | ( wire178  &  wire154  &  nv6886 ) ;
 assign wire34458 = ( (~ ni33)  &  wire244 ) | ( (~ ni29)  &  wire244 ) | ( (~ nv6462)  &  wire244 ) ;
 assign wire34459 = ( (~ ni33)  &  wire251 ) | ( (~ ni29)  &  wire251 ) | ( (~ nv6462)  &  wire251 ) ;
 assign wire34460 = ( (~ ni33)  &  wire183 ) | ( (~ ni29)  &  wire183 ) | ( (~ nv6462)  &  wire183 ) ;
 assign wire34461 = ( wire180  &  nv8372  &  wire154 ) | ( wire152  &  nv8372  &  wire154 ) ;
 assign wire34463 = ( wire3015 ) | ( wire34461 ) | ( n_n4543  &  wire34460 ) ;
 assign wire34464 = ( wire34463 ) | ( wire3185  &  wire34459 ) | ( wire3186  &  wire34459 ) ;
 assign wire34465 = ( wire34464 ) | ( wire3011 ) ;
 assign wire34467 = ( wire2618 ) | ( wire2621 ) | ( wire2624 ) ;
 assign wire34468 = ( wire34467 ) | ( wire197  &  wire34444 ) | ( wire3339  &  wire34444 ) ;
 assign wire34470 = ( wire34468 ) | ( wire3031  &  wire34442 ) | ( wire34440  &  wire34442 ) ;
 assign wire34472 = ( wire2619 ) | ( wire2620 ) | ( wire2622 ) | ( wire34470 ) ;
 assign wire34473 = ( wire3000 ) | ( ni33  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34474 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34475 = ( (~ pi23)  &  (~ pi24)  &  wire189  &  wire34474 ) ;
 assign wire34476 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34477 = ( pi23  &  wire189  &  wire34476 ) | ( pi24  &  wire189  &  wire34476 ) ;
 assign wire34478 = ( (~ pi16)  &  pi23 ) | ( (~ pi16)  &  pi24 ) ;
 assign wire34479 = ( (~ pi17)  &  wire179  &  wire34478 ) ;
 assign wire34480 = ( (~ ni33)  &  wire169 ) | ( (~ ni29)  &  wire169 ) | ( (~ nv6462)  &  wire169 ) ;
 assign wire34481 = ( (~ ni33)  &  wire171 ) | ( (~ ni29)  &  wire171 ) | ( (~ nv6462)  &  wire171 ) ;
 assign wire34482 = ( wire2981 ) | ( wire3326  &  wire34480 ) | ( wire3327  &  wire34480 ) ;
 assign wire34483 = ( wire34482 ) | ( wire3307  &  wire34481 ) | ( wire3308  &  wire34481 ) ;
 assign wire34484 = ( wire2983 ) | ( ni33  &  ni30 ) | ( ni31  &  ni30 ) ;
 assign wire34485 = ( (~ pi16)  &  (~ pi23)  &  (~ pi24) ) ;
 assign wire34486 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34487 = ( (~ pi16)  &  pi23 ) | ( (~ pi16)  &  pi24 ) ;
 assign wire34488 = ( wire2995 ) | ( wire197  &  wire250 ) | ( wire250  &  wire3278 ) ;
 assign wire34489 = ( (~ ni33)  &  wire243 ) | ( (~ ni29)  &  wire243 ) | ( (~ nv6462)  &  wire243 ) ;
 assign wire34490 = ( (~ ni33)  &  wire250 ) | ( (~ ni29)  &  wire250 ) | ( (~ nv6462)  &  wire250 ) ;
 assign wire34491 = ( (~ ni33)  &  wire194 ) | ( (~ ni29)  &  wire194 ) | ( (~ nv6462)  &  wire194 ) ;
 assign wire34492 = ( wire158  &  wire180  &  nv8372 ) | ( wire158  &  wire152  &  nv8372 ) ;
 assign wire34494 = ( wire2990 ) | ( wire34492 ) | ( n_n4611  &  wire34491 ) ;
 assign wire34496 = ( wire2986 ) | ( wire2987 ) | ( wire34494 ) ;
 assign wire34498 = ( wire2629 ) | ( wire2631 ) | ( wire2634 ) ;
 assign wire34499 = ( wire34498 ) | ( wire447  &  wire34487 ) ;
 assign wire34500 = ( wire34499 ) | ( wire197  &  wire34479 ) | ( wire3320  &  wire34479 ) ;
 assign wire34501 = ( wire34500 ) | ( wire197  &  wire34477 ) | ( wire3316  &  wire34477 ) ;
 assign wire34503 = ( wire2632 ) | ( wire891  &  wire34485 ) ;
 assign wire34504 = ( wire2625 ) | ( wire34501 ) | ( (~ wire161)  &  wire673 ) ;
 assign wire34505 = ( n_n3014  &  wire34383 ) | ( n_n3016  &  wire34386 ) ;
 assign wire34507 = ( n_n3016  &  wire34414 ) | ( wire3144  &  wire34414 ) | ( n_n3016  &  wire34438 ) | ( wire3144  &  wire34438 ) ;
 assign wire34508 = ( wire2606 ) | ( n_n3016  &  wire34439 ) | ( wire3144  &  wire34439 ) ;
 assign wire34509 = ( wire2600 ) | ( wire34505 ) | ( wire34507 ) ;
 assign wire34511 = ( wire34508 ) | ( wire34509 ) | ( wire613  &  nv8369 ) ;
 assign wire34513 = ( wire2595 ) | ( wire2597 ) | ( wire34511 ) ;
 assign wire34518 = ( wire2594 ) | ( wire2602 ) | ( wire2604 ) | ( wire34513 ) ;
 assign wire34519 = ( wire2596 ) | ( wire2603 ) | ( wire2607 ) | ( wire2609 ) ;
 assign wire34522 = ( wire34518 ) | ( wire34519 ) | ( wire649  &  wire34397 ) ;
 assign wire34523 = ( wire2608 ) | ( wire34522 ) | ( wire652  &  wire34437 ) ;
 assign wire34525 = ( wire2585 ) | ( wire2889  &  wire34353 ) | ( wire34351  &  wire34353 ) ;
 assign wire34526 = ( wire2587 ) | ( wire161  &  wire268  &  wire597 ) ;
 assign wire34527 = ( wire34525 ) | ( wire2906  &  wire34360 ) | ( wire2907  &  wire34360 ) ;
 assign wire34529 = ( wire2591 ) | ( wire618  &  nv8369 ) ;
 assign wire34530 = ( wire34527 ) | ( wire2886  &  wire34363 ) | ( wire34362  &  wire34363 ) ;
 assign wire34532 = ( wire2586 ) | ( wire34526 ) | ( wire34529 ) | ( wire34530 ) ;
 assign wire34533 = ( (~ ni9)  &  (~ ni10)  &  (~ ni7)  &  ni8 ) ;
 assign wire34534 = ( (~ pi17)  &  pi16  &  (~ pi15) ) ;
 assign wire34536 = ( pi25  &  wire182  &  wire359  &  wire34534 ) ;
 assign wire34537 = ( (~ pi17)  &  pi16  &  (~ pi15) ) ;
 assign wire34540 = ( pi25  &  wire180  &  wire359  &  wire614 ) ;
 assign wire34542 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire359 ) ;
 assign wire34543 = ( pi17  &  pi16  &  (~ pi15)  &  wire359 ) ;
 assign wire34545 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire34547 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire179 ) ;
 assign wire34548 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire34549 = ( pi17  &  pi25  &  (~ pi16)  &  wire180 ) ;
 assign wire34550 = ( wire906 ) | ( n_n4611  &  wire393 ) ;
 assign wire34551 = ( wire2681 ) | ( wire34550 ) | ( wire194  &  wire248 ) ;
 assign wire34553 = ( wire34551 ) | ( wire2659 ) ;
 assign wire34555 = ( wire2654 ) | ( wire2657 ) | ( wire2658 ) | ( wire34553 ) ;
 assign wire34557 = ( wire2655 ) | ( wire2652 ) ;
 assign wire34558 = ( wire2653 ) | ( wire34555 ) | ( wire158  &  wire1326 ) ;
 assign wire34560 = ( pi17  &  pi25  &  (~ pi16)  &  wire180 ) ;
 assign wire34561 = ( pi17  &  pi25  &  (~ pi16)  &  wire178 ) ;
 assign wire34562 = ( (~ pi17)  &  pi25  &  pi16  &  wire182 ) ;
 assign wire34563 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire182 ) ;
 assign wire34564 = ( pi17  &  pi25  &  pi16  &  wire180 ) ;
 assign wire34566 = ( wire1352 ) | ( wire2676 ) | ( n_n4404  &  wire311 ) ;
 assign wire34567 = ( wire34566 ) | ( wire152  &  wire154  &  wire248 ) ;
 assign wire34571 = ( wire575 ) | ( wire957 ) | ( wire2672 ) ;
 assign wire34572 = ( wire2668 ) | ( wire2675 ) | ( n_n4489  &  wire34561 ) ;
 assign wire34573 = ( wire2671 ) | ( wire34567 ) | ( wire34571 ) ;
 assign wire34574 = ( n_n4481  &  wire34560 ) | ( n_n4433  &  wire34562 ) ;
 assign wire34575 = ( n_n4501  &  wire34563 ) | ( n_n4412  &  wire34564 ) ;
 assign wire34579 = ( wire2669 ) | ( wire34575 ) | ( wire154  &  wire1297 ) ;
 assign wire34580 = ( wire2674 ) | ( wire34572 ) | ( wire34573 ) | ( wire34574 ) ;
 assign wire34582 = ( wire1071  &  wire359 ) ;
 assign wire34584 = ( pi17  &  pi16  &  (~ pi15)  &  wire359 ) ;
 assign wire34585 = ( (~ pi15)  &  wire152  &  wire154  &  wire359 ) ;
 assign wire34586 = ( pi16  &  (~ pi15)  &  wire359 ) ;
 assign wire34588 = ( pi19  &  pi20  &  pi16  &  (~ pi15) ) ;
 assign wire34590 = ( (~ pi17)  &  (~ ni14)  &  wire181  &  wire34588 ) ;
 assign wire34591 = ( (~ pi19)  &  pi20  &  (~ ni14) ) ;
 assign wire34593 = ( wire181  &  wire614  &  wire34591 ) ;
 assign wire34594 = ( wire2811 ) | ( pi21  &  n_n3693 ) ;
 assign wire34595 = ( (~ ni14)  &  (~ pi17) ) ;
 assign wire34596 = ( pi19  &  pi20  &  pi16  &  (~ pi15) ) ;
 assign wire34598 = ( pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34600 = ( wire228  &  wire181  &  wire34598 ) ;
 assign wire34602 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34604 = ( (~ pi19)  &  pi20  &  (~ ni14)  &  wire614 ) ;
 assign wire34606 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34608 = ( pi16  &  (~ pi15)  &  (~ ni14)  &  wire228 ) ;
 assign wire34609 = ( pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34610 = ( pi17  &  pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34612 = ( pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34613 = ( (~ pi15)  &  (~ ni14)  &  wire257 ) ;
 assign wire34614 = ( pi17  &  pi16  &  (~ pi15)  &  (~ ni14) ) ;
 assign wire34615 = ( (~ pi15)  &  (~ ni14)  &  wire152  &  wire154 ) ;
 assign wire34617 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire34620 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire34621 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34623 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34624 = ( pi21  &  pi22  &  pi25  &  wire34623 ) ;
 assign wire34626 = ( pi16  &  (~ pi17) ) ;
 assign wire34627 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34628 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire34629 = ( wire2764 ) | ( n_n4404  &  wire311 ) ;
 assign wire34631 = ( wire183  &  wire273 ) | ( pi16  &  wire1320 ) ;
 assign wire34633 = ( wire2812  &  wire34627 ) | ( wire34594  &  wire34627 ) | ( wire2812  &  wire34628 ) | ( wire34594  &  wire34628 ) ;
 assign wire34636 = ( wire2752 ) | ( wire2754 ) | ( wire34629 ) | ( wire34633 ) ;
 assign wire34637 = ( wire2756 ) | ( wire2761 ) | ( wire2762 ) | ( wire34631 ) ;
 assign wire34638 = ( wire34636 ) | ( n_n4433  &  wire181  &  wire34617 ) ;
 assign wire34640 = ( wire34637 ) | ( pi17  &  pi16  &  wire1297 ) ;
 assign wire34642 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire34645 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire34647 = ( pi20  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire34648 = ( pi21  &  pi22  &  pi25  &  wire1293 ) ;
 assign wire34650 = ( (~ pi16)  &  ni30  &  wire156 ) | ( (~ pi16)  &  (~ wire156)  &  nv7447 ) ;
 assign wire34651 = ( pi17  &  (~ pi16)  &  wire766 ) ;
 assign wire34654 = ( wire247  &  wire34650 ) | ( n_n3693  &  wire34651 ) ;
 assign wire34656 = ( wire1352 ) | ( wire2767 ) | ( wire2775 ) | ( wire34654 ) ;
 assign wire34659 = ( wire2770 ) | ( wire34656 ) | ( wire243  &  wire273 ) ;
 assign wire34661 = ( wire1066  &  wire2812 ) | ( wire1066  &  wire34594 ) | ( wire2812  &  wire34645 ) | ( wire34594  &  wire34645 ) ;
 assign wire34663 = ( wire959 ) | ( wire2771 ) | ( wire2778 ) | ( wire2781 ) ;
 assign wire34664 = ( wire2780 ) | ( wire34659 ) | ( wire34661 ) ;
 assign wire34665 = ( wire34663 ) | ( n_n4489  &  wire181  &  wire1066 ) ;
 assign wire34666 = ( wire34664 ) | ( n_n4501  &  wire181  &  wire34642 ) ;
 assign wire34670 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire34671 = ( pi21  &  pi22  &  pi25  &  wire34670 ) ;
 assign wire34673 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire34675 = ( (~ pi17)  &  pi25  &  (~ pi16)  &  wire179 ) ;
 assign wire34676 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire34677 = ( pi21  &  pi22  &  pi25  &  wire34676 ) ;
 assign wire34678 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire34679 = ( pi21  &  pi22  &  pi25  &  wire34678 ) ;
 assign wire34680 = ( (~ pi16)  &  (~ pi17) ) ;
 assign wire34681 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire34682 = ( (~ pi17)  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire34683 = ( (~ pi20)  &  pi25  &  (~ pi16)  &  wire153 ) ;
 assign wire34684 = ( wire1285 ) | ( wire2798 ) | ( wire194  &  wire273 ) ;
 assign wire34686 = ( wire2812  &  wire34681 ) | ( wire34594  &  wire34681 ) | ( wire2812  &  wire34682 ) | ( wire34594  &  wire34682 ) ;
 assign wire34689 = ( wire2785 ) | ( wire2788 ) | ( wire34684 ) ;
 assign wire34690 = ( wire2792 ) | ( wire2794 ) | ( wire34686 ) ;
 assign wire34692 = ( wire2789 ) | ( wire2795 ) | ( wire34689 ) | ( wire34690 ) ;
 assign wire34694 = ( wire2787 ) | ( wire2784 ) ;
 assign wire34695 = ( wire2786 ) | ( wire34692 ) | ( wire158  &  wire1326 ) ;
 assign wire34696 = ( wire2744 ) | ( (~ pi15)  &  (~ ni14)  &  wire906 ) ;
 assign wire34697 = ( wire34696 ) | ( wire273  &  wire34615 ) ;
 assign wire34699 = ( wire2812  &  wire34604 ) | ( wire34594  &  wire34604 ) | ( wire2812  &  wire34608 ) | ( wire34594  &  wire34608 ) ;
 assign wire34702 = ( wire2735 ) | ( wire2736 ) | ( wire2745 ) ;
 assign wire34703 = ( wire2743 ) | ( wire34697 ) | ( wire34699 ) ;
 assign wire34705 = ( wire2739 ) | ( wire2741 ) | ( wire34702 ) | ( wire34703 ) ;
 assign wire34707 = ( wire2734 ) | ( wire1311  &  wire34602 ) ;
 assign wire34708 = ( wire2733 ) | ( wire2742 ) | ( wire34705 ) ;
 assign wire34709 = ( wire34707 ) | ( pi15  &  (~ ni14)  &  n_n4542 ) ;
 assign wire34710 = ( wire34708 ) | ( pi15  &  (~ ni14)  &  n_n4541 ) ;
 assign wire34712 = ( wire209  &  wire34582 ) | ( wire248  &  wire34585 ) ;
 assign wire34714 = ( wire2648 ) | ( wire2646 ) ;
 assign wire34716 = ( wire2640 ) | ( wire2645 ) | ( wire34712 ) | ( wire34714 ) ;
 assign wire34718 = ( wire2639 ) | ( wire1311  &  wire359  &  wire34537 ) ;
 assign wire34719 = ( wire2637 ) | ( wire2641 ) | ( wire34716 ) ;
 assign wire34722 = ( wire2642 ) | ( wire2643 ) | ( wire34718 ) | ( wire34719 ) ;
 assign wire34724 = ( wire2649 ) | ( wire34722 ) | ( nv6450  &  wire618 ) ;
 assign wire34725 = ( (~ ni9)  &  (~ ni10)  &  (~ ni7)  &  (~ ni8) ) ;
 assign wire34726 = ( pi24  &  ni31  &  ni30 ) ;
 assign wire34731 = ( pi21  &  pi22  &  (~ pi24) ) ;
 assign wire34733 = ( (~ pi24)  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34734 = ( (~ pi24)  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34735 = ( pi24  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34739 = ( (~ pi17)  &  (~ pi16)  &  wire179  &  wire369 ) ;
 assign wire34741 = ( (~ pi17)  &  (~ pi16)  &  wire179  &  wire369 ) ;
 assign wire34742 = ( (~ pi17)  &  (~ pi24)  &  wire179  &  wire34741 ) ;
 assign wire34744 = ( pi16  &  wire369  &  wire1114 ) ;
 assign wire34745 = ( wire369  &  pi16 ) ;
 assign wire34748 = ( (~ pi16)  &  pi24  &  wire369 ) ;
 assign wire34749 = ( pi24  &  pi16 ) ;
 assign wire34752 = ( (~ pi16)  &  (~ pi24)  &  wire369 ) ;
 assign wire34754 = ( pi16  &  (~ pi24)  &  wire369 ) ;
 assign wire34755 = ( wire369  &  (~ pi24) ) ;
 assign wire34758 = ( wire369  &  pi24 ) ;
 assign wire34761 = ( (~ pi17)  &  (~ pi16)  &  (~ pi24)  &  wire179 ) ;
 assign wire34763 = ( (~ pi17)  &  (~ pi16)  &  pi24  &  wire182 ) ;
 assign wire34765 = ( pi17  &  (~ pi16)  &  wire336 ) | ( (~ pi17)  &  (~ pi16)  &  wire336 ) ;
 assign wire34766 = ( wire34765 ) | ( wire197  &  wire34761 ) | ( wire3320  &  wire34761 ) ;
 assign wire34767 = ( wire34766 ) | ( wire3001  &  wire34763 ) | ( wire34473  &  wire34763 ) ;
 assign wire34769 = ( wire34767 ) | ( (~ pi16)  &  pi24  &  wire891 ) ;
 assign wire34770 = ( wire2972 ) | ( pi24  &  wire673 ) | ( (~ pi24)  &  wire678 ) ;
 assign wire34771 = ( (~ pi17)  &  pi16  &  (~ pi24)  &  wire182 ) ;
 assign wire34772 = ( (~ pi17)  &  pi16  &  pi24  &  wire182 ) ;
 assign wire34775 = ( pi17  &  pi16  &  wire336 ) | ( (~ pi17)  &  pi16  &  wire336 ) ;
 assign wire34776 = ( wire34775 ) | ( wire197  &  wire34771 ) | ( wire3339  &  wire34771 ) ;
 assign wire34778 = ( wire34776 ) | ( wire3031  &  wire34772 ) | ( wire34440  &  wire34772 ) ;
 assign wire34780 = ( wire3005 ) | ( wire3006 ) | ( wire3008 ) | ( wire34778 ) ;
 assign wire34782 = ( (~ pi17)  &  wire336  &  wire369 ) | ( pi17  &  pi16  &  wire336  &  wire369 ) | ( pi17  &  (~ pi16)  &  wire336  &  wire369 ) ;
 assign wire34783 = ( wire34782 ) | ( nv8638  &  wire613 ) ;
 assign wire34785 = ( wire2911 ) | ( wire2912 ) | ( wire34783 ) ;
 assign wire34790 = ( wire2910 ) | ( wire2915 ) | ( wire2917 ) | ( wire34785 ) ;
 assign wire34791 = ( wire2913 ) | ( wire2916 ) | ( wire2918 ) | ( wire2920 ) ;
 assign wire34794 = ( wire34790 ) | ( wire34791 ) | ( wire649  &  wire34748 ) ;
 assign wire34795 = ( wire2919 ) | ( wire34794 ) | ( wire652  &  wire34758 ) ;
 assign wire34798 = ( wire2893 ) | ( wire2894 ) | ( wire2900 ) ;
 assign wire34801 = ( wire2897 ) | ( wire2899 ) | ( wire2901 ) | ( wire34798 ) ;
 assign wire34803 = ( wire2896 ) | ( wire34801 ) ;
 assign wire34804 = ( wire2895 ) | ( wire2898 ) | ( nv8638  &  wire618 ) ;
 assign wire34806 = ( (~ ni9)  &  ni10  &  (~ ni7)  &  ni8 ) ;
 assign wire34810 = ( wire3122 ) | ( wire912  &  wire3125 ) | ( wire912  &  wire3126 ) ;
 assign wire34813 = ( wire3117 ) | ( wire3118 ) | ( wire34810 ) ;
 assign wire34814 = ( wire3119 ) | ( wire3120 ) | ( wire3121 ) | ( wire34813 ) ;
 assign wire34815 = ( ni8  &  ni7 ) ;
 assign wire34816 = ( (~ ni7)  &  ni9 ) ;
 assign wire34817 = ( pi23  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34819 = ( (~ wire793)  &  wire921  &  wire34817 ) ;
 assign wire34820 = ( (~ pi21)  &  pi23  &  (~ pi24) ) | ( (~ pi22)  &  pi23  &  (~ pi24) ) ;
 assign wire34823 = ( pi21  &  pi22  &  (~ ni8) ) ;
 assign wire34825 = ( (~ wire175)  &  wire264  &  wire160  &  wire34823 ) ;
 assign wire34826 = ( pi21  &  pi22  &  (~ ni8) ) ;
 assign wire34828 = ( (~ wire175)  &  wire264  &  (~ wire160)  &  wire34826 ) ;
 assign wire34830 = ( (~ pi21)  &  pi23  &  (~ ni8) ) | ( (~ pi22)  &  pi23  &  (~ ni8) ) ;
 assign wire34831 = ( (~ wire175)  &  wire264  &  wire34830 ) ;
 assign wire34833 = ( (~ pi23)  &  wire818  &  (~ wire793) ) | ( pi24  &  wire818  &  (~ wire793) ) ;
 assign wire34834 = ( (~ pi23)  &  (~ ni13)  &  (~ ni11)  &  ni12 ) ;
 assign wire34835 = ( (~ ni9)  &  ni10  &  (~ ni8)  &  wire34834 ) ;
 assign wire34837 = ( pi23  &  (~ pi24)  &  wire818  &  (~ wire793) ) ;
 assign wire34838 = ( pi23  &  (~ ni9)  &  ni10  &  (~ ni8) ) ;
 assign wire34839 = ( pi21  &  pi22  &  wire268  &  wire34838 ) ;
 assign wire34841 = ( (~ pi23)  &  wire268  &  (~ wire793) ) | ( pi24  &  wire268  &  (~ wire793) ) ;
 assign wire34843 = ( (~ pi23)  &  (~ ni8)  &  (~ wire175)  &  wire264 ) ;
 assign wire34844 = ( (~ pi21)  &  pi23  &  (~ pi24) ) ;
 assign wire34845 = ( (~ pi22)  &  pi23  &  (~ pi24) ) ;
 assign wire34846 = ( pi21  &  pi22  &  pi23  &  (~ pi24) ) ;
 assign wire34848 = ( ni11  &  (~ ni9)  &  ni10  &  (~ ni8) ) ;
 assign wire34850 = ( (~ pi23)  &  (~ ni9)  &  ni10  &  (~ ni8) ) ;
 assign wire34851 = ( (~ ni9)  &  ni10  &  (~ ni8)  &  wire618 ) ;
 assign wire34853 = ( wire160  &  wire189  &  wire369  &  wire1031 ) ;
 assign wire34855 = ( (~ wire160)  &  wire189  &  wire369  &  wire1031 ) ;
 assign wire34857 = ( (~ wire160)  &  wire213  &  wire369  &  wire698 ) ;
 assign wire34859 = ( wire160  &  wire213  &  wire369  &  wire698 ) ;
 assign wire34860 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire34861 = ( wire34860  &  wire369 ) ;
 assign wire34862 = ( (~ pi17)  &  (~ pi19)  &  pi16 ) | ( (~ pi17)  &  (~ pi20)  &  pi16 ) ;
 assign wire34863 = ( wire34862  &  wire369 ) ;
 assign wire34865 = ( (~ pi16)  &  pi23  &  (~ pi24)  &  wire369 ) ;
 assign wire34866 = ( pi16  &  pi23  &  (~ pi24) ) ;
 assign wire34869 = ( (~ pi16)  &  (~ pi23)  &  wire369 ) | ( (~ pi16)  &  pi24  &  wire369 ) ;
 assign wire34871 = ( pi16  &  (~ pi23)  &  wire369 ) | ( pi16  &  pi24  &  wire369 ) ;
 assign wire34874 = ( pi17  &  (~ pi16)  &  wire369 ) ;
 assign wire34875 = ( pi17  &  pi16  &  wire369 ) ;
 assign wire34876 = ( (~ pi23)  &  wire369 ) | ( pi24  &  wire369 ) ;
 assign wire34877 = ( pi23  &  (~ pi24)  &  wire369 ) ;
 assign wire34879 = ( pi23  &  (~ pi24)  &  wire369 ) ;
 assign wire34880 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34881 = ( pi23  &  (~ pi24)  &  wire213  &  wire34880 ) ;
 assign wire34882 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34883 = ( (~ pi23)  &  wire213  &  wire34882 ) | ( pi24  &  wire213  &  wire34882 ) ;
 assign wire34884 = ( (~ pi17)  &  (~ pi16)  &  (~ wire160)  &  wire182 ) ;
 assign wire34885 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire34886 = ( (~ pi16)  &  (~ pi23) ) | ( (~ pi16)  &  pi24 ) ;
 assign wire34887 = ( (~ pi16)  &  pi23  &  (~ pi24) ) ;
 assign wire34888 = ( (~ pi17)  &  (~ pi19)  &  (~ pi16) ) | ( (~ pi17)  &  pi20  &  (~ pi16) ) ;
 assign wire34890 = ( wire2858 ) | ( wire2861 ) | ( wire2864 ) ;
 assign wire34891 = ( wire34890 ) | ( wire197  &  wire34883 ) | ( wire3320  &  wire34883 ) ;
 assign wire34894 = ( wire2857 ) | ( wire641  &  wire34886 ) ;
 assign wire34895 = ( wire2855 ) | ( wire2860 ) | ( wire2862 ) | ( wire34891 ) ;
 assign wire34897 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34898 = ( (~ pi23)  &  wire189  &  wire34897 ) | ( pi24  &  wire189  &  wire34897 ) ;
 assign wire34899 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34900 = ( pi23  &  (~ pi24)  &  wire189  &  wire34899 ) ;
 assign wire34901 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire34902 = ( pi16  &  pi23  &  (~ pi24) ) ;
 assign wire34904 = ( (~ pi17)  &  (~ pi19)  &  pi16 ) | ( (~ pi17)  &  (~ pi20)  &  pi16 ) ;
 assign wire34906 = ( wire2869 ) | ( wire2872 ) | ( wire2875 ) ;
 assign wire34907 = ( wire34906 ) | ( wire197  &  wire34898 ) | ( wire3339  &  wire34898 ) ;
 assign wire34909 = ( wire34907 ) | ( wire3031  &  wire34900 ) | ( wire34440  &  wire34900 ) ;
 assign wire34911 = ( wire2870 ) | ( wire2871 ) | ( wire2873 ) | ( wire34909 ) ;
 assign wire34912 = ( n_n2546  &  wire34861 ) | ( wire2878  &  wire34861 ) | ( n_n2546  &  wire34863 ) | ( wire2878  &  wire34863 ) ;
 assign wire34914 = ( n_n2546  &  wire34874 ) | ( wire2878  &  wire34874 ) | ( n_n2546  &  wire34875 ) | ( wire2878  &  wire34875 ) ;
 assign wire34916 = ( wire2841 ) | ( wire2842 ) | ( wire34912 ) | ( wire34914 ) ;
 assign wire34917 = ( wire34916 ) | ( wire613  &  nv8777 ) ;
 assign wire34919 = ( wire2831 ) | ( wire2834 ) | ( wire34917 ) ;
 assign wire34924 = ( wire2833 ) | ( wire2838 ) | ( wire2840 ) | ( wire34919 ) ;
 assign wire34925 = ( wire2832 ) | ( wire2839 ) | ( wire2845 ) | ( wire2847 ) ;
 assign wire34928 = ( wire34924 ) | ( wire34925 ) | ( wire649  &  wire34865 ) ;
 assign wire34929 = ( wire2846 ) | ( wire34928 ) | ( wire652  &  wire34879 ) ;
 assign wire34931 = ( (~ ni11)  &  (~ ni9)  &  ni10  &  (~ ni8) ) ;
 assign wire34932 = ( wire2815 ) | ( wire2889  &  wire34819 ) | ( wire34351  &  wire34819 ) ;
 assign wire34934 = ( wire2820 ) | ( n_n3349  &  wire34843 ) | ( n_n3347  &  wire34843 ) ;
 assign wire34935 = ( wire2818 ) | ( wire34932 ) | ( wire597  &  wire34841 ) ;
 assign wire34939 = ( wire2826 ) | ( wire401  &  nv8777  &  wire34848 ) ;
 assign wire34940 = ( wire2816 ) | ( wire2817 ) | ( nv8777  &  wire34851 ) ;
 assign wire34942 = ( wire2819 ) | ( wire34935 ) | ( wire34939 ) ;
 assign wire34943 = ( wire2821 ) | ( wire2822 ) | ( wire34934 ) | ( wire34940 ) ;
 assign wire34945 = ( wire34942 ) | ( wire34943 ) | ( nv8350  &  wire1316 ) ;
 assign wire34947 = ( wire33910  &  wire33911 ) | ( wire33931  &  wire33932 ) ;
 assign wire34950 = ( n_n3349  &  wire33929 ) | ( n_n3347  &  wire33929 ) | ( n_n3349  &  wire33947 ) | ( n_n3347  &  wire33947 ) ;
 assign wire34951 = ( wire2128 ) | ( wire2133 ) | ( wire34947 ) | ( wire34950 ) ;
 assign wire34954 = ( wire34951 ) | ( nv8369  &  wire33945 ) ;
 assign wire34955 = ( wire2129 ) | ( wire2130 ) | ( nv8638  &  wire33952 ) ;
 assign wire34957 = ( wire2134 ) | ( wire2137 ) | ( wire34954 ) | ( wire34955 ) ;
 assign wire34958 = ( wire34957 ) | ( n_n4096  &  wire34008 ) | ( wire34007  &  wire34008 ) ;
 assign wire34959 = ( wire34958 ) | ( wire1150  &  wire34062 ) ;
 assign wire34960 = ( wire34959 ) | ( nv6450  &  wire34348 ) ;
 assign wire34962 = ( wire34960 ) | ( nv8350  &  wire34815 ) | ( nv8350  &  wire34816 ) ;
 assign wire34965 = ( wire2145 ) | ( wire34962 ) | ( n_n4697  &  wire34725 ) ;
 assign wire34966 = ( wire2141 ) | ( wire2143 ) | ( wire2148 ) ;
 assign wire34967 = ( (~ ni2)  &  (~ ni3)  &  wire281 ) ;
 assign wire34968 = ( wire2126 ) | ( wire173  &  wire33864 ) | ( wire1063  &  wire33864 ) ;
 assign wire34971 = ( wire2119 ) | ( wire2120 ) | ( wire34968 ) ;
 assign wire34973 = ( wire2121 ) | ( wire2122 ) | ( wire2124 ) | ( wire34971 ) ;
 assign wire34974 = ( ni3  &  ni31  &  ni30 ) ;
 assign wire34977 = ( ni4  &  ni3  &  ni6 ) ;
 assign wire34981 = ( (~ ni3)  &  wire29371 ) | ( (~ ni3)  &  (~ ni7)  &  n_n983 ) ;
 assign wire34983 = ( ni5  &  (~ ni3) ) ;
 assign wire34984 = ( ni3  &  (~ ni31)  &  (~ ni5) ) | ( ni3  &  (~ ni5)  &  (~ ni6) ) | ( ni3  &  ni31  &  ni5  &  ni6 ) ;
 assign wire34987 = ( wire2111 ) | ( wire2112 ) | ( wire2115 ) | ( wire34984 ) ;
 assign wire34990 = ( wire606 ) | ( (~ wire231)  &  wire1101 ) | ( (~ wire231)  &  wire2001 ) ;
 assign wire34991 = ( wire278  &  wire242 ) | ( wire278  &  wire2003 ) | ( wire278  &  wire2004 ) ;
 assign wire34992 = ( (~ pi17)  &  pi19  &  pi21  &  pi20 ) ;
 assign wire34994 = ( pi16  &  pi15  &  wire289  &  wire34992 ) ;
 assign wire34995 = ( pi21  &  (~ pi22)  &  (~ pi20) ) ;
 assign wire34996 = ( wire607 ) | ( (~ wire229)  &  wire1104 ) | ( (~ wire229)  &  wire2052 ) ;
 assign wire34997 = ( wire327  &  wire242 ) | ( wire327  &  wire2054 ) | ( wire327  &  wire2055 ) ;
 assign wire34998 = ( wire1211 ) | ( (~ ni39)  &  (~ ni36)  &  wire783 ) ;
 assign wire34999 = ( (~ ni32)  &  (~ ni35) ) ;
 assign wire35000 = ( wire398  &  wire835 ) | ( wire835  &  wire2044 ) | ( wire835  &  wire2045 ) ;
 assign wire35001 = ( wire2030 ) | ( wire878 ) ;
 assign wire35003 = ( wire35001 ) | ( wire245  &  n_n1427 ) | ( wire245  &  n_n1426 ) ;
 assign wire35004 = ( (~ pi21)  &  ni32 ) | ( (~ pi21)  &  ni30 ) ;
 assign wire35005 = ( (~ pi21)  &  (~ pi22) ) | ( (~ pi21)  &  (~ ni31) ) | ( (~ pi21)  &  (~ ni29) ) ;
 assign wire35006 = ( wire508 ) | ( wire506  &  n_n1427 ) ;
 assign wire35007 = ( wire508 ) | ( wire2025 ) | ( wire506  &  n_n1427 ) ;
 assign wire35008 = ( pi17  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire35009 = ( wire289  &  wire35008 ) ;
 assign wire35011 = ( (~ ni32)  &  ni35 ) ;
 assign wire35012 = ( wire398  &  wire836 ) | ( wire836  &  n_n1992 ) ;
 assign wire35014 = ( pi16  &  pi15  &  wire289  &  wire381 ) ;
 assign wire35015 = ( (~ ni32)  &  ni31  &  (~ ni30)  &  ni29 ) ;
 assign wire35016 = ( ni32  &  ni38 ) ;
 assign wire35017 = ( wire1213 ) | ( nv9492  &  wire35015 ) ;
 assign wire35020 = ( pi16  &  pi15  &  wire289  &  wire272 ) ;
 assign wire35021 = ( wire1987 ) | ( wire1992 ) | ( wire348  &  wire701 ) ;
 assign wire35023 = ( wire35021 ) | ( wire245  &  n_n1462 ) | ( wire245  &  n_n1463 ) ;
 assign wire35025 = ( (~ pi17)  &  wire289  &  wire182  &  wire226 ) ;
 assign wire35028 = ( wire308 ) | ( pi21  &  wire405 ) | ( (~ pi21)  &  nv9492 ) ;
 assign wire35030 = ( (~ ni32)  &  (~ ni35) ) ;
 assign wire35031 = ( wire398  &  wire835 ) | ( n_n1891  &  wire835 ) ;
 assign wire35033 = ( wire606 ) | ( (~ wire231)  &  wire1104 ) | ( (~ wire231)  &  wire1604 ) ;
 assign wire35034 = ( wire327  &  wire242 ) | ( wire327  &  wire1606 ) | ( wire327  &  wire1607 ) ;
 assign wire35035 = ( wire1385 ) | ( wire877 ) ;
 assign wire35037 = ( wire35035 ) | ( wire245  &  n_n1394 ) | ( wire245  &  n_n1395 ) ;
 assign wire35038 = ( pi16  &  pi15  &  wire289 ) ;
 assign wire35039 = ( wire607 ) | ( (~ wire229)  &  wire1101 ) | ( (~ wire229)  &  wire2083 ) ;
 assign wire35040 = ( wire278  &  wire242 ) | ( wire278  &  wire2085 ) | ( wire278  &  wire2086 ) ;
 assign wire35041 = ( wire1211 ) | ( (~ ni39)  &  (~ ni36)  &  wire780 ) ;
 assign wire35042 = ( (~ ni32)  &  ni35 ) ;
 assign wire35043 = ( wire398  &  wire836 ) | ( wire836  &  wire2107 ) | ( wire836  &  wire2108 ) ;
 assign wire35044 = ( wire2067 ) | ( wire2072 ) | ( wire701  &  wire349 ) ;
 assign wire35046 = ( wire35044 ) | ( wire245  &  n_n1494 ) | ( wire245  &  n_n1495 ) ;
 assign wire35048 = ( wire508 ) | ( wire2062 ) | ( wire506  &  n_n1495 ) ;
 assign wire35051 = ( (~ ni38)  &  (~ ni36)  &  ni32 ) ;
 assign wire35053 = ( ni32  &  (~ ni39) ) ;
 assign wire35054 = ( ni32  &  ni37 ) ;
 assign wire35055 = ( n_n2448  &  wire35051 ) | ( (~ nv401)  &  wire35054 ) ;
 assign wire35056 = ( wire35055 ) | ( ni32  &  nv401  &  nv9262 ) ;
 assign wire35057 = ( wire1938 ) | ( wire1936 ) ;
 assign wire35058 = ( wire1424 ) | ( wire782  &  wire35056 ) | ( wire782  &  wire35057 ) ;
 assign wire35060 = ( (~ ni38)  &  (~ ni36)  &  (~ ni32) ) ;
 assign wire35061 = ( nv758  &  wire293 ) | ( wire266  &  wire349 ) ;
 assign wire35062 = ( wire35061 ) | ( wire245  &  n_n1558 ) ;
 assign wire35063 = ( wire35062 ) | ( wire245  &  wire1426 ) | ( wire245  &  wire35058 ) ;
 assign wire35064 = ( wire508 ) | ( wire506  &  wire1426 ) | ( wire506  &  wire35058 ) ;
 assign wire35065 = ( wire35064 ) | ( wire1417 ) ;
 assign wire35069 = ( (~ ni38)  &  (~ ni36)  &  ni32 ) ;
 assign wire35070 = ( ni39  &  ni32 ) | ( ni38  &  ni32 ) ;
 assign wire35071 = ( ni32  &  ni37 ) ;
 assign wire35072 = ( n_n1966  &  wire35069 ) | ( (~ nv401)  &  wire35071 ) ;
 assign wire35075 = ( wire817  &  (~ pi22) ) ;
 assign wire35076 = ( pi20  &  wire316  &  wire153 ) ;
 assign wire35077 = ( pi20  &  wire293  &  wire153 ) ;
 assign wire35078 = ( pi20  &  wire245  &  wire153 ) ;
 assign wire35079 = ( (~ ni38)  &  (~ ni36)  &  (~ ni32) ) ;
 assign wire35080 = ( pi20  &  wire245  &  wire153 ) ;
 assign wire35081 = ( (~ pi17)  &  (~ pi19)  &  (~ pi21)  &  pi20 ) ;
 assign wire35082 = ( wire1404 ) | ( wire228  &  wire35004 ) | ( wire228  &  wire35005 ) ;
 assign wire35084 = ( wire1403 ) | ( wire35082 ) | ( nv772  &  wire35077 ) ;
 assign wire35085 = ( n_n1528  &  wire35080 ) | ( n_n1528  &  wire35081 ) ;
 assign wire35088 = ( wire1397 ) | ( wire1400 ) | ( wire35084 ) | ( wire35085 ) ;
 assign wire35089 = ( pi16  &  pi15  &  wire289 ) ;
 assign wire35092 = ( wire1705 ) | ( (~ ni38)  &  (~ ni36)  &  n_n1966 ) ;
 assign wire35093 = ( ni38  &  (~ ni37)  &  ni36  &  ni32 ) ;
 assign wire35094 = ( wire1458 ) | ( n_n1566  &  (~ wire782) ) ;
 assign wire35095 = ( wire441  &  wire293 ) | ( wire266  &  wire348 ) ;
 assign wire35096 = ( wire35095 ) | ( wire245  &  n_n1756 ) ;
 assign wire35097 = ( wire35096 ) | ( wire245  &  wire860 ) | ( wire245  &  wire35094 ) ;
 assign wire35098 = ( wire1447 ) | ( wire211  &  n_n1263  &  wire344 ) ;
 assign wire35099 = ( wire1101 ) | ( ni41 ) ;
 assign wire35100 = ( ni38  &  ni36  &  ni32 ) | ( ni38  &  (~ ni35)  &  ni32 ) ;
 assign wire35101 = ( ni35  &  ni32  &  wire269 ) ;
 assign wire35102 = ( wire1901 ) | ( wire1082 ) ;
 assign wire35103 = ( wire1903  &  wire35100 ) | ( wire35099  &  wire35100 ) | ( wire1903  &  wire35101 ) | ( wire35099  &  wire35101 ) ;
 assign wire35105 = ( wire1104 ) | ( ni41 ) ;
 assign wire35106 = ( (~ ni35)  &  ni32  &  wire292 ) ;
 assign wire35107 = ( ni38  &  ni36  &  ni32 ) | ( ni38  &  ni35  &  ni32 ) ;
 assign wire35108 = ( wire1803 ) | ( wire1023 ) ;
 assign wire35109 = ( wire1805  &  wire35106 ) | ( wire35105  &  wire35106 ) | ( wire1805  &  wire35107 ) | ( wire35105  &  wire35107 ) ;
 assign wire35110 = ( (~ ni38)  &  (~ ni36)  &  (~ ni35)  &  (~ ni32) ) ;
 assign wire35111 = ( (~ ni39)  &  (~ ni36)  &  (~ ni35)  &  (~ ni32) ) ;
 assign wire35112 = ( wire1231 ) | ( n_n2466  &  wire35110 ) ;
 assign wire35113 = ( nv9129  &  wire35111 ) | ( ni38  &  (~ ni32)  &  nv9129 ) ;
 assign wire35116 = ( wire878 ) | ( wire1536 ) | ( wire1537 ) | ( wire1538 ) ;
 assign wire35117 = ( wire508 ) | ( wire506  &  wire35108 ) | ( wire506  &  wire35109 ) ;
 assign wire35118 = ( wire35117 ) | ( (~ pi20)  &  n_n1247 ) ;
 assign wire35119 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire35120 = ( ni39  &  (~ ni36)  &  ni35  &  (~ ni32) ) ;
 assign wire35121 = ( (~ ni38)  &  (~ ni36)  &  ni35  &  (~ ni32) ) ;
 assign wire35122 = ( wire1230 ) | ( n_n1984  &  wire35121 ) ;
 assign wire35123 = ( nv9082  &  wire35120 ) | ( ni38  &  (~ ni32)  &  nv9082 ) ;
 assign wire35124 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire35125 = ( (~ ni32)  &  ni31  &  (~ ni30)  &  ni29 ) ;
 assign wire35129 = ( wire272  &  (~ pi16) ) ;
 assign wire35130 = ( (~ pi22)  &  pi21 ) ;
 assign wire35131 = ( wire1466 ) | ( wire35004 ) | ( wire35005 ) ;
 assign wire35133 = ( ni39  &  (~ ni36)  &  (~ ni35)  &  (~ ni32) ) ;
 assign wire35134 = ( (~ ni38)  &  (~ ni36)  &  (~ ni35)  &  (~ ni32) ) ;
 assign wire35135 = ( wire1231 ) | ( n_n1984  &  wire35134 ) ;
 assign wire35136 = ( nv9173  &  wire35133 ) | ( ni38  &  (~ ni32)  &  nv9173 ) ;
 assign wire35137 = ( wire1104 ) | ( ni41 ) ;
 assign wire35138 = ( (~ ni35)  &  ni32  &  wire269 ) ;
 assign wire35139 = ( ni38  &  ni36  &  ni32 ) | ( ni38  &  ni35  &  ni32 ) ;
 assign wire35140 = ( wire1740 ) | ( wire1023 ) ;
 assign wire35141 = ( wire1742  &  wire35138 ) | ( wire35137  &  wire35138 ) | ( wire1742  &  wire35139 ) | ( wire35137  &  wire35139 ) ;
 assign wire35142 = ( wire877 ) | ( wire245  &  wire35140 ) | ( wire245  &  wire35141 ) ;
 assign wire35143 = ( wire1474 ) | ( wire245  &  wire35135 ) | ( wire245  &  wire35136 ) ;
 assign wire35144 = ( wire35143 ) | ( wire35142 ) ;
 assign wire35145 = ( wire1101 ) | ( ni41 ) ;
 assign wire35146 = ( ni38  &  ni36  &  ni32 ) | ( ni38  &  (~ ni35)  &  ni32 ) ;
 assign wire35147 = ( ni35  &  ni32  &  wire292 ) ;
 assign wire35148 = ( wire1853 ) | ( wire1082 ) ;
 assign wire35149 = ( wire1855  &  wire35146 ) | ( wire35145  &  wire35146 ) | ( wire1855  &  wire35147 ) | ( wire35145  &  wire35147 ) ;
 assign wire35150 = ( (~ ni39)  &  (~ ni36)  &  ni35  &  (~ ni32) ) ;
 assign wire35151 = ( (~ ni38)  &  (~ ni36)  &  ni35  &  (~ ni32) ) ;
 assign wire35152 = ( wire1230 ) | ( n_n2466  &  wire35151 ) ;
 assign wire35153 = ( nv9029  &  wire35150 ) | ( ni38  &  (~ ni32)  &  nv9029 ) ;
 assign wire35156 = ( wire975 ) | ( wire1517 ) | ( wire1518 ) | ( wire1519 ) ;
 assign wire35157 = ( wire508 ) | ( wire506  &  wire35148 ) | ( wire506  &  wire35149 ) ;
 assign wire35158 = ( wire35157 ) | ( (~ pi20)  &  n_n1259 ) ;
 assign wire35159 = ( wire974 ) | ( wire245  &  wire35102 ) | ( wire245  &  wire35103 ) ;
 assign wire35160 = ( wire1543 ) | ( wire245  &  wire35122 ) | ( wire245  &  wire35123 ) ;
 assign wire35162 = ( wire1878 ) | ( (~ ni38)  &  (~ ni36)  &  n_n2448 ) ;
 assign wire35163 = ( ni38  &  (~ ni37)  &  ni36  &  ni32 ) ;
 assign wire35164 = ( wire1501 ) | ( n_n1566  &  (~ wire782) ) ;
 assign wire35165 = ( wire293  &  nv628 ) | ( wire266  &  wire349 ) ;
 assign wire35166 = ( wire35165 ) | ( wire245  &  n_n1786 ) ;
 assign wire35167 = ( wire35166 ) | ( wire316  &  nv873 ) ;
 assign wire35168 = ( wire1494 ) | ( wire2065 ) | ( wire218  &  wire34995 ) ;
 assign wire35169 = ( wire508 ) | ( wire1492 ) | ( wire1494 ) ;
 assign wire35170 = ( (~ pi16)  &  wire328 ) | ( (~ pi17)  &  (~ pi16)  &  wire309 ) ;
 assign wire35171 = ( wire35170 ) | ( wire211  &  n_n1253  &  wire698 ) ;
 assign wire35172 = ( n_n1255  &  wire35124 ) | ( n_n1593  &  wire35129 ) ;
 assign wire35174 = ( wire1270 ) | ( wire35171 ) | ( wire35172 ) ;
 assign wire35175 = ( wire35174 ) | ( n_n1111  &  wire35119 ) ;
 assign wire35176 = ( wire1273 ) | ( n_n1119  &  wire698 ) ;
 assign wire35178 = ( wire35176 ) | ( (~ pi16)  &  wire971 ) ;
 assign wire35179 = ( wire1353 ) | ( wire1448 ) | ( wire35098 ) | ( wire35175 ) ;
 assign wire35181 = ( pi17  &  (~ ni29)  &  wire180  &  wire258 ) ;
 assign wire35182 = ( pi20  &  (~ ni29)  &  wire258  &  wire153 ) ;
 assign wire35183 = ( (~ ni32)  &  (~ ni36) ) ;
 assign wire35184 = ( nv9031  &  wire341 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35186 = ( wire841 ) | ( wire1213 ) | ( wire1610 ) ;
 assign wire35187 = ( wire245  &  n_n1824 ) | ( wire245  &  n_n1823 ) ;
 assign wire35188 = ( pi16  &  (~ pi15)  &  wire272 ) ;
 assign wire35189 = ( (~ ni29)  &  wire182  &  wire507 ) ;
 assign wire35190 = ( nv539  &  (~ wire172) ) | ( nv539  &  wire1101 ) | ( nv539  &  wire2001 ) ;
 assign wire35191 = ( wire35190 ) | ( nv590  &  wire1999 ) | ( nv590  &  wire34990 ) ;
 assign wire35192 = ( pi19  &  pi21  &  pi20  &  wire507 ) ;
 assign wire35194 = ( wire1668 ) | ( wire589 ) ;
 assign wire35196 = ( pi19  &  pi20  &  wire507 ) ;
 assign wire35199 = ( wire1662 ) | ( wire1664 ) | ( wire1665 ) | ( wire1666 ) ;
 assign wire35201 = ( nv539  &  (~ wire172) ) | ( nv539  &  wire1101 ) | ( nv539  &  wire2083 ) ;
 assign wire35202 = ( wire35201 ) | ( nv590  &  wire2081 ) | ( nv590  &  wire35039 ) ;
 assign wire35203 = ( ni35  &  wire2101 ) | ( ni35  &  wire35041 ) ;
 assign wire35204 = ( wire341  &  wire780 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35206 = ( wire1959 ) | ( wire1146  &  wire418 ) | ( wire418  &  wire1970 ) ;
 assign wire35208 = ( wire35206 ) | ( wire245  &  n_n2009 ) | ( wire245  &  n_n2010 ) ;
 assign wire35210 = ( wire508 ) | ( wire1951 ) | ( wire1953 ) ;
 assign wire35211 = ( wire361  &  wire1952 ) | ( n_n1301  &  wire1952 ) | ( wire361  &  wire35210 ) | ( n_n1301  &  wire35210 ) ;
 assign wire35212 = ( wire213  &  n_n2007 ) | ( nv783  &  wire35210 ) | ( n_n2007  &  wire35210 ) ;
 assign wire35213 = ( (~ pi17)  &  pi19  &  pi16  &  (~ pi15) ) ;
 assign wire35214 = ( (~ ni35)  &  wire2050 ) | ( (~ ni32)  &  wire2050 ) | ( (~ ni35)  &  wire34996 ) | ( (~ ni32)  &  wire34996 ) ;
 assign wire35215 = ( nv539  &  (~ wire172) ) | ( nv539  &  wire1104 ) | ( nv539  &  wire2052 ) ;
 assign wire35217 = ( (~ ni35)  &  wire2040 ) | ( (~ ni35)  &  wire34998 ) ;
 assign wire35218 = ( wire341  &  wire783 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35221 = ( wire1647 ) | ( wire1649 ) | ( wire245  &  n_n1907 ) ;
 assign wire35223 = ( wire508 ) | ( wire506  &  n_n1908 ) ;
 assign wire35224 = ( wire508 ) | ( wire1643 ) | ( wire506  &  n_n1908 ) ;
 assign wire35225 = ( wire361  &  wire1642 ) | ( n_n1289  &  wire1642 ) | ( wire361  &  wire35224 ) | ( n_n1289  &  wire35224 ) ;
 assign wire35226 = ( wire213  &  n_n1905 ) | ( nv821  &  wire35224 ) | ( n_n1905  &  wire35224 ) ;
 assign wire35227 = ( pi17  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire35228 = ( wire1249 ) | ( wire245  &  wire999 ) | ( wire245  &  wire1941 ) ;
 assign wire35229 = ( wire1928 ) | ( wire245  &  wire35056 ) | ( wire245  &  wire35057 ) ;
 assign wire35231 = ( wire508 ) | ( wire506  &  wire35056 ) | ( wire506  &  wire35057 ) ;
 assign wire35232 = ( wire35231 ) | ( (~ pi20)  &  n_n1311 ) ;
 assign wire35233 = ( wire213  &  n_n2097 ) | ( wire361  &  wire35232 ) | ( n_n2097  &  wire35232 ) ;
 assign wire35234 = ( nv754  &  wire1924 ) | ( n_n1311  &  wire1924 ) | ( nv754  &  wire35232 ) | ( n_n1311  &  wire35232 ) ;
 assign wire35235 = ( (~ pi17)  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire35236 = ( (~ pi22)  &  pi21 ) ;
 assign wire35237 = ( wire1566 ) | ( wire35004 ) | ( wire35005 ) ;
 assign wire35240 = ( wire1579 ) | ( wire589 ) ;
 assign wire35242 = ( (~ ni35)  &  wire1602 ) | ( (~ ni32)  &  wire1602 ) | ( (~ ni35)  &  wire35033 ) | ( (~ ni32)  &  wire35033 ) ;
 assign wire35243 = ( nv539  &  (~ wire172) ) | ( nv539  &  wire1104 ) | ( nv539  &  wire1604 ) ;
 assign wire35245 = ( wire1575 ) | ( wire418  &  wire1142 ) | ( wire418  &  wire1754 ) ;
 assign wire35247 = ( wire35245 ) | ( wire245  &  n_n1858 ) | ( wire245  &  n_n1859 ) ;
 assign wire35248 = ( wire817  &  (~ pi22) ) ;
 assign wire35249 = ( pi20  &  wire316  &  wire153 ) ;
 assign wire35250 = ( pi20  &  wire293  &  wire153 ) ;
 assign wire35251 = ( pi20  &  wire245  &  wire153 ) ;
 assign wire35252 = ( pi20  &  wire245  &  wire153 ) ;
 assign wire35253 = ( (~ pi17)  &  (~ pi19)  &  (~ pi21)  &  pi20 ) ;
 assign wire35254 = ( wire1629 ) | ( wire228  &  wire35004 ) | ( wire228  &  wire35005 ) ;
 assign wire35257 = ( wire1625 ) | ( wire1627 ) | ( wire1628 ) | ( wire35254 ) ;
 assign wire35258 = ( wire1622 ) | ( nv772  &  wire35250 ) ;
 assign wire35261 = ( (~ pi22)  &  (~ ni37)  &  ni36  &  ni32 ) ;
 assign wire35262 = ( wire1689 ) | ( wire1982 ) | ( (~ pi22)  &  (~ ni29) ) ;
 assign wire35264 = ( wire820  &  ni36 ) ;
 assign wire35265 = ( wire1248 ) | ( (~ wire205)  &  wire408  &  wire820 ) ;
 assign wire35268 = ( wire1697 ) | ( wire1699 ) | ( wire1701 ) | ( wire35265 ) ;
 assign wire35271 = ( pi17  &  (~ pi16)  &  (~ ni29)  &  wire180 ) ;
 assign wire35272 = ( ni41  &  nv539 ) | ( nv539  &  (~ wire172) ) | ( nv539  &  nv9050 ) ;
 assign wire35273 = ( (~ ni32)  &  (~ ni36) ) ;
 assign wire35274 = ( wire341  &  wire512 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35275 = ( wire841 ) | ( wire1763 ) | ( nv9066  &  wire266 ) ;
 assign wire35276 = ( wire35275 ) | ( wire316  &  wire6691 ) | ( wire316  &  wire29623 ) ;
 assign wire35277 = ( wire245  &  n_n2143 ) | ( wire245  &  wire1765 ) | ( wire245  &  wire35272 ) ;
 assign wire35278 = ( wire272  &  (~ pi16) ) ;
 assign wire35279 = ( pi20  &  (~ pi16)  &  (~ ni29)  &  wire153 ) ;
 assign wire35280 = ( (~ pi17)  &  (~ pi16)  &  (~ ni29)  &  wire182 ) ;
 assign wire35281 = ( ni35  &  ni32  &  wire269 ) ;
 assign wire35284 = ( wire1892 ) | ( wire1893 ) | ( wire1894 ) | ( wire1895 ) ;
 assign wire35285 = ( (~ pi17)  &  (~ pi16)  &  wire617 ) ;
 assign wire35286 = ( wire341  &  nv9082 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35287 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire35288 = ( wire1798 ) | ( nv539  &  wire1805 ) | ( nv539  &  wire35105 ) ;
 assign wire35289 = ( wire341  &  nv9129 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35290 = ( wire1791 ) | ( wire418  &  wire1142 ) | ( wire418  &  wire1794 ) ;
 assign wire35292 = ( wire35290 ) | ( wire245  &  n_n2228 ) | ( wire245  &  n_n2229 ) ;
 assign wire35294 = ( wire508 ) | ( wire1787 ) | ( wire506  &  n_n2229 ) ;
 assign wire35295 = ( wire213  &  n_n2226 ) | ( wire361  &  wire35294 ) | ( n_n2226  &  wire35294 ) ;
 assign wire35297 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire35298 = ( wire1887 ) | ( wire1146  &  wire418 ) | ( wire418  &  wire1890 ) ;
 assign wire35299 = ( wire245  &  n_n2280 ) | ( wire245  &  wire1896 ) | ( wire245  &  wire35284 ) ;
 assign wire35301 = ( (~ pi17)  &  (~ pi16)  &  wire182 ) ;
 assign wire35303 = ( (~ ni36)  &  ni35  &  ni32  &  nv401 ) ;
 assign wire35304 = ( (~ ni39)  &  (~ ni36)  &  ni35  &  ni32 ) ;
 assign wire35307 = ( nv539  &  wire1855 ) | ( nv539  &  wire35145 ) | ( wire1855  &  wire35304 ) | ( wire35145  &  wire35304 ) ;
 assign wire35308 = ( wire1845 ) | ( wire1847 ) | ( wire1848 ) | ( wire35307 ) ;
 assign wire35309 = ( nv9029  &  wire341 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35310 = ( wire1833 ) | ( wire1146  &  wire418 ) | ( wire418  &  wire1970 ) ;
 assign wire35311 = ( wire1831 ) | ( wire1833 ) | ( wire245  &  n_n2332 ) ;
 assign wire35312 = ( wire1835 ) | ( wire35310 ) | ( wire245  &  n_n2332 ) ;
 assign wire35313 = ( wire508 ) | ( wire506  &  wire1849 ) | ( wire506  &  wire35308 ) ;
 assign wire35314 = ( wire1827 ) | ( wire35313 ) ;
 assign wire35315 = ( wire361  &  n_n1173 ) | ( n_n1341  &  n_n1173 ) ;
 assign wire35316 = ( n_n2327  &  n_n1173 ) | ( n_n1173  &  wire6663 ) | ( n_n1173  &  wire29629 ) ;
 assign wire35317 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire35320 = ( wire308 ) | ( wire1721 ) | ( (~ pi21)  &  n_n2143 ) ;
 assign wire35321 = ( wire341  &  nv9173 ) | ( (~ ni38)  &  ni37  &  wire341 ) ;
 assign wire35322 = ( wire1735 ) | ( nv539  &  wire1742 ) | ( nv539  &  wire35137 ) ;
 assign wire35323 = ( wire1732 ) | ( wire418  &  wire1142 ) | ( wire418  &  wire1754 ) ;
 assign wire35325 = ( wire35323 ) | ( wire245  &  n_n2179 ) | ( wire245  &  n_n2180 ) ;
 assign wire35326 = ( pi21  &  (~ pi22)  &  (~ pi20) ) ;
 assign wire35328 = ( pi21  &  (~ pi22)  &  (~ pi20) ) ;
 assign wire35329 = ( wire1866 ) | ( (~ wire782)  &  wire409  &  wire35326 ) ;
 assign wire35330 = ( pi21  &  pi22  &  (~ pi20)  &  (~ ni29) ) ;
 assign wire35332 = ( wire820  &  ni36 ) ;
 assign wire35333 = ( wire1249 ) | ( (~ wire205)  &  wire820  &  wire409 ) ;
 assign wire35336 = ( wire1872 ) | ( wire1875 ) | ( wire1876 ) | ( wire35333 ) ;
 assign wire35338 = ( wire1860 ) | ( (~ pi20)  &  n_n1351 ) ;
 assign wire35340 = ( wire1680 ) | ( (~ pi16)  &  wire157  &  wire328 ) ;
 assign wire35342 = ( wire1672 ) | ( wire1676 ) ;
 assign wire35343 = ( wire1673 ) | ( wire35340 ) | ( n_n1335  &  wire35285 ) ;
 assign wire35347 = ( wire1674 ) | ( wire1682 ) | ( wire1684 ) ;
 assign wire35348 = ( wire1263 ) | ( wire1671 ) | ( wire35342 ) | ( wire35343 ) ;
 assign wire35351 = ( wire1678 ) | ( wire1683 ) | ( wire35347 ) | ( wire35348 ) ;
 assign wire35352 = ( wire1677 ) | ( wire35315  &  wire35317 ) | ( wire35316  &  wire35317 ) ;
 assign wire35353 = ( wire1557 ) | ( wire157  &  wire258  &  wire328 ) ;
 assign wire35354 = ( wire1548 ) | ( wire35353 ) ;
 assign wire35356 = ( wire1549 ) | ( wire35354 ) | ( wire758  &  wire258 ) ;
 assign wire35359 = ( wire1551 ) | ( wire1552 ) | ( wire35356 ) ;
 assign wire35360 = ( wire1547 ) | ( wire1550 ) | ( wire258  &  wire997 ) ;
 assign wire35363 = ( wire1553 ) | ( wire1556 ) | ( wire35359 ) | ( wire35360 ) ;
 assign wire35365 = ( wire1554 ) | ( wire35363 ) | ( wire258  &  wire972 ) ;
 assign wire35366 = ( wire1555 ) | ( (~ pi15)  &  wire35351 ) | ( (~ pi15)  &  wire35352 ) ;
 assign wire35367 = ( pi17  &  (~ ni29)  &  wire180  &  wire226 ) ;
 assign wire35368 = ( pi20  &  (~ ni29)  &  wire226  &  wire153 ) ;
 assign wire35370 = ( (~ ni29)  &  wire395  &  wire182 ) ;
 assign wire35371 = ( pi19  &  pi21  &  pi20  &  wire395 ) ;
 assign wire35372 = ( pi19  &  pi20  &  wire395 ) ;
 assign wire35373 = ( wire361  &  wire2024 ) | ( n_n1207  &  wire2024 ) | ( wire361  &  wire35007 ) | ( n_n1207  &  wire35007 ) ;
 assign wire35374 = ( wire213  &  n_n1423 ) | ( nv983  &  wire35007 ) | ( n_n1423  &  wire35007 ) ;
 assign wire35375 = ( pi17  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire35377 = ( wire213  &  n_n1491 ) | ( wire361  &  wire35048 ) | ( n_n1491  &  wire35048 ) ;
 assign wire35378 = ( nv963  &  wire2061 ) | ( n_n1219  &  wire2061 ) | ( nv963  &  wire35048 ) | ( n_n1219  &  wire35048 ) ;
 assign wire35379 = ( (~ pi17)  &  pi19  &  pi16  &  pi15 ) ;
 assign wire35380 = ( wire213  &  n_n1555 ) | ( wire361  &  wire35065 ) | ( n_n1555  &  wire35065 ) ;
 assign wire35381 = ( nv942  &  wire1416 ) | ( n_n1229  &  wire1416 ) | ( nv942  &  wire35065 ) | ( n_n1229  &  wire35065 ) ;
 assign wire35382 = ( (~ pi17)  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire35383 = ( pi17  &  (~ pi16)  &  (~ ni29)  &  wire180 ) ;
 assign wire35384 = ( pi20  &  (~ pi16)  &  (~ ni29)  &  wire153 ) ;
 assign wire35386 = ( (~ pi17)  &  (~ pi16)  &  (~ ni29)  &  wire182 ) ;
 assign wire35388 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire35389 = ( n_n1247  &  n_n1111 ) | ( n_n1111  &  wire361 ) ;
 assign wire35390 = ( n_n1649  &  n_n1111 ) | ( n_n1111  &  wire6746 ) | ( n_n1111  &  wire29449 ) ;
 assign wire35391 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire35392 = ( (~ pi17)  &  (~ pi16)  &  wire182 ) ;
 assign wire35393 = ( wire361  &  n_n1119 ) | ( n_n1119  &  wire1516 ) | ( n_n1119  &  wire35156 ) ;
 assign wire35394 = ( n_n1119  &  n_n1259 ) | ( n_n1119  &  wire6667 ) | ( n_n1119  &  wire29466 ) ;
 assign wire35395 = ( (~ pi17)  &  pi19  &  (~ pi16) ) ;
 assign wire35396 = ( wire213  &  n_n1783 ) | ( wire361  &  wire35169 ) | ( n_n1783  &  wire35169 ) ;
 assign wire35397 = ( nv873  &  wire1493 ) | ( n_n1269  &  wire1493 ) | ( nv873  &  wire35169 ) | ( n_n1269  &  wire35169 ) ;
 assign wire35398 = ( wire1440 ) | ( (~ pi16)  &  wire157  &  wire328 ) ;
 assign wire35399 = ( wire35398 ) | ( wire302  &  n_n1253  &  wire617 ) ;
 assign wire35402 = ( wire1431 ) | ( wire1433 ) | ( n_n1255  &  wire35388 ) ;
 assign wire35403 = ( wire1434 ) | ( wire1442 ) | ( wire35399 ) ;
 assign wire35406 = ( wire1432 ) | ( wire1438 ) | ( wire35402 ) | ( wire35403 ) ;
 assign wire35407 = ( wire35406 ) | ( (~ pi16)  &  wire971 ) ;
 assign wire35408 = ( wire1262 ) | ( wire35389  &  wire35391 ) | ( wire35390  &  wire35391 ) ;
 assign wire35411 = ( wire1367 ) | ( wire157  &  wire226  &  wire328 ) ;
 assign wire35412 = ( wire35411 ) | ( wire272  &  wire226  &  wire853 ) ;
 assign wire35414 = ( wire1357 ) | ( wire1362 ) | ( wire35412 ) ;
 assign wire35416 = ( wire1361 ) | ( pi16  &  pi15  &  wire995 ) ;
 assign wire35418 = ( wire1358 ) | ( wire1360 ) | ( wire35416 ) ;
 assign wire35419 = ( wire1364 ) | ( wire1371 ) | ( wire35414 ) ;
 assign wire35421 = ( wire35418 ) | ( wire35419 ) | ( wire226  &  wire970 ) ;
 assign wire35424 = ( wire1363 ) | ( wire1365 ) | ( wire1366 ) | ( wire35421 ) ;
 assign wire35425 = ( wire35424 ) | ( pi15  &  n_n1277 ) ;
 assign wire35426 = ( (~ pi17)  &  pi19  &  pi21  &  pi20 ) ;
 assign wire35427 = ( pi16  &  (~ pi15)  &  wire35426 ) ;
 assign wire35428 = ( pi17  &  (~ pi19)  &  pi16  &  (~ pi15) ) ;
 assign wire35429 = ( pi16  &  (~ pi15)  &  wire381 ) ;
 assign wire35430 = ( pi16  &  (~ pi15)  &  wire272 ) ;
 assign wire35431 = ( (~ pi17)  &  pi16  &  (~ pi15)  &  wire182 ) ;
 assign wire35433 = ( pi17  &  (~ pi19)  &  (~ pi16) ) ;
 assign wire35434 = ( (~ pi17)  &  pi19  &  pi20  &  (~ pi16) ) ;
 assign wire35435 = ( wire272  &  (~ pi16) ) ;
 assign wire35437 = ( wire1238 ) | ( wire1254 ) | ( (~ pi16)  &  wire328 ) ;
 assign wire35439 = ( wire1233 ) | ( wire211  &  wire698  &  n_n1335 ) ;
 assign wire35440 = ( wire1235 ) | ( wire35276  &  wire35435 ) | ( wire35277  &  wire35435 ) ;
 assign wire35443 = ( wire1263 ) | ( wire1251 ) | ( wire35437 ) | ( wire35439 ) ;
 assign wire35445 = ( wire1232 ) | ( wire698  &  n_n1173 ) ;
 assign wire35446 = ( wire1236 ) | ( wire1240 ) | ( wire35440 ) | ( wire35443 ) ;
 assign wire35448 = ( wire1223 ) | ( pi16  &  (~ pi15)  &  wire328 ) ;
 assign wire35449 = ( wire35448 ) | ( wire35186  &  wire35430 ) | ( wire35187  &  wire35430 ) ;
 assign wire35450 = ( wire35449 ) | ( pi16  &  (~ pi15)  &  wire758 ) ;
 assign wire35452 = ( wire1214 ) | ( wire1216 ) | ( wire35450 ) ;
 assign wire35454 = ( wire1218 ) | ( wire35452 ) | ( wire258  &  wire997 ) ;
 assign wire35456 = ( wire1215 ) | ( wire35454 ) | ( wire258  &  wire972 ) ;
 assign wire35458 = ( wire1176 ) | ( wire289  &  wire226  &  wire328 ) ;
 assign wire35461 = ( wire1166 ) | ( wire1168 ) | ( wire1169 ) | ( wire35458 ) ;
 assign wire35464 = ( wire1170 ) | ( wire1172 ) | ( wire1175 ) | ( wire35461 ) ;
 assign wire35466 = ( wire1167 ) | ( wire35464 ) | ( wire970  &  wire35038 ) ;
 assign wire35469 = ( wire1174 ) | ( wire1191 ) | ( wire1202 ) | ( wire35466 ) ;
 assign wire35470 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  pi15 ) ;
 assign wire35471 = ( wire35470  &  wire309 ) ;
 assign wire35473 = ( pi21  &  pi20  &  pi15  &  wire456 ) ;
 assign wire35474 = ( pi21  &  pi22  &  pi20  &  pi15 ) ;
 assign wire35475 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire35474 ) ;
 assign wire35477 = ( (~ pi25)  &  pi15  &  wire456 ) ;
 assign wire35479 = ( pi25  &  pi15  &  wire456 ) ;
 assign wire35481 = ( pi20  &  pi15  &  wire456 ) ;
 assign wire35482 = ( wire700 ) | ( pi20  &  wire308 ) | ( pi20  &  wire1380 ) ;
 assign wire35485 = ( wire561 ) | ( wire562 ) | ( wire563 ) | ( wire35482 ) ;
 assign wire35487 = ( pi17  &  (~ pi19)  &  pi16  &  pi15 ) ;
 assign wire35488 = ( pi17  &  (~ pi16)  &  pi15  &  wire152 ) ;
 assign wire35489 = ( pi17  &  (~ pi16)  &  pi15  &  wire152 ) ;
 assign wire35490 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  pi15 ) ;
 assign wire35491 = ( pi17  &  pi19  &  (~ pi16)  &  pi15 ) ;
 assign wire35492 = ( (~ pi17)  &  pi19  &  wire309 ) ;
 assign wire35493 = ( (~ pi17)  &  pi19  &  pi21  &  pi20 ) ;
 assign wire35494 = ( (~ pi17)  &  pi19  &  wire189 ) ;
 assign wire35495 = ( (~ pi17)  &  pi19  &  pi20 ) ;
 assign wire35496 = ( (~ pi17)  &  pi19  &  (~ pi25) ) ;
 assign wire35497 = ( (~ pi17)  &  (~ pi19)  &  (~ pi25) ) ;
 assign wire35498 = ( wire1322 ) | ( wire191  &  wire309  &  wire259 ) ;
 assign wire35500 = ( n_n1253  &  wire35493 ) | ( n_n1255  &  wire35495 ) ;
 assign wire35502 = ( wire568 ) | ( wire629 ) | ( wire35498 ) | ( wire35500 ) ;
 assign wire35504 = ( wire570 ) | ( n_n1119  &  wire35496 ) ;
 assign wire35505 = ( wire624 ) | ( wire1493  &  wire35497 ) | ( wire35169  &  wire35497 ) ;
 assign wire35506 = ( wire35502 ) | ( wire35504 ) | ( n_n1263  &  wire817 ) ;
 assign wire35507 = ( wire35505 ) | ( wire171  &  wire1454 ) | ( wire171  &  wire35097 ) ;
 assign wire35510 = ( pi15  &  (~ pi16) ) ;
 assign wire35511 = ( (~ pi17)  &  pi19  &  wire309 ) ;
 assign wire35512 = ( (~ pi17)  &  pi19  &  pi21  &  pi20 ) ;
 assign wire35514 = ( (~ pi17)  &  pi19  &  pi20 ) ;
 assign wire35515 = ( wire1322 ) | ( wire191  &  wire309  &  wire259 ) ;
 assign wire35516 = ( wire35515 ) | ( wire308  &  wire35514 ) | ( wire1984  &  wire35514 ) ;
 assign wire35518 = ( wire651 ) | ( wire35088 ) | ( nv952  &  wire35076 ) ;
 assign wire35519 = ( wire709 ) | ( wire35516 ) | ( nv952  &  wire487 ) ;
 assign wire35521 = ( wire710 ) | ( wire35518 ) | ( wire35519 ) ;
 assign wire35522 = ( wire35521 ) | ( wire1027  &  wire35380 ) | ( wire1027  &  wire35381 ) ;
 assign wire35525 = ( (~ pi17)  &  pi19  &  pi16  &  wire309 ) ;
 assign wire35526 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire35527 = ( pi21  &  pi20  &  wire35526 ) ;
 assign wire35528 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire35531 = ( (~ pi17)  &  pi19  &  pi20  &  pi16 ) ;
 assign wire35532 = ( (~ pi17)  &  pi19  &  pi25  &  pi16 ) ;
 assign wire35533 = ( (~ pi17)  &  (~ pi19)  &  pi25  &  pi16 ) ;
 assign wire35535 = ( (~ pi17)  &  pi19  &  pi16 ) ;
 assign wire35536 = ( pi17  &  (~ pi19)  &  pi16  &  wire309 ) ;
 assign wire35537 = ( pi21  &  pi20  &  wire593 ) ;
 assign wire35539 = ( pi17  &  (~ pi19)  &  (~ pi25)  &  pi16 ) ;
 assign wire35540 = ( pi17  &  (~ pi19)  &  pi20  &  pi16 ) ;
 assign wire35541 = ( pi20  &  pi16  &  (~ ni29)  &  wire153 ) ;
 assign wire35542 = ( pi17  &  (~ pi19)  &  pi25  &  pi16 ) ;
 assign wire35544 = ( wire982 ) | ( pi16  &  wire1322 ) ;
 assign wire35545 = ( wire932 ) | ( wire967 ) | ( wire35544 ) ;
 assign wire35547 = ( wire956 ) | ( wire35545 ) | ( wire257  &  wire626 ) ;
 assign wire35549 = ( wire969 ) | ( wire35547 ) | ( pi16  &  wire758 ) ;
 assign wire35553 = ( wire888 ) | ( wire939 ) | ( wire955 ) ;
 assign wire35554 = ( wire823 ) | ( wire825 ) | ( wire938 ) | ( wire35549 ) ;
 assign wire35557 = ( wire879 ) | ( wire925 ) | ( wire35554 ) ;
 assign wire35559 = ( wire944 ) | ( wire945 ) | ( wire35553 ) | ( wire35557 ) ;
 assign wire35562 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire309 ) ;
 assign wire35563 = ( pi21  &  pi20  &  wire456 ) ;
 assign wire35564 = ( pi17  &  (~ pi19)  &  (~ pi16)  &  wire189 ) ;
 assign wire35565 = ( pi17  &  (~ pi19)  &  pi25  &  (~ pi16) ) ;
 assign wire35566 = ( pi17  &  (~ pi19)  &  pi20  &  (~ pi16) ) ;
 assign wire35567 = ( pi17  &  (~ pi19)  &  (~ pi25)  &  (~ pi16) ) ;
 assign wire35568 = ( (~ pi17)  &  (~ pi19)  &  (~ pi25) ) ;
 assign wire35569 = ( (~ pi17)  &  pi19  &  wire309 ) ;
 assign wire35570 = ( (~ pi17)  &  pi19  &  pi21  &  pi20 ) ;
 assign wire35571 = ( (~ pi17)  &  pi19  &  wire189 ) ;
 assign wire35572 = ( (~ pi17)  &  pi19  &  pi25 ) ;
 assign wire35573 = ( (~ pi17)  &  pi19  &  (~ pi25) ) ;
 assign wire35574 = ( (~ pi17)  &  pi19  &  pi20 ) ;
 assign wire35575 = ( (~ pi20)  &  (~ pi25)  &  wire153 ) ;
 assign wire35577 = ( wire1159 ) | ( wire1160 ) | ( wire228  &  n_n1347 ) ;
 assign wire35579 = ( wire1141 ) | ( n_n1335  &  wire35570 ) ;
 assign wire35581 = ( wire1155 ) | ( wire35577 ) | ( wire487  &  wire785 ) ;
 assign wire35584 = ( wire1154 ) | ( wire1157 ) | ( wire35579 ) | ( wire35581 ) ;
 assign wire35585 = ( wire1143 ) | ( wire1156 ) | ( wire1164 ) ;
 assign wire35587 = ( wire1145 ) | ( n_n1173  &  wire35573 ) ;
 assign wire35588 = ( wire35584 ) | ( wire35585 ) | ( wire35587 ) ;
 assign wire35589 = ( wire1136 ) | ( wire309  &  wire456  &  wire259 ) ;
 assign wire35590 = ( wire35589 ) | ( wire295  &  wire1720 ) | ( wire295  &  wire35320 ) ;
 assign wire35593 = ( wire1004 ) | ( wire1042 ) | ( wire1137 ) | ( wire35590 ) ;
 assign wire35595 = ( wire1001 ) | ( wire35593 ) | ( n_n2176  &  wire35564 ) ;
 assign wire35597 = ( wire1040 ) | ( wire1054 ) | ( wire35595 ) ;
 assign wire35599 = ( wire551 ) | ( wire416  &  wire1109 ) | ( wire1109  &  wire35488 ) ;
 assign wire35600 = ( wire35599 ) | ( wire485  &  wire1376 ) | ( wire485  &  wire35028 ) ;
 assign wire35602 = ( n_n1241  &  wire35473 ) | ( n_n1243  &  wire35481 ) ;
 assign wire35603 = ( wire552 ) | ( wire35600 ) | ( wire416  &  wire853 ) ;
 assign wire35606 = ( wire542 ) | ( wire550 ) | ( wire35602 ) | ( wire35603 ) ;
 assign wire35608 = ( wire544 ) | ( wire35606 ) | ( n_n1111  &  wire35477 ) ;
 assign wire35609 = ( wire35608 ) | ( wire35389  &  wire35479 ) | ( wire35390  &  wire35479 ) ;
 assign wire35611 = ( wire548 ) | ( wire35609 ) | ( n_n1813  &  wire35510 ) ;
 assign wire35613 = ( wire558 ) | ( wire35611 ) | ( (~ pi15)  &  n_n2483 ) ;
 assign wire35614 = ( (~ ni9)  &  (~ ni10)  &  (~ ni8)  &  wire175 ) ;
 assign wire35615 = ( (~ ni9)  &  (~ ni8)  &  (~ wire289) ) ;
 assign wire35616 = ( wire538 ) | ( wire559  &  wire35614 ) | ( wire35613  &  wire35614 ) ;
 assign wire35617 = ( wire541 ) | ( wire833  &  wire559 ) | ( wire833  &  wire35613 ) ;
 assign wire35619 = ( (~ ni2)  &  (~ ni3)  &  (~ wire1201)  &  (~ wire35469) ) ;
 assign wire35620 = ( (~ ni2)  &  (~ ni3)  &  ni7 ) ;
 assign wire35621 = ( wire521 ) | ( (~ wire1201)  &  (~ wire35469)  &  wire35620 ) ;
 assign wire35623 = ( ni3  &  ni31  &  ni30 ) ;
 assign wire35626 = ( ni4  &  (~ ni6) ) | ( (~ ni5)  &  (~ ni6) ) ;
 assign wire35628 = ( ni3  &  (~ ni31)  &  (~ ni6) ) ;
 assign wire35629 = ( (~ n_n806)  &  (~ ni3) ) ;
 assign wire35631 = ( ni3  &  ni31  &  ni6 ) | ( ni3  &  (~ ni31)  &  wire35626 ) ;
 assign wire35633 = ( wire497 ) | ( wire511 ) | ( wire35631 ) ;
 assign wire35634 = ( wire35633 ) | ( (~ ni3)  &  ni6  &  (~ n_n806) ) ;
 assign wire35636 = ( ni9  &  (~ ni7) ) | ( (~ ni10)  &  (~ ni7) ) ;
 assign wire35638 = ( ni9  &  (~ ni7) ) | ( ni10  &  (~ ni7) ) ;
 assign wire35640 = ( wire479 ) | ( (~ ni3)  &  (~ ni7)  &  (~ ni8) ) ;
 assign wire35641 = ( pi24  &  (~ ni3)  &  wire35636 ) | ( (~ pi24)  &  (~ ni3)  &  wire35638 ) ;
 assign wire35643 = ( ni4  &  (~ ni36) ) ;
 assign wire35645 = ( ni4  &  ni33  &  ni31 ) ;
 assign wire35648 = ( (~ n_n9245)  &  wire35645 ) | ( ni31  &  (~ n_n9245)  &  wire35643 ) ;
 assign wire35652 = ( (~ ni2)  &  ni3  &  (~ ni6) ) ;
 assign wire35653 = ( (~ ni41)  &  (~ ni33)  &  ni31  &  ni30 ) ;
 assign wire35655 = ( ni32  &  ni5  &  wire35652  &  wire35653 ) ;
 assign wire35656 = ( (~ wire494)  &  (~ wire35640)  &  (~ wire35641)  &  wire35655 ) ;
 assign wire35658 = ( (~ ni2)  &  ni3  &  (~ ni6) ) ;
 assign wire35659 = ( (~ ni33)  &  (~ ni32)  &  ni31  &  ni30 ) ;
 assign wire35661 = ( (~ ni36)  &  ni5  &  wire35658  &  wire35659 ) ;
 assign wire35662 = ( (~ wire494)  &  (~ wire35640)  &  (~ wire35641)  &  wire35661 ) ;
 assign wire35663 = ( (~ ni33)  &  (~ ni5) ) | ( (~ ni31)  &  (~ ni5) ) ;
 assign wire35665 = ( ni31  &  (~ ni30)  &  (~ wire425)  &  wire35663 ) ;
 assign wire35666 = ( (~ wire494)  &  (~ wire35640)  &  (~ wire35641)  &  wire35665 ) ;
 assign wire35667 = ( wire830  &  (~ wire494)  &  (~ wire35640)  &  (~ wire35641) ) ;
 assign wire35670 = ( wire430 ) | ( (~ n_n424)  &  wire35656 ) | ( (~ n_n424)  &  wire35667 ) ;
 assign wire35671 = ( pi24  &  pi23 ) ;
 assign wire35673 = ( (~ ni2)  &  (~ ni4)  &  ni3  &  ni6 ) ;
 assign wire35675 = ( (~ ni2)  &  (~ ni4)  &  ni3  &  (~ ni6) ) ;
 assign wire35678 = ( (~ ni2)  &  ni3  &  ni6 ) ;
 assign wire35679 = ( (~ ni2)  &  ni11  &  (~ ni3) ) ;
 assign wire35680 = ( (~ ni2)  &  ni11  &  (~ ni3) ) ;
 assign wire35681 = ( wire410 ) | ( wire936  &  wire35673 ) ;
 assign wire35682 = ( n_n13958  &  (~ ni33)  &  wire1029 ) | ( n_n13958  &  (~ wire930)  &  wire1029 ) ;
 assign wire35683 = ( (~ wire725)  &  wire35678 ) | ( wire389  &  wire35679 ) ;
 assign wire35684 = ( wire830  &  wire478 ) | ( wire155  &  wire35680 ) ;
 assign wire35685 = ( (~ ni31)  &  wire830 ) | ( (~ ni30)  &  wire830 ) | ( ni5  &  wire830 ) ;
 assign wire35690 = ( wire283 ) | ( wire285 ) | ( wire362 ) | ( wire35681 ) ;
 assign wire35691 = ( wire35682 ) | ( wire35683 ) | ( wire35684 ) | ( wire35685 ) ;
 assign wire35694 = ( pi25  &  (~ ni9)  &  (~ ni7)  &  (~ ni8) ) ;
 assign wire35695 = ( (~ ni2)  &  (~ ni3)  &  (~ ni33) ) | ( (~ ni2)  &  (~ ni3)  &  (~ ni29) ) ;


endmodule

