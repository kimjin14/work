`define CONFIG_SIZE 787512
