module add4 (a,b,z);
	input [3:0] a;
	input [3:0] b;
	output [4:0] z;

	assign z = a+b;
	
endmodule
