module misex3 (
	a, b, c, d, e, f, g, h, 
	i, j, k, l, m, n, r2, s2, p2, q2, 
	t2, u2, j2, k2, h2, i2, n2, o2, l2, m2);

input a;
input b;
input c;
input d;
input e;
input f;
input g;
input h;
input i;
input j;
input k;
input l;
input m;
input n;
output r2;
output s2;
output p2;
output q2;
output t2;
output u2;
output j2;
output k2;
output h2;
output i2;
output n2;
output o2;
output l2;
output m2;
wire n_n1089;
wire n_n842;
wire n_n840;
wire n_n1161;
wire n_n1207;
wire n_n711;
wire n_n713;
wire n_n709;
wire n_n1188;
wire n_n886;
wire wire38;
wire wire46;
wire wire53;
wire wire75;
wire wire84;
wire wire148;
wire wire153;
wire wire172;
wire wire175;
wire wire202;
wire wire224;
wire wire229;
wire wire233;
wire wire393;
wire n_n1177;
wire n_n1165;
wire n_n904;
wire n_n626;
wire n_n671;
wire n_n1101;
wire n_n1229;
wire n_n1193;
wire n_n1344;
wire wire22;
wire wire31;
wire wire45;
wire wire54;
wire wire71;
wire wire101;
wire wire138;
wire wire195;
wire wire232;
wire wire258;
wire wire371;
wire n_n1217;
wire n_n1201;
wire n_n1220;
wire n_n920;
wire n_n918;
wire wire15;
wire wire58;
wire wire82;
wire wire98;
wire wire130;
wire wire220;
wire wire228;
wire wire265;
wire wire390;
wire wire417;
wire n_n1187;
wire n_n996;
wire n_n1155;
wire n_n1171;
wire n_n698;
wire n_n617;
wire n_n730;
wire n_n618;
wire n_n857;
wire n_n933;
wire n_n821;
wire n_n700;
wire n_n824;
wire n_n1792;
wire wire29;
wire wire30;
wire wire34;
wire wire179;
wire wire210;
wire wire255;
wire wire291;
wire wire309;
wire wire380;
wire n_n1069;
wire n_n1104;
wire n_n1203;
wire n_n876;
wire n_n1166;
wire n_n1425;
wire wire74;
wire wire76;
wire wire92;
wire wire112;
wire wire120;
wire wire183;
wire wire184;
wire wire196;
wire wire223;
wire wire230;
wire wire256;
wire n_n841;
wire n_n893;
wire n_n1194;
wire n_n1495;
wire wire33;
wire wire93;
wire wire106;
wire wire156;
wire wire203;
wire wire219;
wire n_n1138;
wire n_n1159;
wire n_n2507;
wire n_n1080;
wire n_n2494;
wire wire116;
wire wire199;
wire wire319;
wire n_n1190;
wire n_n1202;
wire n_n1039;
wire n_n2602;
wire n_n2511;
wire n_n2493;
wire wire157;
wire wire267;
wire n_n1142;
wire n_n949;
wire n_n761;
wire n_n1231;
wire n_n1261;
wire n_n997;
wire n_n1874;
wire wire44;
wire wire57;
wire wire94;
wire wire108;
wire wire200;
wire wire254;
wire wire379;
wire wire387;
wire wire407;
wire wire413;
wire n_n872;
wire n_n838;
wire n_n977;
wire n_n1252;
wire n_n1920;
wire n_n1919;
wire n_n987;
wire n_n1210;
wire n_n1939;
wire n_n988;
wire wire39;
wire wire77;
wire wire89;
wire wire111;
wire wire117;
wire wire135;
wire wire159;
wire wire160;
wire wire164;
wire wire165;
wire wire167;
wire wire386;
wire n_n1022;
wire n_n1573;
wire n_n820;
wire n_n1264;
wire n_n3060;
wire wire14;
wire wire40;
wire wire113;
wire wire208;
wire wire351;
wire n_n1085;
wire n_n1036;
wire n_n1053;
wire n_n619;
wire n_n1653;
wire n_n816;
wire wire21;
wire wire36;
wire wire50;
wire wire207;
wire wire209;
wire wire290;
wire wire315;
wire wire320;
wire n_n1219;
wire n_n2023;
wire wire114;
wire wire127;
wire wire146;
wire wire222;
wire wire263;
wire wire268;
wire wire404;
wire n_n971;
wire n_n1204;
wire n_n973;
wire n_n1072;
wire n_n1028;
wire wire37;
wire wire68;
wire wire384;
wire n_n1160;
wire n_n662;
wire wire282;
wire wire373;
wire n_n1180;
wire n_n1196;
wire wire103;
wire wire204;
wire wire227;
wire wire273;
wire n_n1121;
wire n_n1164;
wire n_n1222;
wire n_n1095;
wire n_n975;
wire wire70;
wire wire221;
wire wire234;
wire wire283;
wire wire285;
wire wire286;
wire wire301;
wire n_n1148;
wire n_n1137;
wire n_n1191;
wire n_n1195;
wire n_n1133;
wire n_n861;
wire n_n1082;
wire n_n1260;
wire n_n819;
wire n_n1131;
wire wire79;
wire wire122;
wire wire158;
wire wire170;
wire wire194;
wire n_n1243;
wire n_n1227;
wire n_n1091;
wire wire95;
wire wire132;
wire wire226;
wire wire395;
wire n_n818;
wire n_n529;
wire n_n670;
wire wire23;
wire wire59;
wire wire96;
wire wire134;
wire wire169;
wire wire398;
wire n_n387;
wire wire72;
wire wire211;
wire wire231;
wire wire137;
wire n_n1118;
wire n_n1216;
wire n_n1056;
wire wire189;
wire n_n868;
wire n_n823;
wire wire259;
wire n_n989;
wire n_n1094;
wire wire249;
wire n_n628;
wire n_n623;
wire wire128;
wire wire396;
wire n_n992;
wire wire118;
wire n_n1146;
wire wire121;
wire n_n1228;
wire n_n1116;
wire n_n1215;
wire n_n1233;
wire n_n940;
wire n_n942;
wire n_n765;
wire n_n822;
wire n_n859;
wire n_n1253;
wire wire248;
wire wire314;
wire wire55;
wire wire149;
wire wire18;
wire wire20;
wire n_n874;
wire n_n605;
wire n_n1084;
wire n_n766;
wire n_n875;
wire n_n871;
wire wire90;
wire n_n235;
wire n_n2572;
wire n_n2953;
wire n_n1167;
wire n_n1083;
wire n_n1189;
wire n_n978;
wire n_n703;
wire n_n864;
wire n_n817;
wire wire197;
wire wire161;
wire wire305;
wire wire399;
wire wire414;
wire wire369;
wire n_n2660;
wire n_n982;
wire wire47;
wire n_n1249;
wire n_n919;
wire n_n694;
wire n_n844;
wire n_n912;
wire wire35;
wire n_n2026;
wire wire56;
wire wire142;
wire wire188;
wire wire216;
wire wire260;
wire n_n747;
wire wire181;
wire wire104;
wire wire293;
wire n_n825;
wire wire43;
wire wire24;
wire wire49;
wire wire109;
wire wire206;
wire wire105;
wire wire152;
wire wire299;
wire wire388;
wire wire65;
wire wire162;
wire wire198;
wire wire377;
wire wire385;
wire wire16;
wire wire25;
wire wire32;
wire wire41;
wire wire60;
wire wire69;
wire wire80;
wire wire81;
wire wire85;
wire wire190;
wire wire115;
wire wire368;
wire wire42;
wire wire61;
wire wire63;
wire wire66;
wire wire140;
wire wire150;
wire wire163;
wire wire173;
wire wire177;
wire wire178;
wire wire180;
wire wire252;
wire wire253;
wire wire269;
wire wire271;
wire wire272;
wire wire274;
wire wire275;
wire wire276;
wire wire277;
wire wire278;
wire wire280;
wire wire281;
wire wire307;
wire wire316;
wire wire317;
wire wire318;
wire wire321;
wire wire322;
wire wire328;
wire wire329;
wire wire330;
wire wire331;
wire wire333;
wire wire334;
wire wire336;
wire wire337;
wire wire338;
wire wire339;
wire wire340;
wire wire341;
wire wire342;
wire wire345;
wire wire347;
wire wire352;
wire wire353;
wire wire354;
wire wire355;
wire wire357;
wire wire359;
wire wire362;
wire wire389;
wire wire424;
wire wire425;
wire wire429;
wire wire430;
wire wire431;
wire wire432;
wire wire433;
wire wire434;
wire wire435;
wire wire440;
wire wire441;
wire wire442;
wire wire443;
wire wire444;
wire wire445;
wire wire446;
wire wire447;
wire wire448;
wire wire449;
wire wire450;
wire wire451;
wire wire452;
wire wire453;
wire wire454;
wire wire455;
wire wire456;
wire wire457;
wire wire458;
wire wire459;
wire wire460;
wire wire461;
wire wire463;
wire wire464;
wire wire465;
wire wire466;
wire wire467;
wire wire468;
wire wire469;
wire wire470;
wire wire471;
wire wire480;
wire wire481;
wire wire482;
wire wire483;
wire wire484;
wire wire485;
wire wire486;
wire wire487;
wire wire488;
wire wire489;
wire wire490;
wire wire491;
wire wire492;
wire wire493;
wire wire494;
wire wire495;
wire wire496;
wire wire499;
wire wire500;
wire wire501;
wire wire502;
wire wire503;
wire wire504;
wire wire505;
wire wire508;
wire wire509;
wire wire510;
wire wire511;
wire wire512;
wire wire513;
wire wire516;
wire wire517;
wire wire520;
wire wire521;
wire wire522;
wire wire523;
wire wire527;
wire wire528;
wire wire532;
wire wire533;
wire wire534;
wire wire535;
wire wire536;
wire wire537;
wire wire539;
wire wire540;
wire wire541;
wire wire542;
wire wire543;
wire wire544;
wire wire545;
wire wire546;
wire wire547;
wire wire548;
wire wire549;
wire wire550;
wire wire551;
wire wire552;
wire wire554;
wire wire565;
wire wire566;
wire wire567;
wire wire568;
wire wire569;
wire wire570;
wire wire571;
wire wire572;
wire wire573;
wire wire575;
wire wire576;
wire wire577;
wire wire579;
wire wire580;
wire wire581;
wire wire583;
wire wire585;
wire wire586;
wire wire587;
wire wire588;
wire wire590;
wire wire593;
wire wire594;
wire wire598;
wire wire610;
wire wire611;
wire wire617;
wire wire618;
wire wire619;
wire wire626;
wire wire627;
wire wire628;
wire wire629;
wire wire630;
wire wire631;
wire wire632;
wire wire633;
wire wire635;
wire wire641;
wire wire642;
wire wire643;
wire wire644;
wire wire645;
wire wire646;
wire wire647;
wire wire649;
wire wire650;
wire wire651;
wire wire652;
wire wire653;
wire wire655;
wire wire657;
wire wire658;
wire wire661;
wire wire663;
wire wire664;
wire wire670;
wire wire671;
wire wire672;
wire wire679;
wire wire680;
wire wire681;
wire wire682;
wire wire683;
wire wire684;
wire wire699;
wire wire700;
wire wire701;
wire wire702;
wire wire703;
wire wire704;
wire wire708;
wire wire709;
wire wire713;
wire wire716;
wire wire717;
wire wire718;
wire wire719;
wire wire724;
wire wire725;
wire wire726;
wire wire727;
wire wire729;
wire wire731;
wire wire732;
wire wire736;
wire wire739;
wire wire743;
wire wire745;
wire wire749;
wire wire750;
wire wire751;
wire wire753;
wire wire754;
wire wire762;
wire wire765;
wire wire766;
wire wire767;
wire wire775;
wire wire776;
wire wire777;
wire wire780;
wire wire781;
wire wire782;
wire wire783;
wire wire784;
wire wire785;
wire wire786;
wire wire787;
wire wire788;
wire wire789;
wire wire790;
wire wire791;
wire wire796;
wire wire797;
wire wire798;
wire wire799;
wire wire802;
wire wire808;
wire wire809;
wire wire810;
wire wire811;
wire wire812;
wire wire813;
wire wire814;
wire wire815;
wire wire816;
wire wire817;
wire wire818;
wire wire821;
wire wire822;
wire wire823;
wire wire826;
wire wire827;
wire wire828;
wire wire829;
wire wire830;
wire wire831;
wire wire832;
wire wire833;
wire wire834;
wire wire835;
wire wire836;
wire wire837;
wire wire841;
wire wire843;
wire wire845;
wire wire849;
wire wire850;
wire wire853;
wire wire854;
wire wire858;
wire wire859;
wire wire860;
wire wire864;
wire wire869;
wire wire871;
wire wire875;
wire wire879;
wire wire880;
wire wire884;
wire wire886;
wire wire895;
wire wire898;
wire wire900;
wire wire901;
wire wire902;
wire wire903;
wire wire904;
wire wire906;
wire wire907;
wire wire908;
wire wire909;
wire wire911;
wire wire912;
wire wire914;
wire wire923;
wire wire924;
wire wire925;
wire wire926;
wire wire927;
wire wire928;
wire wire929;
wire wire931;
wire wire932;
wire wire934;
wire wire935;
wire wire938;
wire wire939;
wire wire940;
wire wire941;
wire wire942;
wire wire943;
wire wire945;
wire wire948;
wire wire951;
wire wire952;
wire wire954;
wire wire960;
wire wire961;
wire wire962;
wire wire963;
wire wire965;
wire wire966;
wire wire967;
wire wire968;
wire wire969;
wire wire970;
wire wire971;
wire wire972;
wire wire973;
wire wire974;
wire wire975;
wire wire976;
wire wire977;
wire wire978;
wire wire980;
wire wire982;
wire wire983;
wire wire985;
wire wire986;
wire wire989;
wire wire990;
wire wire991;
wire wire992;
wire wire993;
wire wire994;
wire wire995;
wire wire997;
wire wire1012;
wire wire1016;
wire wire1018;
wire wire1019;
wire wire1020;
wire wire1021;
wire wire1022;
wire wire1023;
wire wire1024;
wire wire1027;
wire wire1030;
wire wire1031;
wire wire1032;
wire wire1033;
wire wire1034;
wire wire1036;
wire wire1039;
wire wire1042;
wire wire1043;
wire wire1051;
wire wire1052;
wire wire1053;
wire wire1054;
wire wire1055;
wire wire1057;
wire wire1058;
wire wire1059;
wire wire1060;
wire wire1061;
wire wire1062;
wire wire1068;
wire wire1070;
wire wire1071;
wire wire1074;
wire wire1075;
wire wire1076;
wire wire1077;
wire wire1078;
wire wire1079;
wire wire1080;
wire wire1081;
wire wire1082;
wire wire1083;
wire wire1084;
wire wire1096;
wire wire1100;
wire wire1102;
wire wire1106;
wire wire1110;
wire wire1112;
wire wire1113;
wire wire1116;
wire wire1122;
wire wire1123;
wire wire1124;
wire wire1126;
wire wire1128;
wire wire1129;
wire wire1130;
wire wire1131;
wire wire1135;
wire wire1137;
wire wire1138;
wire wire1139;
wire wire1140;
wire wire1141;
wire wire1145;
wire wire1147;
wire wire1148;
wire wire1155;
wire wire1156;
wire wire1157;
wire wire1158;
wire wire1161;
wire wire1162;
wire wire1163;
wire wire1166;
wire wire1167;
wire wire1168;
wire wire1169;
wire wire1170;
wire wire1171;
wire wire1172;
wire wire1173;
wire wire1175;
wire wire1176;
wire wire1185;
wire wire1186;
wire wire1187;
wire wire1188;
wire wire1189;
wire wire1192;
wire wire1193;
wire wire1194;
wire wire1195;
wire wire1196;
wire wire1197;
wire wire1198;
wire wire1200;
wire wire1205;
wire wire5088;
wire wire5091;
wire wire5093;
wire wire5094;
wire wire5095;
wire wire5098;
wire wire5099;
wire wire5108;
wire wire5116;
wire wire5117;
wire wire5120;
wire wire5124;
wire wire5125;
wire wire5126;
wire wire5127;
wire wire5128;
wire wire5129;
wire wire5130;
wire wire5136;
wire wire5137;
wire wire5139;
wire wire5140;
wire wire5144;
wire wire5146;
wire wire5156;
wire wire5159;
wire wire5160;
wire wire5161;
wire wire5162;
wire wire5163;
wire wire5169;
wire wire5170;
wire wire5171;
wire wire5172;
wire wire5175;
wire wire5176;
wire wire5177;
wire wire5179;
wire wire5181;
wire wire5183;
wire wire5184;
wire wire5187;
wire wire5188;
wire wire5190;
wire wire5191;
wire wire5192;
wire wire5194;
wire wire5197;
wire wire5198;
wire wire5199;
wire wire5201;
wire wire5204;
wire wire5205;
wire wire5207;
wire wire5208;
wire wire5209;
wire wire5210;
wire wire5213;
wire wire5215;
wire wire5216;
wire wire5220;
wire wire5226;
wire wire5227;
wire wire5228;
wire wire5232;
wire wire5233;
wire wire5234;
wire wire5237;
wire wire5238;
wire wire5241;
wire wire5242;
wire wire5243;
wire wire5244;
wire wire5246;
wire wire5251;
wire wire5252;
wire wire5253;
wire wire5255;
wire wire5256;
wire wire5257;
wire wire5264;
wire wire5265;
wire wire5266;
wire wire5268;
wire wire5270;
wire wire5271;
wire wire5274;
wire wire5277;
wire wire5279;
wire wire5289;
wire wire5290;
wire wire5291;
wire wire5293;
wire wire5297;
wire wire5298;
wire wire5299;
wire wire5300;
wire wire5305;
wire wire5306;
wire wire5307;
wire wire5309;
wire wire5311;
wire wire5313;
wire wire5314;
wire wire5316;
wire wire5317;
wire wire5318;
wire wire5321;
wire wire5323;
wire wire5325;
wire wire5327;
wire wire5328;
wire wire5329;
wire wire5330;
wire wire5333;
wire wire5356;
wire wire5357;
wire wire5358;
wire wire5359;
wire wire5360;
wire wire5364;
wire wire5367;
wire wire5368;
wire wire5379;
wire wire5382;
wire wire5386;
wire wire5387;
wire wire5388;
wire wire5389;
wire wire5391;
wire wire5394;
wire wire5395;
wire wire5396;
wire wire5397;
wire wire5399;
wire wire5400;
wire wire5406;
wire wire5407;
wire wire5413;
wire wire5414;
wire wire5415;
wire wire5416;
wire wire5418;
wire wire5422;
wire wire5424;
wire wire5431;
wire wire5432;
wire wire5433;
wire wire5435;
wire wire5436;
wire wire5437;
wire wire5443;
wire wire5444;
wire wire5445;
wire wire5446;
wire wire5448;
wire wire5449;
wire wire5451;
wire wire5453;
wire wire5454;
wire wire5456;
wire wire5457;
wire wire5459;
wire wire5460;
wire wire5461;
wire wire5462;
wire wire5463;
wire wire5467;
wire wire5469;
wire wire5474;
wire wire5475;
wire wire5477;
wire wire5479;
wire wire5480;
wire wire5485;
wire wire5486;
wire wire5489;
wire wire5490;
wire wire5493;
wire wire5495;
wire wire5498;
wire wire5499;
wire wire5505;
wire wire5506;
wire wire5507;
wire wire5508;
wire wire5509;
wire wire5513;
wire wire5514;
wire wire5515;
wire wire5517;
wire wire5518;
wire wire5520;
wire wire5521;
wire wire5523;
wire wire5526;
wire wire5529;
wire wire5532;
wire wire5534;
wire wire5557;
wire wire5561;
wire wire5570;
wire wire5572;
wire wire5573;
wire wire5574;
wire wire5575;
wire wire5576;
wire wire5578;
wire wire5579;
wire wire5583;
wire wire5584;
wire wire5585;
wire wire5587;
wire wire5590;
wire wire5592;
wire wire5598;
wire wire5600;
wire wire5601;
wire wire5602;
wire wire5603;
wire wire5605;
wire wire5611;
wire wire5613;
wire wire5615;
wire wire5618;
wire wire5619;
wire wire5620;
wire wire5621;
wire wire5624;
wire wire5629;
wire wire5633;
wire wire5637;
wire wire5639;
wire wire5640;
wire wire5649;
wire wire5650;
wire wire5652;
wire wire5654;
wire wire5659;
wire wire5663;
wire wire5664;
wire wire5666;
wire wire5668;
wire wire5672;
wire wire5674;
wire wire5677;
wire wire5678;
wire wire5679;
wire wire5681;
wire wire5685;
wire wire5686;
wire wire5687;
wire wire5690;
wire wire5693;
wire wire5694;
wire wire5695;
wire wire5696;
wire wire5699;
wire wire5703;
wire wire5704;
wire wire5705;
wire wire5708;
wire wire5709;
wire wire5710;
wire wire5711;
wire wire5715;
wire wire5718;
wire wire5719;
wire wire5720;
wire wire5721;
wire wire5722;
wire wire5726;
wire wire5727;
wire wire5731;
wire wire5732;
wire wire5740;
wire wire5743;
wire wire5744;
wire wire5751;
wire wire5752;
wire wire5753;
wire wire5758;
wire wire5759;
wire wire5760;
wire wire5761;
wire wire5762;
wire wire5763;
wire wire5766;
wire wire5774;
wire wire5775;
wire wire5781;
wire wire5792;
wire wire5793;
wire wire5795;
wire wire5797;
wire wire5798;
wire wire5802;
wire wire5803;
wire wire5804;
wire wire5806;
wire wire5809;
wire wire5810;
wire wire5811;
wire wire5813;
wire wire5814;
wire wire5824;
wire wire5825;
wire wire5826;
wire wire5828;
wire wire5829;
wire wire5830;
wire wire5831;
wire wire5833;
wire wire5834;
wire wire5835;
wire wire5836;
wire wire5837;
wire wire5839;
wire wire5840;
wire wire5841;
wire wire5842;
wire wire5843;
wire wire5846;
wire wire5847;
wire wire5848;
wire wire5849;
wire wire5850;
wire wire5851;
wire wire5857;
wire wire5858;
wire wire5860;
wire wire5864;
wire wire5865;
wire wire5866;
wire wire5867;
wire wire5870;
wire wire5871;
wire wire5873;
wire wire5875;
wire wire5876;
wire wire5877;
wire wire5884;
wire wire5886;
wire wire5888;
wire wire5897;
wire wire5898;
wire wire5899;
wire wire5901;
wire wire5903;
wire wire5904;
wire wire5905;
wire wire5906;
wire wire5912;
wire wire5925;
wire wire5927;
wire wire5928;
wire wire5929;
wire wire5930;
wire wire5934;
wire wire5936;
wire wire5937;
wire wire5938;
wire wire5941;
wire wire5943;
wire wire5944;
wire wire5945;
wire wire5946;
wire wire5951;
wire wire5954;
wire wire5955;
wire wire5958;
wire wire5959;
wire wire5961;
wire wire5962;
wire wire5963;
wire wire5964;
wire wire5967;
wire wire5969;
wire wire5970;
wire wire5971;
wire wire5977;
wire wire5979;
wire wire5981;
wire wire5982;
wire wire5986;
wire wire5990;
wire wire5996;
wire wire5998;
wire wire5999;
wire wire6001;
wire wire6002;
wire wire6005;
wire wire6006;
wire wire6010;
wire wire6012;
wire wire6014;
wire wire6020;
wire wire6022;
wire wire6035;
wire wire6036;
wire wire6037;
wire wire6038;
wire wire6040;
wire wire6041;
wire wire6042;
wire wire6045;
wire wire6047;
wire wire6054;
wire wire6057;
wire wire6062;
wire wire6064;
wire wire6065;
wire wire6066;
wire wire6067;
wire wire6070;
wire wire6071;
wire wire6072;
wire wire6074;
wire wire6076;
wire wire6078;
wire wire6082;
wire wire6085;
wire wire6100;
wire wire6101;
wire wire6102;
wire wire6103;
wire wire6106;
wire wire6107;
wire wire6108;
wire wire6109;
wire wire6112;
wire wire6115;
wire wire6118;
wire wire6119;
wire wire6122;
wire wire6123;
wire wire6125;
wire wire6130;
wire wire6131;
wire wire6132;
wire wire6133;
wire wire6135;
wire wire6138;
wire wire6139;
wire wire6141;
wire wire6142;
wire wire6143;
wire wire6144;
wire wire6145;
wire wire6147;
wire wire6149;
wire wire6150;
wire wire6151;
wire wire6156;
wire wire6158;
wire wire6159;
wire wire6160;
wire wire6161;
wire wire6165;
wire wire6168;
wire wire6169;
wire wire6170;
wire wire6171;
wire wire6176;
wire wire6177;
wire wire6180;
wire wire6183;
wire wire6184;
wire wire6185;
wire wire6187;
wire wire6188;
wire wire6194;
wire wire6195;
wire wire6200;
wire wire6203;
wire wire6204;
wire wire6205;
wire wire6206;
wire wire6207;
wire wire6210;
wire wire6211;
wire wire6213;
wire wire6216;
wire wire6217;
wire wire6220;
wire wire6222;
wire wire6224;
wire wire6225;
wire wire6226;
wire wire6227;
wire wire6230;
wire wire6233;
wire wire6236;
wire wire6238;
wire wire6239;
wire wire6240;
wire wire6241;
wire wire6245;
wire wire6246;
wire wire6248;
wire wire6249;
wire wire6250;
wire wire6251;
wire wire6252;
wire wire6256;
wire wire6257;
wire wire6258;
wire wire6262;
wire wire6263;
wire wire6264;
wire wire6266;
wire wire6268;
wire wire6272;
wire wire6281;
wire wire6282;
wire wire6283;
wire wire6285;
wire wire6286;
wire wire6287;
wire wire6289;
wire wire6290;
wire wire6292;
wire wire6293;
wire wire6297;
wire wire6298;
wire wire6300;
wire wire6301;
wire wire6303;
wire wire6304;
wire wire6306;
wire wire6307;
wire wire6309;
wire wire6310;
wire wire6317;
wire wire6318;
wire wire6322;
wire wire6323;
assign r2 = ( wire5098 ) | ( wire5099 ) | ( wire5139 ) | ( wire5175 ) ;
 assign s2 = ( n_n1344 ) | ( wire5264 ) | ( wire5265 ) | ( wire5268 ) ;
 assign p2 = ( wire5305 ) | ( wire5306 ) | ( wire5307 ) | ( wire5333 ) ;
 assign q2 = ( wire5399 ) | ( wire5400 ) | ( wire5448 ) | ( wire5449 ) ;
 assign t2 = ( n_n1425 ) | ( wire5518 ) | ( wire5521 ) | ( wire5523 ) ;
 assign u2 = ( n_n1495 ) | ( wire5619 ) | ( wire5620 ) | ( wire5624 ) ;
 assign j2 = ( wire5649 ) | ( wire5650 ) | ( wire5654 ) ;
 assign k2 = ( n_n2493 ) | ( wire753 ) | ( wire5668 ) | ( wire5672 ) ;
 assign h2 = ( n_n1874 ) | ( wire5722 ) | ( wire5726 ) ;
 assign i2 = ( wire5809 ) | ( wire5810 ) | ( wire5811 ) ;
 assign n2 = ( n_n1573 ) | ( wire5828 ) | ( wire5829 ) | ( wire5873 ) ;
 assign o2 = ( n_n1653 ) | ( wire5936 ) | ( wire5937 ) | ( wire5938 ) ;
 assign l2 = ( wire6303 ) | ( wire6304 ) | ( wire6306 ) ;
 assign m2 = ( n_n1939 ) | ( wire6322 ) | ( wire6323 ) ;
 assign n_n1089 = ( f  &  (~ g)  &  (~ h) ) ;
 assign n_n842 = ( b  &  (~ c)  &  d ) ;
 assign n_n840 = ( b  &  d  &  (~ e) ) ;
 assign n_n1161 = ( (~ e)  &  g  &  (~ h) ) ;
 assign n_n1207 = ( f  &  g  &  (~ h) ) ;
 assign n_n711 = ( b  &  c  &  e ) ;
 assign n_n713 = ( b  &  c  &  (~ d) ) ;
 assign n_n709 = ( b  &  (~ d)  &  e ) ;
 assign n_n1188 = ( g  &  j  &  (~ k) ) ;
 assign n_n886 = ( e  &  (~ f)  &  h ) ;
 assign wire38 = ( m  &  (~ n)  &  n_n920 ) ;
 assign wire46 = ( (~ g)  &  n_n942 ) | ( g  &  wire20 ) ;
 assign wire53 = ( (~ d)  &  e ) ;
 assign wire75 = ( (~ m)  &  n  &  n_n893 ) ;
 assign wire84 = ( i  &  k  &  (~ m)  &  n ) ;
 assign wire148 = ( i  &  l  &  m  &  (~ n) ) ;
 assign wire153 = ( wire1145 ) | ( (~ d)  &  e  &  n_n1261 ) ;
 assign wire172 = ( (~ i)  &  k  &  (~ m)  &  n ) ;
 assign wire175 = ( (~ e)  &  f  &  (~ g) ) | ( (~ e)  &  (~ f)  &  (~ g) ) ;
 assign wire202 = ( b  &  (~ c)  &  d ) | ( b  &  (~ d)  &  e ) ;
 assign wire224 = ( a  &  b  &  (~ c)  &  f ) ;
 assign wire229 = ( e  &  f  &  g ) | ( e  &  f  &  (~ g) ) ;
 assign wire233 = ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) ;
 assign wire393 = ( (~ f)  &  g  &  (~ h)  &  n_n711 ) | ( (~ f)  &  (~ g)  &  (~ h)  &  n_n711 ) ;
 assign n_n1177 = ( (~ m)  &  n ) ;
 assign n_n1165 = ( (~ m)  &  (~ n) ) ;
 assign n_n904 = ( a  &  (~ c)  &  d ) ;
 assign n_n626 = ( c  &  (~ e)  &  f ) ;
 assign n_n671 = ( (~ b)  &  c  &  f ) ;
 assign n_n1101 = ( (~ c)  &  d  &  f ) ;
 assign n_n1229 = ( c  &  d  &  e ) ;
 assign n_n1193 = ( f  &  g  &  (~ i) ) ;
 assign n_n1344 = ( wire5207 ) | ( wire5208 ) | ( wire5209 ) | ( wire5210 ) ;
 assign wire22 = ( k  &  (~ l)  &  m  &  (~ n) ) ;
 assign wire31 = ( (~ i)  &  l  &  m ) | ( j  &  (~ l)  &  m ) ;
 assign wire45 = ( (~ j)  &  wire22 ) | ( j  &  wire58 ) ;
 assign wire54 = ( (~ j)  &  l  &  m  &  (~ n) ) ;
 assign wire71 = ( (~ f)  &  h ) ;
 assign wire101 = ( wire65 ) | ( h  &  k  &  (~ l) ) ;
 assign wire138 = ( wire22  &  n_n1228 ) | ( wire113  &  n_n1228 ) | ( wire22  &  n_n766 ) ;
 assign wire195 = ( f  &  g  &  j  &  wire58 ) ;
 assign wire232 = ( (~ c) ) | ( (~ d) ) | ( e ) | ( (~ f) ) ;
 assign wire258 = ( (~ e)  &  g  &  n_n904 ) ;
 assign wire371 = ( (~ e)  &  g  &  i  &  n_n904 ) ;
 assign n_n1217 = ( i  &  j  &  k ) ;
 assign n_n1201 = ( f  &  g  &  h ) ;
 assign n_n1220 = ( k  &  m  &  (~ n) ) ;
 assign n_n920 = ( a  &  b  &  (~ c) ) ;
 assign n_n918 = ( a  &  b  &  d ) ;
 assign wire15 = ( a  &  (~ b)  &  c ) | ( (~ a)  &  b  &  (~ d) ) ;
 assign wire58 = ( (~ k)  &  l  &  m  &  (~ n) ) ;
 assign wire82 = ( wire41 ) | ( wire1012 ) | ( n_n1161  &  n_n904 ) ;
 assign wire98 = ( n_n1207  &  wire29 ) | ( n_n918  &  n_n1104 ) ;
 assign wire130 = ( wire228 ) | ( wire265 ) ;
 assign wire220 = ( m  &  (~ n)  &  wire25 ) | ( m  &  (~ n)  &  wire32 ) ;
 assign wire228 = ( j  &  l  &  m  &  (~ n) ) ;
 assign wire265 = ( j  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire390 = ( n_n1193  &  wire228 ) | ( n_n1193  &  wire265 ) ;
 assign wire417 = ( wire228  &  n_n861 ) | ( wire265  &  n_n861 ) ;
 assign n_n1187 = ( m  &  (~ n) ) ;
 assign n_n996 = ( (~ j)  &  k  &  l ) ;
 assign n_n1155 = ( g  &  h  &  (~ i) ) ;
 assign n_n1171 = ( b  &  e  &  (~ f) ) ;
 assign n_n698 = ( (~ a)  &  b  &  e ) ;
 assign n_n617 = ( h  &  j  &  (~ k) ) ;
 assign n_n730 = ( a  &  d  &  (~ e) ) ;
 assign n_n618 = ( h  &  (~ j)  &  k ) ;
 assign n_n857 = ( (~ f)  &  g  &  i ) ;
 assign n_n933 = ( (~ i)  &  j  &  l ) ;
 assign n_n821 = ( (~ g)  &  h  &  (~ i) ) ;
 assign n_n700 = ( (~ c)  &  d  &  (~ e) ) ;
 assign n_n824 = ( f  &  h  &  (~ i) ) ;
 assign n_n1792 = ( wire928 ) | ( wire929 ) | ( wire5406 ) | ( wire5407 ) ;
 assign wire29 = ( a  &  (~ b)  &  c ) | ( a  &  b  &  (~ c) ) | ( (~ a)  &  b  &  (~ d) ) ;
 assign wire30 = ( b  &  d  &  f ) | ( b  &  (~ e)  &  f ) ;
 assign wire34 = ( (~ c)  &  d  &  f ) | ( c  &  (~ d)  &  f ) | ( c  &  (~ e)  &  f ) ;
 assign wire179 = ( n_n996  &  n_n1228 ) | ( n_n1207  &  n_n747 ) ;
 assign wire210 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) | ( (~ b)  &  c  &  (~ e) ) ;
 assign wire255 = ( g  &  (~ h) ) ;
 assign wire291 = ( m  &  (~ n)  &  n_n1201  &  wire15 ) ;
 assign wire309 = ( (~ f)  &  h  &  n_n709 ) ;
 assign wire380 = ( g  &  h  &  (~ i)  &  wire54 ) ;
 assign n_n1069 = ( (~ c)  &  (~ d)  &  e ) ;
 assign n_n1104 = ( (~ f)  &  g  &  (~ h) ) ;
 assign n_n1203 = ( c  &  e  &  (~ f) ) ;
 assign n_n876 = ( a  &  c  &  (~ d) ) ;
 assign n_n1166 = ( (~ h)  &  i  &  (~ j) ) ;
 assign n_n1425 = ( wire871 ) | ( wire5474 ) | ( wire5475 ) ;
 assign wire74 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire76 = ( (~ j)  &  l  &  (~ m)  &  n ) ;
 assign wire92 = ( n_n1233  &  wire20 ) | ( n_n942  &  wire5499 ) ;
 assign wire112 = ( f  &  g ) ;
 assign wire120 = ( a  &  m  &  (~ n) ) ;
 assign wire183 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  l ) | ( j  &  (~ k)  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire184 = ( g  &  n_n842  &  wire71 ) | ( g  &  n_n711  &  wire71 ) | ( (~ g)  &  n_n711  &  wire71 ) ;
 assign wire196 = ( (~ b)  &  f ) ;
 assign wire223 = ( m  &  (~ n)  &  n_n920  &  n_n1233 ) ;
 assign wire230 = ( (~ f)  &  (~ h)  &  i ) | ( g  &  (~ h)  &  i ) ;
 assign wire256 = ( c  &  e ) ;
 assign n_n841 = ( g  &  (~ h)  &  i ) ;
 assign n_n893 = ( i  &  (~ j)  &  l ) ;
 assign n_n1194 = ( f  &  (~ g)  &  h ) ;
 assign n_n1495 = ( wire5583 ) | ( wire5584 ) | ( wire5585 ) ;
 assign wire33 = ( wire22 ) | ( wire113 ) ;
 assign wire93 = ( (~ b)  &  c  &  (~ e) ) | ( (~ b)  &  c  &  f ) | ( b  &  e  &  (~ f) ) ;
 assign wire106 = ( n_n920  &  n_n1194 ) | ( n_n918  &  n_n971 ) ;
 assign wire156 = ( n_n1207  &  n_n920 ) | ( n_n918  &  n_n1104 ) ;
 assign wire203 = ( n_n918  &  n_n857 ) | ( n_n920  &  n_n1228 ) ;
 assign wire219 = ( m  &  (~ n)  &  n_n918  &  n_n1195 ) ;
 assign n_n1138 = ( (~ c)  &  (~ d)  &  (~ f) ) ;
 assign n_n1159 = ( (~ j)  &  (~ k)  &  (~ l) ) ;
 assign n_n2507 = ( wire283  &  n_n1253  &  n_n978  &  n_n1249 ) ;
 assign n_n1080 = ( (~ c)  &  (~ d)  &  (~ e) ) ;
 assign n_n2494 = ( n_n1104  &  n_n973  &  (~ wire118)  &  wire188 ) ;
 assign wire116 = ( wire780 ) | ( n_n1142  &  n_n989  &  wire5639 ) ;
 assign wire199 = ( n_n2602 ) | ( wire777 ) ;
 assign wire319 = ( wire775 ) | ( wire776 ) ;
 assign n_n1190 = ( (~ l)  &  (~ m)  &  (~ n) ) ;
 assign n_n1202 = ( (~ k)  &  (~ m)  &  (~ n) ) ;
 assign n_n1039 = ( (~ f)  &  (~ g)  &  (~ h) ) ;
 assign n_n2602 = ( n_n1207  &  n_n1069  &  (~ wire118)  &  wire188 ) ;
 assign n_n2511 = ( n_n987  &  n_n988  &  wire283  &  n_n978 ) ;
 assign n_n2493 = ( n_n1104  &  n_n975  &  (~ wire118)  &  wire188 ) ;
 assign wire157 = ( wire765 ) | ( n_n1260  &  n_n992  &  wire5659 ) ;
 assign wire267 = ( wire762 ) | ( n_n1215  &  wire5629  &  wire5633 ) ;
 assign n_n1142 = ( (~ g)  &  h  &  i ) ;
 assign n_n949 = ( a  &  (~ b)  &  c ) ;
 assign n_n761 = ( a  &  c  &  e ) ;
 assign n_n1231 = ( (~ e)  &  f  &  g ) ;
 assign n_n1261 = ( a  &  b  &  c ) ;
 assign n_n997 = ( (~ a)  &  b  &  c ) ;
 assign n_n1874 = ( wire751 ) | ( wire5685 ) | ( wire5686 ) | ( wire5687 ) ;
 assign wire44 = ( h  &  wire22 ) | ( (~ g)  &  wire190 ) ;
 assign wire57 = ( (~ c) ) | ( (~ d) ) ;
 assign wire94 = ( n_n1220  &  n_n1194 ) | ( n_n1219  &  n_n822 ) ;
 assign wire108 = ( wire22  &  n_n1083 ) | ( n_n912  &  wire190 ) ;
 assign wire200 = ( n_n1220  &  n_n971 ) | ( n_n1219  &  n_n825 ) ;
 assign wire254 = ( (~ k)  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire379 = ( g  &  (~ j)  &  wire22 ) | ( g  &  j  &  wire58 ) ;
 assign wire387 = ( k  &  m  &  (~ n)  &  n_n1082 ) ;
 assign wire407 = ( (~ g)  &  (~ h)  &  (~ i) ) ;
 assign wire413 = ( a  &  c  &  (~ d)  &  n_n864 ) ;
 assign n_n872 = ( a  &  (~ d)  &  e ) ;
 assign n_n838 = ( b  &  d  &  f ) ;
 assign n_n977 = ( (~ i)  &  j  &  (~ k) ) ;
 assign n_n1252 = ( e  &  f  &  g ) ;
 assign n_n1920 = ( wire5731 ) | ( wire5732 ) | ( wire38  &  wire92 ) ;
 assign n_n1919 = ( wire700 ) | ( wire703 ) | ( wire5740 ) | ( wire5743 ) ;
 assign n_n987 = ( e  &  (~ f)  &  g ) ;
 assign n_n1210 = ( k  &  (~ m)  &  n ) ;
 assign n_n1939 = ( n_n2511 ) | ( n_n2493 ) | ( wire5774 ) | ( wire5775 ) ;
 assign n_n988 = ( (~ b)  &  c  &  d ) ;
 assign wire39 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  l ) | ( i  &  k  &  (~ l) ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire77 = ( k  &  (~ l)  &  (~ m)  &  n ) ;
 assign wire89 = ( f  &  (~ h)  &  i ) | ( f  &  h  &  (~ i) ) | ( f  &  h  &  (~ j) ) ;
 assign wire111 = ( m  &  (~ n)  &  n_n949 ) ;
 assign wire117 = ( n_n1036  &  n_n823 ) | ( n_n1056  &  n_n822 ) ;
 assign wire135 = ( n_n1036  &  n_n1137 ) | ( n_n1056  &  n_n817 ) ;
 assign wire159 = ( n_n872  &  n_n861 ) | ( n_n876  &  n_n864 ) ;
 assign wire160 = ( n_n1082  &  n_n1253 ) | ( n_n1195  &  wire5751 ) ;
 assign wire164 = ( g  &  (~ h)  &  i ) | ( g  &  h  &  (~ i) ) | ( g  &  h  &  (~ j) ) ;
 assign wire165 = ( i  &  (~ j)  &  k ) | ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) | ( i  &  k  &  (~ l) ) ;
 assign wire167 = ( n_n1253  &  wire5752 ) | ( n_n1104  &  wire5753 ) ;
 assign wire386 = ( (~ i)  &  (~ k) ) ;
 assign n_n1022 = ( f  &  h  &  (~ j) ) ;
 assign n_n1573 = ( wire5848 ) | ( wire5849 ) | ( wire5850 ) | ( wire5851 ) ;
 assign n_n820 = ( g  &  h  &  (~ j) ) ;
 assign n_n1264 = ( h  &  i  &  j ) ;
 assign n_n3060 = ( i  &  n_n904  &  wire113  &  wire128 ) ;
 assign wire14 = ( a  &  c  &  e ) | ( a  &  (~ d)  &  e ) ;
 assign wire40 = ( h  &  (~ i)  &  k ) | ( h  &  (~ j)  &  k ) ;
 assign wire113 = ( (~ j)  &  k  &  m  &  (~ n) ) ;
 assign wire208 = ( g  &  n_n1171  &  wire146 ) | ( (~ g)  &  wire30  &  wire146 ) ;
 assign wire351 = ( wire113  &  wire80 ) | ( n_n876  &  wire113  &  n_n859 ) ;
 assign n_n1085 = ( h  &  i  &  (~ j) ) ;
 assign n_n1036 = ( (~ k)  &  (~ m)  &  n ) ;
 assign n_n1053 = ( (~ b)  &  c  &  (~ e) ) ;
 assign n_n619 = ( (~ h)  &  i  &  k ) ;
 assign n_n1653 = ( wire5903 ) | ( wire5904 ) | ( wire5905 ) | ( wire5906 ) ;
 assign n_n816 = ( (~ g)  &  h  &  k ) ;
 assign wire21 = ( (~ j)  &  k  &  (~ m) ) | ( j  &  (~ k)  &  (~ m) ) ;
 assign wire36 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) ;
 assign wire50 = ( wire14  &  n_n971 ) | ( n_n876  &  n_n1082 ) ;
 assign wire207 = ( wire29  &  n_n1194 ) | ( n_n918  &  n_n971 ) ;
 assign wire209 = ( n_n1203  &  n_n1202 ) | ( n_n1202  &  n_n623 ) | ( n_n1036  &  n_n623 ) ;
 assign wire290 = ( g  &  h  &  i  &  (~ n) ) ;
 assign wire315 = ( m  &  (~ n)  &  n_n698 ) ;
 assign wire320 = ( wire5814 ) | ( wire70  &  wire641 ) | ( wire70  &  wire642 ) ;
 assign n_n1219 = ( (~ l)  &  m  &  (~ n) ) ;
 assign n_n2023 = ( wire6168 ) | ( wire6169 ) | ( wire6170 ) | ( wire6171 ) ;
 assign wire114 = ( (~ g)  &  (~ h) ) ;
 assign wire127 = ( (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire146 = ( h  &  (~ j) ) ;
 assign wire222 = ( g  &  h ) ;
 assign wire263 = ( (~ b)  &  (~ m)  &  n ) ;
 assign wire268 = ( (~ c)  &  e  &  (~ f) ) | ( c  &  (~ e)  &  (~ f) ) ;
 assign wire404 = ( (~ b)  &  m  &  (~ n) ) ;
 assign n_n971 = ( (~ f)  &  (~ g)  &  h ) ;
 assign n_n1204 = ( l  &  (~ m)  &  (~ n) ) ;
 assign n_n973 = ( c  &  d  &  (~ e) ) ;
 assign n_n1072 = ( (~ d)  &  (~ e)  &  (~ f) ) ;
 assign n_n1028 = ( (~ e)  &  (~ f)  &  (~ g) ) ;
 assign wire37 = ( h ) | ( i ) ;
 assign wire68 = ( i ) | ( j ) ;
 assign wire384 = ( h  &  (~ i)  &  (~ j) ) ;
 assign n_n1160 = ( (~ e)  &  f  &  (~ h) ) ;
 assign n_n662 = ( (~ f)  &  (~ h)  &  i ) ;
 assign wire282 = ( j  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire373 = ( (~ h)  &  (~ i)  &  (~ j)  &  l ) ;
 assign n_n1180 = ( i  &  (~ j)  &  (~ k) ) ;
 assign n_n1196 = ( (~ e)  &  g  &  h ) ;
 assign wire103 = ( (~ e)  &  (~ f) ) ;
 assign wire204 = ( f ) | ( (~ m) ) | ( n ) ;
 assign wire227 = ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire273 = ( b ) | ( j ) ;
 assign n_n1121 = ( (~ b)  &  e  &  (~ f) ) ;
 assign n_n1164 = ( c  &  (~ e)  &  (~ f) ) ;
 assign n_n1222 = ( (~ k)  &  m  &  (~ n) ) ;
 assign n_n1095 = ( f  &  (~ h)  &  i ) ;
 assign n_n975 = ( (~ c)  &  d  &  e ) ;
 assign wire70 = ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire221 = ( (~ j)  &  k  &  (~ m)  &  n ) ;
 assign wire234 = ( h ) | ( i ) | ( j ) ;
 assign wire283 = ( (~ h)  &  (~ i)  &  j ) ;
 assign wire285 = ( (~ i)  &  (~ k)  &  (~ m)  &  n ) ;
 assign wire286 = ( (~ h)  &  (~ i)  &  (~ m)  &  n ) ;
 assign wire301 = ( (~ k)  &  (~ l)  &  (~ m)  &  n ) ;
 assign n_n1148 = ( e  &  g  &  h ) ;
 assign n_n1137 = ( g  &  h  &  j ) ;
 assign n_n1191 = ( k  &  (~ m)  &  (~ n) ) ;
 assign n_n1195 = ( (~ f)  &  g  &  h ) ;
 assign n_n1133 = ( i  &  (~ j)  &  k ) ;
 assign n_n861 = ( (~ f)  &  g  &  (~ i) ) ;
 assign n_n1082 = ( e  &  (~ g)  &  h ) ;
 assign n_n1260 = ( d  &  e  &  f ) ;
 assign n_n819 = ( (~ g)  &  h  &  (~ j) ) ;
 assign n_n1131 = ( g  &  i  &  k ) ;
 assign wire79 = ( (~ c)  &  d  &  (~ e) ) | ( c  &  e  &  (~ f) ) ;
 assign wire122 = ( (~ h) ) | ( (~ i) ) ;
 assign wire158 = ( (~ c)  &  g  &  h ) | ( (~ f)  &  g  &  h ) ;
 assign wire170 = ( (~ j)  &  (~ m)  &  (~ n) ) ;
 assign wire194 = ( (~ g)  &  h ) ;
 assign n_n1243 = ( (~ i)  &  (~ k)  &  (~ m) ) ;
 assign n_n1227 = ( j  &  (~ k)  &  (~ m) ) ;
 assign n_n1091 = ( (~ c)  &  (~ f)  &  (~ g) ) ;
 assign wire95 = ( c  &  (~ f) ) | ( (~ c)  &  g ) ;
 assign wire132 = ( (~ h)  &  i ) ;
 assign wire226 = ( (~ h)  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire395 = ( (~ c)  &  (~ d) ) | ( (~ c)  &  (~ f) ) ;
 assign n_n818 = ( (~ g)  &  h  &  j ) ;
 assign n_n529 = ( g  &  (~ i)  &  j ) ;
 assign n_n670 = ( h  &  (~ i)  &  j ) ;
 assign wire23 = ( g  &  (~ h)  &  i ) | ( g  &  h  &  (~ i) ) ;
 assign wire59 = ( f  &  (~ h)  &  i ) | ( f  &  h  &  (~ i) ) ;
 assign wire96 = ( (~ k)  &  m  &  (~ n) ) | ( l  &  m  &  (~ n) ) ;
 assign wire134 = ( (~ g)  &  (~ h)  &  i ) | ( (~ g)  &  h  &  (~ i) ) ;
 assign wire169 = ( b  &  e  &  (~ f)  &  n_n841 ) ;
 assign wire398 = ( (~ h)  &  i  &  j ) ;
 assign n_n387 = ( g  &  (~ j)  &  k ) ;
 assign wire72 = ( n_n1219  &  n_n387 ) | ( n_n1220  &  n_n694 ) ;
 assign wire211 = ( (~ g)  &  n_n711  &  wire146 ) | ( g  &  wire146  &  wire47 ) ;
 assign wire231 = ( (~ f)  &  h  &  (~ i) ) | ( (~ f)  &  h  &  (~ j) ) ;
 assign wire137 = ( (~ g) ) | ( (~ j) ) ;
 assign n_n1118 = ( (~ k)  &  (~ l)  &  (~ m) ) ;
 assign n_n1216 = ( l  &  (~ m)  &  n ) ;
 assign n_n1056 = ( (~ l)  &  (~ m)  &  n ) ;
 assign wire189 = ( (~ e)  &  f ) ;
 assign n_n868 = ( j  &  (~ l)  &  m ) ;
 assign n_n823 = ( f  &  h  &  j ) ;
 assign wire259 = ( d  &  (~ e) ) ;
 assign n_n989 = ( j  &  (~ k)  &  l ) ;
 assign n_n1094 = ( (~ g)  &  (~ h)  &  i ) ;
 assign wire249 = ( c  &  (~ d) ) ;
 assign n_n628 = ( c  &  (~ d)  &  f ) ;
 assign n_n623 = ( c  &  f  &  (~ g) ) ;
 assign wire128 = ( (~ e)  &  g ) ;
 assign wire396 = ( b  &  (~ c) ) ;
 assign n_n992 = ( g  &  h  &  i ) ;
 assign wire118 = ( i ) | ( (~ j) ) ;
 assign n_n1146 = ( j  &  k  &  l ) ;
 assign wire121 = ( h  &  k ) ;
 assign n_n1228 = ( f  &  g  &  i ) ;
 assign n_n1116 = ( i  &  k  &  (~ m) ) ;
 assign n_n1215 = ( l  &  m  &  (~ n) ) ;
 assign n_n1233 = ( (~ d)  &  f  &  g ) ;
 assign n_n940 = ( e  &  f  &  (~ g) ) ;
 assign n_n942 = ( h  &  (~ j)  &  l ) ;
 assign n_n765 = ( f  &  g  &  j ) ;
 assign n_n822 = ( f  &  h  &  k ) ;
 assign n_n859 = ( e  &  g  &  i ) ;
 assign n_n1253 = ( b  &  c  &  d ) ;
 assign wire248 = ( (~ m)  &  n  &  n_n1252  &  n_n1253 ) ;
 assign wire314 = ( h  &  (~ i) ) ;
 assign wire55 = ( j  &  (~ k)  &  l ) | ( (~ j)  &  k  &  (~ l) ) ;
 assign wire149 = ( (~ i)  &  j  &  (~ k) ) | ( (~ i)  &  j  &  l ) ;
 assign wire18 = ( i  &  (~ j)  &  k ) | ( i  &  k  &  (~ l) ) ;
 assign wire20 = ( (~ h)  &  i  &  l ) | ( h  &  (~ i)  &  l ) | ( h  &  j  &  (~ l) ) ;
 assign n_n874 = ( i  &  l  &  m ) ;
 assign n_n605 = ( j  &  (~ k)  &  (~ l) ) ;
 assign n_n1084 = ( (~ f)  &  h  &  (~ j) ) ;
 assign n_n766 = ( f  &  g  &  (~ j) ) ;
 assign n_n875 = ( e  &  g  &  (~ h) ) ;
 assign n_n871 = ( (~ i)  &  l  &  m ) ;
 assign wire90 = ( d  &  e ) ;
 assign n_n235 = ( h  &  k  &  (~ l) ) ;
 assign n_n2572 = ( n_n876  &  wire113  &  n_n859 ) ;
 assign n_n2953 = ( n_n698  &  n_n1137  &  wire5830 ) ;
 assign n_n1167 = ( (~ c)  &  e  &  (~ f) ) ;
 assign n_n1083 = ( (~ e)  &  f  &  h ) ;
 assign n_n1189 = ( (~ a)  &  d  &  (~ e) ) ;
 assign n_n978 = ( k  &  l  &  (~ m)  &  n ) ;
 assign n_n703 = ( b  &  (~ e)  &  f ) ;
 assign n_n864 = ( e  &  g  &  (~ i) ) ;
 assign n_n817 = ( g  &  h  &  k ) ;
 assign wire197 = ( g  &  (~ j) ) ;
 assign wire161 = ( (~ k)  &  m  &  (~ n) ) | ( (~ l)  &  m  &  (~ n) ) ;
 assign wire305 = ( (~ c)  &  (~ d)  &  i ) ;
 assign wire399 = ( (~ g)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire414 = ( a  &  c  &  (~ d)  &  n_n859 ) ;
 assign wire369 = ( a  &  c  &  (~ d)  &  e ) ;
 assign n_n2660 = ( g  &  j  &  wire58  &  wire369 ) ;
 assign n_n982 = ( (~ k)  &  l  &  (~ m)  &  n ) ;
 assign wire47 = ( b  &  (~ c)  &  d ) | ( b  &  c  &  (~ d) ) | ( b  &  (~ d)  &  e ) ;
 assign n_n1249 = ( (~ e)  &  (~ f)  &  g ) ;
 assign n_n919 = ( d  &  (~ e)  &  g ) ;
 assign n_n694 = ( g  &  i  &  (~ j) ) ;
 assign n_n844 = ( k  &  (~ l)  &  (~ m) ) ;
 assign n_n912 = ( (~ e)  &  f  &  (~ g) ) ;
 assign wire35 = ( c  &  e  &  (~ f) ) | ( c  &  f  &  (~ g) ) ;
 assign n_n2026 = ( wire6251 ) | ( wire6252 ) | ( wire6256 ) ;
 assign wire56 = ( (~ h)  &  i  &  k ) | ( h  &  j  &  (~ k) ) ;
 assign wire142 = ( k  &  l  &  m  &  (~ n) ) ;
 assign wire188 = ( k  &  l  &  (~ m)  &  (~ n) ) ;
 assign wire216 = ( (~ g)  &  h  &  (~ j) ) | ( (~ g)  &  h  &  k ) | ( g  &  j  &  (~ k) ) ;
 assign wire260 = ( (~ j)  &  l  &  (~ m)  &  (~ n) ) ;
 assign n_n747 = ( i  &  j  &  l ) ;
 assign wire181 = ( wire20 ) | ( (~ i)  &  j  &  (~ k) ) ;
 assign wire104 = ( (~ e)  &  g  &  h ) | ( f  &  g  &  h ) ;
 assign wire293 = ( (~ j)  &  k  &  (~ m)  &  n ) | ( j  &  (~ k)  &  (~ m)  &  n ) ;
 assign n_n825 = ( (~ f)  &  h  &  k ) ;
 assign wire43 = ( (~ a)  &  b  &  (~ d) ) | ( (~ a)  &  b  &  e ) ;
 assign wire24 = ( (~ c)  &  d  &  f ) | ( c  &  (~ e)  &  f ) ;
 assign wire49 = ( (~ i)  &  k  &  (~ m) ) | ( (~ j)  &  k  &  (~ m) ) | ( j  &  (~ k)  &  (~ m) ) ;
 assign wire109 = ( (~ c)  &  d  &  (~ e) ) | ( (~ c)  &  d  &  f ) | ( c  &  (~ e)  &  f ) | ( c  &  e  &  (~ f) ) ;
 assign wire206 = ( (~ g)  &  h  &  i ) | ( g  &  i  &  (~ j) ) ;
 assign wire105 = ( (~ g)  &  h  &  (~ j) ) | ( g  &  j  &  (~ k) ) ;
 assign wire152 = ( (~ l)  &  n_n1187  &  n_n1137 ) | ( l  &  n_n1187  &  wire23 ) ;
 assign wire299 = ( (~ e)  &  g  &  (~ h)  &  n_n904 ) ;
 assign wire388 = ( n_n918  &  n_n1187  &  n_n1231 ) | ( n_n918  &  n_n1187  &  n_n1249 ) ;
 assign wire65 = ( (~ h)  &  i  &  k ) | ( h  &  (~ i)  &  k ) | ( h  &  (~ j)  &  k ) | ( h  &  j  &  (~ k) ) ;
 assign wire162 = ( wire282 ) | ( (~ n_n1264)  &  n_n1191 ) ;
 assign wire198 = ( h  &  j  &  (~ k) ) | ( h  &  k  &  (~ l) ) ;
 assign wire377 = ( (~ f)  &  g  &  h  &  n_n711 ) | ( (~ f)  &  (~ g)  &  h  &  n_n711 ) ;
 assign wire385 = ( (~ f)  &  g  &  h  &  (~ n) ) ;
 assign wire16 = ( a  &  (~ c)  &  d ) | ( a  &  d  &  (~ e) ) ;
 assign wire25 = ( n_n876  &  n_n1148 ) | ( wire14  &  n_n1195 ) ;
 assign wire32 = ( n_n904  &  n_n1201 ) | ( n_n1201  &  n_n730 ) | ( n_n904  &  n_n1196 ) ;
 assign wire41 = ( n_n1104  &  wire14 ) | ( n_n876  &  n_n875 ) ;
 assign wire60 = ( (~ b)  &  c  &  (~ e) ) | ( b  &  e  &  (~ f) ) ;
 assign wire69 = ( wire54  &  n_n1082 ) | ( wire148  &  n_n875 ) ;
 assign wire80 = ( n_n857  &  wire14 ) | ( n_n1228  &  wire16 ) ;
 assign wire81 = ( wire265  &  n_n1155 ) | ( wire58  &  n_n1137 ) ;
 assign wire85 = ( (~ j)  &  m  &  (~ n) ) | ( k  &  m  &  (~ n) ) ;
 assign wire190 = ( h  &  k  &  m  &  (~ n) ) ;
 assign wire115 = ( n_n713  &  n_n886 ) | ( n_n1253  &  n_n1083 ) ;
 assign wire368 = ( e  &  g  &  h  &  (~ n) ) ;
 assign wire42 = ( n_n971  &  n_n1204  &  n_n973  &  wire6310 ) ;
 assign wire61 = ( n_n1165  &  n_n1138  &  n_n1142  &  n_n1146 ) ;
 assign wire63 = ( n_n1138  &  wire254  &  wire407 ) ;
 assign wire66 = ( n_n988  &  n_n1028  &  wire384  &  n_n982 ) ;
 assign wire140 = ( n_n1202  &  (~ wire268)  &  wire6287 ) ;
 assign wire150 = ( m  &  (~ n)  &  n_n1180  &  wire6289 ) ;
 assign wire163 = ( (~ c)  &  (~ d)  &  n_n1155  &  wire127 ) ;
 assign wire173 = ( (~ a)  &  (~ b)  &  m  &  (~ n) ) ;
 assign wire177 = ( (~ b)  &  (~ c)  &  (~ m)  &  n ) ;
 assign wire178 = ( (~ g)  &  (~ h)  &  m  &  (~ n) ) ;
 assign wire180 = ( (~ j)  &  (~ k)  &  (~ l)  &  n_n1219 ) ;
 assign wire252 = ( (~ n_n861)  &  wire395  &  wire6257  &  wire6258 ) ;
 assign wire253 = ( wire6262  &  wire6263 ) ;
 assign wire269 = ( wire395  &  (~ n_n1118)  &  wire6264 ) ;
 assign wire271 = ( wire127  &  (~ n_n765)  &  wire6266 ) ;
 assign wire272 = ( wire254  &  wire6268 ) ;
 assign wire274 = ( h  &  (~ j)  &  (~ wire127)  &  n_n1118 ) ;
 assign wire275 = ( h  &  (~ j)  &  n_n1036  &  n_n1082 ) ;
 assign wire276 = ( g  &  n_n1080  &  wire127 ) | ( h  &  n_n1080  &  wire127 ) ;
 assign wire277 = ( (~ c)  &  e  &  (~ f)  &  wire6272 ) ;
 assign wire278 = ( n_n1194  &  n_n1202  &  n_n819 ) ;
 assign wire280 = ( n_n1202  &  n_n1083  &  n_n694 ) ;
 assign wire281 = ( (~ m)  &  (~ n)  &  wire114  &  n_n1164 ) ;
 assign wire307 = ( (~ n_n912)  &  wire6211  &  wire6216  &  wire6217 ) ;
 assign wire316 = ( (~ wire35)  &  wire6225  &  wire6226  &  wire6227 ) ;
 assign wire317 = ( n_n1190  &  (~ wire127)  &  (~ n_n919)  &  wire6230 ) ;
 assign wire318 = ( (~ e)  &  (~ f)  &  wire234  &  wire6233 ) ;
 assign wire321 = ( (~ i)  &  n_n1165  &  n_n1072  &  n_n1164 ) ;
 assign wire322 = ( (~ m)  &  (~ n)  &  n_n1164  &  wire6236 ) ;
 assign wire328 = ( (~ m)  &  n  &  n_n1069  &  n_n940 ) ;
 assign wire329 = ( (~ g)  &  n_n1072  &  wire85 ) ;
 assign wire330 = ( m  &  (~ n)  &  n_n700  &  n_n1189 ) ;
 assign wire331 = ( (~ l)  &  m  &  (~ n)  &  n_n1189 ) ;
 assign wire333 = ( (~ n_n1171)  &  (~ n_n700)  &  (~ n_n973)  &  wire6177 ) ;
 assign wire334 = ( (~ wire263)  &  wire286  &  n_n1216  &  wire6180 ) ;
 assign wire336 = ( (~ n_n1216)  &  (~ n_n1249)  &  wire6185 ) ;
 assign wire337 = ( wire6187  &  wire6188 ) ;
 assign wire338 = ( (~ wire407)  &  wire170  &  wire226 ) ;
 assign wire339 = ( a  &  j  &  wire399 ) | ( (~ b)  &  j  &  wire399 ) ;
 assign wire340 = ( n_n1210  &  wire286  &  (~ n_n1216) ) ;
 assign wire341 = ( (~ e)  &  wire286  &  (~ n_n1216) ) ;
 assign wire342 = ( n_n1171  &  wire286  &  n_n1056 ) ;
 assign wire345 = ( i  &  (~ m)  &  n  &  n_n1028 ) ;
 assign wire347 = ( (~ d)  &  (~ m)  &  n  &  n_n1121 ) ;
 assign wire352 = ( (~ c)  &  (~ d)  &  f  &  wire6151 ) | ( (~ c)  &  d  &  (~ f)  &  wire6151 ) ;
 assign wire353 = ( j  &  wire232  &  wire399 ) ;
 assign wire354 = ( (~ c)  &  wire286 ) | ( (~ d)  &  wire286 ) ;
 assign wire355 = ( i  &  n_n1072  &  (~ wire204) ) | ( j  &  n_n1072  &  (~ wire204) ) ;
 assign wire357 = ( (~ c)  &  (~ d)  &  n_n1190  &  (~ n_n1091) ) ;
 assign wire359 = ( (~ m)  &  n  &  n_n1028  &  wire68 ) ;
 assign wire362 = ( (~ l)  &  (~ m)  &  n  &  n_n1028 ) ;
 assign wire389 = ( (~ l)  &  (~ m)  &  (~ n)  &  n_n1164 ) ;
 assign wire424 = ( i  &  m  &  (~ n)  &  n_n1039 ) ;
 assign wire425 = ( c  &  (~ g)  &  wire226 ) ;
 assign wire429 = ( n_n1217  &  (~ n_n1260)  &  n_n1215  &  wire6109 ) ;
 assign wire430 = ( n_n1217  &  n_n1215  &  wire6112 ) ;
 assign wire431 = ( n_n1217  &  wire196  &  n_n1264  &  n_n1216 ) ;
 assign wire432 = ( n_n1177  &  wire103  &  n_n1253  &  wire6115 ) ;
 assign wire433 = ( (~ m)  &  n  &  n_n1253  &  wire6118 ) ;
 assign wire434 = ( n_n1227  &  n_n1228  &  wire6119 ) ;
 assign wire435 = ( n_n1177  &  n_n1253  &  wire314  &  n_n1249 ) ;
 assign wire440 = ( n_n1187  &  n_n1261  &  (~ wire222)  &  n_n1260 ) ;
 assign wire441 = ( wire285  &  n_n1253  &  n_n1249 ) ;
 assign wire442 = ( n_n1177  &  n_n1252  &  wire132  &  n_n1253 ) ;
 assign wire443 = ( n_n1022  &  n_n1204  &  wire6072 ) ;
 assign wire444 = ( n_n1187  &  n_n1261  &  (~ n_n1253)  &  wire6074 ) ;
 assign wire445 = ( (~ k)  &  n_n1187  &  n_n1261  &  wire6076 ) ;
 assign wire446 = ( n_n1217  &  n_n1204  &  (~ n_n1091)  &  wire6078 ) ;
 assign wire447 = ( i  &  n_n1207  &  n_n1165  &  n_n1229 ) ;
 assign wire448 = ( n_n1210  &  n_n1253  &  wire6082 ) ;
 assign wire449 = ( n_n1203  &  n_n1202  &  wire384 ) ;
 assign wire450 = ( wire373  &  wire6085 ) ;
 assign wire451 = ( (~ n_n1188)  &  n_n1229  &  n_n1193  &  n_n1190 ) ;
 assign wire452 = ( n_n1217  &  (~ n_n1138)  &  n_n1204  &  wire194 ) ;
 assign wire453 = ( n_n1187  &  n_n1261  &  wire189  &  (~ n_n1253) ) ;
 assign wire454 = ( n_n1229  &  wire170  &  n_n1228 ) ;
 assign wire455 = ( n_n1229  &  n_n1193  &  n_n1204 ) ;
 assign wire456 = ( n_n1229  &  n_n1201  &  n_n1190 ) ;
 assign wire457 = ( n_n1217  &  wire158  &  n_n1215 ) ;
 assign wire458 = ( m  &  (~ n)  &  n_n1188  &  n_n1189 ) ;
 assign wire459 = ( (~ j)  &  n_n1177  &  n_n1252  &  n_n1253 ) ;
 assign wire460 = ( n_n1217  &  n_n1204  &  wire158 ) ;
 assign wire461 = ( (~ n_n1203)  &  n_n1204  &  (~ n_n1227)  &  wire6042 ) ;
 assign wire463 = ( (~ n_n857)  &  wire395  &  wire6047 ) ;
 assign wire464 = ( (~ n)  &  wire114  &  n_n1227  &  (~ n_n1091) ) ;
 assign wire465 = ( n_n1161  &  wire226  &  wire395 ) ;
 assign wire466 = ( (~ g)  &  n_n1204  &  (~ wire95)  &  wire226 ) ;
 assign wire467 = ( g  &  (~ h)  &  n_n1204  &  n_n1243 ) ;
 assign wire468 = ( wire254  &  wire6054 ) ;
 assign wire469 = ( n_n1190  &  wire95  &  wire226 ) ;
 assign wire470 = ( (~ e)  &  (~ h)  &  i  &  wire70 ) ;
 assign wire471 = ( (~ c)  &  d  &  (~ g)  &  wire226 ) ;
 assign wire480 = ( n_n1133  &  wire170  &  wire6005 ) ;
 assign wire481 = ( n_n1159  &  wire170  &  wire6006 ) ;
 assign wire482 = ( (~ n_n1080)  &  n_n861  &  (~ wire79)  &  wire170 ) ;
 assign wire483 = ( n_n1072  &  wire170  &  wire6010 ) ;
 assign wire484 = ( n_n1082  &  wire170  &  wire6012 ) ;
 assign wire485 = ( n_n1131  &  (~ wire79)  &  wire6014 ) ;
 assign wire486 = ( (~ n_n1080)  &  n_n1202  &  n_n861  &  (~ wire79) ) ;
 assign wire487 = ( n_n1165  &  n_n1137  &  n_n1195  &  (~ wire79) ) ;
 assign wire488 = ( n_n1164  &  n_n1191  &  wire6020 ) ;
 assign wire489 = ( m  &  (~ n)  &  n_n1189  &  wire6022 ) ;
 assign wire490 = ( (~ c)  &  d  &  n_n1202  &  n_n819 ) ;
 assign wire491 = ( n_n1159  &  wire158  &  wire170 ) ;
 assign wire492 = ( n_n1177  &  (~ n_n1260)  &  (~ wire122)  &  n_n1146 ) ;
 assign wire493 = ( n_n1177  &  n_n975  &  (~ wire122)  &  n_n1146 ) ;
 assign wire494 = ( m  &  (~ n)  &  n_n1180  &  n_n1195 ) ;
 assign wire495 = ( m  &  (~ n)  &  n_n1180  &  n_n1148 ) ;
 assign wire496 = ( (~ m)  &  n  &  n_n1142  &  n_n1146 ) ;
 assign wire499 = ( n_n1177  &  n_n1121  &  (~ wire70)  &  wire5971 ) ;
 assign wire500 = ( n_n1036  &  wire146  &  (~ wire263)  &  (~ n_n1196) ) ;
 assign wire501 = ( wire54  &  (~ n_n1203)  &  (~ n_n1164)  &  (~ wire234) ) ;
 assign wire502 = ( (~ g)  &  wire85  &  wire5977 ) ;
 assign wire503 = ( (~ b)  &  f  &  (~ h)  &  wire301 ) ;
 assign wire504 = ( (~ m)  &  n  &  n_n1121  &  wire5979 ) ;
 assign wire505 = ( n_n1161  &  wire263  &  wire286 ) ;
 assign wire508 = ( (~ b)  &  wire54  &  (~ wire234) ) ;
 assign wire509 = ( (~ wire204)  &  n_n1121  &  n_n975 ) ;
 assign wire510 = ( (~ b)  &  f  &  (~ h)  &  wire70 ) ;
 assign wire511 = ( (~ g)  &  n_n1187  &  n_n1189  &  wire85 ) ;
 assign wire512 = ( (~ m)  &  n  &  n_n1121  &  wire285 ) ;
 assign wire513 = ( (~ m)  &  n  &  n_n1121  &  wire221 ) ;
 assign wire516 = ( m  &  (~ n)  &  n_n1095  &  n_n1189 ) ;
 assign wire517 = ( (~ h)  &  (~ i)  &  (~ j)  &  wire58 ) ;
 assign wire520 = ( (~ e)  &  h  &  wire263  &  n_n1180 ) ;
 assign wire521 = ( wire373  &  wire5958 ) ;
 assign wire522 = ( m  &  (~ n)  &  n_n1180  &  wire5959 ) ;
 assign wire523 = ( (~ b)  &  (~ j)  &  n_n1036  &  n_n1196 ) ;
 assign wire527 = ( (~ m)  &  n  &  n_n1253  &  wire5964 ) ;
 assign wire528 = ( (~ c)  &  d  &  n_n1190  &  wire5941 ) ;
 assign wire532 = ( wire282  &  wire5946 ) ;
 assign wire533 = ( (~ m)  &  (~ n)  &  n_n1166  &  wire268 ) ;
 assign wire534 = ( i  &  j  &  n_n1161  &  n_n1202 ) ;
 assign wire535 = ( (~ m)  &  (~ n)  &  n_n1159  &  n_n1160 ) ;
 assign wire536 = ( n_n1220  &  n_n730  &  (~ n_n1053)  &  n_n816 ) ;
 assign wire537 = ( n_n700  &  wire21  &  wire290 ) ;
 assign wire539 = ( n_n841  &  n_n1210  &  wire36 ) ;
 assign wire540 = ( wire34  &  n_n1202  &  n_n1264 ) ;
 assign wire541 = ( n_n671  &  n_n1264  &  n_n1036 ) ;
 assign wire542 = ( n_n671  &  n_n1210  &  n_n619 ) ;
 assign wire543 = ( n_n671  &  n_n1210  &  n_n1085 ) ;
 assign wire544 = ( n_n841  &  n_n1210  &  n_n1053 ) ;
 assign wire545 = ( n_n904  &  n_n1220  &  n_n1194 ) ;
 assign wire546 = ( n_n711  &  n_n1142  &  wire70 ) | ( wire30  &  n_n1142  &  wire70 ) ;
 assign wire547 = ( wire34  &  n_n619  &  n_n1191 ) | ( n_n619  &  n_n1191  &  wire35 ) ;
 assign wire548 = ( wire34  &  n_n1085  &  n_n1191 ) | ( n_n1085  &  n_n1191  &  wire35 ) ;
 assign wire549 = ( m  &  (~ n)  &  n_n698  &  n_n816 ) ;
 assign wire550 = ( m  &  (~ n)  &  n_n698  &  n_n618 ) ;
 assign wire551 = ( n_n700  &  n_n841  &  n_n1191 ) ;
 assign wire552 = ( wire36  &  wire70  &  n_n992 ) ;
 assign wire554 = ( n_n709  &  wire230  &  n_n1210 ) ;
 assign wire565 = ( wire22  &  n_n730  &  (~ wire29)  &  wire146 ) ;
 assign wire566 = ( wire22  &  n_n918  &  (~ wire14)  &  wire146 ) ;
 assign wire567 = ( wire22  &  n_n1022  &  wire369 ) ;
 assign wire568 = ( n_n1187  &  n_n996  &  n_n1155  &  n_n698 ) ;
 assign wire569 = ( n_n1053  &  n_n992  &  wire293 ) ;
 assign wire570 = ( n_n1201  &  wire15  &  n_n1187  &  wire5884 ) ;
 assign wire571 = ( n_n1171  &  wire221  &  n_n992 ) | ( wire221  &  n_n992  &  wire47 ) ;
 assign wire572 = ( n_n1187  &  wire25  &  wire5886 ) | ( n_n1187  &  wire32  &  wire5886 ) ;
 assign wire573 = ( n_n1201  &  n_n1187  &  n_n996  &  wire29 ) ;
 assign wire575 = ( wire22  &  wire29  &  n_n1022 ) ;
 assign wire576 = ( wire22  &  wire14  &  n_n1084 ) ;
 assign wire577 = ( n_n904  &  wire22  &  n_n1022 ) ;
 assign wire579 = ( wire221  &  wire642 ) | ( n_n840  &  wire221  &  wire5813 ) ;
 assign wire580 = ( n_n1187  &  n_n996  &  wire25 ) | ( n_n1187  &  n_n996  &  wire32 ) ;
 assign wire581 = ( n_n996  &  wire219 ) | ( n_n996  &  wire1016 ) ;
 assign wire583 = ( g  &  h  &  i  &  wire113 ) ;
 assign wire585 = ( wire22  &  wire210  &  wire14  &  wire197 ) ;
 assign wire586 = ( wire22  &  n_n987  &  wire14  &  wire197 ) ;
 assign wire587 = ( n_n904  &  wire22  &  (~ n_n987)  &  wire197 ) ;
 assign wire588 = ( g  &  (~ j)  &  wire22  &  wire5857 ) ;
 assign wire590 = ( n_n711  &  n_n1142  &  wire70 ) ;
 assign wire593 = ( wire22  &  n_n920  &  n_n766 ) ;
 assign wire594 = ( wire210  &  wire70  &  n_n992 ) ;
 assign wire598 = ( n_n840  &  n_n1210  &  n_n1022 ) ;
 assign wire610 = ( n_n1201  &  n_n1187  &  wire29  &  n_n605 ) ;
 assign wire611 = ( wire299  &  wire5839 ) | ( wire41  &  wire5839 ) | ( wire1012  &  wire5839 ) ;
 assign wire617 = ( n_n1220  &  n_n698  &  n_n841 ) ;
 assign wire618 = ( n_n1187  &  n_n605  &  wire25 ) | ( n_n1187  &  n_n605  &  wire32 ) ;
 assign wire619 = ( n_n918  &  n_n1187  &  n_n1195  &  n_n605 ) ;
 assign wire626 = ( n_n700  &  wire290  &  n_n1227 ) ;
 assign wire627 = ( n_n1155  &  n_n1210  &  wire47 ) | ( n_n1155  &  n_n1210  &  wire60 ) ;
 assign wire628 = ( n_n711  &  n_n821  &  n_n1210 ) | ( n_n821  &  wire30  &  n_n1210 ) ;
 assign wire629 = ( n_n671  &  n_n1264  &  n_n1036 ) ;
 assign wire630 = ( n_n1210  &  n_n820  &  n_n1053 ) ;
 assign wire631 = ( n_n1171  &  n_n1219  &  n_n387 ) ;
 assign wire632 = ( wire30  &  n_n1142  &  wire70 ) ;
 assign wire633 = ( n_n709  &  n_n1210  &  wire231 ) ;
 assign wire635 = ( n_n840  &  n_n824  &  n_n1210 ) ;
 assign wire641 = ( b  &  d  &  (~ e)  &  wire5813 ) ;
 assign wire642 = ( (~ f)  &  h  &  i  &  n_n709 ) ;
 assign wire643 = ( n_n1080  &  n_n1190  &  n_n1039  &  wire386 ) ;
 assign wire644 = ( n_n838  &  (~ n_n1252)  &  n_n1210  &  wire89 ) ;
 assign wire645 = ( (~ g)  &  wire190  &  wire5781 ) ;
 assign wire646 = ( n_n1187  &  n_n949  &  n_n1252  &  wire165 ) ;
 assign wire647 = ( n_n842  &  n_n1210  &  wire164 ) ;
 assign wire649 = ( n_n1187  &  n_n949  &  n_n987  &  wire39 ) ;
 assign wire650 = ( n_n1187  &  n_n949  &  n_n977  &  n_n987 ) ;
 assign wire651 = ( n_n1210  &  n_n988  &  wire89 ) ;
 assign wire652 = ( n_n1217  &  n_n1080  &  n_n971  &  n_n1204 ) ;
 assign wire653 = ( (~ g)  &  wire224  &  wire190 ) ;
 assign wire655 = ( n_n872  &  wire5694 ) | ( wire148  &  n_n1104  &  n_n872 ) ;
 assign wire657 = ( wire111  &  wire743 ) | ( n_n1220  &  wire111  &  n_n1082 ) ;
 assign wire658 = ( n_n876  &  wire743 ) | ( n_n1220  &  n_n876  &  n_n1082 ) ;
 assign wire661 = ( n_n904  &  wire864 ) | ( n_n904  &  n_n940  &  wire190 ) ;
 assign wire663 = ( n_n1187  &  n_n949  &  wire69 ) | ( n_n1187  &  n_n949  &  wire1116 ) ;
 assign wire664 = ( n_n876  &  wire69 ) | ( wire31  &  n_n876  &  wire368 ) ;
 assign wire670 = ( n_n1252  &  wire283  &  wire301  &  n_n1253 ) ;
 assign wire671 = ( n_n1201  &  n_n1069  &  n_n1204  &  n_n1180 ) ;
 assign wire672 = ( n_n1207  &  n_n1229  &  n_n1190  &  n_n977 ) ;
 assign wire679 = ( wire76  &  n_n838  &  n_n1095  &  n_n1094 ) ;
 assign wire680 = ( wire58  &  n_n857  &  n_n872  &  (~ wire137) ) ;
 assign wire681 = ( n_n1161  &  wire84  &  n_n988 ) ;
 assign wire682 = ( n_n988  &  wire77  &  n_n1196 ) ;
 assign wire683 = ( n_n842  &  wire76  &  n_n841 ) ;
 assign wire684 = ( wire22  &  n_n857  &  n_n872 ) | ( n_n857  &  n_n872  &  wire113 ) ;
 assign wire699 = ( n_n904  &  n_n1187  &  wire74  &  n_n1252 ) ;
 assign wire700 = ( n_n904  &  n_n1187  &  n_n1252  &  wire20 ) ;
 assign wire701 = ( n_n904  &  n_n1187  &  n_n940  &  n_n942 ) ;
 assign wire702 = ( n_n1161  &  n_n1177  &  n_n893  &  n_n988 ) ;
 assign wire703 = ( n_n920  &  n_n1187  &  n_n1233  &  wire55 ) ;
 assign wire704 = ( n_n920  &  n_n1187  &  n_n1233  &  wire18 ) ;
 assign wire708 = ( n_n1187  &  n_n949  &  n_n1252  &  wire55 ) ;
 assign wire709 = ( n_n1187  &  n_n949  &  n_n987  &  n_n989 ) ;
 assign wire713 = ( wire417  &  wire1112  &  wire5690 ) | ( wire417  &  wire1113  &  wire5690 ) ;
 assign wire716 = ( wire120  &  wire183  &  n_n1231  &  (~ wire57) ) ;
 assign wire717 = ( wire44  &  (~ wire387)  &  (~ wire743)  &  wire5699 ) ;
 assign wire718 = ( n_n1165  &  n_n1138  &  n_n1142  &  n_n1146 ) ;
 assign wire719 = ( n_n1138  &  wire254  &  wire407 ) ;
 assign wire724 = ( n_n1220  &  n_n997  &  n_n1082 ) ;
 assign wire725 = ( wire390  &  n_n949 ) | ( n_n949  &  wire1068 ) | ( n_n949  &  wire5253 ) ;
 assign wire726 = ( wire58  &  n_n949  &  n_n765 ) ;
 assign wire727 = ( n_n761  &  wire1205 ) | ( (~ f)  &  n_n761  &  wire379 ) ;
 assign wire729 = ( n_n876  &  wire743 ) | ( n_n1220  &  n_n876  &  n_n1082 ) ;
 assign wire731 = ( n_n997  &  wire69 ) | ( wire31  &  n_n997  &  wire368 ) ;
 assign wire732 = ( n_n876  &  wire69 ) | ( wire31  &  n_n876  &  wire368 ) ;
 assign wire736 = ( wire22  &  n_n876  &  n_n859 ) ;
 assign wire739 = ( (~ f)  &  g  &  (~ h)  &  wire148 ) ;
 assign wire743 = ( e  &  h  &  k  &  n_n1219 ) ;
 assign wire745 = ( n_n1187  &  wire74  &  n_n1261  &  wire5674 ) ;
 assign wire749 = ( n_n1201  &  n_n1069  &  n_n1204  &  n_n1180 ) ;
 assign wire750 = ( n_n1187  &  wire74  &  n_n997  &  n_n1233 ) ;
 assign wire751 = ( m  &  (~ n)  &  wire92  &  n_n997 ) ;
 assign wire753 = ( n_n1039  &  wire5663  &  wire5664 ) ;
 assign wire754 = ( n_n1217  &  n_n1069  &  n_n971  &  n_n1204 ) ;
 assign wire762 = ( n_n1229  &  n_n1217  &  n_n1201  &  n_n1204 ) ;
 assign wire765 = ( n_n1252  &  n_n1264  &  n_n1253  &  n_n978 ) ;
 assign wire766 = ( (~ g)  &  n_n1138  &  n_n1159  &  wire226 ) ;
 assign wire767 = ( n_n1217  &  n_n1080  &  n_n971  &  n_n1204 ) ;
 assign wire775 = ( n_n1085  &  n_n1253  &  n_n982  &  n_n1249 ) ;
 assign wire776 = ( n_n1204  &  n_n973  &  n_n1180  &  n_n1195 ) ;
 assign wire777 = ( n_n987  &  n_n988  &  wire398  &  n_n982 ) ;
 assign wire780 = ( n_n1104  &  n_n1204  &  n_n975  &  wire5640 ) ;
 assign wire781 = ( n_n987  &  n_n988  &  n_n1085  &  n_n982 ) ;
 assign wire782 = ( n_n1204  &  n_n1180  &  n_n975  &  n_n1195 ) ;
 assign wire783 = ( n_n1207  &  n_n1165  &  n_n893  &  wire5587 ) ;
 assign wire784 = ( n_n1201  &  n_n1187  &  wire29  &  wire5590 ) ;
 assign wire785 = ( n_n1201  &  n_n1187  &  n_n698  &  wire5592 ) ;
 assign wire786 = ( wire148  &  wire29  &  n_n893  &  n_n1194 ) ;
 assign wire787 = ( wire148  &  n_n698  &  n_n893  &  n_n1194 ) ;
 assign wire788 = ( wire15  &  n_n1194  &  wire5598 ) ;
 assign wire789 = ( n_n1207  &  wire148  &  wire15  &  n_n1228 ) ;
 assign wire790 = ( n_n1187  &  wire25  &  wire5600 ) | ( n_n1187  &  wire32  &  wire5600 ) ;
 assign wire791 = ( n_n918  &  n_n1187  &  n_n1195  &  wire5601 ) ;
 assign wire796 = ( wire76  &  n_n841  &  wire93 ) ;
 assign wire797 = ( wire22  &  wire15  &  n_n1228 ) | ( wire15  &  wire113  &  n_n1228 ) ;
 assign wire798 = ( n_n1177  &  n_n893  &  wire841 ) | ( n_n1177  &  n_n893  &  wire5557 ) ;
 assign wire799 = ( wire371  &  wire33 ) | ( wire33  &  wire414 ) | ( wire33  &  wire80 ) ;
 assign wire802 = ( wire148  &  wire299 ) | ( wire148  &  wire41 ) | ( wire148  &  wire1012 ) ;
 assign wire808 = ( n_n1201  &  wire49  &  wire5526 ) ;
 assign wire809 = ( n_n1201  &  n_n844  &  wire5529 ) ;
 assign wire810 = ( n_n1207  &  n_n1116  &  wire5532 ) ;
 assign wire811 = ( wire58  &  n_n1171  &  wire5534 ) ;
 assign wire812 = ( b  &  (~ c)  &  n_n1148  &  wire293 ) ;
 assign wire813 = ( b  &  (~ c)  &  wire172  &  n_n1148 ) ;
 assign wire814 = ( b  &  (~ c)  &  wire77  &  n_n1148 ) ;
 assign wire815 = ( n_n713  &  n_n1196  &  wire293 ) ;
 assign wire816 = ( n_n840  &  n_n1201  &  wire293 ) ;
 assign wire817 = ( n_n1171  &  wire290  &  n_n868 ) ;
 assign wire818 = ( n_n841  &  wire260  &  wire109 ) ;
 assign wire821 = ( n_n713  &  wire172  &  n_n1196 ) ;
 assign wire822 = ( n_n840  &  wire172  &  n_n1201 ) ;
 assign wire823 = ( wire93  &  n_n1210  &  wire164 ) ;
 assign wire826 = ( n_n713  &  wire77  &  n_n1196 ) ;
 assign wire827 = ( n_n840  &  n_n1201  &  wire77 ) ;
 assign wire828 = ( wire54  &  n_n1171  &  n_n1142 ) ;
 assign wire829 = ( n_n1190  &  n_n817  &  wire24 ) ;
 assign wire830 = ( n_n698  &  n_n1219  &  n_n1131 ) ;
 assign wire831 = ( n_n700  &  n_n1190  &  n_n817 ) ;
 assign wire832 = ( n_n1203  &  n_n1190  &  n_n817 ) ;
 assign wire833 = ( n_n1171  &  n_n1219  &  n_n1131 ) ;
 assign wire834 = ( n_n1202  &  n_n1137  &  wire109 ) ;
 assign wire835 = ( n_n698  &  n_n841  &  n_n1215 ) ;
 assign wire836 = ( wire84  &  wire5557 ) | ( n_n840  &  n_n1207  &  wire84 ) ;
 assign wire837 = ( n_n1171  &  n_n841  &  n_n1215 ) ;
 assign wire841 = ( b  &  d  &  (~ e)  &  n_n1207 ) ;
 assign wire843 = ( (~ n_n1229)  &  wire74  &  wire120  &  wire5480 ) ;
 assign wire845 = ( wire74  &  wire120  &  wire196  &  wire5486 ) ;
 assign wire849 = ( n_n730  &  wire112  &  wire120  &  wire183 ) ;
 assign wire850 = ( wire76  &  n_n1095  &  wire5498 ) ;
 assign wire853 = ( n_n1165  &  n_n1203  &  n_n235 ) | ( n_n1165  &  n_n1203  &  wire65 ) ;
 assign wire854 = ( n_n842  &  wire84  &  n_n1104 ) ;
 assign wire858 = ( wire390  &  n_n730 ) | ( n_n730  &  wire1068 ) | ( n_n730  &  wire5253 ) ;
 assign wire859 = ( n_n920  &  n_n1187  &  wire74  &  n_n1233 ) ;
 assign wire860 = ( n_n876  &  wire864 ) | ( n_n876  &  n_n940  &  wire190 ) ;
 assign wire864 = ( e  &  f  &  h  &  wire22 ) ;
 assign wire869 = ( n_n842  &  n_n1177  &  n_n1252  &  n_n235 ) ;
 assign wire871 = ( wire390  &  wire43 ) | ( wire43  &  wire1068 ) | ( wire43  &  wire5253 ) ;
 assign wire875 = ( n_n1210  &  wire89  &  wire5454 ) ;
 assign wire879 = ( n_n1203  &  n_n1166  &  n_n1204 ) ;
 assign wire880 = ( n_n709  &  n_n1210  &  wire231 ) ;
 assign wire884 = ( n_n709  &  n_n1210  &  n_n662 ) ;
 assign wire886 = ( a  &  d  &  (~ e)  &  wire94 ) ;
 assign wire895 = ( (~ wire15)  &  wire228  &  n_n730  &  wire255 ) ;
 assign wire898 = ( n_n1165  &  n_n1155  &  n_n700  &  n_n1146 ) ;
 assign wire900 = ( n_n1207  &  n_n904  &  wire228  &  n_n1187 ) ;
 assign wire901 = ( n_n1207  &  wire228  &  n_n1187  &  wire29 ) ;
 assign wire902 = ( n_n1207  &  wire228  &  n_n1187  &  n_n698 ) ;
 assign wire903 = ( wire371  &  wire5422 ) | ( wire414  &  wire5422 ) | ( wire80  &  wire5422 ) ;
 assign wire904 = ( n_n1177  &  n_n1155  &  wire210  &  n_n1146 ) ;
 assign wire906 = ( n_n1177  &  n_n821  &  wire30  &  n_n1146 ) ;
 assign wire907 = ( n_n711  &  n_n1177  &  n_n821  &  n_n1146 ) ;
 assign wire908 = ( n_n1177  &  n_n1155  &  n_n1171  &  n_n1146 ) ;
 assign wire909 = ( n_n918  &  n_n1187  &  n_n996  &  n_n857 ) ;
 assign wire911 = ( n_n1187  &  wire380  &  wire25 ) | ( n_n1187  &  wire380  &  wire32 ) ;
 assign wire912 = ( wire54  &  n_n1155  &  wire219 ) | ( wire54  &  n_n1155  &  wire1016 ) ;
 assign wire914 = ( wire228  &  wire41 ) | ( n_n1161  &  n_n904  &  wire228 ) ;
 assign wire923 = ( n_n918  &  wire58  &  (~ wire137)  &  (~ n_n765) ) ;
 assign wire924 = ( n_n904  &  wire58  &  (~ n_n987)  &  (~ wire137) ) ;
 assign wire925 = ( n_n698  &  n_n694  &  wire142 ) ;
 assign wire926 = ( wire15  &  n_n1194  &  wire142 ) ;
 assign wire927 = ( wire54  &  wire15  &  n_n1194 ) ;
 assign wire928 = ( wire106  &  wire142 ) | ( wire50  &  wire142 ) | ( wire142  &  wire5313 ) ;
 assign wire929 = ( wire54  &  wire106 ) | ( wire54  &  wire50 ) | ( wire54  &  wire5313 ) ;
 assign wire931 = ( n_n711  &  (~ wire30)  &  n_n982  &  wire56 ) ;
 assign wire932 = ( n_n1202  &  n_n1137  &  wire5367 ) ;
 assign wire934 = ( n_n700  &  n_n841  &  wire260 ) ;
 assign wire935 = ( n_n1171  &  n_n1215  &  wire216 ) ;
 assign wire938 = ( n_n1171  &  n_n694  &  wire142 ) ;
 assign wire939 = ( n_n1137  &  n_n982  &  wire47 ) ;
 assign wire940 = ( wire30  &  n_n818  &  n_n982 ) ;
 assign wire941 = ( n_n709  &  n_n1084  &  n_n978 ) ;
 assign wire942 = ( n_n840  &  n_n1022  &  n_n978 ) ;
 assign wire943 = ( n_n698  &  n_n1215  &  wire216 ) ;
 assign wire945 = ( n_n1094  &  n_n978  &  n_n703 ) ;
 assign wire948 = ( n_n671  &  n_n618  &  n_n1216 ) ;
 assign wire951 = ( n_n982  &  wire1042 ) | ( n_n840  &  n_n823  &  n_n982 ) ;
 assign wire952 = ( n_n1171  &  n_n841  &  n_n978 ) ;
 assign wire954 = ( n_n619  &  wire960 ) | ( n_n619  &  n_n1216  &  n_n623 ) ;
 assign wire960 = ( wire34  &  n_n1204 ) | ( n_n1204  &  wire35 ) ;
 assign wire961 = ( l  &  (~ m)  &  n  &  n_n623 ) ;
 assign wire962 = ( g  &  (~ h)  &  wire228  &  n_n1171 ) ;
 assign wire963 = ( (~ f)  &  wire58  &  wire14  &  (~ wire137) ) ;
 assign wire965 = ( n_n709  &  wire76  &  n_n662 ) ;
 assign wire966 = ( n_n840  &  wire76  &  n_n1095 ) ;
 assign wire967 = ( wire76  &  n_n841  &  n_n1053 ) ;
 assign wire968 = ( n_n841  &  n_n978  &  wire47 ) ;
 assign wire969 = ( n_n709  &  n_n662  &  n_n978 ) ;
 assign wire970 = ( n_n1053  &  n_n1137  &  n_n982 ) ;
 assign wire971 = ( n_n820  &  n_n1053  &  n_n978 ) ;
 assign wire972 = ( n_n671  &  n_n670  &  n_n978 ) ;
 assign wire973 = ( n_n840  &  n_n1095  &  n_n978 ) ;
 assign wire974 = ( n_n711  &  n_n1094  &  n_n978 ) ;
 assign wire975 = ( n_n841  &  n_n1053  &  n_n978 ) ;
 assign wire976 = ( n_n838  &  n_n1094  &  n_n978 ) ;
 assign wire977 = ( wire76  &  wire980 ) | ( n_n1171  &  wire76  &  n_n841 ) ;
 assign wire978 = ( wire58  &  n_n730  &  n_n765 ) ;
 assign wire980 = ( n_n711  &  n_n1094 ) | ( wire30  &  n_n1094 ) ;
 assign wire982 = ( wire15  &  n_n1194  &  wire5309 ) ;
 assign wire983 = ( n_n1201  &  wire15  &  wire265 ) ;
 assign wire985 = ( n_n1217  &  n_n1220  &  n_n698  &  n_n841 ) ;
 assign wire986 = ( wire106  &  wire5314 ) | ( wire50  &  wire5314 ) | ( wire5313  &  wire5314 ) ;
 assign wire989 = ( wire299  &  wire5317 ) | ( wire41  &  wire5317 ) | ( wire1012  &  wire5317 ) ;
 assign wire990 = ( wire299  &  wire5318 ) | ( wire41  &  wire5318 ) | ( wire1012  &  wire5318 ) ;
 assign wire991 = ( n_n918  &  wire228  &  n_n861 ) | ( n_n918  &  wire265  &  n_n861 ) ;
 assign wire992 = ( n_n1193  &  wire15  &  wire228 ) | ( n_n1193  &  wire15  &  wire265 ) ;
 assign wire993 = ( n_n1193  &  n_n920  &  wire228 ) | ( n_n1193  &  n_n920  &  wire265 ) ;
 assign wire994 = ( wire265  &  n_n698  &  n_n1137 ) ;
 assign wire995 = ( wire265  &  n_n1187  &  wire25 ) | ( wire265  &  n_n1187  &  wire32 ) ;
 assign wire997 = ( wire228  &  wire5289 ) | ( wire228  &  wire14  &  n_n861 ) ;
 assign wire1012 = ( f  &  g  &  (~ h)  &  wire16 ) ;
 assign wire1016 = ( m  &  (~ n)  &  n_n1201  &  n_n920 ) ;
 assign wire1018 = ( wire59  &  wire1039  &  wire5271 ) | ( wire59  &  wire5270  &  wire5271 ) ;
 assign wire1019 = ( wire23  &  wire47  &  wire5274 ) | ( wire23  &  wire60  &  wire5274 ) ;
 assign wire1020 = ( j  &  n_n709  &  n_n1210  &  wire5277 ) ;
 assign wire1021 = ( n_n711  &  wire134  &  wire5279 ) | ( wire30  &  wire134  &  wire5279 ) ;
 assign wire1022 = ( j  &  n_n700  &  n_n1191  &  wire23 ) ;
 assign wire1023 = ( n_n1036  &  n_n1137  &  wire47 ) | ( n_n1036  &  n_n1137  &  wire60 ) ;
 assign wire1024 = ( j  &  n_n840  &  n_n1210  &  wire59 ) ;
 assign wire1027 = ( n_n711  &  n_n1036  &  n_n818 ) | ( wire30  &  n_n1036  &  n_n818 ) ;
 assign wire1030 = ( n_n700  &  n_n1202  &  n_n1137 ) ;
 assign wire1031 = ( wire34  &  n_n1191  &  wire398 ) | ( n_n1191  &  wire398  &  wire35 ) ;
 assign wire1032 = ( wire34  &  n_n1191  &  n_n670 ) | ( n_n1191  &  n_n670  &  wire35 ) ;
 assign wire1033 = ( wire265  &  n_n1171  &  n_n1137 ) ;
 assign wire1034 = ( wire265  &  wire5289 ) | ( wire265  &  wire14  &  n_n861 ) ;
 assign wire1036 = ( n_n617  &  wire1039 ) | ( n_n617  &  wire5270 ) ;
 assign wire1039 = ( (~ m)  &  (~ n)  &  wire34 ) | ( (~ m)  &  (~ n)  &  wire35 ) ;
 assign wire1042 = ( (~ f)  &  h  &  j  &  n_n709 ) ;
 assign wire1043 = ( b  &  d  &  (~ e)  &  n_n823 ) ;
 assign wire1051 = ( n_n1229  &  n_n235  &  wire5246 ) | ( n_n1229  &  wire65  &  wire5246 ) ;
 assign wire1052 = ( n_n1165  &  (~ wire232)  &  n_n235 ) | ( n_n1165  &  (~ wire232)  &  wire65 ) ;
 assign wire1053 = ( n_n1165  &  n_n1101  &  n_n235 ) | ( n_n1165  &  n_n1101  &  wire65 ) ;
 assign wire1054 = ( n_n1177  &  n_n671  &  n_n235 ) | ( n_n1177  &  n_n671  &  wire65 ) ;
 assign wire1055 = ( n_n904  &  wire54  &  wire5220 ) ;
 assign wire1057 = ( wire84  &  wire393 ) | ( wire84  &  n_n1160  &  n_n1253 ) ;
 assign wire1058 = ( wire172  &  wire377 ) | ( wire172  &  wire115 ) ;
 assign wire1059 = ( n_n904  &  wire58  &  n_n765 ) ;
 assign wire1060 = ( n_n626  &  wire5088 ) | ( n_n626  &  n_n816  &  n_n1056 ) ;
 assign wire1061 = ( a  &  (~ c)  &  d  &  wire138 ) ;
 assign wire1062 = ( n_n904  &  wire5253 ) | ( n_n904  &  n_n874  &  wire5252 ) ;
 assign wire1068 = ( i  &  l  &  m  &  wire5252 ) ;
 assign wire1070 = ( n_n1220  &  n_n1082  &  wire5213 ) ;
 assign wire1071 = ( n_n1166  &  n_n1204  &  n_n973  &  n_n1095 ) ;
 assign wire1074 = ( n_n626  &  n_n1210  &  wire134 ) ;
 assign wire1075 = ( n_n626  &  wire76  &  n_n1094 ) ;
 assign wire1076 = ( n_n973  &  n_n1095  &  n_n1191 ) ;
 assign wire1077 = ( n_n1229  &  n_n1166  &  n_n1204  &  n_n662 ) ;
 assign wire1078 = ( n_n1229  &  n_n662  &  n_n1191 ) ;
 assign wire1079 = ( n_n904  &  n_n1220  &  wire5220 ) ;
 assign wire1080 = ( n_n1101  &  n_n1166  &  n_n1204 ) ;
 assign wire1081 = ( n_n671  &  n_n1166  &  n_n1216 ) ;
 assign wire1082 = ( wire293  &  wire377 ) | ( wire293  &  wire115 ) ;
 assign wire1083 = ( wire77  &  wire377 ) | ( wire77  &  wire115 ) ;
 assign wire1084 = ( a  &  (~ c)  &  d  &  wire94 ) ;
 assign wire1096 = ( wire175  &  n_n918  &  n_n1187  &  n_n816 ) ;
 assign wire1100 = ( n_n1187  &  n_n949  &  n_n816  &  wire90 ) ;
 assign wire1102 = ( n_n1187  &  n_n949  &  n_n942  &  n_n912 ) ;
 assign wire1106 = ( wire393  &  n_n1177  &  n_n893 ) | ( n_n1177  &  n_n893  &  wire1110 ) ;
 assign wire1110 = ( (~ e)  &  f  &  (~ h)  &  n_n1253 ) ;
 assign wire1112 = ( wire228  &  n_n864 ) | ( wire265  &  n_n864 ) ;
 assign wire1113 = ( wire22  &  n_n859 ) | ( wire113  &  n_n859 ) ;
 assign wire1116 = ( wire31  &  wire368 ) ;
 assign wire1122 = ( wire84  &  (~ wire175)  &  (~ wire229)  &  wire5140 ) ;
 assign wire1123 = ( (~ g)  &  wire53  &  wire224  &  wire190 ) ;
 assign wire1124 = ( wire76  &  n_n1095  &  wire5144 ) ;
 assign wire1126 = ( g  &  wire233  &  wire1147 ) | ( g  &  wire233  &  wire1148 ) ;
 assign wire1128 = ( n_n711  &  n_n886  &  wire172 ) ;
 assign wire1129 = ( n_n709  &  n_n1188  &  wire148 ) ;
 assign wire1130 = ( n_n1089  &  n_n842  &  wire84 ) ;
 assign wire1131 = ( n_n1161  &  n_n713  &  n_n1177  &  n_n893 ) ;
 assign wire1135 = ( wire76  &  n_n1095  &  n_n1094  &  n_n703 ) ;
 assign wire1137 = ( n_n840  &  wire76  &  n_n1095 ) ;
 assign wire1138 = ( wire153  &  wire72 ) | ( wire153  &  wire1198 ) | ( wire153  &  wire1200 ) ;
 assign wire1139 = ( n_n709  &  wire72 ) | ( n_n709  &  wire1198 ) | ( n_n709  &  wire1200 ) ;
 assign wire1140 = ( wire172  &  wire5116 ) | ( n_n842  &  wire172  &  n_n1201 ) ;
 assign wire1141 = ( wire46  &  wire1147 ) | ( wire46  &  wire1148 ) ;
 assign wire1145 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire1147 = ( (~ d)  &  e  &  n_n1187  &  n_n1261 ) ;
 assign wire1148 = ( (~ e)  &  m  &  (~ n)  &  n_n918 ) ;
 assign wire1155 = ( g  &  n_n711  &  wire172  &  wire71 ) ;
 assign wire1156 = ( n_n709  &  n_n1201  &  wire293 ) ;
 assign wire1157 = ( (~ m)  &  (~ n)  &  n_n626  &  wire198 ) ;
 assign wire1158 = ( n_n709  &  wire172  &  n_n1201 ) ;
 assign wire1161 = ( n_n628  &  wire65  &  wire162 ) ;
 assign wire1162 = ( n_n709  &  n_n1201  &  wire77 ) ;
 assign wire1163 = ( n_n840  &  wire77  &  n_n822 ) ;
 assign wire1166 = ( n_n1191  &  n_n628  &  n_n235 ) ;
 assign wire1167 = ( n_n1229  &  n_n662  &  n_n1191 ) ;
 assign wire1168 = ( g  &  n_n711  &  wire71  &  wire293 ) | ( (~ g)  &  n_n711  &  wire71  &  wire293 ) ;
 assign wire1169 = ( g  &  n_n711  &  wire71  &  wire77 ) | ( (~ g)  &  n_n711  &  wire71  &  wire77 ) ;
 assign wire1170 = ( m  &  (~ n)  &  n_n698  &  n_n816 ) ;
 assign wire1171 = ( n_n1229  &  n_n1190  &  n_n825 ) ;
 assign wire1172 = ( n_n713  &  n_n886  &  wire172 ) ;
 assign wire1173 = ( n_n626  &  n_n1166  &  n_n1204 ) ;
 assign wire1175 = ( wire293  &  wire5116 ) | ( n_n842  &  n_n1201  &  wire293 ) ;
 assign wire1176 = ( wire77  &  wire5116 ) | ( n_n842  &  n_n1201  &  wire77 ) ;
 assign wire1185 = ( n_n709  &  n_n1219  &  n_n825 ) ;
 assign wire1186 = ( n_n821  &  n_n1210  &  n_n703 ) ;
 assign wire1187 = ( n_n840  &  n_n1036  &  n_n823 ) ;
 assign wire1188 = ( n_n709  &  wire228  &  n_n861 ) | ( n_n709  &  wire265  &  n_n861 ) ;
 assign wire1189 = ( n_n1229  &  n_n662  &  wire260 ) ;
 assign wire1192 = ( n_n698  &  n_n1219  &  n_n1137 ) ;
 assign wire1193 = ( n_n1210  &  n_n1094  &  n_n703 ) ;
 assign wire1194 = ( n_n840  &  n_n1210  &  wire89 ) ;
 assign wire1195 = ( n_n698  &  wire72 ) | ( n_n698  &  wire1198 ) | ( n_n698  &  wire1200 ) ;
 assign wire1196 = ( n_n709  &  wire1205 ) | ( (~ f)  &  n_n709  &  wire379 ) ;
 assign wire1197 = ( n_n703  &  wire5088 ) | ( n_n816  &  n_n1056  &  n_n703 ) ;
 assign wire1198 = ( g  &  (~ i)  &  j  &  wire96 ) ;
 assign wire1200 = ( (~ l)  &  m  &  (~ n)  &  n_n1131 ) ;
 assign wire1205 = ( wire22  &  n_n857 ) | ( n_n857  &  wire113 ) ;
 assign wire5088 = ( k  &  n_n1177  &  n_n819 ) | ( (~ k)  &  n_n1177  &  n_n818 ) ;
 assign wire5091 = ( n_n698  &  wire23  &  n_n1215 ) | ( n_n698  &  n_n1215  &  wire105 ) ;
 assign wire5093 = ( wire1185 ) | ( wire1186 ) | ( wire1194 ) ;
 assign wire5094 = ( wire1187 ) | ( wire1189 ) | ( wire5091 ) ;
 assign wire5095 = ( wire1188 ) | ( wire1192 ) | ( wire1193 ) ;
 assign wire5098 = ( wire1195 ) | ( wire1197 ) | ( wire5093 ) ;
 assign wire5099 = ( wire1196 ) | ( wire5094 ) | ( wire5095 ) ;
 assign wire5108 = ( c  &  (~ e)  &  f  &  wire65 ) ;
 assign wire5116 = ( n_n842  &  n_n1194 ) | ( n_n713  &  n_n1196 ) ;
 assign wire5117 = ( n_n709  &  n_n868  &  wire385 ) | ( n_n709  &  n_n871  &  wire385 ) ;
 assign wire5120 = ( n_n709  &  wire54  &  n_n971 ) | ( n_n709  &  n_n1220  &  n_n971 ) ;
 assign wire5124 = ( wire1155 ) | ( n_n1166  &  n_n1204  &  n_n628 ) ;
 assign wire5125 = ( wire1156 ) | ( n_n1229  &  wire71  &  wire162 ) ;
 assign wire5126 = ( wire1169 ) | ( wire1168 ) ;
 assign wire5127 = ( wire1157 ) | ( wire1158 ) | ( wire5117 ) ;
 assign wire5128 = ( wire1162 ) | ( wire1163 ) | ( wire5120 ) ;
 assign wire5129 = ( wire1166 ) | ( wire1167 ) | ( wire1170 ) | ( wire1171 ) ;
 assign wire5130 = ( wire1172 ) | ( wire1173 ) | ( wire162  &  wire5108 ) ;
 assign wire5136 = ( wire1161 ) | ( wire1175 ) | ( wire1176 ) | ( wire5124 ) ;
 assign wire5137 = ( wire5125 ) | ( wire5126 ) | ( wire5127 ) | ( wire5128 ) ;
 assign wire5139 = ( wire5129 ) | ( wire5130 ) | ( wire5136 ) | ( wire5137 ) ;
 assign wire5140 = ( b  &  c  &  (~ d)  &  (~ h) ) ;
 assign wire5144 = ( b  &  (~ c)  &  d ) ;
 assign wire5146 = ( wire202  &  wire76  &  n_n1095 ) ;
 assign wire5156 = ( (~ d)  &  e  &  n_n920  &  n_n1187 ) ;
 assign wire5159 = ( wire1123 ) | ( wire1122 ) ;
 assign wire5160 = ( wire1124 ) | ( n_n1207  &  wire84  &  wire202 ) ;
 assign wire5161 = ( wire84  &  wire393 ) | ( wire393  &  n_n1177  &  n_n893 ) ;
 assign wire5162 = ( wire1135 ) | ( (~ g)  &  wire153  &  wire190 ) ;
 assign wire5163 = ( wire1128 ) | ( wire1129 ) | ( wire1137 ) ;
 assign wire5169 = ( wire1126 ) | ( wire1130 ) | ( wire1131 ) | ( wire1141 ) ;
 assign wire5170 = ( wire1140 ) | ( wire5159 ) | ( wire5160 ) | ( wire5161 ) ;
 assign wire5171 = ( wire1138 ) | ( wire5162 ) | ( wire5163 ) ;
 assign wire5172 = ( wire1139 ) | ( wire46  &  wire5146 ) | ( wire46  &  wire5156 ) ;
 assign wire5175 = ( wire5169 ) | ( wire5170 ) | ( wire5171 ) | ( wire5172 ) ;
 assign wire5176 = ( (~ d)  &  n_n1215 ) | ( (~ e)  &  n_n1215 ) ;
 assign wire5177 = ( m  &  (~ n)  &  n_n918  &  wire105 ) ;
 assign wire5179 = ( (~ m)  &  n  &  n_n713  &  n_n1231 ) ;
 assign wire5181 = ( n_n713  &  n_n1177  &  n_n893  &  n_n1231 ) ;
 assign wire5183 = ( m  &  (~ n)  &  n_n949  &  wire90 ) ;
 assign wire5184 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5187 = ( m  &  (~ n)  &  n_n949  &  wire90 ) ;
 assign wire5188 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5190 = ( m  &  (~ n)  &  n_n949  &  n_n1231 ) ;
 assign wire5191 = ( m  &  (~ n)  &  n_n949  &  wire90 ) ;
 assign wire5192 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5194 = ( m  &  (~ n)  &  n_n949  &  n_n1231 ) ;
 assign wire5197 = ( wire5176  &  wire5177 ) | ( wire20  &  wire5181 ) ;
 assign wire5198 = ( wire1096 ) | ( n_n1187  &  n_n949  &  wire108 ) ;
 assign wire5199 = ( wire1100 ) | ( wire1102 ) | ( wire101  &  wire5179 ) ;
 assign wire5201 = ( wire181  &  wire388 ) | ( wire152  &  wire5190 ) ;
 assign wire5204 = ( wire1112  &  wire5187 ) | ( wire1113  &  wire5187 ) | ( wire1112  &  wire5188 ) | ( wire1113  &  wire5188 ) ;
 assign wire5205 = ( wire69  &  wire5191 ) | ( wire1116  &  wire5191 ) | ( wire69  &  wire5192 ) | ( wire1116  &  wire5192 ) ;
 assign wire5207 = ( wire5199 ) | ( wire379  &  wire5183 ) | ( wire379  &  wire5184 ) ;
 assign wire5208 = ( wire1106 ) | ( wire5201 ) | ( wire152  &  wire299 ) ;
 assign wire5209 = ( wire5197 ) | ( wire5198 ) | ( wire5204 ) ;
 assign wire5210 = ( wire5205 ) | ( wire74  &  wire388 ) | ( wire74  &  wire5194 ) ;
 assign wire5213 = ( (~ a)  &  b  &  d ) ;
 assign wire5215 = ( a  &  (~ c)  &  d  &  (~ e) ) ;
 assign wire5216 = ( (~ a)  &  b  &  d  &  e ) ;
 assign wire5220 = ( (~ e)  &  (~ g)  &  h ) ;
 assign wire5226 = ( n_n1219  &  wire121  &  wire5215 ) | ( n_n1219  &  wire121  &  wire5216 ) ;
 assign wire5227 = ( wire1070 ) | ( wire1071 ) | ( wire1074 ) | ( wire1075 ) ;
 assign wire5228 = ( wire1076 ) | ( wire1077 ) | ( wire1078 ) | ( wire1079 ) ;
 assign wire5232 = ( wire1080 ) | ( wire1081 ) | ( wire1082 ) | ( wire5228 ) ;
 assign wire5233 = ( wire1083 ) | ( wire1084 ) | ( wire5226 ) | ( wire5227 ) ;
 assign wire5234 = ( (~ n)  &  (~ i) ) ;
 assign wire5237 = ( n_n904  &  (~ wire22)  &  wire128  &  wire5234 ) ;
 assign wire5238 = ( a  &  (~ c)  &  d  &  (~ n) ) ;
 assign wire5241 = ( n_n1193  &  (~ wire22)  &  wire5238 ) ;
 assign wire5242 = ( m  &  (~ n) ) ;
 assign wire5243 = ( i  &  n_n904  &  wire128  &  wire5242 ) ;
 assign wire5244 = ( (~ f)  &  h  &  wire54 ) ;
 assign wire5246 = ( (~ f)  &  h  &  (~ m)  &  (~ n) ) ;
 assign wire5251 = ( f  &  g  &  h  &  (~ n) ) ;
 assign wire5252 = ( f  &  g  &  (~ h)  &  (~ n) ) ;
 assign wire5253 = ( wire54  &  n_n1194 ) | ( wire31  &  wire5251 ) ;
 assign wire5255 = ( wire31  &  (~ wire54)  &  wire5237 ) | ( wire31  &  (~ wire54)  &  wire5241 ) ;
 assign wire5256 = ( wire45  &  wire258 ) | ( wire31  &  wire258  &  wire5244 ) ;
 assign wire5257 = ( wire1055 ) | ( wire1059 ) | ( wire101  &  wire5243 ) ;
 assign wire5264 = ( wire1051 ) | ( wire1052 ) | ( wire1053 ) | ( wire1054 ) ;
 assign wire5265 = ( wire1057 ) | ( wire1058 ) | ( wire1060 ) | ( wire1061 ) ;
 assign wire5266 = ( wire1062 ) | ( wire5255 ) | ( wire5256 ) | ( wire5257 ) ;
 assign wire5268 = ( wire5232 ) | ( wire5233 ) | ( wire5266 ) ;
 assign wire5270 = ( (~ m)  &  n  &  n_n671 ) | ( (~ m)  &  n  &  n_n623 ) ;
 assign wire5271 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire5274 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire5277 = ( (~ f)  &  (~ g)  &  (~ h)  &  i ) | ( (~ f)  &  (~ g)  &  h  &  (~ i) ) ;
 assign wire5279 = ( j  &  k  &  (~ m)  &  n ) ;
 assign wire5289 = ( n_n876  &  n_n864 ) | ( n_n1193  &  wire16 ) ;
 assign wire5290 = ( n_n1171  &  n_n529  &  wire96 ) | ( n_n698  &  n_n529  &  wire96 ) ;
 assign wire5291 = ( n_n1220  &  n_n1171  &  n_n818 ) | ( n_n1220  &  n_n698  &  n_n818 ) ;
 assign wire5293 = ( wire58  &  n_n1171  &  n_n841 ) | ( wire58  &  n_n698  &  n_n841 ) ;
 assign wire5297 = ( wire1030 ) | ( wire1033 ) | ( wire5291 ) ;
 assign wire5298 = ( wire1019 ) | ( wire5293 ) ;
 assign wire5299 = ( wire1023 ) | ( n_n1036  &  wire1042 ) | ( n_n1036  &  wire1043 ) ;
 assign wire5300 = ( wire1020 ) | ( wire1021 ) | ( wire1022 ) | ( wire1024 ) ;
 assign wire5305 = ( wire1018 ) | ( wire1027 ) | ( wire5290 ) | ( wire5297 ) ;
 assign wire5306 = ( wire1031 ) | ( wire1032 ) | ( wire1036 ) ;
 assign wire5307 = ( wire1034 ) | ( wire5298 ) | ( wire5299 ) | ( wire5300 ) ;
 assign wire5309 = ( j  &  k  &  m  &  (~ n) ) ;
 assign wire5311 = ( (~ e)  &  g  &  (~ i)  &  n_n904 ) ;
 assign wire5313 = ( n_n904  &  n_n1194 ) | ( n_n730  &  n_n1194 ) | ( n_n904  &  wire5220 ) ;
 assign wire5314 = ( j  &  k  &  m  &  (~ n) ) ;
 assign wire5316 = ( k  &  m  &  (~ n)  &  n_n1217 ) ;
 assign wire5317 = ( wire58  &  i ) ;
 assign wire5318 = ( k  &  m  &  (~ n)  &  n_n1217 ) ;
 assign wire5321 = ( wire985 ) | ( wire994 ) | ( wire130  &  wire5311 ) ;
 assign wire5323 = ( wire993 ) | ( wire265  &  wire219 ) | ( wire265  &  wire1016 ) ;
 assign wire5325 = ( wire98  &  wire5316 ) | ( i  &  wire58  &  wire98 ) ;
 assign wire5327 = ( wire982 ) | ( wire983 ) | ( wire5321 ) | ( wire5323 ) ;
 assign wire5328 = ( wire989 ) | ( wire986 ) ;
 assign wire5329 = ( wire995 ) | ( wire990 ) ;
 assign wire5330 = ( wire991 ) | ( wire992 ) | ( wire997 ) | ( wire5325 ) ;
 assign wire5333 = ( wire5327 ) | ( wire5328 ) | ( wire5329 ) | ( wire5330 ) ;
 assign wire5356 = ( wire963 ) | ( wire76  &  n_n841  &  wire47 ) ;
 assign wire5357 = ( n_n2660 ) | ( wire962 ) | ( wire968 ) ;
 assign wire5358 = ( wire965 ) | ( wire966 ) | ( wire967 ) | ( wire969 ) ;
 assign wire5359 = ( wire970 ) | ( wire971 ) | ( wire972 ) | ( wire973 ) ;
 assign wire5360 = ( wire974 ) | ( wire975 ) | ( wire976 ) | ( wire978 ) ;
 assign wire5364 = ( wire5356 ) | ( wire5357 ) | ( wire5358 ) | ( wire5359 ) ;
 assign wire5367 = ( (~ c)  &  d  &  (~ e)  &  l ) ;
 assign wire5368 = ( k  &  (~ m)  &  n_n670 ) ;
 assign wire5379 = ( n_n700  &  n_n841  &  wire188 ) | ( n_n700  &  n_n820  &  wire188 ) ;
 assign wire5382 = ( n_n671  &  n_n1166  &  n_n1216 ) | ( n_n671  &  n_n1216  &  wire56 ) ;
 assign wire5386 = ( wire932 ) | ( wire934 ) | ( wire943 ) ;
 assign wire5387 = ( wire938 ) | ( wire941 ) | ( wire5379 ) ;
 assign wire5388 = ( wire942 ) | ( wire945 ) | ( wire5382 ) ;
 assign wire5389 = ( wire948 ) | ( wire952 ) | ( wire380  &  wire208 ) ;
 assign wire5391 = ( wire931 ) | ( wire935 ) | ( wire939 ) | ( wire940 ) ;
 assign wire5394 = ( wire951 ) | ( wire5389 ) | ( wire208  &  n_n978 ) ;
 assign wire5395 = ( wire5386 ) | ( wire5387 ) | ( wire5391 ) ;
 assign wire5396 = ( n_n1166  &  wire960 ) | ( n_n1166  &  wire961 ) | ( wire960  &  wire5368 ) | ( wire961  &  wire5368 ) ;
 assign wire5397 = ( wire954 ) | ( wire5388 ) | ( wire211  &  n_n978 ) ;
 assign wire5399 = ( wire977 ) | ( wire5360 ) | ( wire5364 ) | ( wire5396 ) ;
 assign wire5400 = ( wire5394 ) | ( wire5395 ) | ( wire5397 ) ;
 assign wire5406 = ( wire927 ) | ( wire58  &  wire29  &  n_n765 ) ;
 assign wire5407 = ( wire923 ) | ( wire924 ) | ( wire925 ) | ( wire926 ) ;
 assign wire5413 = ( f  &  h  &  (~ i)  &  wire30 ) ;
 assign wire5414 = ( (~ m)  &  n  &  wire34  &  n_n1146 ) ;
 assign wire5415 = ( g  &  n_n709 ) | ( (~ h)  &  n_n709 ) | ( i  &  n_n709 ) ;
 assign wire5416 = ( (~ m)  &  n  &  n_n824  &  n_n1146 ) ;
 assign wire5418 = ( (~ m)  &  n  &  n_n933  &  n_n1146 ) ;
 assign wire5422 = ( m  &  (~ n)  &  n_n996 ) ;
 assign wire5424 = ( m  &  (~ n)  &  wire29 ) ;
 assign wire5431 = ( wire895 ) | ( wire54  &  n_n1155  &  n_n698 ) ;
 assign wire5432 = ( wire5415  &  wire5416 ) | ( wire309  &  wire5418 ) ;
 assign wire5433 = ( wire901 ) | ( wire900 ) ;
 assign wire5435 = ( wire906 ) | ( wire54  &  n_n1155  &  wire291 ) ;
 assign wire5436 = ( wire898 ) | ( wire907 ) | ( wire908 ) | ( wire909 ) ;
 assign wire5437 = ( wire5413  &  wire5414 ) | ( wire179  &  wire5424 ) ;
 assign wire5443 = ( wire912 ) | ( wire5431 ) | ( wire5432 ) | ( wire5433 ) ;
 assign wire5444 = ( wire902 ) | ( wire904 ) | ( wire911 ) | ( wire5435 ) ;
 assign wire5445 = ( n_n617  &  wire960 ) | ( n_n618  &  wire960 ) | ( n_n617  &  wire961 ) | ( n_n618  &  wire961 ) ;
 assign wire5446 = ( wire903 ) | ( wire914 ) | ( wire5436 ) | ( wire5437 ) ;
 assign wire5448 = ( wire5446 ) | ( wire5445 ) ;
 assign wire5449 = ( n_n1792 ) | ( wire5443 ) | ( wire5444 ) ;
 assign wire5451 = ( (~ c)  &  e ) | ( (~ d)  &  e ) ;
 assign wire5453 = ( n_n1166  &  n_n1204  &  wire5451 ) ;
 assign wire5454 = ( (~ b)  &  c  &  e ) ;
 assign wire5456 = ( (~ b)  &  c  &  e ) ;
 assign wire5457 = ( n_n709  &  wire71  &  wire77 ) | ( n_n709  &  wire71  &  wire227 ) ;
 assign wire5459 = ( wire884 ) | ( (~ n_n1069)  &  n_n1095  &  wire5453 ) ;
 assign wire5460 = ( wire875 ) | ( n_n709  &  n_n1210  &  wire164 ) ;
 assign wire5461 = ( wire879 ) | ( wire880 ) | ( wire5457 ) ;
 assign wire5462 = ( wire184  &  wire77 ) | ( wire117  &  wire5456 ) ;
 assign wire5463 = ( n_n709  &  wire135 ) | ( wire94  &  wire43 ) ;
 assign wire5467 = ( wire886 ) | ( wire5459 ) | ( wire5460 ) | ( wire5461 ) ;
 assign wire5469 = ( a  &  (~ b)  &  d  &  f ) ;
 assign wire5474 = ( wire44  &  wire5469 ) | ( (~ n_n842)  &  wire224  &  wire44 ) ;
 assign wire5475 = ( wire869 ) | ( wire138  &  wire43 ) | ( wire195  &  wire43 ) ;
 assign wire5477 = ( b  &  (~ c) ) | ( b  &  (~ e) ) | ( (~ c)  &  (~ f) ) | ( (~ e)  &  (~ f) ) ;
 assign wire5479 = ( (~ n_n709)  &  wire229  &  wire5477 ) ;
 assign wire5480 = ( c  &  e  &  f  &  g ) ;
 assign wire5485 = ( wire229  &  n_n1165  &  (~ n_n1229)  &  (~ n_n1069) ) ;
 assign wire5486 = ( d  &  f  &  g ) ;
 assign wire5489 = ( (~ f)  &  n_n842 ) | ( (~ g)  &  n_n842 ) ;
 assign wire5490 = ( (~ m)  &  n  &  n_n1166  &  n_n893 ) ;
 assign wire5493 = ( (~ m)  &  n  &  n_n842  &  wire229 ) ;
 assign wire5495 = ( (~ b)  &  d  &  f  &  wire120 ) ;
 assign wire5498 = ( (~ b)  &  c  &  e  &  f ) ;
 assign wire5499 = ( (~ d)  &  f  &  (~ g) ) ;
 assign wire5505 = ( wire854 ) | ( wire76  &  n_n1095  &  wire5479 ) ;
 assign wire5506 = ( wire850 ) | ( n_n709  &  wire76  &  wire230 ) ;
 assign wire5507 = ( wire84  &  wire393 ) | ( wire393  &  n_n1177  &  n_n893 ) ;
 assign wire5508 = ( n_n235  &  wire5485 ) | ( wire65  &  wire5485 ) | ( n_n235  &  wire5493 ) | ( wire65  &  wire5493 ) ;
 assign wire5509 = ( wire853 ) | ( n  &  wire184  &  wire49 ) ;
 assign wire5513 = ( wire46  &  wire5495 ) | ( wire46  &  wire5489  &  wire5490 ) ;
 assign wire5514 = ( wire849 ) | ( wire92  &  wire120  &  wire256 ) ;
 assign wire5515 = ( wire859 ) | ( n_n920  &  n_n1187  &  wire92 ) ;
 assign wire5517 = ( wire860 ) | ( wire5505 ) | ( wire5506 ) | ( wire5507 ) ;
 assign wire5518 = ( wire843 ) | ( wire845 ) | ( wire858 ) ;
 assign wire5520 = ( wire5508 ) | ( wire5509 ) | ( wire5515 ) ;
 assign wire5521 = ( wire5462 ) | ( wire5463 ) | ( wire5467 ) | ( wire5517 ) ;
 assign wire5523 = ( wire5513 ) | ( wire5514 ) | ( wire5520 ) ;
 assign wire5526 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire5529 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire5532 = ( c  &  (~ d)  &  e  &  (~ n) ) ;
 assign wire5534 = ( g  &  i  &  j ) ;
 assign wire5557 = ( n_n1161  &  n_n713 ) | ( wire396  &  n_n875 ) ;
 assign wire5561 = ( n_n1220  &  n_n1171  &  wire206 ) | ( n_n1220  &  n_n698  &  wire206 ) ;
 assign wire5570 = ( n_n820  &  n_n1191  &  wire109 ) | ( n_n1191  &  wire23  &  wire109 ) ;
 assign wire5572 = ( wire809 ) | ( wire810 ) | ( wire811 ) | ( wire813 ) ;
 assign wire5573 = ( wire814 ) | ( wire817 ) | ( wire5561 ) ;
 assign wire5574 = ( wire821 ) | ( wire822 ) | ( wire826 ) | ( wire827 ) ;
 assign wire5575 = ( wire828 ) | ( wire829 ) | ( wire830 ) | ( wire831 ) ;
 assign wire5576 = ( wire823 ) | ( wire832 ) | ( wire835 ) ;
 assign wire5578 = ( wire808 ) | ( wire812 ) | ( wire815 ) | ( wire837 ) ;
 assign wire5579 = ( wire816 ) | ( wire818 ) | ( wire5570 ) ;
 assign wire5583 = ( wire836 ) | ( wire5578 ) | ( wire93  &  wire135 ) ;
 assign wire5584 = ( wire833 ) | ( wire834 ) | ( wire5572 ) | ( wire5579 ) ;
 assign wire5585 = ( wire5573 ) | ( wire5574 ) | ( wire5575 ) | ( wire5576 ) ;
 assign wire5587 = ( c  &  (~ d)  &  e ) ;
 assign wire5590 = ( i  &  j  &  (~ k) ) ;
 assign wire5592 = ( i  &  j  &  (~ k) ) ;
 assign wire5598 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5600 = ( i  &  j  &  (~ k) ) ;
 assign wire5601 = ( i  &  j  &  (~ k) ) ;
 assign wire5602 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5603 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5605 = ( (~ i)  &  wire148 ) | ( (~ j)  &  wire148 ) ;
 assign wire5611 = ( wire106  &  wire5602 ) | ( wire148  &  n_n893  &  wire106 ) ;
 assign wire5613 = ( wire148  &  wire156 ) | ( wire33  &  wire203 ) ;
 assign wire5615 = ( wire784 ) | ( wire786 ) | ( wire787 ) | ( wire788 ) ;
 assign wire5618 = ( wire50  &  wire5603 ) | ( wire5313  &  wire5603 ) | ( wire50  &  wire5605 ) | ( wire5313  &  wire5605 ) ;
 assign wire5619 = ( wire783 ) | ( wire785 ) | ( wire798 ) | ( wire799 ) ;
 assign wire5620 = ( wire789 ) | ( wire791 ) | ( wire5611 ) | ( wire5615 ) ;
 assign wire5621 = ( wire790 ) | ( wire796 ) | ( wire797 ) | ( wire5613 ) ;
 assign wire5624 = ( wire802 ) | ( wire5618 ) | ( wire5621 ) ;
 assign wire5629 = ( d  &  f  &  (~ j) ) ;
 assign wire5633 = ( n_n997  &  n_n1222  &  (~ n_n1260)  &  n_n992 ) ;
 assign wire5637 = ( d  &  (~ e)  &  f ) ;
 assign wire5639 = ( m  &  (~ n)  &  n_n997  &  wire5637 ) ;
 assign wire5640 = ( i  &  j  &  (~ k) ) ;
 assign wire5649 = ( n_n2494 ) | ( n_n1215  &  wire5629  &  wire5633 ) ;
 assign wire5650 = ( wire767 ) | ( wire781 ) | ( wire782 ) ;
 assign wire5652 = ( n_n2507 ) | ( wire766 ) | ( wire775 ) | ( wire776 ) ;
 assign wire5654 = ( wire116 ) | ( n_n2602 ) | ( wire777 ) | ( wire5652 ) ;
 assign wire5659 = ( m  &  (~ n)  &  n_n1261  &  n_n1146 ) ;
 assign wire5663 = ( (~ c)  &  (~ d)  &  (~ e)  &  (~ i) ) ;
 assign wire5664 = ( (~ k)  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire5666 = ( n_n2511 ) | ( n_n2602 ) ;
 assign wire5668 = ( wire754 ) | ( wire781 ) | ( wire782 ) ;
 assign wire5672 = ( wire319 ) | ( wire157 ) | ( wire267 ) | ( wire5666 ) ;
 assign wire5674 = ( c  &  d  &  (~ f)  &  g ) ;
 assign wire5677 = ( c  &  d  &  wire120  &  n_n1231 ) ;
 assign wire5678 = ( c  &  d  &  (~ f) ) ;
 assign wire5679 = ( m  &  (~ n)  &  n_n1261  &  wire5678 ) ;
 assign wire5681 = ( c  &  d  &  wire120  &  n_n912 ) ;
 assign wire5685 = ( n_n2602 ) | ( wire749 ) | ( wire181  &  wire5677 ) ;
 assign wire5686 = ( wire745 ) | ( wire46  &  wire5679 ) ;
 assign wire5687 = ( wire750 ) | ( wire46  &  wire5681 ) ;
 assign wire5690 = ( c  &  d  &  wire120 ) ;
 assign wire5693 = ( n_n1220  &  wire120  &  (~ wire57)  &  n_n1082 ) ;
 assign wire5694 = ( wire54  &  n_n971 ) | ( wire31  &  wire385 ) ;
 assign wire5695 = ( c  &  d  &  wire120 ) ;
 assign wire5696 = ( wire69  &  wire5695 ) | ( wire31  &  wire368  &  wire5695 ) ;
 assign wire5699 = ( a  &  b  &  c  &  d ) ;
 assign wire5703 = ( (~ a)  &  b  &  c  &  e ) ;
 assign wire5704 = ( a  &  c  &  (~ d)  &  e ) ;
 assign wire5705 = ( (~ a)  &  b  &  c  &  (~ d) ) ;
 assign wire5708 = ( n_n2660 ) | ( wire736 ) | ( wire108  &  wire5705 ) ;
 assign wire5709 = ( wire718 ) | ( wire719 ) | ( wire724 ) | ( wire726 ) ;
 assign wire5710 = ( wire200  &  wire5693 ) | ( wire379  &  wire5703 ) ;
 assign wire5711 = ( wire138  &  n_n949 ) | ( wire138  &  wire5704 ) ;
 assign wire5715 = ( n_n997  &  wire1112 ) | ( wire413  &  wire1112 ) | ( n_n997  &  wire1113 ) | ( wire413  &  wire1113 ) ;
 assign wire5718 = ( wire5708 ) | ( wire5711 ) | ( n_n949  &  wire94 ) ;
 assign wire5719 = ( wire725 ) | ( wire739  &  wire5696 ) | ( wire5694  &  wire5696 ) ;
 assign wire5720 = ( wire713 ) | ( wire727 ) | ( wire5709 ) ;
 assign wire5721 = ( wire716 ) | ( wire717 ) | ( wire5715 ) ;
 assign wire5722 = ( wire729 ) | ( wire731 ) | ( wire732 ) | ( wire5710 ) ;
 assign wire5726 = ( wire5718 ) | ( wire5719 ) | ( wire5720 ) | ( wire5721 ) ;
 assign wire5727 = ( m  &  (~ n)  &  n_n918  &  wire259 ) ;
 assign wire5731 = ( wire223  &  wire149 ) | ( wire149  &  wire388 ) ;
 assign wire5732 = ( wire708 ) | ( wire709 ) | ( wire46  &  wire5727 ) ;
 assign wire5740 = ( wire701 ) | ( wire702 ) | ( wire704 ) ;
 assign wire5743 = ( wire699 ) | ( wire55  &  wire388 ) | ( wire18  &  wire388 ) ;
 assign wire5744 = ( (~ e)  &  g  &  h  &  n_n988 ) ;
 assign wire5751 = ( b  &  d  &  e ) ;
 assign wire5752 = ( e  &  (~ g)  &  (~ h) ) ;
 assign wire5753 = ( b  &  d  &  e ) ;
 assign wire5758 = ( n_n840  &  wire76  &  n_n1095 ) | ( wire76  &  n_n988  &  n_n1095 ) ;
 assign wire5759 = ( wire228  &  wire159 ) | ( wire22  &  wire159  &  wire197 ) ;
 assign wire5760 = ( n_n2572 ) | ( wire680 ) | ( wire84  &  wire167 ) ;
 assign wire5761 = ( wire681 ) | ( wire682 ) | ( wire683 ) | ( wire684 ) ;
 assign wire5762 = ( n  &  wire160  &  wire49 ) | ( n  &  wire49  &  wire5744 ) ;
 assign wire5763 = ( n_n2660 ) | ( wire679 ) | ( wire736 ) | ( wire5758 ) ;
 assign wire5766 = ( wire5759 ) | ( wire5760 ) | ( wire5763 ) ;
 assign wire5774 = ( wire670 ) | ( wire671 ) | ( wire672 ) ;
 assign wire5775 = ( n_n2507 ) | ( n_n2494 ) | ( wire775 ) | ( wire776 ) ;
 assign wire5781 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire5792 = ( wire265  &  wire159 ) | ( wire75  &  wire167 ) ;
 assign wire5793 = ( wire643 ) | ( wire645 ) | ( wire77  &  wire160 ) ;
 assign wire5795 = ( wire649 ) | ( n_n838  &  (~ n_n1252)  &  wire117 ) ;
 assign wire5797 = ( n_n988  &  wire117 ) | ( n_n842  &  wire135 ) ;
 assign wire5798 = ( wire644 ) | ( wire647 ) | ( wire651 ) | ( wire652 ) ;
 assign wire5802 = ( wire646 ) | ( wire650 ) | ( wire653 ) | ( wire664 ) ;
 assign wire5803 = ( wire661 ) | ( wire5795 ) | ( wire200  &  n_n872 ) ;
 assign wire5804 = ( wire5798 ) | ( wire5797 ) ;
 assign wire5806 = ( wire655 ) | ( wire657 ) | ( wire658 ) | ( wire663 ) ;
 assign wire5809 = ( n_n1919 ) | ( wire5761 ) | ( wire5762 ) | ( wire5766 ) ;
 assign wire5810 = ( n_n1939 ) | ( wire5792 ) | ( wire5793 ) | ( wire5806 ) ;
 assign wire5811 = ( n_n1920 ) | ( wire5802 ) | ( wire5803 ) | ( wire5804 ) ;
 assign wire5813 = ( f  &  h  &  i ) ;
 assign wire5814 = ( n_n709  &  wire70  &  n_n992 ) | ( n_n1171  &  wire70  &  n_n992 ) ;
 assign wire5824 = ( wire626 ) | ( wire629 ) | ( wire630 ) | ( wire633 ) ;
 assign wire5825 = ( wire627 ) | ( n_n698  &  wire72 ) ;
 assign wire5826 = ( wire628 ) | ( wire631 ) | ( wire632 ) | ( wire635 ) ;
 assign wire5828 = ( wire5825 ) | ( n_n1210  &  wire211 ) ;
 assign wire5829 = ( wire320 ) | ( wire5824 ) | ( wire5826 ) ;
 assign wire5830 = ( (~ k)  &  (~ l)  &  m  &  (~ n) ) ;
 assign wire5831 = ( wire54  &  n_n1155 ) | ( n_n529  &  wire142 ) ;
 assign wire5833 = ( (~ n_n1193)  &  (~ n_n1201)  &  n_n918  &  n_n1187 ) ;
 assign wire5834 = ( k  &  m  &  (~ n)  &  n_n1207 ) ;
 assign wire5835 = ( m  &  (~ n)  &  n_n1207  &  wire29 ) ;
 assign wire5836 = ( m  &  (~ n)  &  n_n1201  &  wire29 ) ;
 assign wire5837 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5839 = ( i  &  k  &  m  &  (~ n) ) ;
 assign wire5840 = ( n_n2953 ) | ( wire22  &  wire15  &  n_n766 ) ;
 assign wire5841 = ( wire617 ) | ( wire15  &  n_n1228  &  wire5834 ) ;
 assign wire5842 = ( wire610 ) | ( wire156  &  wire5837 ) ;
 assign wire5843 = ( wire619 ) | ( wire15  &  wire113  &  n_n1228 ) ;
 assign wire5846 = ( wire81  &  wire5833 ) | ( wire5831  &  wire5833 ) | ( wire81  &  wire5835 ) | ( wire5831  &  wire5835 ) ;
 assign wire5847 = ( n_n698  &  wire81 ) | ( n_n698  &  wire5831 ) | ( wire81  &  wire5836 ) | ( wire5831  &  wire5836 ) ;
 assign wire5848 = ( wire5840 ) | ( wire5841 ) | ( wire5842 ) | ( wire5843 ) ;
 assign wire5849 = ( wire611 ) | ( wire220  &  wire81 ) | ( wire220  &  wire5831 ) ;
 assign wire5850 = ( wire618 ) | ( wire82  &  wire81 ) | ( wire82  &  wire5831 ) ;
 assign wire5851 = ( wire5847 ) | ( wire5846 ) ;
 assign wire5857 = ( a  &  b  &  d  &  (~ e) ) ;
 assign wire5858 = ( h  &  i  &  j  &  n_n1202 ) ;
 assign wire5860 = ( n_n1155  &  n_n700  &  n_n1191 ) | ( n_n700  &  n_n820  &  n_n1191 ) ;
 assign wire5864 = ( wire594 ) | ( wire203  &  wire113 ) ;
 assign wire5865 = ( wire587 ) | ( wire588 ) | ( wire5860 ) ;
 assign wire5866 = ( wire593 ) | ( wire598 ) | ( n_n1210  &  wire208 ) ;
 assign wire5867 = ( n_n3060 ) | ( wire585 ) | ( wire586 ) | ( wire590 ) ;
 assign wire5870 = ( wire5864 ) | ( wire5865 ) | ( wire5867 ) ;
 assign wire5871 = ( wire40  &  wire1039 ) | ( wire40  &  wire5270 ) | ( wire1039  &  wire5858 ) | ( wire5270  &  wire5858 ) ;
 assign wire5873 = ( wire351 ) | ( wire5866 ) | ( wire5870 ) | ( wire5871 ) ;
 assign wire5875 = ( h  &  i  &  (~ j)  &  k ) ;
 assign wire5876 = ( wire5875  &  (~ wire104) ) ;
 assign wire5877 = ( n_n711  &  wire293 ) | ( wire30  &  wire293 ) ;
 assign wire5884 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire5886 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire5888 = ( (~ h)  &  (~ k) ) | ( j  &  (~ k) ) ;
 assign wire5897 = ( n_n2953 ) | ( wire567 ) | ( wire575 ) ;
 assign wire5898 = ( wire568 ) | ( wire576 ) | ( wire5876  &  wire5877 ) ;
 assign wire5899 = ( wire571 ) | ( wire219  &  wire5888 ) | ( wire1016  &  wire5888 ) ;
 assign wire5901 = ( wire565 ) | ( wire566 ) | ( wire569 ) | ( wire577 ) ;
 assign wire5903 = ( wire5898 ) | ( wire315  &  wire81 ) | ( wire315  &  wire583 ) ;
 assign wire5904 = ( wire579 ) | ( wire581 ) | ( wire5899 ) ;
 assign wire5905 = ( wire570 ) | ( wire573 ) | ( wire5897 ) | ( wire5901 ) ;
 assign wire5906 = ( wire580 ) | ( wire572 ) ;
 assign wire5912 = ( n_n840  &  wire230  &  n_n1210 ) ;
 assign wire5925 = ( wire540 ) | ( n_n711  &  wire5912 ) | ( wire30  &  wire5912 ) ;
 assign wire5927 = ( wire536 ) | ( wire539 ) | ( wire541 ) | ( wire542 ) ;
 assign wire5928 = ( wire543 ) | ( wire544 ) | ( wire545 ) | ( wire549 ) ;
 assign wire5929 = ( wire550 ) | ( wire551 ) | ( n_n1264  &  wire209 ) ;
 assign wire5930 = ( wire537 ) | ( wire554 ) | ( n_n1220  &  wire50 ) ;
 assign wire5934 = ( wire548 ) | ( n_n1210  &  wire169 ) | ( n_n1210  &  wire980 ) ;
 assign wire5936 = ( wire546 ) | ( wire552 ) | ( wire5925 ) | ( wire5930 ) ;
 assign wire5937 = ( wire320 ) | ( wire547 ) | ( wire5927 ) | ( wire5928 ) ;
 assign wire5938 = ( wire5929 ) | ( wire5934 ) | ( n_n1220  &  wire207 ) ;
 assign wire5941 = ( (~ g)  &  (~ h)  &  (~ k) ) ;
 assign wire5943 = ( e  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire5944 = ( (~ c)  &  d  &  (~ g)  &  (~ h) ) ;
 assign wire5945 = ( c  &  (~ f)  &  (~ h)  &  i ) ;
 assign wire5946 = ( (~ d)  &  g  &  (~ h)  &  i ) ;
 assign wire5951 = ( wire282  &  wire5944 ) | ( wire282  &  wire5945 ) ;
 assign wire5954 = ( wire528 ) | ( wire5951 ) | ( wire373  &  wire5943 ) ;
 assign wire5955 = ( wire532 ) | ( wire533 ) | ( wire534 ) | ( wire535 ) ;
 assign wire5958 = ( d  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire5959 = ( a  &  g  &  h ) | ( (~ b)  &  g  &  h ) ;
 assign wire5961 = ( b  &  (~ f)  &  (~ h)  &  i ) ;
 assign wire5962 = ( (~ b)  &  (~ e)  &  g  &  (~ h) ) ;
 assign wire5963 = ( b  &  e  &  (~ f)  &  (~ h) ) ;
 assign wire5964 = ( (~ e)  &  (~ f)  &  (~ l) ) ;
 assign wire5967 = ( wire227  &  wire5961 ) | ( wire227  &  wire5962 ) ;
 assign wire5969 = ( wire520 ) | ( wire521 ) | ( wire522 ) | ( wire523 ) ;
 assign wire5970 = ( wire527 ) | ( wire5967 ) | ( wire227  &  wire5963 ) ;
 assign wire5971 = ( (~ h)  &  i ) | ( (~ h)  &  (~ j) ) ;
 assign wire5977 = ( (~ a)  &  (~ e)  &  (~ f)  &  (~ g) ) ;
 assign wire5979 = ( e  &  (~ f)  &  h  &  j ) ;
 assign wire5981 = ( (~ i)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire5982 = ( f  &  k  &  m  &  (~ n) ) ;
 assign wire5986 = ( wire22  &  wire283 ) | ( n_n1171  &  wire286 ) ;
 assign wire5990 = ( n_n1187  &  n_n1189  &  wire5981 ) | ( n_n1187  &  n_n1189  &  wire5982 ) ;
 assign wire5996 = ( wire500 ) | ( wire501 ) | ( wire503 ) | ( wire517 ) ;
 assign wire5998 = ( wire508 ) | ( wire509 ) | ( wire510 ) | ( wire512 ) ;
 assign wire5999 = ( wire499 ) | ( wire513 ) | ( wire516 ) | ( wire5986 ) ;
 assign wire6001 = ( wire504 ) | ( wire505 ) | ( wire5990 ) | ( wire5998 ) ;
 assign wire6002 = ( wire502 ) | ( wire511 ) | ( wire5996 ) | ( wire5999 ) ;
 assign wire6005 = ( (~ c)  &  e  &  (~ f) ) | ( c  &  (~ e)  &  (~ f) ) ;
 assign wire6006 = ( c  &  (~ g)  &  h ) ;
 assign wire6010 = ( c  &  i ) | ( d  &  i ) | ( e  &  i ) ;
 assign wire6012 = ( c  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire6014 = ( (~ f)  &  k  &  (~ m)  &  (~ n) ) ;
 assign wire6020 = ( (~ e)  &  (~ f)  &  (~ g)  &  (~ i) ) ;
 assign wire6022 = ( (~ h)  &  (~ k)  &  m  &  (~ n) ) ;
 assign wire6035 = ( wire481 ) | ( wire483 ) | ( wire487 ) ;
 assign wire6036 = ( wire484 ) | ( wire488 ) | ( wire489 ) | ( wire490 ) ;
 assign wire6037 = ( wire491 ) | ( wire492 ) | ( wire493 ) | ( wire494 ) ;
 assign wire6038 = ( wire480 ) | ( wire482 ) | ( wire495 ) | ( wire496 ) ;
 assign wire6040 = ( wire6037 ) | ( wire6036 ) ;
 assign wire6041 = ( wire485 ) | ( wire486 ) | ( wire6035 ) | ( wire6038 ) ;
 assign wire6042 = ( (~ d)  &  (~ f)  &  g  &  (~ h) ) ;
 assign wire6045 = ( f  &  (~ i)  &  k  &  (~ m) ) ;
 assign wire6047 = ( (~ h)  &  i  &  (~ m)  &  (~ n) ) ;
 assign wire6054 = ( c  &  (~ f)  &  (~ h) ) | ( (~ c)  &  g  &  (~ h) ) ;
 assign wire6057 = ( n_n1095  &  n_n1227 ) | ( n_n1203  &  wire226 ) ;
 assign wire6062 = ( n_n1160  &  wire70 ) | ( n_n1161  &  wire285 ) ;
 assign wire6064 = ( wire464 ) | ( wire226  &  (~ wire395)  &  wire6045 ) ;
 assign wire6065 = ( wire463 ) | ( wire465 ) | ( wire466 ) | ( wire467 ) ;
 assign wire6066 = ( wire468 ) | ( wire469 ) | ( wire470 ) | ( wire471 ) ;
 assign wire6067 = ( wire461 ) | ( wire6057 ) | ( wire6062 ) ;
 assign wire6070 = ( wire6064 ) | ( wire6065 ) | ( wire6066 ) | ( wire6067 ) ;
 assign wire6071 = ( wire6001 ) | ( wire6002 ) | ( wire6040 ) | ( wire6041 ) ;
 assign wire6072 = ( c  &  (~ i)  &  (~ k) ) ;
 assign wire6074 = ( (~ l)  &  (~ e) ) ;
 assign wire6076 = ( (~ e)  &  (~ d) ) ;
 assign wire6078 = ( (~ d)  &  h ) | ( (~ e)  &  h ) | ( (~ f)  &  h ) ;
 assign wire6082 = ( (~ e)  &  (~ f)  &  i ) | ( (~ e)  &  (~ f)  &  (~ j) ) ;
 assign wire6085 = ( a  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire6100 = ( wire443 ) | ( wire444 ) | ( wire445 ) | ( wire447 ) ;
 assign wire6101 = ( wire448 ) | ( wire449 ) | ( wire450 ) | ( wire451 ) ;
 assign wire6102 = ( wire452 ) | ( wire453 ) | ( wire454 ) | ( wire455 ) ;
 assign wire6103 = ( wire456 ) | ( wire457 ) | ( wire458 ) | ( wire460 ) ;
 assign wire6106 = ( wire446 ) | ( wire459 ) | ( wire6100 ) | ( wire6103 ) ;
 assign wire6107 = ( (~ e)  &  (~ d) ) ;
 assign wire6108 = ( m  &  (~ n)  &  n_n1261  &  wire6107 ) ;
 assign wire6109 = ( f  &  g  &  h ) ;
 assign wire6112 = ( (~ a)  &  f  &  g  &  h ) ;
 assign wire6115 = ( h  &  j ) | ( i  &  j ) ;
 assign wire6118 = ( (~ e)  &  (~ f)  &  (~ h)  &  (~ j) ) ;
 assign wire6119 = ( c  &  d  &  e  &  (~ n) ) ;
 assign wire6122 = ( m  &  (~ n)  &  n_n1261  &  n_n1260 ) ;
 assign wire6123 = ( (~ b)  &  g  &  h ) ;
 assign wire6125 = ( m ) | ( (~ i)  &  k ) | ( (~ i)  &  l ) | ( (~ k)  &  l ) ;
 assign wire6130 = ( wire440 ) | ( n_n1217  &  n_n1215  &  wire6123 ) ;
 assign wire6131 = ( wire441 ) | ( (~ g)  &  wire85  &  wire6108 ) ;
 assign wire6132 = ( wire435 ) | ( (~ n_n1217)  &  wire6122 ) | ( (~ n_n1215)  &  wire6122 ) ;
 assign wire6133 = ( wire248  &  wire6125 ) | ( wire37  &  (~ n_n1216)  &  wire248 ) ;
 assign wire6135 = ( wire431 ) | ( wire432 ) | ( wire433 ) | ( wire434 ) ;
 assign wire6138 = ( wire429 ) | ( wire430 ) | ( wire442 ) | ( wire6135 ) ;
 assign wire6139 = ( wire6130 ) | ( wire6131 ) | ( wire6132 ) | ( wire6133 ) ;
 assign wire6141 = ( (~ h)  &  i  &  (~ k) ) | ( (~ h)  &  (~ j)  &  (~ k) ) ;
 assign wire6142 = ( (~ h)  &  i  &  (~ k) ) ;
 assign wire6143 = ( (~ h)  &  i  &  (~ k) ) ;
 assign wire6144 = ( (~ i)  &  (~ m)  &  n ) ;
 assign wire6145 = ( n_n1190  &  wire6143 ) | ( n_n1160  &  wire6144 ) ;
 assign wire6147 = ( n_n1056  &  wire6141 ) | ( n_n1219  &  wire6142 ) ;
 assign wire6149 = ( wire6145 ) | ( n_n1089  &  wire127 ) | ( wire127  &  n_n1160 ) ;
 assign wire6150 = ( wire424 ) | ( wire425 ) | ( wire6147 ) ;
 assign wire6151 = ( (~ g)  &  (~ m)  &  (~ n) ) ;
 assign wire6156 = ( c  &  (~ m)  &  n ) | ( d  &  (~ m)  &  n ) ;
 assign wire6158 = ( g  &  (~ m)  &  n ) ;
 assign wire6159 = ( n_n1091  &  wire6156 ) | ( n_n1080  &  wire6158 ) ;
 assign wire6160 = ( wire114  &  wire404 ) | ( n_n1190  &  wire305 ) ;
 assign wire6161 = ( n_n1080  &  (~ wire204) ) | ( wire286  &  wire137 ) ;
 assign wire6165 = ( k  &  n_n1177  &  n_n1028 ) | ( n_n1177  &  n_n1072  &  n_n1028 ) ;
 assign wire6168 = ( wire353 ) | ( n_n1072  &  wire161 ) ;
 assign wire6169 = ( wire352 ) | ( wire354 ) | ( wire355 ) | ( wire389 ) ;
 assign wire6170 = ( wire357 ) | ( wire359 ) | ( wire6165 ) ;
 assign wire6171 = ( wire362 ) | ( wire6159 ) | ( wire6160 ) | ( wire6161 ) ;
 assign wire6176 = ( (~ n_n671)  &  (~ n_n700)  &  (~ n_n1260) ) ;
 assign wire6177 = ( (~ f)  &  (~ g)  &  (~ m)  &  n ) ;
 assign wire6180 = ( f ) | ( (~ b)  &  e ) ;
 assign wire6183 = ( (~ b)  &  (~ m)  &  n  &  wire286 ) ;
 assign wire6184 = ( m  &  (~ n_n1249) ) | ( (~ n)  &  (~ n_n1249) ) | ( (~ n_n1121)  &  (~ n_n1249) ) ;
 assign wire6185 = ( (~ b)  &  (~ f)  &  (~ m)  &  n ) ;
 assign wire6187 = ( (~ c)  &  (~ e)  &  (~ f) ) | ( d  &  (~ e)  &  (~ f) ) ;
 assign wire6188 = ( (~ a)  &  (~ f)  &  m  &  (~ n) ) ;
 assign wire6194 = ( wire407  &  n_n1191 ) | ( wire226  &  wire249 ) ;
 assign wire6195 = ( wire120  &  n_n1039 ) | ( wire120  &  n_n1072 ) ;
 assign wire6200 = ( k  &  n_n1177  &  n_n1028 ) | ( n_n1177  &  n_n1028  &  wire273 ) ;
 assign wire6203 = ( wire334 ) | ( wire404  &  (~ n_n1121)  &  wire6176 ) ;
 assign wire6204 = ( wire333 ) | ( wire336 ) | ( wire6183  &  wire6184 ) ;
 assign wire6205 = ( wire337 ) | ( wire338 ) | ( wire339 ) | ( wire340 ) ;
 assign wire6206 = ( wire341 ) | ( wire342 ) | ( wire6200 ) ;
 assign wire6207 = ( wire345 ) | ( wire347 ) | ( wire6194 ) | ( wire6195 ) ;
 assign wire6210 = ( wire6203 ) | ( wire6204 ) | ( wire6207 ) ;
 assign wire6211 = ( i  &  (~ m)  &  (~ n) ) ;
 assign wire6213 = ( c  &  d ) | ( (~ c)  &  f ) | ( d  &  f ) | ( c  &  (~ f) ) | ( (~ c)  &  g ) | ( d  &  g ) | ( (~ f)  &  g ) ;
 assign wire6216 = ( (~ n_n857)  &  (~ n_n1260)  &  (~ wire35) ) ;
 assign wire6217 = ( (~ n_n766)  &  (~ n_n919)  &  wire6213 ) ;
 assign wire6220 = ( (~ c)  &  (~ f)  &  i ) | ( (~ c)  &  g  &  i ) ;
 assign wire6222 = ( (~ j)  &  k  &  (~ m)  &  (~ n) ) ;
 assign wire6224 = ( (~ n_n857)  &  (~ n_n1260)  &  wire6222 ) ;
 assign wire6225 = ( i  &  j  &  (~ m)  &  (~ n) ) ;
 assign wire6226 = ( c ) | ( (~ d) ) ;
 assign wire6227 = ( c  &  (~ f) ) | ( (~ f)  &  g ) | ( c  &  (~ g) ) | ( f  &  (~ g) ) | ( c  &  (~ j) ) | ( f  &  (~ j) ) | ( g  &  (~ j) ) ;
 assign wire6230 = ( (~ f)  &  (~ c) ) ;
 assign wire6233 = ( (~ a)  &  m  &  (~ n) ) ;
 assign wire6236 = ( (~ d)  &  j ) | ( e  &  j ) | ( (~ g)  &  j ) ;
 assign wire6238 = ( (~ c)  &  (~ d)  &  (~ e)  &  f ) ;
 assign wire6239 = ( (~ a)  &  (~ e)  &  (~ f) ) ;
 assign wire6240 = ( i  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire6241 = ( g  &  (~ l)  &  (~ m)  &  (~ n) ) ;
 assign wire6245 = ( wire170  &  wire6238 ) | ( n_n857  &  wire170  &  wire305 ) ;
 assign wire6246 = ( n_n1091  &  wire6240 ) | ( n_n1167  &  wire6241 ) ;
 assign wire6248 = ( wire331 ) | ( (~ n_n919)  &  wire6220  &  wire6224 ) ;
 assign wire6249 = ( wire316 ) | ( wire161  &  wire6239 ) ;
 assign wire6250 = ( wire317 ) | ( wire318 ) | ( wire329 ) ;
 assign wire6251 = ( wire321 ) | ( wire322 ) | ( wire6245 ) ;
 assign wire6252 = ( wire328 ) | ( wire330 ) | ( wire6246 ) ;
 assign wire6256 = ( wire307 ) | ( wire6248 ) | ( wire6249 ) | ( wire6250 ) ;
 assign wire6257 = ( g ) | ( (~ f)  &  h ) ;
 assign wire6258 = ( (~ i)  &  (~ k)  &  (~ m)  &  (~ n) ) ;
 assign wire6262 = ( h  &  (~ j)  &  (~ k)  &  (~ m) ) ;
 assign wire6263 = ( (~ g)  &  (~ h) ) | ( (~ g)  &  i ) | ( g  &  (~ i) ) | ( (~ h)  &  (~ i) ) | ( g  &  j ) | ( (~ h)  &  j ) | ( i  &  j ) ;
 assign wire6264 = ( (~ g)  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire6266 = ( (~ c)  &  (~ d)  &  g ) ;
 assign wire6268 = ( c  &  (~ g)  &  (~ h) ) | ( f  &  (~ g)  &  (~ h) ) ;
 assign wire6272 = ( h  &  (~ i)  &  (~ m)  &  (~ n) ) ;
 assign wire6281 = ( wire253 ) | ( wire271 ) | ( wire272 ) | ( wire274 ) ;
 assign wire6282 = ( wire275 ) | ( wire276 ) | ( wire277 ) | ( wire278 ) ;
 assign wire6283 = ( wire252 ) | ( wire269 ) | ( wire280 ) | ( wire281 ) ;
 assign wire6285 = ( wire6281 ) | ( wire6282 ) | ( wire6283 ) ;
 assign wire6286 = ( wire6205 ) | ( wire6206 ) | ( wire6210 ) | ( wire6285 ) ;
 assign wire6287 = ( c  &  h  &  (~ j) ) | ( d  &  h  &  (~ j) ) ;
 assign wire6289 = ( (~ c)  &  g  &  h ) | ( (~ d)  &  g  &  h ) ;
 assign wire6290 = ( (~ c)  &  h  &  (~ j) ) | ( (~ d)  &  h  &  (~ j) ) ;
 assign wire6292 = ( wire178 ) | ( n_n1036  &  wire6290 ) ;
 assign wire6293 = ( wire177 ) | ( wire173 ) ;
 assign wire6297 = ( wire140 ) | ( wire6293 ) | ( n_n1022  &  n_n1036 ) ;
 assign wire6298 = ( wire150 ) | ( wire163 ) | ( wire180 ) | ( wire6292 ) ;
 assign wire6300 = ( wire5954 ) | ( wire5955 ) | ( wire5969 ) | ( wire5970 ) ;
 assign wire6301 = ( wire6149 ) | ( wire6150 ) | ( wire6297 ) | ( wire6298 ) ;
 assign wire6303 = ( wire6101 ) | ( wire6102 ) | ( wire6106 ) | ( wire6301 ) ;
 assign wire6304 = ( n_n2023 ) | ( wire6138 ) | ( wire6139 ) | ( wire6300 ) ;
 assign wire6306 = ( n_n2026 ) | ( wire6070 ) | ( wire6071 ) | ( wire6286 ) ;
 assign wire6307 = ( g  &  (~ h)  &  (~ i) ) ;
 assign wire6309 = ( m  &  (~ n)  &  n_n997  &  wire6307 ) ;
 assign wire6310 = ( (~ i)  &  (~ j)  &  (~ k) ) ;
 assign wire6317 = ( wire63 ) | ( n_n996  &  n_n1072  &  wire6309 ) ;
 assign wire6318 = ( wire42 ) | ( wire61 ) | ( wire66 ) ;
 assign wire6322 = ( wire116 ) | ( wire781 ) | ( wire782 ) | ( wire6318 ) ;
 assign wire6323 = ( wire199 ) | ( wire157 ) | ( wire267 ) | ( wire6317 ) ;


endmodule

