module pdc (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, 
	i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, 
	o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, 
	o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, 
	o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, 
	o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_9_;
input i_10_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_14_;
input i_3_;
input i_13_;
input i_4_;
input i_12_;
input i_1_;
input i_11_;
input i_2_;
input i_0_;
input i_15_;
output o_1_;
output o_19_;
output o_2_;
output o_0_;
output o_29_;
output o_39_;
output o_38_;
output o_25_;
output o_12_;
output o_37_;
output o_26_;
output o_11_;
output o_36_;
output o_27_;
output o_14_;
output o_35_;
output o_28_;
output o_13_;
output o_34_;
output o_21_;
output o_16_;
output o_33_;
output o_22_;
output o_15_;
output o_32_;
output o_23_;
output o_18_;
output o_31_;
output o_24_;
output o_17_;
output o_30_;
output o_20_;
output o_10_;
output o_9_;
output o_7_;
output o_8_;
output o_5_;
output o_6_;
output o_3_;
output o_4_;
wire n_n139;
wire n_n151;
wire n_n5686;
wire n_n5231;
wire n_n310;
wire n_n4476;
wire n_n4477;
wire wire394;
wire wire507;
wire wire893;
wire wire937;
wire n_n863;
wire n_n3625;
wire n_n3626;
wire n_n3627;
wire n_n3621;
wire n_n3631;
wire n_n3661;
wire n_n3632;
wire n_n124;
wire n_n123;
wire wire289;
wire wire364;
wire wire535;
wire wire777;
wire wire834;
wire wire939;
wire wire938;
wire n_n106;
wire n_n5678;
wire n_n5671;
wire wire396;
wire wire582;
wire wire583;
wire wire941;
wire wire940;
wire n_n272;
wire n_n118;
wire n_n4442;
wire n_n4439;
wire wire943;
wire n_n231;
wire n_n5792;
wire n_n5794;
wire n_n4203;
wire n_n4206;
wire n_n4306;
wire n_n4807;
wire n_n4223;
wire n_n4224;
wire n_n4303;
wire n_n1;
wire n_n2;
wire n_n2618;
wire wire944;
wire n_n5769;
wire n_n127;
wire n_n4982;
wire wire48;
wire n_n265;
wire n_n268;
wire n_n2550;
wire n_n2545;
wire wire268;
wire wire782;
wire n_n5796;
wire n_n4808;
wire n_n4809;
wire n_n4719;
wire n_n4718;
wire n_n264;
wire n_n153;
wire n_n120;
wire n_n2772;
wire n_n130;
wire n_n110;
wire n_n121;
wire n_n4705;
wire n_n4704;
wire wire949;
wire wire948;
wire n_n5224;
wire n_n4534;
wire n_n4533;
wire n_n4532;
wire n_n4531;
wire n_n4530;
wire n_n3892;
wire n_n4141;
wire n_n4015;
wire n_n4;
wire n_n2789;
wire n_n2795;
wire n_n2840;
wire n_n2839;
wire n_n128;
wire n_n5682;
wire n_n5676;
wire n_n4512;
wire n_n4508;
wire wire216;
wire n_n255;
wire n_n4186;
wire wire392;
wire wire559;
wire wire950;
wire n_n5247;
wire wire926;
wire n_n5797;
wire wire503;
wire n_n4197;
wire n_n4194;
wire n_n5235;
wire n_n163;
wire n_n5693;
wire wire452;
wire wire758;
wire wire923;
wire n_n132;
wire n_n3140;
wire n_n7424;
wire n_n3;
wire n_n3727;
wire n_n3138;
wire n_n3089;
wire n_n3094;
wire n_n152;
wire n_n111;
wire n_n133;
wire n_n3898;
wire n_n3890;
wire n_n3897;
wire n_n3896;
wire n_n57;
wire n_n56;
wire n_n2440;
wire wire955;
wire n_n2060;
wire n_n145;
wire n_n2062;
wire n_n2058;
wire n_n2063;
wire n_n2064;
wire n_n2065;
wire wire169;
wire n_n126;
wire n_n5660;
wire n_n5659;
wire n_n1670;
wire wire581;
wire wire880;
wire n_n1729;
wire n_n1679;
wire n_n1694;
wire n_n1693;
wire wire957;
wire n_n1089;
wire n_n240;
wire n_n380;
wire n_n381;
wire n_n333;
wire n_n746;
wire n_n731;
wire n_n745;
wire wire126;
wire n_n189;
wire n_n5053;
wire n_n241;
wire n_n5061;
wire n_n5062;
wire n_n5020;
wire n_n99;
wire n_n54;
wire n_n186;
wire wire863;
wire n_n4970;
wire wire153;
wire wire200;
wire n_n4926;
wire n_n4315;
wire n_n6;
wire n_n5;
wire n_n4826;
wire n_n4828;
wire n_n4823;
wire wire90;
wire wire584;
wire wire976;
wire n_n4204;
wire n_n4815;
wire n_n4821;
wire n_n4814;
wire n_n4816;
wire wire573;
wire wire60;
wire n_n4834;
wire n_n4961;
wire n_n4966;
wire n_n4967;
wire wire613;
wire wire614;
wire n_n4251;
wire n_n4287;
wire wire99;
wire wire389;
wire wire708;
wire n_n4211;
wire wire166;
wire wire224;
wire wire617;
wire wire673;
wire wire674;
wire n_n4210;
wire n_n4892;
wire n_n4898;
wire n_n4895;
wire wire488;
wire wire878;
wire n_n48;
wire wire51;
wire n_n4179;
wire n_n53;
wire wire40;
wire n_n4168;
wire n_n197;
wire n_n37;
wire wire89;
wire n_n4094;
wire n_n105;
wire n_n47;
wire n_n108;
wire wire67;
wire n_n4174;
wire wire407;
wire wire457;
wire n_n4153;
wire n_n4154;
wire wire456;
wire n_n3964;
wire n_n896;
wire n_n95;
wire n_n76;
wire wire460;
wire wire160;
wire wire409;
wire n_n4920;
wire n_n4907;
wire wire44;
wire wire82;
wire wire635;
wire wire636;
wire n_n3129;
wire n_n11;
wire wire539;
wire wire639;
wire n_n3172;
wire n_n4605;
wire n_n3118;
wire wire640;
wire wire867;
wire n_n3107;
wire n_n3259;
wire n_n3260;
wire n_n3772;
wire n_n3257;
wire n_n3113;
wire n_n2860;
wire n_n3255;
wire wire814;
wire n_n3112;
wire n_n3162;
wire wire68;
wire wire496;
wire wire806;
wire n_n3096;
wire n_n31;
wire n_n10;
wire n_n100;
wire n_n1359;
wire n_n3525;
wire n_n107;
wire wire983;
wire n_n2136;
wire n_n4671;
wire wire252;
wire wire329;
wire n_n2169;
wire n_n12;
wire n_n66;
wire wire164;
wire n_n60;
wire wire985;
wire n_n2081;
wire wire333;
wire n_n2101;
wire wire988;
wire n_n147;
wire n_n94;
wire n_n280;
wire n_n32;
wire n_n80;
wire wire62;
wire n_n4165;
wire n_n42;
wire wire81;
wire n_n1506;
wire wire69;
wire n_n4624;
wire n_n1412;
wire wire990;
wire wire664;
wire wire992;
wire n_n4858;
wire n_n4864;
wire n_n4635;
wire n_n1129;
wire n_n6582;
wire n_n4870;
wire n_n1497;
wire n_n1130;
wire n_n4846;
wire n_n4852;
wire n_n1490;
wire wire998;
wire n_n1095;
wire n_n1132;
wire n_n1133;
wire n_n1505;
wire n_n1096;
wire n_n1542;
wire n_n3827;
wire n_n1135;
wire n_n1097;
wire n_n9;
wire n_n65;
wire wire368;
wire n_n1066;
wire wire114;
wire wire120;
wire wire459;
wire n_n855;
wire n_n3870;
wire wire881;
wire n_n772;
wire wire301;
wire wire461;
wire n_n824;
wire wire670;
wire n_n761;
wire n_n275;
wire n_n266;
wire wire916;
wire n_n260;
wire n_n269;
wire n_n253;
wire n_n229;
wire n_n227;
wire n_n254;
wire n_n274;
wire n_n242;
wire n_n208;
wire n_n207;
wire n_n279;
wire wire911;
wire n_n204;
wire n_n273;
wire n_n177;
wire wire901;
wire n_n84;
wire n_n222;
wire n_n283;
wire n_n247;
wire n_n155;
wire n_n165;
wire n_n142;
wire wire899;
wire n_n223;
wire n_n136;
wire n_n281;
wire wire913;
wire wire896;
wire n_n230;
wire n_n261;
wire n_n278;
wire n_n259;
wire n_n149;
wire n_n271;
wire n_n122;
wire n_n112;
wire wire900;
wire n_n93;
wire wire898;
wire n_n228;
wire wire903;
wire n_n212;
wire wire902;
wire n_n30;
wire n_n221;
wire n_n258;
wire n_n216;
wire n_n220;
wire wire912;
wire n_n7;
wire n_n144;
wire wire905;
wire n_n257;
wire n_n50;
wire n_n267;
wire wire906;
wire n_n46;
wire n_n256;
wire n_n89;
wire wire914;
wire n_n87;
wire n_n282;
wire n_n34;
wire n_n225;
wire n_n270;
wire n_n28;
wire wire897;
wire n_n75;
wire n_n171;
wire n_n21;
wire n_n17;
wire n_n246;
wire n_n236;
wire wire908;
wire n_n40;
wire wire904;
wire n_n102;
wire n_n263;
wire wire907;
wire n_n33;
wire n_n135;
wire n_n78;
wire n_n200;
wire n_n29;
wire n_n64;
wire n_n150;
wire n_n25;
wire n_n70;
wire n_n24;
wire n_n27;
wire n_n20;
wire n_n97;
wire n_n45;
wire n_n52;
wire n_n41;
wire n_n26;
wire n_n23;
wire n_n74;
wire n_n71;
wire n_n69;
wire n_n14;
wire n_n252;
wire n_n63;
wire n_n8;
wire n_n199;
wire n_n18;
wire n_n88;
wire n_n92;
wire n_n98;
wire n_n179;
wire n_n104;
wire n_n38;
wire n_n109;
wire wire1011;
wire n_n5030;
wire n_n5063;
wire wire927;
wire wire254;
wire wire165;
wire n_n4936;
wire n_n6678;
wire wire79;
wire n_n4839;
wire n_n4842;
wire wire1016;
wire n_n4960;
wire n_n4954;
wire n_n4953;
wire n_n4955;
wire wire671;
wire n_n4219;
wire n_n226;
wire n_n61;
wire wire469;
wire n_n4073;
wire wire475;
wire n_n4068;
wire n_n4069;
wire wire77;
wire n_n1363;
wire wire184;
wire n_n3324;
wire n_n6504;
wire n_n1633;
wire n_n4923;
wire wire385;
wire n_n3130;
wire wire686;
wire wire825;
wire n_n3167;
wire wire278;
wire wire1018;
wire n_n3117;
wire n_n3242;
wire wire557;
wire n_n3108;
wire n_n3757;
wire wire739;
wire n_n3110;
wire n_n2852;
wire n_n3109;
wire n_n3155;
wire n_n3519;
wire n_n3520;
wire wire1027;
wire wire1026;
wire n_n81;
wire wire470;
wire n_n3019;
wire n_n2986;
wire n_n3524;
wire wire93;
wire wire185;
wire n_n2148;
wire n_n19;
wire n_n2272;
wire n_n2126;
wire wire135;
wire wire264;
wire wire1031;
wire wire1030;
wire wire466;
wire n_n2104;
wire wire411;
wire n_n2137;
wire n_n2110;
wire n_n2073;
wire n_n2108;
wire wire476;
wire wire1042;
wire n_n1779;
wire n_n58;
wire wire667;
wire wire696;
wire n_n1757;
wire n_n3581;
wire wire700;
wire wire1043;
wire n_n1215;
wire n_n1628;
wire n_n2732;
wire n_n1624;
wire wire1044;
wire n_n1262;
wire wire75;
wire wire579;
wire wire764;
wire n_n1140;
wire wire699;
wire n_n1127;
wire wire1052;
wire n_n1320;
wire n_n1240;
wire n_n4124;
wire wire629;
wire wire631;
wire n_n1242;
wire n_n1243;
wire wire223;
wire wire168;
wire wire1060;
wire n_n852;
wire n_n1058;
wire n_n3604;
wire n_n3610;
wire wire697;
wire wire1061;
wire n_n771;
wire n_n206;
wire wire516;
wire wire1062;
wire n_n825;
wire wire675;
wire wire1064;
wire wire1063;
wire n_n762;
wire n_n13;
wire n_n458;
wire wire1066;
wire n_n374;
wire wire486;
wire n_n2738;
wire n_n462;
wire wire1069;
wire n_n346;
wire n_n203;
wire n_n16;
wire n_n285;
wire n_n43;
wire n_n51;
wire n_n82;
wire n_n68;
wire n_n113;
wire n_n86;
wire n_n79;
wire n_n103;
wire n_n36;
wire n_n284;
wire n_n44;
wire n_n73;
wire n_n72;
wire n_n85;
wire n_n15;
wire wire1071;
wire wire277;
wire n_n4950;
wire n_n4924;
wire wire255;
wire n_n4871;
wire n_n4838;
wire wire111;
wire n_n4730;
wire wire1076;
wire wire1079;
wire n_n6534;
wire n_n4330;
wire n_n4313;
wire wire180;
wire wire70;
wire wire125;
wire wire118;
wire n_n4806;
wire wire709;
wire wire372;
wire wire894;
wire wire141;
wire n_n1341;
wire n_n3974;
wire n_n4090;
wire wire462;
wire wire464;
wire n_n3918;
wire n_n6879;
wire wire1089;
wire n_n3919;
wire n_n3506;
wire wire378;
wire wire455;
wire wire485;
wire wire179;
wire n_n3781;
wire wire676;
wire n_n3184;
wire wire712;
wire n_n3116;
wire n_n4005;
wire wire446;
wire n_n35;
wire n_n4922;
wire n_n4921;
wire n_n4076;
wire n_n3768;
wire n_n2467;
wire wire386;
wire wire484;
wire n_n2439;
wire wire1092;
wire n_n2149;
wire n_n4912;
wire n_n4916;
wire wire327;
wire wire1094;
wire wire191;
wire wire1096;
wire wire1095;
wire wire1097;
wire wire1102;
wire wire641;
wire n_n1756;
wire wire50;
wire wire645;
wire n_n1286;
wire n_n1148;
wire n_n1255;
wire n_n6848;
wire wire479;
wire wire656;
wire n_n1137;
wire n_n62;
wire n_n1157;
wire wire1112;
wire n_n1151;
wire wire1113;
wire n_n1102;
wire n_n1147;
wire n_n4675;
wire n_n4681;
wire n_n1604;
wire wire497;
wire n_n1101;
wire n_n1152;
wire n_n1154;
wire n_n3881;
wire wire784;
wire n_n1103;
wire wire91;
wire wire647;
wire wire1119;
wire n_n803;
wire wire356;
wire n_n850;
wire wire335;
wire wire725;
wire wire1121;
wire wire1120;
wire n_n770;
wire n_n4628;
wire wire727;
wire n_n365;
wire n_n429;
wire n_n343;
wire n_n423;
wire n_n361;
wire n_n363;
wire n_n342;
wire n_n367;
wire n_n369;
wire wire809;
wire wire1128;
wire n_n344;
wire n_n143;
wire n_n116;
wire n_n39;
wire n_n77;
wire n_n67;
wire n_n83;
wire wire1130;
wire wire1132;
wire wire190;
wire n_n4941;
wire n_n4942;
wire wire728;
wire wire729;
wire n_n5685;
wire n_n4416;
wire n_n4418;
wire wire794;
wire n_n4394;
wire n_n4381;
wire n_n3850;
wire wire473;
wire n_n4307;
wire wire124;
wire n_n4929;
wire wire212;
wire wire250;
wire wire1141;
wire n_n4279;
wire n_n3978;
wire n_n1346;
wire n_n884;
wire n_n3908;
wire n_n3778;
wire n_n3229;
wire wire740;
wire wire55;
wire wire741;
wire n_n1555;
wire wire626;
wire n_n3791;
wire wire591;
wire wire736;
wire n_n2815;
wire n_n2982;
wire wire349;
wire wire876;
wire n_n3097;
wire n_n3092;
wire n_n3093;
wire n_n3173;
wire n_n2882;
wire n_n3864;
wire wire780;
wire n_n2702;
wire wire654;
wire wire1149;
wire n_n2398;
wire wire1150;
wire n_n2724;
wire wire1152;
wire wire1156;
wire n_n2133;
wire wire388;
wire wire747;
wire n_n2132;
wire wire391;
wire wire1158;
wire n_n2080;
wire wire1159;
wire n_n2129;
wire wire1161;
wire n_n2079;
wire n_n2274;
wire wire78;
wire wire1163;
wire n_n22;
wire wire49;
wire n_n1217;
wire n_n4687;
wire n_n1284;
wire wire1167;
wire wire1169;
wire n_n1138;
wire wire85;
wire wire750;
wire n_n1433;
wire wire41;
wire wire932;
wire wire1171;
wire n_n1120;
wire n_n1476;
wire n_n1126;
wire n_n1142;
wire n_n1099;
wire n_n3843;
wire wire662;
wire n_n1584;
wire wire706;
wire wire406;
wire n_n952;
wire n_n819;
wire n_n101;
wire wire930;
wire n_n5673;
wire n_n59;
wire n_n148;
wire n_n90;
wire wire1181;
wire wire1187;
wire wire1186;
wire n_n5007;
wire wire936;
wire n_n4938;
wire wire760;
wire wire761;
wire wire762;
wire n_n4728;
wire wire247;
wire wire119;
wire wire763;
wire wire541;
wire wire585;
wire n_n4183;
wire wire376;
wire n_n4770;
wire n_n4160;
wire n_n1645;
wire wire586;
wire wire767;
wire n_n3136;
wire n_n3309;
wire wire463;
wire wire1192;
wire n_n3124;
wire wire681;
wire n_n3123;
wire n_n3099;
wire n_n3101;
wire n_n3587;
wire wire770;
wire wire771;
wire n_n3103;
wire n_n3104;
wire wire553;
wire wire653;
wire wire548;
wire wire773;
wire wire774;
wire wire1194;
wire n_n2665;
wire wire1196;
wire wire1195;
wire wire1198;
wire wire1201;
wire n_n1765;
wire n_n1697;
wire wire690;
wire wire835;
wire n_n1684;
wire n_n1703;
wire n_n1704;
wire n_n1752;
wire n_n1680;
wire wire56;
wire n_n1356;
wire n_n1208;
wire n_n639;
wire wire42;
wire wire694;
wire wire869;
wire n_n1121;
wire n_n876;
wire n_n790;
wire n_n7354;
wire wire743;
wire wire1213;
wire n_n349;
wire n_n7246;
wire wire833;
wire n_n351;
wire n_n385;
wire wire642;
wire wire1217;
wire n_n49;
wire wire590;
wire n_n5051;
wire wire1223;
wire n_n5017;
wire wire1226;
wire n_n5008;
wire wire1229;
wire n_n4729;
wire n_n4633;
wire wire705;
wire wire1230;
wire n_n4261;
wire wire1231;
wire n_n4218;
wire n_n4199;
wire wire140;
wire wire157;
wire n_n1370;
wire n_n4003;
wire wire309;
wire wire571;
wire wire737;
wire wire1234;
wire n_n3928;
wire n_n3659;
wire wire1237;
wire n_n3598;
wire wire208;
wire n_n3209;
wire wire383;
wire wire628;
wire n_n3135;
wire n_n4644;
wire n_n4636;
wire wire317;
wire n_n3121;
wire n_n2890;
wire n_n3122;
wire n_n4632;
wire wire487;
wire wire742;
wire wire931;
wire wire1241;
wire n_n2876;
wire n_n3731;
wire n_n1597;
wire n_n2437;
wire n_n2429;
wire wire271;
wire wire472;
wire n_n1788;
wire n_n1715;
wire wire1250;
wire wire1249;
wire wire1248;
wire n_n1792;
wire wire158;
wire wire1251;
wire n_n1690;
wire n_n1440;
wire wire300;
wire n_n1173;
wire n_n1210;
wire n_n6820;
wire wire1253;
wire wire1254;
wire n_n789;
wire wire320;
wire wire1257;
wire n_n370;
wire wire1259;
wire n_n345;
wire n_n377;
wire n_n464;
wire wire688;
wire wire798;
wire wire1261;
wire n_n347;
wire n_n96;
wire n_n5048;
wire wire315;
wire wire1265;
wire wire1264;
wire wire326;
wire wire1271;
wire n_n5005;
wire n_n4911;
wire wire632;
wire wire198;
wire wire137;
wire wire112;
wire wire80;
wire n_n3736;
wire n_n1339;
wire n_n3579;
wire wire1279;
wire wire204;
wire n_n4674;
wire n_n3703;
wire n_n3127;
wire n_n2875;
wire n_n2145;
wire wire1286;
wire n_n1785;
wire wire1291;
wire wire1290;
wire wire1289;
wire n_n1298;
wire wire687;
wire n_n1212;
wire wire374;
wire wire434;
wire wire799;
wire n_n1123;
wire wire88;
wire n_n3615;
wire wire1305;
wire n_n5664;
wire wire793;
wire wire874;
wire wire1307;
wire wire1311;
wire n_n407;
wire n_n408;
wire n_n340;
wire n_n4736;
wire wire481;
wire wire72;
wire wire273;
wire wire219;
wire n_n4259;
wire wire721;
wire n_n4214;
wire n_n4256;
wire n_n4255;
wire wire465;
wire n_n4774;
wire n_n3786;
wire n_n3782;
wire wire723;
wire wire1320;
wire n_n3382;
wire n_n4676;
wire n_n4686;
wire n_n3722;
wire wire1322;
wire n_n3221;
wire wire1323;
wire n_n3128;
wire wire1326;
wire wire298;
wire wire521;
wire n_n5675;
wire wire1327;
wire n_n2146;
wire wire429;
wire wire1329;
wire wire1330;
wire n_n1774;
wire n_n1710;
wire n_n1536;
wire wire1333;
wire n_n1295;
wire n_n1641;
wire wire1334;
wire n_n4915;
wire wire589;
wire wire679;
wire n_n3884;
wire n_n809;
wire wire1340;
wire wire483;
wire wire1343;
wire wire1345;
wire wire1344;
wire wire1347;
wire wire1346;
wire wire408;
wire wire933;
wire wire1349;
wire wire1348;
wire n_n352;
wire wire1354;
wire wire1357;
wire wire1355;
wire n_n339;
wire wire1359;
wire wire113;
wire n_n4913;
wire n_n4146;
wire n_n3925;
wire n_n3914;
wire n_n3930;
wire n_n3929;
wire n_n3991;
wire n_n3923;
wire wire478;
wire wire1363;
wire n_n3900;
wire n_n3920;
wire n_n3922;
wire n_n3899;
wire n_n3926;
wire n_n3901;
wire wire1368;
wire n_n3404;
wire n_n3486;
wire n_n3403;
wire n_n3372;
wire n_n2713;
wire wire121;
wire wire370;
wire wire493;
wire n_n3371;
wire n_n3398;
wire n_n3397;
wire wire788;
wire n_n3361;
wire n_n3132;
wire n_n2820;
wire n_n2818;
wire wire1371;
wire n_n2798;
wire wire1372;
wire wire1376;
wire n_n2158;
wire wire1378;
wire wire1377;
wire n_n4682;
wire n_n2172;
wire wire98;
wire wire482;
wire wire1379;
wire n_n2093;
wire n_n4666;
wire wire1383;
wire n_n2067;
wire wire425;
wire wire657;
wire n_n1804;
wire wire1387;
wire n_n1092;
wire wire73;
wire n_n1108;
wire n_n1109;
wire wire519;
wire n_n743;
wire n_n742;
wire wire139;
wire wire776;
wire n_n744;
wire wire929;
wire n_n5679;
wire wire1400;
wire wire546;
wire wire634;
wire n_n3915;
wire n_n3406;
wire n_n3932;
wire n_n3904;
wire n_n3806;
wire n_n3408;
wire n_n3374;
wire wire545;
wire n_n3375;
wire wire633;
wire n_n3362;
wire n_n2832;
wire n_n2817;
wire wire533;
wire n_n2797;
wire n_n2792;
wire n_n2793;
wire n_n2796;
wire n_n2140;
wire n_n2099;
wire wire1413;
wire wire1416;
wire n_n2097;
wire n_n2180;
wire wire1423;
wire n_n3770;
wire wire1424;
wire n_n1111;
wire wire276;
wire wire587;
wire wire66;
wire n_n3980;
wire wire1439;
wire n_n3895;
wire wire816;
wire n_n3709;
wire wire1442;
wire n_n2926;
wire wire882;
wire n_n2824;
wire n_n2799;
wire n_n2801;
wire wire1445;
wire n_n2830;
wire n_n2803;
wire n_n2804;
wire wire693;
wire n_n2154;
wire wire1449;
wire n_n2100;
wire wire1450;
wire wire1451;
wire wire823;
wire n_n1124;
wire n_n1093;
wire wire381;
wire n_n5677;
wire wire384;
wire wire621;
wire n_n3913;
wire n_n3133;
wire wire1463;
wire n_n2808;
wire n_n2822;
wire n_n2821;
wire n_n2806;
wire wire792;
wire n_n2155;
wire wire1469;
wire n_n2088;
wire n_n3751;
wire wire380;
wire wire826;
wire wire1475;
wire wire1474;
wire wire101;
wire n_n2827;
wire n_n4914;
wire n_n2813;
wire wire829;
wire wire1483;
wire wire1484;
wire wire330;
wire wire1485;
wire n_n2085;
wire wire1486;
wire wire624;
wire wire1489;
wire wire1488;
wire wire1491;
wire wire1492;
wire n_n834;
wire n_n560;
wire n_n5009;
wire wire716;
wire wire821;
wire n_n2837;
wire n_n2086;
wire n_n2083;
wire n_n1598;
wire wire704;
wire n_n3523;
wire wire1514;
wire n_n1591;
wire wire144;
wire wire877;
wire n_n618;
wire n_n438;
wire wire1517;
wire n_n4781;
wire n_n4733;
wire n_n4773;
wire n_n4680;
wire wire468;
wire wire1528;
wire wire369;
wire wire1530;
wire wire233;
wire wire1540;
wire n_n4489;
wire n_n4677;
wire wire371;
wire wire1545;
wire n_n4598;
wire n_n4585;
wire n_n4555;
wire n_n3711;
wire n_n3710;
wire wire1547;
wire n_n4536;
wire n_n5672;
wire wire1552;
wire n_n3390;
wire n_n3624;
wire n_n3634;
wire n_n3636;
wire wire1555;
wire n_n3550;
wire wire1557;
wire n_n3380;
wire n_n3395;
wire n_n3369;
wire n_n3417;
wire n_n3378;
wire wire597;
wire n_n2597;
wire n_n2598;
wire n_n2579;
wire wire154;
wire n_n1781;
wire n_n785;
wire n_n413;
wire wire471;
wire wire658;
wire n_n359;
wire wire136;
wire n_n4732;
wire wire147;
wire wire1575;
wire n_n4685;
wire wire1577;
wire n_n4556;
wire n_n3638;
wire n_n3650;
wire n_n3629;
wire n_n3424;
wire n_n3379;
wire wire1585;
wire n_n3367;
wire n_n3393;
wire n_n3360;
wire n_n2833;
wire n_n2633;
wire n_n2599;
wire wire812;
wire n_n2580;
wire wire1593;
wire wire1594;
wire n_n1713;
wire wire1597;
wire wire1596;
wire wire1599;
wire wire494;
wire wire1600;
wire n_n1691;
wire wire514;
wire n_n787;
wire n_n749;
wire wire1606;
wire n_n750;
wire n_n409;
wire n_n4545;
wire n_n4548;
wire n_n4549;
wire wire54;
wire wire609;
wire n_n2603;
wire n_n2577;
wire n_n2573;
wire n_n2578;
wire n_n2572;
wire n_n2583;
wire n_n2582;
wire wire1627;
wire n_n1709;
wire wire1630;
wire n_n1688;
wire n_n1706;
wire n_n1705;
wire n_n1687;
wire n_n1711;
wire wire102;
wire n_n1689;
wire wire1637;
wire n_n758;
wire wire275;
wire wire887;
wire wire1640;
wire wire1639;
wire wire1638;
wire wire1641;
wire n_n739;
wire wire1645;
wire wire1648;
wire wire1647;
wire n_n4723;
wire n_n4744;
wire n_n4725;
wire wire672;
wire wire199;
wire n_n3803;
wire n_n4544;
wire n_n4551;
wire n_n3708;
wire n_n4535;
wire wire1657;
wire n_n3364;
wire n_n3386;
wire n_n3385;
wire n_n2835;
wire wire1662;
wire wire1661;
wire n_n707;
wire wire1664;
wire n_n2656;
wire wire1668;
wire n_n1724;
wire wire426;
wire wire134;
wire wire544;
wire wire1669;
wire n_n755;
wire wire1670;
wire n_n756;
wire n_n738;
wire wire403;
wire wire1673;
wire n_n443;
wire wire175;
wire wire1678;
wire wire1677;
wire wire1676;
wire wire292;
wire wire1682;
wire wire1680;
wire wire1679;
wire wire1686;
wire wire1687;
wire n_n3637;
wire n_n3435;
wire n_n3383;
wire wire1693;
wire wire1696;
wire n_n1738;
wire wire379;
wire wire1699;
wire n_n741;
wire n_n740;
wire n_n732;
wire wire1700;
wire wire1703;
wire wire1707;
wire wire1706;
wire n_n3686;
wire wire395;
wire n_n3642;
wire wire400;
wire wire1717;
wire wire182;
wire wire1723;
wire wire132;
wire wire236;
wire wire1730;
wire wire1732;
wire wire123;
wire wire1733;
wire wire1737;
wire n_n431;
wire wire1740;
wire n_n3645;
wire n_n3630;
wire wire1747;
wire wire225;
wire wire1753;
wire wire1752;
wire wire1755;
wire n_n2671;
wire n_n2657;
wire n_n2659;
wire wire1768;
wire n_n1761;
wire n_n1773;
wire wire1773;
wire wire1772;
wire wire1771;
wire wire1776;
wire wire1777;
wire n_n775;
wire n_n4542;
wire n_n4541;
wire wire1786;
wire n_n2433;
wire n_n1753;
wire wire622;
wire wire1793;
wire wire143;
wire wire1794;
wire wire1795;
wire n_n341;
wire wire1797;
wire wire1796;
wire n_n3658;
wire wire117;
wire wire1803;
wire n_n1692;
wire n_n2673;
wire wire1807;
wire n_n2431;
wire wire1812;
wire wire1814;
wire wire1813;
wire wire167;
wire wire1819;
wire wire1825;
wire n_n4539;
wire wire1829;
wire n_n4464;
wire wire879;
wire n_n2428;
wire wire1835;
wire wire1837;
wire wire1836;
wire wire1845;
wire wire1843;
wire wire1842;
wire wire1849;
wire wire43;
wire wire807;
wire wire47;
wire wire52;
wire wire53;
wire wire57;
wire wire58;
wire wire59;
wire wire61;
wire wire63;
wire wire64;
wire wire65;
wire wire71;
wire wire74;
wire wire76;
wire wire83;
wire wire84;
wire wire86;
wire wire87;
wire wire245;
wire wire95;
wire wire96;
wire wire97;
wire wire100;
wire wire103;
wire wire104;
wire wire105;
wire wire453;
wire wire110;
wire wire128;
wire wire130;
wire wire145;
wire wire288;
wire wire148;
wire wire149;
wire wire152;
wire wire161;
wire wire187;
wire wire195;
wire wire196;
wire wire197;
wire wire202;
wire wire203;
wire wire210;
wire wire214;
wire wire215;
wire wire220;
wire wire226;
wire wire227;
wire wire228;
wire wire229;
wire wire230;
wire wire231;
wire wire232;
wire wire235;
wire wire375;
wire wire240;
wire wire241;
wire wire242;
wire wire243;
wire wire246;
wire wire256;
wire wire262;
wire wire263;
wire wire266;
wire wire270;
wire wire274;
wire wire281;
wire wire282;
wire wire285;
wire wire287;
wire wire291;
wire wire294;
wire wire1852;
wire wire299;
wire wire304;
wire wire305;
wire wire306;
wire wire310;
wire wire311;
wire wire1853;
wire wire321;
wire wire325;
wire wire328;
wire wire331;
wire wire338;
wire wire342;
wire wire343;
wire wire345;
wire wire346;
wire wire347;
wire wire348;
wire wire351;
wire wire352;
wire wire357;
wire wire358;
wire wire361;
wire wire362;
wire wire363;
wire wire1855;
wire wire1856;
wire wire397;
wire wire398;
wire wire399;
wire wire405;
wire wire413;
wire wire414;
wire wire419;
wire wire424;
wire wire428;
wire wire431;
wire wire433;
wire wire435;
wire wire436;
wire wire437;
wire wire440;
wire wire441;
wire wire444;
wire wire448;
wire wire454;
wire wire1868;
wire wire1871;
wire wire1873;
wire wire1874;
wire wire1877;
wire wire1878;
wire wire1884;
wire wire1891;
wire wire1892;
wire wire1893;
wire wire1894;
wire wire1896;
wire wire1897;
wire wire1898;
wire wire1899;
wire wire1900;
wire wire1902;
wire wire1903;
wire wire1904;
wire wire1905;
wire wire1910;
wire wire1914;
wire wire1916;
wire wire1917;
wire wire1918;
wire wire1920;
wire wire1923;
wire wire1924;
wire wire1926;
wire wire1927;
wire wire1928;
wire wire1932;
wire wire1936;
wire wire1937;
wire wire1938;
wire wire1939;
wire wire1940;
wire wire1943;
wire wire1945;
wire wire1946;
wire wire1948;
wire wire1950;
wire wire1951;
wire wire1952;
wire wire1953;
wire wire857;
wire wire858;
wire wire1959;
wire wire962;
wire wire966;
wire wire965;
wire wire969;
wire wire968;
wire wire971;
wire wire1037;
wire wire1074;
wire wire1101;
wire wire1124;
wire wire1131;
wire wire1133;
wire wire1135;
wire wire1183;
wire wire1182;
wire wire1199;
wire wire1214;
wire wire1225;
wire wire1317;
wire wire1501;
wire wire1508;
wire wire1529;
wire wire1554;
wire wire1619;
wire wire1649;
wire wire1652;
wire wire1656;
wire wire1705;
wire wire1781;
wire wire1792;
wire wire1822;
wire wire238;
wire wire505;
wire wire510;
wire wire511;
wire wire529;
wire wire543;
wire wire550;
wire wire564;
wire wire580;
wire wire608;
wire wire847;
wire wire850;
wire wire855;
wire wire856;
wire wire862;
wire wire895;
wire wire1964;
wire wire1968;
wire wire1969;
wire wire1970;
wire wire1971;
wire wire1975;
wire wire1976;
wire wire1977;
wire wire1978;
wire wire1984;
wire wire1990;
wire wire1997;
wire wire2001;
wire wire2002;
wire wire2008;
wire wire2011;
wire wire2012;
wire wire2019;
wire wire2022;
wire wire2023;
wire wire2030;
wire wire2034;
wire wire2035;
wire wire2041;
wire wire2059;
wire wire2063;
wire wire2067;
wire wire2072;
wire wire2081;
wire wire2082;
wire wire2089;
wire wire2091;
wire wire2092;
wire wire2103;
wire wire2104;
wire wire2122;
wire wire2126;
wire wire2127;
wire wire2128;
wire wire2129;
wire wire2138;
wire wire2162;
wire wire2163;
wire wire2168;
wire wire2169;
wire wire2170;
wire wire2173;
wire wire2174;
wire wire2176;
wire wire2183;
wire wire2196;
wire wire2200;
wire wire2205;
wire wire2206;
wire wire2225;
wire wire2235;
wire wire2237;
wire wire2239;
wire wire2240;
wire wire2243;
wire wire2246;
wire wire2258;
wire wire2260;
wire wire2263;
wire wire2264;
wire wire2265;
wire wire2267;
wire wire2268;
wire wire2269;
wire wire2277;
wire wire2291;
wire wire2296;
wire wire2299;
wire wire2300;
wire wire2304;
wire wire2305;
wire wire2306;
wire wire2307;
wire wire2308;
wire wire2309;
wire wire2311;
wire wire2324;
wire wire2333;
wire wire2336;
wire wire2344;
wire wire2345;
wire wire2350;
wire wire2353;
wire wire2354;
wire wire2355;
wire wire2356;
wire wire2359;
wire wire2361;
wire wire2363;
wire wire2364;
wire wire2374;
wire wire2377;
wire wire2378;
wire wire2384;
wire wire2385;
wire wire2392;
wire wire2393;
wire wire2398;
wire wire2403;
wire wire2410;
wire wire2425;
wire wire2426;
wire wire2427;
wire wire2428;
wire wire2430;
wire wire2436;
wire wire2437;
wire wire2447;
wire wire2457;
wire wire2458;
wire wire2463;
wire wire2464;
wire wire2465;
wire wire2472;
wire wire2473;
wire wire2474;
wire wire2478;
wire wire2479;
wire wire2486;
wire wire2491;
wire wire2495;
wire wire2496;
wire wire2503;
wire wire2507;
wire wire2508;
wire wire2516;
wire wire2520;
wire wire2521;
wire wire2525;
wire wire2526;
wire wire2532;
wire wire2533;
wire wire2534;
wire wire2542;
wire wire2543;
wire wire2544;
wire wire2545;
wire wire2550;
wire wire2551;
wire wire2560;
wire wire2561;
wire wire2566;
wire wire2571;
wire wire2572;
wire wire2581;
wire wire2583;
wire wire2593;
wire wire2594;
wire wire2596;
wire wire2597;
wire wire2601;
wire wire2602;
wire wire2623;
wire wire2631;
wire wire2637;
wire wire2638;
wire wire2640;
wire wire2652;
wire wire2659;
wire wire2665;
wire wire2672;
wire wire2673;
wire wire2676;
wire wire2686;
wire wire2692;
wire wire2698;
wire wire2699;
wire wire2703;
wire wire2704;
wire wire2708;
wire wire2709;
wire wire2725;
wire wire2726;
wire wire2740;
wire wire2745;
wire wire2774;
wire wire2775;
wire wire2776;
wire wire2777;
wire wire2780;
wire wire2781;
wire wire2784;
wire wire2785;
wire wire2790;
wire wire2798;
wire wire2804;
wire wire2808;
wire wire2811;
wire wire2813;
wire wire2814;
wire wire2822;
wire wire2825;
wire wire2827;
wire wire2830;
wire wire2831;
wire wire2839;
wire wire2842;
wire wire2845;
wire wire2846;
wire wire2854;
wire wire2858;
wire wire2864;
wire wire2874;
wire wire2879;
wire wire2883;
wire wire2885;
wire wire2888;
wire wire2889;
wire wire2893;
wire wire2901;
wire wire2902;
wire wire2906;
wire wire2907;
wire wire2912;
wire wire2913;
wire wire2917;
wire wire2918;
wire wire2919;
wire wire2920;
wire wire2927;
wire wire2928;
wire wire2929;
wire wire2939;
wire wire2942;
wire wire2943;
wire wire2952;
wire wire2960;
wire wire2961;
wire wire2967;
wire wire2972;
wire wire2973;
wire wire2974;
wire wire2975;
wire wire2976;
wire wire2981;
wire wire2982;
wire wire2994;
wire wire2999;
wire wire3000;
wire wire3003;
wire wire3004;
wire wire3005;
wire wire3008;
wire wire3012;
wire wire3018;
wire wire3019;
wire wire3032;
wire wire3033;
wire wire3043;
wire wire3045;
wire wire3056;
wire wire3065;
wire wire3072;
wire wire3080;
wire wire3098;
wire wire3106;
wire wire3109;
wire wire3120;
wire wire3121;
wire wire3145;
wire wire3159;
wire wire3178;
wire wire3179;
wire wire3186;
wire wire3187;
wire wire3190;
wire wire3198;
wire wire3203;
wire wire3211;
wire wire3213;
wire wire3214;
wire wire3215;
wire wire3219;
wire wire3220;
wire wire3221;
wire wire3222;
wire wire3228;
wire wire3232;
wire wire3241;
wire wire3255;
wire wire3256;
wire wire3261;
wire wire3262;
wire wire3270;
wire wire3272;
wire wire3277;
wire wire3282;
wire wire3283;
wire wire3287;
wire wire3288;
wire wire3292;
wire wire3296;
wire wire3297;
wire wire3303;
wire wire3310;
wire wire3316;
wire wire3317;
wire wire3320;
wire wire3324;
wire wire3340;
wire wire3344;
wire wire3345;
wire wire3354;
wire wire3358;
wire wire3360;
wire wire3361;
wire wire3368;
wire wire3370;
wire wire3375;
wire wire3376;
wire wire3382;
wire wire3393;
wire wire3398;
wire wire3400;
wire wire3401;
wire wire3402;
wire wire3409;
wire wire3413;
wire wire3416;
wire wire3419;
wire wire3428;
wire wire3432;
wire wire3440;
wire wire3441;
wire wire3442;
wire wire3447;
wire wire3451;
wire wire3452;
wire wire3469;
wire wire3470;
wire wire3480;
wire wire3489;
wire wire3490;
wire wire3491;
wire wire3496;
wire wire3499;
wire wire3500;
wire wire3507;
wire wire3508;
wire wire3510;
wire wire3518;
wire wire3520;
wire wire3521;
wire wire3528;
wire wire3530;
wire wire3531;
wire wire3533;
wire wire3534;
wire wire3538;
wire wire3541;
wire wire3542;
wire wire3544;
wire wire3550;
wire wire3551;
wire wire3558;
wire wire3562;
wire wire3563;
wire wire3565;
wire wire3572;
wire wire3576;
wire wire3577;
wire wire3578;
wire wire3579;
wire wire3584;
wire wire3585;
wire wire3588;
wire wire3594;
wire wire3595;
wire wire3600;
wire wire3612;
wire wire3613;
wire wire3619;
wire wire3620;
wire wire3626;
wire wire3627;
wire wire3629;
wire wire3636;
wire wire3642;
wire wire3653;
wire wire3660;
wire wire3661;
wire wire3662;
wire wire3664;
wire wire3665;
wire wire3673;
wire wire3674;
wire wire3680;
wire wire3681;
wire wire3682;
wire wire3688;
wire wire3689;
wire wire3698;
wire wire3702;
wire wire3707;
wire wire3708;
wire wire3712;
wire wire3720;
wire wire3725;
wire wire3726;
wire wire3733;
wire wire3736;
wire wire3745;
wire wire3754;
wire wire3755;
wire wire3758;
wire wire3762;
wire wire3764;
wire wire3771;
wire wire3778;
wire wire3790;
wire wire3791;
wire wire3800;
wire wire3821;
wire wire3830;
wire wire3831;
wire wire3837;
wire wire3843;
wire wire3852;
wire wire3860;
wire wire3870;
wire wire3884;
wire wire3889;
wire wire3896;
wire wire3904;
wire wire3924;
wire wire3931;
wire wire3932;
wire wire3943;
wire wire3945;
wire wire3946;
wire wire3967;
wire wire3968;
wire wire3975;
wire wire3976;
wire wire3985;
wire wire3988;
wire wire3989;
wire wire4004;
wire wire4005;
wire wire4016;
wire wire4027;
wire wire4028;
wire wire4035;
wire wire4036;
wire wire4042;
wire wire4043;
wire wire4044;
wire wire4056;
wire wire4059;
wire wire4060;
wire wire4062;
wire wire4071;
wire wire4072;
wire wire4073;
wire wire4076;
wire wire4080;
wire wire4081;
wire wire4089;
wire wire4090;
wire wire4100;
wire wire4117;
wire wire4120;
wire wire4131;
wire wire4159;
wire wire4166;
wire wire4170;
wire wire4183;
wire wire4196;
wire wire4202;
wire wire4234;
wire wire4235;
wire wire4236;
wire wire4248;
wire wire4259;
wire wire4264;
wire wire4267;
wire wire4276;
wire wire4281;
wire wire4285;
wire wire4302;
wire wire4313;
wire wire4319;
wire wire4322;
wire wire4330;
wire wire4344;
wire wire4360;
wire wire4365;
wire wire4373;
wire wire4380;
wire wire4384;
wire wire4391;
wire wire4409;
wire wire4414;
wire wire4417;
wire wire4418;
wire wire4423;
wire wire4435;
wire wire4444;
wire wire4453;
wire wire4463;
wire wire4470;
wire wire4472;
wire wire4478;
wire wire4492;
wire wire4500;
wire wire4506;
wire wire4520;
wire wire4523;
wire wire4524;
wire wire4529;
wire wire4530;
wire wire4551;
wire wire4552;
wire wire4557;
wire wire4558;
wire wire4565;
wire wire4569;
wire wire4570;
wire wire4573;
wire wire4574;
wire wire4586;
wire wire4587;
wire wire4593;
wire wire4602;
wire wire4617;
wire wire4618;
wire wire4636;
wire wire4641;
wire wire4655;
wire wire4656;
wire wire4679;
wire wire4680;
wire wire4684;
wire wire4685;
wire wire4690;
wire wire4691;
wire wire4694;
wire wire4695;
wire wire4696;
wire wire4704;
wire wire4705;
wire wire4710;
wire wire4711;
wire wire4720;
wire wire4726;
wire wire4727;
wire wire4735;
wire wire4745;
wire wire4750;
wire wire4751;
wire wire4756;
wire wire4761;
wire wire4766;
wire wire4789;
wire wire4790;
wire wire4800;
wire wire4805;
wire wire4807;
wire wire4808;
wire wire4817;
wire wire4827;
wire wire4839;
wire wire4844;
wire wire4845;
wire wire4849;
wire wire4856;
wire wire4869;
wire wire4870;
wire wire4871;
wire wire4882;
wire wire4889;
wire wire4890;
wire wire4892;
wire wire4896;
wire wire4899;
wire wire4900;
wire wire4902;
wire wire4905;
wire wire4928;
wire wire4935;
wire wire4939;
wire wire4947;
wire wire4974;
wire wire5002;
wire wire5011;
wire wire5012;
wire wire5013;
wire wire5014;
wire wire5023;
wire wire5031;
wire wire5033;
wire wire5035;
wire wire5036;
wire wire5047;
wire wire5048;
wire wire5053;
wire wire5054;
wire wire5059;
wire wire5060;
wire wire5075;
wire wire5076;
wire wire5091;
wire wire5099;
wire wire5109;
wire wire5115;
wire wire5116;
wire wire5138;
wire wire5140;
wire wire5144;
wire wire5153;
wire wire5160;
wire wire5161;
wire wire5171;
wire wire5184;
wire wire5185;
wire wire5195;
wire wire5205;
wire wire5208;
wire wire5215;
wire wire5219;
wire wire5228;
wire wire5238;
wire wire5239;
wire wire5240;
wire wire5241;
wire wire5242;
wire wire5243;
wire wire5244;
wire wire5245;
wire wire5248;
wire wire5262;
wire wire5268;
wire wire5269;
wire wire5298;
wire wire5299;
wire wire5327;
wire wire5328;
wire wire5336;
wire wire5340;
wire wire5341;
wire wire5343;
wire wire5344;
wire wire5347;
wire wire5348;
wire wire5356;
wire wire5357;
wire wire5361;
wire wire5362;
wire wire5363;
wire wire5368;
wire wire5369;
wire wire5371;
wire wire5372;
wire wire5381;
wire wire5389;
wire wire5390;
wire wire5400;
wire wire5405;
wire wire5408;
wire wire5411;
wire wire5412;
wire wire5413;
wire wire5421;
wire wire5426;
wire wire5430;
wire wire5439;
wire wire5441;
wire wire5442;
wire wire5445;
wire wire5453;
wire wire5457;
wire wire5472;
wire wire5478;
wire wire5485;
wire wire5494;
wire wire5506;
wire wire5509;
wire wire5510;
wire wire5514;
wire wire5515;
wire wire5516;
wire wire5517;
wire wire5544;
wire wire5546;
wire wire5550;
wire wire5552;
wire wire5564;
wire wire5565;
wire wire5569;
wire wire5570;
wire wire5577;
wire wire5587;
wire wire5588;
wire wire5589;
wire wire5590;
wire wire5591;
wire wire5592;
wire wire5595;
wire wire5596;
wire wire5606;
wire wire5607;
wire wire5611;
wire wire5613;
wire wire5617;
wire wire5625;
wire wire5626;
wire wire5629;
wire wire5636;
wire wire5637;
wire wire5640;
wire wire5642;
wire wire5643;
wire wire5650;
wire wire5651;
wire wire5656;
wire wire5657;
wire wire5660;
wire wire5661;
wire wire5671;
wire wire5681;
wire wire5682;
wire wire5683;
wire wire5699;
wire wire5700;
wire wire5709;
wire wire5710;
wire wire5711;
wire wire5718;
wire wire5720;
wire wire5721;
wire wire5725;
wire wire5726;
wire wire5728;
wire wire5733;
wire wire5734;
wire wire5743;
wire wire5744;
wire wire5749;
wire wire5750;
wire wire5754;
wire wire5758;
wire wire5775;
wire wire5778;
wire wire5780;
wire wire5797;
wire wire5812;
wire wire5813;
wire wire5824;
wire wire5834;
wire wire5835;
wire wire5843;
wire wire5844;
wire wire5848;
wire wire5849;
wire wire5850;
wire wire5854;
wire wire5855;
wire wire5861;
wire wire5862;
wire wire5863;
wire wire5874;
wire wire5875;
wire wire5876;
wire wire5877;
wire wire5878;
wire wire5879;
wire wire5880;
wire wire5885;
wire wire5893;
wire wire5900;
wire wire5910;
wire wire5922;
wire wire5923;
wire wire5931;
wire wire5936;
wire wire5941;
wire wire5953;
wire wire5955;
wire wire5957;
wire wire5959;
wire wire5960;
wire wire5973;
wire wire5985;
wire wire5988;
wire wire5990;
wire wire5999;
wire wire6004;
wire wire6008;
wire wire6009;
wire wire6014;
wire wire6020;
wire wire19191;
wire wire19192;
wire wire19194;
wire wire19195;
wire wire19197;
wire wire19198;
wire wire19205;
wire wire19206;
wire wire19207;
wire wire19208;
wire wire19211;
wire wire19212;
wire wire19213;
wire wire19215;
wire wire19216;
wire wire19217;
wire wire19220;
wire wire19221;
wire wire19223;
wire wire19228;
wire wire19230;
wire wire19233;
wire wire19235;
wire wire19236;
wire wire19237;
wire wire19238;
wire wire19239;
wire wire19240;
wire wire19241;
wire wire19243;
wire wire19244;
wire wire19245;
wire wire19246;
wire wire19248;
wire wire19249;
wire wire19250;
wire wire19252;
wire wire19253;
wire wire19254;
wire wire19255;
wire wire19256;
wire wire19258;
wire wire19259;
wire wire19260;
wire wire19261;
wire wire19263;
wire wire19264;
wire wire19265;
wire wire19266;
wire wire19267;
wire wire19269;
wire wire19270;
wire wire19271;
wire wire19274;
wire wire19275;
wire wire19278;
wire wire19279;
wire wire19280;
wire wire19284;
wire wire19285;
wire wire19286;
wire wire19287;
wire wire19288;
wire wire19290;
wire wire19291;
wire wire19292;
wire wire19294;
wire wire19296;
wire wire19297;
wire wire19299;
wire wire19300;
wire wire19301;
wire wire19302;
wire wire19303;
wire wire19305;
wire wire19306;
wire wire19307;
wire wire19308;
wire wire19309;
wire wire19311;
wire wire19313;
wire wire19314;
wire wire19316;
wire wire19318;
wire wire19319;
wire wire19320;
wire wire19323;
wire wire19324;
wire wire19326;
wire wire19327;
wire wire19329;
wire wire19330;
wire wire19331;
wire wire19332;
wire wire19334;
wire wire19337;
wire wire19339;
wire wire19340;
wire wire19341;
wire wire19342;
wire wire19344;
wire wire19345;
wire wire19347;
wire wire19348;
wire wire19350;
wire wire19353;
wire wire19354;
wire wire19355;
wire wire19356;
wire wire19359;
wire wire19363;
wire wire19364;
wire wire19365;
wire wire19369;
wire wire19373;
wire wire19374;
wire wire19377;
wire wire19379;
wire wire19380;
wire wire19381;
wire wire19383;
wire wire19384;
wire wire19385;
wire wire19386;
wire wire19387;
wire wire19391;
wire wire19393;
wire wire19394;
wire wire19395;
wire wire19396;
wire wire19398;
wire wire19400;
wire wire19401;
wire wire19402;
wire wire19403;
wire wire19405;
wire wire19407;
wire wire19408;
wire wire19409;
wire wire19410;
wire wire19413;
wire wire19417;
wire wire19418;
wire wire19420;
wire wire19422;
wire wire19424;
wire wire19426;
wire wire19430;
wire wire19431;
wire wire19435;
wire wire19439;
wire wire19440;
wire wire19442;
wire wire19443;
wire wire19445;
wire wire19446;
wire wire19447;
wire wire19452;
wire wire19453;
wire wire19455;
wire wire19457;
wire wire19458;
wire wire19460;
wire wire19461;
wire wire19465;
wire wire19466;
wire wire19467;
wire wire19469;
wire wire19470;
wire wire19472;
wire wire19473;
wire wire19475;
wire wire19478;
wire wire19480;
wire wire19485;
wire wire19489;
wire wire19490;
wire wire19491;
wire wire19493;
wire wire19495;
wire wire19497;
wire wire19498;
wire wire19499;
wire wire19502;
wire wire19504;
wire wire19506;
wire wire19507;
wire wire19508;
wire wire19511;
wire wire19512;
wire wire19515;
wire wire19516;
wire wire19519;
wire wire19520;
wire wire19522;
wire wire19523;
wire wire19526;
wire wire19528;
wire wire19530;
wire wire19534;
wire wire19535;
wire wire19536;
wire wire19537;
wire wire19539;
wire wire19540;
wire wire19541;
wire wire19544;
wire wire19546;
wire wire19548;
wire wire19549;
wire wire19550;
wire wire19553;
wire wire19554;
wire wire19556;
wire wire19558;
wire wire19559;
wire wire19560;
wire wire19565;
wire wire19566;
wire wire19567;
wire wire19568;
wire wire19571;
wire wire19573;
wire wire19575;
wire wire19576;
wire wire19577;
wire wire19578;
wire wire19579;
wire wire19581;
wire wire19582;
wire wire19586;
wire wire19588;
wire wire19592;
wire wire19593;
wire wire19598;
wire wire19599;
wire wire19601;
wire wire19602;
wire wire19604;
wire wire19605;
wire wire19608;
wire wire19609;
wire wire19610;
wire wire19613;
wire wire19614;
wire wire19617;
wire wire19619;
wire wire19620;
wire wire19622;
wire wire19624;
wire wire19625;
wire wire19626;
wire wire19628;
wire wire19631;
wire wire19632;
wire wire19633;
wire wire19636;
wire wire19638;
wire wire19642;
wire wire19644;
wire wire19645;
wire wire19648;
wire wire19654;
wire wire19655;
wire wire19657;
wire wire19659;
wire wire19661;
wire wire19663;
wire wire19665;
wire wire19668;
wire wire19669;
wire wire19671;
wire wire19674;
wire wire19675;
wire wire19677;
wire wire19682;
wire wire19683;
wire wire19685;
wire wire19687;
wire wire19691;
wire wire19692;
wire wire19693;
wire wire19696;
wire wire19698;
wire wire19701;
wire wire19703;
wire wire19704;
wire wire19705;
wire wire19706;
wire wire19707;
wire wire19709;
wire wire19710;
wire wire19711;
wire wire19712;
wire wire19713;
wire wire19714;
wire wire19717;
wire wire19718;
wire wire19720;
wire wire19723;
wire wire19724;
wire wire19725;
wire wire19727;
wire wire19728;
wire wire19730;
wire wire19732;
wire wire19733;
wire wire19735;
wire wire19736;
wire wire19738;
wire wire19741;
wire wire19742;
wire wire19744;
wire wire19747;
wire wire19749;
wire wire19752;
wire wire19753;
wire wire19754;
wire wire19755;
wire wire19757;
wire wire19758;
wire wire19759;
wire wire19761;
wire wire19763;
wire wire19764;
wire wire19766;
wire wire19768;
wire wire19770;
wire wire19772;
wire wire19773;
wire wire19774;
wire wire19776;
wire wire19778;
wire wire19780;
wire wire19783;
wire wire19784;
wire wire19787;
wire wire19790;
wire wire19791;
wire wire19793;
wire wire19797;
wire wire19798;
wire wire19801;
wire wire19802;
wire wire19803;
wire wire19807;
wire wire19808;
wire wire19810;
wire wire19812;
wire wire19814;
wire wire19817;
wire wire19818;
wire wire19819;
wire wire19821;
wire wire19822;
wire wire19825;
wire wire19826;
wire wire19829;
wire wire19830;
wire wire19831;
wire wire19833;
wire wire19834;
wire wire19835;
wire wire19837;
wire wire19838;
wire wire19842;
wire wire19843;
wire wire19846;
wire wire19847;
wire wire19848;
wire wire19849;
wire wire19852;
wire wire19853;
wire wire19854;
wire wire19855;
wire wire19856;
wire wire19857;
wire wire19859;
wire wire19860;
wire wire19862;
wire wire19864;
wire wire19865;
wire wire19867;
wire wire19868;
wire wire19869;
wire wire19871;
wire wire19872;
wire wire19874;
wire wire19878;
wire wire19881;
wire wire19882;
wire wire19887;
wire wire19888;
wire wire19890;
wire wire19892;
wire wire19893;
wire wire19896;
wire wire19899;
wire wire19900;
wire wire19903;
wire wire19904;
wire wire19906;
wire wire19909;
wire wire19914;
wire wire19916;
wire wire19918;
wire wire19919;
wire wire19921;
wire wire19925;
wire wire19926;
wire wire19927;
wire wire19928;
wire wire19930;
wire wire19931;
wire wire19935;
wire wire19936;
wire wire19938;
wire wire19941;
wire wire19943;
wire wire19944;
wire wire19946;
wire wire19948;
wire wire19949;
wire wire19952;
wire wire19953;
wire wire19954;
wire wire19955;
wire wire19956;
wire wire19957;
wire wire19958;
wire wire19959;
wire wire19961;
wire wire19963;
wire wire19965;
wire wire19967;
wire wire19969;
wire wire19971;
wire wire19973;
wire wire19974;
wire wire19977;
wire wire19978;
wire wire19980;
wire wire19981;
wire wire19984;
wire wire19986;
wire wire19987;
wire wire19988;
wire wire19989;
wire wire19990;
wire wire19996;
wire wire19997;
wire wire19998;
wire wire19999;
wire wire20000;
wire wire20001;
wire wire20002;
wire wire20004;
wire wire20007;
wire wire20008;
wire wire20011;
wire wire20012;
wire wire20015;
wire wire20016;
wire wire20017;
wire wire20020;
wire wire20021;
wire wire20023;
wire wire20027;
wire wire20028;
wire wire20030;
wire wire20031;
wire wire20033;
wire wire20034;
wire wire20038;
wire wire20041;
wire wire20042;
wire wire20045;
wire wire20047;
wire wire20048;
wire wire20051;
wire wire20052;
wire wire20054;
wire wire20055;
wire wire20056;
wire wire20060;
wire wire20061;
wire wire20066;
wire wire20068;
wire wire20070;
wire wire20072;
wire wire20073;
wire wire20075;
wire wire20076;
wire wire20081;
wire wire20083;
wire wire20084;
wire wire20085;
wire wire20086;
wire wire20087;
wire wire20088;
wire wire20089;
wire wire20090;
wire wire20092;
wire wire20093;
wire wire20094;
wire wire20095;
wire wire20096;
wire wire20099;
wire wire20100;
wire wire20101;
wire wire20103;
wire wire20104;
wire wire20107;
wire wire20108;
wire wire20111;
wire wire20113;
wire wire20115;
wire wire20117;
wire wire20119;
wire wire20121;
wire wire20122;
wire wire20125;
wire wire20126;
wire wire20129;
wire wire20131;
wire wire20132;
wire wire20133;
wire wire20134;
wire wire20136;
wire wire20137;
wire wire20141;
wire wire20142;
wire wire20144;
wire wire20145;
wire wire20147;
wire wire20149;
wire wire20150;
wire wire20152;
wire wire20153;
wire wire20155;
wire wire20156;
wire wire20157;
wire wire20160;
wire wire20161;
wire wire20164;
wire wire20166;
wire wire20169;
wire wire20171;
wire wire20173;
wire wire20174;
wire wire20176;
wire wire20179;
wire wire20180;
wire wire20182;
wire wire20184;
wire wire20186;
wire wire20188;
wire wire20190;
wire wire20191;
wire wire20192;
wire wire20193;
wire wire20194;
wire wire20195;
wire wire20199;
wire wire20200;
wire wire20203;
wire wire20205;
wire wire20206;
wire wire20209;
wire wire20212;
wire wire20213;
wire wire20215;
wire wire20216;
wire wire20219;
wire wire20220;
wire wire20224;
wire wire20227;
wire wire20228;
wire wire20232;
wire wire20236;
wire wire20238;
wire wire20240;
wire wire20245;
wire wire20248;
wire wire20253;
wire wire20254;
wire wire20256;
wire wire20257;
wire wire20258;
wire wire20259;
wire wire20262;
wire wire20264;
wire wire20265;
wire wire20268;
wire wire20269;
wire wire20271;
wire wire20273;
wire wire20275;
wire wire20277;
wire wire20278;
wire wire20279;
wire wire20282;
wire wire20284;
wire wire20285;
wire wire20287;
wire wire20289;
wire wire20290;
wire wire20293;
wire wire20297;
wire wire20299;
wire wire20300;
wire wire20301;
wire wire20304;
wire wire20306;
wire wire20307;
wire wire20308;
wire wire20309;
wire wire20310;
wire wire20313;
wire wire20314;
wire wire20315;
wire wire20316;
wire wire20319;
wire wire20323;
wire wire20324;
wire wire20325;
wire wire20330;
wire wire20331;
wire wire20334;
wire wire20336;
wire wire20337;
wire wire20340;
wire wire20341;
wire wire20343;
wire wire20344;
wire wire20346;
wire wire20347;
wire wire20349;
wire wire20350;
wire wire20353;
wire wire20355;
wire wire20356;
wire wire20358;
wire wire20359;
wire wire20362;
wire wire20364;
wire wire20365;
wire wire20366;
wire wire20367;
wire wire20369;
wire wire20370;
wire wire20371;
wire wire20374;
wire wire20376;
wire wire20379;
wire wire20381;
wire wire20382;
wire wire20385;
wire wire20387;
wire wire20390;
wire wire20392;
wire wire20397;
wire wire20400;
wire wire20401;
wire wire20403;
wire wire20404;
wire wire20405;
wire wire20408;
wire wire20409;
wire wire20412;
wire wire20414;
wire wire20415;
wire wire20416;
wire wire20418;
wire wire20419;
wire wire20422;
wire wire20423;
wire wire20424;
wire wire20425;
wire wire20429;
wire wire20430;
wire wire20433;
wire wire20434;
wire wire20435;
wire wire20437;
wire wire20438;
wire wire20441;
wire wire20442;
wire wire20444;
wire wire20445;
wire wire20449;
wire wire20450;
wire wire20452;
wire wire20454;
wire wire20455;
wire wire20457;
wire wire20460;
wire wire20461;
wire wire20463;
wire wire20465;
wire wire20466;
wire wire20467;
wire wire20469;
wire wire20470;
wire wire20471;
wire wire20472;
wire wire20474;
wire wire20475;
wire wire20479;
wire wire20480;
wire wire20482;
wire wire20484;
wire wire20486;
wire wire20488;
wire wire20490;
wire wire20491;
wire wire20492;
wire wire20495;
wire wire20497;
wire wire20499;
wire wire20501;
wire wire20502;
wire wire20505;
wire wire20506;
wire wire20508;
wire wire20510;
wire wire20512;
wire wire20513;
wire wire20514;
wire wire20516;
wire wire20519;
wire wire20520;
wire wire20522;
wire wire20524;
wire wire20525;
wire wire20526;
wire wire20527;
wire wire20528;
wire wire20529;
wire wire20530;
wire wire20532;
wire wire20533;
wire wire20536;
wire wire20537;
wire wire20540;
wire wire20541;
wire wire20542;
wire wire20543;
wire wire20547;
wire wire20548;
wire wire20549;
wire wire20551;
wire wire20553;
wire wire20555;
wire wire20556;
wire wire20557;
wire wire20559;
wire wire20562;
wire wire20566;
wire wire20568;
wire wire20571;
wire wire20573;
wire wire20574;
wire wire20575;
wire wire20576;
wire wire20579;
wire wire20581;
wire wire20583;
wire wire20585;
wire wire20588;
wire wire20590;
wire wire20592;
wire wire20593;
wire wire20595;
wire wire20596;
wire wire20597;
wire wire20600;
wire wire20601;
wire wire20602;
wire wire20604;
wire wire20606;
wire wire20608;
wire wire20609;
wire wire20610;
wire wire20611;
wire wire20614;
wire wire20616;
wire wire20617;
wire wire20620;
wire wire20622;
wire wire20624;
wire wire20625;
wire wire20629;
wire wire20630;
wire wire20633;
wire wire20635;
wire wire20636;
wire wire20637;
wire wire20638;
wire wire20641;
wire wire20642;
wire wire20643;
wire wire20645;
wire wire20646;
wire wire20648;
wire wire20651;
wire wire20652;
wire wire20655;
wire wire20657;
wire wire20658;
wire wire20662;
wire wire20665;
wire wire20667;
wire wire20668;
wire wire20671;
wire wire20675;
wire wire20677;
wire wire20678;
wire wire20682;
wire wire20683;
wire wire20686;
wire wire20688;
wire wire20689;
wire wire20691;
wire wire20692;
wire wire20694;
wire wire20695;
wire wire20696;
wire wire20699;
wire wire20701;
wire wire20703;
wire wire20704;
wire wire20705;
wire wire20706;
wire wire20710;
wire wire20711;
wire wire20712;
wire wire20714;
wire wire20716;
wire wire20718;
wire wire20719;
wire wire20720;
wire wire20721;
wire wire20722;
wire wire20725;
wire wire20728;
wire wire20729;
wire wire20733;
wire wire20737;
wire wire20739;
wire wire20740;
wire wire20742;
wire wire20743;
wire wire20745;
wire wire20746;
wire wire20748;
wire wire20750;
wire wire20751;
wire wire20753;
wire wire20755;
wire wire20756;
wire wire20758;
wire wire20759;
wire wire20760;
wire wire20764;
wire wire20765;
wire wire20767;
wire wire20769;
wire wire20770;
wire wire20772;
wire wire20774;
wire wire20775;
wire wire20776;
wire wire20778;
wire wire20779;
wire wire20781;
wire wire20782;
wire wire20784;
wire wire20785;
wire wire20786;
wire wire20788;
wire wire20791;
wire wire20793;
wire wire20796;
wire wire20797;
wire wire20798;
wire wire20800;
wire wire20802;
wire wire20804;
wire wire20806;
wire wire20807;
wire wire20808;
wire wire20809;
wire wire20814;
wire wire20816;
wire wire20817;
wire wire20819;
wire wire20820;
wire wire20823;
wire wire20824;
wire wire20826;
wire wire20827;
wire wire20831;
wire wire20832;
wire wire20833;
wire wire20836;
wire wire20839;
wire wire20840;
wire wire20842;
wire wire20844;
wire wire20846;
wire wire20847;
wire wire20849;
wire wire20851;
wire wire20853;
wire wire20854;
wire wire20856;
wire wire20858;
wire wire20861;
wire wire20862;
wire wire20865;
wire wire20866;
wire wire20869;
wire wire20870;
wire wire20872;
wire wire20874;
wire wire20875;
wire wire20876;
wire wire20881;
wire wire20882;
wire wire20883;
wire wire20888;
wire wire20889;
wire wire20894;
wire wire20895;
wire wire20897;
wire wire20898;
wire wire20899;
wire wire20900;
wire wire20904;
wire wire20905;
wire wire20907;
wire wire20908;
wire wire20909;
wire wire20912;
wire wire20913;
wire wire20914;
wire wire20917;
wire wire20919;
wire wire20920;
wire wire20923;
wire wire20924;
wire wire20925;
wire wire20926;
wire wire20928;
wire wire20931;
wire wire20933;
wire wire20934;
wire wire20936;
wire wire20938;
wire wire20942;
wire wire20944;
wire wire20946;
wire wire20947;
wire wire20950;
wire wire20952;
wire wire20955;
wire wire20956;
wire wire20958;
wire wire20959;
wire wire20962;
wire wire20964;
wire wire20967;
wire wire20968;
wire wire20971;
wire wire20973;
wire wire20974;
wire wire20975;
wire wire20980;
wire wire20981;
wire wire20982;
wire wire20984;
wire wire20987;
wire wire20988;
wire wire20989;
wire wire20993;
wire wire20994;
wire wire20996;
wire wire20998;
wire wire20999;
wire wire21003;
wire wire21004;
wire wire21006;
wire wire21009;
wire wire21010;
wire wire21013;
wire wire21014;
wire wire21017;
wire wire21019;
wire wire21021;
wire wire21022;
wire wire21023;
wire wire21027;
wire wire21028;
wire wire21030;
wire wire21034;
wire wire21035;
wire wire21038;
wire wire21042;
wire wire21043;
wire wire21046;
wire wire21047;
wire wire21049;
wire wire21051;
wire wire21054;
wire wire21057;
wire wire21059;
wire wire21061;
wire wire21063;
wire wire21065;
wire wire21066;
wire wire21069;
wire wire21070;
wire wire21072;
wire wire21073;
wire wire21074;
wire wire21076;
wire wire21077;
wire wire21081;
wire wire21083;
wire wire21085;
wire wire21089;
wire wire21090;
wire wire21092;
wire wire21093;
wire wire21095;
wire wire21098;
wire wire21101;
wire wire21103;
wire wire21105;
wire wire21108;
wire wire21109;
wire wire21110;
wire wire21113;
wire wire21114;
wire wire21116;
wire wire21118;
wire wire21120;
wire wire21122;
wire wire21125;
wire wire21127;
wire wire21129;
wire wire21131;
wire wire21134;
wire wire21135;
wire wire21136;
wire wire21138;
wire wire21141;
wire wire21142;
wire wire21143;
wire wire21146;
wire wire21148;
wire wire21151;
wire wire21153;
wire wire21154;
wire wire21157;
wire wire21159;
wire wire21160;
wire wire21163;
wire wire21164;
wire wire21165;
wire wire21168;
wire wire21169;
wire wire21170;
wire wire21173;
wire wire21174;
wire wire21175;
wire wire21178;
wire wire21180;
wire wire21182;
wire wire21183;
wire wire21186;
wire wire21188;
wire wire21190;
wire wire21191;
wire wire21193;
wire wire21195;
wire wire21196;
wire wire21197;
wire wire21200;
wire wire21201;
wire wire21203;
wire wire21204;
wire wire21206;
wire wire21208;
wire wire21211;
wire wire21212;
wire wire21213;
wire wire21214;
wire wire21215;
wire wire21217;
wire wire21218;
wire wire21220;
wire wire21221;
wire wire21223;
wire wire21224;
wire wire21225;
wire wire21228;
wire wire21230;
wire wire21231;
wire wire21232;
wire wire21233;
wire wire21234;
wire wire21236;
wire wire21238;
wire wire21240;
wire wire21243;
wire wire21245;
wire wire21247;
wire wire21248;
wire wire21250;
wire wire21252;
wire wire21253;
wire wire21257;
wire wire21258;
wire wire21260;
wire wire21261;
wire wire21263;
wire wire21264;
wire wire21266;
wire wire21268;
wire wire21269;
wire wire21271;
wire wire21272;
wire wire21273;
wire wire21274;
wire wire21276;
wire wire21277;
wire wire21278;
wire wire21279;
wire wire21280;
wire wire21281;
wire wire21284;
wire wire21285;
wire wire21286;
wire wire21288;
wire wire21290;
wire wire21293;
wire wire21296;
wire wire21297;
wire wire21298;
wire wire21299;
wire wire21302;
wire wire21303;
wire wire21306;
wire wire21307;
wire wire21309;
wire wire21310;
wire wire21313;
wire wire21314;
wire wire21315;
wire wire21316;
wire wire21318;
wire wire21322;
wire wire21323;
wire wire21328;
wire wire21329;
wire wire21330;
wire wire21332;
wire wire21333;
wire wire21334;
wire wire21335;
wire wire21337;
wire wire21339;
wire wire21340;
wire wire21341;
wire wire21342;
wire wire21343;
wire wire21345;
wire wire21346;
wire wire21347;
wire wire21348;
wire wire21350;
wire wire21352;
wire wire21353;
wire wire21354;
wire wire21356;
wire wire21359;
wire wire21362;
wire wire21364;
wire wire21365;
wire wire21367;
wire wire21370;
wire wire21371;
wire wire21372;
wire wire21374;
wire wire21377;
wire wire21379;
wire wire21381;
wire wire21383;
wire wire21384;
wire wire21385;
wire wire21387;
wire wire21389;
wire wire21390;
wire wire21391;
wire wire21393;
wire wire21394;
wire wire21396;
wire wire21402;
wire wire21403;
wire wire21404;
wire wire21408;
wire wire21409;
wire wire21414;
wire wire21415;
wire wire21416;
wire wire21417;
wire wire21424;
wire wire21425;
wire wire21426;
wire wire21427;
wire wire21428;
wire wire21431;
wire wire21432;
wire wire21434;
wire wire21435;
wire wire21438;
wire wire21440;
wire wire21442;
wire wire21443;
wire wire21445;
wire wire21446;
wire wire21448;
wire wire21449;
wire wire21453;
wire wire21455;
wire wire21457;
wire wire21458;
wire wire21459;
wire wire21462;
wire wire21463;
wire wire21464;
wire wire21466;
wire wire21467;
wire wire21470;
wire wire21474;
wire wire21477;
wire wire21478;
wire wire21479;
wire wire21482;
wire wire21483;
wire wire21486;
wire wire21487;
wire wire21488;
wire wire21490;
wire wire21491;
wire wire21493;
wire wire21494;
wire wire21497;
wire wire21499;
wire wire21500;
wire wire21501;
wire wire21505;
wire wire21506;
wire wire21507;
wire wire21508;
wire wire21512;
wire wire21514;
wire wire21516;
wire wire21517;
wire wire21521;
wire wire21522;
wire wire21525;
wire wire21529;
wire wire21530;
wire wire21531;
wire wire21533;
wire wire21536;
wire wire21537;
wire wire21538;
wire wire21540;
wire wire21541;
wire wire21544;
wire wire21545;
wire wire21546;
wire wire21549;
wire wire21551;
wire wire21554;
wire wire21555;
wire wire21557;
wire wire21560;
wire wire21561;
wire wire21562;
wire wire21565;
wire wire21566;
wire wire21569;
wire wire21572;
wire wire21574;
wire wire21576;
wire wire21578;
wire wire21579;
wire wire21583;
wire wire21584;
wire wire21586;
wire wire21588;
wire wire21590;
wire wire21593;
wire wire21596;
wire wire21599;
wire wire21600;
wire wire21603;
wire wire21605;
wire wire21608;
wire wire21609;
wire wire21612;
wire wire21614;
wire wire21615;
wire wire21616;
wire wire21620;
wire wire21621;
wire wire21624;
wire wire21626;
wire wire21627;
wire wire21628;
wire wire21631;
wire wire21633;
wire wire21635;
wire wire21636;
wire wire21637;
wire wire21639;
wire wire21640;
wire wire21642;
wire wire21643;
wire wire21646;
wire wire21647;
wire wire21648;
wire wire21649;
wire wire21650;
wire wire21651;
wire wire21652;
wire wire21655;
wire wire21657;
wire wire21658;
wire wire21660;
wire wire21662;
wire wire21663;
wire wire21665;
wire wire21666;
wire wire21668;
wire wire21670;
wire wire21671;
wire wire21673;
wire wire21675;
wire wire21676;
wire wire21677;
wire wire21678;
wire wire21681;
wire wire21683;
wire wire21686;
wire wire21687;
wire wire21690;
wire wire21691;
wire wire21694;
wire wire21695;
wire wire21697;
wire wire21699;
wire wire21700;
wire wire21701;
wire wire21702;
wire wire21705;
wire wire21706;
wire wire21709;
wire wire21711;
wire wire21713;
wire wire21714;
wire wire21715;
wire wire21716;
wire wire21718;
wire wire21719;
wire wire21721;
wire wire21723;
wire wire21724;
wire wire21726;
wire wire21728;
wire wire21729;
wire wire21730;
wire wire21732;
wire wire21733;
wire wire21735;
wire wire21737;
wire wire21739;
wire wire21741;
wire wire21742;
wire wire21743;
wire wire21744;
wire wire21746;
wire wire21748;
wire wire21749;
wire wire21751;
wire wire21752;
wire wire21753;
wire wire21756;
wire wire21757;
wire wire21759;
wire wire21760;
wire wire21761;
wire wire21762;
wire wire21764;
wire wire21766;
wire wire21767;
wire wire21769;
wire wire21770;
wire wire21771;
wire wire21772;
wire wire21775;
wire wire21777;
wire wire21778;
wire wire21780;
wire wire21781;
wire wire21783;
wire wire21784;
wire wire21785;
wire wire21786;
wire wire21789;
wire wire21790;
wire wire21792;
wire wire21794;
wire wire21797;
wire wire21798;
wire wire21799;
wire wire21804;
wire wire21805;
wire wire21807;
wire wire21808;
wire wire21811;
wire wire21813;
wire wire21814;
wire wire21815;
wire wire21817;
wire wire21820;
wire wire21821;
wire wire21823;
wire wire21825;
wire wire21827;
wire wire21828;
wire wire21832;
wire wire21834;
wire wire21837;
wire wire21838;
wire wire21842;
wire wire21844;
wire wire21845;
wire wire21847;
wire wire21849;
wire wire21850;
wire wire21853;
wire wire21855;
wire wire21857;
wire wire21859;
wire wire21860;
wire wire21861;
wire wire21862;
wire wire21864;
wire wire21865;
wire wire21866;
wire wire21867;
wire wire21868;
wire wire21869;
wire wire21872;
wire wire21874;
wire wire21877;
wire wire21881;
wire wire21884;
wire wire21885;
wire wire21888;
wire wire21889;
wire wire21892;
wire wire21893;
wire wire21895;
wire wire21896;
wire wire21900;
wire wire21902;
wire wire21904;
wire wire21907;
wire wire21910;
wire wire21912;
wire wire21913;
wire wire21914;
wire wire21918;
wire wire21920;
wire wire21922;
wire wire21923;
wire wire21925;
wire wire21926;
wire wire21927;
wire wire21928;
wire wire21929;
wire wire21930;
wire wire21933;
wire wire21935;
wire wire21938;
wire wire21939;
wire wire21941;
wire wire21943;
wire wire21944;
wire wire21946;
wire wire21948;
wire wire21950;
wire wire21953;
wire wire21954;
wire wire21956;
wire wire21958;
wire wire21959;
wire wire21960;
wire wire21962;
wire wire21963;
wire wire21965;
wire wire21966;
wire wire21968;
wire wire21969;
wire wire21970;
wire wire21971;
wire wire21973;
wire wire21975;
wire wire21977;
wire wire21979;
wire wire21980;
wire wire21981;
wire wire21982;
wire wire21983;
wire wire21984;
wire wire21985;
wire wire21987;
wire wire21988;
wire wire21991;
wire wire21992;
wire wire21993;
wire wire21995;
wire wire21997;
wire wire21998;
wire wire21999;
wire wire22000;
wire wire22001;
wire wire22002;
wire wire22004;
wire wire22005;
wire wire22007;
wire wire22009;
wire wire22010;
wire wire22012;
wire wire22014;
wire wire22016;
wire wire22017;
wire wire22020;
wire wire22022;
wire wire22024;
wire wire22026;
wire wire22029;
wire wire22033;
wire wire22034;
wire wire22035;
wire wire22039;
wire wire22040;
wire wire22041;
wire wire22043;
wire wire22044;
wire wire22047;
wire wire22048;
wire wire22050;
wire wire22052;
wire wire22053;
wire wire22054;
wire wire22058;
wire wire22059;
wire wire22061;
wire wire22064;
wire wire22066;
wire wire22067;
wire wire22070;
wire wire22071;
wire wire22075;
wire wire22076;
wire wire22079;
wire wire22081;
wire wire22082;
wire wire22083;
wire wire22084;
wire wire22087;
wire wire22088;
wire wire22090;
wire wire22093;
wire wire22095;
wire wire22097;
wire wire22099;
wire wire22101;
wire wire22104;
wire wire22106;
wire wire22108;
wire wire22109;
wire wire22110;
wire wire22112;
wire wire22115;
wire wire22117;
wire wire22119;
wire wire22121;
wire wire22124;
wire wire22125;
wire wire22126;
wire wire22129;
wire wire22130;
wire wire22134;
wire wire22135;
wire wire22136;
wire wire22139;
wire wire22140;
wire wire22142;
wire wire22145;
wire wire22146;
wire wire22148;
wire wire22149;
wire wire22154;
wire wire22157;
wire wire22159;
wire wire22160;
wire wire22162;
wire wire22164;
wire wire22167;
wire wire22168;
wire wire22169;
wire wire22170;
wire wire22171;
wire wire22174;
wire wire22176;
wire wire22181;
wire wire22184;
wire wire22185;
wire wire22187;
wire wire22188;
wire wire22190;
wire wire22193;
wire wire22195;
wire wire22196;
wire wire22197;
wire wire22201;
wire wire22203;
wire wire22206;
wire wire22208;
wire wire22210;
wire wire22211;
wire wire22213;
wire wire22214;
wire wire22217;
wire wire22219;
wire wire22220;
wire wire22227;
wire wire22228;
wire wire22231;
wire wire22232;
wire wire22236;
wire wire22238;
wire wire22240;
wire wire22241;
wire wire22242;
wire wire22244;
wire wire22245;
wire wire22248;
wire wire22249;
wire wire22250;
wire wire22253;
wire wire22255;
wire wire22257;
wire wire22259;
wire wire22262;
wire wire22264;
wire wire22266;
wire wire22270;
wire wire22273;
wire wire22275;
wire wire22276;
wire wire22277;
wire wire22280;
wire wire22282;
wire wire22286;
wire wire22287;
wire wire22290;
wire wire22291;
wire wire22294;
wire wire22298;
wire wire22300;
wire wire22302;
wire wire22304;
wire wire22305;
wire wire22308;
wire wire22309;
wire wire22310;
wire wire22312;
wire wire22314;
wire wire22315;
wire wire22316;
wire wire22317;
wire wire22319;
wire wire22321;
wire wire22322;
wire wire22326;
wire wire22327;
wire wire22328;
wire wire22330;
wire wire22331;
wire wire22332;
wire wire22334;
wire wire22335;
wire wire22336;
wire wire22337;
wire wire22338;
wire wire22340;
wire wire22341;
wire wire22343;
wire wire22345;
wire wire22346;
wire wire22348;
wire wire22351;
wire wire22352;
wire wire22355;
wire wire22356;
wire wire22358;
wire wire22360;
wire wire22361;
wire wire22363;
wire wire22366;
wire wire22368;
wire wire22369;
wire wire22370;
wire wire22372;
wire wire22374;
wire wire22376;
wire wire22378;
wire wire22379;
wire wire22380;
wire wire22382;
wire wire22383;
wire wire22384;
wire wire22387;
wire wire22389;
wire wire22391;
wire wire22393;
wire wire22395;
wire wire22399;
wire wire22400;
wire wire22401;
wire wire22403;
wire wire22404;
wire wire22407;
wire wire22408;
wire wire22409;
wire wire22412;
wire wire22414;
wire wire22415;
wire wire22416;
wire wire22421;
wire wire22426;
wire wire22429;
wire wire22431;
wire wire22432;
wire wire22435;
wire wire22436;
wire wire22438;
wire wire22440;
wire wire22443;
wire wire22446;
wire wire22447;
wire wire22449;
wire wire22451;
wire wire22454;
wire wire22456;
wire wire22457;
wire wire22459;
wire wire22461;
wire wire22463;
wire wire22464;
wire wire22467;
wire wire22468;
wire wire22469;
wire wire22471;
wire wire22473;
wire wire22474;
wire wire22475;
wire wire22476;
wire wire22477;
wire wire22481;
wire wire22483;
wire wire22485;
wire wire22487;
wire wire22488;
wire wire22489;
wire wire22490;
wire wire22491;
wire wire22492;
wire wire22493;
wire wire22494;
wire wire22495;
wire wire22496;
wire wire22502;
wire wire22504;
wire wire22506;
wire wire22510;
wire wire22511;
wire wire22512;
wire wire22513;
wire wire22515;
wire wire22516;
wire wire22518;
wire wire22519;
wire wire22522;
wire wire22523;
wire wire22524;
wire wire22527;
wire wire22531;
wire wire22532;
wire wire22533;
wire wire22535;
wire wire22536;
wire wire22537;
wire wire22538;
wire wire22539;
wire wire22540;
wire wire22541;
wire wire22543;
wire wire22544;
wire wire22546;
wire wire22547;
wire wire22548;
wire wire22551;
wire wire22552;
wire wire22556;
wire wire22557;
wire wire22558;
wire wire22561;
wire wire22562;
wire wire22565;
wire wire22566;
wire wire22567;
wire wire22570;
wire wire22571;
wire wire22572;
wire wire22573;
wire wire22574;
wire wire22575;
wire wire22576;
wire wire22578;
wire wire22581;
wire wire22587;
wire wire22588;
wire wire22590;
wire wire22593;
wire wire22594;
wire wire22596;
wire wire22597;
wire wire22598;
wire wire22599;
wire wire22600;
wire wire22602;
wire wire22605;
wire wire22606;
wire wire22610;
wire wire22611;
wire wire22613;
wire wire22616;
wire wire22618;
wire wire22620;
wire wire22625;
wire wire22626;
wire wire22629;
wire wire22630;
wire wire22631;
wire wire22633;
wire wire22635;
wire wire22636;
wire wire22637;
wire wire22638;
wire wire22639;
wire wire22640;
wire wire22642;
wire wire22643;
wire wire22646;
wire wire22647;
wire wire22648;
wire wire22650;
wire wire22651;
wire wire22652;
wire wire22654;
wire wire22657;
wire wire22658;
wire wire22659;
wire wire22662;
wire wire22663;
wire wire22664;
wire wire22665;
wire wire22667;
wire wire22668;
wire wire22670;
wire wire22672;
wire wire22674;
wire wire22675;
wire wire22676;
wire wire22678;
wire wire22680;
wire wire22681;
wire wire22683;
wire wire22684;
wire wire22685;
wire wire22686;
wire wire22687;
wire wire22689;
wire wire22692;
wire wire22693;
wire wire22695;
wire wire22696;
wire wire22698;
wire wire22700;
wire wire22701;
wire wire22703;
wire wire22704;
wire wire22708;
wire wire22709;
wire wire22710;
wire wire22711;
wire wire22712;
wire wire22714;
wire wire22717;
wire wire22719;
wire wire22720;
wire wire22722;
wire wire22725;
wire wire22727;
wire wire22730;
wire wire22731;
wire wire22732;
wire wire22734;
wire wire22736;
wire wire22740;
wire wire22742;
wire wire22744;
wire wire22746;
wire wire22748;
wire wire22752;
wire wire22754;
wire wire22757;
wire wire22758;
wire wire22761;
wire wire22762;
wire wire22763;
wire wire22764;
wire wire22765;
wire wire22766;
wire wire22769;
wire wire22772;
wire wire22775;
wire wire22776;
wire wire22778;
wire wire22780;
wire wire22781;
wire wire22783;
wire wire22785;
wire wire22786;
wire wire22787;
wire wire22788;
wire wire22792;
wire wire22793;
wire wire22795;
wire wire22796;
wire wire22797;
wire wire22801;
wire wire22803;
wire wire22804;
wire wire22805;
wire wire22806;
wire wire22809;
wire wire22812;
wire wire22814;
wire wire22816;
wire wire22818;
wire wire22820;
wire wire22822;
wire wire22827;
wire wire22829;
wire wire22830;
wire wire22833;
wire wire22835;
wire wire22837;
wire wire22839;
wire wire22841;
wire wire22843;
wire wire22844;
wire wire22847;
assign o_1_ = ( n_n5231 ) | ( n_n310 ) | ( wire19373 ) | ( wire19374 ) ;
 assign o_19_ = ( n_n5231 ) | ( n_n3621 ) | ( wire19592 ) | ( wire19593 ) ;
 assign o_2_ = ( n_n5231 ) | ( wire19601 ) | ( wire19602 ) ;
 assign o_0_ = ( n_n5231 ) | ( wire19622 ) ;
 assign o_29_ = ( n_n5231 ) | ( wire19648 ) ;
 assign o_39_ = ( n_n5231 ) | ( n_n5792 ) | ( wire5408 ) ;
 assign o_38_ = ( n_n5231 ) | ( n_n5794 ) | ( wire5405 ) ;
 assign o_25_ = ( n_n5231 ) | ( n_n4303 ) | ( wire19766 ) ;
 assign o_12_ = ( n_n5231 ) | ( wire19822 ) ;
 assign o_37_ = ( n_n5231 ) | ( n_n4982 ) | ( wire19838 ) ;
 assign o_26_ = ( n_n5231 ) | ( wire19846 ) | ( wire19847 ) ;
 assign o_11_ = ( n_n5231 ) | ( wire5109 ) | ( wire19855 ) | ( wire19860 ) ;
 assign o_36_ = ( n_n5231 ) | ( n_n4718 ) | ( wire19989 ) | ( wire19990 ) ;
 assign o_27_ = ( n_n5231 ) | ( n_n264  &  n_n153  &  n_n120 ) ;
 assign o_14_ = ( n_n5231 ) | ( wire20001 ) | ( wire20002 ) | ( wire20004 ) ;
 assign o_35_ = ( n_n5231 ) | ( n_n4705 ) | ( n_n4704 ) | ( wire20012 ) ;
 assign o_28_ = ( n_n5231 ) | ( n_n5224 ) ;
 assign o_13_ = ( n_n5231 ) | ( n_n2656 ) | ( n_n2657 ) | ( wire20115 ) ;
 assign o_34_ = ( n_n5231 ) | ( n_n4530 ) | ( wire20245 ) ;
 assign o_21_ = ( n_n5231 ) | ( wire20355 ) ;
 assign o_16_ = ( n_n5231 ) | ( n_n2789 ) | ( n_n2795 ) | ( wire20625 ) ;
 assign o_33_ = ( n_n5231 ) | ( n_n4512 ) | ( n_n4508 ) | ( wire20648 ) ;
 assign o_22_ = ( n_n5231 ) | ( n_n4186 ) | ( wire20657 ) | ( wire20658 ) ;
 assign o_15_ = ( n_n5247 ) | ( wire879 ) | ( wire19998 ) | ( wire20665 ) ;
 assign o_32_ = ( n_n5231 ) | ( n_n5797 ) | ( wire20667 ) | ( wire20671 ) ;
 assign o_23_ = ( n_n5231 ) | ( n_n4194 ) | ( wire20753 ) ;
 assign o_18_ = ( n_n5231 ) | ( n_n5235 ) ;
 assign o_31_ = ( n_n5231 ) | ( wire3945 ) | ( wire20919 ) | ( wire20920 ) ;
 assign o_24_ = ( n_n5231 ) | ( wire20924 ) ;
 assign o_17_ = ( n_n5231 ) | ( n_n3089 ) | ( n_n3094 ) | ( wire21154 ) ;
 assign o_30_ = ( n_n5231 ) | ( n_n4464 ) | ( wire21174 ) | ( wire21178 ) ;
 assign o_20_ = ( n_n5231 ) | ( n_n3892 ) | ( n_n3890 ) | ( wire21293 ) ;
 assign o_10_ = ( n_n5231 ) | ( wire21365 ) ;
 assign o_9_ = ( n_n5231 ) | ( n_n2058 ) | ( wire21620 ) | ( wire21621 ) ;
 assign o_7_ = ( n_n5231 ) | ( n_n1670 ) | ( wire21631 ) ;
 assign o_8_ = ( n_n5231 ) | ( n_n1679 ) | ( wire21904 ) ;
 assign o_5_ = ( n_n5231 ) | ( wire22331 ) | ( wire22334 ) ;
 assign o_6_ = ( n_n5247 ) | ( wire2474 ) ;
 assign o_3_ = ( n_n5231 ) | ( n_n333 ) | ( wire22594 ) ;
 assign o_4_ = ( n_n5231 ) | ( n_n731 ) | ( wire22847 ) ;
 assign n_n139 = ( n_n260  &  n_n229  &  n_n165 ) ;
 assign n_n151 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign n_n5686 = ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign n_n5231 = ( wire590 ) | ( n_n5005 ) | ( wire19306 ) | ( wire19359 ) ;
 assign n_n310 = ( wire19365 ) | ( n_n139  &  wire1475 ) ;
 assign n_n4476 = ( wire503 ) | ( wire48  &  n_n152 ) ;
 assign n_n4477 = ( n_n152  &  wire54 ) | ( n_n152  &  wire913  &  n_n220 ) ;
 assign wire394 = ( i_7_  &  i_6_  &  n_n260  &  n_n165 ) ;
 assign wire507 = ( i_7_  &  i_6_  &  wire927 ) | ( (~ i_7_)  &  i_6_  &  wire927 ) | ( i_7_  &  (~ i_6_)  &  wire927 ) | ( (~ i_7_)  &  i_6_  &  wire929 ) | ( i_7_  &  (~ i_6_)  &  wire929 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire929 ) ;
 assign wire893 = ( n_n152  &  n_n111 ) | ( n_n152  &  wire103 ) | ( n_n152  &  wire266 ) ;
 assign wire937 = ( n_n260  &  n_n208  &  n_n165 ) | ( n_n260  &  n_n273  &  n_n165 ) ;
 assign n_n863 = ( wire372 ) | ( wire386 ) | ( wire19380 ) ;
 assign n_n3625 = ( n_n3424 ) | ( n_n3642 ) | ( wire19431 ) | ( wire19435 ) ;
 assign n_n3626 = ( n_n3382 ) | ( wire19445 ) | ( wire19446 ) | ( wire19455 ) ;
 assign n_n3627 = ( n_n3645 ) | ( wire19472 ) | ( wire19473 ) | ( wire19480 ) ;
 assign n_n3621 = ( n_n3629 ) | ( n_n3630 ) | ( wire19530 ) ;
 assign n_n3631 = ( n_n4781 ) | ( n_n3711 ) | ( wire19544 ) | ( wire19546 ) ;
 assign n_n3661 = ( wire383 ) | ( wire19553 ) | ( wire19554 ) ;
 assign n_n3632 = ( n_n3659 ) | ( n_n3658 ) | ( wire19573 ) ;
 assign n_n124 = ( n_n229  &  n_n165  &  n_n284 ) ;
 assign n_n123 = ( n_n208  &  n_n165  &  n_n284 ) ;
 assign wire289 = ( i_7_  &  i_6_ ) | ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) ;
 assign wire364 = ( i_7_  &  i_6_  &  n_n165  &  n_n284 ) ;
 assign wire535 = ( i_7_  &  i_6_  &  n_n264  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign wire777 = ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign wire834 = ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n264 ) ;
 assign wire939 = ( n_n281  &  wire913 ) | ( n_n281  &  wire914 ) | ( n_n281  &  wire907 ) ;
 assign wire938 = ( wire48 ) | ( n_n110 ) | ( (~ i_9_)  &  (~ i_10_) ) ;
 assign n_n106 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign n_n5678 = ( (~ i_7_)  &  (~ i_6_)  &  n_n284  &  n_n116 ) ;
 assign n_n5671 = ( i_7_  &  i_6_  &  n_n264  &  n_n116 ) ;
 assign wire396 = ( n_n208  &  n_n165  &  n_n284 ) | ( n_n273  &  n_n165  &  n_n284 ) ;
 assign wire582 = ( wire777 ) | ( wire880 ) | ( n_n5677 ) | ( n_n5672 ) ;
 assign wire583 = ( wire5453 ) | ( wire19613 ) | ( wire19614 ) ;
 assign wire941 = ( n_n208  &  n_n165  &  n_n284 ) | ( n_n273  &  n_n165  &  n_n284 ) ;
 assign wire940 = ( n_n281  &  wire913 ) | ( n_n281  &  wire914 ) ;
 assign n_n272 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n118 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n4442 = ( wire19624 ) | ( wire19625 ) | ( wire19626 ) ;
 assign n_n4439 = ( n_n5792 ) | ( n_n5794 ) | ( wire5421 ) | ( wire19638 ) ;
 assign wire943 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign n_n231 = ( (~ i_7_)  &  i_6_ ) ;
 assign n_n5792 = ( i_4_  &  n_n231  &  n_n165  &  wire19290 ) ;
 assign n_n5794 = ( i_4_  &  n_n272  &  n_n165  &  wire19290 ) ;
 assign n_n4203 = ( wire573 ) | ( wire5389 ) | ( wire19654 ) | ( wire19655 ) ;
 assign n_n4206 = ( n_n4846 ) | ( n_n4842 ) | ( wire5381 ) | ( wire19659 ) ;
 assign n_n4306 = ( n_n1506 ) | ( n_n4313 ) | ( wire5356 ) | ( wire19677 ) ;
 assign n_n4807 = ( n_n6  &  wire75 ) | ( n_n6  &  wire911  &  n_n228 ) ;
 assign n_n4223 = ( n_n4808 ) | ( n_n4809 ) | ( wire541 ) ;
 assign n_n4224 = ( wire585 ) | ( wire5347 ) | ( wire5348 ) ;
 assign n_n4303 = ( n_n4307 ) | ( wire19717 ) | ( wire19718 ) | ( wire19736 ) ;
 assign n_n1 = ( n_n260  &  n_n273  &  n_n285 ) ;
 assign n_n2 = ( n_n260  &  n_n283  &  n_n285 ) ;
 assign n_n2618 = ( n_n2  &  n_n60 ) | ( n_n1  &  wire118 ) ;
 assign wire944 = ( n_n151 ) | ( wire75 ) | ( n_n206 ) | ( wire72 ) ;
 assign n_n5769 = ( i_7_  &  (~ i_6_)  &  n_n165  &  n_n284 ) ;
 assign n_n127 = ( n_n283  &  n_n165  &  n_n284 ) ;
 assign n_n4982 = ( wire5140 ) | ( wire19834 ) | ( wire19835 ) ;
 assign wire48 = ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n242  &  n_n281 ) ;
 assign n_n265 = ( n_n266  &  n_n285  &  n_n284 ) ;
 assign n_n268 = ( n_n271  &  n_n285  &  n_n284 ) ;
 assign n_n2550 = ( n_n268  &  wire273 ) | ( n_n268  &  wire1326 ) ;
 assign n_n2545 = ( wire5115 ) | ( wire5116 ) | ( wire19849 ) ;
 assign wire268 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire782 = ( n_n265  &  wire200 ) | ( n_n265  &  wire112 ) ;
 assign n_n5796 = ( i_4_  &  n_n155  &  n_n165  &  wire19290 ) ;
 assign n_n4808 = ( n_n5  &  wire75 ) | ( n_n5  &  n_n281  &  wire913 ) ;
 assign n_n4809 = ( n_n5  &  n_n206 ) | ( n_n6  &  wire72 ) ;
 assign n_n4719 = ( n_n4728 ) | ( n_n4729 ) | ( wire19890 ) ;
 assign n_n4718 = ( n_n4723 ) | ( n_n4725 ) | ( wire19980 ) | ( wire19981 ) ;
 assign n_n264 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n153 = ( i_7_  &  i_6_ ) ;
 assign n_n120 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n2772 = ( wire4935 ) | ( wire5453 ) | ( wire19613 ) | ( wire19614 ) ;
 assign n_n130 = ( n_n229  &  n_n165  &  n_n230 ) ;
 assign n_n110 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign n_n121 = ( n_n264  &  n_n165  &  n_n271 ) ;
 assign n_n4705 = ( wire20007 ) | ( n_n124  &  wire1686 ) | ( n_n132  &  wire1686 ) ;
 assign n_n4704 = ( wire20008 ) | ( n_n152  &  wire266 ) | ( n_n152  &  wire1705 ) ;
 assign wire949 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire948 = ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign n_n5224 = ( n_n4416 ) | ( n_n4418 ) | ( wire20033 ) | ( wire20034 ) ;
 assign n_n4534 = ( n_n4548 ) | ( n_n4549 ) | ( wire20129 ) ;
 assign n_n4533 = ( n_n4545 ) | ( n_n4544 ) | ( wire20147 ) ;
 assign n_n4532 = ( n_n4542 ) | ( n_n4541 ) | ( wire20166 ) ;
 assign n_n4531 = ( n_n3173 ) | ( n_n4539 ) | ( wire4679 ) | ( wire20184 ) ;
 assign n_n4530 = ( n_n4536 ) | ( n_n4556 ) | ( n_n4535 ) | ( wire20240 ) ;
 assign n_n3892 = ( n_n3900 ) | ( n_n3899 ) | ( n_n3901 ) ;
 assign n_n4141 = ( n_n3918 ) | ( n_n3919 ) | ( wire20353 ) ;
 assign n_n4015 = ( n_n4  &  wire95 ) | ( n_n4  &  n_n228  &  wire912 ) ;
 assign n_n4 = ( n_n208  &  n_n285  &  n_n284 ) ;
 assign n_n2789 = ( n_n2792 ) | ( n_n2793 ) | ( wire20571 ) ;
 assign n_n2795 = ( n_n2852 ) | ( wire20610 ) | ( wire20611 ) | ( wire20614 ) ;
 assign n_n2840 = ( n_n3727 ) | ( wire4264 ) | ( n_n4  &  n_n9 ) ;
 assign n_n2839 = ( wire4259 ) | ( wire20616 ) | ( wire20617 ) ;
 assign n_n128 = ( n_n165  &  n_n230  &  n_n271 ) ;
 assign n_n5682 = ( (~ i_7_)  &  (~ i_6_)  &  n_n230  &  n_n116 ) ;
 assign n_n5676 = ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n116 ) ;
 assign n_n4512 = ( wire20629 ) | ( wire20630 ) ;
 assign n_n4508 = ( wire826 ) | ( wire4234 ) | ( wire4235 ) | ( wire4236 ) ;
 assign wire216 = ( wire911  &  n_n281 ) | ( n_n281  &  wire912 ) ;
 assign n_n255 = ( n_n260  &  n_n271  &  n_n285 ) ;
 assign n_n4186 = ( wire372 ) | ( wire894 ) | ( wire20651 ) | ( wire20652 ) ;
 assign wire392 = ( n_n255  &  n_n54 ) | ( n_n241  &  n_n105 ) ;
 assign wire559 = ( n_n241  &  n_n216 ) | ( n_n177  &  n_n45 ) ;
 assign wire950 = ( wire902  &  n_n258 ) | ( n_n258  &  wire912 ) ;
 assign n_n5247 = ( wire590 ) | ( n_n5005 ) | ( wire19306 ) | ( wire20662 ) ;
 assign wire926 = ( i_2_  &  (~ i_0_) ) ;
 assign n_n5797 = ( i_4_  &  n_n153  &  n_n165  &  wire19290 ) ;
 assign wire503 = ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n165 ) ;
 assign n_n4197 = ( wire19753 ) | ( wire19754 ) | ( wire19758 ) | ( wire20691 ) ;
 assign n_n4194 = ( n_n4219 ) | ( n_n4199 ) | ( wire20718 ) | ( wire20743 ) ;
 assign n_n5235 = ( n_n3361 ) | ( n_n3360 ) | ( wire20913 ) | ( wire20914 ) ;
 assign n_n163 = ( (~ i_9_)  &  (~ i_10_) ) ;
 assign n_n5693 = ( n_n163  &  n_n273  &  n_n165  &  wire19294 ) ;
 assign wire452 = ( n_n274  &  n_n283  &  n_n165  &  wire19294 ) ;
 assign wire758 = ( n_n274  &  n_n283  &  n_n165  &  wire19296 ) ;
 assign wire923 = ( i_9_  &  (~ i_10_) ) ;
 assign n_n132 = ( n_n283  &  n_n165  &  n_n230 ) ;
 assign n_n3140 = ( n_n4015 ) | ( wire20925 ) | ( wire20926 ) ;
 assign n_n7424 = ( n_n4  &  n_n228  &  wire902 ) ;
 assign n_n3 = ( n_n229  &  n_n285  &  n_n284 ) ;
 assign n_n3727 = ( n_n4  &  n_n60 ) | ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) ;
 assign n_n3138 = ( n_n4005 ) | ( wire446 ) | ( wire20946 ) | ( wire20947 ) ;
 assign n_n3089 = ( n_n3092 ) | ( n_n3093 ) | ( wire21131 ) ;
 assign n_n3094 = ( n_n3107 ) | ( n_n3108 ) | ( wire21148 ) ;
 assign n_n152 = ( n_n260  &  n_n283  &  n_n165 ) ;
 assign n_n111 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign n_n133 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign n_n3898 = ( n_n3918 ) | ( n_n3919 ) | ( wire21186 ) ;
 assign n_n3890 = ( n_n3895 ) | ( wire21220 ) | ( wire21221 ) | ( wire21245 ) ;
 assign n_n3897 = ( n_n3914 ) | ( n_n3915 ) | ( wire21264 ) ;
 assign n_n3896 = ( n_n3913 ) | ( wire3626 ) | ( wire21276 ) | ( wire21290 ) ;
 assign n_n57 = ( n_n266  &  n_n230  &  n_n285 ) ;
 assign n_n56 = ( n_n230  &  n_n271  &  n_n285 ) ;
 assign n_n2440 = ( wire4059 ) | ( wire4060 ) | ( n_n56  &  n_n226 ) ;
 assign wire955 = ( n_n257 ) | ( wire208 ) | ( wire72 ) | ( wire199 ) ;
 assign n_n2060 = ( n_n2073 ) | ( n_n2108 ) | ( wire3510 ) | ( wire21396 ) ;
 assign n_n145 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign n_n2062 = ( n_n2079 ) | ( wire3489 ) | ( wire3490 ) | ( wire21440 ) ;
 assign n_n2058 = ( n_n2067 ) | ( wire21507 ) | ( wire21508 ) | ( wire21514 ) ;
 assign n_n2063 = ( n_n2081 ) | ( n_n2080 ) | ( wire21557 ) ;
 assign n_n2064 = ( n_n2085 ) | ( n_n2083 ) | ( wire21588 ) ;
 assign n_n2065 = ( n_n2088 ) | ( n_n2086 ) | ( wire21612 ) ;
 assign wire169 = ( i_8_  &  n_n231  &  n_n285  &  n_n284 ) | ( (~ i_8_)  &  n_n231  &  n_n285  &  n_n284 ) ;
 assign n_n126 = ( n_n273  &  n_n165  &  n_n284 ) ;
 assign n_n5660 = ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n284 ) ;
 assign n_n5659 = ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n284 ) ;
 assign n_n1670 = ( wire3241 ) | ( n_n127  &  wire299 ) | ( n_n127  &  wire21624 ) ;
 assign wire581 = ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n284  &  n_n116 ) ;
 assign wire880 = ( i_7_  &  i_6_  &  n_n284  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n116 ) ;
 assign n_n1729 = ( wire21635 ) | ( n_n3  &  wire1732 ) ;
 assign n_n1679 = ( n_n1680 ) | ( n_n1689 ) | ( n_n1692 ) | ( wire21881 ) ;
 assign n_n1694 = ( wire2912 ) | ( wire2913 ) | ( wire21885 ) ;
 assign n_n1693 = ( n_n1724 ) | ( wire2901 ) | ( wire2902 ) | ( wire21896 ) ;
 assign wire957 = ( n_n37 ) | ( n_n83 ) | ( wire154 ) | ( wire64 ) ;
 assign n_n1089 = ( n_n1111 ) | ( wire2808 ) | ( wire21999 ) | ( wire22014 ) ;
 assign n_n240 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign n_n380 = ( wire22360 ) | ( wire22361 ) | ( n_n246  &  wire1345 ) ;
 assign n_n381 = ( n_n3  &  wire1347 ) | ( n_n4  &  wire1346 ) ;
 assign n_n333 = ( n_n340 ) | ( n_n339 ) | ( wire22587 ) | ( wire22588 ) ;
 assign n_n746 = ( wire2163 ) | ( wire2168 ) | ( wire2169 ) | ( wire22602 ) ;
 assign n_n731 = ( n_n741 ) | ( n_n740 ) | ( n_n732 ) | ( wire22827 ) ;
 assign n_n745 = ( n_n775 ) | ( wire22839 ) | ( n_n4  &  wire1837 ) ;
 assign wire126 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign n_n189 = ( n_n283  &  n_n230  &  n_n285 ) ;
 assign n_n5053 = ( n_n189  &  wire6004 ) | ( n_n189  &  wire19279 ) | ( n_n189  &  wire19280 ) ;
 assign n_n241 = ( n_n266  &  n_n260  &  n_n285 ) ;
 assign n_n5061 = ( n_n241  &  wire5936 ) | ( n_n241  &  wire19191 ) | ( n_n241  &  wire19192 ) ;
 assign n_n5062 = ( n_n255  &  wire5931 ) | ( n_n255  &  wire19194 ) | ( n_n255  &  wire19195 ) ;
 assign n_n5020 = ( n_n5061 ) | ( n_n5062 ) | ( wire5922 ) | ( wire5923 ) ;
 assign n_n99 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign n_n54 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign n_n186 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire863 = ( n_n57  &  n_n222  &  wire898 ) | ( n_n57  &  wire898  &  n_n258 ) ;
 assign n_n4970 = ( n_n57  &  n_n99 ) | ( n_n57  &  n_n54 ) | ( n_n57  &  n_n186 ) ;
 assign wire153 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign wire200 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n4926 = ( n_n56  &  wire88 ) | ( n_n56  &  n_n222  &  wire908 ) ;
 assign n_n4315 = ( wire5340 ) | ( wire5341 ) | ( wire5343 ) | ( wire5344 ) ;
 assign n_n6 = ( n_n230  &  n_n261  &  n_n285 ) ;
 assign n_n5 = ( n_n230  &  n_n263  &  n_n285 ) ;
 assign n_n4826 = ( n_n5  &  n_n108 ) | ( n_n6  &  wire70 ) ;
 assign n_n4828 = ( n_n5  &  wire66 ) | ( n_n5  &  wire899  &  n_n256 ) ;
 assign n_n4823 = ( n_n6  &  wire73 ) | ( n_n6  &  wire900  &  n_n228 ) ;
 assign wire90 = ( wire19738 ) | ( wire913  &  n_n256 ) ;
 assign wire584 = ( n_n6  &  wire44 ) | ( n_n5  &  n_n65 ) ;
 assign wire976 = ( n_n12 ) | ( n_n70 ) | ( wire79 ) | ( wire73 ) ;
 assign n_n4204 = ( wire5268 ) | ( wire5269 ) | ( wire19741 ) | ( wire19742 ) ;
 assign n_n4815 = ( n_n6  &  wire63 ) | ( n_n6  &  n_n228  &  wire902 ) ;
 assign n_n4821 = ( n_n5  &  wire44 ) | ( n_n6  &  n_n11 ) ;
 assign n_n4814 = ( n_n6  &  n_n60 ) | ( n_n5  &  wire137 ) ;
 assign n_n4816 = ( n_n5  &  wire95 ) | ( n_n5  &  n_n281  &  wire914 ) ;
 assign wire573 = ( n_n6  &  n_n12 ) | ( n_n5  &  wire70 ) ;
 assign wire60 = ( i_15_  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n258 ) ;
 assign n_n4834 = ( n_n110  &  n_n5 ) | ( n_n6  &  wire60 ) ;
 assign n_n4961 = ( wire166  &  n_n266  &  n_n230  &  n_n285 ) ;
 assign n_n4966 = ( wire224  &  n_n230  &  n_n271  &  n_n285 ) ;
 assign n_n4967 = ( n_n57  &  n_n95 ) | ( n_n57  &  n_n49 ) | ( n_n57  &  n_n96 ) ;
 assign wire613 = ( n_n56  &  wire153 ) | ( n_n57  &  wire224 ) ;
 assign wire614 = ( n_n57  &  wire99 ) | ( n_n57  &  wire41 ) ;
 assign n_n4251 = ( wire4761 ) | ( wire5033 ) | ( n_n56  &  wire118 ) ;
 assign n_n4287 = ( n_n5796 ) | ( n_n56  &  wire72 ) ;
 assign wire99 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire389 = ( n_n6  &  n_n220  &  wire904 ) | ( n_n6  &  n_n256  &  wire904 ) ;
 assign wire708 = ( n_n5  &  wire224 ) | ( n_n6  &  n_n96 ) ;
 assign n_n4211 = ( n_n4251 ) | ( wire708 ) | ( wire4196 ) | ( wire20675 ) ;
 assign wire166 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire224 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire617 = ( n_n6  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign wire673 = ( n_n5  &  wire254 ) | ( n_n5  &  wire41 ) ;
 assign wire674 = ( wire153  &  n_n5 ) | ( n_n5  &  wire180 ) ;
 assign n_n4210 = ( wire673 ) | ( wire674 ) | ( wire20677 ) | ( wire20678 ) ;
 assign n_n4892 = ( n_n56  &  wire63 ) | ( n_n56  &  n_n228  &  wire902 ) ;
 assign n_n4898 = ( n_n56  &  n_n11 ) | ( n_n57  &  wire113 ) ;
 assign n_n4895 = ( n_n57  &  n_n60 ) | ( n_n56  &  wire137 ) ;
 assign wire488 = ( wire5035 ) | ( n_n56  &  wire132 ) ;
 assign wire878 = ( wire5031 ) | ( n_n56  &  n_n60 ) | ( n_n56  &  n_n206 ) ;
 assign n_n48 = ( n_n264  &  n_n283  &  n_n285 ) ;
 assign wire51 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign n_n4179 = ( n_n48  &  wire51 ) | ( n_n53  &  n_n105 ) ;
 assign n_n53 = ( n_n264  &  n_n273  &  n_n285 ) ;
 assign wire40 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign n_n4168 = ( n_n53  &  wire40 ) | ( n_n48  &  n_n31 ) ;
 assign n_n197 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign n_n37 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign wire89 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n228  &  n_n282 ) ;
 assign n_n4094 = ( n_n53  &  wire89 ) | ( n_n53  &  wire901  &  n_n222 ) ;
 assign n_n105 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign n_n47 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign n_n108 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire67 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign n_n4174 = ( n_n53  &  wire67 ) | ( n_n48  &  n_n104 ) ;
 assign wire407 = ( n_n264  &  n_n261  &  n_n282  &  n_n285 ) ;
 assign wire457 = ( n_n264  &  n_n247  &  n_n263  &  n_n285 ) ;
 assign n_n4153 = ( wire407 ) | ( wire457 ) | ( n_n53  &  n_n104 ) ;
 assign n_n4154 = ( n_n48  &  wire72 ) | ( n_n48  &  n_n258  &  wire905 ) ;
 assign wire456 = ( n_n53  &  n_n220  &  wire905 ) | ( n_n53  &  wire905  &  n_n256 ) ;
 assign n_n3964 = ( wire4593 ) | ( wire20257 ) | ( wire20385 ) ;
 assign n_n896 = ( n_n4  &  n_n47 ) | ( n_n4  &  n_n93 ) | ( n_n4  &  n_n46 ) ;
 assign n_n95 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n76 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign wire460 = ( n_n57  &  n_n29 ) | ( n_n57  &  wire49 ) | ( n_n57  &  wire88 ) ;
 assign wire160 = ( i_15_  &  n_n247  &  n_n228 ) | ( (~ i_15_)  &  n_n247  &  n_n258 ) ;
 assign wire409 = ( n_n3  &  n_n252 ) | ( n_n3  &  wire898  &  n_n220 ) ;
 assign n_n4920 = ( n_n57  &  wire79 ) | ( n_n57  &  wire905  &  n_n256 ) ;
 assign n_n4907 = ( n_n56  &  n_n108 ) | ( n_n57  &  wire70 ) ;
 assign wire44 = ( (~ i_15_)  &  n_n253  &  n_n281 ) | ( i_15_  &  n_n253  &  n_n220 ) ;
 assign wire82 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign wire635 = ( n_n56  &  wire44 ) | ( n_n56  &  n_n252 ) | ( n_n56  &  n_n15 ) ;
 assign wire636 = ( n_n56  &  wire42 ) | ( n_n56  &  n_n279  &  wire899 ) ;
 assign n_n3129 = ( wire636 ) | ( wire21065 ) | ( wire21069 ) | ( wire21070 ) ;
 assign n_n11 = ( i_14_  &  i_13_  &  i_12_  &  wire912 ) ;
 assign wire539 = ( n_n5  &  n_n281  &  wire904 ) ;
 assign wire639 = ( n_n5  &  wire70 ) | ( n_n5  &  wire898  &  n_n220 ) ;
 assign n_n3172 = ( wire639 ) | ( wire3904 ) | ( wire20950 ) ;
 assign n_n4605 = ( n_n6  &  wire72 ) | ( n_n6  &  n_n258  &  wire905 ) ;
 assign n_n3118 = ( n_n3172 ) | ( wire20955 ) | ( wire20956 ) ;
 assign wire640 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) | ( n_n4  &  wire80 ) ;
 assign wire867 = ( n_n4  &  n_n31 ) | ( n_n4  &  n_n80 ) | ( n_n4  &  wire1959 ) ;
 assign n_n3107 = ( wire867 ) | ( wire3758 ) | ( wire21136 ) ;
 assign n_n3259 = ( n_n1  &  wire453 ) | ( n_n1  &  n_n256  &  wire914 ) ;
 assign n_n3260 = ( n_n1  &  wire245 ) | ( n_n1  &  wire912  &  n_n225 ) ;
 assign n_n3772 = ( n_n1  &  wire61 ) | ( n_n1  &  n_n279  &  wire908 ) ;
 assign n_n3257 = ( n_n2  &  wire245 ) | ( n_n2  &  wire912  &  n_n225 ) ;
 assign n_n3113 = ( n_n3257 ) | ( wire3889 ) | ( wire20959 ) | ( wire20962 ) ;
 assign n_n2860 = ( n_n1  &  n_n223 ) | ( n_n1  &  wire42 ) | ( n_n1  &  wire1923 ) ;
 assign n_n3255 = ( n_n2  &  n_n76 ) | ( n_n1  &  wire82 ) ;
 assign wire814 = ( n_n1  &  n_n76 ) | ( n_n1  &  n_n26 ) | ( n_n1  &  wire80 ) ;
 assign n_n3112 = ( n_n2860 ) | ( wire814 ) | ( wire3884 ) | ( wire20964 ) ;
 assign n_n3162 = ( n_n1  &  n_n49 ) | ( n_n1  &  wire71 ) | ( n_n1  &  wire1877 ) ;
 assign wire68 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign wire496 = ( n_n2  &  n_n95 ) | ( n_n2  &  n_n49 ) | ( n_n2  &  wire71 ) ;
 assign wire806 = ( n_n1  &  n_n179 ) | ( n_n1  &  wire55 ) | ( n_n1  &  wire57 ) ;
 assign n_n3096 = ( n_n3113 ) | ( n_n3112 ) | ( wire20971 ) ;
 assign n_n31 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign n_n10 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign n_n100 = ( n_n260  &  n_n261  &  n_n285 ) ;
 assign n_n1359 = ( n_n4  &  wire19578 ) | ( n_n4  &  n_n222  &  wire906 ) ;
 assign n_n3525 = ( n_n1  &  wire84 ) | ( n_n1  &  n_n279  &  wire913 ) ;
 assign n_n107 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire983 = ( wire48 ) | ( wire62 ) | ( n_n204 ) | ( n_n16 ) ;
 assign n_n2136 = ( wire3358 ) | ( n_n6  &  wire983 ) ;
 assign n_n4671 = ( n_n57  &  wire453 ) | ( n_n57  &  n_n256  &  wire914 ) ;
 assign wire252 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) ;
 assign wire329 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) ;
 assign n_n2169 = ( n_n4671 ) | ( wire21442 ) | ( wire21443 ) ;
 assign n_n12 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign n_n66 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire164 = ( i_8_  &  n_n272  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n272  &  n_n230  &  n_n285 ) ;
 assign n_n60 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire985 = ( n_n281  &  wire903 ) | ( n_n281  &  wire914 ) ;
 assign n_n2081 = ( n_n2136 ) | ( wire3354 ) | ( wire21529 ) | ( wire21533 ) ;
 assign wire333 = ( n_n4  &  n_n220  &  wire905 ) | ( n_n4  &  wire905  &  n_n256 ) ;
 assign n_n2101 = ( wire333 ) | ( wire3541 ) | ( wire3542 ) ;
 assign wire988 = ( wire40 ) | ( n_n171 ) | ( n_n74 ) | ( wire21367 ) ;
 assign n_n147 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire912 ) ;
 assign n_n94 = ( n_n260  &  n_n263  &  n_n285 ) ;
 assign n_n280 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n32 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign n_n80 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign wire62 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign n_n4165 = ( n_n48  &  wire62 ) | ( n_n53  &  n_n216 ) ;
 assign n_n42 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign wire81 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign n_n1506 = ( n_n5  &  n_n42 ) | ( n_n6  &  wire81 ) ;
 assign wire69 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign n_n4624 = ( n_n6  &  n_n197 ) | ( n_n5  &  wire69 ) ;
 assign n_n1412 = ( n_n2  &  n_n32 ) | ( n_n1  &  wire85 ) ;
 assign wire990 = ( wire67 ) | ( n_n135 ) | ( n_n41 ) | ( wire347 ) ;
 assign wire664 = ( n_n3  &  wire911  &  n_n258 ) ;
 assign wire992 = ( wire60 ) | ( n_n18 ) | ( wire123 ) | ( wire100 ) ;
 assign n_n4858 = ( n_n111  &  n_n5 ) | ( n_n6  &  wire49 ) ;
 assign n_n4864 = ( n_n6  &  wire64 ) | ( n_n6  &  n_n279  &  wire907 ) ;
 assign n_n4635 = ( n_n5  &  wire102 ) | ( n_n5  &  n_n279  &  wire914 ) ;
 assign n_n1129 = ( n_n4858 ) | ( n_n4864 ) | ( wire2704 ) | ( wire22106 ) ;
 assign n_n6582 = ( n_n6  &  n_n256  &  wire914 ) ;
 assign n_n4870 = ( n_n111  &  n_n6 ) | ( n_n5  &  wire85 ) ;
 assign n_n1497 = ( n_n6  &  n_n104 ) | ( n_n5  &  wire78 ) ;
 assign n_n1130 = ( wire2698 ) | ( wire2699 ) | ( wire22112 ) ;
 assign n_n4846 = ( n_n6  &  n_n22 ) | ( n_n5  &  wire49 ) ;
 assign n_n4852 = ( n_n5  &  wire19407 ) | ( n_n5  &  n_n256  &  wire897 ) ;
 assign n_n1490 = ( n_n6  &  wire69 ) | ( n_n5  &  n_n103 ) ;
 assign wire998 = ( wire40 ) | ( n_n74 ) | ( wire140 ) | ( wire346 ) ;
 assign n_n1095 = ( n_n1129 ) | ( n_n1130 ) | ( wire22119 ) ;
 assign n_n1132 = ( n_n1240 ) | ( wire22129 ) | ( wire22130 ) ;
 assign n_n1133 = ( n_n1242 ) | ( n_n1243 ) | ( wire22142 ) ;
 assign n_n1505 = ( n_n54  &  n_n5 ) | ( n_n6  &  wire51 ) ;
 assign n_n1096 = ( n_n1132 ) | ( n_n1133 ) | ( wire22148 ) | ( wire22149 ) ;
 assign n_n1542 = ( n_n48  &  n_n22 ) | ( n_n53  &  wire56 ) ;
 assign n_n3827 = ( n_n48  &  wire61 ) | ( n_n48  &  n_n279  &  wire908 ) ;
 assign n_n1135 = ( n_n4165 ) | ( n_n1536 ) | ( wire22157 ) | ( wire22159 ) ;
 assign n_n1097 = ( n_n1135 ) | ( wire2638 ) | ( wire22169 ) | ( wire22176 ) ;
 assign n_n9 = ( i_14_  &  i_13_  &  i_12_  &  wire902 ) ;
 assign n_n65 = ( i_14_  &  i_13_  &  i_12_  &  wire900 ) ;
 assign wire368 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n247  &  n_n228 ) ;
 assign n_n1066 = ( n_n94  &  wire368 ) | ( n_n94  &  n_n88 ) ;
 assign wire114 = ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign wire120 = ( i_15_  &  n_n275  &  n_n225 ) | ( (~ i_15_)  &  n_n275  &  n_n225 ) ;
 assign wire459 = ( n_n31  &  n_n94 ) | ( n_n94  &  n_n80 ) | ( n_n94  &  wire88 ) ;
 assign n_n855 = ( wire459 ) | ( wire22648 ) | ( n_n94  &  wire114 ) ;
 assign n_n3870 = ( n_n100  &  wire19457 ) | ( n_n100  &  n_n222  &  wire897 ) ;
 assign wire881 = ( n_n100  &  wire902  &  n_n258 ) ;
 assign n_n772 = ( n_n855 ) | ( wire2091 ) | ( wire2092 ) | ( wire22654 ) ;
 assign wire301 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n282 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n282 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n282 ) ;
 assign wire461 = ( n_n48  &  n_n88 ) | ( n_n48  &  n_n258  &  wire912 ) ;
 assign n_n824 = ( wire461 ) | ( wire2008 ) | ( n_n53  &  wire301 ) ;
 assign wire670 = ( n_n6  &  n_n105 ) | ( n_n6  &  n_n46 ) | ( n_n6  &  wire19577 ) ;
 assign n_n761 = ( n_n824 ) | ( wire2001 ) | ( wire2002 ) | ( wire22722 ) ;
 assign n_n275 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign n_n266 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign wire916 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_)  &  n_n284 ) ;
 assign n_n260 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n269 = ( i_9_  &  i_10_ ) ;
 assign n_n253 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign n_n229 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n227 = ( n_n229  &  n_n230  &  n_n285 ) ;
 assign n_n254 = ( i_13_  &  i_12_ ) ;
 assign n_n274 = ( (~ i_9_)  &  i_10_ ) ;
 assign n_n242 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign n_n208 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n207 = ( n_n208  &  n_n230  &  n_n285 ) ;
 assign n_n279 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire911 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n204 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign n_n273 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign n_n177 = ( n_n273  &  n_n230  &  n_n285 ) ;
 assign wire901 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n84 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n222 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign n_n283 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n247 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n155 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n165 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n142 = ( n_n260  &  n_n273  &  n_n165 ) ;
 assign wire899 = ( i_9_  &  i_10_  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n223 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign n_n136 = ( n_n260  &  n_n208  &  n_n165 ) ;
 assign n_n281 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire913 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign wire896 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  n_n230 ) ;
 assign n_n230 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n261 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign n_n278 = ( i_13_  &  (~ i_12_) ) ;
 assign n_n259 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign n_n149 = ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign n_n271 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n122 = ( n_n264  &  n_n229  &  n_n165 ) ;
 assign n_n112 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign wire900 = ( (~ i_9_)  &  i_10_  &  i_11_  &  i_15_ ) ;
 assign n_n93 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire898 = ( i_9_  &  i_10_  &  i_11_  &  i_15_ ) ;
 assign n_n228 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign wire903 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  (~ i_15_) ) ;
 assign n_n212 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) ;
 assign wire902 = ( i_9_  &  (~ i_10_)  &  i_11_  &  i_15_ ) ;
 assign n_n30 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n221 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign n_n258 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n216 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign n_n220 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign wire912 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  i_15_ ) ;
 assign n_n7 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n144 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign wire905 = ( i_9_  &  i_10_  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign n_n257 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign n_n50 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign n_n267 = ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign wire906 = ( (~ i_9_)  &  i_10_  &  i_11_  &  (~ i_15_) ) ;
 assign n_n46 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) ;
 assign n_n256 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n89 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign wire914 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign n_n87 = ( i_14_  &  i_13_  &  i_12_  &  wire914 ) ;
 assign n_n282 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n34 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign n_n225 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign n_n270 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign n_n28 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) ;
 assign wire897 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  i_15_ ) ;
 assign n_n75 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) ;
 assign n_n171 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign n_n21 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) ;
 assign n_n17 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign n_n246 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign n_n236 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire903 ) ;
 assign wire908 = ( i_9_  &  (~ i_10_)  &  i_11_  &  (~ i_15_) ) ;
 assign n_n40 = ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire904 = ( i_9_  &  i_10_  &  i_11_  &  (~ i_15_) ) ;
 assign n_n102 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign n_n263 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire907 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  (~ i_15_) ) ;
 assign n_n33 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire907 ) ;
 assign n_n135 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign n_n78 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign n_n200 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n29 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign n_n64 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire900 ) ;
 assign n_n150 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire911 ) ;
 assign n_n25 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign n_n70 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) ;
 assign n_n24 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign n_n27 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n20 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) ;
 assign n_n97 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign n_n45 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign n_n52 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n41 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign n_n26 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) ;
 assign n_n23 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) ;
 assign n_n74 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign n_n71 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) ;
 assign n_n69 = ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign n_n14 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire898 ) ;
 assign n_n252 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign n_n63 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) ;
 assign n_n8 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign n_n199 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign n_n18 = ( i_14_  &  i_13_  &  i_12_  &  wire913 ) ;
 assign n_n88 = ( i_15_  &  n_n222  &  n_n247 ) ;
 assign n_n92 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign n_n98 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) ;
 assign n_n179 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign n_n104 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign n_n38 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) ;
 assign n_n109 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire1011 = ( wire19206 ) | ( n_n283  &  wire384 ) | ( n_n283  &  wire19205 ) ;
 assign n_n5030 = ( n_n124  &  n_n223 ) | ( n_n124  &  wire19239 ) | ( n_n124  &  wire19316 ) ;
 assign n_n5063 = ( wire5910 ) | ( n_n255  &  wire19207 ) | ( n_n255  &  wire19208 ) ;
 assign wire927 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n116 ) ;
 assign wire254 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire165 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n4936 = ( n_n266  &  n_n230  &  wire165  &  n_n285 ) ;
 assign n_n6678 = ( n_n6  &  wire905  &  n_n256 ) ;
 assign wire79 = ( i_15_  &  n_n281  &  n_n259 ) | ( (~ i_15_)  &  n_n259  &  n_n225 ) ;
 assign n_n4839 = ( n_n6  &  wire79 ) | ( n_n6  &  wire905  &  n_n256 ) ;
 assign n_n4842 = ( n_n5  &  n_n76 ) | ( n_n6  &  wire82 ) ;
 assign wire1016 = ( n_n223 ) | ( n_n171 ) | ( wire42 ) | ( wire53 ) ;
 assign n_n4960 = ( n_n266  &  n_n230  &  n_n285  &  wire180 ) ;
 assign n_n4954 = ( n_n57  &  wire55 ) | ( n_n57  &  n_n279  &  wire912 ) ;
 assign n_n4953 = ( n_n57  &  wire57 ) | ( n_n57  &  n_n279  &  wire914 ) ;
 assign n_n4955 = ( n_n56  &  n_n95 ) | ( n_n56  &  n_n49 ) | ( n_n56  &  n_n96 ) ;
 assign wire671 = ( n_n56  &  wire99 ) | ( n_n56  &  wire41 ) ;
 assign n_n4219 = ( wire20705 ) | ( wire20706 ) | ( wire20710 ) ;
 assign n_n226 = ( i_14_  &  i_13_  &  i_12_  &  wire899 ) ;
 assign n_n61 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire908 ) ;
 assign wire469 = ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n259  &  n_n228 ) ;
 assign n_n4073 = ( n_n53  &  wire469 ) | ( n_n53  &  n_n222  &  wire899 ) ;
 assign wire475 = ( n_n53  &  n_n144 ) | ( n_n53  &  n_n281  &  wire905 ) ;
 assign n_n4068 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n9 ) | ( n_n53  &  n_n144 ) ;
 assign n_n4069 = ( n_n53  &  n_n60 ) | ( n_n53  &  n_n8 ) | ( n_n53  &  n_n226 ) ;
 assign wire77 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n1363 = ( n_n3  &  n_n105 ) | ( n_n4  &  wire77 ) ;
 assign wire184 = ( (~ i_15_)  &  n_n247  &  n_n281 ) | ( i_15_  &  n_n247  &  n_n220 ) ;
 assign n_n3324 = ( n_n57  &  n_n9 ) | ( n_n56  &  wire184 ) ;
 assign n_n6504 = ( n_n48  &  n_n258  &  wire912 ) ;
 assign n_n1633 = ( n_n197  &  n_n100 ) | ( n_n94  &  wire69 ) ;
 assign n_n4923 = ( n_n56  &  n_n76 ) | ( n_n57  &  wire82 ) ;
 assign wire385 = ( n_n57  &  wire1856 ) | ( n_n57  &  n_n220  &  wire908 ) ;
 assign n_n3130 = ( wire385 ) | ( wire21073 ) | ( wire21074 ) ;
 assign wire686 = ( n_n94  &  wire912  &  n_n256 ) | ( n_n94  &  wire912  &  n_n225 ) ;
 assign wire825 = ( n_n260  &  n_n263  &  n_n285  &  wire57 ) ;
 assign n_n3167 = ( wire825 ) | ( wire20973 ) | ( wire20974 ) | ( wire20975 ) ;
 assign wire278 = ( i_8_  &  n_n231  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n231  &  n_n230  &  n_n285 ) ;
 assign wire1018 = ( n_n228  &  wire902 ) | ( n_n258  &  wire905 ) ;
 assign n_n3117 = ( n_n3167 ) | ( wire3870 ) | ( wire20984 ) ;
 assign n_n3242 = ( n_n4  &  wire245 ) | ( n_n4  &  wire912  &  n_n225 ) ;
 assign wire557 = ( n_n3  &  n_n95 ) | ( n_n3  &  n_n49 ) | ( n_n3  &  wire71 ) ;
 assign n_n3108 = ( n_n3242 ) | ( wire557 ) | ( wire3754 ) | ( wire3755 ) ;
 assign n_n3757 = ( n_n1  &  wire63 ) | ( n_n1  &  n_n281  &  wire908 ) ;
 assign wire739 = ( n_n2  &  wire899  &  n_n228 ) ;
 assign n_n3110 = ( n_n2550 ) | ( wire3932 ) | ( wire20931 ) ;
 assign n_n2852 = ( n_n4  &  n_n49 ) | ( n_n4  &  wire71 ) | ( n_n4  &  wire20592 ) ;
 assign n_n3109 = ( n_n2852 ) | ( wire20933 ) | ( wire20934 ) | ( wire20936 ) ;
 assign n_n3155 = ( wire20938 ) | ( n_n2  &  wire1932 ) ;
 assign n_n3519 = ( n_n2  &  n_n108 ) | ( n_n1  &  wire70 ) ;
 assign n_n3520 = ( n_n2  &  wire79 ) | ( n_n2  &  wire905  &  n_n256 ) ;
 assign wire1027 = ( wire44 ) | ( n_n11 ) | ( n_n148 ) | ( wire95 ) ;
 assign wire1026 = ( wire160 ) | ( wire44 ) | ( n_n252 ) | ( n_n15 ) ;
 assign n_n81 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign wire470 = ( n_n53  &  n_n33 ) | ( n_n53  &  wire901  &  n_n281 ) ;
 assign n_n3019 = ( n_n53  &  n_n280 ) | ( n_n53  &  n_n33 ) | ( n_n53  &  n_n81 ) ;
 assign n_n2986 = ( n_n4  &  wire79 ) | ( n_n4  &  wire899  &  n_n256 ) ;
 assign n_n3524 = ( n_n1  &  wire19738 ) | ( n_n1  &  wire913  &  n_n256 ) ;
 assign wire93 = ( wire245 ) | ( wire912  &  n_n225 ) ;
 assign wire185 = ( i_8_  &  n_n264  &  n_n155  &  n_n285 ) | ( (~ i_8_)  &  n_n264  &  n_n155  &  n_n285 ) ;
 assign n_n2148 = ( wire3310 ) | ( wire21560 ) | ( wire21561 ) | ( wire21562 ) ;
 assign n_n19 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) ;
 assign n_n2272 = ( n_n53  &  n_n108 ) | ( n_n53  &  n_n70 ) | ( n_n53  &  n_n19 ) ;
 assign n_n2126 = ( n_n2272 ) | ( wire3491 ) | ( wire21417 ) ;
 assign wire135 = ( i_8_  &  n_n260  &  n_n155  &  n_n285 ) | ( (~ i_8_)  &  n_n260  &  n_n155  &  n_n285 ) ;
 assign wire264 = ( i_15_  &  n_n275  &  n_n279 ) | ( (~ i_15_)  &  n_n275  &  n_n279 ) ;
 assign wire1031 = ( n_n281  &  wire905 ) | ( n_n281  &  wire908 ) ;
 assign wire1030 = ( n_n281  &  wire913 ) | ( n_n281  &  wire903 ) ;
 assign wire466 = ( n_n4  &  n_n220  &  wire908 ) | ( n_n4  &  n_n256  &  wire908 ) ;
 assign n_n2104 = ( wire3533 ) | ( wire3534 ) | ( wire21374 ) ;
 assign wire411 = ( n_n6  &  n_n220  &  wire905 ) | ( n_n6  &  wire905  &  n_n256 ) ;
 assign n_n2137 = ( wire411 ) | ( wire3344 ) | ( wire3345 ) ;
 assign n_n2110 = ( wire3528 ) | ( wire21381 ) | ( n_n268  &  wire1484 ) ;
 assign n_n2073 = ( n_n2110 ) | ( wire3521 ) | ( wire21387 ) ;
 assign n_n2108 = ( wire3518 ) | ( wire21390 ) | ( n_n3  &  n_n186 ) ;
 assign wire476 = ( n_n3  &  n_n220  &  wire904 ) | ( n_n3  &  n_n256  &  wire904 ) ;
 assign wire1042 = ( n_n25 ) | ( n_n24 ) | ( wire104 ) | ( wire228 ) ;
 assign n_n1779 = ( wire21842 ) | ( n_n48  &  wire1042 ) ;
 assign n_n58 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign wire667 = ( i_15_  &  n_n94  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n94  &  n_n222  &  n_n247 ) ;
 assign wire696 = ( n_n94  &  wire911  &  n_n281 ) | ( n_n94  &  wire911  &  n_n225 ) ;
 assign n_n1757 = ( wire667 ) | ( wire696 ) | ( wire21686 ) | ( wire21687 ) ;
 assign n_n3581 = ( n_n53  &  wire84 ) | ( n_n53  &  n_n279  &  wire913 ) ;
 assign wire700 = ( n_n207  &  wire913  &  n_n256 ) ;
 assign wire1043 = ( n_n240 ) | ( n_n109 ) | ( wire143 ) | ( wire306 ) ;
 assign n_n1215 = ( wire700 ) | ( wire22079 ) | ( n_n227  &  wire1043 ) ;
 assign n_n1628 = ( n_n94  &  wire514 ) | ( n_n94  &  wire911  &  n_n225 ) ;
 assign n_n2732 = ( n_n100  &  wire52 ) | ( n_n100  &  n_n279  &  wire913 ) ;
 assign n_n1624 = ( n_n197  &  n_n94 ) | ( n_n100  &  wire62 ) ;
 assign wire1044 = ( wire60 ) | ( n_n107 ) | ( wire247 ) | ( wire83 ) ;
 assign n_n1262 = ( n_n53  &  wire68 ) | ( n_n53  &  wire175 ) | ( n_n53  &  wire22257 ) ;
 assign wire75 = ( (~ i_15_)  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n220 ) ;
 assign wire579 = ( n_n264  &  n_n242  &  n_n261  &  n_n285 ) ;
 assign wire764 = ( n_n264  &  n_n259  &  n_n263  &  n_n285 ) ;
 assign n_n1140 = ( n_n1262 ) | ( wire2542 ) | ( wire2543 ) | ( wire22264 ) ;
 assign wire699 = ( n_n6  &  wire66 ) | ( n_n6  &  wire899  &  n_n256 ) ;
 assign n_n1127 = ( n_n4624 ) | ( wire699 ) | ( wire2785 ) | ( wire22020 ) ;
 assign wire1052 = ( wire67 ) | ( n_n135 ) | ( n_n41 ) | ( wire347 ) ;
 assign n_n1320 = ( n_n110  &  n_n4 ) | ( n_n3  &  wire82 ) ;
 assign n_n1240 = ( wire461 ) | ( wire376 ) | ( wire2686 ) | ( wire22121 ) ;
 assign n_n4124 = ( n_n48  &  wire102 ) | ( n_n48  &  n_n279  &  wire914 ) ;
 assign wire629 = ( n_n48  &  n_n281  &  wire912 ) | ( n_n48  &  wire912  &  n_n256 ) ;
 assign wire631 = ( n_n48  &  n_n147 ) | ( n_n53  &  n_n62 ) ;
 assign n_n1242 = ( n_n6879 ) | ( wire679 ) | ( wire2672 ) | ( wire2673 ) ;
 assign n_n1243 = ( wire2665 ) | ( wire22134 ) | ( wire22135 ) | ( wire22136 ) ;
 assign wire223 = ( (~ i_15_)  &  n_n259  &  n_n258 ) | ( i_15_  &  n_n259  &  n_n220 ) ;
 assign wire168 = ( i_8_  &  n_n272  &  n_n260  &  n_n285 ) | ( (~ i_8_)  &  n_n272  &  n_n260  &  n_n285 ) ;
 assign wire1060 = ( n_n221 ) | ( wire469 ) | ( n_n15 ) | ( wire128 ) ;
 assign n_n852 = ( wire22605 ) | ( n_n94  &  wire1060 ) ;
 assign n_n1058 = ( n_n94  &  n_n204 ) | ( n_n94  &  n_n18 ) | ( n_n94  &  n_n203 ) ;
 assign n_n3604 = ( n_n100  &  n_n203 ) | ( n_n100  &  wire20149 ) ;
 assign n_n3610 = ( n_n100  &  wire469 ) | ( n_n100  &  n_n222  &  wire899 ) ;
 assign wire697 = ( n_n94  &  wire911  &  n_n225 ) | ( n_n94  &  wire913  &  n_n225 ) ;
 assign wire1061 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n259  &  n_n225 ) | ( (~ i_15_)  &  n_n259  &  n_n225 ) ;
 assign n_n771 = ( n_n852 ) | ( wire22610 ) | ( wire22611 ) ;
 assign n_n206 = ( i_14_  &  i_13_  &  i_12_  &  wire911 ) ;
 assign wire516 = ( n_n53  &  wire901  &  n_n222 ) | ( n_n53  &  wire901  &  n_n258 ) ;
 assign wire1062 = ( n_n279  &  wire901 ) | ( n_n228  &  wire897 ) ;
 assign n_n825 = ( wire516 ) | ( wire1997 ) | ( wire22725 ) | ( wire22727 ) ;
 assign wire675 = ( n_n48  &  wire898  &  n_n228 ) ;
 assign wire1064 = ( n_n221 ) | ( wire469 ) | ( wire128 ) | ( wire310 ) ;
 assign wire1063 = ( wire901  &  n_n228 ) | ( wire900  &  n_n228 ) ;
 assign n_n762 = ( n_n825 ) | ( wire1990 ) | ( wire22731 ) | ( wire22734 ) ;
 assign n_n13 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign n_n458 = ( wire2436 ) | ( wire2437 ) | ( n_n197  &  n_n94 ) ;
 assign wire1066 = ( n_n258  &  wire914 ) | ( n_n258  &  wire908 ) ;
 assign n_n374 = ( n_n458 ) | ( wire2430 ) | ( wire22372 ) ;
 assign wire486 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n2738 = ( n_n260  &  n_n263  &  n_n285  &  wire140 ) ;
 assign n_n462 = ( wire658 ) | ( n_n707 ) | ( wire2410 ) | ( wire22384 ) ;
 assign wire1069 = ( i_15_  &  n_n258  &  n_n270 ) | ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign n_n346 = ( n_n374 ) | ( wire22382 ) | ( wire22383 ) | ( wire22393 ) ;
 assign n_n203 = ( i_15_  &  n_n242  &  n_n222 ) ;
 assign n_n16 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) ;
 assign n_n285 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n43 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) ;
 assign n_n51 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) ;
 assign n_n82 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) ;
 assign n_n68 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) ;
 assign n_n113 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign n_n86 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) ;
 assign n_n79 = ( i_14_  &  i_13_  &  i_12_  &  wire908 ) ;
 assign n_n103 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) ;
 assign n_n36 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) ;
 assign n_n284 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n44 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) ;
 assign n_n73 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) ;
 assign n_n72 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign n_n85 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) ;
 assign n_n15 = ( i_14_  &  i_13_  &  i_12_  &  wire898 ) ;
 assign wire1071 = ( wire19265 ) | ( wire19266 ) | ( wire19267 ) ;
 assign wire277 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire901 ) ;
 assign n_n4950 = ( n_n230  &  n_n271  &  n_n285  &  wire277 ) ;
 assign n_n4924 = ( n_n56  &  wire80 ) | ( n_n56  &  n_n256  &  wire908 ) ;
 assign wire255 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) ;
 assign n_n4871 = ( n_n230  &  n_n263  &  n_n285  &  wire255 ) ;
 assign n_n4838 = ( n_n5  &  wire60 ) | ( n_n6  &  n_n108 ) ;
 assign wire111 = ( wire42 ) | ( n_n279  &  wire899 ) ;
 assign n_n4730 = ( wire699 ) | ( n_n4838 ) | ( wire5053 ) | ( wire19896 ) ;
 assign wire1076 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign wire1079 = ( n_n264  &  n_n229  &  n_n165 ) | ( n_n264  &  n_n165  &  n_n271 ) ;
 assign n_n6534 = ( n_n6  &  n_n256  &  wire904 ) ;
 assign n_n4330 = ( wire632 ) | ( wire5368 ) | ( wire5369 ) ;
 assign n_n4313 = ( n_n4330 ) | ( wire5361 ) | ( wire5363 ) | ( wire19671 ) ;
 assign wire180 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire70 = ( i_15_  &  n_n253  &  n_n228 ) | ( (~ i_15_)  &  n_n253  &  n_n258 ) ;
 assign wire125 = ( wire66 ) | ( wire899  &  n_n256 ) ;
 assign wire118 = ( i_15_  &  n_n259  &  n_n228 ) | ( (~ i_15_)  &  n_n259  &  n_n258 ) ;
 assign n_n4806 = ( n_n151  &  n_n6 ) | ( n_n5  &  wire118 ) ;
 assign wire709 = ( wire5033 ) | ( n_n56  &  wire118 ) ;
 assign wire372 = ( n_n177  &  n_n200 ) | ( n_n189  &  n_n101 ) ;
 assign wire894 = ( n_n189  &  n_n279  &  wire914 ) ;
 assign wire141 = ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign n_n1341 = ( n_n4  &  wire65 ) | ( n_n4  &  wire902  &  n_n225 ) ;
 assign n_n3974 = ( n_n6504 ) | ( wire470 ) | ( wire376 ) | ( wire4602 ) ;
 assign n_n4090 = ( n_n48  &  wire368 ) | ( n_n48  &  n_n88 ) ;
 assign wire462 = ( n_n48  &  n_n220  &  wire914 ) | ( n_n48  &  n_n256  &  wire914 ) ;
 assign wire464 = ( n_n48  &  n_n85 ) | ( n_n48  &  n_n281  &  wire912 ) ;
 assign n_n3918 = ( n_n3974 ) | ( wire20330 ) | ( wire20331 ) ;
 assign n_n6879 = ( n_n53  &  n_n258  &  wire905 ) ;
 assign wire1089 = ( wire75 ) | ( n_n206 ) | ( wire208 ) | ( wire199 ) ;
 assign n_n3919 = ( n_n4153 ) | ( n_n4154 ) | ( wire20340 ) | ( wire20341 ) ;
 assign n_n3506 = ( n_n4  &  wire42 ) | ( n_n4  &  n_n279  &  wire899 ) ;
 assign wire378 = ( wire4302 ) | ( n_n4  &  wire905  &  n_n256 ) ;
 assign wire455 = ( n_n4  &  n_n222  &  wire900 ) | ( n_n4  &  wire900  &  n_n258 ) ;
 assign wire485 = ( n_n4  &  n_n222  &  wire899 ) | ( n_n4  &  wire899  &  n_n258 ) ;
 assign wire179 = ( wire76 ) | ( n_n279  &  wire900 ) ;
 assign n_n3781 = ( n_n1  &  wire76 ) | ( n_n1  &  n_n279  &  wire900 ) ;
 assign wire676 = ( n_n53  &  n_n226 ) | ( n_n53  &  n_n258  &  wire905 ) ;
 assign n_n3184 = ( n_n4154 ) | ( wire475 ) | ( wire676 ) | ( wire21006 ) ;
 assign wire712 = ( n_n3  &  n_n99 ) | ( n_n3  &  n_n54 ) | ( n_n3  &  wire96 ) ;
 assign n_n3116 = ( wire4472 ) | ( wire20397 ) | ( wire20400 ) | ( wire20987 ) ;
 assign n_n4005 = ( n_n3  &  wire72 ) | ( n_n3  &  n_n258  &  wire905 ) ;
 assign wire446 = ( n_n4  &  n_n144 ) | ( n_n4  &  n_n281  &  wire905 ) ;
 assign n_n35 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign n_n4922 = ( n_n57  &  wire42 ) | ( n_n57  &  n_n279  &  wire899 ) ;
 assign n_n4921 = ( n_n57  &  wire66 ) | ( n_n57  &  wire899  &  n_n256 ) ;
 assign n_n4076 = ( n_n53  &  wire65 ) | ( n_n53  &  wire902  &  n_n225 ) ;
 assign n_n3768 = ( n_n1  &  wire19407 ) | ( n_n1  &  n_n256  &  wire897 ) ;
 assign n_n2467 = ( n_n57  &  n_n99 ) | ( n_n57  &  wire58 ) | ( n_n57  &  wire21296 ) ;
 assign wire386 = ( n_n189  &  n_n102 ) | ( n_n177  &  n_n45 ) ;
 assign wire484 = ( n_n57  &  n_n220  &  wire904 ) | ( n_n57  &  n_n256  &  wire904 ) ;
 assign n_n2439 = ( n_n2467 ) | ( wire3600 ) | ( wire21302 ) | ( wire21303 ) ;
 assign wire1092 = ( n_n66 ) | ( n_n109 ) | ( wire79 ) | ( wire83 ) ;
 assign n_n2149 = ( wire21603 ) | ( n_n48  &  wire1092 ) ;
 assign n_n4912 = ( n_n57  &  wire19738 ) | ( n_n57  &  wire913  &  n_n256 ) ;
 assign n_n4916 = ( n_n56  &  wire19738 ) | ( n_n56  &  wire913  &  n_n256 ) ;
 assign wire327 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) ;
 assign wire1094 = ( i_8_  &  n_n153  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n153  &  n_n230  &  n_n285 ) ;
 assign wire191 = ( i_8_  &  n_n153  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n153  &  n_n230  &  n_n285 ) ;
 assign wire1096 = ( n_n281  &  wire906 ) | ( n_n281  &  wire904 ) ;
 assign wire1095 = ( n_n281  &  wire906 ) | ( n_n281  &  wire914 ) | ( n_n281  &  wire904 ) ;
 assign wire1097 = ( wire167 ) | ( wire210 ) | ( wire235 ) | ( wire399 ) ;
 assign wire1102 = ( wire268 ) | ( wire167 ) | ( wire235 ) | ( wire436 ) ;
 assign wire641 = ( n_n4  &  n_n27 ) | ( n_n4  &  n_n220  &  wire908 ) ;
 assign n_n1756 = ( wire641 ) | ( wire3145 ) | ( wire21690 ) | ( wire21691 ) ;
 assign wire50 = ( (~ i_15_)  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n220 ) ;
 assign wire645 = ( n_n100  &  n_n62 ) | ( n_n100  &  n_n258  &  wire907 ) ;
 assign n_n1286 = ( wire645 ) | ( wire2596 ) | ( wire2597 ) | ( wire22203 ) ;
 assign n_n1148 = ( n_n1286 ) | ( wire2593 ) | ( wire2594 ) ;
 assign n_n1255 = ( wire461 ) | ( wire2516 ) | ( wire22280 ) ;
 assign n_n6848 = ( n_n53  &  wire902  &  n_n258 ) ;
 assign wire479 = ( n_n53  &  n_n220  &  wire908 ) | ( n_n53  &  n_n256  &  wire908 ) ;
 assign wire656 = ( n_n53  &  n_n222  &  wire902 ) | ( n_n53  &  n_n222  &  wire908 ) ;
 assign n_n1137 = ( n_n1255 ) | ( wire22286 ) | ( wire22287 ) ;
 assign n_n62 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign n_n1157 = ( wire2879 ) | ( wire21914 ) | ( wire169  &  n_n10 ) ;
 assign wire1112 = ( n_n58 ) | ( wire75 ) | ( wire223 ) | ( wire63 ) ;
 assign n_n1151 = ( n_n1295 ) | ( n_n1641 ) | ( wire22190 ) | ( wire22193 ) ;
 assign wire1113 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign n_n1102 = ( n_n1151 ) | ( wire22184 ) | ( wire22185 ) | ( wire22201 ) ;
 assign n_n1147 = ( n_n1284 ) | ( wire22219 ) | ( wire22220 ) ;
 assign n_n4675 = ( n_n56  &  wire807 ) | ( n_n56  &  n_n279  &  wire904 ) ;
 assign n_n4681 = ( n_n56  &  n_n42 ) | ( n_n57  &  wire81 ) ;
 assign n_n1604 = ( n_n56  &  n_n54 ) | ( n_n57  &  wire51 ) ;
 assign wire497 = ( n_n56  &  n_n220  &  wire904 ) | ( n_n56  &  n_n256  &  wire904 ) ;
 assign n_n1101 = ( n_n1148 ) | ( n_n1147 ) | ( wire22227 ) | ( wire22228 ) ;
 assign n_n1152 = ( wire798 ) | ( n_n1298 ) | ( wire22236 ) | ( wire22238 ) ;
 assign n_n1154 = ( n_n3615 ) | ( wire874 ) | ( wire2550 ) | ( wire2551 ) ;
 assign n_n3881 = ( wire51  &  n_n100 ) | ( n_n54  &  n_n94 ) ;
 assign wire784 = ( wire166  &  n_n100 ) | ( n_n100  &  wire180 ) ;
 assign n_n1103 = ( n_n1152 ) | ( n_n1154 ) | ( wire22253 ) ;
 assign wire91 = ( wire19457 ) | ( n_n222  &  wire897 ) ;
 assign wire647 = ( n_n6  &  n_n216 ) | ( n_n6  &  n_n203 ) | ( n_n6  &  wire20149 ) ;
 assign wire1119 = ( wire126 ) | ( n_n37 ) | ( wire89 ) | ( wire22783 ) ;
 assign n_n803 = ( wire22785 ) | ( n_n2  &  wire1119 ) ;
 assign wire356 = ( (~ i_14_)  &  i_15_  &  n_n253  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n253  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n253  &  n_n254 ) ;
 assign n_n850 = ( n_n4970 ) | ( wire22613 ) | ( n_n57  &  wire356 ) ;
 assign wire335 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n267 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n267 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n267 ) ;
 assign wire725 = ( n_n100  &  wire899  &  n_n228 ) ;
 assign wire1121 = ( n_n228  &  wire902 ) | ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign wire1120 = ( n_n228  &  wire902 ) | ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign n_n770 = ( n_n850 ) | ( wire2138 ) | ( wire22616 ) | ( wire22620 ) ;
 assign n_n4628 = ( n_n6  &  wire19457 ) | ( n_n6  &  n_n222  &  wire897 ) ;
 assign wire727 = ( n_n5  &  n_n31 ) | ( n_n5  &  n_n80 ) | ( n_n5  &  wire88 ) ;
 assign n_n365 = ( n_n431 ) | ( wire2377 ) | ( wire22409 ) | ( wire22412 ) ;
 assign n_n429 = ( wire2374 ) | ( wire22414 ) | ( wire22415 ) | ( wire22416 ) ;
 assign n_n343 = ( n_n365 ) | ( wire22400 ) | ( wire22401 ) | ( wire22421 ) ;
 assign n_n423 = ( wire2361 ) | ( n_n6  &  wire1645 ) ;
 assign n_n361 = ( wire2355 ) | ( wire2356 ) | ( wire22426 ) ;
 assign n_n363 = ( wire2350 ) | ( wire2353 ) | ( wire2354 ) | ( wire22432 ) ;
 assign n_n342 = ( n_n361 ) | ( n_n363 ) | ( wire22440 ) ;
 assign n_n367 = ( n_n438 ) | ( wire22446 ) | ( wire22447 ) ;
 assign n_n369 = ( n_n443 ) | ( wire2324 ) | ( wire22454 ) | ( wire22457 ) ;
 assign wire809 = ( n_n48  &  wire898  &  n_n258 ) ;
 assign wire1128 = ( wire166 ) | ( n_n113 ) | ( wire57 ) | ( wire22459 ) ;
 assign n_n344 = ( n_n367 ) | ( n_n369 ) | ( wire22463 ) | ( wire22464 ) ;
 assign n_n143 = ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign n_n116 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n39 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) ;
 assign n_n77 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire908 ) ;
 assign n_n67 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign n_n83 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire1130 = ( wire19213 ) | ( n_n275  &  wire1131 ) ;
 assign wire1132 = ( wire5893 ) | ( wire19215 ) | ( wire19216 ) | ( wire19217 ) ;
 assign wire190 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign n_n4941 = ( n_n56  &  wire57 ) | ( n_n56  &  n_n279  &  wire914 ) ;
 assign n_n4942 = ( n_n56  &  wire55 ) | ( n_n56  &  n_n279  &  wire912 ) ;
 assign wire728 = ( n_n56  &  wire157 ) | ( n_n56  &  wire273 ) ;
 assign wire729 = ( n_n57  &  wire277 ) | ( n_n57  &  wire112 ) ;
 assign n_n5685 = ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) ;
 assign n_n4416 = ( wire4889 ) | ( wire20020 ) | ( wire20021 ) ;
 assign n_n4418 = ( wire4882 ) | ( wire20023 ) | ( wire20027 ) ;
 assign wire794 = ( (~ i_7_)  &  i_6_  &  n_n230  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n230  &  n_n116 ) ;
 assign n_n4394 = ( n_n266  &  n_n230  &  n_n285  &  wire247 ) ;
 assign n_n4381 = ( n_n57  &  wire63 ) | ( n_n57  &  n_n281  &  wire908 ) ;
 assign n_n3850 = ( n_n56  &  n_n9 ) | ( n_n57  &  wire132 ) ;
 assign wire473 = ( wire5587 ) | ( n_n57  &  wire137 ) ;
 assign n_n4307 = ( n_n4315 ) | ( wire5336 ) | ( wire19692 ) | ( wire19698 ) ;
 assign wire124 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign n_n4929 = ( n_n266  &  n_n230  &  n_n285  &  wire124 ) ;
 assign wire212 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire250 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire1141 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign n_n4279 = ( n_n4970 ) | ( wire4166 ) | ( wire20712 ) ;
 assign n_n3978 = ( wire4569 ) | ( wire4570 ) | ( wire20273 ) ;
 assign n_n1346 = ( n_n3  &  n_n41 ) | ( n_n4  &  wire78 ) ;
 assign n_n884 = ( n_n4  &  wire88 ) | ( n_n4  &  n_n222  &  wire902 ) ;
 assign n_n3908 = ( n_n884 ) | ( wire3664 ) | ( wire3665 ) | ( wire21228 ) ;
 assign n_n3778 = ( n_n2  &  wire68 ) | ( n_n1  &  n_n42 ) ;
 assign n_n3229 = ( n_n3  &  n_n108 ) | ( n_n4  &  wire70 ) ;
 assign wire740 = ( wire44  &  n_n100 ) | ( n_n100  &  n_n258  &  wire904 ) ;
 assign wire55 = ( i_15_  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n258 ) ;
 assign wire741 = ( n_n48  &  n_n220  &  wire904 ) ;
 assign n_n1555 = ( n_n48  &  n_n95 ) | ( n_n53  &  wire55 ) ;
 assign wire626 = ( n_n53  &  n_n61 ) | ( n_n53  &  wire902  &  n_n220 ) ;
 assign n_n3791 = ( n_n53  &  n_n60 ) | ( n_n53  &  n_n8 ) | ( n_n53  &  n_n61 ) ;
 assign wire591 = ( wire68  &  n_n260  &  n_n273  &  n_n285 ) ;
 assign wire736 = ( n_n4073 ) | ( wire479 ) | ( wire478 ) | ( wire20387 ) ;
 assign n_n2815 = ( n_n3964 ) | ( wire736 ) | ( wire20392 ) ;
 assign n_n2982 = ( n_n4  &  n_n60 ) | ( n_n4  &  n_n8 ) | ( n_n4  &  n_n226 ) ;
 assign wire349 = ( n_n3  &  wire898  &  n_n228 ) ;
 assign wire876 = ( n_n4076 ) | ( wire483 ) | ( n_n4  &  n_n257 ) ;
 assign n_n3097 = ( n_n3116 ) | ( n_n2815 ) | ( wire20996 ) ;
 assign n_n3092 = ( n_n3099 ) | ( n_n3101 ) | ( wire21063 ) ;
 assign n_n3093 = ( n_n3103 ) | ( n_n3104 ) | ( wire21122 ) ;
 assign n_n3173 = ( wire4694 ) | ( wire4695 ) ;
 assign n_n2882 = ( n_n6  &  n_n20 ) | ( n_n6  &  wire79 ) | ( n_n6  &  wire1946 ) ;
 assign n_n3864 = ( n_n100  &  wire63 ) | ( n_n100  &  n_n228  &  wire902 ) ;
 assign wire780 = ( n_n100  &  n_n281  &  wire908 ) ;
 assign n_n2702 = ( n_n106  &  n_n100 ) | ( wire160  &  n_n94 ) ;
 assign wire654 = ( n_n94  &  n_n148 ) | ( n_n94  &  n_n220  &  wire912 ) ;
 assign wire1149 = ( n_n9 ) | ( n_n144 ) | ( wire118 ) | ( wire132 ) ;
 assign n_n2398 = ( n_n94  &  wire1372 ) | ( n_n94  &  wire913  &  n_n220 ) ;
 assign wire1150 = ( wire60 ) | ( n_n204 ) | ( wire247 ) | ( wire210 ) ;
 assign n_n2724 = ( wire160  &  n_n100 ) | ( n_n66  &  n_n94 ) ;
 assign wire1152 = ( n_n66 ) | ( n_n14 ) | ( wire184 ) | ( wire70 ) ;
 assign wire1156 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign n_n2133 = ( wire3340 ) | ( wire21537 ) | ( wire21538 ) ;
 assign wire388 = ( n_n94  &  n_n16 ) | ( n_n94  &  wire911  &  n_n281 ) ;
 assign wire747 = ( wire40  &  n_n94 ) | ( n_n94  &  n_n281  &  wire897 ) ;
 assign n_n2132 = ( wire388 ) | ( wire747 ) | ( wire21540 ) | ( wire21541 ) ;
 assign wire391 = ( n_n100  &  n_n256  &  wire907 ) | ( n_n100  &  n_n225  &  wire907 ) ;
 assign wire1158 = ( n_n281  &  wire913 ) | ( n_n281  &  wire903 ) ;
 assign n_n2080 = ( n_n2133 ) | ( n_n2132 ) | ( wire21549 ) ;
 assign wire1159 = ( wire153 ) | ( wire157 ) | ( wire330 ) | ( wire241 ) ;
 assign n_n2129 = ( wire3518 ) | ( wire21425 ) | ( n_n3  &  n_n186 ) ;
 assign wire1161 = ( n_n109 ) | ( wire79 ) | ( n_n101 ) | ( wire80 ) ;
 assign n_n2079 = ( n_n2129 ) | ( wire21431 ) | ( wire21432 ) ;
 assign n_n2274 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n26 ) | ( n_n53  &  n_n77 ) ;
 assign wire78 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign wire1163 = ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign n_n22 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire49 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) ;
 assign n_n1217 = ( wire2780 ) | ( wire2781 ) | ( wire22022 ) ;
 assign n_n4687 = ( n_n57  &  wire807 ) | ( n_n57  &  n_n279  &  wire904 ) ;
 assign n_n1284 = ( n_n4687 ) | ( wire22213 ) | ( wire22214 ) ;
 assign wire1167 = ( wire81 ) | ( n_n46 ) | ( n_n92 ) | ( wire19578 ) ;
 assign wire1169 = ( n_n113 ) | ( n_n36 ) | ( wire273 ) | ( wire57 ) ;
 assign n_n1138 = ( wire2503 ) | ( wire22294 ) | ( n_n53  &  wire1169 ) ;
 assign wire85 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire901 ) ;
 assign wire750 = ( n_n2  &  wire200 ) | ( n_n2  &  wire112 ) ;
 assign n_n1433 = ( n_n53  &  wire66 ) | ( n_n53  &  wire899  &  n_n256 ) ;
 assign wire41 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire932 = ( n_n2  &  wire901  &  n_n220 ) ;
 assign wire1171 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire907 ) ;
 assign n_n1120 = ( wire750 ) | ( wire22034 ) | ( wire22040 ) | ( wire22041 ) ;
 assign n_n1476 = ( n_n5  &  n_n197 ) | ( n_n6  &  wire62 ) ;
 assign n_n1126 = ( n_n4828 ) | ( n_n1476 ) | ( wire2776 ) | ( wire2777 ) ;
 assign n_n1142 = ( wire589 ) | ( wire2525 ) | ( wire2526 ) | ( wire22270 ) ;
 assign n_n1099 = ( n_n1140 ) | ( n_n1142 ) | ( wire2521 ) | ( wire22277 ) ;
 assign n_n3843 = ( n_n53  &  n_n95 ) | ( n_n48  &  wire81 ) ;
 assign wire662 = ( n_n53  &  wire19385 ) | ( n_n53  &  wire900  &  n_n256 ) ;
 assign n_n1584 = ( n_n57  &  n_n197 ) | ( n_n56  &  wire69 ) ;
 assign wire706 = ( n_n230  &  n_n271  &  wire165  &  n_n285 ) ;
 assign wire406 = ( n_n53  &  n_n222  &  wire899 ) | ( n_n53  &  wire899  &  n_n258 ) ;
 assign n_n952 = ( n_n53  &  n_n197 ) | ( n_n53  &  n_n223 ) | ( n_n53  &  n_n221 ) ;
 assign n_n819 = ( wire1984 ) | ( wire22736 ) | ( wire126  &  n_n5 ) ;
 assign n_n101 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire930 = ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n116 ) ;
 assign n_n5673 = ( (~ i_7_)  &  i_6_  &  n_n264  &  n_n116 ) ;
 assign n_n59 = ( i_14_  &  i_13_  &  i_12_  &  wire897 ) ;
 assign n_n148 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign n_n90 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire1181 = ( wire6020 ) | ( wire19269 ) | ( wire19270 ) | ( wire19271 ) ;
 assign wire1187 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign wire1186 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n5007 = ( n_n5020 ) | ( wire5885 ) | ( wire19223 ) | ( wire19230 ) ;
 assign wire936 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  n_n116 ) ;
 assign n_n4938 = ( n_n266  &  n_n230  &  n_n285  &  wire198 ) ;
 assign wire760 = ( n_n56  &  wire190 ) | ( n_n57  &  wire167 ) ;
 assign wire761 = ( n_n57  &  wire190 ) | ( n_n56  &  wire119 ) ;
 assign wire762 = ( n_n57  &  wire165 ) | ( n_n57  &  wire140 ) ;
 assign n_n4728 = ( wire573 ) | ( wire5075 ) | ( wire5076 ) | ( wire19878 ) ;
 assign wire247 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign wire119 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire763 = ( n_n266  &  n_n230  &  n_n285  &  wire119 ) ;
 assign wire541 = ( n_n5  &  n_n60 ) | ( n_n6  &  wire118 ) ;
 assign wire585 = ( n_n6  &  n_n59 ) | ( n_n5  &  wire132 ) ;
 assign n_n4183 = ( wire579 ) | ( wire764 ) | ( n_n54  &  n_n53 ) ;
 assign wire376 = ( n_n53  &  n_n220  &  wire907 ) | ( n_n53  &  n_n256  &  wire907 ) ;
 assign n_n4770 = ( n_n5  &  wire99 ) | ( n_n5  &  wire254 ) | ( n_n5  &  wire41 ) ;
 assign n_n4160 = ( n_n53  &  wire95 ) | ( n_n53  &  n_n228  &  wire912 ) ;
 assign n_n1645 = ( n_n94  &  wire1279 ) | ( n_n94  &  wire912  &  n_n225 ) ;
 assign wire586 = ( n_n100  &  n_n113 ) | ( n_n100  &  wire102 ) | ( n_n100  &  wire20526 ) ;
 assign wire767 = ( n_n100  &  wire368 ) | ( n_n100  &  n_n41 ) | ( n_n100  &  n_n88 ) ;
 assign n_n3136 = ( wire586 ) | ( wire767 ) | ( wire21098 ) | ( wire21101 ) ;
 assign n_n3309 = ( n_n48  &  n_n108 ) | ( n_n53  &  wire70 ) ;
 assign wire463 = ( n_n48  &  n_n246 ) | ( n_n48  &  n_n228  &  wire912 ) ;
 assign wire1192 = ( wire44 ) | ( n_n70 ) | ( n_n252 ) | ( wire79 ) ;
 assign n_n3124 = ( n_n3309 ) | ( wire20999 ) | ( wire21003 ) | ( wire21004 ) ;
 assign wire681 = ( wire3852 ) | ( n_n48  &  wire912  &  n_n256 ) ;
 assign n_n3123 = ( n_n3184 ) | ( wire681 ) | ( wire21013 ) | ( wire21014 ) ;
 assign n_n3099 = ( n_n3121 ) | ( n_n3122 ) | ( wire21034 ) | ( wire21035 ) ;
 assign n_n3101 = ( n_n3127 ) | ( n_n3128 ) | ( wire21054 ) ;
 assign n_n3587 = ( n_n53  &  wire42 ) | ( n_n53  &  n_n279  &  wire899 ) ;
 assign wire770 = ( n_n48  &  n_n76 ) | ( n_n48  &  n_n26 ) | ( n_n48  &  wire80 ) ;
 assign wire771 = ( n_n48  &  n_n29 ) | ( n_n48  &  wire49 ) | ( n_n48  &  wire88 ) ;
 assign n_n3103 = ( n_n3132 ) | ( n_n3133 ) | ( wire21095 ) ;
 assign n_n3104 = ( n_n3136 ) | ( n_n3135 ) | ( wire21116 ) ;
 assign wire553 = ( n_n56  &  n_n179 ) | ( n_n56  &  wire57 ) | ( n_n56  &  wire20194 ) ;
 assign wire653 = ( n_n57  &  n_n38 ) | ( n_n57  &  wire453 ) | ( n_n57  &  wire1902 ) ;
 assign wire548 = ( n_n94  &  n_n88 ) | ( n_n94  &  n_n258  &  wire912 ) ;
 assign wire773 = ( n_n100  &  wire165 ) | ( n_n100  &  wire140 ) ;
 assign wire774 = ( n_n100  &  n_n220  &  wire907 ) ;
 assign wire1194 = ( n_n113 ) | ( wire157 ) | ( wire57 ) | ( wire20056 ) ;
 assign n_n2665 = ( wire20060 ) | ( wire20061 ) | ( n_n94  &  wire1194 ) ;
 assign wire1196 = ( i_8_  &  n_n272  &  n_n260  &  n_n285 ) | ( (~ i_8_)  &  n_n272  &  n_n260  &  n_n285 ) ;
 assign wire1195 = ( wire911  &  n_n220 ) | ( n_n220  &  wire897 ) ;
 assign wire1198 = ( wire900  &  n_n220 ) | ( wire898  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire1201 = ( n_n25 ) | ( n_n24 ) | ( wire104 ) | ( wire228 ) ;
 assign n_n1765 = ( wire3005 ) | ( n_n5  &  wire1201 ) ;
 assign n_n1697 = ( wire3198 ) | ( wire21660 ) | ( wire21665 ) | ( wire21666 ) ;
 assign wire690 = ( n_n3  &  n_n50 ) | ( n_n3  &  n_n220  &  wire904 ) ;
 assign wire835 = ( wire3186 ) | ( n_n4  &  wire270 ) ;
 assign n_n1684 = ( n_n1697 ) | ( n_n1738 ) | ( wire21657 ) | ( wire21673 ) ;
 assign n_n1703 = ( wire835 ) | ( n_n1753 ) | ( wire3159 ) | ( wire21683 ) ;
 assign n_n1704 = ( n_n1757 ) | ( n_n1756 ) | ( wire21697 ) ;
 assign n_n1752 = ( wire21699 ) | ( wire21700 ) | ( wire21701 ) | ( wire21702 ) ;
 assign n_n1680 = ( n_n1684 ) | ( wire21648 ) | ( wire21649 ) | ( wire21711 ) ;
 assign wire56 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign n_n1356 = ( wire99  &  n_n229  &  n_n285  &  n_n284 ) ;
 assign n_n1208 = ( wire476 ) | ( n_n1356 ) | ( wire22043 ) | ( wire22044 ) ;
 assign n_n639 = ( n_n264  &  n_n273  &  n_n285  &  wire140 ) ;
 assign wire42 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire694 = ( n_n53  &  wire61 ) | ( n_n53  &  n_n281  &  wire902 ) ;
 assign wire869 = ( n_n53  &  n_n222  &  wire902 ) | ( n_n53  &  wire902  &  n_n258 ) ;
 assign n_n1121 = ( n_n1208 ) | ( wire22053 ) | ( wire22054 ) ;
 assign n_n876 = ( n_n4  &  wire469 ) | ( n_n4  &  n_n222  &  wire899 ) ;
 assign n_n790 = ( wire850 ) | ( wire22775 ) | ( wire22776 ) ;
 assign n_n7354 = ( n_n4  &  wire905  &  n_n256 ) ;
 assign wire743 = ( n_n4  &  n_n21 ) | ( n_n4  &  wire899  &  n_n258 ) ;
 assign wire1213 = ( n_n17 ) | ( wire514 ) | ( wire232 ) | ( wire22336 ) ;
 assign n_n349 = ( wire2465 ) | ( wire22338 ) | ( n_n3  &  wire1213 ) ;
 assign n_n7246 = ( n_n3  &  n_n256  &  wire904 ) ;
 assign wire833 = ( wire2463 ) | ( n_n4  &  wire906  &  n_n256 ) ;
 assign n_n351 = ( wire2457 ) | ( wire2458 ) | ( wire22348 ) ;
 assign n_n385 = ( wire22351 ) | ( n_n3  &  wire1257 ) ;
 assign wire642 = ( n_n4  &  n_n79 ) | ( n_n4  &  wire902  &  n_n258 ) ;
 assign wire1217 = ( n_n40 ) | ( wire245 ) | ( wire351 ) | ( wire22352 ) ;
 assign n_n49 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) ;
 assign wire590 = ( n_n5008 ) | ( wire19340 ) | ( wire19341 ) | ( wire19356 ) ;
 assign n_n5051 = ( n_n177  &  wire19284 ) | ( n_n177  &  wire19285 ) ;
 assign wire1223 = ( (~ i_9_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign n_n5017 = ( n_n5053 ) | ( n_n5051 ) | ( wire19288 ) ;
 assign wire1226 = ( i_7_  &  i_8_  &  i_6_ ) | ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n5008 = ( wire5874 ) | ( wire5875 ) | ( wire5876 ) ;
 assign wire1229 = ( n_n112 ) | ( n_n67 ) | ( wire84 ) | ( wire19738 ) ;
 assign n_n4729 = ( wire5268 ) | ( wire5269 ) | ( wire19881 ) | ( wire19882 ) ;
 assign n_n4633 = ( n_n6  &  wire65 ) | ( n_n6  &  wire902  &  n_n225 ) ;
 assign wire705 = ( n_n56  &  wire60 ) | ( n_n57  &  n_n108 ) ;
 assign wire1230 = ( n_n204 ) | ( n_n112 ) | ( wire52 ) | ( wire84 ) ;
 assign n_n4261 = ( wire705 ) | ( n_n56  &  wire1230 ) ;
 assign wire1231 = ( n_n264  &  n_n229  &  n_n165 ) | ( n_n229  &  n_n165  &  n_n230 ) ;
 assign n_n4218 = ( wire20719 ) | ( wire20720 ) | ( wire20721 ) | ( wire20722 ) ;
 assign n_n4199 = ( n_n4214 ) | ( n_n4255 ) | ( wire20729 ) | ( wire20733 ) ;
 assign wire140 = ( i_14_  &  i_13_  &  i_12_  &  wire908 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire157 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire914 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) ;
 assign n_n1370 = ( n_n265  &  n_n32 ) | ( n_n268  &  wire55 ) ;
 assign n_n4003 = ( n_n99  &  n_n53 ) | ( n_n53  &  wire96 ) | ( n_n53  &  wire20297 ) ;
 assign wire309 = ( wire5591 ) | ( wire5592 ) ;
 assign wire571 = ( n_n264  &  n_n275  &  n_n261  &  n_n285 ) ;
 assign wire737 = ( n_n264  &  n_n270  &  n_n263  &  n_n285 ) ;
 assign wire1234 = ( n_n46 ) | ( n_n92 ) | ( wire19577 ) | ( wire19578 ) ;
 assign n_n3928 = ( n_n4003 ) | ( wire20300 ) | ( wire20301 ) | ( wire20304 ) ;
 assign n_n3659 = ( wire5510 ) | ( wire5514 ) | ( wire5515 ) | ( wire19560 ) ;
 assign wire1237 = ( n_n16 ) | ( n_n68 ) | ( wire514 ) | ( wire20155 ) ;
 assign n_n3598 = ( n_n94  &  wire118 ) | ( n_n94  &  wire899  &  n_n220 ) ;
 assign wire208 = ( (~ i_15_)  &  n_n281  &  n_n270 ) | ( i_15_  &  n_n220  &  n_n270 ) ;
 assign n_n3209 = ( n_n3598 ) | ( wire3800 ) | ( wire21083 ) ;
 assign wire383 = ( n_n100  &  wire1855 ) | ( n_n100  &  wire902  &  n_n258 ) ;
 assign wire628 = ( n_n100  &  wire69 ) | ( n_n100  &  n_n78 ) | ( n_n100  &  wire80 ) ;
 assign n_n3135 = ( wire459 ) | ( n_n1633 ) | ( wire3771 ) | ( wire21105 ) ;
 assign n_n4644 = ( n_n6  &  wire368 ) | ( n_n6  &  n_n88 ) ;
 assign n_n4636 = ( n_n5  &  wire368 ) | ( n_n5  &  n_n88 ) ;
 assign wire317 = ( n_n111  &  n_n6 ) | ( n_n6  &  n_n38 ) | ( n_n6  &  wire1853 ) ;
 assign n_n3121 = ( wire317 ) | ( wire4745 ) | ( wire20131 ) | ( wire21019 ) ;
 assign n_n2890 = ( n_n6  &  n_n97 ) | ( n_n6  &  wire71 ) | ( n_n6  &  wire1905 ) ;
 assign n_n3122 = ( n_n2890 ) | ( wire21027 ) | ( wire21028 ) ;
 assign n_n4632 = ( n_n6  &  wire80 ) | ( n_n6  &  wire902  &  n_n256 ) ;
 assign wire487 = ( n_n6  &  n_n31 ) | ( n_n6  &  n_n80 ) | ( n_n6  &  wire88 ) ;
 assign wire742 = ( wire44  &  n_n208  &  n_n285  &  n_n284 ) ;
 assign wire931 = ( n_n208  &  n_n230  &  n_n285  &  wire232 ) ;
 assign wire1241 = ( n_n171 ) | ( n_n23 ) | ( wire56 ) | ( wire20362 ) ;
 assign n_n2876 = ( wire20364 ) | ( n_n207  &  wire1241 ) ;
 assign n_n3731 = ( n_n4  &  wire19407 ) | ( n_n4  &  n_n256  &  wire897 ) ;
 assign n_n1597 = ( n_n57  &  n_n104 ) | ( n_n56  &  wire78 ) ;
 assign n_n2437 = ( wire497 ) | ( n_n1597 ) | ( wire3594 ) | ( wire3595 ) ;
 assign n_n2429 = ( n_n2439 ) | ( n_n2437 ) | ( wire3588 ) | ( wire21318 ) ;
 assign wire271 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign wire472 = ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) ;
 assign n_n1788 = ( wire21723 ) | ( wire21724 ) ;
 assign n_n1715 = ( wire21713 ) | ( wire21714 ) | ( wire21718 ) | ( wire21719 ) ;
 assign wire1250 = ( wire911  &  n_n220 ) | ( wire902  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire1249 = ( wire899  &  n_n220 ) | ( wire902  &  n_n220 ) ;
 assign wire1248 = ( wire901  &  n_n220 ) | ( n_n220  &  wire897 ) ;
 assign n_n1792 = ( wire21729 ) | ( wire21730 ) | ( n_n57  &  wire165 ) ;
 assign wire158 = ( i_15_  &  n_n222  &  n_n282 ) | ( (~ i_15_)  &  n_n222  &  n_n282 ) ;
 assign wire1251 = ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n282 ) | ( (~ i_15_)  &  n_n222  &  n_n282 ) ;
 assign n_n1690 = ( n_n1788 ) | ( n_n1715 ) | ( wire21728 ) | ( wire21739 ) ;
 assign n_n1440 = ( n_n3  &  wire68 ) | ( n_n4  &  n_n42 ) ;
 assign wire300 = ( i_15_  &  n_n281  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n256 ) | ( (~ i_15_)  &  n_n267  &  n_n256 ) ;
 assign n_n1173 = ( n_n1440 ) | ( wire2811 ) | ( n_n4  &  wire300 ) ;
 assign n_n1210 = ( wire466 ) | ( wire2740 ) | ( wire22064 ) ;
 assign n_n6820 = ( n_n94  &  wire911  &  n_n225 ) ;
 assign wire1253 = ( wire899  &  n_n228 ) | ( n_n228  &  wire902 ) ;
 assign wire1254 = ( wire60 ) | ( n_n68 ) | ( wire22765 ) | ( wire22766 ) ;
 assign n_n789 = ( n_n265  &  wire85 ) | ( n_n268  &  wire1254 ) ;
 assign wire320 = ( (~ i_15_)  &  n_n275  &  n_n228 ) | ( i_15_  &  n_n275  &  n_n258 ) ;
 assign wire1257 = ( n_n199 ) | ( n_n73 ) | ( wire320 ) | ( wire22335 ) ;
 assign n_n370 = ( wire2308 ) | ( wire2309 ) | ( n_n13  &  wire191 ) ;
 assign wire1259 = ( wire276 ) | ( wire182 ) | ( wire405 ) | ( wire22477 ) ;
 assign n_n345 = ( n_n370 ) | ( wire2304 ) | ( wire2305 ) | ( wire22481 ) ;
 assign n_n377 = ( wire2296 ) | ( wire22483 ) | ( wire22485 ) | ( wire22487 ) ;
 assign n_n464 = ( wire877 ) | ( wire2277 ) | ( wire22495 ) | ( wire22496 ) ;
 assign wire688 = ( n_n94  &  wire912  &  n_n256 ) | ( n_n94  &  n_n256  &  wire914 ) ;
 assign wire798 = ( n_n260  &  n_n263  &  n_n285  &  wire112 ) ;
 assign wire1261 = ( n_n113 ) | ( wire140 ) | ( wire57 ) | ( wire358 ) ;
 assign n_n347 = ( n_n377 ) | ( wire22493 ) | ( wire22494 ) | ( wire22504 ) ;
 assign n_n96 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) ;
 assign n_n5048 = ( wire5988 ) | ( n_n152  &  wire282 ) | ( n_n152  &  wire19292 ) ;
 assign wire315 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) ;
 assign wire1265 = ( n_n283  &  n_n165  &  wire19294 ) | ( n_n283  &  n_n165  &  wire19296 ) ;
 assign wire1264 = ( n_n273  &  n_n165  &  wire19294 ) | ( n_n273  &  n_n165  &  wire19296 ) ;
 assign wire326 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n281 ) ;
 assign wire1271 = ( (~ i_8_)  &  n_n272 ) | ( i_8_  &  n_n272  &  wire19258 ) | ( i_8_  &  n_n272  &  wire19259 ) ;
 assign n_n5005 = ( wire19260 ) | ( wire19261 ) | ( wire19263 ) ;
 assign n_n4911 = ( n_n110  &  n_n57 ) | ( n_n56  &  wire82 ) ;
 assign wire632 = ( n_n6  &  n_n222  &  wire898 ) | ( n_n6  &  wire898  &  n_n258 ) ;
 assign wire198 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire902 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign wire137 = ( i_15_  &  n_n275  &  n_n228 ) | ( (~ i_15_)  &  n_n275  &  n_n258 ) ;
 assign wire112 = ( i_14_  &  i_13_  &  i_12_  &  wire907 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign wire80 = ( i_15_  &  n_n281  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign n_n3736 = ( n_n4  &  wire80 ) | ( n_n4  &  n_n256  &  wire908 ) ;
 assign n_n1339 = ( n_n4  &  n_n76 ) | ( n_n3  &  wire56 ) ;
 assign n_n3579 = ( n_n53  &  wire44 ) | ( n_n48  &  n_n65 ) ;
 assign wire1279 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire204 = ( wire71 ) | ( n_n256  &  wire904 ) ;
 assign n_n4674 = ( n_n56  &  wire71 ) | ( n_n56  &  n_n256  &  wire904 ) ;
 assign n_n3703 = ( n_n53  &  n_n49 ) | ( n_n53  &  wire71 ) | ( n_n53  &  wire19506 ) ;
 assign n_n3127 = ( n_n3703 ) | ( wire3830 ) | ( wire3831 ) | ( wire21038 ) ;
 assign n_n2875 = ( wire4492 ) | ( wire20366 ) | ( wire20367 ) ;
 assign n_n2145 = ( wire389 ) | ( wire3316 ) | ( wire3317 ) ;
 assign wire1286 = ( n_n99 ) | ( n_n52 ) | ( wire807 ) | ( wire226 ) ;
 assign n_n1785 = ( wire2972 ) | ( wire21832 ) | ( n_n53  &  wire1286 ) ;
 assign wire1291 = ( wire898  &  n_n220 ) | ( n_n220  &  wire912 ) | ( n_n220  &  wire897 ) ;
 assign wire1290 = ( wire902  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire1289 = ( wire901  &  n_n220 ) | ( wire900  &  n_n220 ) ;
 assign n_n1298 = ( wire2566 ) | ( wire22231 ) | ( wire22232 ) ;
 assign wire687 = ( n_n94  &  wire50 ) | ( n_n94  &  wire912  &  n_n256 ) ;
 assign n_n1212 = ( wire825 ) | ( wire687 ) | ( wire22066 ) | ( wire22067 ) ;
 assign wire374 = ( n_n4  &  n_n222  &  wire902 ) | ( n_n4  &  wire902  &  n_n258 ) ;
 assign wire434 = ( n_n100  &  n_n279  &  wire907 ) | ( n_n100  &  n_n228  &  wire907 ) ;
 assign wire799 = ( n_n4  &  wire165 ) | ( n_n4  &  wire140 ) ;
 assign n_n1123 = ( n_n1212 ) | ( wire22075 ) | ( wire22076 ) ;
 assign wire88 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n228  &  n_n270 ) ;
 assign n_n3615 = ( wire20755 ) | ( n_n100  &  wire898  &  n_n258 ) ;
 assign wire1305 = ( n_n41 ) | ( wire41 ) | ( wire175 ) | ( wire229 ) ;
 assign n_n5664 = ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire793 = ( i_7_  &  i_6_  &  n_n230  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n230  &  n_n116 ) ;
 assign wire874 = ( wire22240 ) | ( wire22241 ) | ( wire22242 ) ;
 assign wire1307 = ( n_n281  &  wire913 ) | ( n_n281  &  wire914 ) ;
 assign wire1311 = ( n_n113 ) | ( wire57 ) | ( wire22512 ) | ( wire22513 ) ;
 assign n_n407 = ( wire2258 ) | ( n_n1  &  n_n54 ) | ( n_n1  &  wire41 ) ;
 assign n_n408 = ( wire624 ) | ( wire22522 ) | ( n_n2  &  wire233 ) ;
 assign n_n340 = ( n_n407 ) | ( n_n408 ) | ( wire22524 ) | ( wire22527 ) ;
 assign n_n4736 = ( wire488 ) | ( wire878 ) | ( wire709 ) | ( wire19909 ) ;
 assign wire481 = ( n_n57  &  n_n220  &  wire905 ) | ( n_n57  &  wire905  &  n_n256 ) ;
 assign wire72 = ( (~ i_15_)  &  n_n281  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n220 ) ;
 assign wire273 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire219 = ( wire55 ) | ( n_n279  &  wire912 ) ;
 assign n_n4259 = ( n_n4912 ) | ( n_n4911 ) | ( n_n4913 ) ;
 assign wire721 = ( n_n4916 ) | ( n_n4915 ) | ( n_n4914 ) ;
 assign n_n4214 = ( n_n4259 ) | ( wire721 ) | ( wire20725 ) ;
 assign n_n4256 = ( wire5589 ) | ( wire20121 ) | ( n_n57  &  n_n12 ) ;
 assign n_n4255 = ( wire4756 ) | ( wire5011 ) | ( n_n57  &  wire101 ) ;
 assign wire465 = ( wire5552 ) | ( n_n57  &  wire44 ) ;
 assign n_n4774 = ( wire632 ) | ( wire5613 ) | ( n_n6  &  wire99 ) ;
 assign n_n3786 = ( n_n1  &  n_n95 ) | ( n_n2  &  wire81 ) ;
 assign n_n3782 = ( n_n2  &  n_n42 ) | ( n_n1  &  wire81 ) ;
 assign wire723 = ( n_n2  &  wire19385 ) | ( n_n2  &  wire900  &  n_n256 ) ;
 assign wire1320 = ( n_n93 ) | ( n_n90 ) | ( wire76 ) | ( wire19384 ) ;
 assign n_n3382 = ( n_n3782 ) | ( wire723 ) | ( wire19439 ) | ( wire19440 ) ;
 assign n_n4676 = ( n_n56  &  wire96 ) | ( n_n56  &  n_n222  &  wire904 ) ;
 assign n_n4686 = ( n_n57  &  wire71 ) | ( n_n57  &  n_n256  &  wire904 ) ;
 assign n_n3722 = ( n_n99  &  n_n100 ) | ( n_n100  &  wire96 ) | ( n_n100  &  wire19576 ) ;
 assign wire1322 = ( wire898  &  n_n258 ) | ( wire902  &  n_n258 ) | ( n_n258  &  wire912 ) ;
 assign n_n3221 = ( wire3764 ) | ( wire21108 ) | ( wire21109 ) | ( wire21110 ) ;
 assign wire1323 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n3128 = ( n_n3324 ) | ( n_n4381 ) | ( wire21046 ) | ( wire21047 ) ;
 assign wire1326 = ( n_n179 ) | ( n_n113 ) | ( wire55 ) | ( wire57 ) ;
 assign wire298 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  wire1852 ) ;
 assign wire521 = ( n_n53  &  n_n39 ) | ( n_n53  &  wire245 ) | ( n_n53  &  wire20454 ) ;
 assign n_n5675 = ( i_7_  &  i_6_  &  n_n284  &  n_n116 ) ;
 assign wire1327 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign n_n2146 = ( wire462 ) | ( wire3303 ) | ( wire21565 ) | ( wire21566 ) ;
 assign wire429 = ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) ;
 assign wire1329 = ( wire102 ) | ( wire263 ) | ( wire912  &  n_n256 ) ;
 assign wire1330 = ( wire898  &  n_n220 ) | ( n_n220  &  wire897 ) ;
 assign n_n1774 = ( wire21770 ) | ( wire21771 ) | ( wire21772 ) ;
 assign n_n1710 = ( n_n1774 ) | ( wire3032 ) | ( wire3033 ) ;
 assign n_n1536 = ( wire60  &  n_n48 ) | ( n_n53  &  n_n108 ) ;
 assign wire1333 = ( i_15_  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n228 ) ;
 assign n_n1295 = ( wire747 ) | ( wire22187 ) | ( wire22188 ) ;
 assign n_n1641 = ( n_n100  &  wire69 ) | ( n_n94  &  n_n103 ) ;
 assign wire1334 = ( i_15_  &  n_n247  &  n_n281 ) | ( (~ i_15_)  &  n_n247  &  n_n220 ) ;
 assign n_n4915 = ( n_n110  &  n_n56 ) | ( n_n57  &  wire60 ) ;
 assign wire589 = ( n_n56  &  n_n197 ) | ( n_n57  &  wire62 ) ;
 assign wire679 = ( n_n53  &  n_n144 ) | ( n_n48  &  n_n8 ) ;
 assign n_n3884 = ( n_n100  &  wire19577 ) | ( n_n100  &  n_n228  &  wire906 ) ;
 assign n_n809 = ( wire931 ) | ( wire580 ) | ( wire22796 ) | ( wire22797 ) ;
 assign wire1340 = ( i_15_  &  n_n247  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) | ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire483 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  wire88 ) ;
 assign wire1343 = ( i_15_  &  n_n247  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) | ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire1345 = ( i_8_  &  n_n231  &  n_n285  &  n_n284 ) | ( (~ i_8_)  &  n_n231  &  n_n285  &  n_n284 ) ;
 assign wire1344 = ( wire903  &  n_n258 ) | ( n_n258  &  wire907 ) ;
 assign wire1347 = ( n_n109 ) | ( wire143 ) | ( wire306 ) | ( wire22363 ) ;
 assign wire1346 = ( wire913  &  n_n256 ) | ( n_n258  &  wire904 ) ;
 assign wire408 = ( (~ i_15_)  &  n_n228  &  n_n267 ) | ( i_15_  &  n_n258  &  n_n267 ) ;
 assign wire933 = ( n_n268  &  wire913  &  n_n258 ) ;
 assign wire1349 = ( n_n10 ) | ( n_n83 ) | ( wire233 ) | ( wire414 ) ;
 assign wire1348 = ( n_n52 ) | ( n_n49 ) | ( wire357 ) | ( wire22340 ) ;
 assign n_n352 = ( wire2243 ) | ( wire22533 ) | ( n_n265  &  wire1349 ) ;
 assign wire1354 = ( i_8_  &  n_n260  &  n_n155  &  n_n285 ) | ( (~ i_8_)  &  n_n260  &  n_n155  &  n_n285 ) ;
 assign wire1357 = ( n_n258  &  wire914 ) | ( n_n258  &  wire904 ) ;
 assign wire1355 = ( n_n258  &  wire906 ) | ( n_n258  &  wire907 ) ;
 assign n_n339 = ( n_n352 ) | ( wire22536 ) | ( wire22537 ) | ( wire22544 ) ;
 assign wire1359 = ( n_n133 ) | ( n_n135 ) | ( wire419 ) | ( wire19604 ) ;
 assign wire113 = ( (~ i_15_)  &  n_n281  &  n_n282 ) | ( i_15_  &  n_n220  &  n_n282 ) ;
 assign n_n4913 = ( n_n57  &  wire84 ) | ( n_n57  &  n_n279  &  wire913 ) ;
 assign n_n4146 = ( wire406 ) | ( n_n3587 ) | ( wire478 ) | ( wire20344 ) ;
 assign n_n3925 = ( wire470 ) | ( wire4602 ) | ( wire20253 ) | ( wire20254 ) ;
 assign n_n3914 = ( n_n3964 ) | ( wire3636 ) | ( wire21250 ) ;
 assign n_n3930 = ( wire3707 ) | ( wire3708 ) | ( wire21188 ) ;
 assign n_n3929 = ( wire3702 ) | ( wire21190 ) | ( wire21191 ) ;
 assign n_n3991 = ( n_n48  &  n_n200 ) | ( n_n48  &  wire104 ) | ( n_n48  &  wire20256 ) ;
 assign n_n3923 = ( wire4586 ) | ( wire4587 ) | ( wire20259 ) | ( wire20262 ) ;
 assign wire478 = ( n_n53  &  n_n77 ) | ( n_n53  &  n_n281  &  wire902 ) ;
 assign wire1363 = ( n_n200 ) | ( n_n25 ) | ( wire104 ) | ( wire19457 ) ;
 assign n_n3900 = ( n_n3925 ) | ( n_n3923 ) | ( wire20271 ) ;
 assign n_n3920 = ( n_n3978 ) | ( n_n3980 ) | ( wire20282 ) ;
 assign n_n3922 = ( wire4557 ) | ( wire4558 ) | ( wire20287 ) ;
 assign n_n3899 = ( n_n3920 ) | ( n_n3922 ) | ( wire4552 ) | ( wire20293 ) ;
 assign n_n3926 = ( n_n4174 ) | ( wire4529 ) | ( wire4530 ) | ( wire20310 ) ;
 assign n_n3901 = ( n_n3928 ) | ( n_n3926 ) | ( wire20319 ) ;
 assign wire1368 = ( n_n92 ) | ( n_n43 ) | ( wire59 ) | ( wire19578 ) ;
 assign n_n3404 = ( wire5478 ) | ( wire19581 ) | ( wire19582 ) ;
 assign n_n3486 = ( n_n3610 ) | ( wire4131 ) | ( wire20756 ) ;
 assign n_n3403 = ( n_n3486 ) | ( wire20764 ) | ( wire20765 ) ;
 assign n_n3372 = ( n_n3404 ) | ( n_n3403 ) | ( wire19586 ) | ( wire20770 ) ;
 assign n_n2713 = ( n_n145  &  n_n100 ) | ( n_n94  &  wire225 ) ;
 assign wire121 = ( wire44 ) | ( n_n258  &  wire904 ) ;
 assign wire370 = ( wire863 ) | ( n_n4687 ) | ( wire5506 ) ;
 assign wire493 = ( wire4789 ) | ( n_n94  &  wire130 ) ;
 assign n_n3371 = ( wire20774 ) | ( wire20775 ) | ( wire20781 ) | ( wire20782 ) ;
 assign n_n3398 = ( n_n4915 ) | ( n_n4913 ) | ( wire19935 ) | ( wire19936 ) ;
 assign n_n3397 = ( n_n4912 ) | ( n_n4911 ) | ( n_n4781 ) | ( wire19914 ) ;
 assign wire788 = ( n_n56  &  n_n95 ) | ( n_n56  &  n_n49 ) | ( n_n56  &  wire71 ) ;
 assign n_n3361 = ( n_n3372 ) | ( n_n3371 ) | ( wire20788 ) ;
 assign n_n3132 = ( wire370 ) | ( wire788 ) | ( wire21077 ) | ( wire21081 ) ;
 assign n_n2820 = ( wire411 ) | ( wire647 ) | ( n_n2882 ) | ( wire4500 ) ;
 assign n_n2818 = ( n_n2876 ) | ( n_n2875 ) | ( wire20374 ) ;
 assign wire1371 = ( wire160 ) | ( wire184 ) | ( wire132 ) | ( wire20376 ) ;
 assign n_n2798 = ( n_n2820 ) | ( n_n2818 ) | ( wire20381 ) | ( wire20382 ) ;
 assign wire1372 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) ;
 assign wire1376 = ( wire51 ) | ( n_n93 ) | ( n_n90 ) | ( wire21389 ) ;
 assign n_n2158 = ( wire3398 ) | ( n_n53  &  wire1376 ) ;
 assign wire1378 = ( n_n281  &  wire913 ) | ( n_n281  &  wire905 ) | ( n_n281  &  wire908 ) ;
 assign wire1377 = ( i_8_  &  n_n153  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n153  &  n_n230  &  n_n285 ) ;
 assign n_n4682 = ( n_n56  &  wire19384 ) | ( n_n56  &  n_n281  &  wire900 ) ;
 assign n_n2172 = ( n_n4686 ) | ( wire21445 ) | ( wire21446 ) ;
 assign wire98 = ( wire19384 ) | ( n_n281  &  wire900 ) ;
 assign wire482 = ( i_15_  &  n_n253  &  n_n279 ) | ( (~ i_15_)  &  n_n253  &  n_n279 ) ;
 assign wire1379 = ( i_15_  &  n_n279  &  n_n267 ) | ( (~ i_15_)  &  n_n279  &  n_n267 ) ;
 assign n_n2093 = ( n_n2172 ) | ( wire3452 ) | ( wire21449 ) | ( wire21453 ) ;
 assign n_n4666 = ( n_n57  &  wire86 ) | ( n_n57  &  n_n256  &  wire907 ) ;
 assign wire1383 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign n_n2067 = ( n_n2093 ) | ( wire21462 ) | ( wire21463 ) | ( wire21470 ) ;
 assign wire425 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire897 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire897 ) ;
 assign wire657 = ( n_n94  &  wire228 ) | ( n_n94  &  n_n256  &  wire897 ) ;
 assign n_n1804 = ( wire657 ) | ( wire2939 ) | ( wire21857 ) ;
 assign wire1387 = ( wire51 ) | ( n_n105 ) | ( n_n90 ) | ( wire448 ) ;
 assign n_n1092 = ( n_n1120 ) | ( n_n1121 ) | ( wire2745 ) | ( wire22061 ) ;
 assign wire73 = ( (~ i_15_)  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign n_n1108 = ( wire2858 ) | ( wire21935 ) | ( n_n4  &  wire1491 ) ;
 assign n_n1109 = ( wire2854 ) | ( wire21941 ) | ( n_n4  &  wire1492 ) ;
 assign wire519 = ( n_n3  &  wire40 ) | ( n_n4  &  n_n103 ) ;
 assign n_n743 = ( n_n771 ) | ( n_n770 ) | ( wire22625 ) | ( wire22626 ) ;
 assign n_n742 = ( wire22646 ) | ( wire22647 ) ;
 assign wire139 = ( i_15_  &  n_n267  &  n_n225 ) | ( (~ i_15_)  &  n_n267  &  n_n225 ) ;
 assign wire776 = ( n_n105  &  n_n94 ) | ( n_n94  &  n_n46 ) | ( n_n94  &  wire19577 ) ;
 assign n_n744 = ( n_n772 ) | ( wire22662 ) | ( wire22663 ) | ( wire22670 ) ;
 assign wire929 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n116 ) ;
 assign n_n5679 = ( i_7_  &  i_6_  &  n_n230  &  n_n116 ) ;
 assign wire1400 = ( wire321 ) | ( wire331 ) | ( wire19319 ) | ( wire19320 ) ;
 assign wire546 = ( n_n4  &  n_n13 ) | ( n_n4  &  wire900  &  n_n228 ) ;
 assign wire634 = ( n_n3  &  n_n66 ) | ( n_n4  &  n_n64 ) ;
 assign n_n3915 = ( wire736 ) | ( wire21257 ) | ( wire21258 ) ;
 assign n_n3406 = ( wire4089 ) | ( wire4090 ) | ( n_n3  &  n_n226 ) ;
 assign n_n3932 = ( n_n4015 ) | ( wire3698 ) | ( wire21193 ) ;
 assign n_n3904 = ( n_n3932 ) | ( wire21200 ) | ( wire21201 ) ;
 assign n_n3806 = ( n_n5  &  n_n59 ) | ( n_n6  &  wire208 ) ;
 assign n_n3408 = ( wire546 ) | ( wire5780 ) | ( wire19381 ) ;
 assign n_n3374 = ( n_n3408 ) | ( wire4080 ) | ( wire20793 ) ;
 assign wire545 = ( n_n4  &  n_n204 ) | ( n_n4  &  wire52 ) | ( n_n4  &  wire20579 ) ;
 assign n_n3375 = ( wire545 ) | ( wire4076 ) | ( wire20798 ) ;
 assign wire633 = ( wire19400 ) | ( wire19401 ) | ( n_n3  &  n_n15 ) ;
 assign n_n3362 = ( n_n3374 ) | ( n_n3375 ) | ( wire20804 ) ;
 assign n_n2832 = ( wire460 ) | ( wire653 ) | ( wire4391 ) | ( wire20488 ) ;
 assign n_n2817 = ( wire4472 ) | ( wire20397 ) | ( wire20400 ) | ( wire20403 ) ;
 assign wire533 = ( wire4470 ) | ( n_n4  &  n_n92 ) | ( n_n4  &  wire19578 ) ;
 assign n_n2797 = ( n_n2815 ) | ( n_n2817 ) | ( wire20412 ) ;
 assign n_n2792 = ( n_n2799 ) | ( n_n2801 ) | ( wire20484 ) ;
 assign n_n2793 = ( n_n2803 ) | ( n_n2804 ) | ( wire20553 ) ;
 assign n_n2796 = ( n_n2813 ) | ( wire4319 ) | ( wire20559 ) | ( wire20568 ) ;
 assign n_n2140 = ( wire3292 ) | ( wire21574 ) | ( n_n5  &  wire67 ) ;
 assign n_n2099 = ( wire3370 ) | ( wire21516 ) | ( wire21517 ) ;
 assign wire1413 = ( wire119 ) | ( wire281 ) | ( wire338 ) | ( wire858 ) ;
 assign wire1416 = ( wire153 ) | ( wire255 ) | ( wire241 ) | ( wire242 ) ;
 assign n_n2097 = ( n_n100  &  wire1416 ) | ( n_n94  &  wire1416 ) | ( n_n100  &  wire330 ) ;
 assign n_n2180 = ( wire391 ) | ( wire3419 ) | ( wire21482 ) | ( wire21483 ) ;
 assign wire1423 = ( i_8_  &  n_n260  &  n_n155  &  n_n285 ) | ( (~ i_8_)  &  n_n260  &  n_n155  &  n_n285 ) ;
 assign n_n3770 = ( n_n1  &  n_n76 ) | ( n_n2  &  wire56 ) ;
 assign wire1424 = ( n_n79 ) | ( wire212 ) | ( wire49 ) | ( wire21963 ) ;
 assign n_n1111 = ( wire2798 ) | ( wire2804 ) | ( wire22000 ) | ( wire22007 ) ;
 assign wire276 = ( (~ i_15_)  &  n_n228  &  n_n270 ) | ( i_15_  &  n_n258  &  n_n270 ) ;
 assign wire587 = ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n260 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n260 ) ;
 assign wire66 = ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n225 ) ;
 assign n_n3980 = ( n_n4160 ) | ( wire4565 ) | ( wire20275 ) ;
 assign wire1439 = ( wire368 ) | ( n_n88 ) | ( n_n113 ) | ( wire102 ) ;
 assign n_n3895 = ( n_n3908 ) | ( wire3660 ) | ( wire3661 ) | ( wire21236 ) ;
 assign wire816 = ( n_n56  &  wire903  &  n_n220 ) ;
 assign n_n3709 = ( wire816 ) | ( n_n57  &  wire147 ) | ( n_n57  &  wire19535 ) ;
 assign wire1442 = ( n_n20 ) | ( wire79 ) | ( n_n72 ) | ( wire66 ) ;
 assign n_n2926 = ( n_n100  &  n_n221 ) | ( n_n100  &  wire469 ) | ( n_n100  &  wire1442 ) ;
 assign wire882 = ( n_n53  &  n_n62 ) | ( n_n53  &  n_n281  &  wire907 ) ;
 assign n_n2824 = ( wire4453 ) | ( wire20429 ) | ( wire20430 ) ;
 assign n_n2799 = ( n_n2822 ) | ( n_n2821 ) | ( wire20452 ) ;
 assign n_n2801 = ( n_n2827 ) | ( wire4414 ) | ( wire20469 ) | ( wire20475 ) ;
 assign wire1445 = ( n_n171 ) | ( n_n22 ) | ( wire56 ) | ( wire53 ) ;
 assign n_n2830 = ( n_n4913 ) | ( n_n4914 ) | ( wire4384 ) | ( wire20495 ) ;
 assign n_n2803 = ( n_n2833 ) | ( n_n2835 ) | ( wire4360 ) | ( wire20516 ) ;
 assign n_n2804 = ( n_n2837 ) | ( wire20541 ) | ( wire20542 ) | ( wire20543 ) ;
 assign wire693 = ( n_n57  &  wire19408 ) | ( n_n57  &  wire903  &  n_n256 ) ;
 assign n_n2154 = ( wire479 ) | ( wire478 ) | ( wire3277 ) | ( wire21590 ) ;
 assign wire1449 = ( wire48 ) | ( wire62 ) | ( n_n204 ) | ( n_n16 ) ;
 assign n_n2100 = ( wire3368 ) | ( n_n4  &  wire1449 ) ;
 assign wire1450 = ( n_n281  &  wire903 ) | ( n_n281  &  wire914 ) | ( n_n281  &  wire908 ) ;
 assign wire1451 = ( wire898  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire823 = ( n_n268  &  wire124 ) | ( n_n268  &  wire212 ) ;
 assign n_n1124 = ( n_n1215 ) | ( wire22087 ) | ( wire22088 ) ;
 assign n_n1093 = ( n_n1123 ) | ( n_n1124 ) | ( wire22095 ) ;
 assign wire381 = ( n_n94  &  n_n203 ) | ( n_n94  &  n_n279  &  wire911 ) ;
 assign n_n5677 = ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n116 ) ;
 assign wire384 = ( n_n282  &  wire152 ) | ( i_15_  &  n_n281  &  n_n282 ) ;
 assign wire621 = ( n_n264  &  wire69  &  n_n283  &  n_n285 ) ;
 assign n_n3913 = ( n_n1370 ) | ( wire3619 ) | ( wire3620 ) | ( wire21281 ) ;
 assign n_n3133 = ( n_n3209 ) | ( wire21089 ) | ( wire21090 ) ;
 assign wire1463 = ( wire20573 ) | ( wire20574 ) | ( wire20575 ) | ( wire20576 ) ;
 assign n_n2808 = ( n_n4  &  n_n39 ) | ( n_n4  &  wire1463 ) | ( n_n4  &  wire245 ) ;
 assign n_n2822 = ( wire317 ) | ( wire4444 ) | ( wire20435 ) ;
 assign n_n2821 = ( wire4435 ) | ( wire20437 ) | ( wire20441 ) | ( wire20442 ) ;
 assign n_n2806 = ( n_n7354 ) | ( wire545 ) | ( wire4302 ) | ( wire20583 ) ;
 assign wire792 = ( n_n4  &  n_n171 ) | ( n_n4  &  wire56 ) | ( n_n4  &  wire53 ) ;
 assign n_n2155 = ( wire464 ) | ( wire376 ) | ( wire3272 ) | ( wire21593 ) ;
 assign wire1469 = ( wire67 ) | ( n_n85 ) | ( wire54 ) | ( wire21596 ) ;
 assign n_n2088 = ( n_n2155 ) | ( wire3270 ) | ( n_n53  &  wire1469 ) ;
 assign n_n3751 = ( n_n271  &  n_n285  &  n_n284  &  wire212 ) ;
 assign wire380 = ( n_n94  &  n_n281  &  wire897 ) | ( n_n94  &  n_n256  &  wire897 ) ;
 assign wire826 = ( n_n163  &  n_n260  &  n_n229  &  n_n165 ) ;
 assign wire1475 = ( n_n111 ) | ( n_n108 ) | ( wire54 ) | ( wire103 ) ;
 assign wire1474 = ( n_n260  &  n_n208  &  n_n165 ) | ( n_n260  &  n_n273  &  n_n165 ) ;
 assign wire101 = ( i_15_  &  n_n228  &  n_n282 ) | ( (~ i_15_)  &  n_n258  &  n_n282 ) ;
 assign n_n2827 = ( wire298 ) | ( wire521 ) | ( wire20457 ) ;
 assign n_n4914 = ( n_n57  &  wire52 ) | ( n_n57  &  n_n279  &  wire911 ) ;
 assign n_n2813 = ( n_n3772 ) | ( n_n2603 ) | ( wire395 ) | ( wire20562 ) ;
 assign wire829 = ( n_n1  &  n_n171 ) | ( n_n1  &  wire56 ) | ( n_n1  &  wire53 ) ;
 assign wire1483 = ( wire82 ) | ( n_n73 ) | ( n_n22 ) | ( wire19408 ) ;
 assign wire1484 = ( n_n7 ) | ( n_n38 ) | ( wire453 ) | ( wire21379 ) ;
 assign wire330 = ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n281 ) ;
 assign wire1485 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign n_n2085 = ( n_n2148 ) | ( n_n2146 ) | ( wire21572 ) ;
 assign wire1486 = ( wire40 ) | ( n_n74 ) | ( wire21367 ) | ( wire21551 ) ;
 assign wire624 = ( n_n53  &  wire899  &  n_n256 ) | ( n_n53  &  wire905  &  n_n256 ) ;
 assign wire1489 = ( n_n21 ) | ( n_n72 ) | ( wire66 ) | ( wire343 ) ;
 assign wire1488 = ( n_n112 ) | ( n_n27 ) | ( wire247 ) | ( wire52 ) ;
 assign wire1491 = ( wire200 ) | ( n_n79 ) | ( wire112 ) | ( wire21930 ) ;
 assign wire1492 = ( wire67 ) | ( n_n135 ) | ( wire85 ) | ( wire347 ) ;
 assign n_n834 = ( wire2019 ) | ( wire22710 ) ;
 assign n_n560 = ( n_n264  &  n_n273  &  n_n285  &  wire123 ) ;
 assign n_n5009 = ( wire5834 ) | ( wire5835 ) | ( wire5843 ) | ( wire5844 ) ;
 assign wire716 = ( wire4478 ) | ( n_n4  &  n_n221 ) | ( n_n4  &  wire469 ) ;
 assign wire821 = ( n_n260  &  n_n261  &  wire77  &  n_n285 ) ;
 assign n_n2837 = ( wire586 ) | ( wire4344 ) | ( wire20532 ) | ( wire20533 ) ;
 assign n_n2086 = ( n_n2149 ) | ( wire3261 ) | ( wire3262 ) | ( wire21605 ) ;
 assign n_n2083 = ( n_n2140 ) | ( wire3287 ) | ( wire3288 ) | ( wire21579 ) ;
 assign n_n1598 = ( n_n111  &  n_n57 ) | ( n_n56  &  wire85 ) ;
 assign wire704 = ( n_n56  &  wire200 ) | ( n_n56  &  wire112 ) ;
 assign n_n3523 = ( n_n1  &  n_n110 ) | ( n_n2  &  wire82 ) ;
 assign wire1514 = ( n_n252 ) | ( wire73 ) | ( wire100 ) | ( wire21975 ) ;
 assign n_n1591 = ( n_n57  &  wire69 ) | ( n_n56  &  n_n103 ) ;
 assign wire144 = ( i_15_  &  n_n256  &  n_n282 ) | ( (~ i_15_)  &  n_n256  &  n_n282 ) ;
 assign wire877 = ( n_n100  &  n_n36 ) | ( n_n100  &  n_n35 ) | ( n_n100  &  n_n83 ) ;
 assign n_n618 = ( n_n48  &  n_n41 ) | ( n_n53  &  wire144 ) ;
 assign n_n438 = ( n_n6848 ) | ( n_n618 ) | ( wire2374 ) | ( wire22414 ) ;
 assign wire1517 = ( i_8_  &  n_n264  &  n_n155  &  n_n285 ) | ( (~ i_8_)  &  n_n264  &  n_n155  &  n_n285 ) ;
 assign n_n4781 = ( wire5550 ) | ( wire5552 ) | ( n_n57  &  wire44 ) ;
 assign n_n4733 = ( wire5244 ) | ( wire5245 ) | ( wire19864 ) | ( wire19865 ) ;
 assign n_n4773 = ( wire389 ) | ( wire708 ) | ( n_n5  &  wire166 ) ;
 assign n_n4680 = ( n_n57  &  wire76 ) | ( n_n57  &  n_n279  &  wire900 ) ;
 assign wire468 = ( n_n1  &  wire60 ) | ( n_n1  &  n_n204 ) | ( n_n1  &  wire52 ) ;
 assign wire1528 = ( wire40 ) | ( n_n74 ) | ( wire21367 ) | ( wire21609 ) ;
 assign wire369 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) ;
 assign wire1530 = ( i_15_  &  n_n275  &  n_n279 ) | ( (~ i_15_)  &  n_n275  &  n_n279 ) | ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign wire233 = ( (~ i_15_)  &  n_n228  &  n_n282 ) | ( i_15_  &  n_n258  &  n_n282 ) ;
 assign wire1540 = ( wire40 ) | ( wire899  &  n_n258 ) ;
 assign n_n4489 = ( wire48  &  n_n128 ) | ( n_n130  &  n_n111 ) ;
 assign n_n4677 = ( n_n56  &  wire68 ) | ( n_n57  &  n_n42 ) ;
 assign wire371 = ( n_n279  &  wire913 ) | ( n_n279  &  wire914 ) ;
 assign wire1545 = ( n_n279  &  wire913 ) | ( n_n279  &  wire905 ) | ( n_n279  &  wire914 ) ;
 assign n_n4598 = ( wire20192 ) | ( n_n130  &  n_n163 ) | ( n_n130  &  wire1545 ) ;
 assign n_n4585 = ( wire20117 ) | ( n_n6  &  wire1905 ) ;
 assign n_n4555 = ( wire4655 ) | ( wire20199 ) | ( wire20200 ) ;
 assign n_n3711 = ( wire5546 ) | ( n_n57  &  n_n76 ) | ( n_n57  &  wire1856 ) ;
 assign n_n3710 = ( n_n56  &  n_n73 ) | ( n_n56  &  wire19408 ) | ( n_n56  &  wire19536 ) ;
 assign wire1547 = ( n_n81 ) | ( n_n35 ) | ( wire64 ) | ( wire86 ) ;
 assign n_n4536 = ( n_n4555 ) | ( n_n3711 ) | ( wire20205 ) | ( wire20209 ) ;
 assign n_n5672 = ( i_7_  &  (~ i_6_)  &  n_n264  &  n_n116 ) ;
 assign wire1552 = ( wire190 ) | ( wire124 ) | ( wire212 ) | ( wire119 ) ;
 assign n_n3390 = ( wire674 ) | ( n_n4773 ) | ( wire5629 ) | ( wire19485 ) ;
 assign n_n3624 = ( n_n3638 ) | ( n_n3637 ) | ( wire19398 ) ;
 assign n_n3634 = ( n_n7424 ) | ( n_n3727 ) | ( wire5744 ) | ( wire19405 ) ;
 assign n_n3636 = ( n_n1339 ) | ( wire5733 ) | ( wire5734 ) | ( wire19413 ) ;
 assign wire1555 = ( n_n73 ) | ( wire70 ) | ( n_n22 ) | ( wire19408 ) ;
 assign n_n3550 = ( n_n240  &  n_n227 ) | ( n_n240  &  n_n207 ) | ( n_n227  &  n_n257 ) ;
 assign wire1557 = ( n_n223 ) | ( n_n67 ) | ( wire42 ) | ( wire19738 ) ;
 assign n_n3380 = ( wire468 ) | ( wire5195 ) | ( wire20861 ) | ( wire20862 ) ;
 assign n_n3395 = ( n_n3843 ) | ( n_n3703 ) | ( wire5569 ) | ( wire5570 ) ;
 assign n_n3369 = ( n_n3395 ) | ( wire19511 ) | ( wire19512 ) | ( wire20836 ) ;
 assign n_n3417 = ( wire455 ) | ( n_n3  &  wire43 ) | ( n_n3  &  wire19386 ) ;
 assign n_n3378 = ( wire4071 ) | ( wire4072 ) | ( wire4073 ) | ( wire20809 ) ;
 assign wire597 = ( n_n4  &  wire68 ) | ( n_n4  &  wire1891 ) ;
 assign n_n2597 = ( wire5725 ) | ( wire5726 ) ;
 assign n_n2598 = ( n_n3768 ) | ( wire829 ) | ( n_n2  &  n_n22 ) ;
 assign n_n2579 = ( n_n2598 ) | ( wire5725 ) | ( wire5726 ) | ( wire19768 ) ;
 assign wire154 = ( i_15_  &  n_n281  &  n_n282 ) | ( (~ i_15_)  &  n_n220  &  n_n282 ) ;
 assign n_n1781 = ( wire2975 ) | ( wire2976 ) | ( wire21827 ) | ( wire21828 ) ;
 assign n_n785 = ( n_n896 ) | ( wire712 ) | ( n_n4  &  wire139 ) ;
 assign n_n413 = ( wire434 ) | ( wire22546 ) | ( wire22547 ) | ( wire22548 ) ;
 assign wire471 = ( n_n94  &  n_n279  &  wire903 ) | ( n_n94  &  n_n222  &  wire903 ) ;
 assign wire658 = ( n_n94  &  wire903  &  n_n256 ) | ( n_n94  &  n_n256  &  wire897 ) ;
 assign n_n359 = ( n_n413 ) | ( wire22556 ) | ( wire22557 ) | ( wire22558 ) ;
 assign wire136 = ( wire57 ) | ( n_n279  &  wire912 ) ;
 assign n_n4732 = ( wire5238 ) | ( wire5239 ) | ( wire19899 ) | ( wire19900 ) ;
 assign wire147 = ( wire53 ) | ( n_n279  &  wire897 ) ;
 assign wire1575 = ( n_n279  &  wire913 ) | ( n_n279  &  wire905 ) | ( n_n279  &  wire914 ) ;
 assign n_n4685 = ( n_n57  &  n_n95 ) | ( n_n56  &  wire81 ) ;
 assign wire1577 = ( n_n93 ) | ( n_n44 ) | ( wire76 ) | ( wire19385 ) ;
 assign n_n4556 = ( n_n4680 ) | ( n_n4677 ) | ( wire20219 ) | ( wire20220 ) ;
 assign n_n3638 = ( n_n3417 ) | ( wire597 ) | ( wire19387 ) ;
 assign n_n3650 = ( n_n4774 ) | ( wire5607 ) | ( wire19495 ) ;
 assign n_n3629 = ( n_n3650 ) | ( wire19489 ) | ( wire19490 ) | ( wire19504 ) ;
 assign n_n3424 = ( wire5718 ) | ( wire5720 ) | ( n_n1  &  wire44 ) ;
 assign n_n3379 = ( n_n3424 ) | ( wire20865 ) | ( wire20866 ) ;
 assign wire1585 = ( n_n204 ) | ( n_n112 ) | ( wire52 ) | ( wire84 ) ;
 assign n_n3367 = ( n_n3390 ) | ( wire4042 ) | ( wire4043 ) | ( wire20844 ) ;
 assign n_n3393 = ( wire4027 ) | ( wire4028 ) | ( wire20849 ) ;
 assign n_n3360 = ( n_n3369 ) | ( n_n3367 ) | ( wire20858 ) ;
 assign n_n2833 = ( wire370 ) | ( wire20501 ) | ( wire20502 ) ;
 assign n_n2633 = ( n_n2  &  wire60 ) | ( n_n1  &  n_n108 ) ;
 assign n_n2599 = ( n_n2  &  n_n73 ) | ( n_n2  &  wire19408 ) | ( n_n2  &  wire19424 ) ;
 assign wire812 = ( n_n3772 ) | ( n_n3770 ) | ( wire5711 ) ;
 assign n_n2580 = ( n_n2599 ) | ( wire812 ) | ( wire19770 ) ;
 assign wire1593 = ( n_n281  &  wire913 ) | ( n_n281  &  wire914 ) ;
 assign wire1594 = ( n_n44 ) | ( wire270 ) | ( wire21668 ) | ( wire21834 ) ;
 assign n_n1713 = ( n_n1785 ) | ( wire2967 ) | ( n_n53  &  wire1594 ) ;
 assign wire1597 = ( n_n17 ) | ( wire195 ) | ( wire21748 ) | ( wire21749 ) ;
 assign wire1596 = ( n_n20 ) | ( wire375 ) | ( wire240 ) | ( wire21746 ) ;
 assign wire1599 = ( n_n20 ) | ( wire375 ) | ( wire240 ) | ( wire857 ) ;
 assign wire494 = ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign wire1600 = ( i_15_  &  n_n253  &  n_n222 ) | ( (~ i_15_)  &  n_n253  &  n_n222 ) | ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) ;
 assign n_n1691 = ( wire21766 ) | ( wire21767 ) | ( wire21769 ) ;
 assign wire514 = ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign n_n787 = ( wire862 ) | ( wire895 ) | ( n_n265  &  n_n63 ) ;
 assign n_n749 = ( n_n789 ) | ( n_n787 ) | ( wire855 ) | ( wire856 ) ;
 assign wire1606 = ( wire901  &  n_n228 ) | ( n_n228  &  wire902 ) | ( n_n228  &  wire912 ) ;
 assign n_n750 = ( n_n790 ) | ( wire847 ) | ( wire22778 ) | ( wire22781 ) ;
 assign n_n409 = ( wire22561 ) | ( wire22562 ) | ( wire22565 ) ;
 assign n_n4545 = ( wire317 ) | ( wire4735 ) | ( wire20134 ) ;
 assign n_n4548 = ( n_n4251 ) | ( wire878 ) | ( wire20119 ) ;
 assign n_n4549 = ( n_n4256 ) | ( n_n4255 ) | ( wire20122 ) ;
 assign wire54 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n281 ) ;
 assign wire609 = ( wire5439 ) | ( n_n128  &  n_n220  &  wire914 ) ;
 assign n_n2603 = ( n_n1  &  wire89 ) | ( n_n1  &  n_n83 ) | ( n_n1  &  wire19772 ) ;
 assign n_n2577 = ( wire5720 ) | ( wire5721 ) | ( wire19783 ) | ( wire19784 ) ;
 assign n_n2573 = ( n_n2579 ) | ( n_n2580 ) | ( wire19778 ) ;
 assign n_n2578 = ( n_n2860 ) | ( wire468 ) | ( wire5195 ) | ( wire19787 ) ;
 assign n_n2572 = ( n_n2577 ) | ( n_n2578 ) | ( wire19793 ) ;
 assign n_n2583 = ( n_n3786 ) | ( n_n3782 ) | ( wire19797 ) | ( wire19798 ) ;
 assign n_n2582 = ( wire806 ) | ( wire5171 ) | ( wire19802 ) | ( wire19803 ) ;
 assign wire1627 = ( wire268 ) | ( wire277 ) | ( n_n62 ) | ( wire101 ) ;
 assign n_n1709 = ( n_n1773 ) | ( wire21783 ) | ( wire21784 ) | ( wire21792 ) ;
 assign wire1630 = ( n_n44 ) | ( wire270 ) | ( wire21668 ) | ( wire21794 ) ;
 assign n_n1688 = ( n_n1710 ) | ( n_n1709 ) | ( wire3008 ) | ( wire21799 ) ;
 assign n_n1706 = ( wire2999 ) | ( wire3000 ) | ( wire21808 ) ;
 assign n_n1705 = ( n_n1761 ) | ( wire21813 ) | ( wire21814 ) | ( wire21817 ) ;
 assign n_n1687 = ( n_n1706 ) | ( n_n1705 ) | ( wire21825 ) ;
 assign n_n1711 = ( n_n1779 ) | ( wire2960 ) | ( wire2961 ) | ( wire21847 ) ;
 assign wire102 = ( (~ i_15_)  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n225 ) ;
 assign n_n1689 = ( n_n1713 ) | ( n_n1711 ) | ( wire21855 ) ;
 assign wire1637 = ( n_n221 ) | ( wire469 ) | ( wire22675 ) | ( wire22676 ) ;
 assign n_n758 = ( wire2063 ) | ( wire22678 ) | ( n_n6  &  wire1637 ) ;
 assign wire275 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n270 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n270 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n270 ) ;
 assign wire887 = ( n_n227  &  wire198 ) | ( n_n207  &  wire262 ) ;
 assign wire1640 = ( n_n228  &  wire902 ) | ( n_n228  &  wire912 ) ;
 assign wire1639 = ( wire898  &  n_n228 ) | ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign wire1638 = ( wire901  &  n_n228 ) | ( wire900  &  n_n228 ) ;
 assign wire1641 = ( n_n25 ) | ( wire145 ) | ( wire19457 ) | ( wire22687 ) ;
 assign n_n739 = ( n_n758 ) | ( wire22685 ) | ( wire22686 ) | ( wire22693 ) ;
 assign wire1645 = ( n_n78 ) | ( n_n26 ) | ( wire276 ) | ( wire65 ) ;
 assign wire1648 = ( n_n70 ) | ( n_n109 ) | ( wire143 ) | ( wire1649 ) ;
 assign wire1647 = ( n_n258  &  wire906 ) | ( n_n258  &  wire914 ) | ( n_n258  &  wire904 ) ;
 assign n_n4723 = ( n_n3398 ) | ( wire19930 ) | ( wire19931 ) | ( wire19946 ) ;
 assign n_n4744 = ( wire19959 ) | ( n_n130  &  wire19956 ) | ( n_n130  &  wire19957 ) ;
 assign n_n4725 = ( n_n4744 ) | ( wire19953 ) | ( wire19954 ) | ( wire19967 ) ;
 assign wire672 = ( n_n57  &  wire157 ) | ( n_n57  &  wire273 ) ;
 assign wire199 = ( i_15_  &  n_n228  &  n_n270 ) | ( (~ i_15_)  &  n_n258  &  n_n270 ) ;
 assign n_n3803 = ( n_n6  &  n_n7 ) | ( n_n5  &  wire199 ) ;
 assign n_n4544 = ( wire4726 ) | ( wire20141 ) | ( wire20142 ) ;
 assign n_n4551 = ( n_n4261 ) | ( wire721 ) | ( wire20224 ) ;
 assign n_n3708 = ( n_n4926 ) | ( wire693 ) | ( wire19537 ) ;
 assign n_n4535 = ( n_n3709 ) | ( n_n4551 ) | ( wire20228 ) | ( wire20232 ) ;
 assign wire1657 = ( wire82 ) | ( wire42 ) | ( n_n279  &  wire899 ) ;
 assign n_n3364 = ( n_n3380 ) | ( n_n3379 ) | ( wire20872 ) ;
 assign n_n3386 = ( n_n4807 ) | ( n_n4808 ) | ( wire3989 ) | ( wire20881 ) ;
 assign n_n3385 = ( wire3985 ) | ( wire20882 ) | ( wire20888 ) | ( wire20889 ) ;
 assign n_n2835 = ( n_n2926 ) | ( wire4365 ) | ( wire20508 ) ;
 assign wire1662 = ( wire123 ) | ( wire100 ) | ( wire227 ) | ( wire281 ) ;
 assign wire1661 = ( n_n112 ) | ( wire165 ) | ( wire167 ) | ( wire52 ) ;
 assign n_n707 = ( n_n94  &  n_n212 ) | ( n_n94  &  n_n200 ) | ( n_n94  &  n_n199 ) ;
 assign wire1664 = ( wire190 ) | ( wire124 ) | ( wire212 ) | ( wire119 ) ;
 assign n_n2656 = ( n_n2665 ) | ( wire4827 ) | ( wire20068 ) | ( wire20073 ) ;
 assign wire1668 = ( wire900  &  n_n220 ) | ( n_n220  &  wire912 ) | ( n_n220  &  wire897 ) ;
 assign n_n1724 = ( wire2906 ) | ( wire2907 ) | ( wire21888 ) | ( wire21889 ) ;
 assign wire426 = ( i_15_  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n222 ) ;
 assign wire134 = ( i_15_  &  n_n253  &  n_n225 ) | ( (~ i_15_)  &  n_n253  &  n_n225 ) ;
 assign wire544 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  n_n30 ) ;
 assign wire1669 = ( i_15_  &  n_n259  &  n_n225 ) | ( (~ i_15_)  &  n_n259  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign n_n755 = ( n_n785 ) | ( wire22792 ) | ( wire22793 ) ;
 assign wire1670 = ( wire911  &  n_n228 ) | ( n_n228  &  wire914 ) ;
 assign n_n756 = ( n_n809 ) | ( wire22803 ) | ( wire22804 ) | ( wire22809 ) ;
 assign n_n738 = ( n_n755 ) | ( n_n756 ) | ( wire22814 ) ;
 assign wire403 = ( wire903  &  n_n258 ) | ( n_n258  &  wire914 ) ;
 assign wire1673 = ( n_n258  &  wire905 ) | ( n_n258  &  wire908 ) ;
 assign n_n443 = ( n_n4183 ) | ( wire22451 ) | ( n_n53  &  wire41 ) ;
 assign wire175 = ( i_15_  &  n_n253  &  n_n256 ) | ( (~ i_15_)  &  n_n253  &  n_n256 ) ;
 assign wire1678 = ( n_n258  &  wire905 ) | ( n_n258  &  wire908 ) | ( n_n258  &  wire907 ) ;
 assign wire1677 = ( n_n258  &  wire914 ) | ( n_n258  &  wire908 ) ;
 assign wire1676 = ( wire913  &  n_n258 ) | ( wire903  &  n_n258 ) ;
 assign wire292 = ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire1682 = ( wire913  &  n_n258 ) | ( n_n258  &  wire914 ) | ( n_n258  &  wire908 ) ;
 assign wire1680 = ( n_n258  &  wire905 ) | ( n_n258  &  wire908 ) ;
 assign wire1679 = ( wire903  &  n_n258 ) | ( n_n258  &  wire907 ) ;
 assign wire1686 = ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) | ( n_n220  &  wire914 ) ;
 assign wire1687 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign n_n3637 = ( n_n1440 ) | ( wire5758 ) | ( wire19391 ) | ( wire19393 ) ;
 assign n_n3435 = ( wire20897 ) | ( n_n1  &  wire1877 ) ;
 assign n_n3383 = ( n_n3435 ) | ( wire20904 ) | ( wire20905 ) ;
 assign wire1693 = ( n_n110 ) | ( wire70 ) | ( n_n67 ) | ( wire19738 ) ;
 assign wire1696 = ( i_15_  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign n_n1738 = ( wire21652 ) | ( n_n268  &  wire212 ) | ( n_n268  &  wire1696 ) ;
 assign wire379 = ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire1699 = ( wire139 ) | ( wire19577 ) | ( n_n228  &  wire906 ) ;
 assign n_n741 = ( n_n834 ) | ( wire2011 ) | ( wire22714 ) | ( wire22717 ) ;
 assign n_n740 = ( n_n761 ) | ( n_n762 ) | ( wire22744 ) ;
 assign n_n732 = ( n_n738 ) | ( wire22763 ) | ( wire22764 ) | ( wire22822 ) ;
 assign wire1700 = ( n_n40 ) | ( wire233 ) | ( wire245 ) | ( wire351 ) ;
 assign wire1703 = ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) | ( n_n220  &  wire914 ) ;
 assign wire1707 = ( wire911  &  n_n281 ) | ( wire899  &  n_n281 ) | ( n_n281  &  wire912 ) ;
 assign wire1706 = ( wire911  &  n_n281 ) | ( wire899  &  n_n281 ) | ( n_n281  &  wire912 ) ;
 assign n_n3686 = ( wire5671 ) | ( wire19458 ) | ( n_n5  &  wire208 ) ;
 assign wire395 = ( n_n1  &  n_n29 ) | ( n_n1  &  wire49 ) | ( n_n1  &  wire88 ) ;
 assign n_n3642 = ( wire496 ) | ( wire812 ) | ( wire395 ) | ( wire19426 ) ;
 assign wire400 = ( wire130 ) | ( wire911  &  n_n228 ) ;
 assign wire1717 = ( wire911  &  n_n228 ) | ( n_n228  &  wire897 ) ;
 assign wire182 = ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign wire1723 = ( n_n132 ) | ( n_n260  &  n_n229  &  n_n165 ) ;
 assign wire132 = ( (~ i_15_)  &  n_n275  &  n_n281 ) | ( i_15_  &  n_n275  &  n_n220 ) ;
 assign wire236 = ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) | ( i_15_  &  n_n225  &  n_n270 ) ;
 assign wire1730 = ( wire74 ) | ( wire424 ) | ( wire903  &  n_n220 ) ;
 assign wire1732 = ( n_n25 ) | ( n_n24 ) | ( wire104 ) | ( wire228 ) ;
 assign wire123 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire1733 = ( wire124 ) | ( n_n258  &  wire897 ) ;
 assign wire1737 = ( wire903  &  n_n258 ) | ( n_n258  &  wire905 ) | ( n_n258  &  wire908 ) ;
 assign n_n431 = ( wire2384 ) | ( wire2385 ) | ( wire22403 ) | ( wire22404 ) ;
 assign wire1740 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign n_n3645 = ( wire19465 ) | ( wire19466 ) | ( wire19467 ) ;
 assign n_n3630 = ( n_n3395 ) | ( wire19511 ) | ( wire19512 ) | ( wire19523 ) ;
 assign wire1747 = ( wire165 ) | ( wire140 ) | ( wire198 ) | ( wire167 ) ;
 assign wire225 = ( i_15_  &  n_n242  &  n_n228 ) | ( (~ i_15_)  &  n_n242  &  n_n258 ) ;
 assign wire1753 = ( wire901  &  n_n228 ) | ( wire898  &  n_n228 ) | ( n_n228  &  wire902 ) ;
 assign wire1752 = ( wire901  &  n_n228 ) | ( wire898  &  n_n228 ) | ( n_n228  &  wire912 ) ;
 assign wire1755 = ( (~ i_15_)  &  n_n253  &  n_n279 ) | ( i_15_  &  n_n253  &  n_n256 ) | ( (~ i_15_)  &  n_n253  &  n_n256 ) ;
 assign n_n2671 = ( wire548 ) | ( wire434 ) | ( wire20075 ) | ( wire20076 ) ;
 assign n_n2657 = ( wire20094 ) | ( wire20095 ) ;
 assign n_n2659 = ( wire493 ) | ( n_n2673 ) | ( wire20103 ) | ( wire20104 ) ;
 assign wire1768 = ( n_n221 ) | ( n_n71 ) | ( wire143 ) | ( wire375 ) ;
 assign n_n1761 = ( wire2994 ) | ( n_n5  &  wire1768 ) ;
 assign n_n1773 = ( wire679 ) | ( wire3018 ) | ( wire3019 ) | ( wire21786 ) ;
 assign wire1773 = ( wire901  &  n_n220 ) | ( wire899  &  n_n220 ) | ( wire902  &  n_n220 ) ;
 assign wire1772 = ( wire902  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire1771 = ( wire911  &  n_n220 ) | ( n_n220  &  wire897 ) ;
 assign wire1776 = ( i_8_  &  n_n272  &  n_n230  &  n_n285 ) | ( (~ i_8_)  &  n_n272  &  n_n230  &  n_n285 ) ;
 assign wire1777 = ( n_n228  &  wire902 ) | ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign n_n775 = ( wire510 ) | ( wire511 ) | ( wire22829 ) | ( wire22830 ) ;
 assign n_n4542 = ( wire4710 ) | ( wire20152 ) | ( wire20153 ) ;
 assign n_n4541 = ( wire4704 ) | ( wire4705 ) | ( wire20157 ) ;
 assign wire1786 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign n_n2433 = ( wire481 ) | ( wire589 ) | ( wire3578 ) | ( wire3579 ) ;
 assign n_n1753 = ( wire21675 ) | ( wire21676 ) | ( wire21677 ) | ( wire21678 ) ;
 assign wire622 = ( n_n4  &  n_n107 ) | ( n_n4  &  n_n220  &  wire905 ) ;
 assign wire1793 = ( n_n71 ) | ( n_n44 ) | ( wire143 ) | ( wire21668 ) ;
 assign wire143 = ( (~ i_15_)  &  n_n222  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n256 ) ;
 assign wire1794 = ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n256 ) ;
 assign wire1795 = ( n_n109 ) | ( n_n44 ) | ( wire143 ) | ( wire22341 ) ;
 assign n_n341 = ( n_n359 ) | ( wire22572 ) | ( wire22573 ) | ( wire22581 ) ;
 assign wire1797 = ( n_n279  &  wire913 ) | ( n_n279  &  wire905 ) | ( n_n279  &  wire914 ) ;
 assign wire1796 = ( n_n260  &  n_n229  &  n_n165 ) | ( n_n260  &  n_n283  &  n_n165 ) ;
 assign n_n3658 = ( n_n4682 ) | ( n_n4685 ) | ( wire19565 ) | ( wire19566 ) ;
 assign wire117 = ( wire66 ) | ( n_n222  &  wire905 ) ;
 assign wire1803 = ( (~ i_15_)  &  n_n222  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n225 ) ;
 assign n_n1692 = ( wire21864 ) | ( wire21865 ) | ( wire21874 ) | ( wire21877 ) ;
 assign n_n2673 = ( n_n3598 ) | ( wire380 ) | ( wire471 ) | ( wire20096 ) ;
 assign wire1807 = ( n_n10 ) | ( n_n63 ) | ( wire113 ) | ( wire199 ) ;
 assign n_n2431 = ( wire3572 ) | ( wire3576 ) | ( wire3577 ) | ( wire21330 ) ;
 assign wire1812 = ( n_n99 ) | ( n_n52 ) | ( wire807 ) | ( wire226 ) ;
 assign wire1814 = ( n_n197 ) | ( wire42 ) | ( wire275 ) | ( wire441 ) ;
 assign wire1813 = ( n_n216 ) | ( wire190 ) | ( wire292 ) | ( wire52 ) ;
 assign wire167 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire908 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire908 ) ;
 assign wire1819 = ( n_n93 ) | ( n_n90 ) | ( wire76 ) | ( wire19384 ) ;
 assign wire1825 = ( n_n281  &  wire914 ) | ( n_n281  &  wire907 ) ;
 assign n_n4539 = ( wire4684 ) | ( wire4685 ) | ( wire20176 ) ;
 assign wire1829 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n118 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n118 ) ;
 assign n_n4464 = ( wire3720 ) | ( wire21168 ) | ( n_n127  &  wire1843 ) ;
 assign wire879 = ( (~ i_7_)  &  i_6_  &  wire936 ) | ( i_7_  &  (~ i_6_)  &  wire936 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire936 ) | ( i_7_  &  i_6_  &  wire929 ) | ( (~ i_7_)  &  i_6_  &  wire929 ) | ( i_7_  &  (~ i_6_)  &  wire929 ) ;
 assign n_n2428 = ( wire3558 ) | ( wire21350 ) | ( wire21352 ) ;
 assign wire1835 = ( n_n34 ) | ( wire154 ) | ( wire236 ) | ( wire362 ) ;
 assign wire1837 = ( n_n203 ) | ( wire161 ) | ( wire20149 ) | ( wire22835 ) ;
 assign wire1836 = ( n_n221 ) | ( wire469 ) | ( wire128 ) | ( wire22833 ) ;
 assign wire1845 = ( wire54 ) | ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire1843 = ( wire48 ) | ( n_n110 ) | ( n_n111 ) | ( wire54 ) ;
 assign wire1842 = ( n_n132 ) | ( n_n229  &  n_n165  &  n_n284 ) ;
 assign wire1849 = ( (~ i_15_)  &  n_n222  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n225 ) ;
 assign wire43 = ( wire19385 ) | ( wire900  &  n_n256 ) ;
 assign wire807 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) ;
 assign wire47 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire907 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire907 ) ;
 assign wire52 = ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n228 ) ;
 assign wire53 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire57 = ( (~ i_15_)  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n247  &  n_n228 ) ;
 assign wire58 = ( wire19575 ) | ( wire898  &  n_n225 ) ;
 assign wire59 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire61 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) ;
 assign wire63 = ( (~ i_15_)  &  n_n258  &  n_n270 ) | ( i_15_  &  n_n220  &  n_n270 ) ;
 assign wire64 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire901 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign wire65 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire71 = ( i_15_  &  n_n253  &  n_n281 ) | ( (~ i_15_)  &  n_n253  &  n_n225 ) ;
 assign wire74 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire76 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) ;
 assign wire83 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire84 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) ;
 assign wire86 = ( i_15_  &  n_n281  &  n_n282 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire87 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire245 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n256 ) ;
 assign wire95 = ( (~ i_15_)  &  n_n247  &  n_n258 ) | ( i_15_  &  n_n247  &  n_n220 ) ;
 assign wire96 = ( i_15_  &  n_n253  &  n_n279 ) | ( (~ i_15_)  &  n_n253  &  n_n228 ) ;
 assign wire97 = ( wire514 ) | ( wire911  &  n_n225 ) ;
 assign wire100 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire103 = ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n281  &  n_n259 ) ;
 assign wire104 = ( (~ i_15_)  &  n_n275  &  n_n222 ) | ( i_15_  &  n_n275  &  n_n225 ) ;
 assign wire105 = ( wire20155 ) | ( wire913  &  n_n225 ) ;
 assign wire453 = ( i_15_  &  n_n247  &  n_n281 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign wire110 = ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire128 = ( i_15_  &  n_n259  &  n_n225 ) | ( (~ i_15_)  &  n_n259  &  n_n225 ) ;
 assign wire130 = ( (~ i_15_)  &  n_n242  &  n_n281 ) | ( i_15_  &  n_n242  &  n_n220 ) ;
 assign wire145 = ( i_15_  &  n_n247  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign wire288 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) ;
 assign wire148 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire149 = ( wire21389 ) | ( n_n281  &  wire900 ) ;
 assign wire152 = ( i_13_  &  (~ i_12_) ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire161 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) ;
 assign wire187 = ( i_15_  &  n_n259  &  n_n256 ) | ( (~ i_15_)  &  n_n259  &  n_n256 ) ;
 assign wire195 = ( i_15_  &  n_n242  &  n_n281 ) | ( (~ i_15_)  &  n_n242  &  n_n220 ) ;
 assign wire196 = ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire197 = ( i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire202 = ( wire96 ) | ( n_n222  &  wire898 ) ;
 assign wire203 = ( wire104 ) | ( n_n279  &  wire903 ) ;
 assign wire210 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) ;
 assign wire214 = ( i_14_  &  n_n278  &  n_n259 ) | ( (~ i_14_)  &  i_15_  &  n_n278  &  n_n259 ) ;
 assign wire215 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire220 = ( (~ i_15_)  &  n_n253  &  n_n258 ) | ( i_15_  &  n_n253  &  n_n220 ) ;
 assign wire226 = ( i_15_  &  n_n253  &  n_n281 ) | ( (~ i_15_)  &  n_n253  &  n_n220 ) ;
 assign wire227 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire228 = ( i_15_  &  n_n275  &  n_n281 ) | ( (~ i_15_)  &  n_n275  &  n_n220 ) ;
 assign wire229 = ( i_15_  &  n_n267  &  n_n256 ) | ( (~ i_15_)  &  n_n267  &  n_n256 ) ;
 assign wire230 = ( i_15_  &  n_n281  &  n_n270 ) | ( (~ i_15_)  &  n_n220  &  n_n270 ) ;
 assign wire231 = ( i_15_  &  n_n275  &  n_n256 ) | ( (~ i_15_)  &  n_n275  &  n_n256 ) ;
 assign wire232 = ( (~ i_15_)  &  n_n242  &  n_n228 ) | ( i_15_  &  n_n242  &  n_n258 ) ;
 assign wire235 = ( i_15_  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n279  &  n_n270 ) | ( i_15_  &  n_n281  &  n_n270 ) ;
 assign wire375 = ( i_15_  &  n_n281  &  n_n259 ) | ( (~ i_15_)  &  n_n259  &  n_n220 ) ;
 assign wire240 = ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n225 ) ;
 assign wire241 = ( i_15_  &  n_n279  &  n_n267 ) | ( (~ i_15_)  &  n_n279  &  n_n267 ) | ( i_15_  &  n_n281  &  n_n267 ) ;
 assign wire242 = ( i_15_  &  n_n253  &  n_n279 ) | ( (~ i_15_)  &  n_n253  &  n_n279 ) | ( i_15_  &  n_n253  &  n_n281 ) ;
 assign wire243 = ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) ;
 assign wire246 = ( i_15_  &  n_n228  &  n_n267 ) | ( (~ i_15_)  &  n_n258  &  n_n267 ) ;
 assign wire256 = ( (~ i_15_)  &  n_n281  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign wire262 = ( (~ i_14_)  &  i_15_  &  n_n275  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n275  &  n_n254 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n275  &  n_n254 ) ;
 assign wire263 = ( i_15_  &  n_n247  &  n_n281 ) | ( (~ i_15_)  &  n_n247  &  n_n220 ) ;
 assign wire266 = ( (~ i_9_)  &  (~ i_10_) ) | ( n_n220  &  wire905 ) ;
 assign wire270 = ( i_15_  &  n_n281  &  n_n267 ) | ( (~ i_15_)  &  n_n220  &  n_n267 ) ;
 assign wire274 = ( i_15_  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n222  &  n_n259 ) | ( (~ i_15_)  &  n_n259  &  n_n228 ) ;
 assign wire281 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) ;
 assign wire282 = ( wire19238 ) | ( n_n281  &  wire914 ) ;
 assign wire285 = ( wire19253 ) | ( n_n279  &  wire912 ) ;
 assign wire287 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire291 = ( (~ i_15_)  &  n_n258  &  n_n282 ) | ( i_15_  &  n_n220  &  n_n282 ) ;
 assign wire294 = ( wire103 ) | ( n_n220  &  wire914 ) ;
 assign wire1852 = ( n_n29 ) | ( n_n101 ) | ( wire88 ) | ( wire61 ) ;
 assign wire299 = ( wire54 ) | ( n_n220  &  wire914 ) ;
 assign wire304 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n247 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n247 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n247 ) ;
 assign wire305 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n259 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n259 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n259 ) ;
 assign wire306 = ( (~ i_15_)  &  n_n259  &  n_n228 ) | ( i_15_  &  n_n259  &  n_n258 ) ;
 assign wire310 = ( n_n228  &  wire912 ) | ( n_n228  &  wire897 ) ;
 assign wire311 = ( i_15_  &  n_n253  &  n_n222 ) | ( (~ i_15_)  &  n_n253  &  n_n222 ) | ( (~ i_15_)  &  n_n253  &  n_n228 ) ;
 assign wire1853 = ( n_n113 ) | ( n_n85 ) | ( wire102 ) | ( wire87 ) ;
 assign wire321 = ( n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n281 ) ;
 assign wire325 = ( i_15_  &  n_n242  &  n_n281 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire328 = ( i_9_  &  i_10_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign wire331 = ( wire196 ) | ( i_13_  &  (~ i_12_)  &  n_n247 ) ;
 assign wire338 = ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n281  &  n_n259 ) ;
 assign wire342 = ( i_15_  &  n_n247  &  n_n281 ) | ( i_15_  &  n_n247  &  n_n256 ) | ( (~ i_15_)  &  n_n247  &  n_n256 ) ;
 assign wire343 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n228 ) ;
 assign wire345 = ( i_15_  &  n_n275  &  n_n281 ) | ( i_15_  &  n_n275  &  n_n256 ) | ( (~ i_15_)  &  n_n275  &  n_n256 ) ;
 assign wire346 = ( i_15_  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n228 ) ;
 assign wire347 = ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n247  &  n_n228 ) ;
 assign wire348 = ( (~ i_14_)  &  i_15_  &  n_n254  &  n_n242 ) | ( i_14_  &  (~ i_15_)  &  n_n254  &  n_n242 ) | ( (~ i_14_)  &  (~ i_15_)  &  n_n254  &  n_n242 ) ;
 assign wire351 = ( (~ i_15_)  &  n_n247  &  n_n228 ) | ( i_15_  &  n_n247  &  n_n258 ) ;
 assign wire352 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire357 = ( (~ i_15_)  &  n_n253  &  n_n228 ) | ( i_15_  &  n_n253  &  n_n258 ) ;
 assign wire358 = ( i_15_  &  n_n247  &  n_n256 ) | ( (~ i_15_)  &  n_n247  &  n_n256 ) ;
 assign wire361 = ( i_15_  &  n_n253  &  n_n222 ) | ( (~ i_15_)  &  n_n253  &  n_n222 ) | ( i_15_  &  n_n253  &  n_n225 ) ;
 assign wire362 = ( i_15_  &  n_n222  &  n_n282 ) | ( (~ i_15_)  &  n_n222  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n225 ) ;
 assign wire363 = ( wire226 ) | ( wire898  &  n_n256 ) ;
 assign wire1855 = ( n_n80 ) | ( n_n28 ) | ( wire88 ) | ( wire65 ) ;
 assign wire1856 = ( n_n26 ) | ( n_n101 ) | ( wire80 ) | ( wire61 ) ;
 assign wire397 = ( wire215 ) | ( n_n242  &  n_n222 ) ;
 assign wire398 = ( wire130 ) | ( n_n279  &  wire911 ) ;
 assign wire399 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n242  &  n_n281 ) ;
 assign wire405 = ( (~ i_15_)  &  n_n275  &  n_n279 ) | ( i_15_  &  n_n275  &  n_n256 ) | ( (~ i_15_)  &  n_n275  &  n_n256 ) ;
 assign wire413 = ( i_15_  &  n_n279  &  n_n259 ) | ( (~ i_15_)  &  n_n279  &  n_n259 ) ;
 assign wire414 = ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( i_15_  &  n_n256  &  n_n282 ) | ( (~ i_15_)  &  n_n256  &  n_n282 ) ;
 assign wire419 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire914 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire914 ) ;
 assign wire424 = ( i_15_  &  n_n275  &  n_n222 ) | ( (~ i_15_)  &  n_n275  &  n_n222 ) | ( i_15_  &  n_n275  &  n_n225 ) ;
 assign wire428 = ( i_15_  &  n_n222  &  n_n247 ) | ( (~ i_15_)  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n225 ) ;
 assign wire431 = ( i_15_  &  n_n281  &  n_n270 ) | ( i_15_  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n256  &  n_n270 ) ;
 assign wire433 = ( i_15_  &  n_n222  &  n_n282 ) | ( (~ i_15_)  &  n_n222  &  n_n282 ) | ( (~ i_15_)  &  n_n228  &  n_n282 ) ;
 assign wire435 = ( n_n143 ) | ( wire214 ) ;
 assign wire436 = ( i_15_  &  n_n279  &  n_n282 ) | ( (~ i_15_)  &  n_n279  &  n_n282 ) | ( i_15_  &  n_n281  &  n_n282 ) ;
 assign wire437 = ( i_15_  &  n_n281  &  n_n282 ) | ( i_15_  &  n_n256  &  n_n282 ) | ( (~ i_15_)  &  n_n256  &  n_n282 ) ;
 assign wire440 = ( wire44 ) | ( wire900  &  n_n228 ) ;
 assign wire441 = ( (~ i_15_)  &  n_n279  &  n_n259 ) | ( i_15_  &  n_n259  &  n_n256 ) | ( (~ i_15_)  &  n_n259  &  n_n256 ) ;
 assign wire444 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n256 ) | ( (~ i_15_)  &  n_n247  &  n_n256 ) ;
 assign wire448 = ( i_15_  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n222  &  n_n267 ) | ( (~ i_15_)  &  n_n228  &  n_n267 ) ;
 assign wire454 = ( wire215 ) | ( i_13_  &  (~ i_12_)  &  n_n242 ) ;
 assign wire1868 = ( wire88 ) | ( n_n222  &  wire902 ) | ( wire902  &  n_n258 ) ;
 assign wire1871 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire1873 = ( wire71 ) | ( n_n220  &  wire904 ) | ( n_n256  &  wire904 ) ;
 assign wire1874 = ( n_n228  &  wire912 ) | ( n_n281  &  wire907 ) ;
 assign wire1877 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire1878 = ( n_n44 ) | ( n_n90 ) | ( wire19384 ) | ( wire19385 ) ;
 assign wire1884 = ( n_n179 ) | ( n_n81 ) | ( wire57 ) | ( wire86 ) ;
 assign wire1891 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire1892 = ( n_n93 ) | ( n_n44 ) | ( wire76 ) | ( wire19385 ) ;
 assign wire1893 = ( n_n204 ) | ( n_n112 ) | ( wire52 ) | ( wire84 ) ;
 assign wire1894 = ( wire89 ) | ( n_n35 ) | ( n_n83 ) | ( wire64 ) ;
 assign wire1896 = ( wire69 ) | ( wire80 ) | ( wire902  &  n_n256 ) ;
 assign wire1897 = ( wire44 ) | ( n_n15 ) | ( n_n258  &  wire904 ) ;
 assign wire1898 = ( n_n70 ) | ( n_n20 ) | ( wire79 ) | ( wire66 ) ;
 assign wire1899 = ( n_n26 ) | ( n_n101 ) | ( wire80 ) | ( wire61 ) ;
 assign wire1900 = ( wire89 ) | ( n_n35 ) | ( n_n83 ) | ( wire64 ) ;
 assign wire1902 = ( n_n179 ) | ( n_n39 ) | ( wire57 ) | ( wire245 ) ;
 assign wire1903 = ( n_n200 ) | ( n_n23 ) | ( wire74 ) | ( wire104 ) ;
 assign wire1904 = ( n_n200 ) | ( n_n23 ) | ( wire74 ) | ( wire104 ) ;
 assign wire1905 = ( n_n99 ) | ( n_n51 ) | ( wire96 ) | ( wire19575 ) ;
 assign wire1910 = ( n_n221 ) | ( wire469 ) | ( n_n72 ) | ( wire66 ) ;
 assign wire1914 = ( n_n97 ) | ( n_n51 ) | ( wire71 ) | ( wire19575 ) ;
 assign wire1916 = ( n_n44 ) | ( n_n90 ) | ( wire19384 ) | ( wire19385 ) ;
 assign wire1917 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire1918 = ( wire88 ) | ( n_n222  &  wire902 ) | ( wire902  &  n_n258 ) ;
 assign wire1920 = ( n_n24 ) | ( n_n73 ) | ( wire19407 ) | ( wire19408 ) ;
 assign wire1923 = ( n_n70 ) | ( n_n20 ) | ( wire79 ) | ( wire66 ) ;
 assign wire1924 = ( n_n93 ) | ( n_n44 ) | ( wire76 ) | ( wire19385 ) ;
 assign wire1926 = ( n_n221 ) | ( wire469 ) | ( n_n72 ) | ( wire66 ) ;
 assign wire1927 = ( n_n37 ) | ( wire89 ) | ( n_n82 ) | ( wire47 ) ;
 assign wire1928 = ( n_n99 ) | ( n_n51 ) | ( wire96 ) | ( wire19575 ) ;
 assign wire1932 = ( n_n223 ) | ( n_n20 ) | ( wire42 ) | ( wire66 ) ;
 assign wire1936 = ( wire166 ) | ( wire180 ) ;
 assign wire1937 = ( n_n29 ) | ( n_n101 ) | ( wire88 ) | ( wire61 ) ;
 assign wire1938 = ( n_n223 ) | ( n_n20 ) | ( wire42 ) | ( wire66 ) ;
 assign wire1939 = ( n_n28 ) | ( n_n78 ) | ( wire80 ) | ( wire65 ) ;
 assign wire1940 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire1943 = ( n_n99 ) | ( n_n51 ) | ( wire96 ) | ( wire19575 ) ;
 assign wire1945 = ( n_n38 ) | ( n_n39 ) | ( wire245 ) | ( wire453 ) ;
 assign wire1946 = ( n_n221 ) | ( wire469 ) | ( n_n72 ) | ( wire66 ) ;
 assign wire1948 = ( n_n24 ) | ( n_n73 ) | ( wire19407 ) | ( wire19408 ) ;
 assign wire1950 = ( wire89 ) | ( n_n35 ) | ( n_n83 ) | ( wire64 ) ;
 assign wire1951 = ( n_n204 ) | ( n_n112 ) | ( wire52 ) | ( wire84 ) ;
 assign wire1952 = ( n_n111 ) | ( n_n108 ) | ( wire54 ) | ( wire103 ) ;
 assign wire1953 = ( wire56 ) | ( wire53 ) | ( n_n279  &  wire897 ) ;
 assign wire857 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n225 ) ;
 assign wire858 = ( i_15_  &  n_n275  &  n_n279 ) | ( (~ i_15_)  &  n_n275  &  n_n279 ) | ( i_15_  &  n_n275  &  n_n281 ) ;
 assign wire1959 = ( n_n29 ) | ( n_n101 ) | ( wire88 ) | ( wire61 ) ;
 assign wire962 = ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire966 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire965 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire969 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire968 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire971 = ( (~ i_12_) ) | ( i_13_  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign wire1037 = ( n_n84 ) | ( n_n35 ) | ( wire78 ) | ( wire86 ) ;
 assign wire1074 = ( i_13_  &  (~ i_12_) ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1101 = ( n_n281  &  wire914 ) | ( n_n281  &  wire904 ) | ( n_n281  &  wire907 ) ;
 assign wire1124 = ( n_n89 ) | ( n_n44 ) | ( wire408 ) | ( wire22341 ) ;
 assign wire1131 = ( (~ i_13_) ) | ( (~ i_12_) ) | ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign wire1133 = ( (~ i_14_)  &  i_13_  &  i_12_ ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1135 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1183 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1182 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire1199 = ( wire900  &  n_n220 ) | ( wire898  &  n_n220 ) ;
 assign wire1214 = ( wire514 ) | ( wire232 ) | ( wire911  &  n_n256 ) ;
 assign wire1225 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire1317 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) ;
 assign wire1501 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire1508 = ( wire48 ) | ( wire62 ) | ( n_n204 ) | ( n_n16 ) ;
 assign wire1529 = ( wire40 ) | ( wire21367 ) | ( n_n281  &  wire897 ) ;
 assign wire1554 = ( wire124 ) | ( wire212 ) | ( wire119 ) ;
 assign wire1619 = ( n_n112 ) | ( wire247 ) | ( wire52 ) | ( wire210 ) ;
 assign wire1649 = ( n_n258  &  wire906 ) | ( n_n258  &  wire904 ) ;
 assign wire1652 = ( n_n17 ) | ( n_n67 ) | ( wire514 ) | ( wire232 ) ;
 assign wire1656 = ( n_n204 ) | ( n_n67 ) | ( wire52 ) | ( wire19738 ) ;
 assign wire1705 = ( wire913  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire1781 = ( n_n16 ) | ( n_n68 ) | ( wire514 ) | ( wire20155 ) ;
 assign wire1792 = ( n_n17 ) | ( wire195 ) | ( wire240 ) | ( wire857 ) ;
 assign wire1822 = ( wire84 ) | ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) ;
 assign wire238 = ( n_n3  &  wire368 ) | ( n_n3  &  n_n88 ) | ( n_n3  &  wire22841 ) ;
 assign wire505 = ( wire169  &  wire901  &  n_n228 ) ;
 assign wire510 = ( n_n229  &  n_n285  &  n_n284  &  wire1777 ) ;
 assign wire511 = ( wire169  &  wire911  &  n_n228 ) ;
 assign wire529 = ( n_n3  &  n_n46 ) | ( n_n3  &  wire19577 ) | ( n_n3  &  wire22816 ) ;
 assign wire543 = ( n_n1  &  wire254 ) | ( n_n1  &  wire356 ) ;
 assign wire550 = ( wire224  &  n_n260  &  n_n283  &  n_n285 ) ;
 assign wire564 = ( n_n260  &  n_n263  &  n_n285  &  wire1670 ) ;
 assign wire580 = ( n_n227  &  wire22795 ) | ( n_n227  &  n_n228  &  wire897 ) ;
 assign wire608 = ( i_15_  &  n_n3  &  n_n253  &  n_n225 ) | ( (~ i_15_)  &  n_n3  &  n_n253  &  n_n225 ) ;
 assign wire847 = ( n_n2  &  wire227 ) | ( n_n2  &  wire305 ) ;
 assign wire850 = ( n_n268  &  wire20362 ) | ( n_n268  &  n_n279  &  wire897 ) ;
 assign wire855 = ( n_n268  &  wire368 ) | ( n_n268  &  n_n39 ) | ( n_n268  &  wire55 ) ;
 assign wire856 = ( n_n265  &  wire89 ) | ( n_n265  &  wire22772 ) ;
 assign wire862 = ( n_n4  &  n_n99 ) | ( n_n4  &  n_n54 ) | ( n_n4  &  wire96 ) ;
 assign wire895 = ( n_n268  &  wire310 ) | ( n_n268  &  wire22769 ) ;
 assign wire1964 = ( n_n2  &  wire262 ) | ( n_n2  &  wire304 ) | ( n_n2  &  wire22758 ) ;
 assign wire1968 = ( n_n1  &  wire224 ) | ( n_n1  &  wire335 ) | ( n_n1  &  wire22754 ) ;
 assign wire1969 = ( n_n2  &  wire277 ) | ( n_n2  &  wire356 ) | ( n_n2  &  wire22757 ) ;
 assign wire1970 = ( n_n2  &  wire275 ) | ( n_n2  &  wire348 ) | ( n_n2  &  wire22748 ) ;
 assign wire1971 = ( n_n1  &  wire262 ) | ( n_n1  &  wire305 ) | ( n_n1  &  wire22752 ) ;
 assign wire1975 = ( n_n3  &  wire134 ) | ( n_n3  &  wire901  &  n_n258 ) ;
 assign wire1976 = ( n_n4  &  wire368 ) | ( n_n4  &  n_n88 ) | ( n_n4  &  wire22746 ) ;
 assign wire1977 = ( n_n6  &  n_n41 ) | ( n_n6  &  wire139 ) | ( n_n6  &  wire145 ) ;
 assign wire1978 = ( n_n5  &  n_n104 ) | ( n_n5  &  wire134 ) | ( n_n5  &  wire22740 ) ;
 assign wire1984 = ( wire126  &  n_n6 ) | ( n_n6  &  n_n37 ) | ( n_n6  &  wire89 ) ;
 assign wire1990 = ( n_n53  &  wire161 ) | ( n_n53  &  wire22730 ) ;
 assign wire1997 = ( n_n48  &  n_n228  &  wire902 ) ;
 assign wire2001 = ( n_n99  &  n_n6 ) | ( n_n6  &  wire134 ) | ( n_n6  &  wire96 ) ;
 assign wire2002 = ( n_n5  &  n_n46 ) | ( n_n5  &  wire19577 ) | ( n_n5  &  wire22719 ) ;
 assign wire2008 = ( n_n48  &  wire304 ) | ( n_n48  &  n_n279  &  wire912 ) ;
 assign wire2011 = ( n_n48  &  wire1699 ) | ( n_n48  &  wire22711 ) ;
 assign wire2012 = ( n_n53  &  n_n46 ) | ( n_n53  &  wire139 ) | ( n_n53  &  wire19577 ) ;
 assign wire2019 = ( n_n53  &  wire368 ) | ( n_n53  &  n_n88 ) | ( n_n53  &  wire145 ) ;
 assign wire2022 = ( n_n264  &  n_n283  &  n_n285  &  wire1343 ) ;
 assign wire2023 = ( i_15_  &  n_n53  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n53  &  n_n282  &  n_n225 ) ;
 assign wire2030 = ( n_n48  &  wire120 ) | ( n_n48  &  n_n25 ) | ( n_n48  &  wire19457 ) ;
 assign wire2034 = ( n_n53  &  n_n203 ) | ( n_n53  &  wire128 ) | ( n_n53  &  wire20149 ) ;
 assign wire2035 = ( n_n48  &  n_n203 ) | ( n_n48  &  wire20149 ) | ( n_n48  &  wire22696 ) ;
 assign wire2041 = ( n_n53  &  wire120 ) | ( n_n53  &  n_n25 ) | ( n_n53  &  wire19457 ) ;
 assign wire2059 = ( n_n208  &  n_n230  &  n_n285  &  wire190 ) ;
 assign wire2063 = ( n_n5  &  wire114 ) | ( n_n5  &  n_n216 ) | ( n_n5  &  wire22674 ) ;
 assign wire2067 = ( n_n5  &  n_n203 ) | ( n_n5  &  wire161 ) | ( n_n5  &  wire20149 ) ;
 assign wire2072 = ( n_n99  &  n_n100 ) | ( n_n100  &  wire96 ) | ( n_n100  &  wire22664 ) ;
 assign wire2081 = ( n_n260  &  n_n261  &  n_n285  &  wire1340 ) ;
 assign wire2082 = ( n_n37  &  n_n94 ) | ( wire89  &  n_n94 ) | ( n_n94  &  wire22657 ) ;
 assign wire2089 = ( n_n99  &  n_n94 ) | ( n_n94  &  wire134 ) | ( n_n94  &  wire96 ) ;
 assign wire2091 = ( n_n100  &  n_n80 ) | ( n_n100  &  wire114 ) | ( n_n100  &  wire88 ) ;
 assign wire2092 = ( n_n94  &  n_n25 ) | ( n_n94  &  wire19457 ) | ( n_n94  &  wire22650 ) ;
 assign wire2103 = ( n_n57  &  wire275 ) | ( n_n57  &  wire262 ) ;
 assign wire2104 = ( n_n56  &  wire198 ) | ( n_n56  &  wire262 ) | ( n_n56  &  wire304 ) ;
 assign wire2122 = ( n_n99  &  n_n53 ) | ( n_n53  &  wire96 ) | ( n_n53  &  wire22631 ) ;
 assign wire2126 = ( n_n56  &  wire275 ) | ( n_n56  &  wire22629 ) | ( n_n56  &  wire22630 ) ;
 assign wire2127 = ( n_n57  &  wire305 ) | ( n_n57  &  wire348 ) | ( n_n57  &  wire22629 ) ;
 assign wire2128 = ( n_n56  &  wire301 ) | ( n_n56  &  wire356 ) ;
 assign wire2129 = ( n_n57  &  wire301 ) | ( n_n57  &  wire335 ) | ( n_n57  &  wire304 ) ;
 assign wire2138 = ( n_n230  &  n_n271  &  n_n285  &  wire335 ) ;
 assign wire2162 = ( n_n4  &  wire128 ) | ( n_n4  &  wire911  &  n_n258 ) ;
 assign wire2163 = ( n_n3  &  wire22598 ) | ( n_n3  &  wire22599 ) ;
 assign wire2168 = ( n_n3  &  wire120 ) | ( n_n3  &  wire902  &  n_n258 ) ;
 assign wire2169 = ( n_n4  &  n_n25 ) | ( n_n4  &  wire19457 ) | ( n_n4  &  wire22597 ) ;
 assign wire2170 = ( n_n3  &  n_n25 ) | ( n_n3  &  n_n103 ) | ( n_n3  &  wire19457 ) ;
 assign wire2173 = ( n_n3  &  wire126 ) | ( n_n3  &  n_n37 ) | ( n_n3  &  wire89 ) ;
 assign wire2174 = ( n_n4  &  n_n37 ) | ( n_n4  &  wire89 ) | ( n_n4  &  n_n104 ) ;
 assign wire2176 = ( wire169  &  wire913  &  n_n258 ) ;
 assign wire2183 = ( n_n208  &  n_n285  &  n_n284  &  wire1795 ) ;
 assign wire2196 = ( n_n197  &  n_n227 ) | ( n_n227  &  wire42 ) | ( n_n227  &  wire441 ) ;
 assign wire2200 = ( n_n207  &  n_n212 ) | ( n_n207  &  n_n216 ) | ( n_n207  &  wire52 ) ;
 assign wire2205 = ( n_n4  &  wire65 ) | ( n_n4  &  wire902  &  n_n256 ) ;
 assign wire2206 = ( wire913  &  n_n258  &  wire278 ) ;
 assign wire2225 = ( n_n2  &  wire187 ) | ( n_n2  &  n_n258  &  wire904 ) ;
 assign wire2235 = ( wire1354  &  wire123 ) | ( wire899  &  n_n258  &  wire1354 ) ;
 assign wire2237 = ( n_n1  &  n_n112 ) | ( n_n1  &  wire52 ) | ( n_n1  &  wire110 ) ;
 assign wire2239 = ( n_n1  &  wire187 ) | ( n_n1  &  wire911  &  n_n258 ) ;
 assign wire2240 = ( n_n2  &  n_n112 ) | ( n_n2  &  wire52 ) | ( n_n2  &  wire22535 ) ;
 assign wire2243 = ( n_n268  &  wire403 ) | ( n_n268  &  wire292 ) | ( n_n268  &  wire22531 ) ;
 assign wire2246 = ( n_n1  &  wire175 ) | ( n_n1  &  wire900  &  n_n258 ) ;
 assign wire2258 = ( n_n2  &  n_n34 ) | ( n_n2  &  wire47 ) | ( n_n2  &  wire22519 ) ;
 assign wire2260 = ( n_n1  &  wire124 ) | ( n_n1  &  wire22515 ) | ( n_n1  &  wire22516 ) ;
 assign wire2263 = ( n_n1  &  wire140 ) | ( n_n1  &  wire182 ) ;
 assign wire2264 = ( n_n2  &  wire41 ) | ( n_n2  &  wire175 ) | ( n_n2  &  wire22506 ) ;
 assign wire2265 = ( n_n1  &  wire166 ) | ( n_n1  &  wire358 ) | ( n_n1  &  wire22510 ) ;
 assign wire2267 = ( n_n2  &  wire112 ) | ( n_n2  &  wire144 ) ;
 assign wire2268 = ( n_n1  &  wire112 ) | ( n_n1  &  wire901  &  n_n258 ) ;
 assign wire2269 = ( n_n94  &  n_n104 ) | ( n_n94  &  n_n113 ) | ( n_n94  &  wire57 ) ;
 assign wire2277 = ( i_15_  &  n_n94  &  n_n256  &  n_n282 ) | ( (~ i_15_)  &  n_n94  &  n_n256  &  n_n282 ) ;
 assign wire2291 = ( n_n105  &  n_n94 ) | ( n_n94  &  wire41 ) | ( n_n94  &  wire175 ) ;
 assign wire2296 = ( wire166  &  n_n94 ) | ( n_n94  &  wire229 ) ;
 assign wire2299 = ( n_n57  &  n_n197 ) | ( n_n57  &  wire42 ) | ( n_n57  &  wire22476 ) ;
 assign wire2300 = ( n_n230  &  n_n271  &  n_n285  &  wire1259 ) ;
 assign wire2304 = ( n_n56  &  wire22473 ) | ( n_n56  &  wire22474 ) | ( n_n56  &  wire22475 ) ;
 assign wire2305 = ( n_n57  &  wire22473 ) | ( n_n57  &  wire22474 ) ;
 assign wire2306 = ( n_n57  &  wire276 ) | ( n_n57  &  wire182 ) | ( n_n57  &  wire22471 ) ;
 assign wire2307 = ( n_n56  &  wire53 ) | ( n_n56  &  n_n258  &  wire897 ) ;
 assign wire2308 = ( n_n57  &  n_n246 ) | ( n_n57  &  wire22467 ) | ( n_n57  &  wire22468 ) ;
 assign wire2309 = ( n_n56  &  wire22467 ) | ( n_n56  &  wire22468 ) | ( n_n56  &  wire22469 ) ;
 assign wire2311 = ( n_n48  &  wire41 ) | ( n_n48  &  wire175 ) ;
 assign wire2324 = ( wire166  &  n_n48 ) | ( n_n48  &  wire229 ) ;
 assign wire2333 = ( n_n48  &  wire112 ) | ( n_n48  &  wire144 ) ;
 assign wire2336 = ( wire124  &  wire1517 ) | ( wire1517  &  wire231 ) ;
 assign wire2344 = ( n_n6  &  n_n73 ) | ( n_n6  &  wire320 ) | ( n_n6  &  wire22435 ) ;
 assign wire2345 = ( n_n5  &  wire276 ) | ( n_n5  &  wire22436 ) | ( n_n5  &  wire22438 ) ;
 assign wire2350 = ( n_n5  &  wire233 ) | ( n_n5  &  wire22429 ) | ( n_n5  &  wire22431 ) ;
 assign wire2353 = ( n_n5  &  n_n40 ) | ( n_n5  &  wire245 ) | ( n_n5  &  wire351 ) ;
 assign wire2354 = ( n_n6  &  n_n34 ) | ( n_n6  &  n_n81 ) | ( n_n6  &  wire47 ) ;
 assign wire2355 = ( n_n5  &  wire306 ) | ( n_n5  &  wire1652 ) ;
 assign wire2356 = ( n_n6  &  n_n109 ) | ( n_n6  &  wire143 ) | ( n_n6  &  wire1652 ) ;
 assign wire2359 = ( n_n230  &  n_n261  &  n_n285  &  wire1647 ) ;
 assign wire2361 = ( n_n5  &  wire320 ) | ( n_n5  &  n_n256  &  wire914 ) ;
 assign wire2363 = ( n_n5  &  wire357 ) | ( n_n5  &  wire1124 ) ;
 assign wire2364 = ( n_n6  &  n_n52 ) | ( n_n6  &  wire1124 ) | ( n_n6  &  wire22340 ) ;
 assign wire2374 = ( n_n48  &  wire57 ) | ( n_n48  &  n_n279  &  wire914 ) ;
 assign wire2377 = ( n_n48  &  wire187 ) | ( n_n48  &  wire22407 ) ;
 assign wire2378 = ( n_n53  &  wire112 ) | ( n_n53  &  wire22408 ) ;
 assign wire2384 = ( n_n264  &  n_n283  &  n_n285  &  wire1737 ) ;
 assign wire2385 = ( wire913  &  n_n258  &  wire185 ) ;
 assign wire2392 = ( n_n53  &  n_n112 ) | ( n_n53  &  wire52 ) | ( n_n53  &  wire110 ) ;
 assign wire2393 = ( n_n48  &  wire140 ) | ( n_n48  &  wire182 ) | ( n_n48  &  wire123 ) ;
 assign wire2398 = ( n_n48  &  n_n112 ) | ( n_n48  &  wire52 ) | ( n_n48  &  wire110 ) ;
 assign wire2403 = ( n_n100  &  wire124 ) | ( n_n100  &  wire123 ) | ( n_n100  &  wire22387 ) ;
 assign wire2410 = ( i_15_  &  n_n100  &  n_n256  &  n_n270 ) | ( (~ i_15_)  &  n_n100  &  n_n256  &  n_n270 ) ;
 assign wire2425 = ( n_n56  &  wire357 ) | ( n_n56  &  n_n222  &  wire904 ) ;
 assign wire2426 = ( n_n57  &  wire76 ) | ( n_n57  &  wire229 ) | ( n_n57  &  wire22376 ) ;
 assign wire2427 = ( n_n266  &  n_n230  &  n_n285  &  wire1755 ) ;
 assign wire2428 = ( n_n56  &  wire76 ) | ( n_n56  &  wire229 ) | ( n_n56  &  wire22374 ) ;
 assign wire2430 = ( n_n94  &  wire403 ) | ( n_n94  &  wire110 ) | ( n_n94  &  wire22368 ) ;
 assign wire2436 = ( n_n100  &  wire110 ) | ( n_n100  &  n_n258  &  wire904 ) ;
 assign wire2437 = ( n_n94  &  wire123 ) | ( n_n94  &  wire187 ) ;
 assign wire2447 = ( n_n4  &  n_n81 ) | ( n_n4  &  wire233 ) | ( n_n4  &  wire22355 ) ;
 assign wire2457 = ( n_n3  &  n_n89 ) | ( n_n3  &  wire233 ) | ( n_n3  &  wire22343 ) ;
 assign wire2458 = ( n_n4  &  n_n38 ) | ( n_n4  &  wire351 ) | ( n_n4  &  wire22345 ) ;
 assign wire2463 = ( n_n3  &  n_n52 ) | ( n_n3  &  wire357 ) | ( n_n3  &  wire22340 ) ;
 assign wire2464 = ( n_n4  &  wire906  &  n_n256 ) ;
 assign wire2465 = ( n_n4  &  n_n109 ) | ( n_n4  &  wire143 ) | ( n_n4  &  wire1214 ) ;
 assign wire2472 = ( n_n3  &  n_n78 ) | ( n_n3  &  wire276 ) | ( n_n3  &  wire65 ) ;
 assign wire2473 = ( n_n4  &  n_n199 ) | ( n_n4  &  n_n73 ) | ( n_n4  &  wire22335 ) ;
 assign wire2474 = ( i_3_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire2478 = ( n_n56  &  wire40 ) | ( n_n56  &  n_n74 ) | ( n_n56  &  wire140 ) ;
 assign wire2479 = ( n_n57  &  wire22315 ) | ( n_n57  &  wire22316 ) ;
 assign wire2486 = ( n_n56  &  wire346 ) | ( n_n56  &  wire22309 ) | ( n_n56  &  wire22310 ) ;
 assign wire2491 = ( n_n57  &  wire433 ) | ( n_n57  &  wire22304 ) | ( n_n57  &  wire22305 ) ;
 assign wire2495 = ( wire51  &  n_n53 ) | ( n_n53  &  n_n90 ) | ( n_n53  &  wire448 ) ;
 assign wire2496 = ( wire166  &  n_n48 ) | ( n_n48  &  wire180 ) | ( n_n48  &  wire22298 ) ;
 assign wire2503 = ( n_n48  &  wire433 ) | ( n_n48  &  wire22290 ) | ( n_n48  &  wire22291 ) ;
 assign wire2507 = ( n_n48  &  n_n113 ) | ( n_n48  &  n_n39 ) | ( n_n48  &  wire57 ) ;
 assign wire2508 = ( n_n53  &  n_n79 ) | ( n_n53  &  n_n101 ) | ( n_n53  &  wire61 ) ;
 assign wire2516 = ( n_n53  &  n_n82 ) | ( n_n53  &  wire144 ) | ( n_n53  &  wire47 ) ;
 assign wire2520 = ( n_n57  &  n_n246 ) | ( n_n57  &  wire73 ) | ( n_n57  &  wire220 ) ;
 assign wire2521 = ( n_n56  &  wire22275 ) | ( n_n56  &  wire22276 ) ;
 assign wire2525 = ( n_n57  &  n_n107 ) | ( n_n57  &  n_n112 ) | ( n_n57  &  wire52 ) ;
 assign wire2526 = ( n_n56  &  wire60 ) | ( n_n56  &  n_n18 ) | ( n_n56  &  wire22266 ) ;
 assign wire2532 = ( n_n56  &  n_n147 ) | ( n_n56  &  n_n246 ) | ( n_n56  &  wire291 ) ;
 assign wire2533 = ( n_n57  &  n_n147 ) | ( n_n57  &  wire63 ) | ( n_n57  &  wire291 ) ;
 assign wire2534 = ( n_n56  &  wire223 ) | ( n_n56  &  wire911  &  n_n220 ) ;
 assign wire2542 = ( n_n56  &  n_n240 ) | ( n_n56  &  wire50 ) | ( n_n56  &  wire63 ) ;
 assign wire2543 = ( n_n57  &  wire223 ) | ( n_n57  &  wire22259 ) ;
 assign wire2544 = ( n_n100  &  n_n113 ) | ( n_n100  &  wire102 ) | ( n_n100  &  wire22248 ) ;
 assign wire2545 = ( n_n94  &  wire22249 ) | ( n_n94  &  wire22250 ) ;
 assign wire2550 = ( n_n100  &  n_n50 ) | ( n_n100  &  wire77 ) | ( n_n100  &  wire22244 ) ;
 assign wire2551 = ( n_n94  &  wire81 ) | ( n_n94  &  n_n46 ) | ( n_n94  &  wire22245 ) ;
 assign wire2560 = ( n_n111  &  n_n100 ) | ( n_n100  &  wire158 ) | ( n_n100  &  wire342 ) ;
 assign wire2561 = ( wire200  &  n_n94 ) | ( n_n94  &  wire78 ) | ( n_n94  &  wire85 ) ;
 assign wire2566 = ( n_n100  &  wire154 ) | ( n_n100  &  wire64 ) ;
 assign wire2571 = ( n_n56  &  n_n50 ) | ( n_n56  &  wire300 ) | ( n_n56  &  wire311 ) ;
 assign wire2572 = ( n_n57  &  wire55 ) | ( n_n57  &  n_n228  &  wire914 ) ;
 assign wire2581 = ( n_n94  &  wire63 ) | ( n_n94  &  wire913  &  n_n258 ) ;
 assign wire2583 = ( n_n100  &  n_n58 ) | ( n_n100  &  wire75 ) | ( n_n100  &  wire223 ) ;
 assign wire2593 = ( n_n100  &  wire73 ) | ( n_n100  &  wire220 ) | ( n_n100  &  wire22206 ) ;
 assign wire2594 = ( n_n94  &  wire22210 ) | ( n_n94  &  wire22211 ) ;
 assign wire2596 = ( n_n100  &  wire63 ) | ( n_n100  &  wire903  &  n_n258 ) ;
 assign wire2597 = ( n_n260  &  n_n263  &  n_n285  &  wire50 ) ;
 assign wire2601 = ( n_n260  &  n_n263  &  n_n285  &  wire1113 ) ;
 assign wire2602 = ( n_n100  &  wire22195 ) | ( n_n100  &  wire22196 ) | ( n_n100  &  wire22197 ) ;
 assign wire2623 = ( n_n94  &  wire110 ) | ( n_n94  &  wire232 ) | ( n_n94  &  wire274 ) ;
 assign wire2631 = ( n_n48  &  wire345 ) | ( n_n48  &  wire22170 ) | ( n_n48  &  wire22171 ) ;
 assign wire2637 = ( n_n53  &  wire95 ) | ( n_n53  &  wire220 ) | ( n_n53  &  wire22162 ) ;
 assign wire2638 = ( n_n48  &  wire22167 ) | ( n_n48  &  wire22168 ) ;
 assign wire2640 = ( n_n53  &  wire62 ) | ( n_n53  &  wire911  &  n_n281 ) ;
 assign wire2652 = ( n_n6  &  wire166 ) | ( n_n6  &  n_n50 ) | ( n_n6  &  wire180 ) ;
 assign wire2659 = ( n_n53  &  wire22139 ) | ( n_n53  &  n_n222  &  wire907 ) ;
 assign wire2665 = ( n_n264  &  n_n283  &  n_n285  &  wire50 ) ;
 assign wire2672 = ( n_n48  &  wire75 ) | ( n_n48  &  n_n258  &  wire908 ) ;
 assign wire2673 = ( n_n53  &  wire50 ) | ( n_n53  &  wire913  &  n_n258 ) ;
 assign wire2676 = ( n_n6  &  n_n102 ) | ( n_n6  &  wire807 ) | ( n_n6  &  wire311 ) ;
 assign wire2686 = ( n_n53  &  wire64 ) | ( n_n53  &  n_n279  &  wire907 ) ;
 assign wire2692 = ( n_n6  &  wire345 ) | ( n_n6  &  wire22115 ) ;
 assign wire2698 = ( n_n6  &  n_n113 ) | ( n_n6  &  wire102 ) | ( n_n6  &  wire22108 ) ;
 assign wire2699 = ( n_n5  &  wire22109 ) | ( n_n5  &  wire22110 ) ;
 assign wire2703 = ( n_n5  &  n_n87 ) | ( n_n5  &  wire55 ) | ( n_n5  &  wire342 ) ;
 assign wire2704 = ( n_n6  &  wire165 ) | ( n_n6  &  wire140 ) | ( n_n6  &  wire22104 ) ;
 assign wire2708 = ( n_n5  &  n_n147 ) | ( n_n5  &  n_n246 ) | ( n_n5  &  wire291 ) ;
 assign wire2709 = ( n_n6  &  n_n147 ) | ( n_n6  &  wire63 ) | ( n_n6  &  wire291 ) ;
 assign wire2725 = ( n_n240  &  n_n207 ) | ( n_n207  &  n_n17 ) | ( n_n207  &  wire514 ) ;
 assign wire2726 = ( n_n227  &  wire49 ) | ( n_n227  &  n_n228  &  wire908 ) ;
 assign wire2740 = ( n_n4  &  n_n20 ) | ( n_n4  &  wire42 ) | ( n_n4  &  wire66 ) ;
 assign wire2745 = ( n_n1  &  wire22058 ) | ( n_n1  &  wire22059 ) ;
 assign wire2774 = ( n_n240  &  n_n5 ) | ( n_n5  &  wire50 ) | ( n_n5  &  wire63 ) ;
 assign wire2775 = ( n_n6  &  wire223 ) | ( n_n6  &  wire22033 ) ;
 assign wire2776 = ( n_n5  &  wire220 ) | ( n_n5  &  wire22024 ) | ( n_n5  &  wire22026 ) ;
 assign wire2777 = ( n_n6  &  wire247 ) | ( n_n6  &  wire220 ) | ( n_n6  &  wire22029 ) ;
 assign wire2780 = ( n_n5  &  wire223 ) | ( n_n5  &  wire911  &  n_n220 ) ;
 assign wire2781 = ( n_n207  &  wire425 ) | ( n_n207  &  n_n228  &  wire903 ) ;
 assign wire2784 = ( n_n6  &  wire274 ) | ( n_n6  &  wire899  &  n_n281 ) ;
 assign wire2785 = ( n_n5  &  wire22016 ) | ( n_n5  &  wire22017 ) ;
 assign wire2790 = ( n_n3  &  wire448 ) | ( n_n3  &  wire22009 ) ;
 assign wire2798 = ( n_n268  &  wire95 ) | ( n_n268  &  wire22001 ) | ( n_n268  &  wire22004 ) ;
 assign wire2804 = ( n_n4  &  wire99 ) | ( n_n4  &  wire41 ) ;
 assign wire2808 = ( n_n268  &  wire21997 ) | ( n_n268  &  wire21998 ) ;
 assign wire2811 = ( n_n229  &  n_n285  &  n_n284  &  wire41 ) ;
 assign wire2813 = ( n_n2  &  wire95 ) | ( n_n2  &  wire898  &  n_n220 ) ;
 assign wire2814 = ( n_n1  &  wire95 ) | ( n_n1  &  wire901  &  n_n220 ) ;
 assign wire2822 = ( n_n2  &  wire21983 ) | ( n_n2  &  wire21984 ) | ( n_n2  &  wire21985 ) ;
 assign wire2825 = ( n_n1  &  wire21979 ) | ( n_n1  &  wire21980 ) ;
 assign wire2827 = ( wire75  &  wire1423 ) | ( wire899  &  n_n220  &  wire1423 ) ;
 assign wire2830 = ( n_n2  &  wire63 ) | ( n_n2  &  wire21971 ) ;
 assign wire2831 = ( n_n1  &  n_n257 ) | ( n_n1  &  wire50 ) | ( n_n1  &  wire63 ) ;
 assign wire2839 = ( n_n2  &  wire21958 ) | ( n_n2  &  wire21959 ) | ( n_n2  &  wire21960 ) ;
 assign wire2842 = ( n_n1  &  wire21953 ) | ( n_n1  &  wire21954 ) ;
 assign wire2845 = ( n_n4  &  wire40 ) | ( n_n4  &  n_n74 ) | ( n_n4  &  wire346 ) ;
 assign wire2846 = ( n_n3  &  wire21943 ) | ( n_n3  &  wire21944 ) ;
 assign wire2854 = ( n_n3  &  wire21938 ) | ( n_n3  &  wire21939 ) ;
 assign wire2858 = ( n_n3  &  wire347 ) | ( n_n3  &  wire21929 ) ;
 assign wire2864 = ( n_n4  &  wire95 ) | ( n_n4  &  wire898  &  n_n220 ) ;
 assign wire2874 = ( n_n4  &  wire75 ) | ( n_n4  &  wire50 ) ;
 assign wire2879 = ( n_n3  &  wire95 ) | ( n_n3  &  wire21913 ) ;
 assign wire2883 = ( n_n4  &  n_n68 ) | ( n_n4  &  wire514 ) | ( n_n4  &  wire325 ) ;
 assign wire2885 = ( n_n3  &  wire123 ) | ( n_n3  &  wire100 ) ;
 assign wire2888 = ( wire992  &  n_n208  &  n_n285  &  n_n284 ) ;
 assign wire2889 = ( n_n3  &  wire343 ) | ( n_n3  &  wire431 ) | ( n_n3  &  wire21907 ) ;
 assign wire2893 = ( n_n3  &  n_n88 ) | ( n_n3  &  wire154 ) ;
 assign wire2901 = ( n_n4  &  wire195 ) | ( n_n4  &  wire21892 ) ;
 assign wire2902 = ( n_n3  &  n_n8 ) | ( n_n3  &  wire375 ) | ( n_n3  &  wire21895 ) ;
 assign wire2906 = ( n_n229  &  n_n285  &  n_n284  &  wire1668 ) ;
 assign wire2907 = ( wire169  &  wire901  &  n_n220 ) ;
 assign wire2912 = ( n_n4  &  n_n71 ) | ( n_n4  &  wire143 ) | ( n_n4  &  wire1822 ) ;
 assign wire2913 = ( n_n3  &  wire195 ) | ( n_n3  &  wire230 ) | ( n_n3  &  wire1822 ) ;
 assign wire2917 = ( n_n3  &  n_n80 ) | ( n_n3  &  n_n29 ) | ( n_n3  &  wire61 ) ;
 assign wire2918 = ( n_n4  &  n_n24 ) | ( n_n4  &  wire104 ) | ( n_n4  &  wire228 ) ;
 assign wire2919 = ( n_n94  &  n_n34 ) | ( n_n94  &  wire154 ) | ( n_n94  &  wire263 ) ;
 assign wire2920 = ( n_n260  &  n_n261  &  n_n285  &  wire1835 ) ;
 assign wire2927 = ( n_n100  &  wire21866 ) | ( n_n100  &  wire21867 ) ;
 assign wire2928 = ( n_n94  &  wire363 ) | ( n_n94  &  wire21868 ) | ( n_n94  &  wire21869 ) ;
 assign wire2929 = ( n_n100  &  n_n97 ) | ( n_n100  &  wire226 ) | ( n_n100  &  wire361 ) ;
 assign wire2939 = ( n_n100  &  wire230 ) | ( n_n100  &  wire902  &  n_n256 ) ;
 assign wire2942 = ( n_n53  &  wire61 ) | ( n_n53  &  n_n222  &  wire908 ) ;
 assign wire2943 = ( n_n264  &  n_n283  &  n_n285  &  wire102 ) ;
 assign wire2952 = ( n_n48  &  n_n203 ) | ( n_n48  &  wire230 ) ;
 assign wire2960 = ( n_n48  &  n_n80 ) | ( n_n48  &  n_n29 ) | ( n_n48  &  wire61 ) ;
 assign wire2961 = ( n_n53  &  n_n24 ) | ( n_n53  &  wire104 ) | ( n_n53  &  wire228 ) ;
 assign wire2967 = ( n_n48  &  wire21837 ) | ( n_n48  &  wire21838 ) ;
 assign wire2972 = ( n_n56  &  wire899  &  n_n220 ) ;
 assign wire2973 = ( n_n48  &  n_n37 ) | ( n_n48  &  n_n83 ) | ( n_n48  &  wire64 ) ;
 assign wire2974 = ( n_n53  &  n_n86 ) | ( n_n53  &  wire102 ) | ( n_n53  &  wire263 ) ;
 assign wire2975 = ( n_n53  &  wire64 ) | ( n_n53  &  n_n222  &  wire907 ) ;
 assign wire2976 = ( n_n264  &  n_n283  &  n_n285  &  wire154 ) ;
 assign wire2981 = ( n_n5  &  n_n88 ) | ( n_n5  &  wire154 ) | ( n_n5  &  wire21820 ) ;
 assign wire2982 = ( n_n6  &  wire154 ) | ( n_n6  &  wire21821 ) | ( n_n6  &  wire21823 ) ;
 assign wire2994 = ( n_n6  &  wire195 ) | ( n_n6  &  wire898  &  n_n220 ) ;
 assign wire2999 = ( n_n5  &  n_n203 ) | ( n_n5  &  wire195 ) | ( n_n5  &  wire21804 ) ;
 assign wire3000 = ( n_n6  &  n_n203 ) | ( n_n6  &  wire21805 ) | ( n_n6  &  wire21807 ) ;
 assign wire3003 = ( n_n5  &  n_n80 ) | ( n_n5  &  n_n29 ) | ( n_n5  &  wire61 ) ;
 assign wire3004 = ( n_n6  &  n_n24 ) | ( n_n6  &  wire104 ) | ( n_n6  &  wire228 ) ;
 assign wire3005 = ( n_n6  &  wire230 ) | ( n_n6  &  n_n222  &  wire897 ) ;
 assign wire3008 = ( n_n5  &  wire21797 ) | ( n_n5  &  wire21798 ) ;
 assign wire3012 = ( n_n6  &  n_n52 ) | ( n_n6  &  wire807 ) | ( n_n6  &  wire21789 ) ;
 assign wire3018 = ( n_n53  &  wire21785 ) | ( n_n53  &  n_n222  &  wire907 ) ;
 assign wire3019 = ( wire911  &  n_n220  &  wire185 ) ;
 assign wire3032 = ( n_n53  &  n_n69 ) | ( n_n53  &  wire84 ) | ( n_n53  &  wire21775 ) ;
 assign wire3033 = ( n_n48  &  wire21777 ) | ( n_n48  &  wire21778 ) ;
 assign wire3043 = ( n_n5  &  n_n37 ) | ( n_n5  &  n_n83 ) | ( n_n5  &  wire64 ) ;
 assign wire3045 = ( n_n230  &  n_n271  &  n_n285  &  wire1600 ) ;
 assign wire3056 = ( n_n94  &  n_n78 ) | ( n_n94  &  n_n69 ) | ( n_n94  &  wire230 ) ;
 assign wire3065 = ( n_n260  &  n_n263  &  n_n285  &  wire236 ) ;
 assign wire3072 = ( wire899  &  n_n220  &  wire1196 ) ;
 assign wire3080 = ( n_n230  &  n_n271  &  n_n285  &  wire1251 ) ;
 assign wire3098 = ( n_n230  &  n_n271  &  n_n285  &  wire1250 ) ;
 assign wire3106 = ( n_n56  &  wire100 ) | ( n_n56  &  wire1199 ) ;
 assign wire3109 = ( n_n57  &  wire472 ) | ( n_n57  &  wire100 ) ;
 assign wire3120 = ( n_n1  &  n_n97 ) | ( n_n1  &  wire226 ) | ( n_n1  &  wire361 ) ;
 assign wire3121 = ( n_n2  &  wire21705 ) | ( n_n2  &  wire21706 ) ;
 assign wire3145 = ( n_n4  &  wire61 ) | ( n_n4  &  n_n222  &  wire908 ) ;
 assign wire3159 = ( n_n208  &  n_n285  &  n_n284  &  wire1793 ) ;
 assign wire3178 = ( n_n3  &  n_n44 ) | ( n_n3  &  wire270 ) | ( n_n3  &  wire21668 ) ;
 assign wire3179 = ( n_n4  &  n_n88 ) | ( n_n4  &  n_n44 ) | ( n_n4  &  wire21668 ) ;
 assign wire3186 = ( n_n3  &  n_n99 ) | ( n_n3  &  n_n52 ) | ( n_n3  &  wire807 ) ;
 assign wire3187 = ( n_n208  &  n_n285  &  n_n284  &  wire270 ) ;
 assign wire3190 = ( n_n265  &  wire200 ) | ( n_n265  &  wire158 ) ;
 assign wire3198 = ( n_n268  &  n_n58 ) | ( n_n268  &  wire429 ) | ( n_n268  &  wire21658 ) ;
 assign wire3203 = ( n_n260  &  n_n273  &  n_n285  &  wire1773 ) ;
 assign wire3211 = ( n_n2  &  n_n20 ) | ( n_n2  &  wire375 ) | ( n_n2  &  wire21650 ) ;
 assign wire3213 = ( n_n3  &  n_n37 ) | ( n_n3  &  n_n83 ) | ( n_n3  &  wire64 ) ;
 assign wire3214 = ( n_n4  &  n_n86 ) | ( n_n4  &  wire102 ) | ( n_n4  &  wire263 ) ;
 assign wire3215 = ( n_n2  &  wire424 ) | ( n_n2  &  wire428 ) | ( n_n2  &  wire21643 ) ;
 assign wire3219 = ( n_n1  &  n_n20 ) | ( n_n1  &  wire375 ) | ( n_n1  &  wire1792 ) ;
 assign wire3220 = ( n_n2  &  wire1792 ) | ( n_n2  &  wire21642 ) ;
 assign wire3221 = ( n_n2  &  wire21636 ) | ( n_n2  &  wire21637 ) ;
 assign wire3222 = ( n_n1  &  wire21639 ) | ( n_n1  &  wire21640 ) ;
 assign wire3228 = ( n_n3  &  n_n86 ) | ( n_n3  &  wire102 ) | ( n_n3  &  wire263 ) ;
 assign wire3232 = ( n_n127  &  wire48 ) | ( n_n127  &  wire913  &  n_n220 ) ;
 assign wire3241 = ( n_n273  &  n_n165  &  n_n284  &  wire1825 ) ;
 assign wire3255 = ( n_n48  &  wire1529 ) | ( n_n48  &  wire21608 ) ;
 assign wire3256 = ( n_n264  &  n_n273  &  n_n285  &  wire1528 ) ;
 assign wire3261 = ( n_n48  &  wire1508 ) | ( n_n48  &  n_n279  &  wire899 ) ;
 assign wire3262 = ( n_n53  &  wire1508 ) | ( n_n53  &  n_n279  &  wire905 ) ;
 assign wire3270 = ( n_n48  &  wire21599 ) | ( n_n48  &  wire21600 ) ;
 assign wire3272 = ( i_15_  &  n_n48  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n48  &  n_n279  &  n_n247 ) ;
 assign wire3277 = ( i_15_  &  n_n53  &  n_n279  &  n_n270 ) | ( (~ i_15_)  &  n_n53  &  n_n279  &  n_n270 ) ;
 assign wire3282 = ( n_n186  &  n_n5 ) | ( n_n5  &  wire51 ) | ( n_n5  &  wire21583 ) ;
 assign wire3283 = ( n_n6  &  wire51 ) | ( n_n6  &  wire21584 ) | ( n_n6  &  wire21586 ) ;
 assign wire3287 = ( n_n6  &  n_n84 ) | ( n_n6  &  n_n35 ) | ( n_n6  &  wire86 ) ;
 assign wire3288 = ( n_n5  &  wire78 ) | ( n_n5  &  wire21576 ) | ( n_n5  &  wire21578 ) ;
 assign wire3292 = ( n_n6  &  n_n30 ) | ( n_n6  &  n_n101 ) | ( n_n6  &  wire80 ) ;
 assign wire3296 = ( n_n264  &  n_n273  &  n_n285  &  wire1485 ) ;
 assign wire3297 = ( n_n281  &  wire913  &  wire185 ) ;
 assign wire3303 = ( n_n264  &  n_n283  &  n_n285  &  wire1327 ) ;
 assign wire3310 = ( n_n281  &  wire907  &  wire185 ) ;
 assign wire3316 = ( n_n5  &  n_n93 ) | ( n_n5  &  n_n90 ) | ( n_n5  &  wire21389 ) ;
 assign wire3317 = ( n_n6  &  wire71 ) | ( n_n6  &  n_n279  &  wire904 ) ;
 assign wire3320 = ( n_n5  &  wire21554 ) | ( n_n5  &  wire21555 ) ;
 assign wire3324 = ( n_n260  &  n_n263  &  n_n285  &  wire1158 ) ;
 assign wire3340 = ( n_n207  &  wire21536 ) | ( n_n207  &  wire903  &  n_n225 ) ;
 assign wire3344 = ( wire48  &  n_n5 ) | ( n_n5  &  n_n204 ) | ( n_n5  &  n_n16 ) ;
 assign wire3345 = ( n_n6  &  wire79 ) | ( n_n6  &  n_n279  &  wire905 ) ;
 assign wire3354 = ( n_n5  &  n_n109 ) | ( n_n5  &  wire79 ) | ( n_n5  &  wire83 ) ;
 assign wire3358 = ( n_n5  &  wire62 ) | ( n_n5  &  n_n279  &  wire899 ) ;
 assign wire3360 = ( n_n229  &  n_n285  &  n_n284  &  wire1450 ) ;
 assign wire3361 = ( wire169  &  n_n281  &  wire907 ) ;
 assign wire3368 = ( n_n3  &  wire62 ) | ( n_n3  &  n_n279  &  wire899 ) ;
 assign wire3370 = ( n_n3  &  wire79 ) | ( n_n3  &  n_n279  &  wire905 ) ;
 assign wire3375 = ( n_n100  &  wire157 ) | ( n_n100  &  wire167 ) | ( n_n100  &  wire235 ) ;
 assign wire3376 = ( wire268  &  n_n94 ) | ( n_n94  &  wire157 ) | ( n_n94  &  wire436 ) ;
 assign wire3382 = ( n_n266  &  n_n230  &  n_n285  &  wire1530 ) ;
 assign wire3393 = ( wire1378  &  wire1377 ) ;
 assign wire3398 = ( n_n48  &  wire51 ) | ( n_n48  &  n_n279  &  wire898 ) ;
 assign wire3400 = ( n_n48  &  n_n93 ) | ( n_n48  &  n_n90 ) | ( n_n48  &  wire21389 ) ;
 assign wire3401 = ( n_n53  &  n_n102 ) | ( n_n53  &  wire77 ) | ( n_n53  &  wire71 ) ;
 assign wire3402 = ( n_n230  &  n_n271  &  n_n285  &  wire1095 ) ;
 assign wire3409 = ( i_15_  &  n_n242  &  n_n279  &  wire1094 ) | ( (~ i_15_)  &  n_n242  &  n_n279  &  wire1094 ) ;
 assign wire3413 = ( n_n56  &  n_n70 ) | ( n_n56  &  wire79 ) | ( n_n56  &  wire413 ) ;
 assign wire3416 = ( n_n56  &  wire264 ) | ( n_n56  &  n_n73 ) | ( n_n56  &  wire19408 ) ;
 assign wire3419 = ( n_n260  &  n_n263  &  n_n285  &  wire330 ) ;
 assign wire3428 = ( n_n94  &  wire119 ) | ( n_n94  &  wire167 ) | ( n_n94  &  wire21477 ) ;
 assign wire3432 = ( n_n56  &  n_n81 ) | ( n_n56  &  wire86 ) | ( n_n56  &  wire21464 ) ;
 assign wire3440 = ( n_n100  &  n_n148 ) | ( n_n100  &  wire210 ) | ( n_n100  &  wire399 ) ;
 assign wire3441 = ( n_n94  &  wire21457 ) | ( n_n94  &  wire21458 ) ;
 assign wire3442 = ( n_n281  &  wire903  &  wire168 ) ;
 assign wire3447 = ( n_n94  &  wire281 ) | ( n_n94  &  wire338 ) ;
 assign wire3451 = ( i_15_  &  n_n56  &  n_n253  &  n_n279 ) | ( (~ i_15_)  &  n_n56  &  n_n253  &  n_n279 ) ;
 assign wire3452 = ( n_n57  &  wire19384 ) | ( n_n57  &  n_n281  &  wire900 ) ;
 assign wire3469 = ( n_n1  &  wire255 ) | ( n_n1  &  wire242 ) ;
 assign wire3470 = ( n_n264  &  n_n273  &  n_n285  &  wire1163 ) ;
 assign wire3480 = ( n_n3  &  wire71 ) | ( n_n3  &  n_n279  &  wire904 ) ;
 assign wire3489 = ( n_n260  &  n_n273  &  n_n285  &  wire1159 ) ;
 assign wire3490 = ( n_n2  &  wire241 ) | ( n_n2  &  wire242 ) | ( n_n2  &  wire21424 ) ;
 assign wire3491 = ( n_n2  &  n_n84 ) | ( n_n2  &  n_n35 ) | ( n_n2  &  wire86 ) ;
 assign wire3496 = ( n_n2  &  wire157 ) | ( n_n2  &  wire330 ) | ( n_n2  &  wire21414 ) ;
 assign wire3499 = ( n_n2  &  wire281 ) | ( n_n2  &  wire338 ) | ( n_n2  &  wire1101 ) ;
 assign wire3500 = ( n_n1  &  n_n60 ) | ( n_n1  &  wire210 ) | ( n_n1  &  wire1101 ) ;
 assign wire3507 = ( n_n260  &  n_n283  &  n_n285  &  wire1097 ) ;
 assign wire3508 = ( n_n1  &  wire338 ) | ( n_n1  &  wire399 ) | ( n_n1  &  wire21402 ) ;
 assign wire3510 = ( n_n4  &  n_n179 ) | ( n_n4  &  wire77 ) | ( n_n4  &  wire21393 ) ;
 assign wire3518 = ( n_n4  &  wire51 ) | ( n_n4  &  n_n90 ) | ( n_n4  &  wire21389 ) ;
 assign wire3520 = ( n_n265  &  wire252 ) | ( n_n265  &  n_n81 ) | ( n_n265  &  wire86 ) ;
 assign wire3521 = ( n_n268  &  wire21383 ) | ( n_n268  &  wire21384 ) ;
 assign wire3528 = ( n_n265  &  n_n281  &  wire907 ) ;
 assign wire3530 = ( n_n4  &  wire67 ) | ( n_n4  &  wire1037 ) ;
 assign wire3531 = ( n_n3  &  wire1037 ) | ( n_n3  &  wire21377 ) ;
 assign wire3533 = ( n_n3  &  wire67 ) | ( n_n3  &  n_n279  &  wire897 ) ;
 assign wire3534 = ( n_n4  &  wire80 ) | ( n_n4  &  n_n279  &  wire908 ) ;
 assign wire3538 = ( n_n3  &  wire21370 ) | ( n_n3  &  wire21371 ) ;
 assign wire3541 = ( wire48  &  n_n3 ) | ( n_n3  &  n_n204 ) | ( n_n3  &  n_n16 ) ;
 assign wire3542 = ( n_n4  &  wire79 ) | ( n_n4  &  n_n279  &  wire905 ) ;
 assign wire3544 = ( n_n57  &  n_n7 ) | ( n_n57  &  n_n257 ) | ( n_n57  &  wire72 ) ;
 assign wire3550 = ( n_n57  &  wire44 ) | ( n_n57  &  n_n252 ) | ( n_n57  &  n_n15 ) ;
 assign wire3551 = ( n_n56  &  wire117 ) | ( n_n56  &  wire21353 ) | ( n_n56  &  wire21354 ) ;
 assign wire3558 = ( n_n57  &  wire203 ) | ( n_n57  &  wire21347 ) | ( n_n57  &  wire21348 ) ;
 assign wire3562 = ( n_n56  &  wire21339 ) | ( n_n56  &  wire21340 ) ;
 assign wire3563 = ( n_n57  &  wire21341 ) | ( n_n57  &  wire21342 ) | ( n_n57  &  wire21343 ) ;
 assign wire3565 = ( n_n57  &  wire117 ) | ( n_n57  &  wire21334 ) | ( n_n57  &  wire21335 ) ;
 assign wire3572 = ( n_n56  &  n_n148 ) | ( n_n56  &  wire113 ) | ( n_n56  &  wire21328 ) ;
 assign wire3576 = ( n_n56  &  n_n7 ) | ( n_n56  &  wire50 ) | ( n_n56  &  n_n59 ) ;
 assign wire3577 = ( n_n57  &  wire50 ) | ( n_n57  &  n_n59 ) | ( n_n57  &  wire208 ) ;
 assign wire3578 = ( n_n56  &  wire62 ) | ( n_n56  &  wire21322 ) | ( n_n56  &  wire21323 ) ;
 assign wire3579 = ( n_n57  &  wire21322 ) | ( n_n57  &  wire21323 ) ;
 assign wire3584 = ( n_n57  &  wire246 ) | ( n_n57  &  wire256 ) ;
 assign wire3585 = ( n_n56  &  n_n281  &  wire906 ) ;
 assign wire3588 = ( n_n56  &  wire202 ) | ( n_n56  &  wire21315 ) | ( n_n56  &  wire21316 ) ;
 assign wire3594 = ( n_n56  &  wire21306 ) | ( n_n56  &  wire21307 ) ;
 assign wire3595 = ( n_n57  &  wire21309 ) | ( n_n57  &  wire21310 ) ;
 assign wire3600 = ( n_n56  &  n_n46 ) | ( n_n56  &  wire19577 ) | ( n_n56  &  wire21297 ) ;
 assign wire3612 = ( n_n4  &  n_n99 ) | ( n_n4  &  wire96 ) | ( n_n4  &  wire21284 ) ;
 assign wire3613 = ( n_n3  &  wire21285 ) | ( n_n3  &  wire21286 ) ;
 assign wire3619 = ( n_n268  &  wire21277 ) | ( n_n268  &  wire21278 ) ;
 assign wire3620 = ( n_n265  &  wire21279 ) | ( n_n265  &  wire21280 ) ;
 assign wire3626 = ( n_n268  &  wire21272 ) | ( n_n268  &  wire21273 ) | ( n_n268  &  wire21274 ) ;
 assign wire3627 = ( n_n266  &  n_n285  &  n_n284  &  wire101 ) ;
 assign wire3629 = ( n_n268  &  wire160 ) | ( n_n268  &  n_n59 ) | ( n_n268  &  wire21266 ) ;
 assign wire3636 = ( n_n268  &  n_n73 ) | ( n_n268  &  wire19408 ) | ( n_n268  &  wire21247 ) ;
 assign wire3642 = ( n_n3  &  n_n11 ) | ( n_n3  &  n_n148 ) | ( n_n3  &  wire95 ) ;
 assign wire3653 = ( n_n3  &  n_n99 ) | ( n_n3  &  n_n54 ) | ( n_n3  &  wire96 ) ;
 assign wire3660 = ( n_n3  &  wire78 ) | ( n_n3  &  wire21230 ) | ( n_n3  &  wire21231 ) ;
 assign wire3661 = ( n_n4  &  wire21230 ) | ( n_n4  &  wire21231 ) | ( n_n4  &  wire21232 ) ;
 assign wire3662 = ( n_n4  &  n_n258  &  wire912 ) ;
 assign wire3664 = ( n_n3  &  wire21223 ) | ( n_n3  &  wire21224 ) ;
 assign wire3665 = ( n_n4  &  wire80 ) | ( n_n4  &  wire902  &  n_n256 ) ;
 assign wire3673 = ( n_n4  &  wire40 ) | ( n_n4  &  wire203 ) | ( n_n4  &  wire21217 ) ;
 assign wire3674 = ( n_n3  &  wire203 ) | ( n_n3  &  wire21217 ) | ( n_n3  &  wire21218 ) ;
 assign wire3680 = ( n_n4  &  wire21211 ) | ( n_n4  &  wire21212 ) ;
 assign wire3681 = ( n_n3  &  wire21213 ) | ( n_n3  &  wire21214 ) | ( n_n3  &  wire21215 ) ;
 assign wire3682 = ( n_n3  &  wire97 ) | ( n_n3  &  wire21203 ) | ( n_n3  &  wire21204 ) ;
 assign wire3688 = ( n_n3  &  n_n12 ) | ( n_n3  &  n_n65 ) | ( n_n3  &  wire73 ) ;
 assign wire3689 = ( n_n4  &  wire44 ) | ( n_n4  &  n_n252 ) | ( n_n4  &  n_n15 ) ;
 assign wire3698 = ( n_n3  &  wire113 ) | ( n_n3  &  wire101 ) ;
 assign wire3702 = ( n_n3  &  wire208 ) | ( n_n3  &  wire199 ) ;
 assign wire3707 = ( n_n3  &  n_n7 ) | ( n_n3  &  wire50 ) | ( n_n3  &  n_n59 ) ;
 assign wire3708 = ( n_n4  &  wire50 ) | ( n_n4  &  n_n228  &  wire897 ) ;
 assign wire3712 = ( n_n152  &  n_n220  &  wire914 ) ;
 assign wire3720 = ( n_n139  &  n_n135 ) | ( n_n139  &  wire419 ) | ( n_n139  &  wire19604 ) ;
 assign wire3725 = ( n_n110  &  n_n128 ) | ( n_n128  &  n_n111 ) | ( n_n128  &  wire54 ) ;
 assign wire3726 = ( wire48  &  n_n130 ) | ( n_n130  &  n_n110 ) | ( n_n130  &  wire54 ) ;
 assign wire3733 = ( wire48  &  n_n121 ) | ( n_n110  &  n_n121 ) | ( n_n121  &  wire54 ) ;
 assign wire3736 = ( n_n3  &  n_n9 ) | ( n_n3  &  wire184 ) | ( n_n3  &  wire63 ) ;
 assign wire3745 = ( n_n3  &  wire21141 ) | ( n_n3  &  wire21142 ) ;
 assign wire3754 = ( n_n3  &  wire93 ) | ( n_n3  &  wire136 ) | ( n_n3  &  wire21138 ) ;
 assign wire3755 = ( n_n4  &  n_n111 ) | ( n_n4  &  wire136 ) | ( n_n4  &  wire21138 ) ;
 assign wire3758 = ( n_n3  &  wire21134 ) | ( n_n3  &  wire21135 ) ;
 assign wire3762 = ( n_n3  &  n_n220  &  wire908 ) ;
 assign wire3764 = ( n_n260  &  n_n271  &  n_n285  &  wire1322 ) ;
 assign wire3771 = ( n_n94  &  n_n78 ) | ( n_n94  &  wire80 ) | ( n_n94  &  wire21103 ) ;
 assign wire3778 = ( n_n94  &  n_n97 ) | ( n_n94  &  wire71 ) | ( n_n94  &  wire453 ) ;
 assign wire3790 = ( n_n94  &  n_n14 ) | ( n_n94  &  wire70 ) | ( n_n94  &  wire199 ) ;
 assign wire3791 = ( n_n260  &  n_n261  &  wire184  &  n_n285 ) ;
 assign wire3800 = ( n_n100  &  wire72 ) | ( n_n100  &  n_n258  &  wire905 ) ;
 assign wire3821 = ( n_n264  &  n_n263  &  n_n285  &  wire1323 ) ;
 assign wire3830 = ( n_n48  &  wire68 ) | ( n_n48  &  n_n49 ) | ( n_n48  &  wire71 ) ;
 assign wire3831 = ( n_n53  &  n_n95 ) | ( n_n53  &  n_n179 ) | ( n_n53  &  wire57 ) ;
 assign wire3837 = ( n_n5  &  wire87 ) | ( n_n5  &  wire914  &  n_n225 ) ;
 assign wire3843 = ( n_n48  &  wire63 ) | ( n_n48  &  n_n228  &  wire902 ) ;
 assign wire3852 = ( n_n48  &  n_n179 ) | ( n_n48  &  wire57 ) | ( n_n48  &  wire21009 ) ;
 assign wire3860 = ( n_n264  &  wire44  &  n_n273  &  n_n285 ) ;
 assign wire3870 = ( n_n227  &  wire88 ) | ( n_n227  &  wire306 ) | ( n_n227  &  wire20980 ) ;
 assign wire3884 = ( n_n2  &  n_n29 ) | ( n_n2  &  wire49 ) | ( n_n2  &  wire88 ) ;
 assign wire3889 = ( n_n2  &  n_n179 ) | ( n_n2  &  wire57 ) | ( n_n2  &  wire20958 ) ;
 assign wire3896 = ( n_n5  &  n_n144 ) | ( n_n5  &  wire118 ) | ( n_n5  &  wire199 ) ;
 assign wire3904 = ( n_n6  &  wire160 ) | ( n_n6  &  wire184 ) ;
 assign wire3924 = ( n_n268  &  n_n11 ) | ( n_n268  &  wire157 ) | ( n_n268  &  wire95 ) ;
 assign wire3931 = ( n_n1  &  wire72 ) | ( n_n1  &  n_n228  &  wire902 ) ;
 assign wire3932 = ( n_n2  &  n_n9 ) | ( n_n2  &  wire63 ) | ( n_n2  &  wire20928 ) ;
 assign wire3943 = ( wire396  &  n_n281  &  wire907 ) ;
 assign wire3945 = ( (~ i_9_)  &  (~ i_10_)  &  n_n122 ) | ( (~ i_9_)  &  (~ i_10_)  &  wire20917 ) ;
 assign wire3946 = ( wire923  &  n_n283  &  n_n165  &  wire19294 ) ;
 assign wire3967 = ( n_n5  &  wire100 ) | ( n_n5  &  wire281 ) ;
 assign wire3968 = ( n_n6  &  n_n14 ) | ( n_n6  &  wire70 ) | ( n_n6  &  wire118 ) ;
 assign wire3975 = ( n_n4  &  wire166 ) | ( n_n4  &  wire905  &  n_n225 ) ;
 assign wire3976 = ( n_n94  &  wire130 ) | ( n_n94  &  wire911  &  n_n228 ) ;
 assign wire3985 = ( n_n4  &  wire123 ) | ( n_n4  &  wire100 ) ;
 assign wire3988 = ( n_n207  &  n_n112 ) | ( n_n207  &  wire52 ) | ( n_n207  &  wire20874 ) ;
 assign wire3989 = ( n_n227  &  wire123 ) | ( n_n227  &  wire20875 ) ;
 assign wire4004 = ( n_n1  &  n_n257 ) | ( n_n1  &  n_n226 ) | ( n_n1  &  wire72 ) ;
 assign wire4005 = ( n_n2  &  wire66 ) | ( n_n2  &  wire899  &  n_n256 ) ;
 assign wire4016 = ( n_n48  &  wire44 ) | ( n_n48  &  wire75 ) | ( n_n48  &  n_n206 ) ;
 assign wire4027 = ( wire60  &  n_n53 ) | ( n_n53  &  wire1656 ) ;
 assign wire4028 = ( n_n48  &  wire1656 ) | ( n_n48  &  wire20846 ) ;
 assign wire4035 = ( n_n6  &  wire20839 ) | ( n_n6  &  wire20840 ) ;
 assign wire4036 = ( n_n5  &  wire60 ) | ( n_n5  &  n_n279  &  wire911 ) ;
 assign wire4042 = ( n_n6  &  wire60 ) | ( n_n6  &  n_n204 ) | ( n_n6  &  wire1619 ) ;
 assign wire4043 = ( n_n5  &  wire123 ) | ( n_n5  &  wire227 ) | ( n_n5  &  wire1619 ) ;
 assign wire4044 = ( n_n57  &  wire72 ) | ( n_n57  &  n_n258  &  wire905 ) ;
 assign wire4056 = ( n_n56  &  wire72 ) | ( n_n56  &  n_n258  &  wire905 ) ;
 assign wire4059 = ( n_n151  &  n_n56 ) | ( n_n56  &  wire75 ) | ( n_n56  &  n_n206 ) ;
 assign wire4060 = ( n_n57  &  wire225 ) | ( n_n57  &  wire130 ) ;
 assign wire4062 = ( n_n48  &  wire79 ) | ( n_n48  &  wire905  &  n_n256 ) ;
 assign wire4071 = ( n_n1  &  wire225 ) | ( n_n1  &  wire130 ) ;
 assign wire4072 = ( n_n2  &  wire75 ) | ( n_n2  &  n_n206 ) | ( n_n2  &  wire20806 ) ;
 assign wire4073 = ( n_n268  &  wire20807 ) | ( n_n268  &  wire20808 ) ;
 assign wire4076 = ( n_n3  &  wire20796 ) | ( n_n3  &  wire20797 ) ;
 assign wire4080 = ( n_n3  &  n_n70 ) | ( n_n3  &  wire79 ) | ( n_n3  &  wire20791 ) ;
 assign wire4081 = ( n_n4  &  wire19738 ) | ( n_n4  &  wire913  &  n_n256 ) ;
 assign wire4089 = ( n_n151  &  n_n3 ) | ( n_n3  &  wire75 ) | ( n_n3  &  n_n206 ) ;
 assign wire4090 = ( n_n4  &  wire225 ) | ( n_n4  &  wire130 ) ;
 assign wire4100 = ( n_n100  &  wire118 ) | ( n_n100  &  wire899  &  n_n220 ) ;
 assign wire4117 = ( n_n94  &  n_n20 ) | ( n_n94  &  wire79 ) | ( n_n94  &  wire83 ) ;
 assign wire4120 = ( n_n100  &  wire79 ) | ( n_n100  &  wire899  &  n_n256 ) ;
 assign wire4131 = ( n_n100  &  wire66 ) | ( n_n100  &  n_n222  &  wire905 ) ;
 assign wire4159 = ( wire250  &  wire1231 ) | ( wire899  &  n_n281  &  wire1231 ) ;
 assign wire4166 = ( n_n152  &  wire103 ) | ( n_n152  &  n_n220  &  wire905 ) ;
 assign wire4170 = ( wire250  &  wire1141 ) | ( wire899  &  n_n281  &  wire1141 ) ;
 assign wire4183 = ( n_n6  &  wire57 ) | ( n_n6  &  n_n279  &  wire914 ) ;
 assign wire4196 = ( wire99  &  n_n230  &  n_n261  &  n_n285 ) ;
 assign wire4202 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) ;
 assign wire4234 = ( wire216  &  n_n132 ) | ( wire216  &  wire20637 ) | ( wire216  &  wire20638 ) ;
 assign wire4235 = ( wire899  &  n_n281  &  wire20637 ) | ( wire899  &  n_n281  &  wire20638 ) ;
 assign wire4236 = ( n_n163  &  n_n260  &  n_n283  &  n_n165 ) ;
 assign wire4248 = ( n_n4  &  wire101 ) | ( n_n4  &  n_n281  &  wire914 ) ;
 assign wire4259 = ( n_n151  &  n_n4 ) | ( n_n4  &  wire75 ) | ( n_n4  &  n_n206 ) ;
 assign wire4264 = ( n_n4  &  wire50 ) | ( n_n4  &  n_n59 ) | ( n_n4  &  wire113 ) ;
 assign wire4267 = ( n_n106  &  n_n265 ) | ( n_n265  &  wire268 ) | ( n_n265  &  wire101 ) ;
 assign wire4276 = ( n_n1  &  wire440 ) | ( n_n1  &  wire20601 ) | ( n_n1  &  wire20602 ) ;
 assign wire4281 = ( n_n1  &  wire20595 ) | ( n_n1  &  wire20596 ) | ( n_n1  &  wire20597 ) ;
 assign wire4285 = ( n_n4  &  n_n73 ) | ( n_n4  &  wire19408 ) | ( n_n4  &  wire20585 ) ;
 assign wire4302 = ( n_n4  &  n_n20 ) | ( n_n4  &  wire79 ) | ( n_n4  &  wire66 ) ;
 assign wire4313 = ( n_n1  &  n_n111 ) | ( n_n1  &  n_n32 ) | ( n_n1  &  wire85 ) ;
 assign wire4319 = ( n_n1  &  wire20555 ) | ( n_n1  &  wire20556 ) | ( n_n1  &  wire20557 ) ;
 assign wire4322 = ( n_n57  &  wire20547 ) | ( n_n57  &  wire20548 ) ;
 assign wire4330 = ( n_n100  &  wire19578 ) | ( n_n100  &  n_n222  &  wire906 ) ;
 assign wire4344 = ( n_n100  &  wire20528 ) | ( n_n100  &  wire20529 ) | ( n_n100  &  wire20530 ) ;
 assign wire4360 = ( n_n100  &  wire20512 ) | ( n_n100  &  wire20513 ) | ( n_n100  &  wire20514 ) ;
 assign wire4365 = ( n_n100  &  wire62 ) | ( n_n100  &  n_n15 ) | ( n_n100  &  wire20505 ) ;
 assign wire4373 = ( n_n57  &  n_n42 ) | ( n_n57  &  wire81 ) | ( n_n57  &  wire55 ) ;
 assign wire4380 = ( n_n100  &  wire137 ) | ( n_n100  &  wire113 ) ;
 assign wire4384 = ( n_n57  &  wire20490 ) | ( n_n57  &  wire20491 ) ;
 assign wire4391 = ( n_n57  &  wire85 ) | ( n_n57  &  n_n220  &  wire914 ) ;
 assign wire4409 = ( n_n53  &  wire20470 ) | ( n_n53  &  wire20471 ) | ( n_n53  &  wire20472 ) ;
 assign wire4414 = ( n_n57  &  wire20465 ) | ( n_n57  &  wire20466 ) | ( n_n57  &  wire20467 ) ;
 assign wire4417 = ( n_n57  &  wire75 ) | ( n_n57  &  n_n281  &  wire913 ) ;
 assign wire4418 = ( n_n264  &  n_n261  &  n_n267  &  n_n285 ) ;
 assign wire4423 = ( n_n6  &  wire19578 ) | ( n_n6  &  n_n222  &  wire906 ) ;
 assign wire4435 = ( n_n6  &  wire40 ) | ( n_n6  &  wire899  &  n_n258 ) ;
 assign wire4444 = ( n_n6  &  wire51 ) | ( n_n6  &  n_n41 ) | ( n_n6  &  wire20433 ) ;
 assign wire4453 = ( n_n53  &  wire50 ) | ( n_n53  &  n_n59 ) | ( n_n53  &  wire20423 ) ;
 assign wire4463 = ( n_n53  &  wire20414 ) | ( n_n53  &  wire20415 ) | ( n_n53  &  wire20416 ) ;
 assign wire4470 = ( n_n4  &  wire51 ) | ( n_n4  &  n_n43 ) | ( n_n4  &  wire59 ) ;
 assign wire4472 = ( n_n4  &  wire80 ) | ( n_n4  &  wire902  &  n_n256 ) ;
 assign wire4478 = ( n_n4  &  wire66 ) | ( n_n4  &  n_n222  &  wire905 ) ;
 assign wire4492 = ( n_n207  &  n_n17 ) | ( n_n207  &  wire514 ) | ( n_n207  &  wire20365 ) ;
 assign wire4500 = ( n_n6  &  wire20358 ) | ( n_n6  &  wire20359 ) ;
 assign wire4506 = ( n_n6  &  n_n10 ) | ( n_n6  &  wire137 ) | ( n_n6  &  wire113 ) ;
 assign wire4520 = ( n_n53  &  wire225 ) | ( n_n53  &  wire130 ) ;
 assign wire4523 = ( n_n48  &  wire20313 ) | ( n_n48  &  wire20314 ) ;
 assign wire4524 = ( n_n53  &  wire20315 ) | ( n_n53  &  wire20316 ) ;
 assign wire4529 = ( n_n53  &  wire368 ) | ( n_n53  &  n_n88 ) | ( n_n53  &  wire20306 ) ;
 assign wire4530 = ( n_n48  &  wire20308 ) | ( n_n48  &  wire20309 ) ;
 assign wire4551 = ( n_n53  &  wire246 ) | ( n_n53  &  wire256 ) ;
 assign wire4552 = ( n_n48  &  wire117 ) | ( n_n48  &  wire20289 ) | ( n_n48  &  wire20290 ) ;
 assign wire4557 = ( n_n53  &  wire62 ) | ( n_n53  &  wire105 ) | ( n_n53  &  wire20284 ) ;
 assign wire4558 = ( n_n48  &  n_n16 ) | ( n_n48  &  wire20155 ) | ( n_n48  &  wire20284 ) ;
 assign wire4565 = ( n_n48  &  wire113 ) | ( n_n48  &  wire101 ) ;
 assign wire4569 = ( n_n48  &  n_n7 ) | ( n_n48  &  wire50 ) | ( n_n48  &  n_n59 ) ;
 assign wire4570 = ( n_n53  &  wire50 ) | ( n_n53  &  n_n228  &  wire897 ) ;
 assign wire4573 = ( n_n48  &  n_n65 ) | ( n_n48  &  wire73 ) | ( n_n48  &  wire83 ) ;
 assign wire4574 = ( n_n53  &  wire44 ) | ( n_n53  &  n_n252 ) | ( n_n53  &  n_n15 ) ;
 assign wire4586 = ( n_n48  &  n_n80 ) | ( n_n48  &  wire88 ) | ( n_n48  &  wire20258 ) ;
 assign wire4587 = ( n_n53  &  wire74 ) | ( n_n53  &  wire903  &  n_n225 ) ;
 assign wire4593 = ( n_n53  &  wire66 ) | ( n_n53  &  n_n222  &  wire905 ) ;
 assign wire4602 = ( n_n53  &  n_n34 ) | ( n_n53  &  n_n82 ) | ( n_n53  &  wire47 ) ;
 assign wire4617 = ( i_7_  &  i_6_  &  wire1829 ) | ( (~ i_7_)  &  i_6_  &  wire1829 ) ;
 assign wire4618 = ( i_7_  &  i_6_  &  n_n118  &  n_n284 ) ;
 assign wire4636 = ( n_n132  &  wire1575 ) | ( wire1575  &  wire20213 ) ;
 assign wire4641 = ( wire1797  &  wire1796 ) ;
 assign wire4655 = ( n_n57  &  n_n179 ) | ( n_n57  &  wire57 ) | ( n_n57  &  wire20195 ) ;
 assign wire4656 = ( n_n56  &  wire89 ) | ( n_n56  &  n_n222  &  wire907 ) ;
 assign wire4679 = ( n_n6  &  n_n148 ) | ( n_n6  &  wire246 ) | ( n_n6  &  wire20179 ) ;
 assign wire4680 = ( n_n5  &  wire101 ) | ( n_n5  &  wire20180 ) | ( n_n5  &  wire20182 ) ;
 assign wire4684 = ( n_n5  &  n_n148 ) | ( n_n5  &  wire113 ) | ( n_n5  &  wire20171 ) ;
 assign wire4685 = ( n_n6  &  n_n63 ) | ( n_n6  &  wire199 ) | ( n_n6  &  wire20173 ) ;
 assign wire4690 = ( n_n151  &  n_n5 ) | ( n_n5  &  wire75 ) | ( n_n5  &  n_n206 ) ;
 assign wire4691 = ( n_n6  &  wire225 ) | ( n_n6  &  wire911  &  n_n220 ) ;
 assign wire4694 = ( n_n5  &  n_n20 ) | ( n_n5  &  wire79 ) | ( n_n5  &  wire83 ) ;
 assign wire4695 = ( n_n6  &  wire44 ) | ( n_n6  &  n_n252 ) | ( n_n6  &  n_n15 ) ;
 assign wire4696 = ( n_n5  &  wire20160 ) | ( n_n5  &  wire20161 ) ;
 assign wire4704 = ( n_n5  &  wire62 ) | ( n_n5  &  wire1781 ) ;
 assign wire4705 = ( n_n6  &  wire1781 ) | ( n_n6  &  wire20156 ) ;
 assign wire4710 = ( n_n5  &  n_n203 ) | ( n_n5  &  wire20149 ) | ( n_n5  &  wire20150 ) ;
 assign wire4711 = ( n_n6  &  wire79 ) | ( n_n6  &  wire899  &  n_n256 ) ;
 assign wire4720 = ( n_n6  &  n_n43 ) | ( n_n6  &  wire59 ) | ( n_n6  &  wire20144 ) ;
 assign wire4726 = ( n_n6  &  n_n34 ) | ( n_n6  &  wire86 ) | ( n_n6  &  wire20136 ) ;
 assign wire4727 = ( n_n5  &  wire87 ) | ( n_n5  &  wire914  &  n_n225 ) ;
 assign wire4735 = ( n_n5  &  wire20132 ) | ( n_n5  &  wire20133 ) ;
 assign wire4745 = ( n_n5  &  n_n97 ) | ( n_n5  &  wire77 ) | ( n_n5  &  wire71 ) ;
 assign wire4750 = ( n_n6  &  n_n105 ) | ( n_n6  &  n_n97 ) | ( n_n6  &  wire71 ) ;
 assign wire4751 = ( n_n5  &  wire20125 ) | ( n_n5  &  wire20126 ) ;
 assign wire4756 = ( n_n57  &  wire95 ) | ( n_n57  &  n_n281  &  wire914 ) ;
 assign wire4761 = ( n_n56  &  wire75 ) | ( n_n56  &  n_n281  &  wire913 ) ;
 assign wire4766 = ( n_n151  &  n_n94 ) | ( n_n94  &  n_n206 ) | ( n_n94  &  wire20107 ) ;
 assign wire4789 = ( n_n151  &  n_n100 ) | ( n_n100  &  wire75 ) | ( n_n100  &  n_n206 ) ;
 assign wire4790 = ( n_n260  &  n_n263  &  n_n285  &  wire130 ) ;
 assign wire4800 = ( n_n94  &  wire20089 ) | ( n_n94  &  wire20090 ) ;
 assign wire4805 = ( n_n94  &  wire20086 ) | ( n_n94  &  wire20087 ) ;
 assign wire4807 = ( wire200  &  n_n100 ) | ( n_n100  &  wire157 ) | ( n_n100  &  wire273 ) ;
 assign wire4808 = ( wire268  &  n_n94 ) | ( wire200  &  n_n94 ) | ( n_n94  &  wire277 ) ;
 assign wire4817 = ( n_n94  &  wire190 ) | ( n_n94  &  wire119 ) | ( n_n94  &  wire198 ) ;
 assign wire4827 = ( n_n260  &  n_n261  &  n_n285  &  wire1662 ) ;
 assign wire4839 = ( n_n94  &  n_n63 ) | ( n_n94  &  wire246 ) | ( n_n94  &  wire20051 ) ;
 assign wire4844 = ( n_n100  &  n_n12 ) | ( n_n100  &  n_n65 ) | ( n_n100  &  wire73 ) ;
 assign wire4845 = ( n_n94  &  n_n14 ) | ( n_n94  &  wire70 ) | ( n_n94  &  wire256 ) ;
 assign wire4849 = ( n_n94  &  wire123 ) | ( n_n94  &  wire100 ) | ( n_n94  &  wire227 ) ;
 assign wire4856 = ( n_n60  &  n_n94 ) | ( n_n94  &  n_n9 ) | ( n_n94  &  wire63 ) ;
 assign wire4869 = ( n_n100  &  n_n60 ) | ( n_n100  &  wire137 ) | ( n_n100  &  wire63 ) ;
 assign wire4870 = ( n_n94  &  n_n7 ) | ( n_n94  &  wire50 ) | ( n_n94  &  n_n59 ) ;
 assign wire4871 = ( (~ i_7_)  &  i_6_  &  n_n165  &  wire19294 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19294 ) ;
 assign wire4882 = ( n_n118  &  n_n231  &  n_n264 ) | ( n_n118  &  n_n231  &  n_n230 ) ;
 assign wire4889 = ( wire48  &  n_n128 ) | ( n_n128  &  wire913  &  n_n220 ) ;
 assign wire4890 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) ;
 assign wire4892 = ( n_n163  &  n_n273  &  n_n165  &  wire19296 ) ;
 assign wire4896 = ( wire48  &  wire1079 ) | ( wire913  &  n_n220  &  wire1079 ) ;
 assign wire4899 = ( wire48  &  n_n152 ) | ( n_n152  &  wire913  &  n_n220 ) ;
 assign wire4900 = ( i_7_  &  i_6_  &  n_n165  &  wire19294 ) | ( (~ i_7_)  &  i_6_  &  n_n165  &  wire19294 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19294 ) ;
 assign wire4902 = ( wire48  &  wire1076 ) | ( wire913  &  n_n220  &  wire1076 ) ;
 assign wire4905 = ( wire949  &  n_n128 ) | ( wire949  &  n_n122 ) ;
 assign wire4928 = ( i_7_  &  i_6_  &  n_n118  &  n_n260 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n260 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n260 ) ;
 assign wire4935 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) ;
 assign wire4939 = ( n_n56  &  wire153 ) | ( n_n56  &  wire41 ) ;
 assign wire4947 = ( n_n128  &  wire54 ) | ( n_n128  &  wire913  &  n_n220 ) ;
 assign wire4974 = ( n_n56  &  wire61 ) | ( n_n56  &  n_n279  &  wire908 ) ;
 assign wire5002 = ( n_n57  &  wire95 ) | ( n_n57  &  n_n281  &  wire914 ) ;
 assign wire5011 = ( n_n106  &  n_n56 ) | ( n_n56  &  n_n62 ) | ( n_n56  &  wire101 ) ;
 assign wire5012 = ( n_n266  &  n_n230  &  n_n285  &  wire101 ) ;
 assign wire5013 = ( n_n56  &  wire95 ) | ( n_n56  &  n_n281  &  wire914 ) ;
 assign wire5014 = ( n_n57  &  wire63 ) | ( n_n57  &  n_n228  &  wire902 ) ;
 assign wire5023 = ( n_n56  &  wire75 ) | ( n_n56  &  n_n281  &  wire913 ) ;
 assign wire5031 = ( n_n57  &  wire118 ) | ( n_n57  &  wire72 ) ;
 assign wire5033 = ( n_n151  &  n_n57 ) | ( n_n57  &  wire75 ) | ( n_n57  &  n_n206 ) ;
 assign wire5035 = ( n_n57  &  n_n7 ) | ( n_n57  &  wire50 ) | ( n_n57  &  n_n59 ) ;
 assign wire5036 = ( n_n230  &  n_n271  &  n_n285  &  wire132 ) ;
 assign wire5047 = ( n_n6  &  wire80 ) | ( n_n6  &  n_n256  &  wire908 ) ;
 assign wire5048 = ( n_n5  &  wire57 ) | ( n_n5  &  n_n279  &  wire912 ) ;
 assign wire5053 = ( n_n5  &  wire19892 ) | ( n_n5  &  wire19893 ) ;
 assign wire5054 = ( n_n6  &  wire42 ) | ( n_n6  &  n_n279  &  wire899 ) ;
 assign wire5059 = ( n_n6  &  wire50 ) | ( n_n6  &  n_n281  &  wire903 ) ;
 assign wire5060 = ( n_n5  &  wire63 ) | ( n_n5  &  n_n228  &  wire902 ) ;
 assign wire5075 = ( n_n5  &  n_n12 ) | ( n_n5  &  wire73 ) | ( n_n5  &  wire19874 ) ;
 assign wire5076 = ( n_n6  &  wire95 ) | ( n_n6  &  n_n281  &  wire914 ) ;
 assign wire5091 = ( n_n6  &  wire55 ) | ( n_n6  &  n_n279  &  wire912 ) ;
 assign wire5099 = ( n_n6  &  wire273 ) | ( n_n6  &  wire914  &  n_n225 ) ;
 assign wire5109 = ( n_n268  &  wire19852 ) | ( n_n268  &  wire19853 ) ;
 assign wire5115 = ( n_n265  &  wire101 ) | ( n_n265  &  n_n281  &  wire907 ) ;
 assign wire5116 = ( n_n268  &  n_n11 ) | ( n_n268  &  wire95 ) | ( n_n268  &  wire19848 ) ;
 assign wire5138 = ( n_n124  &  wire48 ) | ( n_n124  &  n_n110 ) | ( n_n124  &  n_n163 ) ;
 assign wire5140 = ( wire48  &  n_n122 ) | ( n_n108  &  n_n122 ) | ( n_n122  &  wire19833 ) ;
 assign wire5144 = ( n_n264  &  n_n163  &  n_n229  &  n_n165 ) ;
 assign wire5153 = ( n_n2  &  wire19817 ) | ( n_n2  &  wire19818 ) ;
 assign wire5160 = ( n_n2  &  wire137 ) | ( n_n2  &  wire132 ) ;
 assign wire5161 = ( n_n1  &  n_n7 ) | ( n_n1  &  wire50 ) | ( n_n1  &  wire19814 ) ;
 assign wire5171 = ( n_n2  &  n_n95 ) | ( n_n2  &  wire85 ) | ( n_n2  &  wire19801 ) ;
 assign wire5184 = ( n_n2  &  n_n11 ) | ( n_n2  &  n_n148 ) | ( n_n2  &  wire95 ) ;
 assign wire5185 = ( n_n1  &  n_n11 ) | ( n_n1  &  wire113 ) | ( n_n1  &  wire19790 ) ;
 assign wire5195 = ( n_n2  &  wire913  &  n_n220 ) ;
 assign wire5205 = ( n_n1  &  n_n148 ) | ( n_n1  &  wire101 ) | ( n_n1  &  wire95 ) ;
 assign wire5208 = ( n_n2  &  wire19773 ) | ( n_n2  &  wire19774 ) ;
 assign wire5215 = ( n_n2  &  wire453 ) | ( n_n2  &  n_n256  &  wire914 ) ;
 assign wire5219 = ( n_n2  &  n_n220  &  wire914 ) ;
 assign wire5228 = ( n_n6  &  wire80 ) | ( n_n6  &  n_n256  &  wire908 ) ;
 assign wire5238 = ( n_n6  &  n_n32 ) | ( n_n6  &  n_n81 ) | ( n_n6  &  wire86 ) ;
 assign wire5239 = ( n_n230  &  n_n263  &  n_n285  &  wire55 ) ;
 assign wire5240 = ( n_n5  &  n_n171 ) | ( n_n5  &  wire56 ) | ( n_n5  &  wire53 ) ;
 assign wire5241 = ( n_n6  &  n_n220  &  wire908 ) ;
 assign wire5242 = ( n_n5  &  n_n73 ) | ( n_n5  &  n_n22 ) | ( n_n5  &  wire19408 ) ;
 assign wire5243 = ( n_n230  &  n_n261  &  n_n285  &  wire56 ) ;
 assign wire5244 = ( n_n6  &  wire89 ) | ( n_n6  &  n_n83 ) | ( n_n6  &  wire85 ) ;
 assign wire5245 = ( n_n5  &  n_n220  &  wire907 ) ;
 assign wire5248 = ( n_n5  &  n_n204 ) | ( n_n5  &  wire52 ) | ( n_n5  &  wire19744 ) ;
 assign wire5262 = ( n_n6  &  wire19738 ) | ( n_n6  &  wire913  &  n_n256 ) ;
 assign wire5268 = ( n_n5  &  wire82 ) | ( n_n5  &  n_n223 ) | ( n_n5  &  wire42 ) ;
 assign wire5269 = ( n_n6  &  wire913  &  n_n220 ) ;
 assign wire5298 = ( n_n56  &  wire19711 ) | ( n_n56  &  wire19712 ) ;
 assign wire5299 = ( n_n57  &  wire19713 ) | ( n_n57  &  wire19714 ) ;
 assign wire5327 = ( n_n56  &  wire160 ) | ( n_n56  &  n_n60 ) | ( n_n56  &  wire63 ) ;
 assign wire5328 = ( n_n57  &  n_n144 ) | ( n_n57  &  wire118 ) | ( n_n57  &  wire19693 ) ;
 assign wire5336 = ( n_n56  &  wire100 ) | ( n_n56  &  wire210 ) | ( n_n56  &  wire19691 ) ;
 assign wire5340 = ( n_n57  &  wire160 ) | ( n_n57  &  n_n66 ) | ( n_n57  &  wire19682 ) ;
 assign wire5341 = ( n_n56  &  wire246 ) | ( n_n56  &  wire19683 ) | ( n_n56  &  wire19685 ) ;
 assign wire5343 = ( n_n56  &  n_n14 ) | ( n_n56  &  wire70 ) | ( n_n56  &  wire256 ) ;
 assign wire5344 = ( n_n57  &  n_n12 ) | ( n_n57  &  n_n65 ) | ( n_n57  &  wire73 ) ;
 assign wire5347 = ( n_n6  &  wire50 ) | ( n_n6  &  n_n281  &  wire903 ) ;
 assign wire5348 = ( n_n5  &  wire63 ) | ( n_n5  &  n_n228  &  wire902 ) ;
 assign wire5356 = ( n_n6  &  n_n42 ) | ( n_n6  &  wire43 ) | ( n_n6  &  wire19674 ) ;
 assign wire5357 = ( n_n5  &  wire43 ) | ( n_n5  &  wire19674 ) | ( n_n5  &  wire19675 ) ;
 assign wire5361 = ( n_n6  &  n_n102 ) | ( n_n6  &  wire807 ) | ( n_n6  &  wire71 ) ;
 assign wire5362 = ( n_n56  &  wire225 ) | ( n_n56  &  wire130 ) ;
 assign wire5363 = ( n_n151  &  n_n57 ) | ( n_n57  &  wire75 ) | ( n_n57  &  wire19668 ) ;
 assign wire5368 = ( n_n56  &  n_n145 ) | ( n_n56  &  n_n144 ) | ( n_n56  &  wire118 ) ;
 assign wire5369 = ( n_n6  &  wire96 ) | ( n_n6  &  n_n222  &  wire904 ) ;
 assign wire5371 = ( n_n5  &  n_n49 ) | ( n_n5  &  wire71 ) | ( n_n5  &  wire19661 ) ;
 assign wire5372 = ( n_n6  &  wire55 ) | ( n_n6  &  wire453 ) | ( n_n6  &  wire19663 ) ;
 assign wire5381 = ( n_n5  &  n_n101 ) | ( n_n5  &  wire61 ) | ( n_n5  &  wire19657 ) ;
 assign wire5389 = ( n_n5  &  wire101 ) | ( n_n5  &  wire901  &  n_n220 ) ;
 assign wire5390 = ( n_n6  &  wire95 ) | ( n_n6  &  n_n281  &  wire914 ) ;
 assign wire5400 = ( n_n6  &  wire113 ) | ( n_n6  &  wire101 ) ;
 assign wire5405 = ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19294 ) ;
 assign wire5408 = ( (~ i_7_)  &  i_6_  &  n_n165  &  wire19294 ) ;
 assign wire5411 = ( i_7_  &  i_6_  &  wire943 ) | ( i_7_  &  (~ i_6_)  &  wire943 ) ;
 assign wire5412 = ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n284 ) ;
 assign wire5413 = ( i_7_  &  i_6_  &  n_n118  &  n_n284 ) ;
 assign wire5421 = ( n_n152  &  wire54 ) | ( n_n152  &  n_n220  &  wire914 ) ;
 assign wire5426 = ( n_n130  &  wire54 ) | ( n_n121  &  wire54 ) | ( n_n122  &  wire54 ) ;
 assign wire5430 = ( wire54  &  wire1687 ) | ( n_n220  &  wire914  &  wire1687 ) ;
 assign wire5439 = ( wire923  &  n_n283  &  n_n165  &  wire19294 ) ;
 assign wire5441 = ( wire923  &  n_n283  &  n_n165  &  wire19296 ) ;
 assign wire5442 = ( n_n163  &  n_n273  &  n_n165  &  wire19296 ) ;
 assign wire5445 = ( n_n124  &  n_n111 ) | ( n_n124  &  wire103 ) | ( n_n124  &  wire266 ) ;
 assign wire5453 = ( i_7_  &  i_6_  &  n_n118  &  n_n264 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n264 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n264 ) ;
 assign wire5457 = ( n_n127  &  wire419 ) | ( n_n127  &  wire19605 ) | ( n_n127  &  wire19608 ) ;
 assign wire5472 = ( n_n94  &  wire19578 ) | ( n_n94  &  n_n222  &  wire906 ) ;
 assign wire5478 = ( n_n94  &  n_n43 ) | ( n_n94  &  wire59 ) | ( n_n94  &  wire19579 ) ;
 assign wire5485 = ( n_n94  &  n_n78 ) | ( n_n94  &  wire80 ) | ( n_n94  &  wire19567 ) ;
 assign wire5494 = ( n_n94  &  n_n281  &  wire908 ) ;
 assign wire5506 = ( n_n57  &  wire96 ) | ( n_n57  &  n_n222  &  wire904 ) ;
 assign wire5509 = ( n_n100  &  n_n7 ) | ( n_n100  &  wire50 ) | ( n_n100  &  n_n59 ) ;
 assign wire5510 = ( n_n94  &  wire137 ) | ( n_n94  &  wire132 ) | ( n_n94  &  wire19558 ) ;
 assign wire5514 = ( n_n100  &  wire246 ) | ( n_n100  &  wire256 ) ;
 assign wire5515 = ( n_n94  &  n_n65 ) | ( n_n94  &  wire73 ) | ( n_n94  &  wire19556 ) ;
 assign wire5516 = ( n_n94  &  n_n25 ) | ( n_n94  &  wire19457 ) | ( n_n94  &  wire19548 ) ;
 assign wire5517 = ( n_n100  &  wire80 ) | ( n_n100  &  wire902  &  n_n256 ) ;
 assign wire5544 = ( n_n56  &  wire61 ) | ( n_n56  &  n_n279  &  wire908 ) ;
 assign wire5546 = ( n_n230  &  n_n271  &  n_n285  &  wire56 ) ;
 assign wire5550 = ( n_n57  &  wire73 ) | ( n_n57  &  wire900  &  n_n228 ) ;
 assign wire5552 = ( n_n56  &  n_n12 ) | ( n_n56  &  n_n65 ) | ( n_n56  &  wire73 ) ;
 assign wire5564 = ( n_n48  &  wire68 ) | ( n_n48  &  n_n49 ) | ( n_n48  &  wire71 ) ;
 assign wire5565 = ( n_n53  &  n_n42 ) | ( n_n53  &  n_n90 ) | ( n_n53  &  wire19384 ) ;
 assign wire5569 = ( n_n53  &  wire81 ) | ( n_n53  &  n_n93 ) | ( n_n53  &  wire76 ) ;
 assign wire5570 = ( n_n48  &  wire19507 ) | ( n_n48  &  wire19508 ) ;
 assign wire5577 = ( n_n56  &  wire63 ) | ( n_n56  &  n_n281  &  wire908 ) ;
 assign wire5587 = ( n_n56  &  n_n7 ) | ( n_n56  &  wire50 ) | ( n_n56  &  n_n59 ) ;
 assign wire5588 = ( n_n266  &  n_n230  &  n_n285  &  wire137 ) ;
 assign wire5589 = ( n_n56  &  wire44 ) | ( n_n56  &  wire70 ) ;
 assign wire5590 = ( n_n57  &  n_n281  &  wire906 ) ;
 assign wire5591 = ( n_n264  &  n_n253  &  n_n263  &  n_n285 ) ;
 assign wire5592 = ( n_n264  &  n_n261  &  n_n267  &  n_n285 ) ;
 assign wire5595 = ( n_n48  &  wire19497 ) | ( n_n48  &  wire19498 ) ;
 assign wire5596 = ( n_n53  &  wire53 ) | ( n_n53  &  n_n279  &  wire897 ) ;
 assign wire5606 = ( n_n53  &  wire137 ) | ( n_n53  &  wire132 ) ;
 assign wire5607 = ( n_n48  &  wire44 ) | ( n_n48  &  wire19491 ) | ( n_n48  &  wire19493 ) ;
 assign wire5611 = ( wire99  &  n_n230  &  n_n261  &  n_n285 ) ;
 assign wire5613 = ( n_n6  &  wire41 ) | ( n_n6  &  n_n279  &  wire898 ) ;
 assign wire5617 = ( n_n53  &  wire70 ) | ( n_n53  &  wire903  &  n_n220 ) ;
 assign wire5625 = ( n_n48  &  n_n12 ) | ( n_n48  &  wire70 ) | ( n_n48  &  wire73 ) ;
 assign wire5626 = ( n_n53  &  n_n12 ) | ( n_n53  &  n_n65 ) | ( n_n53  &  wire73 ) ;
 assign wire5629 = ( wire224  &  n_n230  &  n_n261  &  n_n285 ) ;
 assign wire5636 = ( n_n230  &  n_n261  &  n_n285  &  wire1552 ) ;
 assign wire5637 = ( n_n5  &  wire140 ) | ( n_n5  &  wire198 ) | ( n_n5  &  wire1554 ) ;
 assign wire5640 = ( n_n80  &  n_n227 ) | ( wire114  &  n_n227 ) | ( n_n227  &  wire88 ) ;
 assign wire5642 = ( n_n5  &  wire50 ) | ( n_n5  &  n_n281  &  wire903 ) ;
 assign wire5643 = ( n_n6  &  wire50 ) | ( n_n6  &  n_n228  &  wire897 ) ;
 assign wire5650 = ( n_n5  &  wire165 ) | ( n_n5  &  wire167 ) ;
 assign wire5651 = ( n_n6  &  n_n14 ) | ( n_n6  &  wire70 ) | ( n_n6  &  wire199 ) ;
 assign wire5656 = ( n_n5  &  wire246 ) | ( n_n5  &  wire256 ) ;
 assign wire5657 = ( n_n6  &  n_n12 ) | ( n_n6  &  wire73 ) | ( n_n6  &  wire19469 ) ;
 assign wire5660 = ( n_n4  &  wire166 ) | ( n_n4  &  n_n225  &  wire908 ) ;
 assign wire5661 = ( n_n94  &  wire50 ) | ( n_n94  &  n_n281  &  wire903 ) ;
 assign wire5671 = ( wire120  &  n_n207 ) | ( n_n207  &  n_n25 ) | ( n_n207  &  wire19457 ) ;
 assign wire5681 = ( n_n4  &  wire153 ) | ( n_n4  &  wire180 ) ;
 assign wire5682 = ( n_n229  &  wire254  &  n_n285  &  n_n284 ) ;
 assign wire5683 = ( n_n229  &  n_n285  &  n_n284  &  wire1786 ) ;
 assign wire5699 = ( n_n1  &  wire70 ) | ( n_n1  &  n_n228  &  wire902 ) ;
 assign wire5700 = ( n_n2  &  n_n220  &  wire908 ) ;
 assign wire5709 = ( n_n2  &  wire44 ) | ( n_n2  &  wire70 ) ;
 assign wire5710 = ( n_n1  &  n_n281  &  wire906 ) ;
 assign wire5711 = ( n_n1  &  wire80 ) | ( n_n1  &  n_n256  &  wire908 ) ;
 assign wire5718 = ( n_n1  &  wire73 ) | ( n_n1  &  wire900  &  n_n228 ) ;
 assign wire5720 = ( n_n2  &  n_n12 ) | ( n_n2  &  n_n65 ) | ( n_n2  &  wire73 ) ;
 assign wire5721 = ( wire44  &  n_n260  &  n_n273  &  n_n285 ) ;
 assign wire5725 = ( n_n2  &  n_n29 ) | ( n_n2  &  wire49 ) | ( n_n2  &  wire88 ) ;
 assign wire5726 = ( n_n1  &  n_n73 ) | ( n_n1  &  n_n22 ) | ( n_n1  &  wire19408 ) ;
 assign wire5728 = ( n_n3  &  wire19417 ) | ( n_n3  &  wire19418 ) ;
 assign wire5733 = ( n_n3  &  wire19409 ) | ( n_n3  &  wire19410 ) ;
 assign wire5734 = ( n_n4  &  wire61 ) | ( n_n4  &  n_n279  &  wire908 ) ;
 assign wire5743 = ( n_n4  &  wire137 ) | ( n_n4  &  wire132 ) ;
 assign wire5744 = ( n_n3  &  n_n60 ) | ( n_n3  &  wire63 ) | ( n_n3  &  wire19403 ) ;
 assign wire5749 = ( n_n1  &  wire137 ) | ( n_n1  &  wire132 ) ;
 assign wire5750 = ( n_n2  &  n_n60 ) | ( n_n2  &  wire63 ) | ( n_n2  &  wire19395 ) ;
 assign wire5754 = ( n_n4  &  wire88 ) | ( n_n4  &  n_n222  &  wire908 ) ;
 assign wire5758 = ( n_n4  &  wire19384 ) | ( n_n4  &  n_n281  &  wire900 ) ;
 assign wire5775 = ( n_n3  &  wire81 ) | ( n_n3  &  n_n93 ) | ( n_n3  &  wire76 ) ;
 assign wire5778 = ( n_n268  &  n_n7 ) | ( n_n268  &  wire50 ) | ( n_n268  &  wire119 ) ;
 assign wire5780 = ( n_n3  &  n_n12 ) | ( n_n3  &  n_n65 ) | ( n_n3  &  wire73 ) ;
 assign wire5797 = ( n_n139  &  wire48 ) | ( n_n139  &  wire913  &  n_n220 ) ;
 assign wire5812 = ( i_7_  &  i_6_  &  n_n118  &  n_n260 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n260 ) ;
 assign wire5813 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire5824 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire19350 ) ;
 assign wire5834 = ( n_n223  &  n_n122 ) | ( n_n122  &  wire214 ) | ( n_n122  &  wire19344 ) ;
 assign wire5835 = ( n_n123  &  wire19347 ) | ( n_n123  &  wire19348 ) ;
 assign wire5843 = ( n_n124  &  n_n253 ) | ( n_n124  &  n_n143 ) | ( n_n124  &  wire214 ) ;
 assign wire5844 = ( n_n123  &  wire19342 ) | ( n_n123  &  n_n282  &  wire1074 ) ;
 assign wire5848 = ( n_n128  &  n_n147 ) | ( n_n128  &  wire328 ) | ( n_n128  &  wire19237 ) ;
 assign wire5849 = ( n_n127  &  wire397 ) | ( n_n127  &  wire19334 ) | ( n_n127  &  wire19337 ) ;
 assign wire5850 = ( n_n266  &  n_n165  &  n_n230 ) ;
 assign wire5854 = ( n_n127  &  wire72 ) | ( n_n127  &  wire352 ) | ( n_n127  &  wire19332 ) ;
 assign wire5855 = ( n_n273  &  n_n165  &  n_n284  &  wire384 ) ;
 assign wire5861 = ( n_n130  &  wire19329 ) | ( n_n130  &  wire19330 ) ;
 assign wire5862 = ( n_n208  &  n_n165  &  n_n230 ) ;
 assign wire5863 = ( n_n124  &  n_n150 ) | ( n_n124  &  wire326 ) | ( n_n124  &  wire19244 ) ;
 assign wire5874 = ( n_n264  &  n_n165  &  wire1226 ) ;
 assign wire5875 = ( n_n121  &  wire398 ) | ( n_n121  &  wire19308 ) | ( n_n121  &  wire19309 ) ;
 assign wire5876 = ( n_n122  &  wire19313 ) | ( n_n122  &  wire19314 ) ;
 assign wire5877 = ( n_n271  &  n_n285  &  n_n284  &  wire1186 ) ;
 assign wire5878 = ( n_n266  &  n_n285  &  n_n284  &  wire1187 ) ;
 assign wire5879 = ( (~ i_9_)  &  n_n264  &  n_n263  &  n_n285 ) ;
 assign wire5880 = ( i_9_  &  n_n264  &  n_n261  &  n_n285 ) ;
 assign wire5885 = ( n_n227  &  wire65 ) | ( n_n227  &  wire19220 ) | ( n_n227  &  wire19221 ) ;
 assign wire5893 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire1133 ) ;
 assign wire5900 = ( n_n207  &  wire19211 ) | ( n_n207  &  wire911  &  n_n228 ) ;
 assign wire5910 = ( i_6_  &  n_n264  &  n_n285 ) ;
 assign wire5922 = ( n_n241  &  wire19197 ) | ( n_n241  &  wire19198 ) ;
 assign wire5923 = ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n285 ) ;
 assign wire5931 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire969 ) ;
 assign wire5936 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire966 ) ;
 assign wire5941 = ( n_n130  &  n_n281  &  wire905 ) ;
 assign wire5953 = ( n_n132  &  n_n223 ) | ( n_n132  &  wire214 ) | ( n_n132  &  wire19252 ) ;
 assign wire5955 = ( n_n139  &  n_n150 ) | ( n_n139  &  wire326 ) | ( n_n139  &  wire19244 ) ;
 assign wire5957 = ( n_n142  &  wire19248 ) | ( n_n142  &  wire19249 ) ;
 assign wire5959 = ( n_n139  &  wire435 ) | ( n_n139  &  wire19240 ) | ( n_n139  &  wire19241 ) ;
 assign wire5960 = ( n_n283  &  n_n165  &  n_n230  &  wire326 ) ;
 assign wire5973 = ( i_6_  &  n_n165  &  wire19296 ) | ( i_7_  &  (~ i_6_)  &  n_n165  &  wire19296 ) ;
 assign wire5985 = ( i_9_  &  n_n273  &  n_n230  &  n_n285 ) ;
 assign wire5988 = ( i_5_  &  i_3_  &  n_n165  &  wire19291 ) ;
 assign wire5990 = ( n_n283  &  n_n230  &  n_n285  &  wire1223 ) ;
 assign wire5999 = ( (~ i_9_)  &  i_10_  &  i_12_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire6004 = ( i_9_  &  i_10_  &  i_12_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  i_11_ ) ;
 assign wire6008 = ( (~ i_11_)  &  wire923  &  n_n207 ) | ( i_11_  &  wire923  &  (~ n_n254)  &  n_n207 ) ;
 assign wire6009 = ( n_n189  &  wire6014 ) | ( n_n189  &  wire19274 ) | ( n_n189  &  wire19275 ) ;
 assign wire6014 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire197 ) ;
 assign wire6020 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire1183 ) ;
 assign wire19191 = ( wire913  &  n_n258 ) | ( wire903  &  n_n258 ) ;
 assign wire19192 = ( n_n267  &  wire965 ) | ( (~ i_15_)  &  n_n258  &  n_n267 ) ;
 assign wire19194 = ( (~ i_9_) ) | ( n_n258  &  wire914 ) ;
 assign wire19195 = ( n_n258  &  wire908 ) | ( n_n247  &  wire968 ) ;
 assign wire19197 = ( i_9_ ) | ( n_n258  &  wire907 ) ;
 assign wire19198 = ( i_11_  &  n_n163  &  wire148 ) | ( (~ i_11_)  &  n_n163  &  wire971 ) ;
 assign wire19205 = ( i_9_ ) | ( (~ i_9_)  &  i_10_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19206 = ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire19207 = ( n_n258  &  wire905 ) | ( n_n258  &  wire904 ) ;
 assign wire19208 = ( i_11_  &  n_n269  &  n_n256 ) | ( (~ i_11_)  &  n_n269  &  n_n256 ) | ( i_11_  &  n_n269  &  wire288 ) | ( (~ i_11_)  &  n_n269  &  wire288 ) ;
 assign wire19211 = ( n_n242  &  n_n225 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign wire19212 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire19213 = ( wire19212 ) | ( n_n228  &  wire903 ) ;
 assign wire19215 = ( i_9_  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  n_n256 ) ;
 assign wire19216 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire19217 = ( wire899  &  n_n228 ) | ( n_n258  &  wire908 ) ;
 assign wire19220 = ( n_n247 ) | ( wire911  &  n_n258 ) ;
 assign wire19221 = ( n_n242  &  wire148 ) | ( n_n270  &  wire1135 ) ;
 assign wire19223 = ( wire5900 ) | ( n_n227  &  wire1130 ) | ( n_n227  &  wire1132 ) ;
 assign wire19228 = ( wire5877 ) | ( wire5878 ) | ( wire5879 ) | ( wire5880 ) ;
 assign wire19230 = ( n_n5063 ) | ( wire19228 ) | ( wire916  &  wire1011 ) ;
 assign wire19233 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  n_n279 ) ;
 assign wire19235 = ( wire331 ) | ( wire19233 ) | ( wire911  &  n_n281 ) ;
 assign wire19236 = ( wire321 ) | ( wire454 ) | ( (~ i_9_)  &  (~ i_10_) ) ;
 assign wire19237 = ( i_12_  &  n_n247 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  n_n247 ) ;
 assign wire19238 = ( n_n267 ) | ( n_n279  &  wire912 ) ;
 assign wire19239 = ( n_n270 ) | ( n_n281  &  wire905 ) ;
 assign wire19240 = ( n_n253 ) | ( wire19237 ) | ( n_n220  &  wire912 ) ;
 assign wire19241 = ( n_n223 ) | ( n_n148 ) | ( wire19238 ) | ( wire19239 ) ;
 assign wire19243 = ( wire5960 ) | ( n_n136  &  wire19235 ) | ( n_n136  &  wire19236 ) ;
 assign wire19244 = ( i_12_  &  n_n242 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  n_n242 ) ;
 assign wire19245 = ( n_n253 ) | ( wire19237 ) | ( n_n220  &  wire912 ) ;
 assign wire19246 = ( n_n223 ) | ( n_n143 ) | ( wire214 ) | ( wire19239 ) ;
 assign wire19248 = ( wire331 ) | ( wire19233 ) | ( wire911  &  n_n281 ) ;
 assign wire19249 = ( wire321 ) | ( wire454 ) | ( (~ i_9_)  &  (~ i_10_) ) ;
 assign wire19250 = ( wire5955 ) | ( n_n152  &  wire19245 ) | ( n_n152  &  wire19246 ) ;
 assign wire19252 = ( wire196 ) | ( wire352 ) | ( n_n281  &  wire905 ) ;
 assign wire19253 = ( i_14_  &  n_n247  &  n_n278 ) | ( (~ i_14_)  &  i_15_  &  n_n247  &  n_n278 ) ;
 assign wire19254 = ( (~ i_9_)  &  (~ i_10_) ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign wire19255 = ( wire19254 ) | ( n_n281  &  wire914 ) ;
 assign wire19256 = ( wire19244 ) | ( wire19255 ) | ( wire911  &  n_n220 ) ;
 assign wire19258 = ( (~ i_9_) ) | ( i_9_  &  i_10_ ) | ( n_n281  &  wire912 ) ;
 assign wire19259 = ( wire196 ) | ( n_n247  &  wire152 ) ;
 assign wire19260 = ( wire5941 ) | ( n_n132  &  wire285 ) | ( n_n132  &  wire19256 ) ;
 assign wire19261 = ( wire5953 ) | ( n_n273  &  wire896 ) | ( wire896  &  wire1271 ) ;
 assign wire19263 = ( wire5957 ) | ( wire5959 ) | ( wire19243 ) | ( wire19250 ) ;
 assign wire19264 = ( i_9_  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire19265 = ( n_n275  &  n_n220 ) | ( n_n225  &  n_n270 ) ;
 assign wire19266 = ( wire19264 ) | ( wire899  &  n_n258 ) ;
 assign wire19267 = ( n_n228  &  wire908 ) | ( n_n259  &  wire148 ) ;
 assign wire19269 = ( n_n267 ) | ( wire903  &  n_n258 ) ;
 assign wire19270 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign wire19271 = ( n_n242  &  wire1182 ) | ( i_15_  &  n_n242  &  n_n222 ) ;
 assign wire19274 = ( n_n143 ) | ( n_n253  &  n_n281 ) ;
 assign wire19275 = ( n_n279  &  wire899 ) | ( n_n279  &  wire898 ) ;
 assign wire19278 = ( n_n207  &  wire1071 ) | ( n_n207  &  wire1181 ) ;
 assign wire19279 = ( n_n253  &  n_n278 ) | ( n_n279  &  wire902 ) ;
 assign wire19280 = ( n_n279  &  wire912 ) | ( wire197  &  wire962 ) ;
 assign wire19284 = ( i_11_  &  n_n163  &  n_n281 ) | ( (~ i_11_)  &  n_n163  &  n_n281 ) | ( i_11_  &  n_n163  &  n_n278 ) | ( (~ i_11_)  &  n_n163  &  n_n278 ) ;
 assign wire19285 = ( wire5999 ) | ( n_n279  &  wire901 ) | ( n_n279  &  wire897 ) ;
 assign wire19286 = ( n_n149 ) | ( n_n279  &  wire911 ) ;
 assign wire19287 = ( n_n279  &  wire900 ) | ( wire197  &  wire1225 ) ;
 assign wire19288 = ( wire5990 ) | ( n_n177  &  wire19286 ) | ( n_n177  &  wire19287 ) ;
 assign wire19290 = ( i_3_  &  i_5_ ) ;
 assign wire19291 = ( i_7_  &  i_6_  &  (~ i_4_) ) ;
 assign wire19292 = ( wire326 ) | ( wire19244 ) | ( wire911  &  n_n220 ) ;
 assign wire19294 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire19296 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire19297 = ( wire5985 ) | ( i_9_  &  i_10_  &  wire1265 ) | ( (~ i_9_)  &  (~ i_10_)  &  wire1265 ) ;
 assign wire19299 = ( i_7_  &  i_8_  &  (~ i_6_) ) | ( i_7_  &  (~ i_8_)  &  (~ i_6_)  &  wire1317 ) ;
 assign wire19300 = ( (~ i_7_)  &  (~ i_6_) ) | ( (~ i_7_)  &  i_8_  &  i_6_ ) | ( (~ i_7_)  &  (~ i_8_)  &  i_6_  &  wire315 ) ;
 assign wire19301 = ( i_5_  &  i_3_  &  (~ i_4_)  &  n_n165 ) ;
 assign wire19302 = ( wire5973 ) | ( wire19299  &  wire19301 ) | ( wire19300  &  wire19301 ) ;
 assign wire19303 = ( wire19297 ) | ( wire19302 ) | ( wire315  &  wire1264 ) ;
 assign wire19305 = ( n_n5017 ) | ( wire6008 ) | ( wire6009 ) | ( wire19278 ) ;
 assign wire19306 = ( n_n5007 ) | ( n_n5048 ) | ( wire19303 ) | ( wire19305 ) ;
 assign wire19307 = ( (~ i_9_)  &  (~ i_10_) ) | ( n_n279  &  wire912 ) ;
 assign wire19308 = ( wire328 ) | ( wire19237 ) | ( n_n220  &  wire912 ) ;
 assign wire19309 = ( wire397 ) | ( wire19307 ) | ( n_n281  &  wire914 ) ;
 assign wire19311 = ( n_n242  &  n_n222 ) | ( i_15_  &  n_n242  &  n_n279 ) ;
 assign wire19313 = ( wire196 ) | ( wire215 ) | ( n_n281  &  wire913 ) ;
 assign wire19314 = ( n_n150 ) | ( n_n179 ) | ( wire19253 ) | ( wire19311 ) ;
 assign wire19316 = ( n_n147 ) | ( n_n148 ) | ( wire19237 ) | ( wire19238 ) ;
 assign wire19318 = ( i_9_  &  i_10_ ) | ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) ;
 assign wire19319 = ( wire287 ) | ( wire911  &  n_n281 ) ;
 assign wire19320 = ( wire19318 ) | ( n_n242  &  wire152 ) ;
 assign wire19323 = ( wire5863 ) | ( n_n126  &  wire1400 ) ;
 assign wire19324 = ( wire397 ) | ( wire19307 ) | ( n_n281  &  wire914 ) ;
 assign wire19326 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  i_12_  &  (~ i_11_) ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19327 = ( wire352 ) | ( n_n281  &  wire913 ) | ( n_n281  &  wire914 ) ;
 assign wire19329 = ( n_n223 ) | ( n_n150 ) | ( wire214 ) | ( wire19311 ) ;
 assign wire19330 = ( n_n179 ) | ( wire19253 ) | ( wire19326 ) | ( wire19327 ) ;
 assign wire19331 = ( wire5862 ) | ( n_n128  &  wire398 ) | ( n_n128  &  wire19324 ) ;
 assign wire19332 = ( n_n222  &  n_n259 ) | ( i_15_  &  n_n279  &  n_n259 ) ;
 assign wire19334 = ( n_n222  &  n_n247 ) | ( i_15_  &  n_n279  &  n_n247 ) ;
 assign wire19337 = ( n_n204 ) | ( wire184 ) | ( wire130 ) | ( wire196 ) ;
 assign wire19339 = ( wire5848 ) | ( wire5850 ) | ( wire5854 ) | ( wire5855 ) ;
 assign wire19340 = ( n_n5030 ) | ( wire5849 ) | ( wire19323 ) ;
 assign wire19341 = ( wire5861 ) | ( wire19331 ) | ( wire19339 ) ;
 assign wire19342 = ( wire287 ) | ( wire901  &  n_n281 ) ;
 assign wire19344 = ( wire352 ) | ( n_n281  &  wire905 ) | ( n_n281  &  wire914 ) ;
 assign wire19345 = ( i_9_  &  i_10_ ) | ( i_9_  &  (~ i_10_)  &  i_11_ ) | ( i_9_  &  (~ i_10_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire19347 = ( wire215 ) | ( wire152  &  wire1501 ) ;
 assign wire19348 = ( wire19345 ) | ( wire911  &  n_n281 ) | ( n_n281  &  wire912 ) ;
 assign wire19350 = ( i_5_  &  (~ i_6_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire19353 = ( i_6_  &  n_n230 ) | ( i_7_  &  i_6_  &  n_n260 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260 ) | ( i_7_  &  (~ i_6_)  &  n_n230 ) ;
 assign wire19354 = ( (~ i_6_)  &  n_n264 ) | ( (~ i_7_)  &  i_6_  &  n_n264 ) | ( i_7_  &  i_6_  &  n_n284 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n284 ) ;
 assign wire19355 = ( wire5824 ) | ( n_n120  &  wire19353 ) | ( n_n120  &  wire19354 ) ;
 assign wire19356 = ( n_n5009 ) | ( wire19355 ) ;
 assign wire19359 = ( i_1_  &  i_2_ ) | ( i_2_  &  (~ i_0_) ) | ( i_3_  &  i_1_  &  (~ i_2_)  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire19363 = ( wire5812 ) | ( wire289  &  n_n118  &  n_n230 ) ;
 assign wire19364 = ( n_n5664 ) | ( n_n5679 ) | ( wire587 ) ;
 assign wire19365 = ( wire826 ) | ( n_n281  &  wire914  &  wire1474 ) ;
 assign wire19369 = ( n_n5686 ) | ( wire394 ) | ( n_n151  &  wire937 ) ;
 assign wire19373 = ( n_n4476 ) | ( wire893 ) | ( wire19363 ) | ( wire19364 ) ;
 assign wire19374 = ( n_n4477 ) | ( wire507 ) | ( wire5797 ) | ( wire19369 ) ;
 assign wire19377 = ( n_n54  &  n_n100 ) | ( n_n241  &  n_n103 ) ;
 assign wire19379 = ( wire386 ) | ( wire372 ) ;
 assign wire19380 = ( wire392 ) | ( wire19377 ) | ( n_n255  &  n_n31 ) ;
 assign wire19381 = ( n_n4  &  wire44 ) | ( n_n4  &  wire900  &  n_n220 ) ;
 assign wire19383 = ( n_n4  &  n_n95 ) | ( n_n4  &  n_n49 ) | ( n_n4  &  wire71 ) ;
 assign wire19384 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) ;
 assign wire19385 = ( (~ i_15_)  &  n_n279  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) ;
 assign wire19386 = ( n_n90 ) | ( wire19384 ) | ( n_n220  &  wire906 ) ;
 assign wire19387 = ( wire5775 ) | ( wire19383 ) | ( n_n268  &  n_n59 ) ;
 assign wire19391 = ( n_n4  &  wire1924 ) | ( n_n3  &  wire1940 ) ;
 assign wire19393 = ( wire557 ) | ( wire374 ) | ( wire5754 ) ;
 assign wire19394 = ( n_n281  &  wire903 ) | ( n_n228  &  wire902 ) ;
 assign wire19395 = ( wire50 ) | ( wire19394 ) | ( n_n228  &  wire897 ) ;
 assign wire19396 = ( wire5749 ) | ( n_n268  &  wire190 ) | ( n_n268  &  wire124 ) ;
 assign wire19398 = ( n_n3751 ) | ( wire5750 ) | ( wire5778 ) | ( wire19396 ) ;
 assign wire19400 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n252 ) ;
 assign wire19401 = ( n_n3  &  n_n14 ) | ( n_n3  &  n_n281  &  wire904 ) ;
 assign wire19402 = ( n_n281  &  wire903 ) | ( n_n228  &  wire902 ) ;
 assign wire19403 = ( wire50 ) | ( wire19402 ) | ( n_n228  &  wire897 ) ;
 assign wire19405 = ( wire349 ) | ( wire5743 ) | ( wire19400 ) | ( wire19401 ) ;
 assign wire19407 = ( (~ i_15_)  &  n_n275  &  n_n279 ) | ( i_15_  &  n_n275  &  n_n225 ) ;
 assign wire19408 = ( i_15_  &  n_n275  &  n_n281 ) | ( (~ i_15_)  &  n_n275  &  n_n225 ) ;
 assign wire19409 = ( n_n22 ) | ( wire19407 ) | ( n_n256  &  wire897 ) ;
 assign wire19410 = ( n_n171 ) | ( n_n73 ) | ( wire53 ) | ( wire19408 ) ;
 assign wire19413 = ( n_n3731 ) | ( n_n3736 ) | ( wire792 ) ;
 assign wire19417 = ( n_n29 ) | ( n_n26 ) | ( wire80 ) | ( wire88 ) ;
 assign wire19418 = ( n_n76 ) | ( wire49 ) | ( n_n101 ) | ( wire61 ) ;
 assign wire19420 = ( n_n3408 ) | ( wire5728 ) | ( n_n4  &  wire1555 ) ;
 assign wire19422 = ( n_n3634 ) | ( n_n3636 ) | ( wire19420 ) ;
 assign wire19424 = ( n_n171 ) | ( n_n24 ) | ( wire53 ) | ( wire19407 ) ;
 assign wire19426 = ( n_n3778 ) | ( n_n2  &  wire1871 ) ;
 assign wire19430 = ( wire5699 ) | ( n_n2  &  wire1899 ) ;
 assign wire19431 = ( n_n3757 ) | ( wire5700 ) | ( wire5709 ) | ( wire5710 ) ;
 assign wire19435 = ( n_n2597 ) | ( n_n2598 ) | ( n_n2599 ) | ( wire19430 ) ;
 assign wire19439 = ( n_n1  &  n_n49 ) | ( n_n1  &  wire71 ) | ( n_n1  &  wire1916 ) ;
 assign wire19440 = ( n_n3781 ) | ( n_n3786 ) | ( n_n2  &  wire1320 ) ;
 assign wire19442 = ( n_n3  &  wire99 ) | ( n_n3  &  n_n95 ) | ( n_n3  &  n_n49 ) ;
 assign wire19443 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n15 ) ;
 assign wire19445 = ( n_n3727 ) | ( wire409 ) | ( wire546 ) | ( wire19443 ) ;
 assign wire19446 = ( wire5681 ) | ( wire5682 ) | ( wire5683 ) | ( wire19442 ) ;
 assign wire19447 = ( n_n4  &  n_n228  &  wire902 ) | ( n_n53  &  n_n228  &  wire902 ) ;
 assign wire19452 = ( wire634 ) | ( n_n1  &  wire68 ) | ( n_n1  &  wire1877 ) ;
 assign wire19453 = ( n_n3791 ) | ( n_n2274 ) | ( n_n639 ) | ( wire19447 ) ;
 assign wire19455 = ( wire694 ) | ( wire544 ) | ( wire19452 ) | ( wire19453 ) ;
 assign wire19457 = ( i_15_  &  n_n275  &  n_n279 ) | ( (~ i_15_)  &  n_n275  &  n_n228 ) ;
 assign wire19458 = ( n_n31  &  n_n227 ) | ( n_n207  &  n_n103 ) ;
 assign wire19460 = ( n_n4  &  n_n93 ) | ( n_n94  &  n_n24 ) ;
 assign wire19461 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n30 ) | ( n_n4  &  n_n26 ) ;
 assign wire19465 = ( wire455 ) | ( wire374 ) | ( wire19461 ) ;
 assign wire19466 = ( wire799 ) | ( wire471 ) | ( wire19460 ) ;
 assign wire19467 = ( wire747 ) | ( wire5660 ) | ( wire5661 ) ;
 assign wire19469 = ( wire900  &  n_n228 ) | ( n_n281  &  wire904 ) ;
 assign wire19470 = ( n_n5  &  n_n66 ) | ( n_n5  &  n_n14 ) | ( n_n5  &  wire70 ) ;
 assign wire19472 = ( wire19470 ) | ( wire5651 ) ;
 assign wire19473 = ( n_n3806 ) | ( wire5650 ) | ( wire5656 ) | ( wire5657 ) ;
 assign wire19475 = ( n_n9  &  n_n227 ) | ( n_n9  &  n_n207 ) | ( n_n227  &  n_n59 ) | ( n_n207  &  n_n59 ) ;
 assign wire19478 = ( n_n3803 ) | ( wire5640 ) | ( wire5642 ) ;
 assign wire19480 = ( n_n3686 ) | ( wire5643 ) | ( wire19475 ) | ( wire19478 ) ;
 assign wire19485 = ( wire153  &  n_n6 ) | ( n_n6  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign wire19489 = ( n_n3827 ) | ( wire771 ) | ( n_n3579 ) ;
 assign wire19490 = ( wire770 ) | ( wire5617 ) | ( wire5625 ) | ( wire5626 ) ;
 assign wire19491 = ( n_n281  &  wire903 ) | ( n_n228  &  wire902 ) ;
 assign wire19493 = ( n_n60 ) | ( wire50 ) | ( n_n59 ) | ( wire63 ) ;
 assign wire19495 = ( n_n3791 ) | ( wire5606 ) | ( n_n53  &  n_n9 ) ;
 assign wire19497 = ( wire56 ) | ( wire19407 ) | ( n_n256  &  wire897 ) ;
 assign wire19498 = ( n_n171 ) | ( n_n73 ) | ( wire53 ) | ( wire19408 ) ;
 assign wire19499 = ( n_n53  &  n_n220  &  wire908 ) | ( n_n53  &  n_n256  &  wire908 ) ;
 assign wire19502 = ( wire478 ) | ( wire19499 ) | ( n_n53  &  wire1948 ) ;
 assign wire19504 = ( n_n1542 ) | ( wire5595 ) | ( wire5596 ) | ( wire19502 ) ;
 assign wire19506 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire19507 = ( n_n93 ) | ( wire76 ) | ( n_n220  &  wire906 ) ;
 assign wire19508 = ( n_n44 ) | ( n_n90 ) | ( wire19384 ) | ( wire19385 ) ;
 assign wire19511 = ( wire662 ) | ( n_n48  &  wire1917 ) ;
 assign wire19512 = ( wire5565 ) | ( wire5564 ) ;
 assign wire19515 = ( wire5591 ) | ( wire5592 ) | ( n_n57  &  n_n9 ) ;
 assign wire19516 = ( wire571 ) | ( wire737 ) | ( n_n53  &  wire68 ) ;
 assign wire19519 = ( wire5589 ) | ( wire19516 ) | ( n_n57  &  n_n12 ) ;
 assign wire19520 = ( n_n4381 ) | ( n_n3850 ) | ( wire5577 ) | ( wire19515 ) ;
 assign wire19522 = ( wire741 ) | ( wire869 ) | ( n_n53  &  wire1852 ) ;
 assign wire19523 = ( wire473 ) | ( wire19519 ) | ( wire19520 ) | ( wire19522 ) ;
 assign wire19526 = ( n_n5  &  wire255 ) | ( n_n5  &  wire190 ) ;
 assign wire19528 = ( n_n4770 ) | ( wire19526 ) | ( n_n6  &  wire1747 ) ;
 assign wire19530 = ( n_n3390 ) | ( wire5636 ) | ( wire5637 ) | ( wire19528 ) ;
 assign wire19534 = ( n_n4675 ) | ( n_n4676 ) | ( n_n57  &  wire1878 ) ;
 assign wire19535 = ( wire56 ) | ( wire19407 ) | ( n_n256  &  wire897 ) ;
 assign wire19536 = ( n_n171 ) | ( n_n24 ) | ( wire53 ) | ( wire19407 ) ;
 assign wire19537 = ( n_n57  &  n_n22 ) | ( n_n56  &  wire49 ) ;
 assign wire19539 = ( n_n56  &  n_n76 ) | ( n_n57  &  wire70 ) ;
 assign wire19540 = ( wire460 ) | ( wire19539 ) ;
 assign wire19541 = ( n_n4924 ) | ( wire788 ) | ( wire5544 ) ;
 assign wire19544 = ( n_n3709 ) | ( n_n4680 ) | ( n_n4677 ) | ( wire19534 ) ;
 assign wire19546 = ( n_n3710 ) | ( n_n3708 ) | ( wire19540 ) | ( wire19541 ) ;
 assign wire19548 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) ;
 assign wire19549 = ( n_n94  &  n_n75 ) | ( n_n100  &  n_n103 ) ;
 assign wire19550 = ( n_n94  &  n_n24 ) | ( n_n94  &  n_n74 ) | ( n_n94  &  wire77 ) ;
 assign wire19553 = ( wire471 ) | ( wire19549 ) | ( wire19550 ) ;
 assign wire19554 = ( n_n1641 ) | ( wire5516 ) | ( wire5517 ) ;
 assign wire19556 = ( wire898  &  n_n228 ) | ( n_n281  &  wire906 ) ;
 assign wire19558 = ( wire44 ) | ( n_n9 ) | ( n_n252 ) | ( wire63 ) ;
 assign wire19559 = ( n_n100  &  n_n60 ) | ( n_n100  &  n_n9 ) | ( n_n100  &  wire63 ) ;
 assign wire19560 = ( wire19559 ) | ( wire5509 ) ;
 assign wire19565 = ( n_n4681 ) | ( n_n4686 ) | ( n_n56  &  wire1892 ) ;
 assign wire19566 = ( wire863 ) | ( n_n4687 ) | ( wire5494 ) | ( wire5506 ) ;
 assign wire19567 = ( wire69 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire19568 = ( wire40  &  n_n100 ) | ( n_n100  &  wire898  &  n_n228 ) ;
 assign wire19571 = ( n_n100  &  wire91 ) | ( n_n100  &  wire121 ) | ( n_n100  &  wire1903 ) ;
 assign wire19573 = ( wire459 ) | ( wire5485 ) | ( wire19568 ) | ( wire19571 ) ;
 assign wire19575 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire19576 = ( n_n97 ) | ( n_n51 ) | ( wire71 ) | ( wire19575 ) ;
 assign wire19577 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire19578 = ( (~ i_15_)  &  n_n279  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) ;
 assign wire19579 = ( wire51 ) | ( wire71 ) | ( wire898  &  n_n256 ) ;
 assign wire19581 = ( n_n3884 ) | ( n_n94  &  wire1943 ) ;
 assign wire19582 = ( n_n3881 ) | ( n_n105  &  n_n100 ) | ( n_n100  &  wire1368 ) ;
 assign wire19586 = ( n_n3722 ) | ( wire776 ) | ( wire821 ) | ( wire5472 ) ;
 assign wire19588 = ( n_n863 ) | ( n_n3661 ) | ( n_n3404 ) | ( wire19586 ) ;
 assign wire19592 = ( n_n3625 ) | ( n_n3626 ) | ( n_n3624 ) | ( wire19422 ) ;
 assign wire19593 = ( n_n3627 ) | ( n_n3631 ) | ( n_n3632 ) | ( wire19588 ) ;
 assign wire19598 = ( wire535 ) | ( wire289  &  n_n118  &  n_n264 ) ;
 assign wire19599 = ( wire364 ) | ( wire777 ) | ( wire834 ) ;
 assign wire19601 = ( wire19598 ) | ( wire19599 ) | ( n_n123  &  wire939 ) ;
 assign wire19602 = ( n_n124  &  wire938 ) | ( n_n124  &  wire1952 ) ;
 assign wire19604 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire913 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire913 ) ;
 assign wire19605 = ( (~ i_9_)  &  (~ i_10_) ) | ( wire911  &  n_n281 ) ;
 assign wire19608 = ( n_n107 ) | ( n_n135 ) | ( wire250 ) | ( wire19604 ) ;
 assign wire19609 = ( wire364 ) | ( n_n5769 ) | ( n_n124  &  wire48 ) ;
 assign wire19610 = ( wire19609 ) | ( n_n124  &  n_n110 ) | ( n_n124  &  wire54 ) ;
 assign wire19613 = ( n_n118  &  n_n264  &  n_n155 ) | ( n_n118  &  n_n155  &  n_n284 ) ;
 assign wire19614 = ( i_7_  &  i_6_  &  n_n118  &  n_n284 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n284 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n284 ) ;
 assign wire19617 = ( n_n5678 ) | ( n_n5671 ) | ( wire396  &  wire940 ) ;
 assign wire19619 = ( wire5453 ) | ( wire19613 ) | ( wire19614 ) | ( wire19617 ) ;
 assign wire19620 = ( wire582 ) | ( wire5445 ) | ( n_n106  &  wire941 ) ;
 assign wire19622 = ( wire5457 ) | ( wire19610 ) | ( wire19619 ) | ( wire19620 ) ;
 assign wire19624 = ( n_n5693 ) | ( n_n130  &  n_n220  &  wire914 ) ;
 assign wire19625 = ( n_n5797 ) | ( wire5441 ) | ( wire5442 ) ;
 assign wire19626 = ( wire5439 ) | ( n_n128  &  n_n111 ) | ( n_n128  &  wire54 ) ;
 assign wire19628 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire19631 = ( wire19628 ) | ( wire793 ) ;
 assign wire19632 = ( n_n5792 ) | ( n_n5794 ) | ( wire880 ) | ( n_n5672 ) ;
 assign wire19633 = ( n_n139  &  n_n111 ) | ( n_n132  &  wire54 ) ;
 assign wire19636 = ( n_n121  &  n_n111 ) | ( n_n132  &  n_n111 ) | ( n_n111  &  n_n122 ) ;
 assign wire19638 = ( n_n5797 ) | ( n_n139  &  wire54 ) ;
 assign wire19642 = ( n_n5671 ) | ( wire5412 ) | ( wire5413 ) ;
 assign wire19644 = ( wire5411 ) | ( wire19631 ) | ( wire19632 ) | ( wire19642 ) ;
 assign wire19645 = ( wire5426 ) | ( wire5430 ) | ( wire19633 ) | ( wire19636 ) ;
 assign wire19648 = ( n_n4442 ) | ( n_n4439 ) | ( wire19644 ) | ( wire19645 ) ;
 assign wire19654 = ( wire5390 ) | ( wire5400 ) | ( n_n5  &  wire1874 ) ;
 assign wire19655 = ( n_n4815 ) | ( n_n4821 ) | ( n_n4814 ) | ( n_n4816 ) ;
 assign wire19657 = ( n_n29 ) | ( n_n26 ) | ( wire80 ) | ( wire88 ) ;
 assign wire19659 = ( n_n6  &  wire1016 ) | ( n_n6  &  wire1920 ) ;
 assign wire19661 = ( wire807 ) | ( n_n279  &  wire904 ) | ( n_n220  &  wire904 ) ;
 assign wire19663 = ( n_n179 ) | ( n_n39 ) | ( wire57 ) | ( wire245 ) ;
 assign wire19665 = ( n_n6582 ) | ( n_n4870 ) | ( n_n5  &  wire1894 ) ;
 assign wire19668 = ( wire911  &  n_n228 ) | ( n_n281  &  wire905 ) ;
 assign wire19669 = ( n_n6  &  n_n220  &  wire904 ) | ( n_n6  &  n_n256  &  wire904 ) ;
 assign wire19671 = ( wire5362 ) | ( wire19669 ) | ( n_n5  &  wire81 ) ;
 assign wire19674 = ( n_n93 ) | ( n_n90 ) | ( wire76 ) | ( wire19384 ) ;
 assign wire19675 = ( wire68 ) | ( wire96 ) | ( n_n222  &  wire904 ) ;
 assign wire19677 = ( wire5357 ) | ( wire5371 ) | ( wire5372 ) | ( wire19665 ) ;
 assign wire19682 = ( wire184 ) | ( wire70 ) | ( wire898  &  n_n220 ) ;
 assign wire19683 = ( wire901  &  n_n228 ) | ( n_n281  &  wire904 ) ;
 assign wire19685 = ( wire113 ) | ( wire281 ) | ( n_n258  &  wire907 ) ;
 assign wire19687 = ( wire60 ) | ( n_n204 ) | ( n_n112 ) | ( wire52 ) ;
 assign wire19691 = ( wire247 ) | ( wire123 ) | ( wire227 ) ;
 assign wire19692 = ( n_n57  &  wire247 ) | ( n_n57  &  wire210 ) | ( n_n57  &  wire19687 ) ;
 assign wire19693 = ( n_n62 ) | ( wire101 ) | ( n_n281  &  wire907 ) ;
 assign wire19696 = ( n_n3324 ) | ( n_n4381 ) | ( wire5587 ) | ( wire5588 ) ;
 assign wire19698 = ( n_n3850 ) | ( wire5327 ) | ( wire5328 ) | ( wire19696 ) ;
 assign wire19701 = ( wire268  &  n_n57 ) | ( n_n57  &  wire198 ) ;
 assign wire19703 = ( n_n4941 ) | ( n_n4942 ) | ( wire762 ) ;
 assign wire19704 = ( wire728 ) | ( wire19701 ) | ( n_n57  &  wire167 ) ;
 assign wire19705 = ( n_n56  &  wire190 ) | ( n_n57  &  wire124 ) ;
 assign wire19706 = ( n_n56  &  wire124 ) | ( n_n57  &  wire212 ) ;
 assign wire19707 = ( n_n56  &  wire212 ) | ( n_n57  &  wire119 ) ;
 assign wire19709 = ( wire19706 ) | ( wire19705 ) ;
 assign wire19710 = ( wire761 ) | ( wire19707 ) | ( n_n56  &  wire198 ) ;
 assign wire19711 = ( wire60 ) | ( wire140 ) | ( n_n279  &  wire911 ) ;
 assign wire19712 = ( wire167 ) | ( wire52 ) | ( n_n279  &  wire913 ) ;
 assign wire19713 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire19714 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire19717 = ( wire706 ) | ( wire481 ) | ( wire5298 ) | ( wire5299 ) ;
 assign wire19718 = ( wire19703 ) | ( wire19704 ) | ( wire19709 ) | ( wire19710 ) ;
 assign wire19720 = ( n_n56  &  wire254 ) | ( n_n57  &  wire180 ) ;
 assign wire19723 = ( wire19720 ) | ( n_n57  &  wire153 ) | ( n_n57  &  wire166 ) ;
 assign wire19724 = ( n_n4954 ) | ( n_n4953 ) | ( n_n4955 ) | ( wire671 ) ;
 assign wire19725 = ( n_n57  &  wire200 ) | ( n_n56  &  wire277 ) ;
 assign wire19727 = ( wire704 ) | ( n_n57  &  wire157 ) | ( n_n57  &  wire273 ) ;
 assign wire19728 = ( wire729 ) | ( wire19725 ) | ( wire268  &  n_n56 ) ;
 assign wire19730 = ( n_n56  &  wire224 ) | ( n_n56  &  wire180 ) ;
 assign wire19732 = ( n_n4970 ) | ( wire614 ) | ( n_n56  &  wire166 ) ;
 assign wire19733 = ( n_n4967 ) | ( wire613 ) | ( wire19730 ) ;
 assign wire19735 = ( wire19723 ) | ( wire19724 ) | ( wire19727 ) | ( wire19728 ) ;
 assign wire19736 = ( wire19732 ) | ( wire19733 ) | ( wire19735 ) ;
 assign wire19738 = ( i_15_  &  n_n242  &  n_n281 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) ;
 assign wire19741 = ( wire5262 ) | ( n_n5  &  wire976 ) ;
 assign wire19742 = ( n_n4826 ) | ( n_n4828 ) | ( n_n4823 ) | ( wire584 ) ;
 assign wire19744 = ( n_n112 ) | ( n_n67 ) | ( wire84 ) | ( wire19738 ) ;
 assign wire19747 = ( n_n4834 ) | ( n_n4839 ) | ( n_n6  &  wire1893 ) ;
 assign wire19749 = ( wire699 ) | ( n_n4838 ) | ( wire5248 ) | ( wire19747 ) ;
 assign wire19752 = ( n_n6  &  wire1937 ) | ( n_n5  &  wire1945 ) ;
 assign wire19753 = ( n_n4858 ) | ( n_n4864 ) | ( n_n5  &  wire1884 ) ;
 assign wire19754 = ( n_n4852 ) | ( wire5228 ) | ( wire5244 ) | ( wire5245 ) ;
 assign wire19755 = ( wire5238 ) | ( wire5239 ) | ( wire5242 ) | ( wire5243 ) ;
 assign wire19757 = ( wire19754 ) | ( wire19753 ) ;
 assign wire19758 = ( wire5240 ) | ( wire5241 ) | ( wire19752 ) | ( wire19755 ) ;
 assign wire19759 = ( n_n4807 ) | ( n_n4806 ) | ( n_n5  &  wire72 ) ;
 assign wire19761 = ( n_n4223 ) | ( n_n4224 ) | ( wire19759 ) ;
 assign wire19763 = ( n_n4204 ) | ( wire19749 ) | ( wire19761 ) ;
 assign wire19764 = ( n_n4203 ) | ( n_n4206 ) | ( wire19757 ) | ( wire19758 ) ;
 assign wire19766 = ( n_n4306 ) | ( wire19763 ) | ( wire19764 ) ;
 assign wire19768 = ( n_n3255 ) | ( n_n2  &  wire1899 ) ;
 assign wire19770 = ( wire395 ) | ( wire5215 ) | ( n_n2  &  n_n111 ) ;
 assign wire19772 = ( n_n81 ) | ( n_n35 ) | ( wire64 ) | ( wire86 ) ;
 assign wire19773 = ( wire55 ) | ( wire64 ) | ( n_n279  &  wire907 ) ;
 assign wire19774 = ( n_n179 ) | ( n_n81 ) | ( wire57 ) | ( wire86 ) ;
 assign wire19776 = ( n_n3257 ) | ( n_n1412 ) | ( n_n1  &  n_n32 ) ;
 assign wire19778 = ( n_n2603 ) | ( wire5208 ) | ( wire19776 ) ;
 assign wire19780 = ( n_n106  &  n_n2 ) | ( n_n2  &  n_n62 ) | ( n_n2  &  wire101 ) ;
 assign wire19783 = ( n_n3523 ) | ( n_n2  &  wire1932 ) ;
 assign wire19784 = ( n_n3525 ) | ( n_n3519 ) | ( n_n3520 ) | ( n_n3524 ) ;
 assign wire19787 = ( n_n2633 ) | ( n_n2  &  wire90 ) | ( n_n2  &  wire1951 ) ;
 assign wire19790 = ( n_n9 ) | ( n_n65 ) | ( wire73 ) | ( wire63 ) ;
 assign wire19791 = ( wire5184 ) | ( wire5709 ) | ( n_n1  &  n_n12 ) ;
 assign wire19793 = ( wire5185 ) | ( wire5205 ) | ( wire19780 ) | ( wire19791 ) ;
 assign wire19797 = ( wire723 ) | ( n_n1  &  wire1916 ) ;
 assign wire19798 = ( n_n3781 ) | ( n_n3778 ) | ( n_n2  &  wire1819 ) ;
 assign wire19801 = ( wire89 ) | ( n_n83 ) | ( n_n49 ) | ( wire71 ) ;
 assign wire19802 = ( n_n1  &  n_n111 ) | ( n_n1  &  n_n38 ) | ( n_n1  &  wire453 ) ;
 assign wire19803 = ( n_n3260 ) | ( n_n2  &  wire1871 ) ;
 assign wire19807 = ( n_n106  &  n_n2 ) | ( n_n1  &  wire68 ) ;
 assign wire19808 = ( wire19807 ) | ( n_n2  &  wire200 ) | ( n_n2  &  wire112 ) ;
 assign wire19810 = ( n_n3162 ) | ( wire19808 ) | ( n_n2  &  wire1627 ) ;
 assign wire19812 = ( n_n2583 ) | ( n_n2582 ) | ( wire19810 ) ;
 assign wire19814 = ( n_n228  &  wire897 ) | ( n_n281  &  wire908 ) ;
 assign wire19817 = ( wire75 ) | ( wire72 ) | ( n_n281  &  wire913 ) ;
 assign wire19818 = ( n_n9 ) | ( n_n206 ) | ( wire118 ) | ( wire63 ) ;
 assign wire19819 = ( n_n2618 ) | ( n_n1  &  wire944 ) ;
 assign wire19821 = ( wire5153 ) | ( wire5160 ) | ( wire5161 ) | ( wire19819 ) ;
 assign wire19822 = ( n_n2573 ) | ( n_n2572 ) | ( wire19812 ) | ( wire19821 ) ;
 assign wire19825 = ( wire758 ) | ( n_n122  &  n_n220  &  wire914 ) ;
 assign wire19826 = ( n_n5678 ) | ( n_n5671 ) | ( wire5144 ) ;
 assign wire19829 = ( wire583 ) | ( wire5441 ) | ( wire5442 ) | ( wire19825 ) ;
 assign wire19830 = ( wire582 ) | ( wire19826 ) | ( n_n121  &  wire1359 ) ;
 assign wire19831 = ( wire54 ) | ( wire266 ) | ( wire913  &  n_n220 ) ;
 assign wire19833 = ( wire54 ) | ( wire103 ) | ( wire913  &  n_n220 ) ;
 assign wire19834 = ( wire364 ) | ( n_n124  &  wire1952 ) ;
 assign wire19835 = ( wire5138 ) | ( n_n127  &  wire294 ) | ( n_n127  &  wire19831 ) ;
 assign wire19837 = ( n_n5769 ) | ( n_n127  &  wire48 ) ;
 assign wire19838 = ( wire19829 ) | ( wire19830 ) | ( wire19837 ) ;
 assign wire19842 = ( n_n207  &  n_n257 ) | ( n_n207  &  n_n228  &  wire902 ) ;
 assign wire19843 = ( n_n9  &  n_n227 ) | ( n_n227  &  n_n59 ) | ( n_n207  &  n_n59 ) ;
 assign wire19846 = ( n_n3550 ) | ( wire19842 ) | ( n_n207  &  wire1813 ) ;
 assign wire19847 = ( wire887 ) | ( wire19843 ) | ( n_n227  &  wire1814 ) ;
 assign wire19848 = ( wire913  &  n_n258 ) | ( n_n228  &  wire897 ) ;
 assign wire19849 = ( n_n265  &  n_n62 ) | ( n_n268  &  n_n148 ) ;
 assign wire19852 = ( wire60 ) | ( n_n204 ) | ( n_n112 ) | ( wire52 ) ;
 assign wire19853 = ( wire190 ) | ( wire119 ) | ( wire210 ) ;
 assign wire19854 = ( n_n265  &  wire277 ) | ( n_n268  &  wire247 ) ;
 assign wire19855 = ( wire19854 ) | ( n_n268  &  wire124 ) | ( n_n268  &  wire212 ) ;
 assign wire19856 = ( wire50 ) | ( wire157 ) | ( n_n281  &  wire903 ) ;
 assign wire19857 = ( n_n265  &  wire268 ) | ( n_n265  &  wire200 ) | ( n_n265  &  wire112 ) ;
 assign wire19859 = ( wire19857 ) | ( n_n268  &  wire400 ) | ( n_n268  &  wire19856 ) ;
 assign wire19860 = ( n_n2550 ) | ( n_n2545 ) | ( wire19859 ) ;
 assign wire19862 = ( n_n5796 ) | ( n_n6  &  n_n256  &  wire914 ) ;
 assign wire19864 = ( n_n5  &  n_n81 ) | ( n_n5  &  wire86 ) | ( n_n5  &  wire1894 ) ;
 assign wire19865 = ( n_n4864 ) | ( n_n4870 ) | ( wire5099 ) | ( wire19862 ) ;
 assign wire19867 = ( wire153  &  n_n6 ) | ( n_n6  &  n_n113 ) | ( n_n6  &  wire57 ) ;
 assign wire19868 = ( wire617 ) | ( wire5091 ) | ( n_n5  &  wire255 ) ;
 assign wire19869 = ( n_n4770 ) | ( wire19867 ) ;
 assign wire19871 = ( wire632 ) | ( wire5611 ) | ( wire5613 ) | ( wire19868 ) ;
 assign wire19872 = ( wire674 ) | ( n_n4773 ) | ( wire5629 ) | ( wire19869 ) ;
 assign wire19874 = ( n_n70 ) | ( wire79 ) | ( n_n62 ) | ( wire101 ) ;
 assign wire19878 = ( n_n4826 ) | ( n_n4823 ) | ( wire584 ) | ( n_n4821 ) ;
 assign wire19881 = ( n_n6  &  n_n67 ) | ( n_n6  &  wire1893 ) | ( n_n6  &  wire19738 ) ;
 assign wire19882 = ( n_n4834 ) | ( n_n5  &  wire125 ) | ( n_n5  &  wire1229 ) ;
 assign wire19887 = ( wire5060 ) | ( wire5400 ) | ( n_n5  &  wire1874 ) ;
 assign wire19888 = ( n_n4815 ) | ( n_n4814 ) | ( n_n4816 ) | ( wire541 ) ;
 assign wire19890 = ( wire585 ) | ( wire5059 ) | ( wire19887 ) | ( wire19888 ) ;
 assign wire19892 = ( n_n29 ) | ( n_n26 ) | ( wire80 ) | ( wire88 ) ;
 assign wire19893 = ( n_n204 ) | ( n_n101 ) | ( wire52 ) | ( wire61 ) ;
 assign wire19896 = ( n_n4839 ) | ( n_n4842 ) | ( wire5054 ) ;
 assign wire19899 = ( wire5048 ) | ( n_n6  &  wire1937 ) ;
 assign wire19900 = ( n_n4858 ) | ( wire5047 ) | ( n_n5  &  wire1945 ) ;
 assign wire19903 = ( n_n6  &  n_n171 ) | ( n_n6  &  wire53 ) | ( n_n6  &  wire1920 ) ;
 assign wire19904 = ( n_n4846 ) | ( n_n4852 ) | ( wire5242 ) | ( wire5243 ) ;
 assign wire19906 = ( wire5240 ) | ( wire5241 ) | ( wire19903 ) | ( wire19904 ) ;
 assign wire19909 = ( n_n4287 ) | ( n_n4892 ) | ( wire5023 ) ;
 assign wire19914 = ( n_n4907 ) | ( n_n56  &  wire111 ) | ( n_n56  &  wire1898 ) ;
 assign wire19916 = ( n_n57  &  n_n11 ) | ( n_n56  &  n_n11 ) | ( n_n57  &  wire113 ) ;
 assign wire19918 = ( wire5013 ) | ( wire5014 ) | ( wire5589 ) | ( wire5590 ) ;
 assign wire19919 = ( n_n4895 ) | ( wire5002 ) | ( wire19916 ) ;
 assign wire19921 = ( wire5011 ) | ( wire5012 ) | ( wire19918 ) | ( wire19919 ) ;
 assign wire19925 = ( wire268  &  n_n56 ) | ( n_n56  &  wire157 ) | ( n_n56  &  wire273 ) ;
 assign wire19926 = ( n_n4941 ) | ( n_n4942 ) | ( wire729 ) ;
 assign wire19927 = ( wire19925 ) | ( wire268  &  n_n57 ) | ( n_n57  &  wire200 ) ;
 assign wire19928 = ( n_n56  &  wire124 ) | ( n_n56  &  wire212 ) ;
 assign wire19930 = ( wire761 ) | ( n_n57  &  wire165 ) | ( n_n57  &  wire140 ) ;
 assign wire19931 = ( wire760 ) | ( wire19928 ) | ( n_n57  &  wire198 ) ;
 assign wire19935 = ( n_n4914 ) | ( n_n56  &  wire1585 ) ;
 assign wire19936 = ( n_n4920 ) | ( n_n4921 ) | ( n_n4916 ) | ( wire705 ) ;
 assign wire19938 = ( n_n5796 ) | ( n_n56  &  wire49 ) ;
 assign wire19941 = ( n_n57  &  wire124 ) | ( n_n57  &  wire212 ) ;
 assign wire19943 = ( n_n4926 ) | ( n_n4923 ) | ( wire19938 ) ;
 assign wire19944 = ( n_n4924 ) | ( n_n4922 ) | ( wire19941 ) ;
 assign wire19946 = ( wire763 ) | ( wire4974 ) | ( wire19943 ) | ( wire19944 ) ;
 assign wire19948 = ( wire48 ) | ( n_n110 ) | ( n_n108 ) | ( wire103 ) ;
 assign wire19949 = ( n_n5796 ) | ( n_n272  &  n_n260  &  n_n165 ) ;
 assign wire19952 = ( n_n57  &  wire99 ) | ( n_n57  &  wire41 ) ;
 assign wire19953 = ( n_n4970 ) | ( n_n4966 ) | ( n_n4967 ) | ( wire19949 ) ;
 assign wire19954 = ( wire19952 ) | ( n_n152  &  wire299 ) | ( n_n152  &  wire19948 ) ;
 assign wire19955 = ( wire54 ) | ( wire913  &  n_n220 ) | ( n_n220  &  wire905 ) ;
 assign wire19956 = ( wire48 ) | ( n_n220  &  wire905 ) ;
 assign wire19957 = ( wire54 ) | ( wire103 ) | ( wire913  &  n_n220 ) ;
 assign wire19958 = ( wire394 ) | ( n_n139  &  wire48 ) | ( wire48  &  n_n132 ) ;
 assign wire19959 = ( wire19958 ) | ( wire1723  &  wire294 ) | ( wire1723  &  wire19955 ) ;
 assign wire19961 = ( wire452 ) | ( n_n5796 ) ;
 assign wire19963 = ( wire5812 ) | ( wire5813 ) | ( wire19364 ) | ( wire19961 ) ;
 assign wire19965 = ( n_n5686 ) | ( n_n5693 ) | ( wire609 ) | ( wire4947 ) ;
 assign wire19967 = ( wire507 ) | ( n_n4489 ) | ( wire19963 ) | ( wire19965 ) ;
 assign wire19969 = ( n_n57  &  wire153 ) | ( n_n57  &  wire166 ) ;
 assign wire19971 = ( n_n56  &  wire254 ) | ( n_n57  &  wire180 ) ;
 assign wire19973 = ( wire19969 ) | ( n_n56  &  wire166 ) | ( n_n56  &  wire180 ) ;
 assign wire19974 = ( wire4939 ) | ( wire19971 ) | ( n_n57  &  wire224 ) ;
 assign wire19977 = ( n_n56  &  wire200 ) | ( n_n56  &  wire99 ) | ( n_n56  &  wire112 ) ;
 assign wire19978 = ( n_n4954 ) | ( n_n4953 ) | ( wire672 ) ;
 assign wire19980 = ( n_n4955 ) | ( n_n4950 ) | ( wire19977 ) | ( wire19978 ) ;
 assign wire19981 = ( wire19926 ) | ( wire19927 ) | ( wire19973 ) | ( wire19974 ) ;
 assign wire19984 = ( n_n5796 ) | ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) ;
 assign wire19986 = ( n_n4806 ) | ( wire19984 ) | ( n_n5  &  wire72 ) ;
 assign wire19987 = ( n_n4808 ) | ( n_n4809 ) | ( wire19986 ) ;
 assign wire19988 = ( n_n4733 ) | ( wire19871 ) | ( wire19872 ) | ( wire19987 ) ;
 assign wire19989 = ( n_n4719 ) | ( n_n4730 ) | ( n_n4732 ) | ( wire19906 ) ;
 assign wire19990 = ( n_n4736 ) | ( n_n3397 ) | ( wire19921 ) | ( wire19988 ) ;
 assign wire19996 = ( i_3_  &  n_n116 ) | ( n_n155  &  n_n230  &  n_n116 ) ;
 assign wire19997 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire19998 = ( wire19997 ) | ( wire19996 ) ;
 assign wire19999 = ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire20000 = ( i_3_  &  n_n118 ) | ( n_n118  &  n_n260  &  n_n155 ) ;
 assign wire20001 = ( wire20000 ) | ( wire535 ) ;
 assign wire20002 = ( wire777 ) | ( n_n5675 ) | ( wire4928 ) | ( wire19999 ) ;
 assign wire20004 = ( n_n2772 ) | ( wire879 ) | ( wire19996 ) | ( wire19997 ) ;
 assign wire20007 = ( n_n127  &  n_n111 ) | ( n_n127  &  n_n108 ) | ( n_n108  &  n_n122 ) ;
 assign wire20008 = ( n_n127  &  n_n110 ) | ( n_n139  &  wire1703 ) ;
 assign wire20011 = ( n_n130  &  wire948 ) | ( n_n130  &  n_n111 ) | ( n_n121  &  n_n111 ) ;
 assign wire20012 = ( wire4905 ) | ( wire20011 ) | ( n_n110  &  n_n121 ) ;
 assign wire20015 = ( n_n139  &  n_n110 ) | ( wire48  &  n_n132 ) ;
 assign wire20016 = ( wire4900 ) | ( n_n139  &  wire48 ) ;
 assign wire20017 = ( wire48  &  n_n130 ) | ( n_n110  &  n_n132 ) ;
 assign wire20020 = ( wire4892 ) | ( n_n130  &  wire913  &  n_n220 ) ;
 assign wire20021 = ( n_n5693 ) | ( wire452 ) | ( wire758 ) | ( wire4890 ) ;
 assign wire20023 = ( n_n118  &  n_n264  &  n_n155 ) | ( n_n118  &  n_n155  &  n_n284 ) ;
 assign wire20027 = ( n_n5659 ) | ( n_n5673 ) | ( n_n5664 ) | ( wire587 ) ;
 assign wire20028 = ( n_n264  &  n_n155  &  n_n116 ) | ( n_n260  &  n_n155  &  n_n116 ) ;
 assign wire20030 = ( wire794 ) | ( wire581 ) ;
 assign wire20031 = ( n_n5685 ) | ( wire4871 ) | ( wire20028 ) ;
 assign wire20033 = ( wire4902 ) | ( wire20015 ) | ( wire20030 ) | ( wire20031 ) ;
 assign wire20034 = ( wire4896 ) | ( wire4899 ) | ( wire20016 ) | ( wire20017 ) ;
 assign wire20038 = ( n_n10  &  n_n100 ) | ( n_n100  &  n_n63 ) | ( n_n100  &  n_n62 ) ;
 assign wire20041 = ( n_n2702 ) | ( wire654 ) | ( n_n100  &  wire1149 ) ;
 assign wire20042 = ( wire4856 ) | ( wire4869 ) | ( wire4870 ) | ( wire20038 ) ;
 assign wire20045 = ( n_n133  &  n_n94 ) | ( n_n94  &  n_n17 ) | ( n_n94  &  n_n68 ) ;
 assign wire20047 = ( n_n2732 ) | ( n_n2398 ) | ( wire20045 ) ;
 assign wire20048 = ( wire4849 ) | ( n_n100  &  wire1150 ) ;
 assign wire20051 = ( wire113 ) | ( wire281 ) | ( n_n258  &  wire907 ) ;
 assign wire20052 = ( n_n2724 ) | ( n_n100  &  wire1152 ) ;
 assign wire20054 = ( wire4839 ) | ( wire4844 ) | ( wire4845 ) | ( wire20052 ) ;
 assign wire20055 = ( wire20041 ) | ( wire20042 ) | ( wire20047 ) | ( wire20048 ) ;
 assign wire20056 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire912 ) ;
 assign wire20060 = ( wire686 ) | ( wire391 ) | ( wire548 ) | ( wire774 ) ;
 assign wire20061 = ( wire773 ) | ( n_n100  &  wire198 ) | ( n_n100  &  wire167 ) ;
 assign wire20066 = ( n_n94  &  n_n204 ) | ( n_n94  &  n_n216 ) | ( n_n94  &  n_n203 ) ;
 assign wire20068 = ( wire20066 ) | ( n_n94  &  wire140 ) | ( n_n94  &  wire1661 ) ;
 assign wire20070 = ( n_n94  &  n_n75 ) | ( n_n94  &  n_n24 ) | ( n_n94  &  n_n74 ) ;
 assign wire20072 = ( n_n707 ) | ( wire4817 ) | ( wire20070 ) ;
 assign wire20073 = ( wire20072 ) | ( n_n100  &  wire1664 ) ;
 assign wire20075 = ( n_n100  &  n_n81 ) | ( n_n94  &  n_n39 ) ;
 assign wire20076 = ( n_n100  &  n_n33 ) | ( n_n94  &  wire57 ) ;
 assign wire20081 = ( n_n37  &  n_n100 ) | ( n_n100  &  n_n84 ) | ( n_n100  &  n_n104 ) ;
 assign wire20083 = ( wire877 ) | ( wire20081 ) | ( n_n94  &  wire112 ) ;
 assign wire20084 = ( wire4808 ) | ( wire4807 ) ;
 assign wire20085 = ( wire153 ) | ( wire57 ) | ( n_n279  &  wire914 ) ;
 assign wire20086 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire898 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire20087 = ( i_14_  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire904 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire904 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire904 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire904 ) ;
 assign wire20088 = ( n_n100  &  wire219 ) | ( n_n100  &  wire1936 ) | ( n_n100  &  wire20085 ) ;
 assign wire20089 = ( i_14_  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire906 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire20090 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire900 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire900 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire900 ) ;
 assign wire20092 = ( wire255 ) | ( wire254 ) ;
 assign wire20093 = ( wire99 ) | ( wire224 ) | ( wire41 ) ;
 assign wire20094 = ( wire4800 ) | ( n_n100  &  wire20092 ) | ( n_n100  &  wire20093 ) ;
 assign wire20095 = ( wire4805 ) | ( wire20083 ) | ( wire20084 ) | ( wire20088 ) ;
 assign wire20096 = ( n_n94  &  n_n73 ) | ( n_n94  &  n_n281  &  wire905 ) ;
 assign wire20099 = ( n_n110  &  n_n94 ) | ( n_n100  &  n_n104 ) ;
 assign wire20100 = ( n_n100  &  n_n84 ) | ( n_n94  &  n_n68 ) ;
 assign wire20101 = ( n_n133  &  n_n94 ) | ( n_n94  &  n_n16 ) | ( n_n94  &  n_n22 ) ;
 assign wire20103 = ( n_n2713 ) | ( wire20100 ) ;
 assign wire20104 = ( wire381 ) | ( wire20099 ) | ( wire20101 ) ;
 assign wire20107 = ( n_n281  &  wire903 ) | ( wire911  &  n_n220 ) ;
 assign wire20108 = ( n_n10  &  n_n100 ) | ( n_n147  &  n_n94 ) ;
 assign wire20111 = ( wire4766 ) | ( wire20108 ) | ( n_n100  &  n_n63 ) ;
 assign wire20113 = ( n_n2702 ) | ( wire687 ) | ( n_n2671 ) | ( wire20111 ) ;
 assign wire20115 = ( n_n2659 ) | ( wire20054 ) | ( wire20055 ) | ( wire20113 ) ;
 assign wire20117 = ( n_n54  &  n_n6 ) | ( n_n56  &  wire72 ) ;
 assign wire20119 = ( n_n4892 ) | ( n_n4895 ) | ( wire5035 ) | ( wire5036 ) ;
 assign wire20121 = ( n_n57  &  n_n11 ) | ( n_n57  &  n_n65 ) | ( n_n57  &  wire73 ) ;
 assign wire20122 = ( n_n4898 ) | ( wire5013 ) | ( wire5014 ) ;
 assign wire20125 = ( n_n46 ) | ( n_n92 ) | ( wire19577 ) | ( wire19578 ) ;
 assign wire20126 = ( wire51 ) | ( n_n105 ) | ( n_n43 ) | ( wire59 ) ;
 assign wire20129 = ( wire389 ) | ( n_n4585 ) | ( wire4750 ) | ( wire4751 ) ;
 assign wire20131 = ( n_n6  &  wire368 ) | ( n_n6  &  n_n41 ) | ( n_n6  &  n_n88 ) ;
 assign wire20132 = ( wire89 ) | ( wire901  &  n_n222 ) | ( wire901  &  n_n258 ) ;
 assign wire20133 = ( n_n34 ) | ( n_n82 ) | ( wire47 ) | ( wire86 ) ;
 assign wire20134 = ( n_n1497 ) | ( n_n6  &  wire1927 ) ;
 assign wire20136 = ( wire88 ) | ( n_n222  &  wire902 ) | ( wire902  &  n_n258 ) ;
 assign wire20137 = ( n_n5  &  wire67 ) | ( n_n5  &  n_n258  &  wire912 ) ;
 assign wire20141 = ( n_n4635 ) | ( wire20137 ) | ( n_n6  &  wire78 ) ;
 assign wire20142 = ( n_n4633 ) | ( n_n4636 ) | ( n_n4632 ) | ( wire4727 ) ;
 assign wire20144 = ( n_n46 ) | ( n_n92 ) | ( wire19577 ) | ( wire19578 ) ;
 assign wire20145 = ( n_n1505 ) | ( n_n5  &  wire1928 ) ;
 assign wire20147 = ( wire4720 ) | ( wire4745 ) | ( wire20131 ) | ( wire20145 ) ;
 assign wire20149 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n228 ) ;
 assign wire20150 = ( n_n216 ) | ( wire88 ) | ( n_n222  &  wire902 ) ;
 assign wire20152 = ( wire4711 ) | ( n_n5  &  wire1939 ) ;
 assign wire20153 = ( n_n4624 ) | ( wire411 ) | ( n_n6  &  wire1946 ) ;
 assign wire20155 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire911 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire911 ) ;
 assign wire20156 = ( n_n203 ) | ( wire20149 ) | ( wire911  &  n_n258 ) ;
 assign wire20157 = ( n_n1476 ) | ( n_n5  &  wire1926 ) ;
 assign wire20160 = ( n_n25 ) | ( n_n23 ) | ( wire74 ) | ( wire19457 ) ;
 assign wire20161 = ( wire40 ) | ( n_n31 ) | ( n_n200 ) | ( wire104 ) ;
 assign wire20164 = ( n_n6  &  wire40 ) | ( n_n6  &  n_n103 ) | ( n_n6  &  wire1904 ) ;
 assign wire20166 = ( n_n1490 ) | ( n_n4628 ) | ( wire4696 ) | ( wire20164 ) ;
 assign wire20169 = ( n_n4806 ) | ( wire4690 ) | ( n_n5  &  wire72 ) ;
 assign wire20171 = ( n_n11 ) | ( n_n7 ) | ( wire50 ) | ( wire95 ) ;
 assign wire20173 = ( n_n10 ) | ( wire50 ) | ( n_n59 ) | ( wire113 ) ;
 assign wire20174 = ( n_n6  &  n_n226 ) | ( n_n5  &  wire208 ) ;
 assign wire20176 = ( n_n3806 ) | ( n_n3803 ) | ( wire20174 ) ;
 assign wire20179 = ( wire95 ) | ( wire256 ) | ( n_n228  &  wire912 ) ;
 assign wire20180 = ( wire898  &  n_n228 ) | ( n_n281  &  wire906 ) ;
 assign wire20182 = ( wire44 ) | ( n_n65 ) | ( n_n252 ) | ( wire73 ) ;
 assign wire20184 = ( n_n4605 ) | ( wire4680 ) | ( wire4691 ) | ( wire20169 ) ;
 assign wire20186 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) ;
 assign wire20188 = ( i_7_  &  i_6_  &  n_n230  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n230  &  n_n116 ) ;
 assign wire20190 = ( n_n5673 ) | ( n_n5675 ) | ( wire20188 ) ;
 assign wire20191 = ( n_n5677 ) | ( wire20186 ) | ( n_n128  &  wire371 ) ;
 assign wire20192 = ( n_n122  &  n_n109 ) | ( n_n121  &  wire371 ) | ( n_n122  &  wire371 ) ;
 assign wire20193 = ( n_n111  &  n_n56 ) | ( n_n56  &  n_n38 ) | ( n_n56  &  wire453 ) ;
 assign wire20194 = ( wire55 ) | ( wire245 ) | ( wire912  &  n_n225 ) ;
 assign wire20195 = ( wire55 ) | ( wire245 ) | ( wire912  &  n_n225 ) ;
 assign wire20199 = ( n_n4671 ) | ( wire4656 ) | ( n_n56  &  n_n95 ) ;
 assign wire20200 = ( n_n4675 ) | ( n_n4674 ) | ( n_n4676 ) | ( n_n1598 ) ;
 assign wire20203 = ( n_n57  &  n_n32 ) | ( n_n56  &  n_n32 ) | ( n_n57  &  wire85 ) ;
 assign wire20205 = ( n_n56  &  wire1547 ) | ( n_n57  &  wire1950 ) ;
 assign wire20206 = ( wire460 ) | ( n_n4666 ) | ( wire20193 ) | ( wire20203 ) ;
 assign wire20209 = ( wire553 ) | ( n_n3710 ) | ( wire20206 ) ;
 assign wire20212 = ( wire826 ) | ( n_n57  &  n_n99 ) | ( n_n57  &  n_n54 ) ;
 assign wire20213 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign wire20215 = ( wire4636 ) | ( n_n57  &  n_n52 ) | ( n_n57  &  wire96 ) ;
 assign wire20216 = ( n_n4687 ) | ( n_n4686 ) | ( wire4641 ) | ( wire20212 ) ;
 assign wire20219 = ( n_n4685 ) | ( n_n57  &  wire1878 ) ;
 assign wire20220 = ( n_n4681 ) | ( n_n56  &  wire98 ) | ( n_n56  &  wire1577 ) ;
 assign wire20224 = ( n_n4920 ) | ( n_n4922 ) | ( n_n4921 ) ;
 assign wire20227 = ( n_n4923 ) | ( n_n56  &  wire1898 ) ;
 assign wire20228 = ( n_n4907 ) | ( wire636 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire20232 = ( n_n4259 ) | ( wire465 ) | ( n_n3708 ) | ( wire20227 ) ;
 assign wire20236 = ( n_n5671 ) | ( n_n5659 ) | ( wire4618 ) ;
 assign wire20238 = ( wire4617 ) | ( wire20190 ) | ( wire20191 ) | ( wire20236 ) ;
 assign wire20240 = ( n_n4598 ) | ( wire20215 ) | ( wire20216 ) | ( wire20238 ) ;
 assign wire20245 = ( n_n4534 ) | ( n_n4533 ) | ( n_n4532 ) | ( n_n4531 ) ;
 assign wire20248 = ( n_n48  &  n_n258  &  wire912 ) | ( n_n48  &  wire912  &  n_n256 ) ;
 assign wire20253 = ( wire462 ) | ( wire464 ) | ( wire376 ) | ( wire20248 ) ;
 assign wire20254 = ( n_n4094 ) | ( n_n4124 ) | ( n_n4090 ) | ( wire483 ) ;
 assign wire20256 = ( n_n25 ) | ( n_n23 ) | ( wire74 ) | ( wire19457 ) ;
 assign wire20257 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n20 ) | ( n_n53  &  n_n19 ) ;
 assign wire20258 = ( n_n28 ) | ( n_n78 ) | ( wire80 ) | ( wire65 ) ;
 assign wire20259 = ( n_n53  &  n_n197 ) | ( n_n48  &  wire69 ) ;
 assign wire20262 = ( n_n4168 ) | ( n_n4073 ) | ( wire4593 ) | ( wire20257 ) ;
 assign wire20264 = ( n_n48  &  n_n258  &  wire897 ) | ( n_n53  &  n_n258  &  wire897 ) ;
 assign wire20265 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n78 ) | ( n_n53  &  n_n26 ) ;
 assign wire20268 = ( wire478 ) | ( wire20265 ) | ( n_n48  &  wire40 ) ;
 assign wire20269 = ( wire20264 ) | ( n_n53  &  wire141 ) | ( n_n53  &  wire1363 ) ;
 assign wire20271 = ( n_n3991 ) | ( wire20268 ) | ( wire20269 ) ;
 assign wire20273 = ( n_n53  &  n_n8 ) | ( n_n53  &  n_n281  &  wire908 ) ;
 assign wire20275 = ( n_n53  &  n_n148 ) | ( n_n53  &  wire901  &  n_n228 ) ;
 assign wire20277 = ( n_n53  &  n_n61 ) | ( n_n53  &  n_n228  &  wire902 ) ;
 assign wire20278 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n148 ) ;
 assign wire20279 = ( n_n48  &  n_n11 ) | ( n_n48  &  n_n147 ) | ( n_n48  &  n_n246 ) ;
 assign wire20282 = ( wire882 ) | ( wire20277 ) | ( wire20278 ) | ( wire20279 ) ;
 assign wire20284 = ( n_n203 ) | ( n_n68 ) | ( wire514 ) | ( wire20149 ) ;
 assign wire20285 = ( n_n48  &  wire911  &  n_n258 ) | ( n_n48  &  wire899  &  n_n258 ) ;
 assign wire20287 = ( wire456 ) | ( n_n4165 ) | ( wire20285 ) ;
 assign wire20289 = ( n_n20 ) | ( wire79 ) | ( n_n281  &  wire906 ) ;
 assign wire20290 = ( wire44 ) | ( n_n221 ) | ( n_n252 ) | ( wire469 ) ;
 assign wire20293 = ( wire675 ) | ( wire4551 ) | ( wire4573 ) | ( wire4574 ) ;
 assign wire20297 = ( n_n97 ) | ( n_n51 ) | ( wire71 ) | ( wire19575 ) ;
 assign wire20299 = ( wire571 ) | ( n_n48  &  wire900  &  n_n258 ) ;
 assign wire20300 = ( wire737 ) | ( wire5591 ) | ( wire5592 ) ;
 assign wire20301 = ( wire407 ) | ( wire457 ) | ( n_n53  &  wire77 ) ;
 assign wire20304 = ( n_n4183 ) | ( wire20299 ) | ( n_n48  &  wire1234 ) ;
 assign wire20306 = ( n_n113 ) | ( n_n85 ) | ( wire102 ) | ( wire87 ) ;
 assign wire20307 = ( n_n220  &  wire904 ) | ( n_n256  &  wire904 ) | ( n_n220  &  wire907 ) | ( n_n256  &  wire907 ) ;
 assign wire20308 = ( n_n37 ) | ( wire89 ) | ( n_n82 ) | ( wire47 ) ;
 assign wire20309 = ( wire86 ) | ( wire20307 ) | ( wire901  &  n_n256 ) ;
 assign wire20310 = ( n_n53  &  wire901  &  n_n258 ) | ( n_n53  &  n_n258  &  wire912 ) ;
 assign wire20313 = ( n_n97 ) | ( n_n51 ) | ( wire71 ) | ( wire19575 ) ;
 assign wire20314 = ( n_n99 ) | ( n_n43 ) | ( wire59 ) | ( wire96 ) ;
 assign wire20315 = ( wire51 ) | ( wire19578 ) | ( n_n222  &  wire906 ) ;
 assign wire20316 = ( n_n46 ) | ( n_n43 ) | ( wire59 ) | ( wire19577 ) ;
 assign wire20319 = ( n_n4179 ) | ( wire809 ) | ( wire4523 ) | ( wire4524 ) ;
 assign wire20323 = ( n_n48  &  n_n11 ) | ( n_n53  &  n_n63 ) ;
 assign wire20324 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n246 ) ;
 assign wire20325 = ( n_n106  &  n_n53 ) | ( n_n48  &  n_n86 ) ;
 assign wire20330 = ( wire631 ) | ( wire462 ) | ( wire464 ) | ( wire20323 ) ;
 assign wire20331 = ( n_n4124 ) | ( n_n4090 ) | ( wire20324 ) | ( wire20325 ) ;
 assign wire20334 = ( n_n48  &  n_n226 ) | ( n_n48  &  n_n281  &  wire913 ) ;
 assign wire20336 = ( n_n53  &  n_n226 ) | ( n_n53  &  n_n281  &  wire903 ) ;
 assign wire20337 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n144 ) | ( n_n53  &  n_n257 ) ;
 assign wire20340 = ( wire4520 ) | ( wire20334 ) | ( wire20337 ) ;
 assign wire20341 = ( n_n4094 ) | ( wire20336 ) | ( n_n48  &  wire1089 ) ;
 assign wire20343 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n70 ) | ( n_n53  &  n_n19 ) ;
 assign wire20344 = ( n_n53  &  n_n220  &  wire908 ) | ( n_n53  &  n_n256  &  wire908 ) ;
 assign wire20346 = ( n_n53  &  n_n60 ) | ( n_n48  &  n_n148 ) ;
 assign wire20347 = ( n_n53  &  n_n108 ) | ( n_n53  &  n_n257 ) | ( n_n53  &  n_n226 ) ;
 assign wire20349 = ( wire20347 ) | ( n_n4068 ) ;
 assign wire20350 = ( wire626 ) | ( n_n1433 ) | ( wire20343 ) | ( wire20346 ) ;
 assign wire20353 = ( wire298 ) | ( n_n4146 ) | ( wire20349 ) | ( wire20350 ) ;
 assign wire20355 = ( n_n4141 ) | ( n_n3900 ) | ( n_n3899 ) | ( n_n3901 ) ;
 assign wire20356 = ( n_n6  &  n_n60 ) | ( n_n6  &  n_n9 ) | ( n_n6  &  wire63 ) ;
 assign wire20358 = ( wire44 ) | ( n_n252 ) | ( n_n68 ) | ( wire514 ) ;
 assign wire20359 = ( wire62 ) | ( n_n16 ) | ( n_n15 ) | ( wire20155 ) ;
 assign wire20362 = ( (~ i_14_)  &  i_15_  &  n_n275  &  n_n254 ) | ( i_14_  &  (~ i_15_)  &  n_n275  &  n_n254 ) ;
 assign wire20364 = ( n_n151  &  n_n6 ) | ( n_n207  &  wire232 ) ;
 assign wire20365 = ( wire913  &  n_n258 ) | ( n_n228  &  wire897 ) ;
 assign wire20366 = ( n_n207  &  n_n67 ) | ( n_n207  &  n_n258  &  wire905 ) ;
 assign wire20367 = ( n_n9  &  n_n207 ) | ( n_n100  &  n_n104 ) ;
 assign wire20369 = ( n_n4  &  n_n31 ) | ( n_n10  &  n_n100 ) ;
 assign wire20370 = ( n_n100  &  n_n279  &  wire901 ) | ( n_n100  &  wire901  &  n_n228 ) ;
 assign wire20371 = ( n_n106  &  n_n100 ) | ( n_n100  &  n_n33 ) | ( n_n100  &  n_n81 ) ;
 assign wire20374 = ( wire434 ) | ( wire20369 ) | ( wire20370 ) | ( wire20371 ) ;
 assign wire20376 = ( wire901  &  n_n228 ) | ( n_n281  &  wire906 ) ;
 assign wire20379 = ( n_n6  &  n_n226 ) | ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) ;
 assign wire20381 = ( wire20379 ) | ( n_n6  &  wire1371 ) ;
 assign wire20382 = ( n_n4823 ) | ( n_n4605 ) | ( wire4506 ) | ( wire20356 ) ;
 assign wire20385 = ( n_n53  &  n_n108 ) | ( n_n53  &  n_n70 ) | ( n_n53  &  n_n61 ) ;
 assign wire20387 = ( n_n53  &  n_n78 ) | ( n_n53  &  wire899  &  n_n258 ) ;
 assign wire20390 = ( n_n1  &  wire68 ) | ( n_n53  &  n_n257 ) ;
 assign wire20392 = ( n_n4068 ) | ( n_n4069 ) | ( wire20390 ) ;
 assign wire20397 = ( n_n4  &  n_n197 ) | ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) ;
 assign wire20400 = ( n_n1341 ) | ( n_n884 ) | ( n_n876 ) | ( wire4478 ) ;
 assign wire20401 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n108 ) | ( n_n4  &  n_n70 ) ;
 assign wire20403 = ( n_n896 ) | ( n_n2986 ) | ( wire20401 ) ;
 assign wire20404 = ( n_n4  &  n_n13 ) | ( n_n4  &  wire900  &  n_n220 ) ;
 assign wire20405 = ( n_n4  &  n_n9 ) | ( n_n4  &  n_n281  &  wire906 ) ;
 assign wire20408 = ( wire20405 ) | ( n_n4  &  n_n65 ) | ( n_n4  &  n_n61 ) ;
 assign wire20409 = ( wire446 ) | ( n_n2982 ) | ( wire20404 ) ;
 assign wire20412 = ( wire876 ) | ( wire533 ) | ( wire20408 ) | ( wire20409 ) ;
 assign wire20414 = ( wire60 ) | ( wire19738 ) | ( wire913  &  n_n256 ) ;
 assign wire20415 = ( n_n12 ) | ( n_n204 ) | ( wire73 ) | ( wire52 ) ;
 assign wire20416 = ( n_n110 ) | ( wire44 ) | ( n_n65 ) | ( wire70 ) ;
 assign wire20418 = ( n_n53  &  n_n148 ) | ( n_n53  &  wire901  &  n_n228 ) ;
 assign wire20419 = ( n_n53  &  n_n10 ) | ( n_n53  &  n_n220  &  wire905 ) ;
 assign wire20422 = ( n_n3581 ) | ( n_n4160 ) | ( wire20418 ) | ( wire20419 ) ;
 assign wire20423 = ( wire75 ) | ( n_n206 ) | ( n_n281  &  wire913 ) ;
 assign wire20424 = ( wire407 ) | ( n_n53  &  n_n228  &  wire902 ) ;
 assign wire20425 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n7 ) | ( n_n53  &  n_n144 ) ;
 assign wire20429 = ( wire516 ) | ( wire676 ) | ( wire882 ) | ( wire20424 ) ;
 assign wire20430 = ( n_n3791 ) | ( wire20425 ) | ( n_n53  &  wire1900 ) ;
 assign wire20433 = ( n_n34 ) | ( n_n43 ) | ( wire59 ) | ( wire86 ) ;
 assign wire20434 = ( n_n6  &  wire368 ) | ( n_n6  &  n_n88 ) | ( n_n6  &  n_n104 ) ;
 assign wire20435 = ( wire20434 ) | ( n_n6  &  wire1927 ) ;
 assign wire20437 = ( n_n6  &  wire69 ) | ( n_n6  &  n_n258  &  wire897 ) ;
 assign wire20438 = ( n_n6  &  n_n25 ) | ( n_n6  &  wire78 ) | ( n_n6  &  wire19457 ) ;
 assign wire20441 = ( n_n6  &  wire1868 ) | ( n_n6  &  wire1904 ) ;
 assign wire20442 = ( n_n4633 ) | ( n_n4632 ) | ( wire20438 ) ;
 assign wire20444 = ( n_n54  &  n_n6 ) | ( n_n53  &  n_n32 ) ;
 assign wire20445 = ( n_n53  &  n_n63 ) | ( n_n53  &  n_n258  &  wire907 ) ;
 assign wire20449 = ( wire389 ) | ( wire882 ) | ( wire20444 ) | ( wire20445 ) ;
 assign wire20450 = ( wire670 ) | ( n_n3019 ) | ( wire4423 ) ;
 assign wire20452 = ( n_n2890 ) | ( wire20449 ) | ( wire20450 ) ;
 assign wire20454 = ( wire453 ) | ( n_n220  &  wire914 ) | ( n_n256  &  wire914 ) ;
 assign wire20455 = ( n_n53  &  n_n37 ) | ( n_n53  &  n_n32 ) | ( n_n53  &  n_n104 ) ;
 assign wire20457 = ( n_n3019 ) | ( wire20455 ) | ( n_n53  &  wire1900 ) ;
 assign wire20460 = ( wire4418 ) | ( wire571 ) ;
 assign wire20461 = ( wire407 ) | ( wire579 ) | ( n_n53  &  wire68 ) ;
 assign wire20463 = ( n_n281  &  wire903 ) | ( n_n228  &  wire902 ) ;
 assign wire20465 = ( wire113 ) | ( wire72 ) ;
 assign wire20466 = ( wire101 ) | ( wire20463 ) | ( n_n281  &  wire914 ) ;
 assign wire20467 = ( n_n206 ) | ( wire118 ) | ( wire50 ) | ( n_n59 ) ;
 assign wire20469 = ( n_n4381 ) | ( wire4417 ) | ( wire20460 ) | ( wire20461 ) ;
 assign wire20470 = ( wire81 ) | ( n_n220  &  wire904 ) ;
 assign wire20471 = ( n_n93 ) | ( n_n90 ) | ( wire76 ) | ( wire19384 ) ;
 assign wire20472 = ( n_n42 ) | ( n_n179 ) | ( wire55 ) | ( wire57 ) ;
 assign wire20474 = ( n_n53  &  wire204 ) | ( n_n53  &  wire43 ) | ( n_n53  &  wire19506 ) ;
 assign wire20475 = ( wire20474 ) | ( wire4409 ) ;
 assign wire20479 = ( n_n1433 ) | ( wire478 ) | ( wire20343 ) | ( wire20344 ) ;
 assign wire20480 = ( n_n53  &  wire1445 ) | ( n_n53  &  wire1948 ) ;
 assign wire20482 = ( wire406 ) | ( n_n3587 ) | ( wire20479 ) | ( wire20480 ) ;
 assign wire20484 = ( n_n2824 ) | ( wire4463 ) | ( wire20422 ) | ( wire20482 ) ;
 assign wire20486 = ( n_n57  &  n_n32 ) | ( n_n57  &  n_n81 ) | ( n_n57  &  wire86 ) ;
 assign wire20488 = ( wire20486 ) | ( n_n57  &  wire1950 ) ;
 assign wire20490 = ( wire60 ) | ( wire73 ) | ( n_n281  &  wire906 ) ;
 assign wire20491 = ( n_n110 ) | ( wire44 ) | ( n_n65 ) | ( wire70 ) ;
 assign wire20492 = ( n_n57  &  n_n108 ) | ( n_n57  &  n_n11 ) | ( n_n57  &  wire95 ) ;
 assign wire20495 = ( n_n4920 ) | ( n_n4912 ) | ( wire20492 ) ;
 assign wire20497 = ( n_n100  &  n_n60 ) | ( n_n100  &  n_n258  &  wire907 ) ;
 assign wire20499 = ( n_n57  &  n_n95 ) | ( n_n151  &  n_n100 ) ;
 assign wire20501 = ( n_n57  &  n_n93 ) | ( n_n57  &  wire76 ) | ( n_n57  &  wire1878 ) ;
 assign wire20502 = ( n_n4686 ) | ( wire4373 ) | ( wire20499 ) ;
 assign wire20505 = ( n_n16 ) | ( n_n68 ) | ( wire514 ) | ( wire20155 ) ;
 assign wire20506 = ( n_n100  &  wire83 ) | ( n_n100  &  wire911  &  n_n258 ) ;
 assign wire20508 = ( n_n3604 ) | ( wire740 ) | ( wire20506 ) ;
 assign wire20510 = ( wire901  &  n_n228 ) | ( n_n281  &  wire906 ) ;
 assign wire20512 = ( wire20510 ) | ( wire132 ) ;
 assign wire20513 = ( n_n257 ) | ( wire75 ) | ( n_n206 ) | ( wire72 ) ;
 assign wire20514 = ( wire160 ) | ( n_n65 ) | ( wire184 ) | ( wire73 ) ;
 assign wire20516 = ( wire725 ) | ( n_n3864 ) | ( wire4380 ) | ( wire20497 ) ;
 assign wire20519 = ( n_n100  &  n_n25 ) | ( n_n100  &  n_n103 ) | ( n_n100  &  wire19457 ) ;
 assign wire20520 = ( n_n241  &  wire901  &  n_n258 ) | ( n_n241  &  n_n258  &  wire897 ) ;
 assign wire20522 = ( n_n241  &  n_n105 ) | ( n_n54  &  n_n100 ) ;
 assign wire20524 = ( wire20520 ) | ( n_n177  &  n_n112 ) | ( n_n177  &  n_n35 ) ;
 assign wire20525 = ( wire559 ) | ( wire20522 ) | ( n_n177  &  n_n200 ) ;
 assign wire20526 = ( wire67 ) | ( wire87 ) | ( wire914  &  n_n225 ) ;
 assign wire20527 = ( n_n258  &  wire912 ) | ( wire901  &  n_n225 ) ;
 assign wire20528 = ( wire51 ) | ( n_n222  &  wire907 ) ;
 assign wire20529 = ( wire368 ) | ( n_n88 ) | ( wire20527 ) ;
 assign wire20530 = ( n_n34 ) | ( n_n43 ) | ( wire59 ) | ( wire86 ) ;
 assign wire20532 = ( n_n100  &  n_n279  &  wire907 ) | ( n_n100  &  n_n228  &  wire907 ) ;
 assign wire20533 = ( n_n37  &  n_n100 ) | ( n_n100  &  n_n84 ) | ( n_n100  &  n_n104 ) ;
 assign wire20536 = ( n_n100  &  n_n220  &  wire907 ) | ( n_n100  &  n_n256  &  wire907 ) ;
 assign wire20537 = ( n_n100  &  wire77 ) | ( n_n100  &  wire900  &  n_n258 ) ;
 assign wire20540 = ( n_n3884 ) | ( wire4330 ) | ( wire20536 ) | ( wire20537 ) ;
 assign wire20541 = ( wire383 ) | ( n_n100  &  wire202 ) | ( n_n100  &  wire19576 ) ;
 assign wire20542 = ( wire628 ) | ( wire20519 ) | ( wire20524 ) | ( wire20525 ) ;
 assign wire20543 = ( wire20540 ) | ( n_n100  &  wire1540 ) | ( n_n100  &  wire1903 ) ;
 assign wire20547 = ( wire56 ) | ( wire19407 ) | ( n_n256  &  wire897 ) ;
 assign wire20548 = ( wire82 ) | ( n_n171 ) | ( n_n22 ) | ( wire53 ) ;
 assign wire20549 = ( n_n4922 ) | ( n_n4921 ) | ( wire693 ) ;
 assign wire20551 = ( wire385 ) | ( wire4322 ) | ( wire20549 ) ;
 assign wire20553 = ( n_n2832 ) | ( n_n2830 ) | ( wire20551 ) ;
 assign wire20555 = ( wire81 ) | ( n_n220  &  wire904 ) ;
 assign wire20556 = ( n_n179 ) | ( n_n90 ) | ( wire57 ) | ( wire19384 ) ;
 assign wire20557 = ( n_n42 ) | ( n_n44 ) | ( wire55 ) | ( wire19385 ) ;
 assign wire20559 = ( n_n1  &  wire179 ) | ( n_n1  &  wire204 ) | ( n_n1  &  wire1877 ) ;
 assign wire20562 = ( n_n3259 ) | ( n_n3260 ) | ( wire4313 ) ;
 assign wire20566 = ( n_n1  &  wire1483 ) | ( n_n1  &  wire1953 ) ;
 assign wire20568 = ( n_n2860 ) | ( wire814 ) | ( n_n3768 ) | ( wire20566 ) ;
 assign wire20571 = ( n_n2798 ) | ( n_n2797 ) | ( n_n2796 ) ;
 assign wire20573 = ( n_n38 ) | ( n_n35 ) | ( wire64 ) | ( wire453 ) ;
 assign wire20574 = ( n_n111 ) | ( wire85 ) | ( n_n90 ) | ( wire19384 ) ;
 assign wire20575 = ( wire89 ) | ( n_n81 ) | ( n_n83 ) | ( wire86 ) ;
 assign wire20576 = ( n_n42 ) | ( n_n179 ) | ( wire55 ) | ( wire57 ) ;
 assign wire20579 = ( wire60 ) | ( wire84 ) | ( n_n279  &  wire913 ) ;
 assign wire20581 = ( n_n4  &  n_n108 ) | ( n_n4  &  wire44 ) | ( n_n4  &  n_n65 ) ;
 assign wire20583 = ( wire20581 ) | ( n_n4  &  wire111 ) | ( n_n4  &  wire1693 ) ;
 assign wire20585 = ( wire903  &  n_n220 ) | ( n_n220  &  wire907 ) ;
 assign wire20588 = ( wire485 ) | ( n_n3731 ) | ( wire4285 ) ;
 assign wire20590 = ( wire640 ) | ( wire867 ) | ( wire792 ) | ( wire20588 ) ;
 assign wire20592 = ( n_n102 ) | ( n_n52 ) | ( wire807 ) | ( wire96 ) ;
 assign wire20593 = ( n_n281  &  wire903 ) | ( n_n228  &  wire902 ) ;
 assign wire20595 = ( wire113 ) | ( wire72 ) ;
 assign wire20596 = ( wire75 ) | ( wire20593 ) | ( n_n281  &  wire913 ) ;
 assign wire20597 = ( n_n206 ) | ( wire118 ) | ( wire50 ) | ( n_n59 ) ;
 assign wire20600 = ( wire782 ) | ( n_n3757 ) | ( n_n265  &  wire277 ) ;
 assign wire20601 = ( n_n11 ) | ( n_n148 ) | ( wire101 ) | ( wire95 ) ;
 assign wire20602 = ( n_n110 ) | ( n_n12 ) | ( wire70 ) | ( wire73 ) ;
 assign wire20604 = ( n_n1  &  n_n108 ) | ( n_n1  &  n_n112 ) | ( n_n1  &  wire84 ) ;
 assign wire20606 = ( n_n3524 ) | ( wire468 ) | ( wire20604 ) ;
 assign wire20608 = ( n_n4  &  n_n95 ) | ( n_n265  &  n_n62 ) ;
 assign wire20609 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n47 ) | ( n_n4  &  wire68 ) ;
 assign wire20610 = ( wire20609 ) | ( wire20608 ) ;
 assign wire20611 = ( wire4267 ) | ( n_n4  &  wire1924 ) ;
 assign wire20614 = ( wire4276 ) | ( wire4281 ) | ( wire20600 ) | ( wire20606 ) ;
 assign wire20616 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n258  &  wire905 ) ;
 assign wire20617 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n7 ) | ( n_n4  &  n_n144 ) ;
 assign wire20620 = ( n_n4  &  n_n12 ) | ( n_n4  &  n_n64 ) | ( n_n4  &  n_n13 ) ;
 assign wire20622 = ( n_n4015 ) | ( wire4248 ) | ( wire20620 ) ;
 assign wire20624 = ( n_n2840 ) | ( n_n2839 ) | ( wire20622 ) ;
 assign wire20625 = ( n_n2808 ) | ( n_n2806 ) | ( wire20590 ) | ( wire20624 ) ;
 assign wire20629 = ( n_n121  &  wire216 ) | ( n_n132  &  n_n107 ) ;
 assign wire20630 = ( n_n122  &  wire1707 ) | ( n_n130  &  wire1706 ) ;
 assign wire20633 = ( n_n118  &  n_n260  &  n_n155 ) | ( n_n118  &  n_n155  &  n_n284 ) ;
 assign wire20635 = ( wire20633 ) | ( n_n118  &  n_n264  &  n_n155 ) ;
 assign wire20636 = ( n_n5664 ) | ( n_n272  &  wire930 ) | ( n_n272  &  wire1740 ) ;
 assign wire20637 = ( n_n260  &  n_n229  &  n_n165 ) | ( n_n229  &  n_n165  &  n_n284 ) ;
 assign wire20638 = ( n_n260  &  n_n283  &  n_n165 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign wire20641 = ( n_n260  &  n_n155  &  n_n116 ) | ( n_n155  &  n_n284  &  n_n116 ) ;
 assign wire20642 = ( n_n264  &  n_n155  &  n_n116 ) | ( n_n155  &  n_n230  &  n_n116 ) ;
 assign wire20643 = ( n_n272  &  n_n260  &  n_n116 ) | ( n_n272  &  n_n230  &  n_n116 ) ;
 assign wire20645 = ( wire20643 ) | ( wire20642 ) ;
 assign wire20646 = ( n_n5676 ) | ( wire20641 ) | ( n_n128  &  wire216 ) ;
 assign wire20648 = ( wire20635 ) | ( wire20636 ) | ( wire20645 ) | ( wire20646 ) ;
 assign wire20651 = ( n_n177  &  n_n112 ) | ( n_n189  &  n_n109 ) ;
 assign wire20652 = ( n_n189  &  n_n102 ) | ( n_n177  &  n_n35 ) ;
 assign wire20655 = ( n_n255  &  n_n197 ) | ( n_n241  &  n_n103 ) ;
 assign wire20657 = ( wire559 ) | ( n_n255  &  wire950 ) ;
 assign wire20658 = ( wire392 ) | ( wire20655 ) | ( n_n241  &  n_n104 ) ;
 assign wire20662 = ( i_1_  &  i_2_  &  i_0_ ) | ( i_3_  &  i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire20665 = ( wire535 ) | ( wire777 ) | ( wire926 ) | ( n_n5675 ) ;
 assign wire20667 = ( n_n153  &  n_n260  &  n_n165 ) | ( n_n153  &  n_n165  &  n_n284 ) ;
 assign wire20668 = ( n_n272  &  n_n260  &  n_n165 ) | ( n_n272  &  n_n165  &  n_n284 ) ;
 assign wire20671 = ( n_n5796 ) | ( wire4202 ) | ( wire20668 ) ;
 assign wire20675 = ( n_n4287 ) | ( wire389 ) | ( wire632 ) | ( wire5613 ) ;
 assign wire20677 = ( wire153  &  n_n6 ) | ( n_n6  &  wire224 ) ;
 assign wire20678 = ( n_n6  &  wire166 ) | ( n_n5  &  wire166 ) | ( n_n6  &  wire180 ) ;
 assign wire20682 = ( n_n4895 ) | ( wire5013 ) | ( wire5014 ) ;
 assign wire20683 = ( n_n4892 ) | ( n_n4898 ) | ( wire5035 ) | ( wire5036 ) ;
 assign wire20686 = ( n_n4210 ) | ( wire878 ) | ( wire20682 ) | ( wire20683 ) ;
 assign wire20688 = ( n_n5  &  wire99 ) | ( n_n5  &  wire1894 ) ;
 assign wire20689 = ( n_n4870 ) | ( n_n4871 ) | ( wire4183 ) | ( wire5091 ) ;
 assign wire20691 = ( wire5099 ) | ( wire19862 ) | ( wire20688 ) | ( wire20689 ) ;
 assign wire20692 = ( n_n5796 ) | ( n_n56  &  wire49 ) ;
 assign wire20694 = ( n_n57  &  wire190 ) | ( n_n57  &  wire212 ) ;
 assign wire20695 = ( n_n56  &  wire124 ) | ( n_n56  &  wire212 ) ;
 assign wire20696 = ( n_n57  &  wire119 ) | ( n_n56  &  wire119 ) ;
 assign wire20699 = ( n_n4926 ) | ( n_n4929 ) | ( wire20692 ) | ( wire20696 ) ;
 assign wire20701 = ( n_n56  &  wire224 ) | ( n_n56  &  wire180 ) ;
 assign wire20703 = ( wire614 ) | ( n_n57  &  wire166 ) | ( n_n56  &  wire166 ) ;
 assign wire20704 = ( n_n4967 ) | ( wire613 ) | ( wire20701 ) ;
 assign wire20705 = ( n_n57  &  wire153 ) | ( n_n56  &  wire254 ) ;
 assign wire20706 = ( n_n57  &  wire180 ) | ( n_n57  &  wire273 ) ;
 assign wire20710 = ( n_n4954 ) | ( n_n4953 ) | ( n_n4955 ) | ( wire671 ) ;
 assign wire20711 = ( n_n132  &  n_n107 ) | ( n_n139  &  wire250 ) ;
 assign wire20712 = ( n_n5796 ) | ( n_n139  &  wire899  &  n_n281 ) ;
 assign wire20714 = ( n_n5796 ) | ( n_n132  &  wire250 ) ;
 assign wire20716 = ( wire4159 ) | ( wire4170 ) | ( wire20711 ) | ( wire20714 ) ;
 assign wire20718 = ( n_n4279 ) | ( wire20703 ) | ( wire20704 ) | ( wire20716 ) ;
 assign wire20719 = ( n_n56  &  wire200 ) | ( n_n56  &  wire277 ) ;
 assign wire20720 = ( wire268  &  n_n57 ) | ( n_n57  &  wire200 ) ;
 assign wire20721 = ( wire268  &  n_n56 ) | ( n_n57  &  wire277 ) ;
 assign wire20722 = ( n_n57  &  wire157 ) | ( n_n57  &  wire112 ) | ( n_n56  &  wire112 ) ;
 assign wire20725 = ( n_n56  &  n_n223 ) | ( n_n56  &  wire42 ) | ( n_n56  &  wire1898 ) ;
 assign wire20728 = ( n_n4923 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire20729 = ( n_n4920 ) | ( n_n4907 ) | ( n_n4922 ) | ( n_n4921 ) ;
 assign wire20733 = ( n_n4261 ) | ( n_n4256 ) | ( wire465 ) | ( wire20728 ) ;
 assign wire20737 = ( n_n56  &  wire157 ) | ( n_n56  &  wire273 ) ;
 assign wire20739 = ( n_n4936 ) | ( n_n4941 ) | ( n_n4942 ) | ( n_n4938 ) ;
 assign wire20740 = ( wire760 ) | ( wire20737 ) | ( n_n57  &  wire140 ) ;
 assign wire20742 = ( n_n4218 ) | ( wire20694 ) | ( wire20695 ) | ( wire20699 ) ;
 assign wire20743 = ( wire20739 ) | ( wire20740 ) | ( wire20742 ) ;
 assign wire20745 = ( n_n5796 ) | ( n_n6  &  wire75 ) | ( n_n6  &  n_n206 ) ;
 assign wire20746 = ( n_n4806 ) | ( wire20745 ) | ( n_n5  &  wire72 ) ;
 assign wire20748 = ( n_n4223 ) | ( n_n4224 ) | ( wire20746 ) ;
 assign wire20750 = ( n_n4204 ) | ( wire19749 ) | ( wire20748 ) ;
 assign wire20751 = ( n_n4203 ) | ( n_n4206 ) | ( n_n4211 ) | ( wire20686 ) ;
 assign wire20753 = ( n_n4197 ) | ( wire20750 ) | ( wire20751 ) ;
 assign wire20755 = ( n_n177  &  n_n112 ) | ( n_n189  &  n_n109 ) ;
 assign wire20756 = ( n_n197  &  n_n100 ) | ( n_n94  &  wire77 ) ;
 assign wire20758 = ( n_n94  &  n_n216 ) | ( n_n94  &  wire913  &  n_n220 ) ;
 assign wire20759 = ( n_n100  &  n_n216 ) | ( n_n94  &  n_n17 ) ;
 assign wire20760 = ( n_n133  &  n_n94 ) | ( n_n94  &  n_n16 ) | ( n_n94  &  n_n67 ) ;
 assign wire20764 = ( wire20758 ) | ( wire20760 ) | ( n_n100  &  wire83 ) ;
 assign wire20765 = ( n_n1628 ) | ( n_n1058 ) | ( wire4120 ) | ( wire20759 ) ;
 assign wire20767 = ( n_n255  &  n_n197 ) | ( n_n241  &  n_n216 ) ;
 assign wire20769 = ( wire20755 ) | ( wire20767 ) | ( n_n54  &  n_n100 ) ;
 assign wire20770 = ( wire392 ) | ( wire386 ) | ( wire20769 ) ;
 assign wire20772 = ( wire44  &  n_n100 ) | ( n_n100  &  n_n252 ) | ( n_n100  &  n_n15 ) ;
 assign wire20774 = ( n_n100  &  wire1237 ) | ( n_n94  &  wire1910 ) ;
 assign wire20775 = ( n_n1624 ) | ( n_n3604 ) | ( wire4117 ) | ( wire20772 ) ;
 assign wire20776 = ( n_n145  &  n_n94 ) | ( n_n94  &  n_n144 ) | ( n_n94  &  wire118 ) ;
 assign wire20778 = ( wire20776 ) | ( wire44  &  n_n94 ) | ( n_n94  &  n_n252 ) ;
 assign wire20779 = ( n_n2713 ) | ( wire4100 ) | ( wire5514 ) | ( wire5515 ) ;
 assign wire20781 = ( n_n4682 ) | ( n_n4685 ) | ( wire19565 ) | ( wire20778 ) ;
 assign wire20782 = ( wire370 ) | ( wire4789 ) | ( wire4790 ) | ( wire20779 ) ;
 assign wire20784 = ( n_n57  &  wire82 ) | ( n_n57  &  n_n223 ) | ( n_n57  &  wire42 ) ;
 assign wire20785 = ( wire20784 ) | ( wire788 ) ;
 assign wire20786 = ( n_n4680 ) | ( n_n4677 ) | ( wire19534 ) | ( wire20785 ) ;
 assign wire20788 = ( n_n3398 ) | ( n_n3397 ) | ( wire20786 ) ;
 assign wire20791 = ( n_n223 ) | ( n_n20 ) | ( wire42 ) | ( wire66 ) ;
 assign wire20793 = ( n_n1320 ) | ( n_n3229 ) | ( wire4081 ) ;
 assign wire20796 = ( n_n112 ) | ( n_n67 ) | ( wire84 ) | ( wire19738 ) ;
 assign wire20797 = ( n_n110 ) | ( wire60 ) | ( n_n204 ) | ( wire52 ) ;
 assign wire20798 = ( wire4302 ) | ( n_n4  &  n_n108 ) | ( n_n4  &  n_n70 ) ;
 assign wire20800 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n258  &  wire905 ) ;
 assign wire20802 = ( n_n4005 ) | ( wire446 ) | ( wire20800 ) ;
 assign wire20804 = ( n_n3406 ) | ( wire633 ) | ( wire20802 ) ;
 assign wire20806 = ( n_n257 ) | ( wire72 ) | ( n_n281  &  wire913 ) ;
 assign wire20807 = ( wire60 ) | ( n_n204 ) | ( n_n112 ) | ( wire52 ) ;
 assign wire20808 = ( wire130 ) | ( wire210 ) | ( wire911  &  n_n228 ) ;
 assign wire20809 = ( n_n2  &  n_n226 ) | ( n_n268  &  wire247 ) ;
 assign wire20814 = ( wire557 ) | ( n_n3506 ) | ( wire485 ) | ( wire933 ) ;
 assign wire20816 = ( n_n1440 ) | ( wire5758 ) | ( wire19391 ) | ( wire20814 ) ;
 assign wire20817 = ( n_n3417 ) | ( wire597 ) | ( wire5775 ) | ( wire19383 ) ;
 assign wire20819 = ( n_n3378 ) | ( wire20816 ) | ( wire20817 ) ;
 assign wire20820 = ( n_n110  &  n_n53 ) | ( n_n48  &  wire82 ) ;
 assign wire20823 = ( n_n3309 ) | ( n_n3579 ) | ( n_n48  &  wire1938 ) ;
 assign wire20824 = ( wire4062 ) | ( wire5625 ) | ( wire5626 ) | ( wire20820 ) ;
 assign wire20826 = ( wire764 ) | ( n_n53  &  wire68 ) ;
 assign wire20827 = ( wire579 ) | ( n_n57  &  wire899  &  n_n228 ) ;
 assign wire20831 = ( wire406 ) | ( wire4044 ) | ( n_n48  &  n_n95 ) ;
 assign wire20832 = ( wire309 ) | ( wire4056 ) | ( wire20826 ) | ( wire20827 ) ;
 assign wire20833 = ( n_n1433 ) | ( n_n3587 ) | ( wire5589 ) | ( wire5590 ) ;
 assign wire20836 = ( n_n2440 ) | ( wire20831 ) | ( wire20832 ) | ( wire20833 ) ;
 assign wire20839 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire20840 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire899 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire20842 = ( wire411 ) | ( wire4036 ) | ( n_n5  &  wire255 ) ;
 assign wire20844 = ( n_n4770 ) | ( wire4035 ) | ( wire20842 ) ;
 assign wire20846 = ( wire84 ) | ( n_n279  &  wire913 ) | ( wire913  &  n_n220 ) ;
 assign wire20847 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n70 ) | ( n_n53  &  n_n19 ) ;
 assign wire20849 = ( n_n3581 ) | ( n_n1536 ) | ( wire20847 ) ;
 assign wire20851 = ( n_n53  &  n_n226 ) | ( n_n53  &  n_n258  &  wire905 ) ;
 assign wire20853 = ( n_n4154 ) | ( wire475 ) | ( wire20851 ) ;
 assign wire20854 = ( wire4016 ) | ( wire4520 ) | ( wire20334 ) ;
 assign wire20856 = ( n_n4774 ) | ( wire20853 ) | ( wire20854 ) ;
 assign wire20858 = ( n_n3393 ) | ( wire20823 ) | ( wire20824 ) | ( wire20856 ) ;
 assign wire20861 = ( n_n3523 ) | ( n_n2  &  wire1951 ) ;
 assign wire20862 = ( n_n3525 ) | ( n_n3524 ) | ( n_n2  &  wire1557 ) ;
 assign wire20865 = ( wire4005 ) | ( wire5709 ) | ( n_n1  &  n_n12 ) ;
 assign wire20866 = ( n_n3519 ) | ( n_n3520 ) | ( wire4004 ) ;
 assign wire20869 = ( n_n2  &  wire1871 ) | ( n_n2  &  wire1873 ) ;
 assign wire20870 = ( n_n1  &  wire1657 ) | ( n_n1  &  wire1923 ) ;
 assign wire20872 = ( n_n3778 ) | ( n_n2633 ) | ( wire20869 ) | ( wire20870 ) ;
 assign wire20874 = ( i_15_  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire20875 = ( i_15_  &  n_n259  &  n_n258 ) | ( i_15_  &  n_n259  &  n_n256 ) | ( (~ i_15_)  &  n_n259  &  n_n256 ) ;
 assign wire20876 = ( n_n207  &  n_n257 ) | ( n_n5  &  wire72 ) ;
 assign wire20881 = ( n_n4806 ) | ( n_n3550 ) | ( wire3988 ) | ( wire20876 ) ;
 assign wire20882 = ( n_n4  &  n_n197 ) | ( n_n4  &  n_n223 ) | ( n_n4  &  n_n221 ) ;
 assign wire20883 = ( n_n110  &  n_n94 ) | ( n_n4  &  n_n93 ) ;
 assign wire20888 = ( wire455 ) | ( wire388 ) | ( wire381 ) | ( wire20883 ) ;
 assign wire20889 = ( wire333 ) | ( n_n6820 ) | ( wire3975 ) | ( wire3976 ) ;
 assign wire20894 = ( wire639 ) | ( wire3967 ) | ( wire5656 ) | ( wire5657 ) ;
 assign wire20895 = ( n_n4809 ) | ( wire539 ) | ( wire3968 ) | ( wire20894 ) ;
 assign wire20897 = ( n_n1  &  wire68 ) | ( n_n53  &  n_n257 ) ;
 assign wire20898 = ( n_n53  &  n_n107 ) | ( n_n4  &  n_n257 ) ;
 assign wire20899 = ( n_n53  &  wire899  &  n_n228 ) | ( n_n53  &  wire899  &  n_n256 ) ;
 assign wire20900 = ( n_n145  &  n_n53 ) | ( n_n53  &  n_n144 ) | ( n_n53  &  n_n71 ) ;
 assign wire20904 = ( wire634 ) | ( wire20898 ) | ( wire20900 ) ;
 assign wire20905 = ( n_n2272 ) | ( n_n952 ) | ( n_n560 ) | ( wire20899 ) ;
 assign wire20907 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n144 ) | ( n_n4  &  n_n226 ) ;
 assign wire20908 = ( wire409 ) | ( wire546 ) | ( wire19443 ) | ( wire20907 ) ;
 assign wire20909 = ( wire5681 ) | ( wire5682 ) | ( wire5683 ) | ( wire19442 ) ;
 assign wire20912 = ( n_n3382 ) | ( n_n3383 ) | ( wire20908 ) | ( wire20909 ) ;
 assign wire20913 = ( n_n3364 ) | ( n_n3386 ) | ( n_n3385 ) | ( wire20895 ) ;
 assign wire20914 = ( n_n3362 ) | ( wire20819 ) | ( wire20912 ) ;
 assign wire20917 = ( n_n229  &  n_n165  &  n_n284 ) | ( n_n283  &  n_n165  &  n_n284 ) ;
 assign wire20919 = ( wire3946 ) | ( wire758 ) ;
 assign wire20920 = ( n_n5693 ) | ( wire452 ) | ( wire5441 ) | ( wire5442 ) ;
 assign wire20923 = ( wire48 ) | ( n_n110 ) | ( n_n108 ) | ( wire103 ) ;
 assign wire20924 = ( wire3943 ) | ( n_n132  &  wire299 ) | ( n_n132  &  wire20923 ) ;
 assign wire20925 = ( n_n3  &  n_n66 ) | ( n_n4  &  n_n148 ) ;
 assign wire20926 = ( n_n3  &  wire160 ) | ( n_n3  &  n_n14 ) | ( n_n3  &  n_n252 ) ;
 assign wire20928 = ( wire184 ) | ( wire72 ) | ( n_n258  &  wire905 ) ;
 assign wire20931 = ( n_n2618 ) | ( n_n3757 ) | ( wire739 ) | ( wire3931 ) ;
 assign wire20933 = ( n_n4  &  n_n95 ) | ( n_n268  &  n_n148 ) ;
 assign wire20934 = ( n_n4  &  wire68 ) | ( n_n3  &  wire68 ) ;
 assign wire20936 = ( wire3924 ) | ( n_n3  &  wire1940 ) ;
 assign wire20938 = ( n_n1  &  n_n108 ) | ( n_n2  &  wire82 ) ;
 assign wire20942 = ( n_n1  &  wire1027 ) | ( n_n2  &  wire1026 ) ;
 assign wire20944 = ( n_n3155 ) | ( n_n3519 ) | ( n_n3520 ) | ( wire20942 ) ;
 assign wire20946 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n258  &  wire905 ) ;
 assign wire20947 = ( n_n3  &  n_n226 ) | ( n_n3  &  n_n281  &  wire908 ) ;
 assign wire20950 = ( n_n5  &  n_n66 ) | ( n_n5  &  n_n228  &  wire912 ) ;
 assign wire20952 = ( n_n6  &  n_n226 ) | ( n_n6  &  n_n281  &  wire908 ) ;
 assign wire20955 = ( n_n4605 ) | ( wire20952 ) | ( n_n5  &  wire208 ) ;
 assign wire20956 = ( n_n4815 ) | ( n_n4816 ) | ( wire3896 ) ;
 assign wire20958 = ( wire55 ) | ( wire453 ) | ( n_n256  &  wire914 ) ;
 assign wire20959 = ( n_n1  &  n_n111 ) | ( n_n1  &  n_n38 ) | ( n_n1  &  wire453 ) ;
 assign wire20962 = ( n_n3260 ) | ( n_n3772 ) | ( wire395 ) | ( wire5219 ) ;
 assign wire20964 = ( n_n3255 ) | ( n_n2  &  wire1899 ) ;
 assign wire20967 = ( n_n1  &  n_n95 ) | ( n_n2  &  wire68 ) ;
 assign wire20968 = ( wire20967 ) | ( n_n2  &  wire1871 ) ;
 assign wire20971 = ( n_n3162 ) | ( wire496 ) | ( wire806 ) | ( wire20968 ) ;
 assign wire20973 = ( n_n4  &  n_n31 ) | ( n_n147  &  n_n94 ) ;
 assign wire20974 = ( n_n94  &  n_n88 ) | ( n_n94  &  n_n258  &  wire914 ) ;
 assign wire20975 = ( n_n11  &  n_n94 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  n_n39 ) ;
 assign wire20980 = ( n_n109 ) | ( n_n77 ) | ( wire49 ) | ( wire143 ) ;
 assign wire20981 = ( n_n227  &  n_n28 ) | ( n_n94  &  n_n41 ) ;
 assign wire20982 = ( n_n145  &  n_n5 ) | ( n_n227  &  n_n70 ) ;
 assign wire20984 = ( wire20981 ) | ( wire20982 ) | ( wire278  &  wire1018 ) ;
 assign wire20987 = ( wire333 ) | ( n_n2986 ) | ( wire712 ) ;
 assign wire20988 = ( n_n3  &  n_n66 ) | ( n_n4  &  n_n9 ) ;
 assign wire20989 = ( n_n4  &  n_n61 ) | ( n_n3  &  n_n15 ) ;
 assign wire20993 = ( wire409 ) | ( wire476 ) | ( wire446 ) | ( wire20988 ) ;
 assign wire20994 = ( n_n2982 ) | ( wire20989 ) | ( n_n3  &  wire1914 ) ;
 assign wire20996 = ( wire876 ) | ( wire20993 ) | ( wire20994 ) ;
 assign wire20998 = ( n_n48  &  n_n15 ) | ( n_n53  &  n_n148 ) ;
 assign wire20999 = ( n_n53  &  n_n108 ) | ( n_n48  &  wire82 ) ;
 assign wire21003 = ( wire463 ) | ( wire3860 ) | ( n_n48  &  wire1938 ) ;
 assign wire21004 = ( n_n4160 ) | ( wire20998 ) | ( n_n48  &  wire1192 ) ;
 assign wire21006 = ( n_n48  &  n_n226 ) | ( n_n48  &  n_n281  &  wire908 ) ;
 assign wire21009 = ( (~ i_15_)  &  n_n279  &  n_n247 ) | ( i_15_  &  n_n247  &  n_n225 ) ;
 assign wire21010 = ( wire457 ) | ( n_n53  &  n_n228  &  wire902 ) ;
 assign wire21013 = ( n_n3791 ) | ( n_n48  &  n_n147 ) | ( n_n48  &  n_n148 ) ;
 assign wire21014 = ( wire461 ) | ( wire3843 ) | ( wire21010 ) ;
 assign wire21017 = ( n_n5  &  n_n41 ) | ( n_n5  &  n_n113 ) | ( n_n5  &  wire102 ) ;
 assign wire21019 = ( n_n4636 ) | ( wire3837 ) | ( wire21017 ) ;
 assign wire21021 = ( n_n54  &  n_n6 ) | ( n_n48  &  n_n148 ) ;
 assign wire21022 = ( n_n48  &  n_n220  &  wire914 ) | ( n_n48  &  n_n256  &  wire914 ) ;
 assign wire21023 = ( n_n54  &  n_n5 ) | ( n_n48  &  n_n147 ) ;
 assign wire21027 = ( wire389 ) | ( wire464 ) | ( wire463 ) | ( wire21021 ) ;
 assign wire21028 = ( wire21022 ) | ( wire21023 ) | ( n_n5  &  wire1928 ) ;
 assign wire21030 = ( n_n5  &  wire67 ) | ( n_n6  &  wire69 ) ;
 assign wire21034 = ( n_n4624 ) | ( n_n4633 ) | ( n_n5  &  wire1939 ) ;
 assign wire21035 = ( wire727 ) | ( n_n4632 ) | ( wire487 ) | ( wire21030 ) ;
 assign wire21038 = ( n_n1555 ) | ( n_n48  &  wire1917 ) ;
 assign wire21042 = ( n_n56  &  n_n226 ) | ( n_n57  &  n_n148 ) ;
 assign wire21043 = ( wire3821 ) | ( n_n56  &  wire160 ) ;
 assign wire21046 = ( wire5031 ) | ( wire21043 ) | ( n_n56  &  n_n60 ) ;
 assign wire21047 = ( n_n4892 ) | ( wire4056 ) | ( wire20826 ) | ( wire21042 ) ;
 assign wire21049 = ( n_n48  &  n_n220  &  wire914 ) | ( n_n48  &  n_n256  &  wire914 ) ;
 assign wire21051 = ( wire461 ) | ( wire464 ) | ( wire21049 ) ;
 assign wire21054 = ( wire681 ) | ( wire298 ) | ( wire521 ) | ( wire21051 ) ;
 assign wire21057 = ( n_n3587 ) | ( wire478 ) | ( wire20344 ) ;
 assign wire21059 = ( n_n3827 ) | ( n_n1433 ) | ( wire406 ) | ( wire20343 ) ;
 assign wire21061 = ( wire770 ) | ( wire771 ) | ( wire21057 ) | ( wire21059 ) ;
 assign wire21063 = ( n_n3124 ) | ( n_n3123 ) | ( wire21061 ) ;
 assign wire21065 = ( n_n57  &  n_n108 ) | ( n_n56  &  wire82 ) ;
 assign wire21066 = ( n_n57  &  wire44 ) | ( n_n57  &  n_n11 ) | ( n_n57  &  wire95 ) ;
 assign wire21069 = ( n_n56  &  wire1897 ) | ( n_n56  &  wire1898 ) ;
 assign wire21070 = ( n_n4920 ) | ( n_n4907 ) | ( wire21066 ) ;
 assign wire21072 = ( n_n56  &  n_n29 ) | ( n_n56  &  wire49 ) | ( n_n56  &  wire88 ) ;
 assign wire21073 = ( n_n4923 ) | ( n_n4924 ) | ( wire5544 ) ;
 assign wire21074 = ( n_n4922 ) | ( n_n4921 ) | ( wire21072 ) ;
 assign wire21076 = ( n_n57  &  n_n95 ) | ( n_n145  &  n_n94 ) ;
 assign wire21077 = ( n_n56  &  wire68 ) | ( n_n57  &  wire55 ) ;
 assign wire21081 = ( n_n4675 ) | ( n_n4676 ) | ( n_n4686 ) | ( wire21076 ) ;
 assign wire21083 = ( n_n100  &  n_n226 ) | ( n_n94  &  wire208 ) ;
 assign wire21085 = ( n_n94  &  n_n246 ) | ( n_n94  &  n_n228  &  wire912 ) ;
 assign wire21089 = ( wire780 ) | ( wire654 ) | ( wire3791 ) | ( wire21085 ) ;
 assign wire21090 = ( n_n3864 ) | ( n_n2724 ) | ( wire3790 ) ;
 assign wire21092 = ( n_n197  &  n_n94 ) | ( n_n100  &  wire83 ) ;
 assign wire21093 = ( wire21092 ) | ( n_n94  &  wire1910 ) ;
 assign wire21095 = ( n_n2926 ) | ( wire4117 ) | ( wire20772 ) | ( wire21093 ) ;
 assign wire21098 = ( n_n94  &  n_n41 ) | ( n_n94  &  wire77 ) | ( n_n94  &  n_n86 ) ;
 assign wire21101 = ( n_n1066 ) | ( n_n1645 ) | ( wire3778 ) ;
 assign wire21103 = ( wire67 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21105 = ( n_n31  &  n_n100 ) | ( n_n100  &  wire1855 ) | ( n_n100  &  wire1896 ) ;
 assign wire21108 = ( n_n255  &  n_n197 ) | ( n_n189  &  n_n109 ) ;
 assign wire21109 = ( n_n189  &  n_n279  &  wire914 ) | ( n_n189  &  n_n279  &  wire904 ) ;
 assign wire21110 = ( n_n54  &  n_n100 ) | ( n_n189  &  n_n101 ) ;
 assign wire21113 = ( n_n54  &  n_n94 ) | ( n_n100  &  wire77 ) ;
 assign wire21114 = ( wire21113 ) | ( n_n94  &  wire1943 ) ;
 assign wire21116 = ( n_n3722 ) | ( n_n3221 ) | ( wire21114 ) ;
 assign wire21118 = ( wire460 ) | ( wire20193 ) | ( n_n111  &  n_n57 ) ;
 assign wire21120 = ( wire553 ) | ( wire653 ) | ( wire21118 ) ;
 assign wire21122 = ( n_n3129 ) | ( n_n3130 ) | ( wire21120 ) ;
 assign wire21125 = ( wire411 ) | ( n_n5  &  n_n197 ) | ( n_n5  &  wire1926 ) ;
 assign wire21127 = ( n_n2882 ) | ( wire4694 ) | ( wire4695 ) | ( wire21125 ) ;
 assign wire21129 = ( n_n3118 ) | ( n_n3117 ) | ( wire21127 ) ;
 assign wire21131 = ( n_n3096 ) | ( n_n3097 ) | ( wire21129 ) ;
 assign wire21134 = ( n_n29 ) | ( n_n26 ) | ( wire80 ) | ( wire88 ) ;
 assign wire21135 = ( n_n111 ) | ( wire49 ) | ( n_n101 ) | ( wire61 ) ;
 assign wire21136 = ( wire640 ) | ( wire485 ) | ( n_n3  &  n_n76 ) ;
 assign wire21138 = ( wire55 ) | ( wire453 ) | ( n_n256  &  wire914 ) ;
 assign wire21141 = ( wire82 ) | ( wire42 ) | ( n_n279  &  wire899 ) ;
 assign wire21142 = ( n_n70 ) | ( n_n20 ) | ( wire79 ) | ( wire66 ) ;
 assign wire21143 = ( n_n4  &  n_n108 ) | ( n_n3  &  n_n15 ) ;
 assign wire21146 = ( n_n3506 ) | ( n_n3229 ) | ( wire742 ) | ( wire21143 ) ;
 assign wire21148 = ( n_n7354 ) | ( wire3745 ) | ( wire4302 ) | ( wire21146 ) ;
 assign wire21151 = ( n_n3727 ) | ( wire3736 ) | ( n_n4  &  n_n9 ) ;
 assign wire21153 = ( n_n3140 ) | ( n_n3138 ) | ( wire21151 ) ;
 assign wire21154 = ( n_n3110 ) | ( n_n3109 ) | ( wire20944 ) | ( wire21153 ) ;
 assign wire21157 = ( n_n110  &  n_n122 ) | ( n_n111  &  n_n122 ) | ( n_n122  &  wire54 ) ;
 assign wire21159 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire21160 = ( n_n5682 ) | ( wire21159 ) | ( n_n121  &  n_n111 ) ;
 assign wire21163 = ( n_n4489 ) | ( wire3733 ) | ( wire21157 ) | ( wire21160 ) ;
 assign wire21164 = ( n_n5769 ) | ( wire48  &  n_n132 ) ;
 assign wire21165 = ( wire364 ) | ( n_n124  &  wire48 ) | ( wire48  &  n_n122 ) ;
 assign wire21168 = ( wire21164 ) | ( wire21165 ) | ( wire1845  &  wire1842 ) ;
 assign wire21169 = ( wire535 ) | ( n_n118  &  n_n260  &  n_n155 ) ;
 assign wire21170 = ( wire777 ) | ( n_n5675 ) | ( wire4928 ) | ( wire19999 ) ;
 assign wire21173 = ( n_n2772 ) | ( wire879 ) | ( wire21169 ) | ( wire21170 ) ;
 assign wire21174 = ( wire3725 ) | ( wire3726 ) | ( wire21163 ) | ( wire21173 ) ;
 assign wire21175 = ( wire394 ) | ( n_n139  &  wire911  &  n_n281 ) ;
 assign wire21178 = ( n_n4476 ) | ( n_n4477 ) | ( wire3712 ) | ( wire21175 ) ;
 assign wire21180 = ( n_n4  &  n_n108 ) | ( n_n48  &  n_n148 ) ;
 assign wire21182 = ( wire21180 ) | ( n_n4  &  n_n223 ) | ( n_n4  &  wire42 ) ;
 assign wire21183 = ( wire640 ) | ( wire455 ) | ( wire485 ) ;
 assign wire21186 = ( wire867 ) | ( wire378 ) | ( wire21182 ) | ( wire21183 ) ;
 assign wire21188 = ( n_n4  &  n_n8 ) | ( n_n4  &  n_n281  &  wire908 ) ;
 assign wire21190 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n258  &  wire905 ) ;
 assign wire21191 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n7 ) | ( n_n4  &  n_n144 ) ;
 assign wire21193 = ( n_n4  &  n_n148 ) | ( n_n4  &  wire901  &  n_n228 ) ;
 assign wire21195 = ( n_n4  &  n_n64 ) | ( n_n4  &  n_n281  &  wire906 ) ;
 assign wire21196 = ( n_n3  &  n_n15 ) | ( n_n3  &  n_n281  &  wire904 ) ;
 assign wire21197 = ( n_n3  &  n_n14 ) | ( n_n3  &  n_n252 ) | ( n_n3  &  wire83 ) ;
 assign wire21200 = ( wire546 ) | ( wire3688 ) | ( wire21195 ) ;
 assign wire21201 = ( wire3689 ) | ( wire21196 ) | ( wire21197 ) ;
 assign wire21203 = ( wire69 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21204 = ( n_n78 ) | ( n_n203 ) | ( wire80 ) | ( wire20149 ) ;
 assign wire21206 = ( n_n4  &  n_n197 ) | ( n_n3  &  n_n216 ) ;
 assign wire21208 = ( wire333 ) | ( n_n2986 ) | ( wire21206 ) ;
 assign wire21211 = ( n_n203 ) | ( n_n68 ) | ( wire514 ) | ( wire20149 ) ;
 assign wire21212 = ( wire62 ) | ( n_n216 ) | ( n_n16 ) | ( wire20155 ) ;
 assign wire21213 = ( wire62 ) | ( wire899  &  n_n258 ) ;
 assign wire21214 = ( n_n221 ) | ( n_n20 ) | ( wire79 ) | ( wire469 ) ;
 assign wire21215 = ( n_n16 ) | ( n_n72 ) | ( wire66 ) | ( wire20155 ) ;
 assign wire21217 = ( n_n25 ) | ( n_n23 ) | ( wire74 ) | ( wire19457 ) ;
 assign wire21218 = ( wire88 ) | ( n_n222  &  wire902 ) | ( wire902  &  n_n258 ) ;
 assign wire21220 = ( wire716 ) | ( wire3674 ) | ( wire3682 ) | ( wire21208 ) ;
 assign wire21221 = ( wire519 ) | ( wire3673 ) | ( wire3680 ) | ( wire3681 ) ;
 assign wire21223 = ( n_n113 ) | ( n_n85 ) | ( wire102 ) | ( wire87 ) ;
 assign wire21224 = ( wire67 ) | ( wire368 ) | ( n_n88 ) | ( n_n103 ) ;
 assign wire21225 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n31 ) | ( n_n4  &  n_n26 ) ;
 assign wire21228 = ( n_n1341 ) | ( n_n1346 ) | ( wire21225 ) ;
 assign wire21230 = ( wire89 ) | ( wire901  &  n_n222 ) | ( wire901  &  n_n258 ) ;
 assign wire21231 = ( n_n34 ) | ( n_n82 ) | ( wire47 ) | ( wire86 ) ;
 assign wire21232 = ( wire67 ) | ( wire87 ) | ( wire914  &  n_n225 ) ;
 assign wire21233 = ( wire476 ) | ( wire3662 ) | ( n_n3  &  wire1914 ) ;
 assign wire21234 = ( wire3653 ) | ( n_n4  &  wire1439 ) ;
 assign wire21236 = ( n_n1359 ) | ( wire4470 ) | ( wire21233 ) | ( wire21234 ) ;
 assign wire21238 = ( n_n4  &  n_n61 ) | ( n_n4  &  n_n228  &  wire902 ) ;
 assign wire21240 = ( wire3642 ) | ( n_n4  &  n_n10 ) | ( n_n4  &  wire113 ) ;
 assign wire21243 = ( n_n4005 ) | ( n_n3930 ) | ( wire21238 ) | ( wire21240 ) ;
 assign wire21245 = ( n_n3929 ) | ( n_n3406 ) | ( n_n3904 ) | ( wire21243 ) ;
 assign wire21247 = ( n_n171 ) | ( n_n24 ) | ( wire53 ) | ( wire19407 ) ;
 assign wire21248 = ( n_n53  &  n_n257 ) | ( n_n268  &  wire56 ) ;
 assign wire21250 = ( n_n4068 ) | ( n_n4069 ) | ( wire21248 ) ;
 assign wire21252 = ( n_n4  &  n_n257 ) | ( n_n4  &  n_n228  &  wire902 ) ;
 assign wire21253 = ( n_n4  &  n_n145 ) | ( n_n3  &  n_n14 ) ;
 assign wire21257 = ( wire349 ) | ( wire546 ) | ( wire634 ) | ( wire19400 ) ;
 assign wire21258 = ( n_n4076 ) | ( wire483 ) | ( wire21252 ) | ( wire21253 ) ;
 assign wire21260 = ( n_n4  &  n_n226 ) | ( n_n4  &  n_n281  &  wire908 ) ;
 assign wire21261 = ( n_n4  &  n_n144 ) | ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) ;
 assign wire21263 = ( wire557 ) | ( wire21260 ) | ( wire21261 ) ;
 assign wire21264 = ( n_n1440 ) | ( wire5758 ) | ( wire19391 ) | ( wire21263 ) ;
 assign wire21266 = ( wire913  &  n_n258 ) | ( n_n220  &  wire912 ) ;
 assign wire21268 = ( n_n265  &  n_n62 ) | ( n_n268  &  n_n148 ) ;
 assign wire21269 = ( n_n106  &  n_n265 ) | ( n_n4  &  n_n54 ) ;
 assign wire21271 = ( n_n281  &  wire913 ) | ( n_n220  &  wire914 ) ;
 assign wire21272 = ( wire21271 ) | ( wire50 ) ;
 assign wire21273 = ( n_n38 ) | ( n_n39 ) | ( wire245 ) | ( wire453 ) ;
 assign wire21274 = ( n_n179 ) | ( n_n206 ) | ( wire57 ) | ( wire20107 ) ;
 assign wire21276 = ( wire3627 ) | ( wire3629 ) | ( wire21268 ) | ( wire21269 ) ;
 assign wire21277 = ( wire60 ) | ( wire19738 ) | ( wire913  &  n_n256 ) ;
 assign wire21278 = ( n_n204 ) | ( n_n112 ) | ( wire52 ) | ( wire84 ) ;
 assign wire21279 = ( wire85 ) | ( wire64 ) | ( n_n279  &  wire907 ) ;
 assign wire21280 = ( wire89 ) | ( n_n81 ) | ( n_n83 ) | ( wire86 ) ;
 assign wire21281 = ( n_n268  &  wire913  &  n_n220 ) | ( n_n268  &  wire903  &  n_n220 ) ;
 assign wire21284 = ( n_n97 ) | ( n_n51 ) | ( wire71 ) | ( wire19575 ) ;
 assign wire21285 = ( wire51 ) | ( wire19578 ) | ( n_n222  &  wire906 ) ;
 assign wire21286 = ( n_n46 ) | ( n_n43 ) | ( wire59 ) | ( wire19577 ) ;
 assign wire21288 = ( n_n896 ) | ( n_n1363 ) | ( n_n4  &  n_n105 ) ;
 assign wire21290 = ( wire3612 ) | ( wire3613 ) | ( wire21288 ) ;
 assign wire21293 = ( n_n3898 ) | ( n_n3897 ) | ( n_n3896 ) ;
 assign wire21296 = ( wire71 ) | ( wire96 ) | ( wire898  &  n_n256 ) ;
 assign wire21297 = ( n_n92 ) | ( wire19578 ) | ( wire900  &  n_n258 ) ;
 assign wire21298 = ( n_n57  &  n_n54 ) | ( n_n177  &  n_n112 ) ;
 assign wire21299 = ( n_n189  &  n_n109 ) | ( n_n177  &  n_n35 ) ;
 assign wire21302 = ( wire21299 ) | ( wire21298 ) ;
 assign wire21303 = ( wire372 ) | ( wire894 ) | ( wire386 ) | ( wire484 ) ;
 assign wire21306 = ( wire89 ) | ( wire901  &  n_n222 ) | ( wire901  &  n_n258 ) ;
 assign wire21307 = ( n_n34 ) | ( n_n82 ) | ( wire47 ) | ( wire86 ) ;
 assign wire21309 = ( n_n113 ) | ( n_n85 ) | ( wire102 ) | ( wire87 ) ;
 assign wire21310 = ( wire67 ) | ( wire368 ) | ( n_n41 ) | ( n_n88 ) ;
 assign wire21313 = ( n_n92 ) | ( wire19578 ) | ( wire900  &  n_n258 ) ;
 assign wire21314 = ( n_n46 ) | ( n_n43 ) | ( wire59 ) | ( wire19577 ) ;
 assign wire21315 = ( wire51 ) | ( wire71 ) | ( wire898  &  n_n256 ) ;
 assign wire21316 = ( n_n43 ) | ( n_n51 ) | ( wire59 ) | ( wire19575 ) ;
 assign wire21318 = ( n_n1604 ) | ( n_n57  &  wire21313 ) | ( n_n57  &  wire21314 ) ;
 assign wire21322 = ( n_n203 ) | ( wire20149 ) | ( wire911  &  n_n258 ) ;
 assign wire21323 = ( n_n16 ) | ( n_n68 ) | ( wire514 ) | ( wire20155 ) ;
 assign wire21328 = ( wire101 ) | ( wire95 ) | ( n_n228  &  wire912 ) ;
 assign wire21329 = ( n_n57  &  n_n11 ) | ( n_n57  &  n_n148 ) | ( n_n57  &  wire95 ) ;
 assign wire21330 = ( wire21329 ) | ( n_n57  &  wire1807 ) ;
 assign wire21332 = ( wire65 ) | ( wire902  &  n_n258 ) | ( wire902  &  n_n225 ) ;
 assign wire21333 = ( n_n80 ) | ( n_n78 ) | ( wire80 ) | ( wire88 ) ;
 assign wire21334 = ( wire40 ) | ( wire79 ) | ( wire899  &  n_n256 ) ;
 assign wire21335 = ( n_n221 ) | ( n_n23 ) | ( wire469 ) | ( wire74 ) ;
 assign wire21337 = ( n_n1584 ) | ( n_n56  &  wire21332 ) | ( n_n56  &  wire21333 ) ;
 assign wire21339 = ( n_n113 ) | ( n_n85 ) | ( wire102 ) | ( wire87 ) ;
 assign wire21340 = ( wire67 ) | ( wire368 ) | ( n_n41 ) | ( n_n88 ) ;
 assign wire21341 = ( wire78 ) | ( wire902  &  n_n258 ) ;
 assign wire21342 = ( n_n37 ) | ( wire89 ) | ( n_n80 ) | ( wire88 ) ;
 assign wire21343 = ( n_n34 ) | ( n_n82 ) | ( wire47 ) | ( wire86 ) ;
 assign wire21345 = ( wire40 ) | ( wire19457 ) | ( n_n222  &  wire897 ) ;
 assign wire21346 = ( n_n200 ) | ( n_n23 ) | ( wire74 ) | ( wire104 ) ;
 assign wire21347 = ( n_n103 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21348 = ( n_n78 ) | ( n_n25 ) | ( wire80 ) | ( wire19457 ) ;
 assign wire21350 = ( n_n1591 ) | ( n_n56  &  wire21345 ) | ( n_n56  &  wire21346 ) ;
 assign wire21352 = ( wire3562 ) | ( wire3563 ) | ( wire3565 ) | ( wire21337 ) ;
 assign wire21353 = ( wire79 ) | ( wire83 ) | ( wire899  &  n_n256 ) ;
 assign wire21354 = ( n_n65 ) | ( n_n221 ) | ( wire469 ) | ( wire73 ) ;
 assign wire21356 = ( wire635 ) | ( wire3550 ) | ( wire3584 ) | ( wire3585 ) ;
 assign wire21359 = ( n_n2433 ) | ( n_n2431 ) | ( wire3551 ) | ( wire21356 ) ;
 assign wire21362 = ( wire3544 ) | ( n_n57  &  wire899  &  n_n228 ) ;
 assign wire21364 = ( n_n2440 ) | ( wire21362 ) | ( n_n56  &  wire955 ) ;
 assign wire21365 = ( n_n2429 ) | ( n_n2428 ) | ( wire21359 ) | ( wire21364 ) ;
 assign wire21367 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign wire21370 = ( wire69 ) | ( wire80 ) | ( n_n279  &  wire908 ) ;
 assign wire21371 = ( wire40 ) | ( n_n30 ) | ( n_n74 ) | ( wire21367 ) ;
 assign wire21372 = ( n_n4  &  wire988 ) | ( n_n4  &  n_n279  &  wire899 ) ;
 assign wire21374 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n30 ) | ( n_n4  &  n_n26 ) ;
 assign wire21377 = ( n_n85 ) | ( wire54 ) | ( n_n279  &  wire912 ) ;
 assign wire21379 = ( n_n281  &  wire913 ) | ( n_n220  &  wire914 ) ;
 assign wire21381 = ( n_n4  &  n_n186 ) | ( n_n268  &  n_n148 ) ;
 assign wire21383 = ( i_15_  &  n_n242  &  n_n279 ) | ( (~ i_15_)  &  n_n242  &  n_n279 ) | ( i_15_  &  n_n279  &  n_n247 ) | ( (~ i_15_)  &  n_n279  &  n_n247 ) ;
 assign wire21384 = ( n_n73 ) | ( n_n67 ) | ( wire19408 ) | ( wire19738 ) ;
 assign wire21385 = ( n_n268  &  n_n110 ) | ( n_n265  &  n_n32 ) ;
 assign wire21387 = ( wire3520 ) | ( wire21385 ) | ( n_n268  &  n_n22 ) ;
 assign wire21389 = ( (~ i_14_)  &  i_13_  &  i_12_  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire21390 = ( n_n3  &  wire51 ) | ( n_n4  &  n_n93 ) ;
 assign wire21391 = ( wire71 ) | ( n_n279  &  wire900 ) | ( n_n279  &  wire904 ) ;
 assign wire21393 = ( n_n102 ) | ( n_n85 ) | ( wire54 ) | ( wire71 ) ;
 assign wire21394 = ( wire476 ) | ( n_n3  &  wire149 ) | ( n_n3  &  wire21391 ) ;
 assign wire21396 = ( n_n2104 ) | ( wire3530 ) | ( wire3531 ) | ( wire21394 ) ;
 assign wire21402 = ( wire119 ) | ( wire281 ) | ( wire858 ) ;
 assign wire21403 = ( n_n1  &  n_n145 ) | ( n_n1  &  wire1030 ) | ( n_n2  &  wire1030 ) ;
 assign wire21404 = ( n_n268  &  wire264 ) | ( n_n2  &  wire1031 ) ;
 assign wire21408 = ( wire21403 ) | ( wire21404 ) | ( n_n12  &  wire135 ) ;
 assign wire21409 = ( wire3500 ) | ( wire3499 ) ;
 assign wire21414 = ( wire268 ) | ( wire119 ) | ( wire858 ) ;
 assign wire21415 = ( wire3496 ) | ( n_n1  &  wire1102 ) ;
 assign wire21416 = ( wire3507 ) | ( wire3508 ) | ( wire21408 ) | ( wire21409 ) ;
 assign wire21417 = ( n_n53  &  n_n281  &  wire905 ) | ( n_n53  &  n_n281  &  wire908 ) ;
 assign wire21424 = ( wire153 ) | ( wire255 ) | ( wire436 ) ;
 assign wire21425 = ( n_n4  &  n_n108 ) | ( n_n4  &  n_n93 ) | ( n_n4  &  n_n70 ) ;
 assign wire21426 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n66 ) ;
 assign wire21427 = ( n_n4  &  n_n223 ) | ( n_n4  &  n_n281  &  wire908 ) ;
 assign wire21428 = ( n_n4  &  n_n145 ) | ( n_n4  &  n_n76 ) | ( n_n4  &  n_n26 ) ;
 assign wire21431 = ( wire476 ) | ( wire21426 ) | ( wire21428 ) ;
 assign wire21432 = ( wire3480 ) | ( wire21427 ) | ( n_n4  &  wire1161 ) ;
 assign wire21434 = ( n_n53  &  wire899  &  n_n281 ) | ( n_n53  &  n_n281  &  wire902 ) ;
 assign wire21435 = ( n_n2  &  wire78 ) | ( n_n2  &  n_n281  &  wire907 ) ;
 assign wire21438 = ( n_n2274 ) | ( wire3469 ) | ( wire21434 ) ;
 assign wire21440 = ( n_n2126 ) | ( wire3470 ) | ( wire21435 ) | ( wire21438 ) ;
 assign wire21442 = ( n_n111  &  n_n57 ) | ( n_n56  &  n_n95 ) ;
 assign wire21443 = ( n_n56  &  wire252 ) | ( n_n57  &  wire329 ) ;
 assign wire21445 = ( n_n100  &  n_n281  &  wire905 ) | ( n_n94  &  n_n281  &  wire905 ) ;
 assign wire21446 = ( n_n151  &  wire168 ) | ( n_n57  &  wire482 ) ;
 assign wire21448 = ( n_n57  &  n_n95 ) | ( n_n56  &  n_n42 ) ;
 assign wire21449 = ( n_n57  &  n_n42 ) | ( n_n57  &  wire1379 ) | ( n_n56  &  wire1379 ) ;
 assign wire21453 = ( n_n4674 ) | ( n_n4682 ) | ( wire3451 ) | ( wire21448 ) ;
 assign wire21455 = ( n_n100  &  n_n12 ) | ( n_n100  &  n_n66 ) | ( n_n12  &  n_n94 ) ;
 assign wire21457 = ( n_n281  &  wire904 ) | ( n_n281  &  wire907 ) ;
 assign wire21458 = ( n_n281  &  wire914 ) | ( n_n281  &  wire908 ) ;
 assign wire21459 = ( n_n100  &  n_n281  &  wire908 ) | ( n_n100  &  n_n281  &  wire907 ) ;
 assign wire21462 = ( n_n2398 ) | ( wire3441 ) | ( wire3442 ) | ( wire21459 ) ;
 assign wire21463 = ( wire3440 ) | ( wire3447 ) | ( wire21455 ) ;
 assign wire21464 = ( wire329 ) | ( wire453 ) | ( n_n256  &  wire914 ) ;
 assign wire21466 = ( n_n111  &  n_n56 ) | ( n_n57  &  n_n32 ) | ( n_n56  &  n_n32 ) ;
 assign wire21467 = ( n_n57  &  n_n81 ) | ( n_n57  &  wire1383 ) | ( n_n57  &  wire86 ) ;
 assign wire21470 = ( n_n2169 ) | ( wire3432 ) | ( wire21466 ) | ( wire21467 ) ;
 assign wire21474 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire897 ) ;
 assign wire21477 = ( wire327 ) | ( wire235 ) | ( wire21474 ) ;
 assign wire21478 = ( n_n94  &  n_n200 ) | ( n_n94  &  wire911  &  n_n281 ) ;
 assign wire21479 = ( wire21478 ) | ( n_n100  &  wire1413 ) ;
 assign wire21482 = ( n_n100  &  n_n279  &  wire901 ) | ( n_n100  &  n_n279  &  wire907 ) ;
 assign wire21483 = ( n_n100  &  n_n32 ) | ( n_n100  &  wire901  &  n_n281 ) ;
 assign wire21486 = ( n_n57  &  n_n76 ) | ( n_n57  &  n_n26 ) | ( n_n57  &  wire80 ) ;
 assign wire21487 = ( n_n110  &  n_n57 ) | ( n_n57  &  n_n67 ) | ( n_n57  &  wire19738 ) ;
 assign wire21488 = ( n_n110  &  n_n56 ) | ( n_n57  &  n_n108 ) ;
 assign wire21490 = ( n_n56  &  n_n108 ) | ( n_n57  &  n_n148 ) ;
 assign wire21491 = ( n_n106  &  n_n57 ) | ( n_n106  &  n_n56 ) | ( n_n57  &  wire1096 ) ;
 assign wire21493 = ( n_n4916 ) | ( wire3409 ) | ( wire21488 ) | ( wire21491 ) ;
 assign wire21494 = ( wire3402 ) | ( wire3413 ) | ( wire21487 ) | ( wire21490 ) ;
 assign wire21497 = ( n_n186  &  n_n53 ) | ( n_n7  &  wire191 ) ;
 assign wire21499 = ( wire3393 ) | ( wire3400 ) | ( wire3401 ) | ( wire21497 ) ;
 assign wire21500 = ( n_n56  &  n_n76 ) | ( n_n57  &  n_n22 ) ;
 assign wire21501 = ( n_n56  &  wire369 ) | ( n_n56  &  wire903  &  n_n220 ) ;
 assign wire21505 = ( n_n4920 ) | ( n_n4924 ) | ( wire693 ) | ( wire21500 ) ;
 assign wire21506 = ( wire3382 ) | ( wire3416 ) | ( wire21486 ) | ( wire21501 ) ;
 assign wire21507 = ( wire21506 ) | ( wire21505 ) ;
 assign wire21508 = ( n_n2158 ) | ( wire21493 ) | ( wire21494 ) | ( wire21499 ) ;
 assign wire21512 = ( n_n2180 ) | ( wire3375 ) | ( wire3376 ) ;
 assign wire21514 = ( n_n2097 ) | ( wire3428 ) | ( wire21479 ) | ( wire21512 ) ;
 assign wire21516 = ( n_n4  &  n_n281  &  wire904 ) | ( n_n3  &  n_n281  &  wire904 ) ;
 assign wire21517 = ( n_n4  &  n_n12 ) | ( n_n3  &  n_n12 ) | ( n_n3  &  wire83 ) ;
 assign wire21521 = ( n_n4  &  n_n281  &  wire914 ) | ( n_n4  &  n_n281  &  wire908 ) ;
 assign wire21522 = ( n_n4  &  n_n281  &  wire903 ) | ( n_n4  &  n_n281  &  wire905 ) ;
 assign wire21525 = ( wire3360 ) | ( wire3361 ) | ( wire21521 ) | ( wire21522 ) ;
 assign wire21529 = ( n_n6  &  n_n12 ) | ( n_n5  &  n_n12 ) | ( n_n6  &  n_n66 ) | ( n_n5  &  n_n66 ) ;
 assign wire21530 = ( n_n6  &  n_n281  &  wire905 ) | ( n_n6  &  n_n281  &  wire908 ) ;
 assign wire21531 = ( n_n5  &  n_n60 ) | ( n_n6  &  wire985 ) | ( n_n5  &  wire985 ) ;
 assign wire21533 = ( wire21530 ) | ( wire21531 ) | ( n_n106  &  wire164 ) ;
 assign wire21536 = ( n_n279  &  wire913 ) | ( n_n279  &  wire897 ) ;
 assign wire21537 = ( n_n145  &  n_n5 ) | ( n_n207  &  n_n67 ) ;
 assign wire21538 = ( n_n151  &  wire164 ) | ( n_n227  &  wire1156 ) ;
 assign wire21540 = ( n_n94  &  n_n200 ) | ( n_n227  &  n_n70 ) ;
 assign wire21541 = ( n_n94  &  n_n204 ) | ( n_n227  &  n_n109 ) ;
 assign wire21544 = ( n_n110  &  n_n94 ) | ( n_n4  &  n_n30 ) ;
 assign wire21545 = ( n_n100  &  n_n279  &  wire901 ) | ( n_n100  &  n_n279  &  wire907 ) ;
 assign wire21546 = ( n_n106  &  n_n100 ) | ( n_n100  &  n_n33 ) | ( n_n100  &  n_n81 ) ;
 assign wire21549 = ( wire3324 ) | ( wire21544 ) | ( wire21545 ) | ( wire21546 ) ;
 assign wire21551 = ( n_n279  &  wire899 ) | ( n_n279  &  wire897 ) ;
 assign wire21554 = ( wire69 ) | ( wire80 ) | ( n_n279  &  wire908 ) ;
 assign wire21555 = ( wire40 ) | ( n_n30 ) | ( n_n74 ) | ( wire21367 ) ;
 assign wire21557 = ( n_n2137 ) | ( wire3320 ) | ( n_n6  &  wire1486 ) ;
 assign wire21560 = ( n_n53  &  n_n281  &  wire905 ) | ( n_n53  &  n_n281  &  wire908 ) ;
 assign wire21561 = ( n_n48  &  n_n281  &  wire914 ) | ( n_n53  &  n_n281  &  wire914 ) ;
 assign wire21562 = ( n_n48  &  n_n60 ) | ( n_n48  &  n_n7 ) | ( n_n53  &  n_n7 ) ;
 assign wire21565 = ( n_n106  &  n_n53 ) | ( n_n48  &  n_n148 ) ;
 assign wire21566 = ( n_n186  &  n_n6 ) | ( n_n48  &  n_n135 ) ;
 assign wire21569 = ( n_n145  &  n_n48 ) | ( n_n53  &  n_n280 ) ;
 assign wire21572 = ( wire376 ) | ( wire3296 ) | ( wire3297 ) | ( wire21569 ) ;
 assign wire21574 = ( n_n6  &  wire69 ) | ( n_n5  &  n_n171 ) ;
 assign wire21576 = ( n_n279  &  wire901 ) | ( n_n279  &  wire912 ) ;
 assign wire21578 = ( n_n85 ) | ( n_n35 ) | ( wire54 ) | ( wire86 ) ;
 assign wire21579 = ( n_n111  &  n_n6 ) | ( n_n6  &  n_n38 ) | ( n_n6  &  wire78 ) ;
 assign wire21583 = ( wire77 ) | ( wire71 ) | ( n_n279  &  wire904 ) ;
 assign wire21584 = ( n_n279  &  wire900 ) | ( n_n279  &  wire912 ) ;
 assign wire21586 = ( n_n85 ) | ( n_n90 ) | ( wire54 ) | ( wire21389 ) ;
 assign wire21588 = ( n_n2145 ) | ( wire3282 ) | ( wire3283 ) ;
 assign wire21590 = ( n_n111  &  n_n48 ) | ( n_n48  &  n_n171 ) | ( n_n48  &  n_n38 ) ;
 assign wire21593 = ( n_n53  &  n_n280 ) | ( n_n53  &  n_n33 ) | ( n_n53  &  n_n35 ) ;
 assign wire21596 = ( n_n279  &  wire901 ) | ( n_n279  &  wire912 ) ;
 assign wire21599 = ( wire78 ) | ( wire71 ) | ( n_n279  &  wire904 ) ;
 assign wire21600 = ( n_n84 ) | ( wire77 ) | ( n_n35 ) | ( wire86 ) ;
 assign wire21603 = ( n_n48  &  n_n12 ) | ( n_n53  &  n_n12 ) | ( n_n53  &  n_n66 ) ;
 assign wire21605 = ( wire456 ) | ( n_n53  &  n_n107 ) | ( n_n53  &  n_n19 ) ;
 assign wire21608 = ( wire80 ) | ( n_n279  &  wire902 ) | ( n_n279  &  wire908 ) ;
 assign wire21609 = ( n_n279  &  wire899 ) | ( n_n279  &  wire897 ) ;
 assign wire21612 = ( n_n2154 ) | ( wire621 ) | ( wire3255 ) | ( wire3256 ) ;
 assign wire21614 = ( n_n151  &  n_n4 ) | ( n_n151  &  n_n3 ) | ( n_n3  &  n_n145 ) ;
 assign wire21615 = ( n_n2101 ) | ( wire3538 ) | ( wire21372 ) | ( wire21614 ) ;
 assign wire21616 = ( n_n2099 ) | ( n_n2100 ) | ( wire21525 ) | ( wire21615 ) ;
 assign wire21620 = ( n_n2060 ) | ( wire21415 ) | ( wire21416 ) | ( wire21616 ) ;
 assign wire21621 = ( n_n2062 ) | ( n_n2063 ) | ( n_n2064 ) | ( n_n2065 ) ;
 assign wire21624 = ( n_n108 ) | ( wire103 ) | ( (~ i_9_)  &  (~ i_10_) ) ;
 assign wire21626 = ( i_7_  &  i_6_  &  n_n118  &  n_n284 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n284 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n284 ) ;
 assign wire21627 = ( i_7_  &  i_6_  &  n_n284  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n284  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n284  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n284  &  n_n116 ) ;
 assign wire21628 = ( n_n5769 ) | ( n_n5660 ) | ( n_n151  &  n_n126 ) ;
 assign wire21631 = ( wire3232 ) | ( wire21626 ) | ( wire21627 ) | ( wire21628 ) ;
 assign wire21633 = ( n_n4  &  n_n80 ) | ( n_n4  &  n_n29 ) | ( n_n4  &  wire61 ) ;
 assign wire21635 = ( n_n4  &  n_n76 ) | ( n_n4  &  n_n25 ) | ( n_n4  &  n_n27 ) ;
 assign wire21636 = ( wire154 ) | ( wire361 ) | ( wire901  &  n_n256 ) ;
 assign wire21637 = ( wire226 ) | ( wire362 ) | ( wire898  &  n_n256 ) ;
 assign wire21639 = ( wire87 ) | ( wire362 ) | ( n_n220  &  wire914 ) ;
 assign wire21640 = ( n_n42 ) | ( wire59 ) | ( wire243 ) | ( wire428 ) ;
 assign wire21642 = ( wire236 ) | ( wire230 ) | ( wire902  &  n_n256 ) ;
 assign wire21643 = ( n_n111 ) | ( n_n22 ) | ( wire74 ) | ( wire87 ) ;
 assign wire21646 = ( n_n34 ) | ( n_n22 ) | ( wire154 ) | ( wire74 ) ;
 assign wire21647 = ( n_n78 ) | ( wire236 ) | ( wire230 ) | ( wire424 ) ;
 assign wire21648 = ( wire3215 ) | ( n_n1  &  wire21646 ) | ( n_n1  &  wire21647 ) ;
 assign wire21649 = ( wire3219 ) | ( wire3220 ) | ( wire3221 ) | ( wire3222 ) ;
 assign wire21650 = ( wire901  &  n_n220 ) | ( wire898  &  n_n220 ) ;
 assign wire21651 = ( n_n1  &  n_n64 ) | ( n_n2  &  n_n64 ) | ( n_n1  &  wire1451 ) ;
 assign wire21652 = ( n_n2  &  n_n144 ) | ( n_n268  &  n_n22 ) ;
 assign wire21655 = ( n_n2  &  wire1772 ) | ( n_n1  &  wire1771 ) | ( n_n2  &  wire1771 ) ;
 assign wire21657 = ( wire3203 ) | ( wire3211 ) | ( wire21651 ) | ( wire21655 ) ;
 assign wire21658 = ( wire911  &  n_n220 ) | ( n_n220  &  wire914 ) ;
 assign wire21660 = ( n_n265  &  n_n32 ) | ( n_n268  &  wire273 ) ;
 assign wire21662 = ( n_n268  &  n_n110 ) | ( n_n265  &  n_n62 ) ;
 assign wire21663 = ( n_n3  &  n_n47 ) | ( n_n268  &  n_n147 ) ;
 assign wire21665 = ( wire21662 ) | ( wire21663 ) | ( n_n268  &  wire247 ) ;
 assign wire21666 = ( wire3190 ) | ( n_n4  &  wire1812 ) ;
 assign wire21668 = ( (~ i_15_)  &  n_n222  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) ;
 assign wire21670 = ( wire690 ) | ( wire3178 ) | ( n_n4  &  n_n47 ) ;
 assign wire21671 = ( wire3179 ) | ( wire3213 ) | ( wire3214 ) ;
 assign wire21673 = ( wire3186 ) | ( wire3187 ) | ( wire21670 ) | ( wire21671 ) ;
 assign wire21675 = ( n_n4  &  n_n64 ) | ( n_n53  &  n_n27 ) ;
 assign wire21676 = ( n_n53  &  n_n76 ) | ( n_n3  &  n_n14 ) ;
 assign wire21677 = ( n_n4  &  n_n144 ) | ( n_n53  &  n_n78 ) ;
 assign wire21678 = ( n_n53  &  n_n80 ) | ( n_n53  &  n_n28 ) | ( n_n53  &  n_n29 ) ;
 assign wire21681 = ( n_n4  &  n_n8 ) | ( n_n4  &  n_n222  &  wire900 ) ;
 assign wire21683 = ( wire690 ) | ( wire622 ) | ( wire21681 ) ;
 assign wire21686 = ( n_n94  &  n_n203 ) | ( n_n94  &  wire913  &  n_n220 ) ;
 assign wire21687 = ( n_n94  &  n_n58 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  n_n39 ) ;
 assign wire21690 = ( n_n147  &  n_n94 ) | ( n_n4  &  n_n80 ) ;
 assign wire21691 = ( n_n4  &  n_n221 ) | ( n_n94  &  n_n150 ) ;
 assign wire21694 = ( n_n227  &  n_n28 ) | ( n_n94  &  n_n199 ) ;
 assign wire21695 = ( n_n227  &  wire143 ) | ( n_n207  &  wire1794 ) ;
 assign wire21697 = ( wire657 ) | ( wire21694 ) | ( wire21695 ) ;
 assign wire21699 = ( n_n53  &  wire899  &  n_n281 ) | ( n_n53  &  wire899  &  n_n256 ) ;
 assign wire21700 = ( n_n53  &  n_n8 ) | ( n_n53  &  n_n222  &  wire899 ) ;
 assign wire21701 = ( n_n53  &  wire899  &  n_n220 ) | ( n_n53  &  n_n220  &  wire905 ) ;
 assign wire21702 = ( n_n2  &  n_n37 ) | ( n_n53  &  wire1849 ) ;
 assign wire21705 = ( wire154 ) | ( wire64 ) | ( n_n222  &  wire907 ) ;
 assign wire21706 = ( wire59 ) | ( wire243 ) | ( n_n220  &  wire906 ) ;
 assign wire21709 = ( wire932 ) | ( n_n1752 ) | ( wire3120 ) | ( wire3121 ) ;
 assign wire21711 = ( n_n1703 ) | ( n_n1704 ) | ( wire21709 ) ;
 assign wire21713 = ( n_n56  &  n_n22 ) | ( n_n57  &  wire426 ) ;
 assign wire21714 = ( n_n57  &  wire212 ) | ( n_n56  &  wire212 ) ;
 assign wire21715 = ( i_15_  &  n_n242  &  n_n222 ) | ( (~ i_15_)  &  n_n242  &  n_n222 ) | ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) ;
 assign wire21716 = ( n_n57  &  wire903  &  n_n220 ) | ( n_n57  &  n_n220  &  wire905 ) ;
 assign wire21718 = ( wire21716 ) | ( n_n56  &  n_n76 ) | ( n_n56  &  wire165 ) ;
 assign wire21719 = ( wire3109 ) | ( n_n56  &  wire247 ) | ( n_n56  &  wire21715 ) ;
 assign wire21721 = ( n_n56  &  n_n108 ) | ( n_n57  &  wire1198 ) ;
 assign wire21723 = ( n_n57  &  wire271 ) | ( n_n56  &  wire472 ) ;
 assign wire21724 = ( n_n110  &  n_n57 ) | ( n_n110  &  n_n56 ) | ( n_n57  &  wire247 ) ;
 assign wire21726 = ( n_n57  &  wire1249 ) | ( n_n57  &  wire1248 ) | ( n_n56  &  wire1248 ) ;
 assign wire21728 = ( wire3098 ) | ( wire3106 ) | ( wire21721 ) | ( wire21726 ) ;
 assign wire21729 = ( n_n111  &  n_n56 ) | ( n_n57  &  n_n76 ) ;
 assign wire21730 = ( n_n56  &  wire426 ) | ( n_n57  &  wire379 ) ;
 assign wire21732 = ( n_n57  &  n_n220  &  wire914 ) | ( n_n57  &  n_n220  &  wire907 ) ;
 assign wire21733 = ( n_n56  &  n_n32 ) | ( n_n57  &  wire158 ) ;
 assign wire21735 = ( n_n57  &  wire200 ) | ( n_n56  &  wire273 ) ;
 assign wire21737 = ( wire21732 ) | ( wire21735 ) | ( n_n56  &  wire200 ) ;
 assign wire21739 = ( n_n1792 ) | ( wire3080 ) | ( wire21733 ) | ( wire21737 ) ;
 assign wire21741 = ( n_n56  &  n_n95 ) | ( n_n57  &  wire429 ) ;
 assign wire21742 = ( n_n56  &  wire99 ) | ( n_n57  &  wire273 ) ;
 assign wire21743 = ( n_n57  &  n_n99 ) | ( n_n94  &  n_n8 ) ;
 assign wire21744 = ( n_n57  &  n_n52 ) | ( wire168  &  wire1195 ) ;
 assign wire21746 = ( wire901  &  n_n220 ) | ( wire898  &  n_n220 ) ;
 assign wire21748 = ( wire898  &  n_n220 ) | ( n_n220  &  wire912 ) ;
 assign wire21749 = ( wire901  &  n_n220 ) | ( wire902  &  n_n220 ) ;
 assign wire21751 = ( n_n147  &  n_n94 ) | ( n_n100  &  n_n64 ) | ( n_n94  &  n_n64 ) ;
 assign wire21752 = ( wire3072 ) | ( wire21743 ) | ( wire21744 ) | ( wire21751 ) ;
 assign wire21753 = ( n_n100  &  wire1597 ) | ( n_n94  &  wire1596 ) ;
 assign wire21756 = ( n_n94  &  wire911  &  n_n281 ) | ( n_n94  &  wire911  &  n_n256 ) ;
 assign wire21757 = ( n_n110  &  n_n94 ) | ( n_n94  &  n_n203 ) | ( n_n94  &  n_n68 ) ;
 assign wire21759 = ( wire3056 ) | ( wire21756 ) | ( wire21757 ) ;
 assign wire21760 = ( wire3065 ) | ( n_n100  &  wire1599 ) | ( n_n100  &  wire1730 ) ;
 assign wire21761 = ( n_n57  &  n_n95 ) | ( n_n56  &  n_n42 ) ;
 assign wire21762 = ( n_n57  &  wire494 ) | ( n_n57  &  n_n220  &  wire906 ) ;
 assign wire21764 = ( n_n57  &  wire99 ) | ( n_n57  &  wire180 ) ;
 assign wire21766 = ( wire21761 ) | ( wire21764 ) | ( n_n56  &  wire180 ) ;
 assign wire21767 = ( wire3045 ) | ( wire21741 ) | ( wire21742 ) | ( wire21762 ) ;
 assign wire21769 = ( wire21752 ) | ( wire21753 ) | ( wire21759 ) | ( wire21760 ) ;
 assign wire21770 = ( n_n48  &  n_n147 ) | ( n_n53  &  n_n8 ) ;
 assign wire21771 = ( n_n53  &  n_n147 ) | ( n_n48  &  n_n62 ) | ( n_n53  &  n_n62 ) ;
 assign wire21772 = ( n_n48  &  n_n64 ) | ( n_n53  &  n_n64 ) | ( n_n48  &  wire1330 ) ;
 assign wire21775 = ( n_n203 ) | ( wire195 ) | ( wire898  &  n_n220 ) ;
 assign wire21777 = ( n_n69 ) | ( wire84 ) | ( wire375 ) ;
 assign wire21778 = ( n_n221 ) | ( n_n71 ) | ( wire143 ) | ( wire195 ) ;
 assign wire21780 = ( n_n53  &  n_n32 ) | ( n_n53  &  wire901  &  n_n281 ) ;
 assign wire21781 = ( n_n48  &  n_n88 ) | ( n_n48  &  n_n220  &  wire914 ) ;
 assign wire21783 = ( wire21780 ) | ( n_n48  &  wire102 ) ;
 assign wire21784 = ( wire629 ) | ( wire21781 ) | ( n_n53  &  n_n34 ) ;
 assign wire21785 = ( wire901  &  n_n225 ) | ( n_n220  &  wire897 ) ;
 assign wire21786 = ( n_n53  &  n_n37 ) | ( n_n48  &  n_n144 ) ;
 assign wire21789 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire898 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire898 ) ;
 assign wire21790 = ( n_n5  &  n_n47 ) | ( n_n6  &  n_n95 ) ;
 assign wire21792 = ( wire631 ) | ( wire3012 ) | ( wire21790 ) ;
 assign wire21794 = ( i_15_  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n267 ) ;
 assign wire21797 = ( wire807 ) | ( wire270 ) | ( n_n222  &  wire904 ) ;
 assign wire21798 = ( n_n99 ) | ( n_n44 ) | ( wire226 ) | ( wire21668 ) ;
 assign wire21799 = ( wire3043 ) | ( n_n6  &  wire1329 ) | ( n_n6  &  wire1630 ) ;
 assign wire21804 = ( n_n69 ) | ( wire84 ) | ( wire230 ) ;
 assign wire21805 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire899 ) ;
 assign wire21807 = ( n_n71 ) | ( n_n69 ) | ( wire143 ) | ( wire84 ) ;
 assign wire21808 = ( wire3003 ) | ( wire3004 ) | ( n_n6  &  n_n108 ) ;
 assign wire21811 = ( n_n6  &  wire1290 ) | ( n_n6  &  wire1289 ) | ( n_n5  &  wire1289 ) ;
 assign wire21813 = ( n_n5  &  n_n8 ) | ( n_n6  &  n_n58 ) ;
 assign wire21814 = ( n_n80  &  n_n227 ) | ( n_n144  &  wire1776 ) ;
 assign wire21815 = ( wire164  &  n_n150 ) | ( n_n207  &  wire425 ) ;
 assign wire21817 = ( wire21811 ) | ( wire21815 ) | ( n_n5  &  wire1291 ) ;
 assign wire21820 = ( wire102 ) | ( wire263 ) | ( wire912  &  n_n256 ) ;
 assign wire21821 = ( wire901  &  n_n222 ) | ( n_n222  &  wire902 ) ;
 assign wire21823 = ( n_n29 ) | ( n_n83 ) | ( wire61 ) | ( wire64 ) ;
 assign wire21825 = ( n_n1765 ) | ( wire2981 ) | ( wire2982 ) ;
 assign wire21827 = ( n_n53  &  wire901  &  n_n222 ) | ( n_n53  &  wire901  &  n_n281 ) ;
 assign wire21828 = ( n_n53  &  n_n32 ) | ( n_n48  &  n_n88 ) ;
 assign wire21832 = ( n_n48  &  n_n47 ) | ( n_n57  &  n_n150 ) ;
 assign wire21834 = ( i_15_  &  n_n222  &  n_n247 ) | ( i_15_  &  n_n222  &  n_n267 ) ;
 assign wire21837 = ( wire807 ) | ( wire270 ) | ( n_n222  &  wire904 ) ;
 assign wire21838 = ( n_n99 ) | ( n_n44 ) | ( wire226 ) | ( wire21668 ) ;
 assign wire21842 = ( n_n53  &  n_n76 ) | ( n_n53  &  n_n25 ) | ( n_n53  &  n_n27 ) ;
 assign wire21844 = ( n_n53  &  n_n221 ) | ( n_n53  &  n_n220  &  wire905 ) ;
 assign wire21845 = ( n_n53  &  n_n107 ) | ( n_n53  &  n_n20 ) | ( n_n53  &  wire1803 ) ;
 assign wire21847 = ( wire2952 ) | ( wire21844 ) | ( wire21845 ) ;
 assign wire21849 = ( n_n111  &  n_n48 ) | ( n_n53  &  n_n80 ) ;
 assign wire21850 = ( n_n48  &  n_n281  &  wire912 ) | ( n_n48  &  wire912  &  n_n256 ) ;
 assign wire21853 = ( wire2942 ) | ( wire2943 ) | ( wire21849 ) | ( wire21850 ) ;
 assign wire21855 = ( n_n1781 ) | ( wire2973 ) | ( wire2974 ) | ( wire21853 ) ;
 assign wire21857 = ( n_n94  &  wire425 ) | ( n_n94  &  n_n222  &  wire903 ) ;
 assign wire21859 = ( i_7_  &  i_6_  &  n_n118  &  n_n260 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n260 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n260 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n260 ) ;
 assign wire21860 = ( i_7_  &  i_6_  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n260  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n260  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n260  &  n_n116 ) ;
 assign wire21861 = ( wire21859 ) | ( n_n142  &  wire1593 ) ;
 assign wire21862 = ( wire503 ) | ( wire21860 ) | ( wire48  &  n_n152 ) ;
 assign wire21864 = ( wire2929 ) | ( wire893 ) ;
 assign wire21865 = ( n_n4477 ) | ( wire21861 ) | ( wire21862 ) ;
 assign wire21866 = ( wire59 ) | ( wire243 ) | ( n_n220  &  wire906 ) ;
 assign wire21867 = ( wire87 ) | ( wire428 ) | ( n_n220  &  wire914 ) ;
 assign wire21868 = ( wire59 ) | ( wire243 ) | ( n_n220  &  wire906 ) ;
 assign wire21869 = ( wire362 ) | ( wire361 ) ;
 assign wire21872 = ( n_n94  &  wire912  &  n_n256 ) | ( n_n94  &  wire912  &  n_n225 ) ;
 assign wire21874 = ( wire667 ) | ( wire2919 ) | ( wire21872 ) ;
 assign wire21877 = ( n_n1804 ) | ( wire2920 ) | ( wire2927 ) | ( wire2928 ) ;
 assign wire21881 = ( n_n1690 ) | ( n_n1691 ) | ( n_n1688 ) | ( n_n1687 ) ;
 assign wire21884 = ( n_n4  &  n_n108 ) | ( n_n4  &  n_n107 ) | ( n_n4  &  n_n221 ) ;
 assign wire21885 = ( wire2917 ) | ( wire2918 ) | ( wire21884 ) ;
 assign wire21888 = ( n_n4  &  wire900  &  n_n220 ) | ( n_n4  &  wire902  &  n_n220 ) ;
 assign wire21889 = ( n_n4  &  n_n147 ) | ( n_n3  &  n_n14 ) ;
 assign wire21892 = ( wire898  &  n_n220 ) | ( n_n220  &  wire897 ) ;
 assign wire21893 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire899 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire899 ) ;
 assign wire21895 = ( wire143 ) | ( wire21893 ) | ( wire899  &  n_n225 ) ;
 assign wire21896 = ( n_n4  &  n_n144 ) | ( n_n4  &  n_n150 ) | ( n_n3  &  n_n150 ) ;
 assign wire21900 = ( wire2893 ) | ( n_n4  &  wire957 ) ;
 assign wire21902 = ( n_n1729 ) | ( wire3228 ) | ( wire21633 ) | ( wire21900 ) ;
 assign wire21904 = ( n_n1694 ) | ( n_n1693 ) | ( wire21902 ) ;
 assign wire21907 = ( n_n133 ) | ( wire62 ) | ( n_n112 ) | ( wire84 ) ;
 assign wire21910 = ( wire333 ) | ( wire664 ) | ( wire485 ) | ( wire3762 ) ;
 assign wire21912 = ( n_n4  &  n_n252 ) | ( n_n3  &  wire83 ) ;
 assign wire21913 = ( wire903  &  n_n258 ) | ( wire901  &  n_n220 ) ;
 assign wire21914 = ( n_n4  &  n_n8 ) | ( n_n4  &  n_n61 ) | ( n_n4  &  n_n62 ) ;
 assign wire21918 = ( n_n4  &  n_n257 ) | ( n_n4  &  wire899  &  n_n220 ) ;
 assign wire21920 = ( wire2874 ) | ( wire21918 ) | ( n_n3  &  wire1112 ) ;
 assign wire21922 = ( n_n3  &  n_n252 ) | ( n_n3  &  wire898  &  n_n220 ) ;
 assign wire21923 = ( n_n4  &  n_n64 ) | ( n_n3  &  n_n64 ) | ( n_n4  &  n_n13 ) | ( n_n3  &  n_n13 ) ;
 assign wire21925 = ( wire2864 ) | ( wire21922 ) | ( wire21923 ) ;
 assign wire21926 = ( n_n1320 ) | ( wire2883 ) | ( wire2885 ) | ( wire21912 ) ;
 assign wire21927 = ( n_n1157 ) | ( wire21920 ) | ( wire21925 ) ;
 assign wire21928 = ( wire2888 ) | ( wire2889 ) | ( wire21910 ) | ( wire21926 ) ;
 assign wire21929 = ( wire67 ) | ( n_n135 ) | ( n_n39 ) | ( wire245 ) ;
 assign wire21930 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire902 ) | ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  wire902 ) ;
 assign wire21933 = ( n_n4  &  n_n31 ) | ( n_n4  &  n_n80 ) | ( n_n4  &  n_n26 ) ;
 assign wire21935 = ( n_n1341 ) | ( n_n1346 ) | ( wire21933 ) ;
 assign wire21938 = ( n_n82 ) | ( wire47 ) | ( n_n220  &  wire907 ) ;
 assign wire21939 = ( wire85 ) | ( wire437 ) | ( n_n228  &  wire907 ) ;
 assign wire21941 = ( n_n3242 ) | ( wire476 ) | ( n_n1356 ) | ( wire3662 ) ;
 assign wire21943 = ( wire124 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21944 = ( wire212 ) | ( wire49 ) | ( n_n228  &  wire908 ) ;
 assign wire21946 = ( wire2845 ) | ( wire519 ) ;
 assign wire21948 = ( n_n3731 ) | ( n_n1339 ) | ( wire2846 ) | ( wire21946 ) ;
 assign wire21950 = ( n_n1108 ) | ( n_n1109 ) | ( wire21948 ) ;
 assign wire21953 = ( wire112 ) | ( wire65 ) | ( wire902  &  n_n225 ) ;
 assign wire21954 = ( wire200 ) | ( n_n79 ) | ( wire78 ) | ( wire49 ) ;
 assign wire21956 = ( n_n1412 ) | ( n_n2  &  wire990 ) | ( n_n2  &  wire93 ) ;
 assign wire21958 = ( wire99 ) | ( n_n220  &  wire904 ) | ( n_n256  &  wire904 ) ;
 assign wire21959 = ( wire41 ) | ( wire47 ) | ( wire901  &  n_n225 ) ;
 assign wire21960 = ( wire85 ) | ( wire437 ) | ( n_n228  &  wire907 ) ;
 assign wire21962 = ( n_n1  &  wire1052 ) | ( n_n1  &  n_n39 ) | ( n_n1  &  wire245 ) ;
 assign wire21963 = ( i_14_  &  i_13_  &  i_12_  &  wire903 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire903 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire903 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire903 ) ;
 assign wire21965 = ( wire40 ) | ( n_n281  &  wire897 ) | ( n_n258  &  wire897 ) ;
 assign wire21966 = ( wire431 ) | ( wire346 ) ;
 assign wire21968 = ( n_n3768 ) | ( n_n3770 ) | ( n_n2  &  wire1424 ) ;
 assign wire21969 = ( wire21968 ) | ( n_n1  &  wire21965 ) | ( n_n1  &  wire21966 ) ;
 assign wire21970 = ( wire2839 ) | ( wire2842 ) | ( wire21956 ) | ( wire21962 ) ;
 assign wire21971 = ( (~ i_15_)  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n220 ) ;
 assign wire21973 = ( n_n2  &  n_n257 ) | ( n_n268  &  wire56 ) ;
 assign wire21975 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire21977 = ( (~ i_15_)  &  n_n253  &  n_n258 ) | ( i_15_  &  n_n253  &  n_n220 ) ;
 assign wire21979 = ( wire514 ) | ( wire325 ) | ( wire911  &  n_n225 ) ;
 assign wire21980 = ( wire60 ) | ( n_n18 ) | ( wire73 ) | ( wire21977 ) ;
 assign wire21981 = ( n_n3523 ) | ( n_n2  &  wire1514 ) ;
 assign wire21982 = ( i_14_  &  i_13_  &  i_12_  &  wire905 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire905 ) | ( i_14_  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  wire905 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire905 ) ;
 assign wire21983 = ( n_n216 ) | ( wire84 ) | ( n_n279  &  wire913 ) ;
 assign wire21984 = ( n_n133 ) | ( wire62 ) | ( n_n28 ) | ( wire65 ) ;
 assign wire21985 = ( wire431 ) | ( wire343 ) ;
 assign wire21987 = ( n_n3255 ) | ( n_n1  &  wire100 ) | ( n_n1  &  wire21982 ) ;
 assign wire21988 = ( n_n1  &  n_n10 ) | ( n_n2  &  n_n10 ) | ( n_n2  &  n_n62 ) ;
 assign wire21991 = ( wire2813 ) | ( wire2814 ) | ( wire2830 ) | ( wire2831 ) ;
 assign wire21992 = ( wire2827 ) | ( wire21973 ) | ( wire21988 ) | ( wire21991 ) ;
 assign wire21993 = ( wire2822 ) | ( wire2825 ) | ( wire21981 ) | ( wire21987 ) ;
 assign wire21995 = ( n_n82 ) | ( n_n36 ) | ( wire85 ) | ( wire47 ) ;
 assign wire21997 = ( n_n133 ) | ( wire62 ) | ( n_n112 ) | ( wire84 ) ;
 assign wire21998 = ( wire40 ) | ( wire343 ) | ( wire911  &  n_n258 ) ;
 assign wire21999 = ( wire823 ) | ( n_n265  &  wire437 ) | ( n_n265  &  wire21995 ) ;
 assign wire22000 = ( n_n4  &  wire68 ) | ( n_n265  &  n_n62 ) ;
 assign wire22001 = ( wire903  &  n_n258 ) | ( wire911  &  n_n220 ) ;
 assign wire22002 = ( n_n220  &  wire914 ) | ( n_n256  &  wire914 ) | ( n_n220  &  wire897 ) ;
 assign wire22004 = ( wire57 ) | ( wire22002 ) | ( n_n279  &  wire914 ) ;
 assign wire22005 = ( n_n268  &  n_n240 ) | ( n_n265  &  n_n10 ) ;
 assign wire22007 = ( n_n1370 ) | ( wire22005 ) | ( n_n268  &  wire273 ) ;
 assign wire22009 = ( wire51 ) | ( n_n44 ) | ( n_n90 ) | ( wire19385 ) ;
 assign wire22010 = ( n_n4  &  n_n105 ) | ( n_n4  &  n_n47 ) | ( n_n4  &  n_n46 ) ;
 assign wire22012 = ( n_n1359 ) | ( n_n1363 ) | ( wire22010 ) ;
 assign wire22014 = ( n_n1173 ) | ( wire2790 ) | ( wire22012 ) ;
 assign wire22016 = ( wire165 ) | ( wire514 ) | ( wire911  &  n_n225 ) ;
 assign wire22017 = ( wire60 ) | ( wire325 ) | ( wire913  &  n_n228 ) ;
 assign wire22020 = ( n_n4834 ) | ( wire411 ) | ( wire2784 ) ;
 assign wire22022 = ( n_n6  &  wire75 ) | ( n_n207  &  n_n103 ) ;
 assign wire22024 = ( (~ i_15_)  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign wire22026 = ( wire83 ) | ( wire274 ) | ( wire899  &  n_n281 ) ;
 assign wire22029 = ( n_n112 ) | ( n_n246 ) | ( wire73 ) | ( wire52 ) ;
 assign wire22033 = ( (~ i_15_)  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n220 ) ;
 assign wire22034 = ( n_n53  &  n_n257 ) | ( n_n2  &  wire85 ) ;
 assign wire22035 = ( n_n53  &  wire899  &  n_n281 ) | ( n_n53  &  wire899  &  n_n220 ) ;
 assign wire22039 = ( n_n1  &  wire41 ) | ( n_n2  &  wire1171 ) ;
 assign wire22040 = ( wire456 ) | ( wire626 ) | ( wire591 ) | ( wire932 ) ;
 assign wire22041 = ( n_n1433 ) | ( wire22035 ) | ( wire22039 ) ;
 assign wire22043 = ( n_n4  &  n_n258  &  wire906 ) | ( n_n4  &  n_n258  &  wire908 ) ;
 assign wire22044 = ( n_n4  &  wire899  &  n_n220 ) | ( n_n4  &  wire902  &  n_n220 ) ;
 assign wire22047 = ( n_n4  &  n_n64 ) | ( n_n4  &  n_n258  &  wire905 ) ;
 assign wire22048 = ( n_n53  &  n_n222  &  wire899 ) | ( n_n53  &  wire899  &  n_n258 ) ;
 assign wire22050 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n80 ) | ( n_n53  &  wire42 ) ;
 assign wire22052 = ( n_n53  &  n_n27 ) | ( n_n53  &  wire140 ) | ( n_n53  &  wire61 ) ;
 assign wire22053 = ( wire409 ) | ( wire479 ) | ( wire22050 ) ;
 assign wire22054 = ( wire22047 ) | ( wire22048 ) | ( wire22052 ) ;
 assign wire22058 = ( wire300 ) | ( wire19578 ) | ( n_n222  &  wire906 ) ;
 assign wire22059 = ( wire99 ) | ( wire81 ) | ( n_n46 ) | ( wire77 ) ;
 assign wire22061 = ( n_n3778 ) | ( n_n2  &  wire1387 ) | ( n_n2  &  wire43 ) ;
 assign wire22064 = ( n_n4  &  n_n222  &  wire899 ) | ( n_n4  &  wire899  &  n_n258 ) ;
 assign wire22066 = ( n_n10  &  n_n100 ) | ( n_n94  &  n_n39 ) ;
 assign wire22067 = ( n_n94  &  n_n150 ) | ( n_n94  &  n_n258  &  wire914 ) ;
 assign wire22070 = ( n_n147  &  n_n94 ) | ( n_n100  &  n_n81 ) ;
 assign wire22071 = ( n_n110  &  n_n94 ) | ( n_n100  &  n_n104 ) ;
 assign wire22075 = ( wire696 ) | ( wire548 ) | ( wire374 ) | ( wire434 ) ;
 assign wire22076 = ( wire799 ) | ( wire22070 ) | ( wire22071 ) ;
 assign wire22079 = ( n_n207  &  n_n257 ) | ( n_n227  &  n_n70 ) ;
 assign wire22081 = ( n_n227  &  n_n28 ) | ( n_n94  &  n_n203 ) ;
 assign wire22082 = ( n_n94  &  n_n279  &  wire903 ) | ( n_n94  &  n_n222  &  wire903 ) ;
 assign wire22083 = ( n_n227  &  n_n257 ) | ( n_n207  &  wire232 ) ;
 assign wire22084 = ( wire40  &  n_n94 ) | ( n_n94  &  n_n24 ) | ( n_n94  &  n_n74 ) ;
 assign wire22087 = ( wire22081 ) | ( wire22082 ) | ( wire22084 ) ;
 assign wire22088 = ( wire2725 ) | ( wire2726 ) | ( wire22083 ) ;
 assign wire22090 = ( n_n4  &  n_n46 ) | ( n_n4  &  wire899  &  n_n281 ) ;
 assign wire22093 = ( n_n1359 ) | ( wire333 ) | ( wire455 ) | ( wire22090 ) ;
 assign wire22095 = ( n_n1173 ) | ( n_n1210 ) | ( wire22093 ) ;
 assign wire22097 = ( wire2709 ) | ( wire2708 ) ;
 assign wire22099 = ( n_n1217 ) | ( wire2774 ) | ( wire2775 ) | ( wire22097 ) ;
 assign wire22101 = ( n_n1127 ) | ( n_n1126 ) | ( wire22099 ) ;
 assign wire22104 = ( wire78 ) | ( wire433 ) | ( wire901  &  n_n281 ) ;
 assign wire22106 = ( wire2703 ) | ( n_n5  &  n_n113 ) | ( n_n5  &  wire102 ) ;
 assign wire22108 = ( wire55 ) | ( wire87 ) | ( n_n228  &  wire914 ) ;
 assign wire22109 = ( wire200 ) | ( wire807 ) | ( n_n279  &  wire904 ) ;
 assign wire22110 = ( wire77 ) | ( wire112 ) | ( n_n281  &  wire898 ) ;
 assign wire22112 = ( n_n4870 ) | ( n_n1497 ) | ( n_n6  &  n_n38 ) ;
 assign wire22115 = ( n_n212 ) | ( n_n200 ) | ( wire56 ) | ( wire104 ) ;
 assign wire22117 = ( n_n4846 ) | ( n_n4852 ) | ( n_n1490 ) ;
 assign wire22119 = ( wire2692 ) | ( wire22117 ) | ( n_n5  &  wire998 ) ;
 assign wire22121 = ( n_n53  &  n_n280 ) | ( n_n48  &  n_n87 ) ;
 assign wire22124 = ( n_n54  &  n_n6 ) | ( n_n53  &  n_n10 ) ;
 assign wire22125 = ( n_n48  &  n_n220  &  wire914 ) | ( n_n48  &  n_n256  &  wire914 ) ;
 assign wire22126 = ( n_n48  &  n_n246 ) | ( n_n48  &  n_n135 ) | ( n_n48  &  n_n86 ) ;
 assign wire22129 = ( wire631 ) | ( wire22124 ) | ( wire22126 ) ;
 assign wire22130 = ( n_n4124 ) | ( wire2676 ) | ( wire22125 ) ;
 assign wire22134 = ( n_n53  &  n_n61 ) | ( n_n53  &  wire902  &  n_n220 ) ;
 assign wire22135 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n246 ) ;
 assign wire22136 = ( n_n48  &  n_n147 ) | ( n_n48  &  n_n62 ) | ( n_n53  &  n_n62 ) ;
 assign wire22139 = ( wire911  &  n_n220 ) | ( n_n228  &  wire907 ) ;
 assign wire22140 = ( n_n53  &  n_n37 ) | ( n_n48  &  wire223 ) ;
 assign wire22142 = ( n_n4153 ) | ( wire2659 ) | ( wire22140 ) ;
 assign wire22145 = ( wire300 ) | ( wire19578 ) | ( n_n222  &  wire906 ) ;
 assign wire22146 = ( wire81 ) | ( wire311 ) | ( n_n228  &  wire906 ) ;
 assign wire22148 = ( wire389 ) | ( n_n1506 ) | ( n_n1505 ) ;
 assign wire22149 = ( wire2652 ) | ( n_n5  &  wire22145 ) | ( n_n5  &  wire22146 ) ;
 assign wire22154 = ( n_n53  &  n_n197 ) | ( n_n53  &  n_n107 ) | ( n_n53  &  n_n221 ) ;
 assign wire22157 = ( wire624 ) | ( wire22154 ) | ( n_n48  &  wire69 ) ;
 assign wire22159 = ( n_n53  &  wire1489 ) | ( n_n48  &  wire1488 ) ;
 assign wire22160 = ( n_n48  &  wire82 ) | ( n_n48  &  n_n228  &  wire905 ) ;
 assign wire22162 = ( (~ i_15_)  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign wire22164 = ( n_n220  &  wire905 ) | ( n_n258  &  wire907 ) ;
 assign wire22167 = ( wire66 ) | ( wire22164 ) | ( n_n222  &  wire905 ) ;
 assign wire22168 = ( n_n107 ) | ( wire73 ) | ( wire187 ) | ( wire220 ) ;
 assign wire22169 = ( n_n3581 ) | ( wire2637 ) | ( wire2640 ) | ( wire22160 ) ;
 assign wire22170 = ( i_15_  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n222  &  n_n270 ) | ( (~ i_15_)  &  n_n228  &  n_n270 ) ;
 assign wire22171 = ( n_n212 ) | ( n_n200 ) | ( wire56 ) | ( wire104 ) ;
 assign wire22174 = ( n_n3827 ) | ( n_n53  &  wire124 ) | ( n_n53  &  wire212 ) ;
 assign wire22176 = ( n_n4168 ) | ( n_n1542 ) | ( wire2631 ) | ( wire22174 ) ;
 assign wire22181 = ( n_n110  &  n_n94 ) | ( n_n133  &  n_n94 ) | ( n_n94  &  n_n203 ) ;
 assign wire22184 = ( n_n1628 ) | ( n_n2732 ) | ( wire2623 ) ;
 assign wire22185 = ( n_n1624 ) | ( wire22181 ) | ( n_n100  &  wire1044 ) ;
 assign wire22187 = ( n_n94  &  n_n199 ) | ( n_n94  &  n_n225  &  wire897 ) ;
 assign wire22188 = ( n_n94  &  n_n200 ) | ( n_n94  &  n_n24 ) | ( n_n94  &  wire1333 ) ;
 assign wire22190 = ( n_n94  &  n_n38 ) | ( n_n94  &  n_n86 ) | ( n_n94  &  wire1334 ) ;
 assign wire22193 = ( n_n1645 ) | ( wire773 ) | ( n_n100  &  wire49 ) ;
 assign wire22195 = ( n_n22 ) | ( wire66 ) | ( wire899  &  n_n256 ) ;
 assign wire22196 = ( wire104 ) | ( wire274 ) | ( n_n279  &  wire903 ) ;
 assign wire22197 = ( wire56 ) | ( wire345 ) | ( n_n228  &  wire903 ) ;
 assign wire22201 = ( n_n1633 ) | ( n_n2738 ) | ( wire2601 ) | ( wire2602 ) ;
 assign wire22203 = ( n_n94  &  n_n246 ) | ( n_n94  &  n_n220  &  wire912 ) ;
 assign wire22206 = ( (~ i_15_)  &  n_n247  &  n_n258 ) | ( i_15_  &  n_n247  &  n_n220 ) ;
 assign wire22208 = ( (~ i_15_)  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign wire22210 = ( wire66 ) | ( wire22208 ) | ( wire899  &  n_n256 ) ;
 assign wire22211 = ( n_n107 ) | ( wire83 ) | ( wire220 ) | ( wire291 ) ;
 assign wire22213 = ( n_n57  &  n_n222  &  wire898 ) | ( n_n57  &  wire898  &  n_n258 ) ;
 assign wire22214 = ( n_n94  &  wire223 ) | ( n_n57  &  wire486 ) ;
 assign wire22217 = ( n_n57  &  n_n50 ) | ( n_n94  &  n_n150 ) ;
 assign wire22219 = ( wire484 ) | ( wire2581 ) | ( wire22217 ) ;
 assign wire22220 = ( wire2583 ) | ( n_n56  &  wire1167 ) ;
 assign wire22227 = ( n_n4960 ) | ( n_n4675 ) | ( n_n4681 ) | ( n_n1604 ) ;
 assign wire22228 = ( n_n4961 ) | ( wire497 ) | ( wire2571 ) | ( wire2572 ) ;
 assign wire22231 = ( n_n100  &  n_n279  &  wire907 ) | ( n_n100  &  n_n256  &  wire907 ) ;
 assign wire22232 = ( n_n94  &  n_n87 ) | ( n_n94  &  n_n41 ) | ( n_n94  &  n_n88 ) ;
 assign wire22236 = ( n_n100  &  n_n36 ) | ( n_n100  &  wire901  &  n_n258 ) ;
 assign wire22238 = ( wire2561 ) | ( wire2560 ) ;
 assign wire22240 = ( n_n255  &  n_n197 ) | ( n_n241  &  n_n104 ) ;
 assign wire22241 = ( n_n189  &  n_n113 ) | ( n_n177  &  n_n35 ) ;
 assign wire22242 = ( n_n241  &  n_n216 ) | ( n_n255  &  n_n41 ) ;
 assign wire22244 = ( wire807 ) | ( wire311 ) | ( n_n279  &  wire904 ) ;
 assign wire22245 = ( wire300 ) | ( wire19578 ) | ( n_n222  &  wire906 ) ;
 assign wire22248 = ( wire81 ) | ( wire55 ) | ( n_n228  &  wire914 ) ;
 assign wire22249 = ( n_n102 ) | ( wire807 ) | ( n_n220  &  wire906 ) ;
 assign wire22250 = ( wire77 ) | ( wire311 ) | ( n_n281  &  wire898 ) ;
 assign wire22253 = ( n_n3881 ) | ( wire784 ) | ( wire2544 ) | ( wire2545 ) ;
 assign wire22255 = ( i_15_  &  n_n253  &  n_n281 ) | ( (~ i_15_)  &  n_n253  &  n_n228 ) ;
 assign wire22257 = ( wire19575 ) | ( wire22255 ) | ( wire898  &  n_n225 ) ;
 assign wire22259 = ( (~ i_15_)  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n220 ) ;
 assign wire22262 = ( wire407 ) | ( wire457 ) | ( n_n57  &  wire75 ) ;
 assign wire22264 = ( wire579 ) | ( wire764 ) | ( wire2534 ) | ( wire22262 ) ;
 assign wire22266 = ( wire514 ) | ( wire325 ) | ( wire911  &  n_n225 ) ;
 assign wire22270 = ( n_n4921 ) | ( n_n4394 ) | ( wire481 ) | ( n_n4915 ) ;
 assign wire22273 = ( (~ i_15_)  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n220  &  n_n267 ) ;
 assign wire22275 = ( wire66 ) | ( wire274 ) | ( wire899  &  n_n256 ) ;
 assign wire22276 = ( n_n107 ) | ( wire83 ) | ( wire220 ) | ( wire22273 ) ;
 assign wire22277 = ( wire2520 ) | ( wire2532 ) | ( wire2533 ) ;
 assign wire22280 = ( n_n53  &  n_n32 ) | ( n_n53  &  wire901  &  n_n281 ) ;
 assign wire22282 = ( n_n53  &  n_n281  &  wire902 ) | ( n_n53  &  wire902  &  n_n258 ) ;
 assign wire22286 = ( wire479 ) | ( wire656 ) | ( wire2507 ) ;
 assign wire22287 = ( wire629 ) | ( wire462 ) | ( wire2508 ) | ( wire22282 ) ;
 assign wire22290 = ( i_15_  &  n_n253  &  n_n281 ) | ( i_15_  &  n_n253  &  n_n256 ) | ( (~ i_15_)  &  n_n253  &  n_n256 ) ;
 assign wire22291 = ( n_n280 ) | ( n_n35 ) | ( wire78 ) | ( wire64 ) ;
 assign wire22294 = ( n_n4174 ) | ( wire516 ) | ( n_n1555 ) ;
 assign wire22298 = ( wire68 ) | ( n_n98 ) | ( n_n51 ) | ( wire19575 ) ;
 assign wire22300 = ( wire2495 ) | ( n_n53  &  n_n44 ) | ( n_n53  &  wire19385 ) ;
 assign wire22302 = ( n_n4179 ) | ( n_n3843 ) | ( wire2496 ) | ( wire22300 ) ;
 assign wire22304 = ( n_n113 ) | ( n_n35 ) | ( wire102 ) | ( wire64 ) ;
 assign wire22305 = ( wire78 ) | ( wire342 ) | ( wire901  &  n_n281 ) ;
 assign wire22308 = ( n_n1597 ) | ( n_n1598 ) | ( wire704 ) ;
 assign wire22309 = ( n_n87 ) | ( n_n24 ) | ( wire55 ) | ( wire19407 ) ;
 assign wire22310 = ( wire102 ) | ( wire342 ) | ( n_n279  &  wire914 ) ;
 assign wire22312 = ( n_n111  &  n_n56 ) | ( n_n57  &  wire49 ) ;
 assign wire22314 = ( wire762 ) | ( n_n1591 ) | ( wire22312 ) ;
 assign wire22315 = ( wire104 ) | ( wire274 ) | ( n_n279  &  wire903 ) ;
 assign wire22316 = ( wire56 ) | ( wire345 ) | ( n_n228  &  wire903 ) ;
 assign wire22317 = ( n_n57  &  n_n22 ) | ( n_n56  &  wire49 ) ;
 assign wire22319 = ( wire2478 ) | ( wire22317 ) ;
 assign wire22321 = ( n_n1584 ) | ( wire706 ) | ( wire2479 ) | ( wire22319 ) ;
 assign wire22322 = ( wire2486 ) | ( wire2491 ) | ( wire22308 ) | ( wire22314 ) ;
 assign wire22326 = ( n_n1137 ) | ( n_n1138 ) | ( n_n1099 ) | ( wire22302 ) ;
 assign wire22327 = ( n_n1095 ) | ( n_n1096 ) | ( wire22321 ) | ( wire22322 ) ;
 assign wire22328 = ( n_n1097 ) | ( n_n1102 ) | ( n_n1101 ) | ( n_n1103 ) ;
 assign wire22330 = ( wire21969 ) | ( wire21970 ) | ( wire21992 ) | ( wire21993 ) ;
 assign wire22331 = ( n_n1089 ) | ( wire21927 ) | ( wire21928 ) | ( wire21950 ) ;
 assign wire22332 = ( n_n1092 ) | ( n_n1093 ) | ( wire22101 ) | ( wire22330 ) ;
 assign wire22334 = ( wire22326 ) | ( wire22327 ) | ( wire22328 ) | ( wire22332 ) ;
 assign wire22335 = ( (~ i_15_)  &  n_n275  &  n_n279 ) | ( i_15_  &  n_n275  &  n_n256 ) ;
 assign wire22336 = ( wire913  &  n_n256 ) | ( n_n256  &  wire908 ) ;
 assign wire22337 = ( n_n4  &  n_n197 ) | ( n_n4  &  n_n21 ) | ( n_n4  &  n_n70 ) ;
 assign wire22338 = ( wire2472 ) | ( wire2473 ) | ( wire22337 ) ;
 assign wire22340 = ( (~ i_15_)  &  n_n253  &  n_n279 ) | ( i_15_  &  n_n253  &  n_n256 ) ;
 assign wire22341 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire906 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire906 ) ;
 assign wire22343 = ( n_n34 ) | ( n_n44 ) | ( wire47 ) | ( wire22341 ) ;
 assign wire22345 = ( n_n40 ) | ( n_n44 ) | ( wire245 ) | ( wire22341 ) ;
 assign wire22346 = ( n_n4  &  n_n46 ) | ( n_n4  &  wire900  &  n_n258 ) ;
 assign wire22348 = ( n_n7246 ) | ( wire2463 ) | ( wire2464 ) | ( wire22346 ) ;
 assign wire22351 = ( n_n4  &  wire320 ) | ( n_n4  &  n_n256  &  wire908 ) ;
 assign wire22352 = ( n_n256  &  wire914 ) | ( n_n256  &  wire907 ) ;
 assign wire22355 = ( n_n34 ) | ( n_n78 ) | ( wire47 ) | ( wire65 ) ;
 assign wire22356 = ( wire642 ) | ( n_n3  &  wire1217 ) ;
 assign wire22358 = ( n_n385 ) | ( wire2447 ) | ( wire22356 ) ;
 assign wire22360 = ( n_n4  &  n_n258  &  wire906 ) | ( n_n4  &  n_n258  &  wire908 ) ;
 assign wire22361 = ( n_n3  &  n_n252 ) | ( n_n4  &  wire1344 ) | ( n_n3  &  wire1344 ) ;
 assign wire22363 = ( n_n258  &  wire906 ) | ( wire905  &  n_n256 ) ;
 assign wire22366 = ( n_n258  &  wire904 ) | ( n_n258  &  wire907 ) ;
 assign wire22368 = ( wire52 ) | ( wire22366 ) | ( n_n279  &  wire913 ) ;
 assign wire22369 = ( n_n100  &  wire911  &  n_n258 ) | ( n_n100  &  n_n258  &  wire907 ) ;
 assign wire22370 = ( n_n100  &  n_n13 ) | ( n_n94  &  n_n13 ) | ( n_n100  &  wire1066 ) ;
 assign wire22372 = ( n_n2732 ) | ( wire22369 ) | ( wire22370 ) ;
 assign wire22374 = ( (~ i_15_)  &  n_n279  &  n_n267 ) | ( i_15_  &  n_n258  &  n_n267 ) ;
 assign wire22376 = ( (~ i_15_)  &  n_n279  &  n_n267 ) | ( i_15_  &  n_n258  &  n_n267 ) ;
 assign wire22378 = ( n_n57  &  n_n54 ) | ( n_n94  &  n_n61 ) ;
 assign wire22379 = ( n_n100  &  n_n257 ) | ( n_n94  &  n_n257 ) | ( n_n100  &  n_n236 ) ;
 assign wire22380 = ( n_n240  &  wire168 ) | ( n_n57  &  wire486 ) ;
 assign wire22382 = ( wire22378 ) | ( wire22379 ) | ( wire22380 ) ;
 assign wire22383 = ( wire2425 ) | ( wire2426 ) | ( wire2427 ) | ( wire2428 ) ;
 assign wire22384 = ( n_n100  &  n_n258  &  wire897 ) | ( n_n94  &  n_n258  &  wire897 ) ;
 assign wire22387 = ( i_15_  &  n_n275  &  n_n256 ) | ( (~ i_15_)  &  n_n275  &  n_n256 ) | ( i_15_  &  n_n259  &  n_n256 ) | ( (~ i_15_)  &  n_n259  &  n_n256 ) ;
 assign wire22389 = ( n_n197  &  n_n100 ) | ( n_n94  &  n_n216 ) ;
 assign wire22391 = ( wire22389 ) | ( n_n94  &  wire1069 ) | ( n_n94  &  wire140 ) ;
 assign wire22393 = ( n_n462 ) | ( wire2403 ) | ( wire22391 ) ;
 assign wire22395 = ( n_n48  &  wire911  &  n_n258 ) | ( n_n53  &  wire911  &  n_n258 ) ;
 assign wire22399 = ( n_n48  &  n_n197 ) | ( n_n53  &  n_n197 ) | ( n_n53  &  wire123 ) ;
 assign wire22400 = ( wire22399 ) | ( wire2392 ) ;
 assign wire22401 = ( wire624 ) | ( wire2393 ) | ( wire2398 ) | ( wire22395 ) ;
 assign wire22403 = ( n_n48  &  n_n246 ) | ( n_n53  &  n_n61 ) ;
 assign wire22404 = ( n_n53  &  wire903  &  n_n258 ) | ( n_n53  &  n_n258  &  wire905 ) ;
 assign wire22407 = ( n_n258  &  wire904 ) | ( n_n258  &  wire907 ) ;
 assign wire22408 = ( n_n258  &  wire914 ) | ( n_n258  &  wire904 ) ;
 assign wire22409 = ( n_n53  &  n_n10 ) | ( n_n48  &  n_n13 ) | ( n_n53  &  n_n13 ) ;
 assign wire22412 = ( n_n4153 ) | ( n_n618 ) | ( wire2378 ) ;
 assign wire22414 = ( n_n48  &  wire912  &  n_n256 ) | ( n_n48  &  n_n256  &  wire914 ) ;
 assign wire22415 = ( n_n54  &  n_n6 ) | ( n_n53  &  n_n10 ) ;
 assign wire22416 = ( n_n48  &  n_n246 ) | ( n_n6  &  n_n98 ) ;
 assign wire22421 = ( n_n6534 ) | ( n_n429 ) | ( wire2363 ) | ( wire2364 ) ;
 assign wire22426 = ( n_n6678 ) | ( wire2359 ) | ( n_n5  &  wire1648 ) ;
 assign wire22429 = ( n_n256  &  wire904 ) | ( n_n256  &  wire907 ) ;
 assign wire22431 = ( n_n34 ) | ( n_n52 ) | ( wire47 ) | ( wire22340 ) ;
 assign wire22432 = ( n_n6  &  wire1700 ) | ( n_n6  &  n_n256  &  wire914 ) ;
 assign wire22435 = ( wire306 ) | ( wire22335 ) | ( n_n222  &  wire903 ) ;
 assign wire22436 = ( wire903  &  n_n256 ) | ( n_n256  &  wire908 ) ;
 assign wire22438 = ( n_n78 ) | ( n_n199 ) | ( wire65 ) | ( wire22335 ) ;
 assign wire22440 = ( n_n423 ) | ( wire2344 ) | ( wire2345 ) ;
 assign wire22443 = ( n_n48  &  n_n31 ) | ( n_n53  &  n_n26 ) ;
 assign wire22446 = ( n_n48  &  n_n103 ) | ( n_n53  &  n_n103 ) | ( n_n53  &  wire140 ) ;
 assign wire22447 = ( wire2336 ) | ( wire22443 ) | ( n_n53  &  n_n78 ) ;
 assign wire22449 = ( n_n53  &  wire112 ) | ( n_n53  &  wire901  &  n_n258 ) ;
 assign wire22451 = ( wire407 ) | ( wire457 ) | ( n_n56  &  n_n257 ) ;
 assign wire22454 = ( n_n48  &  n_n105 ) | ( n_n53  &  n_n105 ) | ( n_n53  &  wire175 ) ;
 assign wire22456 = ( n_n56  &  wire1677 ) | ( n_n57  &  wire1676 ) | ( n_n56  &  wire1676 ) ;
 assign wire22457 = ( wire22456 ) | ( n_n57  &  wire1678 ) ;
 assign wire22459 = ( i_15_  &  n_n247  &  n_n256 ) | ( (~ i_15_)  &  n_n247  &  n_n256 ) | ( i_15_  &  n_n267  &  n_n256 ) | ( (~ i_15_)  &  n_n267  &  n_n256 ) ;
 assign wire22461 = ( n_n53  &  n_n41 ) | ( n_n48  &  n_n104 ) ;
 assign wire22463 = ( wire2311 ) | ( wire22461 ) | ( n_n54  &  n_n48 ) ;
 assign wire22464 = ( wire2333 ) | ( wire22449 ) | ( n_n53  &  wire1128 ) ;
 assign wire22467 = ( wire292 ) | ( n_n258  &  wire904 ) ;
 assign wire22468 = ( wire52 ) | ( wire441 ) | ( wire911  &  n_n258 ) ;
 assign wire22469 = ( wire42 ) | ( wire899  &  n_n258 ) | ( n_n258  &  wire907 ) ;
 assign wire22471 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire22473 = ( wire57 ) | ( wire414 ) | ( n_n258  &  wire912 ) ;
 assign wire22474 = ( wire233 ) | ( wire444 ) | ( n_n222  &  wire907 ) ;
 assign wire22475 = ( (~ i_15_)  &  n_n253  &  n_n279 ) | ( i_15_  &  n_n253  &  n_n256 ) | ( (~ i_15_)  &  n_n253  &  n_n256 ) ;
 assign wire22476 = ( wire53 ) | ( wire405 ) | ( n_n258  &  wire897 ) ;
 assign wire22477 = ( i_14_  &  i_13_  &  (~ i_12_)  &  wire908 ) | ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  wire908 ) ;
 assign wire22481 = ( wire2299 ) | ( wire2300 ) | ( wire2306 ) | ( wire2307 ) ;
 assign wire22483 = ( wire166  &  n_n100 ) | ( n_n100  &  wire900  &  n_n258 ) ;
 assign wire22485 = ( wire20755 ) | ( n_n54  &  n_n100 ) | ( n_n54  &  n_n94 ) ;
 assign wire22487 = ( wire2291 ) | ( n_n100  &  wire1305 ) ;
 assign wire22488 = ( wire54 ) | ( wire266 ) | ( wire913  &  n_n220 ) ;
 assign wire22489 = ( i_7_  &  i_6_  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  i_6_  &  n_n118  &  n_n230 ) | ( i_7_  &  (~ i_6_)  &  n_n118  &  n_n230 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n118  &  n_n230 ) ;
 assign wire22490 = ( i_7_  &  i_6_  &  n_n230  &  n_n116 ) | ( (~ i_7_)  &  i_6_  &  n_n230  &  n_n116 ) | ( i_7_  &  (~ i_6_)  &  n_n230  &  n_n116 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n230  &  n_n116 ) ;
 assign wire22491 = ( wire22489 ) | ( n_n136  &  wire1307 ) ;
 assign wire22492 = ( wire394 ) | ( wire22490 ) | ( n_n139  &  wire48 ) ;
 assign wire22493 = ( wire22240 ) | ( wire22241 ) | ( wire22242 ) | ( wire22491 ) ;
 assign wire22494 = ( wire22492 ) | ( n_n139  &  wire294 ) | ( n_n139  &  wire22488 ) ;
 assign wire22495 = ( n_n94  &  n_n41 ) | ( n_n100  &  n_n81 ) ;
 assign wire22496 = ( n_n100  &  wire901  &  n_n258 ) | ( n_n100  &  wire901  &  n_n256 ) ;
 assign wire22502 = ( wire881 ) | ( wire688 ) | ( wire798 ) | ( wire2269 ) ;
 assign wire22504 = ( n_n464 ) | ( wire22502 ) | ( n_n100  &  wire1261 ) ;
 assign wire22506 = ( wire901  &  n_n258 ) | ( wire898  &  n_n258 ) ;
 assign wire22510 = ( n_n41 ) | ( n_n113 ) | ( wire57 ) | ( wire229 ) ;
 assign wire22511 = ( wire2264 ) | ( wire2267 ) | ( wire2268 ) ;
 assign wire22512 = ( wire902  &  n_n258 ) | ( n_n258  &  wire912 ) ;
 assign wire22513 = ( i_15_  &  n_n275  &  n_n256 ) | ( (~ i_15_)  &  n_n275  &  n_n256 ) | ( i_15_  &  n_n247  &  n_n256 ) | ( (~ i_15_)  &  n_n247  &  n_n256 ) ;
 assign wire22515 = ( wire902  &  n_n258 ) | ( n_n258  &  wire897 ) ;
 assign wire22516 = ( i_11_  &  i_15_  &  n_n163  &  n_n256 ) | ( (~ i_11_)  &  i_15_  &  n_n163  &  n_n256 ) | ( i_11_  &  (~ i_15_)  &  n_n163  &  n_n256 ) | ( (~ i_11_)  &  (~ i_15_)  &  n_n163  &  n_n256 ) ;
 assign wire22518 = ( wire2263 ) | ( n_n2  &  wire1311 ) | ( n_n2  &  wire1733 ) ;
 assign wire22519 = ( i_14_  &  (~ i_13_)  &  i_12_  &  wire907 ) | ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  wire907 ) ;
 assign wire22522 = ( n_n53  &  n_n257 ) | ( n_n53  &  n_n61 ) | ( n_n53  &  wire123 ) ;
 assign wire22523 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n256 ) | ( (~ i_15_)  &  n_n267  &  n_n256 ) ;
 assign wire22524 = ( wire2246 ) | ( n_n2  &  wire166 ) | ( n_n2  &  wire22523 ) ;
 assign wire22527 = ( wire2260 ) | ( wire2265 ) | ( wire22511 ) | ( wire22518 ) ;
 assign wire22531 = ( wire57 ) | ( wire444 ) | ( n_n258  &  wire912 ) ;
 assign wire22532 = ( n_n268  &  n_n240 ) | ( n_n3  &  wire408 ) ;
 assign wire22533 = ( wire22532 ) | ( n_n4  &  wire1348 ) ;
 assign wire22535 = ( i_15_  &  n_n242  &  n_n258 ) | ( i_15_  &  n_n242  &  n_n256 ) | ( (~ i_15_)  &  n_n242  &  n_n256 ) ;
 assign wire22536 = ( wire2235 ) | ( n_n2  &  wire140 ) | ( n_n2  &  wire182 ) ;
 assign wire22537 = ( wire2237 ) | ( wire2239 ) | ( wire2240 ) ;
 assign wire22538 = ( n_n1  &  n_n236 ) | ( n_n1  &  wire1673 ) | ( n_n2  &  wire1673 ) ;
 assign wire22539 = ( n_n1  &  n_n240 ) | ( n_n2  &  n_n240 ) | ( n_n2  &  wire403 ) ;
 assign wire22540 = ( n_n216 ) | ( n_n103 ) | ( wire52 ) | ( wire53 ) ;
 assign wire22541 = ( n_n1  &  wire1357 ) | ( n_n1  &  wire1355 ) | ( n_n2  &  wire1355 ) ;
 assign wire22543 = ( wire2225 ) | ( wire22538 ) | ( wire22539 ) | ( wire22541 ) ;
 assign wire22544 = ( wire22543 ) | ( n_n268  &  wire405 ) | ( n_n268  &  wire22540 ) ;
 assign wire22546 = ( n_n10  &  n_n100 ) | ( n_n94  &  n_n41 ) ;
 assign wire22547 = ( n_n100  &  n_n81 ) | ( n_n94  &  n_n86 ) ;
 assign wire22548 = ( n_n94  &  wire57 ) | ( n_n94  &  wire903  &  n_n258 ) ;
 assign wire22551 = ( n_n207  &  n_n257 ) | ( n_n94  &  n_n246 ) ;
 assign wire22552 = ( n_n4  &  n_n26 ) | ( n_n100  &  n_n104 ) ;
 assign wire22556 = ( wire22552 ) | ( wire22551 ) ;
 assign wire22557 = ( wire743 ) | ( wire2205 ) | ( n_n227  &  n_n257 ) ;
 assign wire22558 = ( wire642 ) | ( wire471 ) | ( wire658 ) | ( wire2206 ) ;
 assign wire22561 = ( n_n53  &  n_n197 ) | ( n_n4  &  n_n257 ) ;
 assign wire22562 = ( n_n53  &  n_n26 ) | ( n_n3  &  n_n252 ) ;
 assign wire22565 = ( n_n53  &  n_n31 ) | ( n_n53  &  n_n78 ) | ( n_n53  &  wire140 ) ;
 assign wire22566 = ( n_n240  &  n_n6 ) | ( n_n207  &  n_n103 ) ;
 assign wire22567 = ( n_n5  &  n_n257 ) | ( n_n227  &  wire276 ) ;
 assign wire22570 = ( n_n6  &  wire1680 ) | ( n_n6  &  wire1679 ) | ( n_n5  &  wire1679 ) ;
 assign wire22571 = ( n_n207  &  wire292 ) | ( n_n5  &  wire1682 ) ;
 assign wire22572 = ( wire2196 ) | ( wire22570 ) ;
 assign wire22573 = ( wire2200 ) | ( wire22566 ) | ( wire22567 ) | ( wire22571 ) ;
 assign wire22574 = ( n_n4  &  wire900  &  n_n258 ) | ( n_n4  &  n_n258  &  wire906 ) ;
 assign wire22575 = ( n_n4  &  n_n61 ) | ( n_n4  &  n_n228  &  wire906 ) ;
 assign wire22576 = ( n_n4  &  n_n70 ) | ( n_n3  &  n_n49 ) ;
 assign wire22578 = ( wire22574 ) | ( wire22575 ) | ( wire22576 ) ;
 assign wire22581 = ( wire833 ) | ( n_n409 ) | ( wire2183 ) | ( wire22578 ) ;
 assign wire22587 = ( n_n346 ) | ( n_n343 ) | ( n_n341 ) ;
 assign wire22588 = ( n_n342 ) | ( n_n344 ) | ( n_n345 ) | ( n_n347 ) ;
 assign wire22590 = ( n_n4  &  n_n257 ) | ( n_n3  &  n_n257 ) | ( n_n3  &  n_n61 ) ;
 assign wire22593 = ( n_n380 ) | ( n_n381 ) | ( wire2176 ) | ( wire22590 ) ;
 assign wire22594 = ( n_n349 ) | ( n_n351 ) | ( wire22358 ) | ( wire22593 ) ;
 assign wire22596 = ( n_n4  &  n_n80 ) | ( n_n4  &  wire114 ) | ( n_n4  &  wire88 ) ;
 assign wire22597 = ( i_15_  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n225 ) | ( (~ i_15_)  &  n_n275  &  n_n225 ) ;
 assign wire22598 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign wire22599 = ( n_n80 ) | ( n_n203 ) | ( wire88 ) | ( wire20149 ) ;
 assign wire22600 = ( n_n4  &  n_n197 ) | ( n_n3  &  n_n216 ) ;
 assign wire22602 = ( n_n876 ) | ( wire2162 ) | ( wire22600 ) ;
 assign wire22605 = ( n_n100  &  n_n65 ) | ( n_n94  &  n_n65 ) | ( n_n100  &  n_n15 ) ;
 assign wire22606 = ( n_n94  &  wire911  &  n_n258 ) | ( n_n94  &  wire899  &  n_n258 ) ;
 assign wire22610 = ( wire697 ) | ( n_n100  &  n_n216 ) | ( n_n100  &  wire1061 ) ;
 assign wire22611 = ( n_n1058 ) | ( n_n3604 ) | ( n_n3610 ) | ( wire22606 ) ;
 assign wire22613 = ( n_n94  &  n_n226 ) | ( n_n100  &  n_n206 ) | ( n_n94  &  n_n206 ) ;
 assign wire22616 = ( n_n100  &  n_n63 ) | ( n_n94  &  n_n63 ) | ( n_n100  &  n_n226 ) ;
 assign wire22618 = ( n_n100  &  wire1121 ) | ( n_n94  &  wire1120 ) ;
 assign wire22620 = ( wire22618 ) | ( n_n57  &  wire224 ) | ( n_n56  &  wire224 ) ;
 assign wire22625 = ( n_n4954 ) | ( wire2128 ) | ( n_n56  &  wire254 ) ;
 assign wire22626 = ( wire2129 ) | ( n_n57  &  wire277 ) | ( n_n56  &  wire277 ) ;
 assign wire22629 = ( wire60 ) | ( wire227 ) | ( n_n279  &  wire911 ) ;
 assign wire22630 = ( wire348 ) | ( wire305 ) ;
 assign wire22631 = ( i_15_  &  n_n253  &  n_n258 ) | ( i_15_  &  n_n253  &  n_n225 ) | ( (~ i_15_)  &  n_n253  &  n_n225 ) ;
 assign wire22633 = ( wire571 ) | ( wire737 ) | ( n_n48  &  n_n105 ) ;
 assign wire22635 = ( wire5591 ) | ( wire5592 ) | ( n_n56  &  n_n9 ) ;
 assign wire22636 = ( n_n57  &  n_n226 ) | ( n_n56  &  n_n226 ) | ( n_n57  &  wire1717 ) | ( n_n56  &  wire1717 ) ;
 assign wire22637 = ( n_n57  &  n_n11 ) | ( n_n57  &  n_n65 ) | ( n_n56  &  n_n65 ) ;
 assign wire22638 = ( n_n57  &  wire1753 ) | ( n_n56  &  wire1752 ) ;
 assign wire22639 = ( wire22635 ) | ( wire22636 ) | ( wire22637 ) ;
 assign wire22640 = ( wire2122 ) | ( wire22633 ) | ( wire22638 ) ;
 assign wire22642 = ( n_n56  &  n_n179 ) | ( n_n56  &  wire190 ) | ( n_n56  &  wire55 ) ;
 assign wire22643 = ( n_n57  &  wire190 ) | ( n_n57  &  wire198 ) ;
 assign wire22646 = ( wire2103 ) | ( wire2104 ) | ( wire22642 ) | ( wire22643 ) ;
 assign wire22647 = ( wire2126 ) | ( wire2127 ) | ( wire22639 ) | ( wire22640 ) ;
 assign wire22648 = ( n_n100  &  wire120 ) | ( n_n100  &  wire899  &  n_n258 ) ;
 assign wire22650 = ( i_15_  &  n_n275  &  n_n225 ) | ( (~ i_15_)  &  n_n275  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign wire22651 = ( n_n100  &  n_n103 ) | ( n_n94  &  n_n39 ) ;
 assign wire22652 = ( n_n31  &  n_n100 ) | ( n_n94  &  n_n103 ) ;
 assign wire22654 = ( n_n3870 ) | ( wire22651 ) | ( wire22652 ) ;
 assign wire22657 = ( i_15_  &  n_n258  &  n_n282 ) | ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire22658 = ( n_n94  &  n_n41 ) | ( n_n100  &  n_n36 ) ;
 assign wire22659 = ( n_n37  &  n_n100 ) | ( n_n100  &  n_n84 ) | ( n_n100  &  n_n104 ) ;
 assign wire22662 = ( n_n1066 ) | ( wire2082 ) | ( wire22658 ) ;
 assign wire22663 = ( wire767 ) | ( wire2081 ) | ( wire2089 ) | ( wire22659 ) ;
 assign wire22664 = ( i_15_  &  n_n253  &  n_n225 ) | ( (~ i_15_)  &  n_n253  &  n_n225 ) | ( i_15_  &  n_n267  &  n_n225 ) | ( (~ i_15_)  &  n_n267  &  n_n225 ) ;
 assign wire22665 = ( n_n105  &  n_n100 ) | ( n_n54  &  n_n94 ) ;
 assign wire22667 = ( n_n3884 ) | ( wire22665 ) | ( n_n94  &  wire139 ) ;
 assign wire22668 = ( wire2072 ) | ( wire776 ) ;
 assign wire22670 = ( wire19379 ) | ( wire19380 ) | ( wire22667 ) | ( wire22668 ) ;
 assign wire22672 = ( n_n6  &  wire120 ) | ( n_n6  &  n_n25 ) | ( n_n6  &  wire19457 ) ;
 assign wire22674 = ( wire469 ) | ( wire128 ) | ( n_n222  &  wire899 ) ;
 assign wire22675 = ( wire898  &  n_n228 ) | ( wire899  &  n_n258 ) ;
 assign wire22676 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n259  &  n_n225 ) | ( (~ i_15_)  &  n_n259  &  n_n225 ) ;
 assign wire22678 = ( wire647 ) | ( wire2067 ) | ( n_n5  &  n_n197 ) ;
 assign wire22680 = ( n_n6  &  wire899  &  n_n228 ) | ( n_n6  &  n_n228  &  wire897 ) ;
 assign wire22681 = ( n_n6  &  n_n206 ) | ( n_n5  &  n_n206 ) | ( n_n5  &  wire1253 ) ;
 assign wire22683 = ( n_n6  &  wire1640 ) | ( n_n6  &  wire1638 ) | ( n_n5  &  wire1638 ) ;
 assign wire22684 = ( n_n227  &  wire275 ) | ( n_n5  &  wire1639 ) ;
 assign wire22685 = ( wire887 ) | ( wire22683 ) ;
 assign wire22686 = ( wire2059 ) | ( wire22680 ) | ( wire22681 ) | ( wire22684 ) ;
 assign wire22687 = ( i_15_  &  n_n275  &  n_n258 ) | ( i_15_  &  n_n275  &  n_n225 ) | ( (~ i_15_)  &  n_n275  &  n_n225 ) ;
 assign wire22689 = ( n_n6  &  wire114 ) | ( n_n6  &  n_n258  &  wire897 ) ;
 assign wire22692 = ( wire22672 ) | ( n_n5  &  wire1641 ) | ( n_n5  &  wire1918 ) ;
 assign wire22693 = ( n_n4636 ) | ( wire487 ) | ( wire22689 ) | ( wire22692 ) ;
 assign wire22695 = ( n_n48  &  n_n31 ) | ( n_n48  &  n_n80 ) | ( n_n48  &  wire88 ) ;
 assign wire22696 = ( i_15_  &  n_n242  &  n_n225 ) | ( (~ i_15_)  &  n_n242  &  n_n225 ) | ( i_15_  &  n_n225  &  n_n270 ) | ( (~ i_15_)  &  n_n225  &  n_n270 ) ;
 assign wire22698 = ( n_n53  &  n_n197 ) | ( n_n48  &  n_n216 ) | ( n_n53  &  n_n216 ) ;
 assign wire22700 = ( wire2035 ) | ( wire2034 ) ;
 assign wire22701 = ( n_n4073 ) | ( wire2041 ) | ( wire22695 ) | ( wire22698 ) ;
 assign wire22703 = ( n_n53  &  wire114 ) | ( n_n48  &  n_n103 ) | ( n_n53  &  n_n103 ) ;
 assign wire22704 = ( n_n48  &  n_n41 ) | ( n_n53  &  n_n104 ) ;
 assign wire22708 = ( n_n4094 ) | ( n_n4090 ) | ( wire2023 ) | ( wire22704 ) ;
 assign wire22709 = ( wire483 ) | ( wire2022 ) | ( wire2030 ) | ( wire22703 ) ;
 assign wire22710 = ( n_n48  &  n_n37 ) | ( n_n48  &  wire89 ) | ( n_n48  &  n_n104 ) ;
 assign wire22711 = ( wire134 ) | ( wire96 ) | ( n_n222  &  wire898 ) ;
 assign wire22712 = ( n_n53  &  wire900  &  n_n258 ) | ( n_n53  &  n_n258  &  wire912 ) ;
 assign wire22714 = ( wire2012 ) | ( wire22712 ) | ( n_n54  &  n_n48 ) ;
 assign wire22717 = ( wire22700 ) | ( wire22701 ) | ( wire22708 ) | ( wire22709 ) ;
 assign wire22719 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) | ( (~ i_15_)  &  n_n267  &  n_n225 ) ;
 assign wire22720 = ( n_n54  &  n_n6 ) | ( n_n53  &  n_n63 ) ;
 assign wire22722 = ( wire670 ) | ( wire22720 ) | ( n_n48  &  n_n11 ) ;
 assign wire22725 = ( n_n48  &  wire899  &  n_n228 ) | ( n_n53  &  wire899  &  n_n228 ) ;
 assign wire22727 = ( n_n48  &  n_n206 ) | ( n_n53  &  n_n206 ) | ( n_n53  &  wire1062 ) ;
 assign wire22730 = ( wire898  &  n_n228 ) | ( n_n228  &  wire912 ) ;
 assign wire22731 = ( n_n53  &  n_n9 ) | ( n_n48  &  n_n15 ) ;
 assign wire22732 = ( n_n48  &  n_n197 ) | ( n_n48  &  wire1063 ) | ( n_n53  &  wire1063 ) ;
 assign wire22734 = ( wire22732 ) | ( n_n48  &  wire1064 ) ;
 assign wire22736 = ( n_n5  &  n_n41 ) | ( n_n6  &  n_n104 ) ;
 assign wire22740 = ( n_n99 ) | ( n_n37 ) | ( wire89 ) | ( wire96 ) ;
 assign wire22742 = ( n_n4644 ) | ( wire1977 ) | ( n_n54  &  n_n5 ) ;
 assign wire22744 = ( n_n819 ) | ( wire1978 ) | ( wire22742 ) ;
 assign wire22746 = ( i_15_  &  n_n247  &  n_n258 ) | ( i_15_  &  n_n247  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign wire22748 = ( wire60 ) | ( wire198 ) | ( n_n279  &  wire911 ) ;
 assign wire22752 = ( wire60 ) | ( n_n204 ) | ( wire227 ) | ( wire348 ) ;
 assign wire22754 = ( wire55 ) | ( wire304 ) | ( n_n279  &  wire912 ) ;
 assign wire22757 = ( wire301 ) | ( wire254 ) | ( wire335 ) ;
 assign wire22758 = ( wire190 ) | ( wire55 ) | ( n_n279  &  wire912 ) ;
 assign wire22761 = ( wire198 ) | ( wire190 ) ;
 assign wire22762 = ( wire301 ) | ( wire277 ) | ( wire275 ) ;
 assign wire22763 = ( wire1964 ) | ( n_n1  &  wire22761 ) | ( n_n1  &  wire22762 ) ;
 assign wire22764 = ( wire1968 ) | ( wire1969 ) | ( wire1970 ) | ( wire1971 ) ;
 assign wire22765 = ( n_n279  &  wire911 ) | ( wire903  &  n_n225 ) ;
 assign wire22766 = ( i_14_  &  i_13_  &  i_12_  &  wire913 ) | ( (~ i_14_)  &  i_13_  &  i_12_  &  wire913 ) ;
 assign wire22769 = ( i_14_  &  n_n254  &  wire911 ) | ( (~ i_14_)  &  n_n254  &  wire914 ) ;
 assign wire22772 = ( i_15_  &  n_n282  &  n_n225 ) | ( (~ i_15_)  &  n_n282  &  n_n225 ) ;
 assign wire22775 = ( n_n1  &  wire899  &  n_n228 ) | ( n_n2  &  wire899  &  n_n228 ) ;
 assign wire22776 = ( wire135  &  n_n206 ) | ( n_n268  &  wire56 ) ;
 assign wire22778 = ( n_n1  &  n_n65 ) | ( n_n2  &  n_n65 ) | ( n_n1  &  n_n15 ) ;
 assign wire22780 = ( n_n1  &  n_n59 ) | ( n_n2  &  n_n59 ) | ( n_n1  &  wire1606 ) ;
 assign wire22781 = ( wire22780 ) | ( n_n2  &  n_n15 ) | ( n_n2  &  wire1606 ) ;
 assign wire22783 = ( i_14_  &  i_13_  &  i_12_  &  wire901 ) | ( i_14_  &  (~ i_13_)  &  i_12_  &  wire901 ) ;
 assign wire22785 = ( n_n53  &  wire899  &  n_n228 ) | ( n_n53  &  n_n228  &  wire902 ) ;
 assign wire22786 = ( n_n4  &  n_n9 ) | ( n_n4  &  wire900  &  n_n258 ) ;
 assign wire22787 = ( n_n4  &  wire899  &  n_n228 ) | ( n_n4  &  wire900  &  n_n228 ) ;
 assign wire22788 = ( n_n4  &  n_n197 ) | ( n_n3  &  n_n15 ) ;
 assign wire22792 = ( wire608 ) | ( wire22786 ) | ( n_n4  &  wire1669 ) ;
 assign wire22793 = ( n_n876 ) | ( wire544 ) | ( wire22787 ) | ( wire22788 ) ;
 assign wire22795 = ( (~ i_15_)  &  n_n259  &  n_n228 ) | ( i_15_  &  n_n259  &  n_n258 ) ;
 assign wire22796 = ( n_n9  &  n_n207 ) | ( n_n94  &  n_n203 ) ;
 assign wire22797 = ( n_n9  &  n_n227 ) | ( n_n207  &  n_n59 ) ;
 assign wire22801 = ( n_n94  &  n_n204 ) | ( n_n100  &  n_n84 ) ;
 assign wire22803 = ( wire548 ) | ( n_n100  &  n_n104 ) | ( n_n100  &  n_n36 ) ;
 assign wire22804 = ( wire697 ) | ( wire22801 ) | ( n_n100  &  n_n33 ) ;
 assign wire22805 = ( n_n4  &  n_n31 ) | ( n_n94  &  n_n39 ) ;
 assign wire22806 = ( n_n11  &  n_n94 ) | ( n_n100  &  n_n63 ) ;
 assign wire22809 = ( n_n884 ) | ( wire564 ) | ( wire22805 ) | ( wire22806 ) ;
 assign wire22812 = ( wire543 ) | ( n_n53  &  wire275 ) | ( n_n53  &  wire305 ) ;
 assign wire22814 = ( n_n803 ) | ( n_n952 ) | ( wire550 ) | ( wire22812 ) ;
 assign wire22816 = ( i_15_  &  n_n258  &  n_n267 ) | ( i_15_  &  n_n267  &  n_n225 ) | ( (~ i_15_)  &  n_n267  &  n_n225 ) ;
 assign wire22818 = ( wire529 ) | ( n_n4  &  n_n105 ) | ( n_n4  &  wire134 ) ;
 assign wire22820 = ( n_n785 ) | ( wire1975 ) | ( wire1976 ) | ( wire22818 ) ;
 assign wire22822 = ( n_n749 ) | ( n_n750 ) | ( wire22820 ) ;
 assign wire22827 = ( n_n743 ) | ( n_n742 ) | ( n_n744 ) | ( n_n739 ) ;
 assign wire22829 = ( n_n4  &  wire899  &  n_n228 ) | ( n_n4  &  n_n228  &  wire902 ) ;
 assign wire22830 = ( n_n3  &  n_n226 ) | ( n_n4  &  n_n59 ) ;
 assign wire22833 = ( wire900  &  n_n228 ) | ( wire899  &  n_n258 ) ;
 assign wire22835 = ( wire898  &  n_n228 ) | ( n_n228  &  wire912 ) ;
 assign wire22837 = ( n_n4  &  n_n65 ) | ( n_n3  &  n_n15 ) ;
 assign wire22839 = ( wire505 ) | ( wire22837 ) | ( n_n3  &  wire1836 ) ;
 assign wire22841 = ( i_15_  &  n_n247  &  n_n258 ) | ( i_15_  &  n_n247  &  n_n225 ) | ( (~ i_15_)  &  n_n247  &  n_n225 ) ;
 assign wire22843 = ( wire238 ) | ( n_n4  &  wire126 ) | ( n_n4  &  n_n31 ) ;
 assign wire22844 = ( wire2170 ) | ( wire2173 ) | ( wire2174 ) | ( wire22596 ) ;
 assign wire22847 = ( n_n746 ) | ( n_n745 ) | ( wire22843 ) | ( wire22844 ) ;


endmodule

