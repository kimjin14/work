module des (
	pcount_3_, pdata_22_, pdata_35_, pdata_48_, pinreg_1_, poutreg_51_, pcount_2_, pdata_10_, 
	pdata_21_, pdata_36_, pdata_47_, pinreg_0_, poutreg_52_, poutreg_63_, pcount_1_, pdata_8_, pdata_24_, pdata_37_, 
	pdata_46_, pdata_59_, poutreg_40_, poutreg_53_, poutreg_62_, pcount_0_, pdata_9_, pdata_23_, pdata_38_, pdata_45_, 
	poutreg_54_, poutreg_61_, pdata_6_, pdata_26_, pdata_31_, pdata_44_, pinreg_5_, poutreg_55_, pdata_7_, pdata_25_, 
	pdata_32_, pdata_43_, pinreg_4_, poutreg_30_, poutreg_56_, pdata_4_, pdata_28_, pdata_33_, pdata_42_, pinreg_3_, 
	poutreg_57_, pdata_5_, pdata_27_, pdata_34_, pdata_41_, pinreg_2_, poutreg_58_, pd_20_, pdata_17_, pdata_40_, 
	pinreg_9_, poutreg_0_, poutreg_33_, poutreg_46_, pc_20_, pd_10_, pdata_18_, pinreg_8_, poutreg_1_, poutreg_34_, 
	poutreg_45_, preset_0_, pc_21_, pd_11_, pd_22_, pdata_15_, pinreg_7_, poutreg_31_, poutreg_48_, pc_22_, 
	pd_12_, pd_21_, pdata_16_, pdata_30_, pinreg_6_, poutreg_32_, poutreg_47_, pc_12_, pdata_13_, poutreg_19_, 
	poutreg_37_, poutreg_42_, poutreg_60_, pc_11_, pdata_14_, poutreg_38_, poutreg_41_, pc_10_, pdata_11_, pdata_20_, 
	poutreg_35_, poutreg_44_, pdata_12_, poutreg_29_, poutreg_36_, poutreg_43_, poutreg_50_, pc_9_, pc_16_, pc_27_, 
	pd_8_, pd_17_, pdata_in_4_, pinreg_30_, pinreg_41_, pinreg_52_, poutreg_8_, poutreg_15_, poutreg_28_, pc_15_, 
	pd_9_, pd_18_, pd_27_, pdata_in_3_, pinreg_31_, pinreg_40_, pinreg_53_, poutreg_9_, poutreg_16_, poutreg_27_, 
	pc_14_, pd_19_, pdata_60_, pdata_in_6_, pinreg_32_, pinreg_43_, pinreg_50_, poutreg_6_, poutreg_17_, poutreg_26_, 
	poutreg_39_, pc_13_, pdata_in_5_, pinreg_33_, pinreg_42_, pinreg_51_, poutreg_7_, poutreg_18_, poutreg_25_, pc_5_, 
	pc_23_, pd_4_, pd_13_, pd_24_, pinreg_12_, pinreg_23_, poutreg_4_, poutreg_11_, poutreg_24_, pc_6_, 
	pc_19_, pc_24_, pd_5_, pd_14_, pd_23_, pdata_50_, pdata_in_7_, pencrypt_0_, pinreg_13_, pinreg_22_, 
	poutreg_5_, poutreg_12_, poutreg_23_, poutreg_49_, pc_7_, pc_18_, pc_25_, pd_6_, pd_15_, pd_26_, 
	pdata_19_, pinreg_10_, pinreg_21_, pload_key_0_, poutreg_2_, poutreg_13_, poutreg_22_, pc_8_, pc_17_, pc_26_, 
	pd_7_, pd_16_, pd_25_, pinreg_11_, pinreg_20_, poutreg_3_, poutreg_14_, poutreg_21_, pc_1_, pd_0_, 
	pdata_2_, pdata_53_, pinreg_16_, pinreg_27_, pinreg_38_, pinreg_49_, poutreg_20_, poutreg_59_, pc_2_, pd_1_, 
	pdata_3_, pdata_29_, pdata_54_, pinreg_17_, pinreg_26_, pinreg_39_, pinreg_48_, pc_3_, pd_2_, pdata_0_, 
	pdata_51_, pinreg_14_, pinreg_25_, pc_4_, pd_3_, pdata_1_, pdata_52_, pencrypt_mode_0_, pinreg_15_, pinreg_24_, 
	poutreg_10_, pdata_39_, pdata_57_, pdata_62_, pdata_in_0_, pinreg_34_, pinreg_45_, pdata_58_, pdata_61_, pinreg_35_, 
	pinreg_44_, pdata_55_, pdata_in_2_, pinreg_18_, pinreg_29_, pinreg_36_, pinreg_47_, pinreg_54_, pc_0_, pdata_49_, 
	pdata_56_, pdata_63_, pdata_in_1_, pinreg_19_, pinreg_28_, pinreg_37_, pinreg_46_, pinreg_55_, pc_new_6_, pc_new_19_, 
	pd_new_5_, pdata_new_14_, pdata_new_27_, pinreg_new_6_, pinreg_new_19_, poutreg_new_9_, pc_new_7_, pd_new_6_, pd_new_19_, pdata_new_13_, 
	pdata_new_28_, pdata_new_39_, pinreg_new_5_, pinreg_new_18_, poutreg_new_19_, pc_new_4_, pd_new_3_, pdata_new_9_, pdata_new_12_, pdata_new_25_, 
	pinreg_new_8_, pinreg_new_17_, poutreg_new_7_, pc_new_5_, pd_new_4_, pdata_new_11_, pdata_new_26_, pinreg_new_7_, pinreg_new_16_, poutreg_new_8_, 
	pc_new_2_, pd_new_1_, pdata_new_10_, pdata_new_36_, pinreg_new_2_, pinreg_new_15_, poutreg_new_16_, pc_new_3_, pd_new_2_, pdata_new_35_, 
	pinreg_new_1_, pinreg_new_14_, poutreg_new_15_, pc_new_0_, pdata_new_29_, pdata_new_38_, pinreg_new_4_, pinreg_new_13_, poutreg_new_18_, pc_new_1_, 
	pd_new_0_, pdata_new_37_, pinreg_new_3_, pinreg_new_12_, poutreg_new_17_, pc_new_11_, pc_new_22_, pd_new_12_, pd_new_23_, pcount_new_0_, 
	pdata_new_3_, pdata_new_45_, pdata_new_58_, pinreg_new_22_, pinreg_new_33_, pinreg_new_44_, pinreg_new_55_, poutreg_new_1_, poutreg_new_25_, poutreg_new_38_, 
	poutreg_new_61_, pc_new_12_, pc_new_21_, pd_new_11_, pd_new_24_, pdata_new_4_, pdata_new_46_, pdata_new_57_, pinreg_new_23_, pinreg_new_32_, 
	pinreg_new_45_, pinreg_new_54_, poutreg_new_2_, poutreg_new_26_, poutreg_new_37_, poutreg_new_62_, pc_new_13_, pc_new_24_, pd_new_14_, pd_new_21_, 
	pcount_new_2_, pdata_new_1_, pdata_new_47_, pdata_new_56_, pinreg_new_0_, pinreg_new_24_, pinreg_new_35_, pinreg_new_42_, pinreg_new_53_, poutreg_new_27_, 
	poutreg_new_36_, poutreg_new_49_, poutreg_new_50_, poutreg_new_63_, pc_new_14_, pc_new_23_, pd_new_13_, pd_new_22_, pcount_new_1_, pdata_new_2_, 
	pdata_new_48_, pdata_new_55_, pinreg_new_25_, pinreg_new_34_, pinreg_new_43_, pinreg_new_52_, poutreg_new_0_, poutreg_new_28_, poutreg_new_35_, pc_new_15_, 
	pc_new_26_, pd_new_16_, pd_new_27_, pdata_new_7_, pdata_new_49_, pinreg_new_26_, pinreg_new_37_, pinreg_new_48_, poutreg_new_5_, poutreg_new_29_, 
	poutreg_new_47_, poutreg_new_52_, pc_new_16_, pc_new_25_, pd_new_15_, pcount_new_3_, pdata_new_8_, pinreg_new_27_, pinreg_new_36_, pinreg_new_49_, 
	poutreg_new_6_, poutreg_new_48_, poutreg_new_51_, pc_new_17_, pd_new_18_, pd_new_25_, pdata_new_5_, pinreg_new_28_, pinreg_new_39_, pinreg_new_46_, 
	poutreg_new_3_, poutreg_new_45_, poutreg_new_54_, pc_new_18_, pc_new_27_, pd_new_17_, pd_new_26_, pdata_new_6_, pdata_new_59_, pinreg_new_29_, 
	pinreg_new_38_, pinreg_new_47_, poutreg_new_4_, poutreg_new_39_, poutreg_new_46_, poutreg_new_53_, poutreg_new_60_, pdata_new_50_, pdata_new_63_, poutreg_new_30_, 
	poutreg_new_43_, poutreg_new_56_, poutreg_new_44_, poutreg_new_55_, pdata_new_61_, pencrypt_mode_new_0_, poutreg_new_41_, poutreg_new_58_, pdata_new_40_, pdata_new_62_, 
	poutreg_new_20_, poutreg_new_42_, poutreg_new_57_, pdata_new_41_, pdata_new_54_, pinreg_new_40_, pinreg_new_51_, poutreg_new_21_, poutreg_new_34_, pd_new_20_, 
	pdata_new_0_, pdata_new_42_, pdata_new_53_, pdata_new_60_, pinreg_new_41_, pinreg_new_50_, poutreg_new_22_, poutreg_new_33_, poutreg_new_40_, poutreg_new_59_, 
	pc_new_20_, pd_new_10_, pdata_new_43_, pdata_new_52_, pinreg_new_20_, pinreg_new_31_, poutreg_new_23_, poutreg_new_32_, pc_new_10_, pdata_new_44_, 
	pdata_new_51_, pinreg_new_21_, pinreg_new_30_, poutreg_new_24_, poutreg_new_31_, pdata_new_32_, pinreg_new_11_, poutreg_new_12_, pdata_new_20_, pdata_new_31_, 
	pinreg_new_10_, poutreg_new_11_, pdata_new_34_, poutreg_new_14_, pdata_new_19_, pdata_new_33_, poutreg_new_13_, pd_new_9_, pdata_new_18_, pdata_new_23_, 
	pdata_new_17_, pdata_new_24_, pinreg_new_9_, pc_new_8_, pd_new_7_, pdata_new_16_, pdata_new_21_, pdata_new_30_, poutreg_new_10_, pc_new_9_, 
	pd_new_8_, pdata_new_15_, pdata_new_22_);

input pcount_3_;
input pdata_22_;
input pdata_35_;
input pdata_48_;
input pinreg_1_;
input poutreg_51_;
input pcount_2_;
input pdata_10_;
input pdata_21_;
input pdata_36_;
input pdata_47_;
input pinreg_0_;
input poutreg_52_;
input poutreg_63_;
input pcount_1_;
input pdata_8_;
input pdata_24_;
input pdata_37_;
input pdata_46_;
input pdata_59_;
input poutreg_40_;
input poutreg_53_;
input poutreg_62_;
input pcount_0_;
input pdata_9_;
input pdata_23_;
input pdata_38_;
input pdata_45_;
input poutreg_54_;
input poutreg_61_;
input pdata_6_;
input pdata_26_;
input pdata_31_;
input pdata_44_;
input pinreg_5_;
input poutreg_55_;
input pdata_7_;
input pdata_25_;
input pdata_32_;
input pdata_43_;
input pinreg_4_;
input poutreg_30_;
input poutreg_56_;
input pdata_4_;
input pdata_28_;
input pdata_33_;
input pdata_42_;
input pinreg_3_;
input poutreg_57_;
input pdata_5_;
input pdata_27_;
input pdata_34_;
input pdata_41_;
input pinreg_2_;
input poutreg_58_;
input pd_20_;
input pdata_17_;
input pdata_40_;
input pinreg_9_;
input poutreg_0_;
input poutreg_33_;
input poutreg_46_;
input pc_20_;
input pd_10_;
input pdata_18_;
input pinreg_8_;
input poutreg_1_;
input poutreg_34_;
input poutreg_45_;
input preset_0_;
input pc_21_;
input pd_11_;
input pd_22_;
input pdata_15_;
input pinreg_7_;
input poutreg_31_;
input poutreg_48_;
input pc_22_;
input pd_12_;
input pd_21_;
input pdata_16_;
input pdata_30_;
input pinreg_6_;
input poutreg_32_;
input poutreg_47_;
input pc_12_;
input pdata_13_;
input poutreg_19_;
input poutreg_37_;
input poutreg_42_;
input poutreg_60_;
input pc_11_;
input pdata_14_;
input poutreg_38_;
input poutreg_41_;
input pc_10_;
input pdata_11_;
input pdata_20_;
input poutreg_35_;
input poutreg_44_;
input pdata_12_;
input poutreg_29_;
input poutreg_36_;
input poutreg_43_;
input poutreg_50_;
input pc_9_;
input pc_16_;
input pc_27_;
input pd_8_;
input pd_17_;
input pdata_in_4_;
input pinreg_30_;
input pinreg_41_;
input pinreg_52_;
input poutreg_8_;
input poutreg_15_;
input poutreg_28_;
input pc_15_;
input pd_9_;
input pd_18_;
input pd_27_;
input pdata_in_3_;
input pinreg_31_;
input pinreg_40_;
input pinreg_53_;
input poutreg_9_;
input poutreg_16_;
input poutreg_27_;
input pc_14_;
input pd_19_;
input pdata_60_;
input pdata_in_6_;
input pinreg_32_;
input pinreg_43_;
input pinreg_50_;
input poutreg_6_;
input poutreg_17_;
input poutreg_26_;
input poutreg_39_;
input pc_13_;
input pdata_in_5_;
input pinreg_33_;
input pinreg_42_;
input pinreg_51_;
input poutreg_7_;
input poutreg_18_;
input poutreg_25_;
input pc_5_;
input pc_23_;
input pd_4_;
input pd_13_;
input pd_24_;
input pinreg_12_;
input pinreg_23_;
input poutreg_4_;
input poutreg_11_;
input poutreg_24_;
input pc_6_;
input pc_19_;
input pc_24_;
input pd_5_;
input pd_14_;
input pd_23_;
input pdata_50_;
input pdata_in_7_;
input pencrypt_0_;
input pinreg_13_;
input pinreg_22_;
input poutreg_5_;
input poutreg_12_;
input poutreg_23_;
input poutreg_49_;
input pc_7_;
input pc_18_;
input pc_25_;
input pd_6_;
input pd_15_;
input pd_26_;
input pdata_19_;
input pinreg_10_;
input pinreg_21_;
input pload_key_0_;
input poutreg_2_;
input poutreg_13_;
input poutreg_22_;
input pc_8_;
input pc_17_;
input pc_26_;
input pd_7_;
input pd_16_;
input pd_25_;
input pinreg_11_;
input pinreg_20_;
input poutreg_3_;
input poutreg_14_;
input poutreg_21_;
input pc_1_;
input pd_0_;
input pdata_2_;
input pdata_53_;
input pinreg_16_;
input pinreg_27_;
input pinreg_38_;
input pinreg_49_;
input poutreg_20_;
input poutreg_59_;
input pc_2_;
input pd_1_;
input pdata_3_;
input pdata_29_;
input pdata_54_;
input pinreg_17_;
input pinreg_26_;
input pinreg_39_;
input pinreg_48_;
input pc_3_;
input pd_2_;
input pdata_0_;
input pdata_51_;
input pinreg_14_;
input pinreg_25_;
input pc_4_;
input pd_3_;
input pdata_1_;
input pdata_52_;
input pencrypt_mode_0_;
input pinreg_15_;
input pinreg_24_;
input poutreg_10_;
input pdata_39_;
input pdata_57_;
input pdata_62_;
input pdata_in_0_;
input pinreg_34_;
input pinreg_45_;
input pdata_58_;
input pdata_61_;
input pinreg_35_;
input pinreg_44_;
input pdata_55_;
input pdata_in_2_;
input pinreg_18_;
input pinreg_29_;
input pinreg_36_;
input pinreg_47_;
input pinreg_54_;
input pc_0_;
input pdata_49_;
input pdata_56_;
input pdata_63_;
input pdata_in_1_;
input pinreg_19_;
input pinreg_28_;
input pinreg_37_;
input pinreg_46_;
input pinreg_55_;
output pc_new_6_;
output pc_new_19_;
output pd_new_5_;
output pdata_new_14_;
output pdata_new_27_;
output pinreg_new_6_;
output pinreg_new_19_;
output poutreg_new_9_;
output pc_new_7_;
output pd_new_6_;
output pd_new_19_;
output pdata_new_13_;
output pdata_new_28_;
output pdata_new_39_;
output pinreg_new_5_;
output pinreg_new_18_;
output poutreg_new_19_;
output pc_new_4_;
output pd_new_3_;
output pdata_new_9_;
output pdata_new_12_;
output pdata_new_25_;
output pinreg_new_8_;
output pinreg_new_17_;
output poutreg_new_7_;
output pc_new_5_;
output pd_new_4_;
output pdata_new_11_;
output pdata_new_26_;
output pinreg_new_7_;
output pinreg_new_16_;
output poutreg_new_8_;
output pc_new_2_;
output pd_new_1_;
output pdata_new_10_;
output pdata_new_36_;
output pinreg_new_2_;
output pinreg_new_15_;
output poutreg_new_16_;
output pc_new_3_;
output pd_new_2_;
output pdata_new_35_;
output pinreg_new_1_;
output pinreg_new_14_;
output poutreg_new_15_;
output pc_new_0_;
output pdata_new_29_;
output pdata_new_38_;
output pinreg_new_4_;
output pinreg_new_13_;
output poutreg_new_18_;
output pc_new_1_;
output pd_new_0_;
output pdata_new_37_;
output pinreg_new_3_;
output pinreg_new_12_;
output poutreg_new_17_;
output pc_new_11_;
output pc_new_22_;
output pd_new_12_;
output pd_new_23_;
output pcount_new_0_;
output pdata_new_3_;
output pdata_new_45_;
output pdata_new_58_;
output pinreg_new_22_;
output pinreg_new_33_;
output pinreg_new_44_;
output pinreg_new_55_;
output poutreg_new_1_;
output poutreg_new_25_;
output poutreg_new_38_;
output poutreg_new_61_;
output pc_new_12_;
output pc_new_21_;
output pd_new_11_;
output pd_new_24_;
output pdata_new_4_;
output pdata_new_46_;
output pdata_new_57_;
output pinreg_new_23_;
output pinreg_new_32_;
output pinreg_new_45_;
output pinreg_new_54_;
output poutreg_new_2_;
output poutreg_new_26_;
output poutreg_new_37_;
output poutreg_new_62_;
output pc_new_13_;
output pc_new_24_;
output pd_new_14_;
output pd_new_21_;
output pcount_new_2_;
output pdata_new_1_;
output pdata_new_47_;
output pdata_new_56_;
output pinreg_new_0_;
output pinreg_new_24_;
output pinreg_new_35_;
output pinreg_new_42_;
output pinreg_new_53_;
output poutreg_new_27_;
output poutreg_new_36_;
output poutreg_new_49_;
output poutreg_new_50_;
output poutreg_new_63_;
output pc_new_14_;
output pc_new_23_;
output pd_new_13_;
output pd_new_22_;
output pcount_new_1_;
output pdata_new_2_;
output pdata_new_48_;
output pdata_new_55_;
output pinreg_new_25_;
output pinreg_new_34_;
output pinreg_new_43_;
output pinreg_new_52_;
output poutreg_new_0_;
output poutreg_new_28_;
output poutreg_new_35_;
output pc_new_15_;
output pc_new_26_;
output pd_new_16_;
output pd_new_27_;
output pdata_new_7_;
output pdata_new_49_;
output pinreg_new_26_;
output pinreg_new_37_;
output pinreg_new_48_;
output poutreg_new_5_;
output poutreg_new_29_;
output poutreg_new_47_;
output poutreg_new_52_;
output pc_new_16_;
output pc_new_25_;
output pd_new_15_;
output pcount_new_3_;
output pdata_new_8_;
output pinreg_new_27_;
output pinreg_new_36_;
output pinreg_new_49_;
output poutreg_new_6_;
output poutreg_new_48_;
output poutreg_new_51_;
output pc_new_17_;
output pd_new_18_;
output pd_new_25_;
output pdata_new_5_;
output pinreg_new_28_;
output pinreg_new_39_;
output pinreg_new_46_;
output poutreg_new_3_;
output poutreg_new_45_;
output poutreg_new_54_;
output pc_new_18_;
output pc_new_27_;
output pd_new_17_;
output pd_new_26_;
output pdata_new_6_;
output pdata_new_59_;
output pinreg_new_29_;
output pinreg_new_38_;
output pinreg_new_47_;
output poutreg_new_4_;
output poutreg_new_39_;
output poutreg_new_46_;
output poutreg_new_53_;
output poutreg_new_60_;
output pdata_new_50_;
output pdata_new_63_;
output poutreg_new_30_;
output poutreg_new_43_;
output poutreg_new_56_;
output poutreg_new_44_;
output poutreg_new_55_;
output pdata_new_61_;
output pencrypt_mode_new_0_;
output poutreg_new_41_;
output poutreg_new_58_;
output pdata_new_40_;
output pdata_new_62_;
output poutreg_new_20_;
output poutreg_new_42_;
output poutreg_new_57_;
output pdata_new_41_;
output pdata_new_54_;
output pinreg_new_40_;
output pinreg_new_51_;
output poutreg_new_21_;
output poutreg_new_34_;
output pd_new_20_;
output pdata_new_0_;
output pdata_new_42_;
output pdata_new_53_;
output pdata_new_60_;
output pinreg_new_41_;
output pinreg_new_50_;
output poutreg_new_22_;
output poutreg_new_33_;
output poutreg_new_40_;
output poutreg_new_59_;
output pc_new_20_;
output pd_new_10_;
output pdata_new_43_;
output pdata_new_52_;
output pinreg_new_20_;
output pinreg_new_31_;
output poutreg_new_23_;
output poutreg_new_32_;
output pc_new_10_;
output pdata_new_44_;
output pdata_new_51_;
output pinreg_new_21_;
output pinreg_new_30_;
output poutreg_new_24_;
output poutreg_new_31_;
output pdata_new_32_;
output pinreg_new_11_;
output poutreg_new_12_;
output pdata_new_20_;
output pdata_new_31_;
output pinreg_new_10_;
output poutreg_new_11_;
output pdata_new_34_;
output poutreg_new_14_;
output pdata_new_19_;
output pdata_new_33_;
output poutreg_new_13_;
output pd_new_9_;
output pdata_new_18_;
output pdata_new_23_;
output pdata_new_17_;
output pdata_new_24_;
output pinreg_new_9_;
output pc_new_8_;
output pd_new_7_;
output pdata_new_16_;
output pdata_new_21_;
output pdata_new_30_;
output poutreg_new_10_;
output pc_new_9_;
output pd_new_8_;
output pdata_new_15_;
output pdata_new_22_;
wire wire254;
wire n_n1327;
wire wire340;
wire wire341;
wire wire342;
wire wire343;
wire wire514;
wire wire348;
wire wire351;
wire wire352;
wire wire355;
wire wire359;
wire wire392;
wire wire362;
wire wire364;
wire wire366;
wire wire367;
wire wire368;
wire wire369;
wire wire370;
wire wire371;
wire wire577;
wire n_n1709;
wire n_n1710;
wire n_n1712;
wire n_n1708;
wire n_n1707;
wire n_n1696;
wire n_n1699;
wire n_n1700;
wire n_n1695;
wire n_n1715;
wire n_n1714;
wire n_n1716;
wire n_n1713;
wire n_n1718;
wire n_n1723;
wire n_n1724;
wire n_n1720;
wire n_n1719;
wire n_n1726;
wire n_n1728;
wire n_n1725;
wire n_n1730;
wire n_n1697;
wire n_n1702;
wire n_n1704;
wire n_n1706;
wire n_n1329;
wire wire616;
wire n_n1684;
wire n_n1686;
wire n_n1727;
wire n_n1705;
wire n_n1701;
wire wire264;
wire wire275;
wire wire325;
wire wire465;
wire wire512;
wire wire568;
wire wire594;
wire n_n1711;
wire n_n1703;
wire n_n1690;
wire n_n1722;
wire n_n1687;
wire n_n1688;
wire n_n1683;
wire n_n1685;
wire n_n1698;
wire n_n1721;
wire n_n1729;
wire n_n1717;
wire wire462;
wire wire620;
wire n_n1753;
wire n_n1694;
wire wire333;
wire wire393;
wire wire423;
wire wire592;
wire wire626;
wire n_n1736;
wire wire280;
wire wire297;
wire wire396;
wire wire424;
wire wire470;
wire wire475;
wire wire531;
wire n_n1691;
wire n_n1693;
wire n_n1692;
wire wire247;
wire wire270;
wire wire323;
wire wire328;
wire wire398;
wire wire507;
wire wire525;
wire wire537;
wire wire630;
wire n_n1689;
wire wire277;
wire wire467;
wire wire471;
wire wire634;
wire wire632;
wire wire631;
wire wire307;
wire wire463;
wire wire636;
wire n_n1742;
wire wire278;
wire wire306;
wire wire315;
wire wire472;
wire wire518;
wire wire335;
wire wire401;
wire wire402;
wire wire417;
wire wire529;
wire wire541;
wire wire584;
wire wire646;
wire wire645;
wire wire289;
wire wire336;
wire wire485;
wire wire552;
wire wire321;
wire wire322;
wire wire405;
wire wire523;
wire wire533;
wire wire606;
wire wire312;
wire wire431;
wire wire508;
wire wire549;
wire wire654;
wire wire653;
wire wire245;
wire wire305;
wire wire313;
wire wire324;
wire wire407;
wire wire517;
wire wire528;
wire wire655;
wire wire496;
wire n_n1758;
wire wire662;
wire wire268;
wire wire320;
wire wire664;
wire wire669;
wire wire666;
wire wire279;
wire wire309;
wire wire380;
wire wire409;
wire wire432;
wire wire468;
wire wire476;
wire wire574;
wire wire673;
wire wire672;
wire wire263;
wire wire285;
wire wire286;
wire wire331;
wire wire678;
wire wire677;
wire wire284;
wire wire379;
wire wire411;
wire wire505;
wire wire540;
wire wire680;
wire wire273;
wire wire274;
wire wire469;
wire wire558;
wire wire684;
wire wire683;
wire wire316;
wire wire338;
wire wire439;
wire wire506;
wire wire543;
wire wire588;
wire wire283;
wire wire304;
wire wire420;
wire wire504;
wire wire579;
wire wire310;
wire wire433;
wire wire534;
wire wire535;
wire wire689;
wire wire688;
wire wire246;
wire wire271;
wire wire585;
wire wire692;
wire wire691;
wire wire267;
wire wire473;
wire wire696;
wire n_n1731;
wire wire302;
wire wire426;
wire wire474;
wire wire503;
wire wire526;
wire wire536;
wire n_n1737;
wire wire265;
wire wire381;
wire wire701;
wire wire700;
wire wire301;
wire wire308;
wire wire524;
wire wire546;
wire wire477;
wire wire582;
wire wire705;
wire wire295;
wire wire413;
wire wire708;
wire wire559;
wire wire710;
wire wire709;
wire wire509;
wire wire516;
wire wire261;
wire wire262;
wire wire532;
wire wire598;
wire wire519;
wire wire269;
wire wire515;
wire wire480;
wire wire481;
wire wire555;
wire wire513;
wire wire595;
wire wire712;
wire wire713;
wire wire303;
wire wire510;
wire wire715;
wire wire714;
wire wire716;
wire wire586;
wire wire294;
wire wire604;
wire wire562;
wire wire319;
wire wire717;
wire wire718;
wire wire539;
wire wire719;
wire wire520;
wire wire527;
wire wire427;
wire wire725;
wire wire726;
wire wire484;
wire wire729;
wire wire428;
wire wire732;
wire wire569;
wire wire567;
wire wire734;
wire wire735;
wire wire736;
wire wire737;
wire wire738;
wire wire740;
wire wire739;
wire wire742;
wire wire743;
wire wire745;
wire wire744;
wire wire747;
wire wire749;
wire wire751;
wire wire750;
wire wire511;
wire wire591;
wire wire603;
wire wire619;
wire wire618;
wire wire624;
wire wire623;
wire wire635;
wire wire639;
wire wire638;
wire wire643;
wire wire650;
wire wire649;
wire wire663;
wire wire667;
wire wire670;
wire wire676;
wire wire682;
wire wire687;
wire wire697;
wire wire706;
wire wire722;
wire wire724;
wire wire327;
wire wire329;
wire wire330;
wire wire332;
wire wire339;
wire wire374;
wire wire376;
wire wire377;
wire wire378;
wire wire382;
wire wire383;
wire wire384;
wire wire404;
wire wire414;
wire wire415;
wire wire416;
wire wire418;
wire wire419;
wire wire422;
wire wire425;
wire wire429;
wire wire430;
wire wire435;
wire wire436;
wire wire451;
wire wire452;
wire wire453;
wire wire454;
wire wire455;
wire wire456;
wire wire492;
wire wire756;
wire wire770;
wire wire771;
wire wire772;
wire wire773;
wire wire774;
wire wire775;
wire wire787;
wire wire791;
wire wire792;
wire wire793;
wire wire794;
wire wire795;
wire wire796;
wire wire798;
wire wire799;
wire wire800;
wire wire801;
wire wire802;
wire wire803;
wire wire810;
wire wire820;
wire wire824;
wire wire825;
wire wire827;
wire wire828;
wire wire831;
wire wire833;
wire wire835;
wire wire836;
wire wire842;
wire wire846;
wire wire847;
wire wire848;
wire wire849;
wire wire850;
wire wire851;
wire wire862;
wire wire863;
wire wire866;
wire wire883;
wire wire889;
wire wire892;
wire wire894;
wire wire904;
wire wire905;
wire wire908;
wire wire909;
wire wire934;
wire wire935;
wire wire937;
wire wire944;
wire wire954;
wire wire955;
wire wire956;
wire wire957;
wire wire958;
wire wire962;
wire wire963;
wire wire964;
wire wire975;
wire wire976;
wire wire977;
wire wire995;
wire wire1000;
wire wire1001;
wire wire1002;
wire wire1004;
wire wire1005;
wire wire1012;
wire wire1021;
wire wire1025;
wire wire1047;
wire wire1049;
wire wire1050;
wire wire1056;
wire wire1057;
wire wire1062;
wire wire1063;
wire wire1064;
wire wire1065;
wire wire1066;
wire wire1067;
wire wire1069;
wire wire1070;
wire wire1071;
wire wire1072;
wire wire1073;
wire wire1074;
wire wire1076;
wire wire1077;
wire wire1078;
wire wire1079;
wire wire1080;
wire wire1081;
wire wire1083;
wire wire1084;
wire wire1085;
wire wire1086;
wire wire1087;
wire wire1088;
wire wire1093;
wire wire1098;
wire wire1099;
wire wire1101;
wire wire1102;
wire wire1111;
wire wire1112;
wire wire1113;
wire wire1114;
wire wire1126;
wire wire1127;
wire wire1128;
wire wire1129;
wire wire1130;
wire wire1131;
wire wire1133;
wire wire1134;
wire wire1135;
wire wire1136;
wire wire1137;
wire wire1138;
wire wire1140;
wire wire1141;
wire wire1142;
wire wire1143;
wire wire1144;
wire wire1145;
wire wire1152;
wire wire1156;
wire wire1180;
wire wire1181;
wire wire1182;
wire wire1184;
wire wire1185;
wire wire1186;
wire wire1187;
wire wire1188;
wire wire1189;
wire wire1191;
wire wire1192;
wire wire1193;
wire wire1194;
wire wire1195;
wire wire1196;
wire wire1198;
wire wire1199;
wire wire1200;
wire wire1201;
wire wire1202;
wire wire1203;
wire wire1211;
wire wire1216;
wire wire1220;
wire wire1221;
wire wire1222;
wire wire1229;
wire wire1238;
wire wire1242;
wire wire1243;
wire wire1244;
wire wire1245;
wire wire1246;
wire wire1249;
wire wire1250;
wire wire1253;
wire wire1254;
wire wire1257;
wire wire1258;
wire wire1259;
wire wire1260;
wire wire1261;
wire wire1262;
wire wire1264;
wire wire1265;
wire wire1266;
wire wire1267;
wire wire1268;
wire wire1269;
wire wire1271;
wire wire1272;
wire wire1273;
wire wire1274;
wire wire1275;
wire wire1276;
wire wire1278;
wire wire1279;
wire wire1280;
wire wire1281;
wire wire1282;
wire wire1283;
wire wire1291;
wire wire1301;
wire wire1319;
wire wire1324;
wire wire1325;
wire wire1326;
wire wire1327;
wire wire1331;
wire wire1341;
wire wire1342;
wire wire1343;
wire wire1344;
wire wire1345;
wire wire1346;
wire wire1348;
wire wire1349;
wire wire1350;
wire wire1351;
wire wire1352;
wire wire1353;
wire wire1355;
wire wire1356;
wire wire1357;
wire wire1358;
wire wire1359;
wire wire1360;
wire wire1362;
wire wire1363;
wire wire1364;
wire wire1365;
wire wire1366;
wire wire1367;
wire wire1380;
wire wire1383;
wire wire1384;
wire wire1385;
wire wire1386;
wire wire1389;
wire wire1390;
wire wire1391;
wire wire1392;
wire wire1397;
wire wire1399;
wire wire1411;
wire wire1412;
wire wire1413;
wire wire1418;
wire wire1420;
wire wire1421;
wire wire1425;
wire wire1426;
wire wire1427;
wire wire1428;
wire wire1429;
wire wire1430;
wire wire1434;
wire wire1435;
wire wire1436;
wire wire1437;
wire wire1438;
wire wire1439;
wire wire1440;
wire wire1441;
wire wire1442;
wire wire1443;
wire wire1444;
wire wire1445;
wire wire1446;
wire wire1447;
wire wire1474;
wire wire1475;
wire wire1476;
wire wire1477;
wire wire1478;
wire wire1483;
wire wire1484;
wire wire1494;
wire wire1495;
wire wire1496;
wire wire1498;
wire wire1501;
wire wire1503;
wire wire1505;
wire wire1508;
wire wire1509;
wire wire1510;
wire wire1519;
wire wire1521;
wire wire1522;
wire wire1523;
wire wire1524;
wire wire1525;
wire wire1526;
wire wire1528;
wire wire1529;
wire wire1530;
wire wire1531;
wire wire1532;
wire wire1533;
wire wire1535;
wire wire1536;
wire wire1537;
wire wire1538;
wire wire1539;
wire wire1540;
wire wire1542;
wire wire1543;
wire wire1544;
wire wire1545;
wire wire1546;
wire wire1547;
wire wire1556;
wire wire1559;
wire wire1560;
wire wire1561;
wire wire1562;
wire wire1574;
wire wire1576;
wire wire1597;
wire wire1598;
wire wire1599;
wire wire1600;
wire wire1601;
wire wire1602;
wire wire1607;
wire wire1617;
wire wire1618;
wire wire1619;
wire wire1620;
wire wire1621;
wire wire1625;
wire wire1626;
wire wire1630;
wire wire1631;
wire wire1632;
wire wire1633;
wire wire1634;
wire wire1647;
wire wire1651;
wire wire1652;
wire wire1653;
wire wire1654;
wire wire1655;
wire wire1656;
wire wire1657;
wire wire1659;
wire wire1660;
wire wire1666;
wire wire1667;
wire wire1668;
wire wire1669;
wire wire1670;
wire wire1671;
wire wire1673;
wire wire1674;
wire wire1675;
wire wire1676;
wire wire1677;
wire wire1678;
wire wire1680;
wire wire1681;
wire wire1682;
wire wire1683;
wire wire1684;
wire wire1685;
wire wire1687;
wire wire1688;
wire wire1689;
wire wire1690;
wire wire1691;
wire wire1692;
wire wire1695;
wire wire1698;
wire wire1699;
wire wire1704;
wire wire1705;
wire wire1706;
wire wire1707;
wire wire1708;
wire wire1709;
wire wire1714;
wire wire1716;
wire wire1723;
wire wire1741;
wire wire1742;
wire wire1744;
wire wire1745;
wire wire1746;
wire wire1747;
wire wire1753;
wire wire1754;
wire wire1756;
wire wire1758;
wire wire1759;
wire wire1760;
wire wire1761;
wire wire1766;
wire wire1767;
wire wire1768;
wire wire1769;
wire wire1770;
wire wire1771;
wire wire1773;
wire wire1774;
wire wire1775;
wire wire1776;
wire wire1777;
wire wire1778;
wire wire1780;
wire wire1781;
wire wire1782;
wire wire1783;
wire wire1784;
wire wire1785;
wire wire1787;
wire wire1788;
wire wire1789;
wire wire1790;
wire wire1791;
wire wire1792;
wire wire1805;
wire wire1806;
wire wire1807;
wire wire1808;
wire wire1809;
wire wire1810;
wire wire1813;
wire wire1814;
wire wire1815;
wire wire1816;
wire wire1817;
wire wire1818;
wire wire1819;
wire wire1829;
wire wire1830;
wire wire1834;
wire wire1835;
wire wire1836;
wire wire1837;
wire wire1838;
wire wire1839;
wire wire1841;
wire wire1842;
wire wire1857;
wire wire1858;
wire wire1859;
wire wire1860;
wire wire1861;
wire wire1862;
wire wire1864;
wire wire1865;
wire wire1866;
wire wire1867;
wire wire1868;
wire wire1869;
wire wire1882;
wire wire1883;
wire wire1884;
wire wire1885;
wire wire1886;
wire wire1887;
wire wire1894;
wire wire1895;
wire wire1896;
wire wire1897;
wire wire1902;
wire wire1903;
wire wire1904;
wire wire1905;
wire wire1906;
wire wire1913;
wire wire1914;
wire wire1917;
wire wire1918;
wire wire1919;
wire wire1920;
wire wire1921;
wire wire1922;
wire wire1923;
wire wire1925;
wire wire1929;
wire wire1930;
wire wire1949;
wire wire1953;
wire wire1955;
wire wire1956;
wire wire1962;
wire wire1964;
wire wire1969;
wire wire1970;
wire wire1973;
wire wire1977;
wire wire1978;
wire wire1979;
wire wire1980;
wire wire1981;
wire wire1982;
wire wire1983;
wire wire1996;
wire wire1997;
wire wire1998;
wire wire1999;
wire wire2000;
wire wire2001;
wire wire2003;
wire wire2004;
wire wire2005;
wire wire2006;
wire wire2007;
wire wire2008;
wire wire2017;
wire wire2021;
wire wire2022;
wire wire2023;
wire wire2025;
wire wire2026;
wire wire2027;
wire wire2032;
wire wire2033;
wire wire2034;
wire wire2035;
wire wire2036;
wire wire2037;
wire wire2038;
wire wire2039;
wire wire2040;
wire wire2041;
wire wire2044;
wire wire2046;
wire wire2048;
wire wire2049;
wire wire2050;
wire wire2051;
wire wire2066;
wire wire2067;
wire wire2068;
wire wire2069;
wire wire2070;
wire wire2071;
wire wire2073;
wire wire2074;
wire wire2075;
wire wire2076;
wire wire2077;
wire wire2078;
wire wire2091;
wire wire2092;
wire wire2093;
wire wire2094;
wire wire2095;
wire wire2096;
wire wire2098;
wire wire2099;
wire wire2100;
wire wire2101;
wire wire2102;
wire wire2103;
wire wire2110;
wire wire2111;
wire wire2112;
wire wire2113;
wire wire2123;
wire wire2124;
wire wire2125;
wire wire2127;
wire wire2143;
wire wire2144;
wire wire2145;
wire wire2146;
wire wire2147;
wire wire2148;
wire wire2150;
wire wire2151;
wire wire2152;
wire wire2153;
wire wire2154;
wire wire2155;
wire wire2162;
wire wire2167;
wire wire2169;
wire wire2175;
wire wire2182;
wire wire2184;
wire wire2195;
wire wire2198;
wire wire2202;
wire wire2208;
wire wire2209;
wire wire2210;
wire wire2211;
wire wire2212;
wire wire2214;
wire wire2218;
wire wire2219;
wire wire2222;
wire wire2223;
wire wire2224;
wire wire2225;
wire wire2227;
wire wire2228;
wire wire2231;
wire wire2232;
wire wire2249;
wire wire2250;
wire wire2251;
wire wire2252;
wire wire2253;
wire wire2254;
wire wire2256;
wire wire2257;
wire wire2258;
wire wire2259;
wire wire2260;
wire wire2261;
wire wire2263;
wire wire2264;
wire wire2265;
wire wire2266;
wire wire2267;
wire wire2268;
wire wire2275;
wire wire2276;
wire wire2277;
wire wire2278;
wire wire2293;
wire wire2294;
wire wire2295;
wire wire2304;
wire wire2306;
wire wire2309;
wire wire2311;
wire wire2334;
wire wire2335;
wire wire2336;
wire wire2337;
wire wire2338;
wire wire2339;
wire wire2341;
wire wire2342;
wire wire2343;
wire wire2344;
wire wire2345;
wire wire2346;
wire wire2348;
wire wire2349;
wire wire2350;
wire wire2351;
wire wire2352;
wire wire2353;
wire wire7710;
wire wire7711;
wire wire7712;
wire wire7714;
wire wire7717;
wire wire7719;
wire wire7722;
wire wire7724;
wire wire7727;
wire wire7729;
wire wire7731;
wire wire7732;
wire wire7733;
wire wire7738;
wire wire7741;
wire wire7744;
wire wire7745;
wire wire7747;
wire wire7748;
wire wire7751;
wire wire7752;
wire wire7753;
wire wire7755;
wire wire7757;
wire wire7760;
wire wire7762;
wire wire7765;
wire wire7767;
wire wire7770;
wire wire7771;
wire wire7772;
wire wire7775;
wire wire7776;
wire wire7783;
wire wire7785;
wire wire7786;
wire wire7787;
wire wire7791;
wire wire7793;
wire wire7794;
wire wire7795;
wire wire7799;
wire wire7800;
wire wire7802;
wire wire7805;
wire wire7807;
wire wire7810;
wire wire7816;
wire wire7819;
wire wire7820;
wire wire7822;
wire wire7825;
wire wire7827;
wire wire7830;
wire wire7831;
wire wire7833;
wire wire7836;
wire wire7838;
wire wire7841;
wire wire7844;
wire wire7845;
wire wire7846;
wire wire7850;
wire wire7852;
wire wire7853;
wire wire7856;
wire wire7857;
wire wire7860;
wire wire7863;
wire wire7865;
wire wire7866;
wire wire7867;
wire wire7871;
wire wire7872;
wire wire7873;
wire wire7875;
wire wire7878;
wire wire7880;
wire wire7883;
wire wire7884;
wire wire7894;
wire wire7898;
wire wire7900;
wire wire7901;
wire wire7902;
wire wire7905;
wire wire7908;
wire wire7912;
wire wire7919;
wire wire7920;
wire wire7923;
wire wire7925;
wire wire7928;
wire wire7929;
wire wire7931;
wire wire7934;
wire wire7936;
wire wire7939;
wire wire7943;
wire wire7946;
wire wire7948;
wire wire7949;
wire wire7952;
wire wire7953;
wire wire7960;
wire wire7962;
wire wire7966;
wire wire7967;
wire wire7969;
wire wire7971;
wire wire7974;
wire wire7976;
wire wire7979;
wire wire7981;
wire wire7984;
wire wire7986;
wire wire7989;
wire wire7996;
wire wire8000;
wire wire8001;
wire wire8004;
wire wire8005;
wire wire8006;
wire wire8008;
wire wire8009;
wire wire8010;
wire wire8013;
wire wire8018;
wire wire8019;
wire wire8023;
wire wire8026;
wire wire8028;
wire wire8031;
wire wire8033;
wire wire8036;
wire wire8038;
wire wire8041;
wire wire8047;
wire wire8048;
wire wire8049;
wire wire8053;
wire wire8054;
wire wire8055;
wire wire8057;
wire wire8058;
wire wire8060;
wire wire8062;
wire wire8063;
wire wire8066;
wire wire8067;
wire wire8074;
wire wire8075;
wire wire8077;
wire wire8078;
wire wire8080;
wire wire8081;
wire wire8084;
wire wire8088;
wire wire8089;
wire wire8091;
wire wire8092;
wire wire8096;
wire wire8097;
wire wire8099;
wire wire8102;
wire wire8104;
wire wire8107;
wire wire8109;
wire wire8112;
wire wire8114;
wire wire8117;
wire wire8125;
wire wire8130;
wire wire8131;
wire wire8134;
wire wire8138;
wire wire8139;
wire wire8140;
wire wire8143;
wire wire8144;
wire wire8150;
wire wire8153;
wire wire8154;
wire wire8155;
wire wire8160;
wire wire8162;
wire wire8163;
wire wire8165;
wire wire8166;
wire wire8168;
wire wire8169;
wire wire8170;
wire wire8175;
wire wire8176;
wire wire8178;
wire wire8179;
wire wire8181;
wire wire8184;
wire wire8186;
wire wire8189;
wire wire8191;
wire wire8194;
wire wire8196;
wire wire8199;
wire wire8202;
wire wire8204;
wire wire8206;
wire wire8207;
wire wire8210;
wire wire8211;
wire wire8212;
wire wire8215;
wire wire8217;
wire wire8218;
wire wire8219;
wire wire8221;
wire wire8223;
wire wire8226;
wire wire8228;
wire wire8231;
wire wire8233;
wire wire8236;
wire wire8238;
wire wire8241;
wire wire8245;
wire wire8246;
wire wire8247;
wire wire8250;
wire wire8253;
wire wire8254;
wire wire8258;
wire wire8259;
wire wire8263;
wire wire8264;
wire wire8265;
wire wire8266;
wire wire8267;
wire wire8268;
wire wire8270;
wire wire8273;
wire wire8275;
wire wire8278;
wire wire8280;
wire wire8283;
wire wire8284;
wire wire8285;
wire wire8289;
wire wire8290;
wire wire8291;
wire wire8293;
wire wire8294;
wire wire8296;
wire wire8298;
wire wire8301;
wire wire8303;
wire wire8306;
wire wire8308;
wire wire8311;
wire wire8312;
wire wire8319;
wire wire8320;
wire wire8322;
wire wire8323;
wire wire8326;
wire wire8327;
wire wire8328;
wire wire8330;
wire wire8333;
wire wire8335;
wire wire8338;
wire wire8340;
wire wire8343;
wire wire8345;
wire wire8348;
wire wire8350;
wire wire8352;
wire wire8353;
wire wire8355;
wire wire8356;
wire wire8358;
wire wire8359;
wire wire8360;
wire wire8361;
wire wire8362;
wire wire8364;
wire wire8367;
wire wire8370;
wire wire8371;
wire wire8374;
wire wire8375;
wire wire8376;
wire wire8377;
wire wire8378;
wire wire8382;
wire wire8383;
wire wire8385;
wire wire8389;
wire wire8393;
wire wire8396;
wire wire8397;
wire wire8400;
wire wire8402;
wire wire8403;
wire wire8404;
wire wire8406;
wire wire8407;
wire wire8413;
wire wire8414;
wire wire8416;
wire wire8417;
wire wire8418;
wire wire8420;
wire wire8421;
wire wire8423;
wire wire8424;
wire wire8428;
wire wire8429;
wire wire8432;
wire wire8433;
wire wire8435;
wire wire8437;
wire wire8439;
wire wire8440;
wire wire8441;
wire wire8443;
wire wire8444;
wire wire8446;
wire wire8449;
wire wire8457;
wire wire8459;
wire wire8460;
wire wire8461;
wire wire8462;
wire wire8464;
wire wire8467;
wire wire8469;
wire wire8472;
wire wire8473;
wire wire8474;
wire wire8476;
wire wire8479;
wire wire8480;
wire wire8481;
wire wire8482;
wire wire8483;
wire wire8484;
wire wire8485;
wire wire8487;
wire wire8490;
wire wire8492;
wire wire8495;
wire wire8497;
wire wire8500;
wire wire8501;
wire wire8503;
wire wire8506;
wire wire8508;
wire wire8511;
assign pc_new_6_ = ( wire2350 ) | ( wire2351 ) | ( wire7717 ) ;
 assign pc_new_19_ = ( wire2343 ) | ( wire2344 ) | ( wire7722 ) ;
 assign pd_new_5_ = ( wire2336 ) | ( wire2337 ) | ( wire7727 ) ;
 assign pdata_new_14_ = ( pinreg_3_  &  n_n1327 ) | ( pdata_46_  &  (~ n_n1327) ) ;
 assign pdata_new_27_ = ( pinreg_31_  &  n_n1327 ) | ( pdata_59_  &  (~ n_n1327) ) ;
 assign pinreg_new_6_ = ( (~ pcount_0_)  &  pinreg_6_ ) | ( pcount_0_  &  pdata_in_6_  &  (~ wire577) ) ;
 assign pinreg_new_19_ = ( (~ pcount_0_)  &  pinreg_19_ ) | ( pcount_0_  &  pinreg_11_  &  (~ wire577) ) ;
 assign poutreg_new_9_ = ( wire7755 ) | ( n_n1327  &  wire340 ) ;
 assign pc_new_7_ = ( wire2265 ) | ( wire2266 ) | ( wire7760 ) ;
 assign pd_new_6_ = ( wire2258 ) | ( wire2259 ) | ( wire7765 ) ;
 assign pd_new_19_ = ( wire2251 ) | ( wire2252 ) | ( wire7770 ) ;
 assign pdata_new_13_ = ( pinreg_11_  &  n_n1327 ) | ( pdata_45_  &  (~ n_n1327) ) ;
 assign pdata_new_28_ = ( pinreg_23_  &  n_n1327 ) | ( pdata_60_  &  (~ n_n1327) ) ;
 assign pdata_new_39_ = ( pdata_in_0_  &  n_n1327 ) | ( (~ n_n1327)  &  wire341 ) ;
 assign pinreg_new_5_ = ( (~ pcount_0_)  &  pinreg_5_ ) | ( pcount_0_  &  pdata_in_5_  &  (~ wire577) ) ;
 assign pinreg_new_18_ = ( (~ pcount_0_)  &  pinreg_18_ ) | ( pcount_0_  &  pinreg_10_  &  (~ wire577) ) ;
 assign poutreg_new_19_ = ( wire7800 ) | ( n_n1327  &  wire342 ) ;
 assign pc_new_4_ = ( wire2152 ) | ( wire2153 ) | ( wire7805 ) ;
 assign pd_new_3_ = ( wire2145 ) | ( wire2146 ) | ( wire7810 ) ;
 assign pdata_new_9_ = ( pinreg_43_  &  n_n1327 ) | ( pdata_41_  &  (~ n_n1327) ) ;
 assign pdata_new_12_ = ( pinreg_19_  &  n_n1327 ) | ( pdata_44_  &  (~ n_n1327) ) ;
 assign pdata_new_25_ = ( pinreg_47_  &  n_n1327 ) | ( pdata_57_  &  (~ n_n1327) ) ;
 assign pinreg_new_8_ = ( (~ pcount_0_)  &  pinreg_8_ ) | ( pinreg_0_  &  pcount_0_  &  (~ wire577) ) ;
 assign pinreg_new_17_ = ( (~ pcount_0_)  &  pinreg_17_ ) | ( pcount_0_  &  pinreg_9_  &  (~ wire577) ) ;
 assign poutreg_new_7_ = ( wire7820 ) | ( n_n1327  &  wire343 ) ;
 assign pc_new_5_ = ( wire2100 ) | ( wire2101 ) | ( wire7825 ) ;
 assign pd_new_4_ = ( wire2093 ) | ( wire2094 ) | ( wire7830 ) ;
 assign pdata_new_11_ = ( pinreg_27_  &  n_n1327 ) | ( pdata_43_  &  (~ n_n1327) ) ;
 assign pdata_new_26_ = ( pinreg_39_  &  n_n1327 ) | ( pdata_58_  &  (~ n_n1327) ) ;
 assign pinreg_new_7_ = ( (~ pcount_0_)  &  pinreg_7_ ) | ( pcount_0_  &  pdata_in_7_  &  (~ wire577) ) ;
 assign pinreg_new_16_ = ( (~ pcount_0_)  &  pinreg_16_ ) | ( pcount_0_  &  pinreg_8_  &  (~ wire577) ) ;
 assign poutreg_new_8_ = ( wire7831 ) | ( (~ pcount_0_)  &  poutreg_8_ ) ;
 assign pc_new_2_ = ( wire2075 ) | ( wire2076 ) | ( wire7836 ) ;
 assign pd_new_1_ = ( wire2068 ) | ( wire2069 ) | ( wire7841 ) ;
 assign pdata_new_10_ = ( pinreg_35_  &  n_n1327 ) | ( pdata_42_  &  (~ n_n1327) ) ;
 assign pdata_new_36_ = ( wire2017 ) | ( pinreg_16_  &  n_n1327 ) ;
 assign pinreg_new_2_ = ( (~ pcount_0_)  &  pinreg_2_ ) | ( pcount_0_  &  pdata_in_2_  &  (~ wire577) ) ;
 assign pinreg_new_15_ = ( (~ pcount_0_)  &  pinreg_15_ ) | ( pcount_0_  &  pinreg_7_  &  (~ wire577) ) ;
 assign poutreg_new_16_ = ( wire7873 ) | ( (~ pcount_0_)  &  poutreg_16_ ) ;
 assign pc_new_3_ = ( wire2005 ) | ( wire2006 ) | ( wire7878 ) ;
 assign pd_new_2_ = ( wire1998 ) | ( wire1999 ) | ( wire7883 ) ;
 assign pdata_new_35_ = ( wire1949 ) | ( pinreg_24_  &  n_n1327 ) ;
 assign pinreg_new_1_ = ( pinreg_1_  &  (~ pcount_0_) ) | ( pcount_0_  &  pdata_in_1_  &  (~ wire577) ) ;
 assign pinreg_new_14_ = ( (~ pcount_0_)  &  pinreg_14_ ) | ( pcount_0_  &  pinreg_6_  &  (~ wire577) ) ;
 assign poutreg_new_15_ = ( wire7923 ) | ( (~ pdata_30_)  &  n_n1327  &  n_n1736 ) | ( pdata_30_  &  n_n1327  &  (~ n_n1736) ) ;
 assign pc_new_0_ = ( wire1884 ) | ( wire1885 ) | ( wire7928 ) ;
 assign pdata_new_29_ = ( pinreg_15_  &  n_n1327 ) | ( pdata_61_  &  (~ n_n1327) ) ;
 assign pdata_new_38_ = ( pinreg_0_  &  n_n1327 ) | ( (~ n_n1327)  &  wire340 ) ;
 assign pinreg_new_4_ = ( (~ pcount_0_)  &  pinreg_4_ ) | ( pcount_0_  &  pdata_in_4_  &  (~ wire577) ) ;
 assign pinreg_new_13_ = ( (~ pcount_0_)  &  pinreg_13_ ) | ( pcount_0_  &  pinreg_5_  &  (~ wire577) ) ;
 assign poutreg_new_18_ = ( wire7929 ) | ( (~ pcount_0_)  &  poutreg_18_ ) ;
 assign pc_new_1_ = ( wire1866 ) | ( wire1867 ) | ( wire7934 ) ;
 assign pd_new_0_ = ( wire1859 ) | ( wire1860 ) | ( wire7939 ) ;
 assign pdata_new_37_ = ( pinreg_8_  &  n_n1327 ) | ( (~ pdata_5_)  &  (~ n_n1327)  &  n_n1737 ) | ( pdata_5_  &  (~ n_n1327)  &  (~ n_n1737) ) ;
 assign pinreg_new_3_ = ( (~ pcount_0_)  &  pinreg_3_ ) | ( pcount_0_  &  pdata_in_3_  &  (~ wire577) ) ;
 assign pinreg_new_12_ = ( (~ pcount_0_)  &  pinreg_12_ ) | ( pcount_0_  &  pinreg_4_  &  (~ wire577) ) ;
 assign poutreg_new_17_ = ( wire7969 ) | ( (~ pdata_5_)  &  n_n1327  &  n_n1737 ) | ( pdata_5_  &  n_n1327  &  (~ n_n1737) ) ;
 assign pc_new_11_ = ( wire1789 ) | ( wire1790 ) | ( wire7974 ) ;
 assign pc_new_22_ = ( wire1782 ) | ( wire1783 ) | ( wire7979 ) ;
 assign pd_new_12_ = ( wire1775 ) | ( wire1776 ) | ( wire7984 ) ;
 assign pd_new_23_ = ( wire1768 ) | ( wire1769 ) | ( wire7989 ) ;
 assign pcount_new_0_ = ( (~ pcount_0_)  &  (~ preset_0_) ) ;
 assign pdata_new_3_ = ( pinreg_25_  &  n_n1327 ) | ( pdata_35_  &  (~ n_n1327) ) ;
 assign pdata_new_45_ = ( pinreg_10_  &  n_n1327 ) | ( (~ n_n1327)  &  wire342 ) ;
 assign pdata_new_58_ = ( pinreg_38_  &  n_n1327 ) | ( (~ n_n1327)  &  wire348 ) ;
 assign pinreg_new_22_ = ( (~ pcount_0_)  &  pinreg_22_ ) | ( pcount_0_  &  pinreg_14_  &  (~ wire577) ) ;
 assign pinreg_new_33_ = ( (~ pcount_0_)  &  pinreg_33_ ) | ( pcount_0_  &  pinreg_25_  &  (~ wire577) ) ;
 assign pinreg_new_44_ = ( (~ pcount_0_)  &  pinreg_44_ ) | ( pcount_0_  &  pinreg_36_  &  (~ wire577) ) ;
 assign pinreg_new_55_ = ( (~ pcount_0_)  &  pinreg_55_ ) | ( pcount_0_  &  pinreg_47_  &  (~ wire577) ) ;
 assign poutreg_new_1_ = ( wire8008 ) | ( n_n1327  &  wire341 ) ;
 assign poutreg_new_25_ = ( wire1723 ) | ( wire8009 ) ;
 assign poutreg_new_38_ = ( wire8010 ) | ( (~ pcount_0_)  &  poutreg_38_ ) ;
 assign poutreg_new_61_ = ( wire1695 ) | ( (~ pdata_16_)  &  n_n1327  &  n_n1758 ) | ( pdata_16_  &  n_n1327  &  (~ n_n1758) ) ;
 assign pc_new_12_ = ( wire1689 ) | ( wire1690 ) | ( wire8026 ) ;
 assign pc_new_21_ = ( wire1682 ) | ( wire1683 ) | ( wire8031 ) ;
 assign pd_new_11_ = ( wire1675 ) | ( wire1676 ) | ( wire8036 ) ;
 assign pd_new_24_ = ( wire1668 ) | ( wire1669 ) | ( wire8041 ) ;
 assign pdata_new_4_ = ( pinreg_17_  &  n_n1327 ) | ( pdata_36_  &  (~ n_n1327) ) ;
 assign pdata_new_46_ = ( wire1647 ) | ( pinreg_2_  &  n_n1327 ) ;
 assign pdata_new_57_ = ( pinreg_46_  &  n_n1327 ) | ( (~ n_n1327)  &  wire351 ) ;
 assign pinreg_new_23_ = ( (~ pcount_0_)  &  pinreg_23_ ) | ( pcount_0_  &  pinreg_15_  &  (~ wire577) ) ;
 assign pinreg_new_32_ = ( (~ pcount_0_)  &  pinreg_32_ ) | ( pcount_0_  &  pinreg_24_  &  (~ wire577) ) ;
 assign pinreg_new_45_ = ( (~ pcount_0_)  &  pinreg_45_ ) | ( pcount_0_  &  pinreg_37_  &  (~ wire577) ) ;
 assign pinreg_new_54_ = ( (~ pcount_0_)  &  pinreg_54_ ) | ( pcount_0_  &  pinreg_46_  &  (~ wire577) ) ;
 assign poutreg_new_2_ = ( wire8080 ) | ( (~ pcount_0_)  &  poutreg_2_ ) ;
 assign poutreg_new_26_ = ( wire8081 ) | ( (~ pcount_0_)  &  poutreg_26_ ) ;
 assign poutreg_new_37_ = ( wire8097 ) | ( n_n1327  &  wire352 ) ;
 assign poutreg_new_62_ = ( poutreg_62_  &  (~ pcount_0_) ) | ( pcount_0_  &  pdata_56_  &  wire577 ) ;
 assign pc_new_13_ = ( wire1544 ) | ( wire1545 ) | ( wire8102 ) ;
 assign pc_new_24_ = ( wire1537 ) | ( wire1538 ) | ( wire8107 ) ;
 assign pd_new_14_ = ( wire1530 ) | ( wire1531 ) | ( wire8112 ) ;
 assign pd_new_21_ = ( wire1523 ) | ( wire1524 ) | ( wire8117 ) ;
 assign pcount_new_2_ = ( pcount_2_  &  (~ pcount_1_)  &  wire514 ) | ( pcount_2_  &  (~ pcount_0_)  &  wire514 ) | ( (~ pcount_2_)  &  pcount_1_  &  pcount_0_  &  wire514 ) ;
 assign pdata_new_1_ = ( pinreg_41_  &  n_n1327 ) | ( pdata_33_  &  (~ n_n1327) ) ;
 assign pdata_new_47_ = ( pdata_in_2_  &  n_n1327 ) | ( (~ pdata_15_)  &  (~ n_n1327)  &  n_n1731 ) | ( pdata_15_  &  (~ n_n1327)  &  (~ n_n1731) ) ;
 assign pdata_new_56_ = ( pinreg_54_  &  n_n1327 ) | ( (~ n_n1327)  &  wire355 ) ;
 assign pinreg_new_0_ = ( pinreg_0_  &  (~ pcount_0_) ) | ( pcount_0_  &  pdata_in_0_  &  (~ wire577) ) ;
 assign pinreg_new_24_ = ( (~ pcount_0_)  &  pinreg_24_ ) | ( pcount_0_  &  pinreg_16_  &  (~ wire577) ) ;
 assign pinreg_new_35_ = ( (~ pcount_0_)  &  pinreg_35_ ) | ( pcount_0_  &  pinreg_27_  &  (~ wire577) ) ;
 assign pinreg_new_42_ = ( (~ pcount_0_)  &  pinreg_42_ ) | ( pcount_0_  &  pinreg_34_  &  (~ wire577) ) ;
 assign pinreg_new_53_ = ( (~ pcount_0_)  &  pinreg_53_ ) | ( pcount_0_  &  pinreg_45_  &  (~ wire577) ) ;
 assign poutreg_new_27_ = ( wire8168 ) | ( (~ pdata_12_)  &  n_n1327  &  n_n1742 ) | ( pdata_12_  &  n_n1327  &  (~ n_n1742) ) ;
 assign poutreg_new_36_ = ( wire8169 ) | ( (~ pcount_0_)  &  poutreg_36_ ) ;
 assign poutreg_new_49_ = ( wire8178 ) | ( (~ pdata_1_)  &  n_n1327  &  n_n1753 ) | ( pdata_1_  &  n_n1327  &  (~ n_n1753) ) ;
 assign poutreg_new_50_ = ( wire8179 ) | ( (~ pcount_0_)  &  poutreg_50_ ) ;
 assign poutreg_new_63_ = ( poutreg_63_  &  (~ pcount_0_) ) | ( n_n1327  &  wire355 ) ;
 assign pc_new_14_ = ( wire1364 ) | ( wire1365 ) | ( wire8184 ) ;
 assign pc_new_23_ = ( wire1357 ) | ( wire1358 ) | ( wire8189 ) ;
 assign pd_new_13_ = ( wire1350 ) | ( wire1351 ) | ( wire8194 ) ;
 assign pd_new_22_ = ( wire1343 ) | ( wire1344 ) | ( wire8199 ) ;
 assign pcount_new_1_ = ( (~ pcount_1_)  &  pcount_0_  &  wire514 ) | ( pcount_1_  &  (~ pcount_0_)  &  wire514 ) ;
 assign pdata_new_2_ = ( pinreg_33_  &  n_n1327 ) | ( pdata_34_  &  (~ n_n1327) ) ;
 assign pdata_new_48_ = ( pinreg_52_  &  n_n1327 ) | ( (~ pdata_16_)  &  (~ n_n1327)  &  n_n1758 ) | ( pdata_16_  &  (~ n_n1327)  &  (~ n_n1758) ) ;
 assign pdata_new_55_ = ( wire1319 ) | ( pdata_in_4_  &  n_n1327 ) ;
 assign pinreg_new_25_ = ( (~ pcount_0_)  &  pinreg_25_ ) | ( pcount_0_  &  pinreg_17_  &  (~ wire577) ) ;
 assign pinreg_new_34_ = ( (~ pcount_0_)  &  pinreg_34_ ) | ( pcount_0_  &  pinreg_26_  &  (~ wire577) ) ;
 assign pinreg_new_43_ = ( (~ pcount_0_)  &  pinreg_43_ ) | ( pcount_0_  &  pinreg_35_  &  (~ wire577) ) ;
 assign pinreg_new_52_ = ( (~ pcount_0_)  &  pinreg_52_ ) | ( pcount_0_  &  pinreg_44_  &  (~ wire577) ) ;
 assign poutreg_new_0_ = ( wire8211 ) | ( (~ pcount_0_)  &  poutreg_0_ ) ;
 assign poutreg_new_28_ = ( wire8212 ) | ( (~ pcount_0_)  &  poutreg_28_ ) ;
 assign poutreg_new_35_ = ( wire8221 ) | ( n_n1327  &  wire359 ) ;
 assign pc_new_15_ = ( wire1280 ) | ( wire1281 ) | ( wire8226 ) ;
 assign pc_new_26_ = ( wire1273 ) | ( wire1274 ) | ( wire8231 ) ;
 assign pd_new_16_ = ( wire1266 ) | ( wire1267 ) | ( wire8236 ) ;
 assign pd_new_27_ = ( wire1259 ) | ( wire1260 ) | ( wire8241 ) ;
 assign pdata_new_7_ = ( pdata_in_1_  &  n_n1327 ) | ( pdata_39_  &  (~ n_n1327) ) ;
 assign pdata_new_49_ = ( wire1238 ) | ( pinreg_44_  &  n_n1327 ) ;
 assign pinreg_new_26_ = ( (~ pcount_0_)  &  pinreg_26_ ) | ( pcount_0_  &  pinreg_18_  &  (~ wire577) ) ;
 assign pinreg_new_37_ = ( (~ pcount_0_)  &  pinreg_37_ ) | ( pcount_0_  &  pinreg_29_  &  (~ wire577) ) ;
 assign pinreg_new_48_ = ( (~ pcount_0_)  &  pinreg_48_ ) | ( pcount_0_  &  pinreg_40_  &  (~ wire577) ) ;
 assign poutreg_new_5_ = ( wire1229 ) | ( wire8254 ) ;
 assign poutreg_new_29_ = ( wire1211 ) | ( wire8266 ) ;
 assign poutreg_new_47_ = ( wire8267 ) | ( n_n1327  &  wire348 ) ;
 assign poutreg_new_52_ = ( wire8268 ) | ( poutreg_52_  &  (~ pcount_0_) ) ;
 assign pc_new_16_ = ( wire1200 ) | ( wire1201 ) | ( wire8273 ) ;
 assign pc_new_25_ = ( wire1193 ) | ( wire1194 ) | ( wire8278 ) ;
 assign pd_new_15_ = ( wire1186 ) | ( wire1187 ) | ( wire8283 ) ;
 assign pcount_new_3_ = ( wire1180 ) | ( wire1181 ) ;
 assign pdata_new_8_ = ( pinreg_51_  &  n_n1327 ) | ( pdata_40_  &  (~ n_n1327) ) ;
 assign pinreg_new_27_ = ( (~ pcount_0_)  &  pinreg_27_ ) | ( pcount_0_  &  pinreg_19_  &  (~ wire577) ) ;
 assign pinreg_new_36_ = ( (~ pcount_0_)  &  pinreg_36_ ) | ( pcount_0_  &  pinreg_28_  &  (~ wire577) ) ;
 assign pinreg_new_49_ = ( (~ pcount_0_)  &  pinreg_49_ ) | ( pcount_0_  &  pinreg_41_  &  (~ wire577) ) ;
 assign poutreg_new_6_ = ( wire8284 ) | ( (~ pcount_0_)  &  poutreg_6_ ) ;
 assign poutreg_new_48_ = ( wire8285 ) | ( (~ pcount_0_)  &  poutreg_48_ ) ;
 assign poutreg_new_51_ = ( wire8296 ) | ( n_n1327  &  wire362 ) ;
 assign pc_new_17_ = ( wire1142 ) | ( wire1143 ) | ( wire8301 ) ;
 assign pd_new_18_ = ( wire1135 ) | ( wire1136 ) | ( wire8306 ) ;
 assign pd_new_25_ = ( wire1128 ) | ( wire1129 ) | ( wire8311 ) ;
 assign pdata_new_5_ = ( pinreg_9_  &  n_n1327 ) | ( pdata_37_  &  (~ n_n1327) ) ;
 assign pinreg_new_28_ = ( (~ pcount_0_)  &  pinreg_28_ ) | ( pcount_0_  &  pinreg_20_  &  (~ wire577) ) ;
 assign pinreg_new_39_ = ( (~ pcount_0_)  &  pinreg_39_ ) | ( pcount_0_  &  pinreg_31_  &  (~ wire577) ) ;
 assign pinreg_new_46_ = ( (~ pcount_0_)  &  pinreg_46_ ) | ( pcount_0_  &  pinreg_38_  &  (~ wire577) ) ;
 assign poutreg_new_3_ = ( wire8312 ) | ( (~ pdata_15_)  &  n_n1327  &  n_n1731 ) | ( pdata_15_  &  n_n1327  &  (~ n_n1731) ) ;
 assign poutreg_new_45_ = ( wire1093 ) | ( wire8327 ) ;
 assign poutreg_new_54_ = ( wire8328 ) | ( (~ pcount_0_)  &  poutreg_54_ ) ;
 assign pc_new_18_ = ( wire1085 ) | ( wire1086 ) | ( wire8333 ) ;
 assign pc_new_27_ = ( wire1078 ) | ( wire1079 ) | ( wire8338 ) ;
 assign pd_new_17_ = ( wire1071 ) | ( wire1072 ) | ( wire8343 ) ;
 assign pd_new_26_ = ( wire1064 ) | ( wire1065 ) | ( wire8348 ) ;
 assign pdata_new_6_ = ( pinreg_1_  &  n_n1327 ) | ( pdata_38_  &  (~ n_n1327) ) ;
 assign pdata_new_59_ = ( pinreg_30_  &  n_n1327 ) | ( (~ n_n1327)  &  wire364 ) ;
 assign pinreg_new_29_ = ( (~ pcount_0_)  &  pinreg_29_ ) | ( pcount_0_  &  pinreg_21_  &  (~ wire577) ) ;
 assign pinreg_new_38_ = ( (~ pcount_0_)  &  pinreg_38_ ) | ( pcount_0_  &  pinreg_30_  &  (~ wire577) ) ;
 assign pinreg_new_47_ = ( (~ pcount_0_)  &  pinreg_47_ ) | ( pcount_0_  &  pinreg_39_  &  (~ wire577) ) ;
 assign poutreg_new_4_ = ( wire8358 ) | ( (~ pcount_0_)  &  poutreg_4_ ) ;
 assign poutreg_new_39_ = ( wire8359 ) | ( n_n1327  &  wire364 ) ;
 assign poutreg_new_46_ = ( wire8360 ) | ( (~ pcount_0_)  &  poutreg_46_ ) ;
 assign poutreg_new_53_ = ( wire1025 ) | ( wire8361 ) ;
 assign poutreg_new_60_ = ( (~ pcount_0_)  &  poutreg_60_ ) | ( pdata_48_  &  pcount_0_  &  wire577 ) ;
 assign pdata_new_50_ = ( wire1021 ) | ( pinreg_36_  &  n_n1327 ) ;
 assign pdata_new_63_ = ( pdata_in_6_  &  n_n1327 ) | ( (~ n_n1327)  &  wire343 ) ;
 assign poutreg_new_30_ = ( wire8362 ) | ( (~ pcount_0_)  &  poutreg_30_ ) ;
 assign poutreg_new_43_ = ( wire995 ) | ( wire8375 ) ;
 assign poutreg_new_56_ = ( (~ pcount_0_)  &  poutreg_56_ ) | ( pcount_0_  &  pdata_32_  &  wire577 ) ;
 assign poutreg_new_44_ = ( wire8376 ) | ( (~ pcount_0_)  &  poutreg_44_ ) ;
 assign poutreg_new_55_ = ( wire8377 ) | ( n_n1327  &  wire351 ) ;
 assign pdata_new_61_ = ( pinreg_14_  &  n_n1327 ) | ( (~ n_n1327)  &  wire366 ) ;
 assign pencrypt_mode_new_0_ = ( pencrypt_0_  &  n_n1327 ) | ( pencrypt_mode_0_  &  (~ n_n1327) ) ;
 assign poutreg_new_41_ = ( wire8397 ) | ( n_n1327  &  wire367 ) ;
 assign poutreg_new_58_ = ( (~ pcount_0_)  &  poutreg_58_ ) | ( pcount_0_  &  pdata_40_  &  wire577 ) ;
 assign pdata_new_40_ = ( pinreg_50_  &  n_n1327 ) | ( (~ n_n1327)  &  wire368 ) ;
 assign pdata_new_62_ = ( pinreg_6_  &  n_n1327 ) | ( (~ pdata_30_)  &  (~ n_n1327)  &  n_n1736 ) | ( pdata_30_  &  (~ n_n1327)  &  (~ n_n1736) ) ;
 assign poutreg_new_20_ = ( wire8406 ) | ( (~ pcount_0_)  &  poutreg_20_ ) ;
 assign poutreg_new_42_ = ( wire8407 ) | ( (~ pcount_0_)  &  poutreg_42_ ) ;
 assign poutreg_new_57_ = ( (~ pcount_0_)  &  poutreg_57_ ) | ( n_n1327  &  wire369 ) ;
 assign pdata_new_41_ = ( pinreg_42_  &  n_n1327 ) | ( (~ n_n1327)  &  wire362 ) ;
 assign pdata_new_54_ = ( pinreg_4_  &  n_n1327 ) | ( (~ n_n1327)  &  wire370 ) ;
 assign pinreg_new_40_ = ( (~ pcount_0_)  &  pinreg_40_ ) | ( pcount_0_  &  pinreg_32_  &  (~ wire577) ) ;
 assign pinreg_new_51_ = ( (~ pcount_0_)  &  pinreg_51_ ) | ( pcount_0_  &  pinreg_43_  &  (~ wire577) ) ;
 assign poutreg_new_21_ = ( wire8443 ) | ( n_n1327  &  wire371 ) ;
 assign poutreg_new_34_ = ( wire8444 ) | ( (~ pcount_0_)  &  poutreg_34_ ) ;
 assign pd_new_20_ = ( wire848 ) | ( wire849 ) | ( wire8449 ) ;
 assign pdata_new_0_ = ( pinreg_49_  &  n_n1327 ) | ( pdata_32_  &  (~ n_n1327) ) ;
 assign pdata_new_42_ = ( wire842 ) | ( pinreg_34_  &  n_n1327 ) ;
 assign pdata_new_53_ = ( pinreg_12_  &  n_n1327 ) | ( (~ n_n1327)  &  wire371 ) ;
 assign pdata_new_60_ = ( wire820 ) | ( pinreg_22_  &  n_n1327 ) ;
 assign pinreg_new_41_ = ( (~ pcount_0_)  &  pinreg_41_ ) | ( pcount_0_  &  pinreg_33_  &  (~ wire577) ) ;
 assign pinreg_new_50_ = ( (~ pcount_0_)  &  pinreg_50_ ) | ( pcount_0_  &  pinreg_42_  &  (~ wire577) ) ;
 assign poutreg_new_22_ = ( wire8460 ) | ( (~ pcount_0_)  &  poutreg_22_ ) ;
 assign poutreg_new_33_ = ( wire810 ) | ( wire8461 ) ;
 assign poutreg_new_40_ = ( wire8462 ) | ( poutreg_40_  &  (~ pcount_0_) ) ;
 assign poutreg_new_59_ = ( (~ pcount_0_)  &  poutreg_59_ ) | ( n_n1327  &  wire368 ) ;
 assign pc_new_20_ = ( wire800 ) | ( wire801 ) | ( wire8467 ) ;
 assign pd_new_10_ = ( wire793 ) | ( wire794 ) | ( wire8472 ) ;
 assign pdata_new_43_ = ( pinreg_26_  &  n_n1327 ) | ( (~ n_n1327)  &  wire359 ) ;
 assign pdata_new_52_ = ( wire787 ) | ( pinreg_20_  &  n_n1327 ) ;
 assign pinreg_new_20_ = ( (~ pcount_0_)  &  pinreg_20_ ) | ( pcount_0_  &  pinreg_12_  &  (~ wire577) ) ;
 assign pinreg_new_31_ = ( (~ pcount_0_)  &  pinreg_31_ ) | ( pcount_0_  &  pinreg_23_  &  (~ wire577) ) ;
 assign poutreg_new_23_ = ( wire8473 ) | ( n_n1327  &  wire366 ) ;
 assign poutreg_new_32_ = ( wire8474 ) | ( (~ pcount_0_)  &  poutreg_32_ ) ;
 assign pc_new_10_ = ( wire772 ) | ( wire773 ) | ( wire8479 ) ;
 assign pdata_new_44_ = ( pinreg_18_  &  n_n1327 ) | ( (~ pdata_12_)  &  (~ n_n1327)  &  n_n1742 ) | ( pdata_12_  &  (~ n_n1327)  &  (~ n_n1742) ) ;
 assign pdata_new_51_ = ( pinreg_28_  &  n_n1327 ) | ( (~ n_n1327)  &  wire352 ) ;
 assign pinreg_new_21_ = ( (~ pcount_0_)  &  pinreg_21_ ) | ( pcount_0_  &  pinreg_13_  &  (~ wire577) ) ;
 assign pinreg_new_30_ = ( (~ pcount_0_)  &  pinreg_30_ ) | ( pcount_0_  &  pinreg_22_  &  (~ wire577) ) ;
 assign poutreg_new_24_ = ( wire8480 ) | ( (~ pcount_0_)  &  poutreg_24_ ) ;
 assign poutreg_new_31_ = ( wire756 ) | ( wire8481 ) ;
 assign pdata_new_32_ = ( pinreg_48_  &  n_n1327 ) | ( (~ n_n1327)  &  wire369 ) ;
 assign pinreg_new_11_ = ( (~ pcount_0_)  &  pinreg_11_ ) | ( pcount_0_  &  pinreg_3_  &  (~ wire577) ) ;
 assign poutreg_new_12_ = ( wire8482 ) | ( (~ pcount_0_)  &  poutreg_12_ ) ;
 assign pdata_new_20_ = ( pinreg_21_  &  n_n1327 ) | ( pdata_52_  &  (~ n_n1327) ) ;
 assign pdata_new_31_ = ( pdata_in_7_  &  n_n1327 ) | ( pdata_63_  &  (~ n_n1327) ) ;
 assign pinreg_new_10_ = ( (~ pcount_0_)  &  pinreg_10_ ) | ( pcount_0_  &  pinreg_2_  &  (~ wire577) ) ;
 assign poutreg_new_11_ = ( wire492 ) | ( wire8483 ) ;
 assign pdata_new_34_ = ( pinreg_32_  &  n_n1327 ) | ( (~ n_n1327)  &  wire367 ) ;
 assign poutreg_new_14_ = ( wire8484 ) | ( (~ pcount_0_)  &  poutreg_14_ ) ;
 assign pdata_new_19_ = ( pinreg_29_  &  n_n1327 ) | ( pdata_51_  &  (~ n_n1327) ) ;
 assign pdata_new_33_ = ( pinreg_40_  &  n_n1327 ) | ( (~ pdata_1_)  &  (~ n_n1327)  &  n_n1753 ) | ( pdata_1_  &  (~ n_n1327)  &  (~ n_n1753) ) ;
 assign poutreg_new_13_ = ( wire8485 ) | ( n_n1327  &  wire370 ) ;
 assign pd_new_9_ = ( wire453 ) | ( wire454 ) | ( wire8490 ) ;
 assign pdata_new_18_ = ( pinreg_37_  &  n_n1327 ) | ( pdata_50_  &  (~ n_n1327) ) ;
 assign pdata_new_23_ = ( pdata_in_5_  &  n_n1327 ) | ( pdata_55_  &  (~ n_n1327) ) ;
 assign pdata_new_17_ = ( pinreg_45_  &  n_n1327 ) | ( pdata_49_  &  (~ n_n1327) ) ;
 assign pdata_new_24_ = ( pinreg_55_  &  n_n1327 ) | ( pdata_56_  &  (~ n_n1327) ) ;
 assign pinreg_new_9_ = ( (~ pcount_0_)  &  pinreg_9_ ) | ( pinreg_1_  &  pcount_0_  &  (~ wire577) ) ;
 assign pc_new_8_ = ( wire429 ) | ( wire430 ) | ( wire8495 ) ;
 assign pd_new_7_ = ( wire415 ) | ( wire416 ) | ( wire8500 ) ;
 assign pdata_new_16_ = ( pinreg_53_  &  n_n1327 ) | ( pdata_48_  &  (~ n_n1327) ) ;
 assign pdata_new_21_ = ( pinreg_13_  &  n_n1327 ) | ( pdata_53_  &  (~ n_n1327) ) ;
 assign pdata_new_30_ = ( pinreg_7_  &  n_n1327 ) | ( pdata_62_  &  (~ n_n1327) ) ;
 assign poutreg_new_10_ = ( wire8501 ) | ( (~ pcount_0_)  &  poutreg_10_ ) ;
 assign pc_new_9_ = ( wire378 ) | ( wire382 ) | ( wire8506 ) ;
 assign pd_new_8_ = ( wire330 ) | ( wire332 ) | ( wire8511 ) ;
 assign pdata_new_15_ = ( pdata_in_3_  &  n_n1327 ) | ( pdata_47_  &  (~ n_n1327) ) ;
 assign pdata_new_22_ = ( pinreg_5_  &  n_n1327 ) | ( pdata_54_  &  (~ n_n1327) ) ;
 assign wire254 = ( (~ preset_0_)  &  (~ pload_key_0_)  &  n_n1327  &  wire616 ) ;
 assign n_n1327 = ( pcount_3_  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) ;
 assign wire340 = ( (~ pdata_6_)  &  wire7751 ) | ( (~ pdata_6_)  &  wire7752 ) | ( (~ pdata_6_)  &  wire7753 ) | ( pdata_6_  &  (~ wire7751)  &  (~ wire7752)  &  (~ wire7753) ) ;
 assign wire341 = ( (~ pdata_7_)  &  wire7785 ) | ( (~ pdata_7_)  &  wire7786 ) | ( (~ pdata_7_)  &  wire7787 ) | ( pdata_7_  &  (~ wire7785)  &  (~ wire7786)  &  (~ wire7787) ) ;
 assign wire342 = ( (~ pdata_13_)  &  wire277 ) | ( (~ pdata_13_)  &  wire2162 ) | ( (~ pdata_13_)  &  wire7799 ) | ( pdata_13_  &  (~ wire277)  &  (~ wire2162)  &  (~ wire7799) ) ;
 assign wire343 = ( (~ pdata_31_)  &  wire278 ) | ( (~ pdata_31_)  &  wire7816 ) | ( (~ pdata_31_)  &  wire7819 ) | ( pdata_31_  &  (~ wire278)  &  (~ wire7816)  &  (~ wire7819) ) ;
 assign wire514 = ( (~ preset_0_)  &  (~ pload_key_0_) ) | ( (~ preset_0_)  &  (~ n_n1327) ) ;
 assign wire348 = ( (~ pdata_26_)  &  wire8004 ) | ( (~ pdata_26_)  &  wire8005 ) | ( (~ pdata_26_)  &  wire8006 ) | ( pdata_26_  &  (~ wire8004)  &  (~ wire8005)  &  (~ wire8006) ) ;
 assign wire351 = ( (~ pdata_25_)  &  wire279 ) | ( (~ pdata_25_)  &  wire8077 ) | ( (~ pdata_25_)  &  wire8078 ) | ( pdata_25_  &  (~ wire279)  &  (~ wire8077)  &  (~ wire8078) ) ;
 assign wire352 = ( (~ pdata_19_)  &  wire279 ) | ( (~ pdata_19_)  &  wire8092 ) | ( (~ pdata_19_)  &  wire8096 ) | ( pdata_19_  &  (~ wire279)  &  (~ wire8092)  &  (~ wire8096) ) ;
 assign wire355 = ( (~ pdata_24_)  &  wire8138 ) | ( (~ pdata_24_)  &  wire8139 ) | ( (~ pdata_24_)  &  wire8140 ) | ( pdata_24_  &  (~ wire8138)  &  (~ wire8139)  &  (~ wire8140) ) ;
 assign wire359 = ( (~ pdata_11_)  &  wire278 ) | ( (~ pdata_11_)  &  wire8218 ) | ( (~ pdata_11_)  &  wire8219 ) | ( pdata_11_  &  (~ wire278)  &  (~ wire8218)  &  (~ wire8219) ) ;
 assign wire392 = ( (~ pcount_3_)  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) ;
 assign wire362 = ( (~ pdata_9_)  &  wire279 ) | ( (~ pdata_9_)  &  wire8293 ) | ( (~ pdata_9_)  &  wire8294 ) | ( pdata_9_  &  (~ wire279)  &  (~ wire8293)  &  (~ wire8294) ) ;
 assign wire364 = ( (~ pdata_27_)  &  wire322 ) | ( (~ pdata_27_)  &  wire1049 ) | ( (~ pdata_27_)  &  wire8356 ) | ( pdata_27_  &  (~ wire322)  &  (~ wire1049)  &  (~ wire8356) ) ;
 assign wire366 = ( (~ pdata_29_)  &  wire323 ) | ( (~ pdata_29_)  &  wire975 ) | ( (~ pdata_29_)  &  wire8385 ) | ( pdata_29_  &  (~ wire323)  &  (~ wire975)  &  (~ wire8385) ) ;
 assign wire367 = ( (~ pdata_2_)  &  wire277 ) | ( (~ pdata_2_)  &  wire8393 ) | ( (~ pdata_2_)  &  wire8396 ) | ( pdata_2_  &  (~ wire277)  &  (~ wire8393)  &  (~ wire8396) ) ;
 assign wire368 = ( (~ pdata_8_)  &  wire275 ) | ( (~ pdata_8_)  &  wire8403 ) | ( (~ pdata_8_)  &  wire8404 ) | ( pdata_8_  &  (~ wire275)  &  (~ wire8403)  &  (~ wire8404) ) ;
 assign wire369 = ( (~ pdata_0_)  &  wire8416 ) | ( (~ pdata_0_)  &  wire8417 ) | ( (~ pdata_0_)  &  wire8418 ) | ( pdata_0_  &  (~ wire8416)  &  (~ wire8417)  &  (~ wire8418) ) ;
 assign wire370 = ( (~ pdata_22_)  &  wire275 ) | ( (~ pdata_22_)  &  wire8428 ) | ( (~ pdata_22_)  &  wire8429 ) | ( pdata_22_  &  (~ wire275)  &  (~ wire8428)  &  (~ wire8429) ) ;
 assign wire371 = ( (~ pdata_21_)  &  wire278 ) | ( (~ pdata_21_)  &  wire8440 ) | ( (~ pdata_21_)  &  wire8441 ) | ( pdata_21_  &  (~ wire278)  &  (~ wire8440)  &  (~ wire8441) ) ;
 assign wire577 = ( pcount_3_  &  pcount_2_  &  pcount_1_ ) ;
 assign n_n1709 = ( (~ pdata_42_)  &  pc_3_ ) | ( pdata_42_  &  (~ pc_3_) ) ;
 assign n_n1710 = ( (~ pdata_41_)  &  pc_11_ ) | ( pdata_41_  &  (~ pc_11_) ) ;
 assign n_n1712 = ( (~ pc_22_)  &  pdata_39_ ) | ( pc_22_  &  (~ pdata_39_) ) ;
 assign n_n1708 = ( (~ pdata_43_)  &  pc_25_ ) | ( pdata_43_  &  (~ pc_25_) ) ;
 assign n_n1707 = ( (~ pdata_44_)  &  pc_7_ ) | ( pdata_44_  &  (~ pc_7_) ) ;
 assign n_n1696 = ( (~ pd_18_)  &  pdata_51_ ) | ( pd_18_  &  (~ pdata_51_) ) ;
 assign n_n1699 = ( (~ pdata_48_)  &  pd_23_ ) | ( pdata_48_  &  (~ pd_23_) ) ;
 assign n_n1700 = ( (~ pdata_47_)  &  pd_12_ ) | ( pdata_47_  &  (~ pd_12_) ) ;
 assign n_n1695 = ( (~ pd_26_)  &  pdata_52_ ) | ( pd_26_  &  (~ pdata_52_) ) ;
 assign n_n1715 = ( (~ pd_16_)  &  pdata_54_ ) | ( pd_16_  &  (~ pdata_54_) ) ;
 assign n_n1714 = ( (~ pd_4_)  &  pdata_55_ ) | ( pd_4_  &  (~ pdata_55_) ) ;
 assign n_n1716 = ( (~ pd_22_)  &  pdata_53_ ) | ( pd_22_  &  (~ pdata_53_) ) ;
 assign n_n1713 = ( (~ pd_19_)  &  pdata_56_ ) | ( pd_19_  &  (~ pdata_56_) ) ;
 assign n_n1718 = ( (~ pd_1_)  &  pdata_51_ ) | ( pd_1_  &  (~ pdata_51_) ) ;
 assign n_n1723 = ( (~ pd_20_)  &  pdata_56_ ) | ( pd_20_  &  (~ pdata_56_) ) ;
 assign n_n1724 = ( (~ pd_15_)  &  pdata_55_ ) | ( pd_15_  &  (~ pdata_55_) ) ;
 assign n_n1720 = ( (~ pdata_59_)  &  pd_5_ ) | ( pdata_59_  &  (~ pd_5_) ) ;
 assign n_n1719 = ( (~ pdata_60_)  &  pd_24_ ) | ( pdata_60_  &  (~ pd_24_) ) ;
 assign n_n1726 = ( (~ pd_0_)  &  pdata_63_ ) | ( pd_0_  &  (~ pdata_63_) ) ;
 assign n_n1728 = ( (~ pd_21_)  &  pdata_61_ ) | ( pd_21_  &  (~ pdata_61_) ) ;
 assign n_n1725 = ( (~ pdata_32_)  &  pd_3_ ) | ( pdata_32_  &  (~ pd_3_) ) ;
 assign n_n1730 = ( (~ pdata_59_)  &  pd_17_ ) | ( pdata_59_  &  (~ pd_17_) ) ;
 assign n_n1697 = ( (~ pd_8_)  &  pdata_50_ ) | ( pd_8_  &  (~ pdata_50_) ) ;
 assign n_n1702 = ( (~ pdata_35_)  &  pc_0_ ) | ( pdata_35_  &  (~ pc_0_) ) ;
 assign n_n1704 = ( (~ pdata_33_)  &  pc_10_ ) | ( pdata_33_  &  (~ pc_10_) ) ;
 assign n_n1706 = ( (~ pc_13_)  &  pdata_63_ ) | ( pc_13_  &  (~ pdata_63_) ) ;
 assign n_n1329 = ( pcount_3_  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) | ( (~ pcount_3_)  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) | ( pcount_3_  &  pcount_2_  &  pcount_1_  &  (~ pcount_0_) ) | ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_) ) ;
 assign wire616 = ( (~ pencrypt_0_)  &  pencrypt_mode_0_ ) | ( pencrypt_0_  &  (~ pencrypt_mode_0_) ) ;
 assign n_n1684 = ( (~ pdata_37_)  &  pc_14_ ) | ( pdata_37_  &  (~ pc_14_) ) ;
 assign n_n1686 = ( (~ pdata_35_)  &  pc_2_ ) | ( pdata_35_  &  (~ pc_2_) ) ;
 assign n_n1727 = ( (~ pd_7_)  &  pdata_62_ ) | ( pd_7_  &  (~ pdata_62_) ) ;
 assign n_n1705 = ( (~ pdata_32_)  &  pc_16_ ) | ( pdata_32_  &  (~ pc_16_) ) ;
 assign n_n1701 = ( (~ pdata_36_)  &  pc_4_ ) | ( pdata_36_  &  (~ pc_4_) ) ;
 assign wire264 = ( (~ pdata_35_)  &  pdata_36_  &  pc_4_  &  pc_0_ ) | ( pdata_35_  &  (~ pdata_36_)  &  pc_4_  &  pc_0_ ) | ( pdata_35_  &  pdata_36_  &  (~ pc_4_)  &  pc_0_ ) | ( (~ pdata_35_)  &  (~ pdata_36_)  &  (~ pc_4_)  &  pc_0_ ) | ( pdata_35_  &  pdata_36_  &  pc_4_  &  (~ pc_0_) ) | ( (~ pdata_35_)  &  (~ pdata_36_)  &  pc_4_  &  (~ pc_0_) ) | ( (~ pdata_35_)  &  pdata_36_  &  (~ pc_4_)  &  (~ pc_0_) ) | ( pdata_35_  &  (~ pdata_36_)  &  (~ pc_4_)  &  (~ pc_0_) ) ;
 assign wire275 = ( wire1922 ) | ( wire1923 ) | ( wire8013 ) ;
 assign wire325 = ( pc_13_  &  pdata_63_  &  n_n1705 ) | ( (~ pc_13_)  &  (~ pdata_63_)  &  n_n1705 ) | ( (~ pc_13_)  &  pdata_63_  &  (~ n_n1705)  &  n_n1703 ) | ( pc_13_  &  (~ pdata_63_)  &  (~ n_n1705)  &  n_n1703 ) ;
 assign wire465 = ( wire1913 ) | ( wire1914 ) | ( (~ wire496)  &  wire734 ) ;
 assign wire512 = ( pdata_35_  &  (~ pdata_36_)  &  pc_4_  &  pc_0_ ) | ( pdata_35_  &  pdata_36_  &  (~ pc_4_)  &  pc_0_ ) | ( (~ pdata_35_)  &  (~ pdata_36_)  &  pc_4_  &  (~ pc_0_) ) | ( (~ pdata_35_)  &  pdata_36_  &  (~ pc_4_)  &  (~ pc_0_) ) ;
 assign wire568 = ( pdata_33_  &  (~ pdata_34_)  &  pc_10_  &  pc_23_ ) | ( (~ pdata_33_)  &  (~ pdata_34_)  &  (~ pc_10_)  &  pc_23_ ) | ( pdata_33_  &  pdata_34_  &  pc_10_  &  (~ pc_23_) ) | ( (~ pdata_33_)  &  pdata_34_  &  (~ pc_10_)  &  (~ pc_23_) ) ;
 assign wire594 = ( (~ pdata_33_)  &  pdata_34_  &  pc_10_  &  pc_23_ ) | ( pdata_33_  &  pdata_34_  &  (~ pc_10_)  &  pc_23_ ) | ( (~ pdata_33_)  &  (~ pdata_34_)  &  pc_10_  &  (~ pc_23_) ) | ( pdata_33_  &  (~ pdata_34_)  &  (~ pc_10_)  &  (~ pc_23_) ) ;
 assign n_n1711 = ( (~ pdata_40_)  &  pc_18_ ) | ( pdata_40_  &  (~ pc_18_) ) ;
 assign n_n1703 = ( (~ pdata_34_)  &  pc_23_ ) | ( pdata_34_  &  (~ pc_23_) ) ;
 assign n_n1690 = ( (~ pdata_47_)  &  pc_12_ ) | ( pdata_47_  &  (~ pc_12_) ) ;
 assign n_n1722 = ( (~ pd_10_)  &  pdata_57_ ) | ( pd_10_  &  (~ pdata_57_) ) ;
 assign n_n1687 = ( (~ pdata_40_)  &  pc_9_ ) | ( pdata_40_  &  (~ pc_9_) ) ;
 assign n_n1688 = ( (~ pc_20_)  &  pdata_39_ ) | ( pc_20_  &  (~ pdata_39_) ) ;
 assign n_n1683 = ( (~ pdata_38_)  &  pc_5_ ) | ( pdata_38_  &  (~ pc_5_) ) ;
 assign n_n1685 = ( (~ pdata_36_)  &  pc_27_ ) | ( pdata_36_  &  (~ pc_27_) ) ;
 assign n_n1698 = ( (~ pd_2_)  &  pdata_49_ ) | ( pd_2_  &  (~ pdata_49_) ) ;
 assign n_n1721 = ( (~ pd_27_)  &  pdata_58_ ) | ( pd_27_  &  (~ pdata_58_) ) ;
 assign n_n1729 = ( (~ pdata_60_)  &  pd_13_ ) | ( pdata_60_  &  (~ pd_13_) ) ;
 assign n_n1717 = ( (~ pd_11_)  &  pdata_52_ ) | ( pd_11_  &  (~ pdata_52_) ) ;
 assign wire462 = ( wire1397 ) | ( wire1399 ) | ( wire533  &  wire732 ) ;
 assign wire620 = ( wire1383 ) | ( wire1384 ) | ( wire1385 ) | ( wire1386 ) ;
 assign n_n1753 = ( wire1380 ) | ( wire8153 ) | ( wire8154 ) | ( wire8176 ) ;
 assign n_n1694 = ( (~ pdata_43_)  &  pc_15_ ) | ( pdata_43_  &  (~ pc_15_) ) ;
 assign wire333 = ( wire1929 ) | ( wire1930 ) | ( wire532  &  wire717 ) ;
 assign wire393 = ( wire1923 ) | ( wire594  &  wire532  &  wire520 ) ;
 assign wire423 = ( pdata_34_  &  pc_23_  &  wire319 ) | ( (~ pdata_34_)  &  (~ pc_23_)  &  wire319 ) ;
 assign wire592 = ( pdata_35_  &  pdata_36_  &  pc_4_  &  pc_0_ ) | ( pdata_35_  &  (~ pdata_36_)  &  (~ pc_4_)  &  pc_0_ ) | ( (~ pdata_35_)  &  pdata_36_  &  pc_4_  &  (~ pc_0_) ) | ( (~ pdata_35_)  &  (~ pdata_36_)  &  (~ pc_4_)  &  (~ pc_0_) ) ;
 assign wire626 = ( wire423 ) | ( wire1904 ) | ( wire1905 ) | ( wire1906 ) ;
 assign n_n1736 = ( wire393 ) | ( wire1895 ) | ( wire7919 ) | ( wire7920 ) ;
 assign wire280 = ( pd_0_  &  pdata_63_  &  (~ n_n1730)  &  wire511 ) | ( (~ pd_0_)  &  (~ pdata_63_)  &  (~ n_n1730)  &  wire511 ) ;
 assign wire297 = ( pdata_32_  &  (~ pd_7_)  &  pd_3_  &  pdata_62_ ) | ( (~ pdata_32_)  &  (~ pd_7_)  &  (~ pd_3_)  &  pdata_62_ ) | ( pdata_32_  &  pd_7_  &  pd_3_  &  (~ pdata_62_) ) | ( (~ pdata_32_)  &  pd_7_  &  (~ pd_3_)  &  (~ pdata_62_) ) ;
 assign wire396 = ( (~ pdata_60_)  &  pd_13_  &  wire265  &  wire7853 ) | ( pdata_60_  &  (~ pd_13_)  &  wire265  &  wire7853 ) ;
 assign wire424 = ( (~ pd_0_)  &  pdata_63_  &  wire562  &  wire7863 ) | ( pd_0_  &  (~ pdata_63_)  &  wire562  &  wire7863 ) ;
 assign wire470 = ( wire2038 ) | ( wire2039 ) | ( wire2040 ) | ( wire2041 ) ;
 assign wire475 = ( wire2035 ) | ( wire2036 ) | ( wire2037 ) ;
 assign wire531 = ( pdata_32_  &  pd_7_  &  pd_3_  &  pdata_62_ ) | ( (~ pdata_32_)  &  pd_7_  &  (~ pd_3_)  &  pdata_62_ ) | ( pdata_32_  &  (~ pd_7_)  &  pd_3_  &  (~ pdata_62_) ) | ( (~ pdata_32_)  &  (~ pd_7_)  &  (~ pd_3_)  &  (~ pdata_62_) ) ;
 assign n_n1691 = ( (~ pdata_46_)  &  pc_19_ ) | ( pdata_46_  &  (~ pc_19_) ) ;
 assign n_n1693 = ( (~ pdata_44_)  &  pc_6_ ) | ( pdata_44_  &  (~ pc_6_) ) ;
 assign n_n1692 = ( (~ pdata_45_)  &  pc_26_ ) | ( pdata_45_  &  (~ pc_26_) ) ;
 assign wire247 = ( pdata_44_  &  pdata_42_  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  (~ pc_7_)  &  pc_3_ ) | ( pdata_44_  &  (~ pdata_42_)  &  (~ pc_7_)  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  (~ pdata_42_)  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  pdata_42_  &  (~ pc_7_)  &  (~ pc_3_) ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign wire270 = ( (~ pdata_43_)  &  pdata_41_  &  pc_11_  &  pc_25_ ) | ( pdata_43_  &  (~ pdata_41_)  &  pc_11_  &  pc_25_ ) | ( pdata_43_  &  pdata_41_  &  (~ pc_11_)  &  pc_25_ ) | ( (~ pdata_43_)  &  (~ pdata_41_)  &  (~ pc_11_)  &  pc_25_ ) | ( pdata_43_  &  pdata_41_  &  pc_11_  &  (~ pc_25_) ) | ( (~ pdata_43_)  &  (~ pdata_41_)  &  pc_11_  &  (~ pc_25_) ) | ( (~ pdata_43_)  &  pdata_41_  &  (~ pc_11_)  &  (~ pc_25_) ) | ( pdata_43_  &  (~ pdata_41_)  &  (~ pc_11_)  &  (~ pc_25_) ) ;
 assign wire323 = ( wire473 ) | ( wire474 ) | ( wire480 ) ;
 assign wire328 = ( pdata_43_  &  pc_22_  &  pc_25_  &  pdata_39_ ) | ( (~ pdata_43_)  &  (~ pc_22_)  &  pc_25_  &  pdata_39_ ) | ( (~ pdata_43_)  &  pc_22_  &  (~ pc_25_)  &  pdata_39_ ) | ( pdata_43_  &  (~ pc_22_)  &  (~ pc_25_)  &  pdata_39_ ) | ( (~ pdata_43_)  &  pc_22_  &  pc_25_  &  (~ pdata_39_) ) | ( pdata_43_  &  (~ pc_22_)  &  pc_25_  &  (~ pdata_39_) ) | ( pdata_43_  &  pc_22_  &  (~ pc_25_)  &  (~ pdata_39_) ) | ( (~ pdata_43_)  &  (~ pc_22_)  &  (~ pc_25_)  &  (~ pdata_39_) ) ;
 assign wire398 = ( wire1839 ) | ( (~ n_n1710)  &  wire1841 ) | ( (~ n_n1710)  &  wire1842 ) ;
 assign wire507 = ( (~ pdata_44_)  &  (~ pdata_42_)  &  pc_7_  &  pc_3_ ) | ( pdata_44_  &  (~ pdata_42_)  &  (~ pc_7_)  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  pdata_42_  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign wire525 = ( (~ pdata_44_)  &  pdata_42_  &  pc_7_  &  pc_3_ ) | ( pdata_44_  &  pdata_42_  &  (~ pc_7_)  &  pc_3_ ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  (~ pdata_42_)  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign wire537 = ( (~ pdata_40_)  &  pc_22_  &  pc_18_  &  pdata_39_ ) | ( pdata_40_  &  pc_22_  &  (~ pc_18_)  &  pdata_39_ ) | ( (~ pdata_40_)  &  (~ pc_22_)  &  pc_18_  &  (~ pdata_39_) ) | ( pdata_40_  &  (~ pc_22_)  &  (~ pc_18_)  &  (~ pdata_39_) ) ;
 assign wire630 = ( (~ pdata_41_)  &  pc_11_  &  n_n1708  &  n_n1711 ) | ( pdata_41_  &  (~ pc_11_)  &  n_n1708  &  n_n1711 ) | ( (~ pdata_41_)  &  pc_11_  &  (~ n_n1708)  &  (~ n_n1711) ) | ( pdata_41_  &  (~ pc_11_)  &  (~ n_n1708)  &  (~ n_n1711) ) ;
 assign n_n1689 = ( (~ pdata_48_)  &  pc_1_ ) | ( pdata_48_  &  (~ pc_1_) ) ;
 assign wire277 = ( wire2228 ) | ( wire7775 ) | ( wire539  &  wire726 ) ;
 assign wire467 = ( wire2218 ) | ( wire2219 ) | ( wire304  &  wire735 ) ;
 assign wire471 = ( wire2212 ) | ( wire2214 ) | ( wire527  &  wire738 ) ;
 assign wire634 = ( wire2208 ) | ( wire2209 ) | ( wire2210 ) | ( wire2211 ) ;
 assign wire632 = ( wire2202 ) | ( (~ n_n1700)  &  wire304  &  wire303 ) ;
 assign wire631 = ( pd_8_  &  pd_18_  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  (~ pd_18_)  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  (~ pdata_50_)  &  pdata_51_ ) | ( pd_8_  &  (~ pd_18_)  &  (~ pdata_50_)  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  (~ pd_18_)  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  pd_18_  &  (~ pdata_50_)  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  (~ pd_18_)  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire307 = ( pdata_38_  &  pc_20_  &  pc_5_  &  pdata_39_ ) | ( (~ pdata_38_)  &  pc_20_  &  (~ pc_5_)  &  pdata_39_ ) | ( pdata_38_  &  (~ pc_20_)  &  pc_5_  &  (~ pdata_39_) ) | ( (~ pdata_38_)  &  (~ pc_20_)  &  (~ pc_5_)  &  (~ pdata_39_) ) ;
 assign wire463 = ( wire1425 ) | ( wire1426 ) | ( wire1427 ) | ( wire1428 ) ;
 assign wire636 = ( (~ n_n1686)  &  (~ n_n1687)  &  (~ n_n1688)  &  n_n1683 ) | ( n_n1686  &  n_n1687  &  n_n1688  &  (~ n_n1683) ) ;
 assign n_n1742 = ( wire1411 ) | ( wire8153 ) | ( wire8154 ) | ( wire8166 ) ;
 assign wire278 = ( wire401 ) | ( wire2127 ) | ( wire510  &  wire714 ) ;
 assign wire306 = ( (~ pd_20_)  &  pd_27_  &  pdata_58_  &  pdata_56_ ) | ( (~ pd_20_)  &  (~ pd_27_)  &  (~ pdata_58_)  &  pdata_56_ ) | ( pd_20_  &  pd_27_  &  pdata_58_  &  (~ pdata_56_) ) | ( pd_20_  &  (~ pd_27_)  &  (~ pdata_58_)  &  (~ pdata_56_) ) ;
 assign wire315 = ( (~ pd_10_)  &  pdata_60_  &  pd_24_  &  pdata_57_ ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  (~ pd_24_)  &  pdata_57_ ) | ( pd_10_  &  pdata_60_  &  pd_24_  &  (~ pdata_57_) ) | ( pd_10_  &  (~ pdata_60_)  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire472 = ( wire510  &  wire740 ) | ( wire541  &  wire739 ) ;
 assign wire518 = ( pd_10_  &  (~ pd_15_)  &  pdata_57_  &  pdata_55_ ) | ( (~ pd_10_)  &  (~ pd_15_)  &  (~ pdata_57_)  &  pdata_55_ ) | ( pd_10_  &  pd_15_  &  pdata_57_  &  (~ pdata_55_) ) | ( (~ pd_10_)  &  pd_15_  &  (~ pdata_57_)  &  (~ pdata_55_) ) ;
 assign wire335 = ( wire2309 ) | ( wire2311 ) | ( wire294  &  wire718 ) ;
 assign wire401 = ( wire2304 ) | ( wire2306 ) | ( wire559  &  wire725 ) ;
 assign wire402 = ( pd_27_  &  pdata_58_  &  wire315  &  wire7738 ) | ( (~ pd_27_)  &  (~ pdata_58_)  &  wire315  &  wire7738 ) ;
 assign wire417 = ( (~ pdata_59_)  &  pd_5_ ) | ( pdata_59_  &  (~ pd_5_) ) | ( (~ pd_15_)  &  pdata_55_ ) | ( pd_15_  &  (~ pdata_55_) ) ;
 assign wire529 = ( (~ pd_10_)  &  (~ pdata_60_)  &  pd_24_  &  pdata_57_ ) | ( (~ pd_10_)  &  pdata_60_  &  (~ pd_24_)  &  pdata_57_ ) | ( pd_10_  &  (~ pdata_60_)  &  pd_24_  &  (~ pdata_57_) ) | ( pd_10_  &  pdata_60_  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire541 = ( pd_10_  &  (~ pdata_60_)  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  pdata_60_  &  (~ pd_24_)  &  pdata_57_ ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  pdata_60_  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire584 = ( (~ pdata_59_)  &  (~ pd_20_)  &  pd_5_  &  pdata_56_ ) | ( pdata_59_  &  (~ pd_20_)  &  (~ pd_5_)  &  pdata_56_ ) | ( (~ pdata_59_)  &  pd_20_  &  pd_5_  &  (~ pdata_56_) ) | ( pdata_59_  &  pd_20_  &  (~ pd_5_)  &  (~ pdata_56_) ) ;
 assign wire646 = ( pd_15_  &  pdata_55_  &  (~ n_n1720)  &  n_n1721 ) | ( (~ pd_15_)  &  (~ pdata_55_)  &  (~ n_n1720)  &  n_n1721 ) | ( pd_15_  &  pdata_55_  &  n_n1720  &  (~ n_n1721) ) | ( (~ pd_15_)  &  (~ pdata_55_)  &  n_n1720  &  (~ n_n1721) ) | ( (~ pd_15_)  &  pdata_55_  &  (~ n_n1720)  &  (~ n_n1721) ) | ( pd_15_  &  (~ pdata_55_)  &  (~ n_n1720)  &  (~ n_n1721) ) ;
 assign wire645 = ( n_n1723  &  n_n1721  &  wire7731 ) | ( n_n1723  &  (~ n_n1721)  &  wire7744 ) ;
 assign wire289 = ( (~ pdata_48_)  &  pd_23_  &  (~ pd_26_)  &  pdata_52_ ) | ( pdata_48_  &  (~ pd_23_)  &  (~ pd_26_)  &  pdata_52_ ) | ( (~ pdata_48_)  &  pd_23_  &  pd_26_  &  (~ pdata_52_) ) | ( pdata_48_  &  (~ pd_23_)  &  pd_26_  &  (~ pdata_52_) ) ;
 assign wire336 = ( wire2182 ) | ( wire2184 ) | ( (~ wire420)  &  wire719 ) ;
 assign wire485 = ( wire289  &  wire283 ) ;
 assign wire552 = ( (~ pd_8_)  &  pd_18_  &  pdata_50_  &  pdata_51_ ) | ( pd_8_  &  pd_18_  &  (~ pdata_50_)  &  pdata_51_ ) | ( (~ pd_8_)  &  (~ pd_18_)  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  (~ pd_18_)  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire321 = ( (~ pdata_38_)  &  pc_20_  &  pc_5_  &  pdata_39_ ) | ( pdata_38_  &  pc_20_  &  (~ pc_5_)  &  pdata_39_ ) | ( (~ pdata_38_)  &  (~ pc_20_)  &  pc_5_  &  (~ pdata_39_) ) | ( pdata_38_  &  (~ pc_20_)  &  (~ pc_5_)  &  (~ pdata_39_) ) ;
 assign wire322 = ( wire462 ) | ( wire463 ) | ( wire1435 ) | ( wire8150 ) ;
 assign wire405 = ( wire1444 ) | ( wire1445 ) | ( wire1446 ) | ( wire1447 ) ;
 assign wire523 = ( (~ pdata_38_)  &  (~ pc_20_)  &  pc_5_  &  pdata_39_ ) | ( pdata_38_  &  (~ pc_20_)  &  (~ pc_5_)  &  pdata_39_ ) | ( (~ pdata_38_)  &  pc_20_  &  pc_5_  &  (~ pdata_39_) ) | ( pdata_38_  &  pc_20_  &  (~ pc_5_)  &  (~ pdata_39_) ) ;
 assign wire533 = ( pdata_37_  &  pdata_40_  &  pc_9_  &  pc_14_ ) | ( pdata_37_  &  (~ pdata_40_)  &  (~ pc_9_)  &  pc_14_ ) | ( (~ pdata_37_)  &  pdata_40_  &  pc_9_  &  (~ pc_14_) ) | ( (~ pdata_37_)  &  (~ pdata_40_)  &  (~ pc_9_)  &  (~ pc_14_) ) ;
 assign wire606 = ( pdata_36_  &  pc_27_  &  wire320 ) | ( (~ pdata_36_)  &  (~ pc_27_)  &  wire320 ) ;
 assign wire312 = ( pdata_43_  &  pc_25_  &  wire525 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire525 ) ;
 assign wire431 = ( (~ pdata_41_)  &  pc_11_  &  wire247  &  wire302 ) | ( pdata_41_  &  (~ pc_11_)  &  wire247  &  wire302 ) ;
 assign wire508 = ( pdata_44_  &  pdata_42_  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  (~ pc_7_)  &  pc_3_ ) | ( pdata_44_  &  (~ pdata_42_)  &  pc_7_  &  (~ pc_3_) ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign wire549 = ( (~ pdata_40_)  &  (~ pc_22_)  &  pc_18_  &  pdata_39_ ) | ( pdata_40_  &  (~ pc_22_)  &  (~ pc_18_)  &  pdata_39_ ) | ( (~ pdata_40_)  &  pc_22_  &  pc_18_  &  (~ pdata_39_) ) | ( pdata_40_  &  pc_22_  &  (~ pc_18_)  &  (~ pdata_39_) ) ;
 assign wire654 = ( (~ n_n1709)  &  (~ n_n1712)  &  (~ n_n1711) ) | ( n_n1709  &  (~ n_n1710)  &  n_n1712  &  n_n1711 ) | ( n_n1709  &  n_n1710  &  (~ n_n1712)  &  n_n1711 ) | ( n_n1709  &  n_n1710  &  n_n1712  &  (~ n_n1711) ) ;
 assign wire653 = ( (~ pdata_41_)  &  pc_11_  &  (~ n_n1711) ) | ( pdata_41_  &  (~ pc_11_)  &  (~ n_n1711) ) | ( pdata_41_  &  pc_11_  &  (~ n_n1712)  &  n_n1711 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  (~ n_n1712)  &  n_n1711 ) ;
 assign wire245 = ( (~ pd_4_)  &  pd_1_  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  (~ pd_1_)  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  (~ pdata_51_)  &  pdata_55_ ) | ( (~ pd_4_)  &  (~ pd_1_)  &  (~ pdata_51_)  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  (~ pd_1_)  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  pd_1_  &  (~ pdata_51_)  &  (~ pdata_55_) ) | ( pd_4_  &  (~ pd_1_)  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire305 = ( pd_11_  &  pd_16_  &  pdata_54_  &  pdata_52_ ) | ( pd_11_  &  (~ pd_16_)  &  (~ pdata_54_)  &  pdata_52_ ) | ( (~ pd_11_)  &  pd_16_  &  pdata_54_  &  (~ pdata_52_) ) | ( (~ pd_11_)  &  (~ pd_16_)  &  (~ pdata_54_)  &  (~ pdata_52_) ) ;
 assign wire313 = ( (~ pd_22_)  &  (~ pd_19_)  &  pdata_53_  &  pdata_56_ ) | ( pd_22_  &  (~ pd_19_)  &  (~ pdata_53_)  &  pdata_56_ ) | ( (~ pd_22_)  &  pd_19_  &  pdata_53_  &  (~ pdata_56_) ) | ( pd_22_  &  pd_19_  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire324 = ( wire469 ) | ( wire477 ) | ( wire481 ) ;
 assign wire407 = ( wire1969 ) | ( wire1970 ) | ( wire528  &  wire729 ) ;
 assign wire517 = ( pd_22_  &  pd_19_  &  pdata_53_  &  pdata_56_ ) | ( (~ pd_22_)  &  pd_19_  &  (~ pdata_53_)  &  pdata_56_ ) | ( pd_22_  &  (~ pd_19_)  &  pdata_53_  &  (~ pdata_56_) ) | ( (~ pd_22_)  &  (~ pd_19_)  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire528 = ( (~ pd_4_)  &  (~ pd_1_)  &  pdata_51_  &  pdata_55_ ) | ( (~ pd_4_)  &  pd_1_  &  (~ pdata_51_)  &  pdata_55_ ) | ( pd_4_  &  (~ pd_1_)  &  pdata_51_  &  (~ pdata_55_) ) | ( pd_4_  &  pd_1_  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire655 = ( (~ n_n1714)  &  (~ n_n1716)  &  (~ n_n1713) ) | ( (~ n_n1714)  &  (~ n_n1716)  &  (~ n_n1718) ) | ( (~ n_n1714)  &  (~ n_n1713)  &  (~ n_n1718) ) ;
 assign wire496 = ( pdata_36_  &  pc_4_ ) | ( (~ pdata_36_)  &  (~ pc_4_) ) | ( pdata_35_  &  pc_0_ ) | ( (~ pdata_35_)  &  (~ pc_0_) ) ;
 assign n_n1758 = ( wire275 ) | ( wire1699 ) | ( wire8018 ) | ( wire8019 ) ;
 assign wire662 = ( wire892 ) | ( wire894 ) | ( (~ n_n1703)  &  wire663 ) ;
 assign wire268 = ( pdata_35_  &  pdata_37_  &  pc_14_  &  pc_2_ ) | ( (~ pdata_35_)  &  (~ pdata_37_)  &  pc_14_  &  pc_2_ ) | ( (~ pdata_35_)  &  pdata_37_  &  (~ pc_14_)  &  pc_2_ ) | ( pdata_35_  &  (~ pdata_37_)  &  (~ pc_14_)  &  pc_2_ ) | ( (~ pdata_35_)  &  pdata_37_  &  pc_14_  &  (~ pc_2_) ) | ( pdata_35_  &  (~ pdata_37_)  &  pc_14_  &  (~ pc_2_) ) | ( pdata_35_  &  pdata_37_  &  (~ pc_14_)  &  (~ pc_2_) ) | ( (~ pdata_35_)  &  (~ pdata_37_)  &  (~ pc_14_)  &  (~ pc_2_) ) ;
 assign wire320 = ( (~ pdata_37_)  &  pdata_40_  &  pc_9_  &  pc_14_ ) | ( (~ pdata_37_)  &  (~ pdata_40_)  &  (~ pc_9_)  &  pc_14_ ) | ( pdata_37_  &  pdata_40_  &  pc_9_  &  (~ pc_14_) ) | ( pdata_37_  &  (~ pdata_40_)  &  (~ pc_9_)  &  (~ pc_14_) ) ;
 assign wire664 = ( pdata_35_  &  pc_2_  &  n_n1688  &  n_n1683 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  n_n1688  &  n_n1683 ) | ( (~ pdata_35_)  &  pc_2_  &  n_n1688  &  (~ n_n1683) ) | ( pdata_35_  &  (~ pc_2_)  &  n_n1688  &  (~ n_n1683) ) ;
 assign wire669 = ( wire2175 ) | ( wire7795 ) | ( (~ n_n1699)  &  wire670 ) ;
 assign wire666 = ( wire2167 ) | ( wire2169 ) | ( n_n1700  &  wire667 ) ;
 assign wire279 = ( wire1630 ) | ( wire1631 ) | ( wire1632 ) | ( wire8062 ) ;
 assign wire309 = ( (~ pdata_48_)  &  (~ pdata_44_)  &  pc_6_  &  pc_1_ ) | ( (~ pdata_48_)  &  pdata_44_  &  (~ pc_6_)  &  pc_1_ ) | ( pdata_48_  &  (~ pdata_44_)  &  pc_6_  &  (~ pc_1_) ) | ( pdata_48_  &  pdata_44_  &  (~ pc_6_)  &  (~ pc_1_) ) ;
 assign wire380 = ( pdata_46_  &  pc_19_  &  n_n1692  &  wire285 ) | ( (~ pdata_46_)  &  (~ pc_19_)  &  n_n1692  &  wire285 ) ;
 assign wire409 = ( pdata_44_  &  pc_6_  &  wire286  &  wire8088 ) | ( (~ pdata_44_)  &  (~ pc_6_)  &  wire286  &  wire8088 ) ;
 assign wire432 = ( (~ pdata_48_)  &  pc_1_  &  wire310  &  wire301 ) | ( pdata_48_  &  (~ pc_1_)  &  wire310  &  wire301 ) ;
 assign wire468 = ( wire1574 ) | ( wire1576 ) | ( wire309  &  wire736 ) ;
 assign wire476 = ( wire524  &  wire745 ) | ( wire535  &  wire744 ) ;
 assign wire574 = ( (~ pdata_45_)  &  (~ pdata_43_)  &  pc_15_  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_43_  &  (~ pc_15_)  &  pc_26_ ) | ( pdata_45_  &  (~ pdata_43_)  &  pc_15_  &  (~ pc_26_) ) | ( pdata_45_  &  pdata_43_  &  (~ pc_15_)  &  (~ pc_26_) ) ;
 assign wire673 = ( n_n1690  &  n_n1694  &  (~ n_n1691)  &  (~ n_n1692) ) | ( (~ n_n1690)  &  (~ n_n1694)  &  (~ n_n1691)  &  (~ n_n1692) ) ;
 assign wire672 = ( (~ n_n1690)  &  (~ n_n1691)  &  n_n1693 ) | ( (~ n_n1690)  &  (~ n_n1691)  &  (~ n_n1689) ) | ( n_n1690  &  n_n1691  &  n_n1693  &  (~ n_n1689) ) ;
 assign wire263 = ( pdata_45_  &  pdata_43_  &  pc_15_  &  pc_26_ ) | ( (~ pdata_45_)  &  (~ pdata_43_)  &  pc_15_  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_43_  &  (~ pc_15_)  &  pc_26_ ) | ( pdata_45_  &  (~ pdata_43_)  &  (~ pc_15_)  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_43_  &  pc_15_  &  (~ pc_26_) ) | ( pdata_45_  &  (~ pdata_43_)  &  pc_15_  &  (~ pc_26_) ) | ( pdata_45_  &  pdata_43_  &  (~ pc_15_)  &  (~ pc_26_) ) | ( (~ pdata_45_)  &  (~ pdata_43_)  &  (~ pc_15_)  &  (~ pc_26_) ) ;
 assign wire285 = ( (~ pdata_47_)  &  pdata_43_  &  pc_12_  &  pc_15_ ) | ( pdata_47_  &  pdata_43_  &  (~ pc_12_)  &  pc_15_ ) | ( (~ pdata_47_)  &  (~ pdata_43_)  &  pc_12_  &  (~ pc_15_) ) | ( pdata_47_  &  (~ pdata_43_)  &  (~ pc_12_)  &  (~ pc_15_) ) ;
 assign wire286 = ( pdata_45_  &  (~ pdata_43_)  &  pc_15_  &  pc_26_ ) | ( pdata_45_  &  pdata_43_  &  (~ pc_15_)  &  pc_26_ ) | ( (~ pdata_45_)  &  (~ pdata_43_)  &  pc_15_  &  (~ pc_26_) ) | ( (~ pdata_45_)  &  pdata_43_  &  (~ pc_15_)  &  (~ pc_26_) ) ;
 assign wire331 = ( pdata_47_  &  pc_12_  &  (~ n_n1691) ) | ( (~ pdata_47_)  &  (~ pc_12_)  &  (~ n_n1691) ) | ( (~ pdata_47_)  &  pc_12_  &  n_n1691  &  n_n1689 ) | ( pdata_47_  &  (~ pc_12_)  &  n_n1691  &  n_n1689 ) ;
 assign wire678 = ( n_n1691  &  (~ n_n1693)  &  n_n1692 ) | ( n_n1691  &  (~ n_n1693)  &  (~ n_n1689) ) | ( (~ n_n1693)  &  n_n1692  &  (~ n_n1689) ) ;
 assign wire677 = ( (~ n_n1690)  &  n_n1691  &  n_n1693  &  n_n1689 ) | ( n_n1690  &  (~ n_n1691)  &  n_n1693  &  (~ n_n1689) ) ;
 assign wire284 = ( pd_4_  &  pd_1_  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  (~ pd_1_)  &  (~ pdata_51_)  &  pdata_55_ ) | ( (~ pd_4_)  &  pd_1_  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  (~ pd_1_)  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire379 = ( (~ pd_16_)  &  pdata_54_  &  wire313  &  wire284 ) | ( pd_16_  &  (~ pdata_54_)  &  wire313  &  wire284 ) ;
 assign wire411 = ( wire1111 ) | ( wire1112 ) | ( wire1113 ) | ( wire1114 ) ;
 assign wire505 = ( (~ pd_4_)  &  pd_1_  &  pdata_51_  &  pdata_55_ ) | ( (~ pd_4_)  &  (~ pd_1_)  &  (~ pdata_51_)  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  pdata_51_  &  (~ pdata_55_) ) | ( pd_4_  &  (~ pd_1_)  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire540 = ( pd_11_  &  (~ pd_16_)  &  pdata_54_  &  pdata_52_ ) | ( pd_11_  &  pd_16_  &  (~ pdata_54_)  &  pdata_52_ ) | ( (~ pd_11_)  &  (~ pd_16_)  &  pdata_54_  &  (~ pdata_52_) ) | ( (~ pd_11_)  &  pd_16_  &  (~ pdata_54_)  &  (~ pdata_52_) ) ;
 assign wire680 = ( n_n1715  &  (~ n_n1713)  &  n_n1717 ) | ( (~ n_n1715)  &  n_n1716  &  (~ n_n1713)  &  (~ n_n1717) ) ;
 assign wire273 = ( wire407 ) | ( wire411 ) | ( wire8364 ) ;
 assign wire274 = ( (~ pd_19_)  &  pd_16_  &  pdata_54_  &  pdata_56_ ) | ( pd_19_  &  (~ pd_16_)  &  pdata_54_  &  pdata_56_ ) | ( pd_19_  &  pd_16_  &  (~ pdata_54_)  &  pdata_56_ ) | ( (~ pd_19_)  &  (~ pd_16_)  &  (~ pdata_54_)  &  pdata_56_ ) | ( pd_19_  &  pd_16_  &  pdata_54_  &  (~ pdata_56_) ) | ( (~ pd_19_)  &  (~ pd_16_)  &  pdata_54_  &  (~ pdata_56_) ) | ( (~ pd_19_)  &  pd_16_  &  (~ pdata_54_)  &  (~ pdata_56_) ) | ( pd_19_  &  (~ pd_16_)  &  (~ pdata_54_)  &  (~ pdata_56_) ) ;
 assign wire469 = ( wire1981 ) | ( wire1982 ) | ( wire1983 ) ;
 assign wire558 = ( pd_22_  &  (~ pd_19_)  &  pdata_53_  &  pdata_56_ ) | ( (~ pd_22_)  &  (~ pd_19_)  &  (~ pdata_53_)  &  pdata_56_ ) | ( pd_22_  &  pd_19_  &  pdata_53_  &  (~ pdata_56_) ) | ( (~ pd_22_)  &  pd_19_  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire684 = ( n_n1715  &  n_n1714  &  n_n1718  &  n_n1717 ) | ( n_n1715  &  (~ n_n1714)  &  (~ n_n1718)  &  (~ n_n1717) ) ;
 assign wire683 = ( n_n1715  &  (~ n_n1716)  &  n_n1713  &  (~ n_n1717) ) | ( (~ n_n1715)  &  n_n1716  &  (~ n_n1713)  &  (~ n_n1717) ) ;
 assign wire316 = ( (~ pd_0_)  &  pdata_63_  &  wire562 ) | ( pd_0_  &  (~ pdata_63_)  &  wire562 ) ;
 assign wire338 = ( wire1758 ) | ( wire1759 ) | ( wire1760 ) | ( wire1761 ) ;
 assign wire439 = ( wire297  &  wire7996 ) ;
 assign wire506 = ( pdata_59_  &  (~ pd_21_)  &  pd_17_  &  pdata_61_ ) | ( (~ pdata_59_)  &  (~ pd_21_)  &  (~ pd_17_)  &  pdata_61_ ) | ( pdata_59_  &  pd_21_  &  pd_17_  &  (~ pdata_61_) ) | ( (~ pdata_59_)  &  pd_21_  &  (~ pd_17_)  &  (~ pdata_61_) ) ;
 assign wire543 = ( pd_21_  &  pdata_60_  &  pd_13_  &  pdata_61_ ) | ( pd_21_  &  (~ pdata_60_)  &  (~ pd_13_)  &  pdata_61_ ) | ( (~ pd_21_)  &  pdata_60_  &  pd_13_  &  (~ pdata_61_) ) | ( (~ pd_21_)  &  (~ pdata_60_)  &  (~ pd_13_)  &  (~ pdata_61_) ) ;
 assign wire588 = ( (~ pdata_32_)  &  pd_7_  &  pd_3_  &  pdata_62_ ) | ( pdata_32_  &  pd_7_  &  (~ pd_3_)  &  pdata_62_ ) | ( (~ pdata_32_)  &  (~ pd_7_)  &  pd_3_  &  (~ pdata_62_) ) | ( pdata_32_  &  (~ pd_7_)  &  (~ pd_3_)  &  (~ pdata_62_) ) ;
 assign wire283 = ( pd_8_  &  pd_18_  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  (~ pdata_50_)  &  pdata_51_ ) | ( pd_8_  &  (~ pd_18_)  &  pdata_50_  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  (~ pd_18_)  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire304 = ( (~ pdata_48_)  &  pd_23_  &  pd_26_  &  pdata_52_ ) | ( pdata_48_  &  (~ pd_23_)  &  pd_26_  &  pdata_52_ ) | ( (~ pdata_48_)  &  pd_23_  &  (~ pd_26_)  &  (~ pdata_52_) ) | ( pdata_48_  &  (~ pd_23_)  &  (~ pd_26_)  &  (~ pdata_52_) ) ;
 assign wire420 = ( (~ pdata_47_)  &  pd_12_ ) | ( pdata_47_  &  (~ pd_12_) ) | ( pd_2_  &  pdata_49_ ) | ( (~ pd_2_)  &  (~ pdata_49_) ) ;
 assign wire504 = ( pd_8_  &  (~ pd_18_)  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  (~ pd_18_)  &  (~ pdata_50_)  &  pdata_51_ ) | ( pd_8_  &  pd_18_  &  pdata_50_  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  pd_18_  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire579 = ( (~ pdata_47_)  &  pd_12_  &  (~ pd_2_)  &  pdata_49_ ) | ( pdata_47_  &  (~ pd_12_)  &  (~ pd_2_)  &  pdata_49_ ) | ( (~ pdata_47_)  &  pd_12_  &  pd_2_  &  (~ pdata_49_) ) | ( pdata_47_  &  (~ pd_12_)  &  pd_2_  &  (~ pdata_49_) ) ;
 assign wire310 = ( (~ pdata_45_)  &  pdata_44_  &  pc_6_  &  pc_26_ ) | ( (~ pdata_45_)  &  (~ pdata_44_)  &  (~ pc_6_)  &  pc_26_ ) | ( pdata_45_  &  pdata_44_  &  pc_6_  &  (~ pc_26_) ) | ( pdata_45_  &  (~ pdata_44_)  &  (~ pc_6_)  &  (~ pc_26_) ) ;
 assign wire433 = ( pdata_47_  &  pc_12_  &  wire309  &  wire286 ) | ( (~ pdata_47_)  &  (~ pc_12_)  &  wire309  &  wire286 ) ;
 assign wire534 = ( (~ pdata_47_)  &  pdata_46_  &  pc_12_  &  pc_19_ ) | ( pdata_47_  &  pdata_46_  &  (~ pc_12_)  &  pc_19_ ) | ( (~ pdata_47_)  &  (~ pdata_46_)  &  pc_12_  &  (~ pc_19_) ) | ( pdata_47_  &  (~ pdata_46_)  &  (~ pc_12_)  &  (~ pc_19_) ) ;
 assign wire535 = ( (~ pdata_43_)  &  pc_15_  &  wire310 ) | ( pdata_43_  &  (~ pc_15_)  &  wire310 ) ;
 assign wire689 = ( (~ n_n1690)  &  (~ n_n1691)  &  n_n1689 ) | ( (~ n_n1690)  &  n_n1691  &  (~ n_n1689) ) | ( n_n1690  &  (~ n_n1691)  &  n_n1693  &  (~ n_n1689) ) ;
 assign wire688 = ( n_n1691  &  (~ n_n1693)  &  (~ n_n1692) ) | ( n_n1691  &  n_n1692  &  n_n1689 ) | ( n_n1691  &  (~ n_n1692)  &  (~ n_n1689) ) ;
 assign wire246 = ( pdata_59_  &  pd_5_  &  pd_15_  &  pdata_55_ ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  pd_15_  &  pdata_55_ ) | ( (~ pdata_59_)  &  pd_5_  &  (~ pd_15_)  &  pdata_55_ ) | ( pdata_59_  &  (~ pd_5_)  &  (~ pd_15_)  &  pdata_55_ ) | ( (~ pdata_59_)  &  pd_5_  &  pd_15_  &  (~ pdata_55_) ) | ( pdata_59_  &  (~ pd_5_)  &  pd_15_  &  (~ pdata_55_) ) | ( pdata_59_  &  pd_5_  &  (~ pd_15_)  &  (~ pdata_55_) ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  (~ pd_15_)  &  (~ pdata_55_) ) ;
 assign wire271 = ( (~ pd_10_)  &  pdata_60_  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  (~ pdata_60_)  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  pdata_60_  &  (~ pd_24_)  &  pdata_57_ ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  (~ pd_24_)  &  pdata_57_ ) | ( pd_10_  &  pdata_60_  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  pdata_60_  &  (~ pd_24_)  &  (~ pdata_57_) ) | ( pd_10_  &  (~ pdata_60_)  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire585 = ( pd_20_  &  pd_27_  &  pdata_58_  &  pdata_56_ ) | ( pd_20_  &  (~ pd_27_)  &  (~ pdata_58_)  &  pdata_56_ ) | ( (~ pd_20_)  &  pd_27_  &  pdata_58_  &  (~ pdata_56_) ) | ( (~ pd_20_)  &  (~ pd_27_)  &  (~ pdata_58_)  &  (~ pdata_56_) ) ;
 assign wire692 = ( n_n1723  &  n_n1724  &  (~ n_n1720)  &  n_n1721 ) | ( n_n1723  &  (~ n_n1724)  &  n_n1720  &  (~ n_n1721) ) ;
 assign wire691 = ( n_n1723  &  n_n1724  &  n_n1720  &  (~ n_n1721) ) | ( (~ n_n1723)  &  n_n1724  &  (~ n_n1720)  &  (~ n_n1721) ) ;
 assign wire267 = ( pdata_41_  &  pc_11_  &  n_n1712  &  n_n1711 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  n_n1712  &  n_n1711 ) | ( (~ pdata_41_)  &  pc_11_  &  (~ n_n1712)  &  n_n1711 ) | ( pdata_41_  &  (~ pc_11_)  &  (~ n_n1712)  &  n_n1711 ) | ( (~ pdata_41_)  &  pc_11_  &  n_n1712  &  (~ n_n1711) ) | ( pdata_41_  &  (~ pc_11_)  &  n_n1712  &  (~ n_n1711) ) ;
 assign wire473 = ( wire1508 ) | ( wire1509 ) | ( wire1510 ) ;
 assign wire696 = ( wire1503 ) | ( wire1505 ) | ( n_n1708  &  wire697 ) ;
 assign n_n1731 = ( wire7952 ) | ( wire7953 ) | ( wire8130 ) | ( wire8131 ) ;
 assign wire302 = ( pdata_40_  &  pc_22_  &  pc_18_  &  pdata_39_ ) | ( (~ pdata_40_)  &  pc_22_  &  (~ pc_18_)  &  pdata_39_ ) | ( pdata_40_  &  (~ pc_22_)  &  pc_18_  &  (~ pdata_39_) ) | ( (~ pdata_40_)  &  (~ pc_22_)  &  (~ pc_18_)  &  (~ pdata_39_) ) ;
 assign wire426 = ( (~ pdata_40_)  &  pc_18_  &  wire7943  &  wire7962 ) | ( pdata_40_  &  (~ pc_18_)  &  wire7943  &  wire7962 ) ;
 assign wire474 = ( wire1818 ) | ( wire1819 ) | ( wire508  &  wire742 ) ;
 assign wire503 = ( pdata_41_  &  (~ pdata_40_)  &  pc_11_  &  pc_18_ ) | ( (~ pdata_41_)  &  (~ pdata_40_)  &  (~ pc_11_)  &  pc_18_ ) | ( pdata_41_  &  pdata_40_  &  pc_11_  &  (~ pc_18_) ) | ( (~ pdata_41_)  &  pdata_40_  &  (~ pc_11_)  &  (~ pc_18_) ) ;
 assign wire526 = ( pdata_40_  &  (~ pc_22_)  &  pc_18_  &  pdata_39_ ) | ( (~ pdata_40_)  &  (~ pc_22_)  &  (~ pc_18_)  &  pdata_39_ ) | ( pdata_40_  &  pc_22_  &  pc_18_  &  (~ pdata_39_) ) | ( (~ pdata_40_)  &  pc_22_  &  (~ pc_18_)  &  (~ pdata_39_) ) ;
 assign wire536 = ( pdata_44_  &  (~ pdata_42_)  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  (~ pc_7_)  &  pc_3_ ) | ( pdata_44_  &  pdata_42_  &  pc_7_  &  (~ pc_3_) ) | ( (~ pdata_44_)  &  pdata_42_  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign n_n1737 = ( wire7952 ) | ( wire7953 ) | ( wire7966 ) | ( wire7967 ) ;
 assign wire265 = ( (~ pdata_59_)  &  pd_21_  &  pd_17_  &  pdata_61_ ) | ( pdata_59_  &  (~ pd_21_)  &  pd_17_  &  pdata_61_ ) | ( pdata_59_  &  pd_21_  &  (~ pd_17_)  &  pdata_61_ ) | ( (~ pdata_59_)  &  (~ pd_21_)  &  (~ pd_17_)  &  pdata_61_ ) | ( pdata_59_  &  pd_21_  &  pd_17_  &  (~ pdata_61_) ) | ( (~ pdata_59_)  &  (~ pd_21_)  &  pd_17_  &  (~ pdata_61_) ) | ( (~ pdata_59_)  &  pd_21_  &  (~ pd_17_)  &  (~ pdata_61_) ) | ( pdata_59_  &  (~ pd_21_)  &  (~ pd_17_)  &  (~ pdata_61_) ) ;
 assign wire381 = ( pd_0_  &  pdata_63_  &  wire531  &  wire506 ) | ( (~ pd_0_)  &  (~ pdata_63_)  &  wire531  &  wire506 ) ;
 assign wire701 = ( (~ n_n1726)  &  n_n1728  &  n_n1730  &  n_n1729 ) | ( (~ n_n1726)  &  (~ n_n1728)  &  (~ n_n1730)  &  n_n1729 ) | ( n_n1726  &  (~ n_n1728)  &  n_n1730  &  (~ n_n1729) ) | ( n_n1726  &  n_n1728  &  (~ n_n1730)  &  (~ n_n1729) ) ;
 assign wire700 = ( n_n1728  &  n_n1730  &  n_n1729 ) | ( (~ n_n1726)  &  (~ n_n1728)  &  (~ n_n1730)  &  (~ n_n1729) ) ;
 assign wire301 = ( pdata_47_  &  pdata_46_  &  pc_12_  &  pc_19_ ) | ( (~ pdata_47_)  &  pdata_46_  &  (~ pc_12_)  &  pc_19_ ) | ( pdata_47_  &  (~ pdata_46_)  &  pc_12_  &  (~ pc_19_) ) | ( (~ pdata_47_)  &  (~ pdata_46_)  &  (~ pc_12_)  &  (~ pc_19_) ) ;
 assign wire308 = ( pdata_48_  &  (~ pdata_46_)  &  pc_19_  &  pc_1_ ) | ( pdata_48_  &  pdata_46_  &  (~ pc_19_)  &  pc_1_ ) | ( (~ pdata_48_)  &  (~ pdata_46_)  &  pc_19_  &  (~ pc_1_) ) | ( (~ pdata_48_)  &  pdata_46_  &  (~ pc_19_)  &  (~ pc_1_) ) ;
 assign wire524 = ( pdata_45_  &  pdata_44_  &  pc_6_  &  pc_26_ ) | ( pdata_45_  &  (~ pdata_44_)  &  (~ pc_6_)  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_44_  &  pc_6_  &  (~ pc_26_) ) | ( (~ pdata_45_)  &  (~ pdata_44_)  &  (~ pc_6_)  &  (~ pc_26_) ) ;
 assign wire546 = ( (~ pdata_46_)  &  pc_19_  &  wire309 ) | ( pdata_46_  &  (~ pc_19_)  &  wire309 ) ;
 assign wire477 = ( wire1977 ) | ( wire1978 ) | ( wire1979 ) | ( wire1980 ) ;
 assign wire582 = ( pd_19_  &  (~ pd_16_)  &  pdata_54_  &  pdata_56_ ) | ( pd_19_  &  pd_16_  &  (~ pdata_54_)  &  pdata_56_ ) | ( (~ pd_19_)  &  (~ pd_16_)  &  pdata_54_  &  (~ pdata_56_) ) | ( (~ pd_19_)  &  pd_16_  &  (~ pdata_54_)  &  (~ pdata_56_) ) ;
 assign wire705 = ( wire835 ) | ( wire836 ) | ( (~ n_n1717)  &  wire706 ) ;
 assign wire295 = ( pd_7_  &  (~ pd_0_)  &  pdata_62_  &  pdata_63_ ) | ( (~ pd_7_)  &  (~ pd_0_)  &  (~ pdata_62_)  &  pdata_63_ ) | ( pd_7_  &  pd_0_  &  pdata_62_  &  (~ pdata_63_) ) | ( (~ pd_7_)  &  pd_0_  &  (~ pdata_62_)  &  (~ pdata_63_) ) ;
 assign wire413 = ( wire2048 ) | ( wire2049 ) | ( wire2050 ) | ( wire2051 ) ;
 assign wire708 = ( wire280 ) | ( wire1753 ) | ( wire1754 ) | ( wire1756 ) ;
 assign wire559 = ( (~ pdata_59_)  &  pd_5_  &  wire306 ) | ( pdata_59_  &  (~ pd_5_)  &  wire306 ) ;
 assign wire710 = ( n_n1723  &  n_n1724  &  (~ n_n1722) ) | ( n_n1723  &  (~ n_n1722)  &  (~ n_n1721) ) | ( (~ n_n1723)  &  (~ n_n1724)  &  (~ n_n1722)  &  n_n1721 ) ;
 assign wire709 = ( n_n1723  &  (~ n_n1719)  &  n_n1722  &  n_n1721 ) | ( n_n1723  &  n_n1719  &  n_n1722  &  (~ n_n1721) ) ;
 assign wire509 = ( pd_4_  &  (~ pd_1_)  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  (~ pdata_51_)  &  pdata_55_ ) | ( (~ pd_4_)  &  (~ pd_1_)  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  pd_1_  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire516 = ( pdata_48_  &  pd_23_  &  (~ pd_26_)  &  pdata_52_ ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  (~ pd_26_)  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  pd_26_  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  pd_26_  &  (~ pdata_52_) ) ;
 assign wire261 = ( (~ pdata_48_)  &  pd_23_  &  pd_26_  &  pdata_52_ ) | ( pdata_48_  &  (~ pd_23_)  &  pd_26_  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  (~ pd_26_)  &  pdata_52_ ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  (~ pd_26_)  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  pd_26_  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  pd_26_  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  pd_23_  &  (~ pd_26_)  &  (~ pdata_52_) ) | ( pdata_48_  &  (~ pd_23_)  &  (~ pd_26_)  &  (~ pdata_52_) ) ;
 assign wire262 = ( (~ pdata_47_)  &  pd_12_  &  pd_18_  &  pdata_51_ ) | ( pdata_47_  &  (~ pd_12_)  &  pd_18_  &  pdata_51_ ) | ( pdata_47_  &  pd_12_  &  (~ pd_18_)  &  pdata_51_ ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  (~ pd_18_)  &  pdata_51_ ) | ( pdata_47_  &  pd_12_  &  pd_18_  &  (~ pdata_51_) ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  pd_18_  &  (~ pdata_51_) ) | ( (~ pdata_47_)  &  pd_12_  &  (~ pd_18_)  &  (~ pdata_51_) ) | ( pdata_47_  &  (~ pd_12_)  &  (~ pd_18_)  &  (~ pdata_51_) ) ;
 assign wire532 = ( (~ pdata_35_)  &  pdata_36_  &  pc_4_  &  pc_0_ ) | ( (~ pdata_35_)  &  (~ pdata_36_)  &  (~ pc_4_)  &  pc_0_ ) | ( pdata_35_  &  pdata_36_  &  pc_4_  &  (~ pc_0_) ) | ( pdata_35_  &  (~ pdata_36_)  &  (~ pc_4_)  &  (~ pc_0_) ) ;
 assign wire598 = ( (~ pdata_35_)  &  (~ pdata_37_)  &  pc_14_  &  pc_2_ ) | ( (~ pdata_35_)  &  pdata_37_  &  (~ pc_14_)  &  pc_2_ ) | ( pdata_35_  &  (~ pdata_37_)  &  pc_14_  &  (~ pc_2_) ) | ( pdata_35_  &  pdata_37_  &  (~ pc_14_)  &  (~ pc_2_) ) ;
 assign wire519 = ( pdata_34_  &  (~ pc_13_)  &  pc_23_  &  pdata_63_ ) | ( (~ pdata_34_)  &  (~ pc_13_)  &  (~ pc_23_)  &  pdata_63_ ) | ( pdata_34_  &  pc_13_  &  pc_23_  &  (~ pdata_63_) ) | ( (~ pdata_34_)  &  pc_13_  &  (~ pc_23_)  &  (~ pdata_63_) ) ;
 assign wire269 = ( (~ pdata_34_)  &  pc_13_  &  pc_23_  &  pdata_63_ ) | ( pdata_34_  &  (~ pc_13_)  &  pc_23_  &  pdata_63_ ) | ( pdata_34_  &  pc_13_  &  (~ pc_23_)  &  pdata_63_ ) | ( (~ pdata_34_)  &  (~ pc_13_)  &  (~ pc_23_)  &  pdata_63_ ) | ( pdata_34_  &  pc_13_  &  pc_23_  &  (~ pdata_63_) ) | ( (~ pdata_34_)  &  (~ pc_13_)  &  pc_23_  &  (~ pdata_63_) ) | ( (~ pdata_34_)  &  pc_13_  &  (~ pc_23_)  &  (~ pdata_63_) ) | ( pdata_34_  &  (~ pc_13_)  &  (~ pc_23_)  &  (~ pdata_63_) ) ;
 assign wire515 = ( pdata_43_  &  (~ pdata_41_)  &  pc_11_  &  pc_25_ ) | ( pdata_43_  &  pdata_41_  &  (~ pc_11_)  &  pc_25_ ) | ( (~ pdata_43_)  &  (~ pdata_41_)  &  pc_11_  &  (~ pc_25_) ) | ( (~ pdata_43_)  &  pdata_41_  &  (~ pc_11_)  &  (~ pc_25_) ) ;
 assign wire480 = ( wire1829 ) | ( wire1830 ) | ( wire515  &  wire749 ) ;
 assign wire481 = ( wire1973 ) | ( wire505  &  wire750 ) ;
 assign wire555 = ( (~ pd_11_)  &  pd_16_  &  pdata_54_  &  pdata_52_ ) | ( (~ pd_11_)  &  (~ pd_16_)  &  (~ pdata_54_)  &  pdata_52_ ) | ( pd_11_  &  pd_16_  &  pdata_54_  &  (~ pdata_52_) ) | ( pd_11_  &  (~ pd_16_)  &  (~ pdata_54_)  &  (~ pdata_52_) ) ;
 assign wire513 = ( (~ pdata_34_)  &  (~ pc_13_)  &  pc_23_  &  pdata_63_ ) | ( pdata_34_  &  (~ pc_13_)  &  (~ pc_23_)  &  pdata_63_ ) | ( (~ pdata_34_)  &  pc_13_  &  pc_23_  &  (~ pdata_63_) ) | ( pdata_34_  &  pc_13_  &  (~ pc_23_)  &  (~ pdata_63_) ) ;
 assign wire595 = ( (~ pdata_32_)  &  pdata_33_  &  pc_10_  &  pc_16_ ) | ( (~ pdata_32_)  &  (~ pdata_33_)  &  (~ pc_10_)  &  pc_16_ ) | ( pdata_32_  &  pdata_33_  &  pc_10_  &  (~ pc_16_) ) | ( pdata_32_  &  (~ pdata_33_)  &  (~ pc_10_)  &  (~ pc_16_) ) ;
 assign wire712 = ( n_n1706  &  (~ n_n1705)  &  n_n1703  &  wire592 ) | ( (~ n_n1706)  &  (~ n_n1705)  &  (~ n_n1703)  &  wire592 ) ;
 assign wire713 = ( (~ pd_21_)  &  pdata_61_  &  n_n1730  &  n_n1729 ) | ( pd_21_  &  (~ pdata_61_)  &  n_n1730  &  n_n1729 ) | ( pd_21_  &  pdata_61_  &  (~ n_n1730)  &  n_n1729 ) | ( (~ pd_21_)  &  (~ pdata_61_)  &  (~ n_n1730)  &  n_n1729 ) ;
 assign wire303 = ( (~ pd_8_)  &  (~ pd_18_)  &  pdata_50_  &  pdata_51_ ) | ( pd_8_  &  (~ pd_18_)  &  (~ pdata_50_)  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  pd_18_  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire510 = ( (~ pdata_59_)  &  pd_20_  &  pd_5_  &  pdata_56_ ) | ( pdata_59_  &  pd_20_  &  (~ pd_5_)  &  pdata_56_ ) | ( (~ pdata_59_)  &  (~ pd_20_)  &  pd_5_  &  (~ pdata_56_) ) | ( pdata_59_  &  (~ pd_20_)  &  (~ pd_5_)  &  (~ pdata_56_) ) ;
 assign wire715 = ( n_n1724  &  (~ n_n1720)  &  n_n1719  &  n_n1722 ) | ( (~ n_n1724)  &  (~ n_n1720)  &  n_n1719  &  (~ n_n1722) ) ;
 assign wire714 = ( n_n1724  &  (~ n_n1719)  &  n_n1722  &  n_n1721 ) | ( (~ n_n1724)  &  (~ n_n1719)  &  (~ n_n1722)  &  n_n1721 ) ;
 assign wire716 = ( (~ pdata_47_)  &  pc_12_  &  n_n1694  &  n_n1692 ) | ( pdata_47_  &  (~ pc_12_)  &  n_n1694  &  n_n1692 ) | ( pdata_47_  &  pc_12_  &  (~ n_n1694)  &  n_n1692 ) | ( (~ pdata_47_)  &  (~ pc_12_)  &  (~ n_n1694)  &  n_n1692 ) ;
 assign wire586 = ( pdata_59_  &  pd_5_  &  (~ pd_15_)  &  pdata_55_ ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  (~ pd_15_)  &  pdata_55_ ) | ( pdata_59_  &  pd_5_  &  pd_15_  &  (~ pdata_55_) ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  pd_15_  &  (~ pdata_55_) ) ;
 assign wire294 = ( (~ pd_27_)  &  pdata_58_  &  wire7731 ) | ( pd_27_  &  (~ pdata_58_)  &  wire7731 ) ;
 assign wire604 = ( pdata_38_  &  (~ pc_20_)  &  pc_5_  &  pdata_39_ ) | ( (~ pdata_38_)  &  (~ pc_20_)  &  (~ pc_5_)  &  pdata_39_ ) | ( pdata_38_  &  pc_20_  &  pc_5_  &  (~ pdata_39_) ) | ( (~ pdata_38_)  &  pc_20_  &  (~ pc_5_)  &  (~ pdata_39_) ) ;
 assign wire562 = ( (~ pdata_32_)  &  (~ pd_7_)  &  pd_3_  &  pdata_62_ ) | ( pdata_32_  &  (~ pd_7_)  &  (~ pd_3_)  &  pdata_62_ ) | ( (~ pdata_32_)  &  pd_7_  &  pd_3_  &  (~ pdata_62_) ) | ( pdata_32_  &  pd_7_  &  (~ pd_3_)  &  (~ pdata_62_) ) ;
 assign wire319 = ( (~ pdata_32_)  &  pc_16_  &  pc_13_  &  pdata_63_ ) | ( pdata_32_  &  (~ pc_16_)  &  pc_13_  &  pdata_63_ ) | ( (~ pdata_32_)  &  pc_16_  &  (~ pc_13_)  &  (~ pdata_63_) ) | ( pdata_32_  &  (~ pc_16_)  &  (~ pc_13_)  &  (~ pdata_63_) ) ;
 assign wire717 = ( (~ n_n1704)  &  n_n1706  &  n_n1705  &  n_n1703 ) | ( n_n1704  &  (~ n_n1706)  &  n_n1705  &  n_n1703 ) ;
 assign wire718 = ( pd_20_  &  pdata_56_  &  n_n1720  &  n_n1719 ) | ( (~ pd_20_)  &  (~ pdata_56_)  &  n_n1720  &  n_n1719 ) | ( (~ pd_20_)  &  pdata_56_  &  n_n1720  &  (~ n_n1719) ) | ( pd_20_  &  (~ pdata_56_)  &  n_n1720  &  (~ n_n1719) ) ;
 assign wire539 = ( (~ pdata_47_)  &  pd_12_  &  pd_2_  &  pdata_49_ ) | ( pdata_47_  &  (~ pd_12_)  &  pd_2_  &  pdata_49_ ) | ( (~ pdata_47_)  &  pd_12_  &  (~ pd_2_)  &  (~ pdata_49_) ) | ( pdata_47_  &  (~ pd_12_)  &  (~ pd_2_)  &  (~ pdata_49_) ) ;
 assign wire719 = ( n_n1696  &  (~ n_n1699)  &  n_n1695  &  (~ n_n1697) ) | ( (~ n_n1696)  &  (~ n_n1699)  &  (~ n_n1695)  &  (~ n_n1697) ) ;
 assign wire520 = ( pdata_32_  &  pc_16_  &  pc_13_  &  pdata_63_ ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  pc_13_  &  pdata_63_ ) | ( pdata_32_  &  pc_16_  &  (~ pc_13_)  &  (~ pdata_63_) ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  (~ pc_13_)  &  (~ pdata_63_) ) ;
 assign wire527 = ( pdata_48_  &  pd_23_  &  pd_26_  &  pdata_52_ ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  pd_26_  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  (~ pd_26_)  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  (~ pd_26_)  &  (~ pdata_52_) ) ;
 assign wire427 = ( wire315  &  (~ wire417) ) ;
 assign wire725 = ( pd_15_  &  pdata_55_  &  n_n1719  &  n_n1722 ) | ( (~ pd_15_)  &  (~ pdata_55_)  &  n_n1719  &  n_n1722 ) | ( (~ pd_15_)  &  pdata_55_  &  (~ n_n1719)  &  (~ n_n1722) ) | ( pd_15_  &  (~ pdata_55_)  &  (~ n_n1719)  &  (~ n_n1722) ) ;
 assign wire726 = ( n_n1696  &  n_n1699  &  n_n1695  &  (~ n_n1697) ) | ( (~ n_n1696)  &  n_n1699  &  (~ n_n1695)  &  (~ n_n1697) ) ;
 assign wire484 = ( pdata_37_  &  pc_14_  &  n_n1686  &  wire523 ) | ( (~ pdata_37_)  &  (~ pc_14_)  &  n_n1686  &  wire523 ) ;
 assign wire729 = ( (~ n_n1715)  &  (~ n_n1716)  &  n_n1713  &  n_n1717 ) | ( (~ n_n1715)  &  (~ n_n1716)  &  (~ n_n1713)  &  (~ n_n1717) ) ;
 assign wire428 = ( wire306  &  wire7744 ) ;
 assign wire732 = ( (~ n_n1686)  &  n_n1688  &  (~ n_n1683)  &  n_n1685 ) | ( n_n1686  &  (~ n_n1688)  &  n_n1683  &  (~ n_n1685) ) ;
 assign wire569 = ( pdata_37_  &  (~ pdata_40_)  &  pc_9_  &  pc_14_ ) | ( pdata_37_  &  pdata_40_  &  (~ pc_9_)  &  pc_14_ ) | ( (~ pdata_37_)  &  (~ pdata_40_)  &  pc_9_  &  (~ pc_14_) ) | ( (~ pdata_37_)  &  pdata_40_  &  (~ pc_9_)  &  (~ pc_14_) ) ;
 assign wire567 = ( (~ pdata_33_)  &  (~ pdata_34_)  &  pc_10_  &  pc_23_ ) | ( pdata_33_  &  (~ pdata_34_)  &  (~ pc_10_)  &  pc_23_ ) | ( (~ pdata_33_)  &  pdata_34_  &  pc_10_  &  (~ pc_23_) ) | ( pdata_33_  &  pdata_34_  &  (~ pc_10_)  &  (~ pc_23_) ) ;
 assign wire734 = ( (~ n_n1704)  &  (~ n_n1706)  &  n_n1705  &  n_n1703 ) | ( (~ n_n1704)  &  n_n1706  &  n_n1705  &  (~ n_n1703) ) ;
 assign wire735 = ( n_n1696  &  n_n1700  &  n_n1697  &  n_n1698 ) | ( (~ n_n1696)  &  (~ n_n1700)  &  n_n1697  &  n_n1698 ) ;
 assign wire736 = ( n_n1690  &  n_n1694  &  (~ n_n1691)  &  n_n1692 ) | ( n_n1690  &  (~ n_n1694)  &  (~ n_n1691)  &  (~ n_n1692) ) ;
 assign wire737 = ( (~ pd_4_)  &  pd_1_  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  (~ pd_1_)  &  pdata_51_  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  (~ pdata_51_)  &  pdata_55_ ) | ( (~ pd_4_)  &  (~ pd_1_)  &  (~ pdata_51_)  &  pdata_55_ ) | ( pd_4_  &  pd_1_  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  (~ pd_1_)  &  pdata_51_  &  (~ pdata_55_) ) | ( (~ pd_4_)  &  pd_1_  &  (~ pdata_51_)  &  (~ pdata_55_) ) | ( pd_4_  &  (~ pd_1_)  &  (~ pdata_51_)  &  (~ pdata_55_) ) ;
 assign wire738 = ( (~ n_n1696)  &  (~ n_n1700)  &  n_n1697  &  n_n1698 ) | ( n_n1696  &  n_n1700  &  n_n1697  &  (~ n_n1698) ) ;
 assign wire740 = ( (~ n_n1724)  &  (~ n_n1719)  &  n_n1722  &  n_n1721 ) | ( n_n1724  &  (~ n_n1719)  &  (~ n_n1722)  &  n_n1721 ) ;
 assign wire739 = ( (~ n_n1723)  &  n_n1724  &  (~ n_n1720)  &  n_n1721 ) | ( (~ n_n1723)  &  (~ n_n1724)  &  (~ n_n1720)  &  (~ n_n1721) ) ;
 assign wire742 = ( (~ n_n1710)  &  n_n1712  &  (~ n_n1708)  &  n_n1711 ) | ( n_n1710  &  (~ n_n1712)  &  (~ n_n1708)  &  n_n1711 ) ;
 assign wire743 = ( pdata_32_  &  pd_7_  &  pd_3_  &  pdata_62_ ) | ( (~ pdata_32_)  &  (~ pd_7_)  &  pd_3_  &  pdata_62_ ) | ( (~ pdata_32_)  &  pd_7_  &  (~ pd_3_)  &  pdata_62_ ) | ( pdata_32_  &  (~ pd_7_)  &  (~ pd_3_)  &  pdata_62_ ) | ( (~ pdata_32_)  &  pd_7_  &  pd_3_  &  (~ pdata_62_) ) | ( pdata_32_  &  (~ pd_7_)  &  pd_3_  &  (~ pdata_62_) ) | ( pdata_32_  &  pd_7_  &  (~ pd_3_)  &  (~ pdata_62_) ) | ( (~ pdata_32_)  &  (~ pd_7_)  &  (~ pd_3_)  &  (~ pdata_62_) ) ;
 assign wire745 = ( (~ n_n1690)  &  (~ n_n1694)  &  (~ n_n1691)  &  n_n1689 ) | ( n_n1690  &  (~ n_n1694)  &  (~ n_n1691)  &  (~ n_n1689) ) ;
 assign wire744 = ( pdata_47_  &  pc_12_  &  n_n1691  &  n_n1689 ) | ( (~ pdata_47_)  &  (~ pc_12_)  &  n_n1691  &  n_n1689 ) | ( (~ pdata_47_)  &  pc_12_  &  n_n1691  &  (~ n_n1689) ) | ( pdata_47_  &  (~ pc_12_)  &  n_n1691  &  (~ n_n1689) ) ;
 assign wire747 = ( (~ n_n1723)  &  n_n1724  &  (~ n_n1720)  &  n_n1721 ) | ( (~ n_n1723)  &  (~ n_n1724)  &  n_n1720  &  (~ n_n1721) ) ;
 assign wire749 = ( n_n1709  &  (~ n_n1712)  &  n_n1707  &  n_n1711 ) | ( n_n1709  &  (~ n_n1712)  &  (~ n_n1707)  &  (~ n_n1711) ) ;
 assign wire751 = ( pd_22_  &  pd_19_  &  pdata_53_  &  pdata_56_ ) | ( (~ pd_22_)  &  (~ pd_19_)  &  pdata_53_  &  pdata_56_ ) | ( (~ pd_22_)  &  pd_19_  &  (~ pdata_53_)  &  pdata_56_ ) | ( pd_22_  &  (~ pd_19_)  &  (~ pdata_53_)  &  pdata_56_ ) | ( (~ pd_22_)  &  pd_19_  &  pdata_53_  &  (~ pdata_56_) ) | ( pd_22_  &  (~ pd_19_)  &  pdata_53_  &  (~ pdata_56_) ) | ( pd_22_  &  pd_19_  &  (~ pdata_53_)  &  (~ pdata_56_) ) | ( (~ pd_22_)  &  (~ pd_19_)  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire750 = ( (~ n_n1715)  &  (~ n_n1716)  &  n_n1713  &  (~ n_n1717) ) | ( n_n1715  &  (~ n_n1716)  &  (~ n_n1713)  &  (~ n_n1717) ) ;
 assign wire511 = ( pd_21_  &  (~ pdata_60_)  &  pd_13_  &  pdata_61_ ) | ( pd_21_  &  pdata_60_  &  (~ pd_13_)  &  pdata_61_ ) | ( (~ pd_21_)  &  (~ pdata_60_)  &  pd_13_  &  (~ pdata_61_) ) | ( (~ pd_21_)  &  pdata_60_  &  (~ pd_13_)  &  (~ pdata_61_) ) ;
 assign wire591 = ( (~ pdata_35_)  &  pdata_32_  &  pc_16_  &  pc_0_ ) | ( (~ pdata_35_)  &  (~ pdata_32_)  &  (~ pc_16_)  &  pc_0_ ) | ( pdata_35_  &  pdata_32_  &  pc_16_  &  (~ pc_0_) ) | ( pdata_35_  &  (~ pdata_32_)  &  (~ pc_16_)  &  (~ pc_0_) ) ;
 assign wire603 = ( (~ pdata_35_)  &  pc_2_  &  n_n1687  &  wire604 ) | ( pdata_35_  &  (~ pc_2_)  &  n_n1687  &  wire604 ) ;
 assign wire619 = ( n_n1706  &  (~ n_n1705)  &  (~ n_n1703) ) | ( n_n1704  &  (~ n_n1706)  &  n_n1705  &  n_n1703 ) ;
 assign wire618 = ( wire944 ) | ( wire520  &  wire567 ) ;
 assign wire624 = ( (~ n_n1684)  &  n_n1686  &  n_n1688  &  n_n1683 ) | ( n_n1684  &  n_n1686  &  (~ n_n1688)  &  n_n1683 ) | ( (~ n_n1684)  &  (~ n_n1686)  &  (~ n_n1688)  &  n_n1683 ) ;
 assign wire623 = ( (~ pdata_37_)  &  pdata_40_  &  pc_9_  &  pc_14_ ) | ( pdata_37_  &  (~ pdata_40_)  &  pc_9_  &  pc_14_ ) | ( pdata_37_  &  pdata_40_  &  (~ pc_9_)  &  pc_14_ ) | ( (~ pdata_37_)  &  (~ pdata_40_)  &  (~ pc_9_)  &  pc_14_ ) | ( pdata_37_  &  pdata_40_  &  pc_9_  &  (~ pc_14_) ) | ( (~ pdata_37_)  &  (~ pdata_40_)  &  pc_9_  &  (~ pc_14_) ) | ( (~ pdata_37_)  &  pdata_40_  &  (~ pc_9_)  &  (~ pc_14_) ) | ( pdata_37_  &  (~ pdata_40_)  &  (~ pc_9_)  &  (~ pc_14_) ) ;
 assign wire635 = ( (~ pd_8_)  &  pd_18_  &  pdata_50_  &  pdata_51_ ) | ( pd_8_  &  (~ pd_18_)  &  pdata_50_  &  pdata_51_ ) | ( pd_8_  &  pd_18_  &  (~ pdata_50_)  &  pdata_51_ ) | ( (~ pd_8_)  &  (~ pd_18_)  &  (~ pdata_50_)  &  pdata_51_ ) | ( pd_8_  &  pd_18_  &  pdata_50_  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  (~ pd_18_)  &  pdata_50_  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  pd_18_  &  (~ pdata_50_)  &  (~ pdata_51_) ) | ( pd_8_  &  (~ pd_18_)  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire639 = ( n_n1687  &  n_n1688  &  n_n1683 ) | ( (~ n_n1684)  &  (~ n_n1687)  &  (~ n_n1688)  &  n_n1683 ) ;
 assign wire638 = ( pdata_40_  &  pc_9_ ) | ( (~ pdata_40_)  &  (~ pc_9_) ) | ( pdata_37_  &  pc_14_ ) | ( (~ pdata_37_)  &  (~ pc_14_) ) ;
 assign wire643 = ( (~ n_n1723)  &  (~ n_n1724)  &  n_n1722 ) | ( (~ n_n1723)  &  n_n1724  &  (~ n_n1722)  &  n_n1721 ) | ( n_n1723  &  (~ n_n1724)  &  (~ n_n1722)  &  n_n1721 ) ;
 assign wire650 = ( (~ n_n1696)  &  (~ n_n1695)  &  (~ n_n1697) ) | ( n_n1699  &  (~ n_n1695)  &  (~ n_n1697) ) ;
 assign wire649 = ( pd_8_  &  pd_18_  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  (~ pd_18_)  &  pdata_50_  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  (~ pdata_50_)  &  pdata_51_ ) | ( pd_8_  &  (~ pd_18_)  &  (~ pdata_50_)  &  pdata_51_ ) | ( (~ pd_8_)  &  pd_18_  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  (~ pd_18_)  &  pdata_50_  &  (~ pdata_51_) ) | ( pd_8_  &  pd_18_  &  (~ pdata_50_)  &  (~ pdata_51_) ) | ( (~ pd_8_)  &  (~ pd_18_)  &  (~ pdata_50_)  &  (~ pdata_51_) ) ;
 assign wire663 = ( (~ n_n1702)  &  n_n1706  &  n_n1705 ) | ( n_n1702  &  n_n1706  &  (~ n_n1701) ) | ( n_n1702  &  (~ n_n1706)  &  (~ n_n1705)  &  n_n1701 ) | ( (~ n_n1702)  &  (~ n_n1706)  &  (~ n_n1705)  &  (~ n_n1701) ) ;
 assign wire667 = ( n_n1696  &  n_n1699  &  n_n1695  &  (~ n_n1697) ) | ( (~ n_n1696)  &  n_n1699  &  (~ n_n1695)  &  (~ n_n1697) ) ;
 assign wire670 = ( (~ n_n1696)  &  n_n1700  &  n_n1695  &  n_n1697 ) | ( n_n1696  &  (~ n_n1700)  &  n_n1695  &  n_n1697 ) | ( (~ n_n1696)  &  (~ n_n1700)  &  (~ n_n1695)  &  n_n1697 ) | ( (~ n_n1696)  &  n_n1700  &  (~ n_n1695)  &  (~ n_n1697) ) ;
 assign wire676 = ( n_n1690  &  (~ n_n1694)  &  n_n1693 ) | ( n_n1690  &  (~ n_n1693)  &  n_n1689 ) ;
 assign wire682 = ( n_n1715  &  (~ n_n1716)  &  n_n1713  &  n_n1717 ) | ( (~ n_n1715)  &  n_n1716  &  (~ n_n1713)  &  n_n1717 ) ;
 assign wire687 = ( n_n1699  &  n_n1695  &  (~ n_n1697) ) | ( n_n1696  &  (~ n_n1699)  &  n_n1695  &  n_n1697 ) | ( n_n1696  &  n_n1699  &  (~ n_n1695)  &  n_n1697 ) ;
 assign wire697 = ( n_n1709  &  (~ n_n1710)  &  (~ n_n1707)  &  n_n1711 ) | ( (~ n_n1709)  &  (~ n_n1710)  &  (~ n_n1707)  &  (~ n_n1711) ) ;
 assign wire706 = ( n_n1715  &  n_n1714  &  n_n1718 ) | ( n_n1715  &  (~ n_n1714)  &  n_n1713  &  (~ n_n1718) ) | ( (~ n_n1715)  &  (~ n_n1714)  &  (~ n_n1713)  &  (~ n_n1718) ) ;
 assign wire722 = ( n_n1702  &  (~ n_n1706)  &  (~ n_n1705)  &  n_n1701 ) | ( (~ n_n1702)  &  n_n1706  &  n_n1705  &  (~ n_n1701) ) ;
 assign wire724 = ( pdata_44_  &  pdata_42_  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  pc_7_  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  (~ pc_7_)  &  pc_3_ ) | ( pdata_44_  &  (~ pdata_42_)  &  (~ pc_7_)  &  pc_3_ ) | ( (~ pdata_44_)  &  pdata_42_  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  (~ pdata_42_)  &  pc_7_  &  (~ pc_3_) ) | ( pdata_44_  &  pdata_42_  &  (~ pc_7_)  &  (~ pc_3_) ) | ( (~ pdata_44_)  &  (~ pdata_42_)  &  (~ pc_7_)  &  (~ pc_3_) ) ;
 assign wire327 = ( pd_6_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire329 = ( pd_10_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire330 = ( pd_7_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire332 = ( pd_9_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire339 = ( pinreg_53_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire374 = ( pencrypt_0_  &  pinreg_45_  &  n_n1327  &  wire7712 ) ;
 assign wire376 = ( pc_7_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire377 = ( pc_11_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire378 = ( pc_8_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire382 = ( pc_10_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire383 = ( pinreg_41_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire384 = ( pinreg_33_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire404 = ( pd_5_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire414 = ( pd_9_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire415 = ( pd_6_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire416 = ( pd_8_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire418 = ( pdata_in_6_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire419 = ( pinreg_53_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire422 = ( pc_6_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire425 = ( pc_10_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire429 = ( pc_7_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire430 = ( pc_9_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire435 = ( (~ pencrypt_0_)  &  pinreg_49_  &  n_n1327  &  wire7712 ) ;
 assign wire436 = ( pinreg_41_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire451 = ( pd_7_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire452 = ( pd_11_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire453 = ( pd_8_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire454 = ( pd_10_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire455 = ( (~ pencrypt_0_)  &  pinreg_45_  &  n_n1327  &  wire7712 ) ;
 assign wire456 = ( pencrypt_0_  &  pinreg_37_  &  n_n1327  &  wire7712 ) ;
 assign wire492 = ( (~ pdata_14_)  &  n_n1327  &  wire8053 ) | ( (~ pdata_14_)  &  n_n1327  &  wire8054 ) | ( pdata_14_  &  n_n1327  &  (~ wire8053)  &  (~ wire8054) ) ;
 assign wire756 = ( (~ pdata_28_)  &  n_n1327  &  wire273 ) | ( (~ pdata_28_)  &  n_n1327  &  wire8459 ) | ( pdata_28_  &  n_n1327  &  (~ wire273)  &  (~ wire8459) ) ;
 assign wire770 = ( pc_8_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire771 = ( pc_12_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire772 = ( pc_9_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire773 = ( pc_11_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire774 = ( pinreg_33_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire775 = ( pencrypt_0_  &  pinreg_25_  &  n_n1327  &  wire7712 ) ;
 assign wire787 = ( (~ pdata_20_)  &  (~ n_n1327)  &  wire8264 ) | ( (~ pdata_20_)  &  (~ n_n1327)  &  wire8265 ) | ( pdata_20_  &  (~ n_n1327)  &  (~ wire8264)  &  (~ wire8265) ) ;
 assign wire791 = ( pd_8_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire792 = ( pd_12_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire793 = ( pd_9_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire794 = ( pd_11_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire795 = ( (~ pencrypt_0_)  &  pinreg_37_  &  n_n1327  &  wire7712 ) ;
 assign wire796 = ( pencrypt_0_  &  pinreg_29_  &  n_n1327  &  wire7712 ) ;
 assign wire798 = ( pc_18_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire799 = ( pc_22_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire800 = ( pc_19_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire801 = ( pc_21_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire802 = ( (~ pencrypt_0_)  &  pinreg_18_  &  n_n1327  &  wire7712 ) ;
 assign wire803 = ( pencrypt_0_  &  pinreg_10_  &  n_n1327  &  wire7712 ) ;
 assign wire810 = ( (~ pdata_3_)  &  n_n1327  &  wire324 ) | ( (~ pdata_3_)  &  n_n1327  &  wire7905 ) | ( pdata_3_  &  n_n1327  &  (~ wire324)  &  (~ wire7905) ) ;
 assign wire820 = ( (~ pdata_28_)  &  (~ n_n1327)  &  wire273 ) | ( (~ pdata_28_)  &  (~ n_n1327)  &  wire8459 ) | ( pdata_28_  &  (~ n_n1327)  &  (~ wire273)  &  (~ wire8459) ) ;
 assign wire824 = ( n_n1716  &  wire284  &  wire582 ) | ( n_n1716  &  wire582  &  wire831 ) ;
 assign wire825 = ( n_n1714  &  wire305  &  wire313 ) | ( n_n1714  &  wire313  &  wire833 ) ;
 assign wire827 = ( (~ n_n1715)  &  n_n1717  &  wire284  &  wire558 ) ;
 assign wire828 = ( n_n1715  &  n_n1717  &  wire528  &  wire7884 ) ;
 assign wire831 = ( pd_11_  &  pd_4_  &  pdata_52_  &  pdata_55_ ) | ( (~ pd_11_)  &  pd_4_  &  (~ pdata_52_)  &  pdata_55_ ) | ( pd_11_  &  (~ pd_4_)  &  pdata_52_  &  (~ pdata_55_) ) | ( (~ pd_11_)  &  (~ pd_4_)  &  (~ pdata_52_)  &  (~ pdata_55_) ) ;
 assign wire833 = ( pd_11_  &  pd_1_  &  pdata_51_  &  pdata_52_ ) | ( pd_11_  &  (~ pd_1_)  &  (~ pdata_51_)  &  pdata_52_ ) | ( (~ pd_11_)  &  pd_1_  &  pdata_51_  &  (~ pdata_52_) ) | ( (~ pd_11_)  &  (~ pd_1_)  &  (~ pdata_51_)  &  (~ pdata_52_) ) ;
 assign wire835 = ( (~ pd_11_)  &  pdata_52_  &  wire245  &  wire582 ) | ( pd_11_  &  (~ pdata_52_)  &  wire245  &  wire582 ) ;
 assign wire836 = ( (~ pd_19_)  &  pdata_56_  &  wire305  &  wire509 ) | ( pd_19_  &  (~ pdata_56_)  &  wire305  &  wire509 ) ;
 assign wire842 = ( (~ pdata_10_)  &  (~ n_n1327)  &  wire273 ) | ( (~ pdata_10_)  &  (~ n_n1327)  &  wire8374 ) | ( pdata_10_  &  (~ n_n1327)  &  (~ wire273)  &  (~ wire8374) ) ;
 assign wire846 = ( pd_18_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire847 = ( pd_22_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire848 = ( pd_19_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire849 = ( pd_21_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire850 = ( (~ pencrypt_0_)  &  pinreg_20_  &  n_n1327  &  wire7712 ) ;
 assign wire851 = ( pinreg_12_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire862 = ( (~ n_n1723)  &  (~ n_n1721)  &  wire586  &  wire8433 ) ;
 assign wire863 = ( (~ n_n1724)  &  n_n1720  &  wire306  &  wire271 ) ;
 assign wire866 = ( (~ n_n1723)  &  (~ n_n1721)  &  wire315  &  wire7738 ) ;
 assign wire883 = ( (~ pdata_32_)  &  pc_16_  &  wire7912  &  wire8420 ) | ( pdata_32_  &  (~ pc_16_)  &  wire7912  &  wire8420 ) ;
 assign wire889 = ( (~ pdata_34_)  &  pc_23_  &  wire591  &  wire8421 ) | ( pdata_34_  &  (~ pc_23_)  &  wire591  &  wire8421 ) ;
 assign wire892 = ( wire512  &  wire8424 ) ;
 assign wire894 = ( pdata_32_  &  pc_16_  &  wire592  &  wire513 ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  wire592  &  wire513 ) ;
 assign wire904 = ( (~ n_n1694)  &  n_n1692  &  wire309  &  wire301 ) ;
 assign wire905 = ( n_n1694  &  n_n1689  &  wire310  &  wire534 ) ;
 assign wire908 = ( wire263  &  wire301  &  wire8057 ) ;
 assign wire909 = ( (~ n_n1690)  &  (~ n_n1694)  &  wire310  &  wire308 ) ;
 assign wire934 = ( (~ pdata_32_)  &  pc_16_  &  wire512  &  wire594 ) | ( pdata_32_  &  (~ pc_16_)  &  wire512  &  wire594 ) ;
 assign wire935 = ( n_n1705  &  (~ n_n1701)  &  wire568  &  wire7912 ) ;
 assign wire937 = ( n_n1702  &  n_n1701  &  wire619 ) | ( n_n1702  &  (~ n_n1701)  &  wire618 ) ;
 assign wire944 = ( (~ pdata_32_)  &  pdata_34_  &  pc_16_  &  pc_23_ ) | ( pdata_32_  &  pdata_34_  &  (~ pc_16_)  &  pc_23_ ) | ( (~ pdata_32_)  &  (~ pdata_34_)  &  pc_16_  &  (~ pc_23_) ) | ( pdata_32_  &  (~ pdata_34_)  &  (~ pc_16_)  &  (~ pc_23_) ) ;
 assign wire954 = ( (~ pd_8_)  &  pdata_50_  &  wire289  &  wire579 ) | ( pd_8_  &  (~ pdata_50_)  &  wire289  &  wire579 ) ;
 assign wire955 = ( wire304  &  wire420  &  wire504 ) ;
 assign wire956 = ( (~ n_n1698)  &  wire962 ) | ( (~ n_n1698)  &  wire963 ) | ( (~ n_n1698)  &  wire964 ) ;
 assign wire957 = ( (~ n_n1700)  &  wire485 ) | ( (~ n_n1700)  &  n_n1698  &  wire687 ) ;
 assign wire958 = ( wire283  &  wire579  &  wire7772 ) ;
 assign wire962 = ( wire303  &  wire8389 ) ;
 assign wire963 = ( (~ pd_8_)  &  pdata_50_  &  wire262  &  wire527 ) | ( pd_8_  &  (~ pdata_50_)  &  wire262  &  wire527 ) ;
 assign wire964 = ( pdata_47_  &  pd_12_  &  wire552  &  wire304 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire552  &  wire304 ) ;
 assign wire975 = ( wire654  &  wire8378 ) ;
 assign wire976 = ( wire270  &  wire507  &  wire549 ) ;
 assign wire977 = ( n_n1712  &  n_n1711  &  wire508  &  wire7943 ) ;
 assign wire995 = ( (~ pdata_10_)  &  n_n1327  &  wire273 ) | ( (~ pdata_10_)  &  n_n1327  &  wire8374 ) | ( pdata_10_  &  n_n1327  &  (~ wire273)  &  (~ wire8374) ) ;
 assign wire1000 = ( wire305  &  wire528  &  wire558 ) ;
 assign wire1001 = ( (~ pd_16_)  &  pdata_54_  &  wire528  &  wire8367 ) | ( pd_16_  &  (~ pdata_54_)  &  wire528  &  wire8367 ) ;
 assign wire1002 = ( pd_22_  &  pdata_53_  &  wire284  &  wire274 ) | ( (~ pd_22_)  &  (~ pdata_53_)  &  wire284  &  wire274 ) ;
 assign wire1004 = ( pd_19_  &  pdata_56_  &  wire684 ) | ( (~ pd_19_)  &  (~ pdata_56_)  &  wire684 ) ;
 assign wire1005 = ( n_n1715  &  n_n1717  &  wire313  &  wire284 ) ;
 assign wire1012 = ( wire313  &  wire509  &  wire555 ) ;
 assign wire1021 = ( (~ pdata_18_)  &  (~ n_n1327)  &  wire324 ) | ( (~ pdata_18_)  &  (~ n_n1327)  &  wire8326 ) | ( pdata_18_  &  (~ n_n1327)  &  (~ wire324)  &  (~ wire8326) ) ;
 assign wire1025 = ( (~ pdata_17_)  &  n_n1327  &  wire322 ) | ( (~ pdata_17_)  &  n_n1327  &  wire8253 ) | ( pdata_17_  &  n_n1327  &  (~ wire322)  &  (~ wire8253) ) ;
 assign wire1047 = ( n_n1687  &  (~ n_n1685)  &  wire321  &  wire268 ) ;
 assign wire1049 = ( (~ pdata_36_)  &  pc_27_  &  wire8352 ) | ( pdata_36_  &  (~ pc_27_)  &  wire8352 ) | ( (~ pdata_36_)  &  pc_27_  &  wire8353 ) | ( pdata_36_  &  (~ pc_27_)  &  wire8353 ) ;
 assign wire1050 = ( pdata_35_  &  pc_2_  &  wire307  &  wire320 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  wire307  &  wire320 ) ;
 assign wire1056 = ( (~ pdata_40_)  &  pc_9_  &  wire523  &  wire8144 ) | ( pdata_40_  &  (~ pc_9_)  &  wire523  &  wire8144 ) ;
 assign wire1057 = ( pdata_35_  &  pc_2_  &  n_n1687  &  wire307 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  n_n1687  &  wire307 ) ;
 assign wire1062 = ( pd_24_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1063 = ( pd_0_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1064 = ( pd_25_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1065 = ( pd_27_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1066 = ( pinreg_3_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1067 = ( pdata_in_3_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1069 = ( pd_15_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1070 = ( pd_19_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1071 = ( pd_16_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1072 = ( pd_18_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1073 = ( (~ pencrypt_0_)  &  pinreg_44_  &  n_n1327  &  wire7712 ) ;
 assign wire1074 = ( pencrypt_0_  &  pinreg_36_  &  n_n1327  &  wire7712 ) ;
 assign wire1076 = ( pc_25_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1077 = ( pc_1_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1078 = ( pc_26_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1079 = ( pc_0_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1080 = ( (~ pencrypt_0_)  &  pinreg_27_  &  n_n1327  &  wire7712 ) ;
 assign wire1081 = ( pencrypt_0_  &  pinreg_48_  &  n_n1327  &  wire7712 ) ;
 assign wire1083 = ( pc_16_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1084 = ( pc_20_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1085 = ( pc_17_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1086 = ( pc_19_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1087 = ( (~ pencrypt_0_)  &  pinreg_34_  &  n_n1327  &  wire7712 ) ;
 assign wire1088 = ( pencrypt_0_  &  pinreg_26_  &  n_n1327  &  wire7712 ) ;
 assign wire1093 = ( (~ pdata_18_)  &  n_n1327  &  wire324 ) | ( (~ pdata_18_)  &  n_n1327  &  wire8326 ) | ( pdata_18_  &  n_n1327  &  (~ wire324)  &  (~ wire8326) ) ;
 assign wire1098 = ( pd_1_  &  pdata_51_  &  wire313  &  wire540 ) | ( (~ pd_1_)  &  (~ pdata_51_)  &  wire313  &  wire540 ) ;
 assign wire1099 = ( wire245  &  wire305  &  wire517 ) ;
 assign wire1101 = ( n_n1718  &  wire8320 ) | ( (~ n_n1714)  &  n_n1718  &  wire682 ) ;
 assign wire1102 = ( (~ n_n1715)  &  n_n1717  &  wire505  &  wire558 ) ;
 assign wire1111 = ( wire517  &  wire509  &  wire555 ) ;
 assign wire1112 = ( wire305  &  wire313  &  wire284 ) ;
 assign wire1113 = ( (~ n_n1715)  &  n_n1717  &  wire505  &  wire7884 ) ;
 assign wire1114 = ( n_n1715  &  n_n1717  &  wire528  &  wire558 ) ;
 assign wire1126 = ( pd_23_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1127 = ( pd_27_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1128 = ( pd_24_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1129 = ( pd_26_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1130 = ( (~ pencrypt_0_)  &  pinreg_11_  &  n_n1327  &  wire7712 ) ;
 assign wire1131 = ( pinreg_3_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1133 = ( pd_16_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1134 = ( pd_20_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1135 = ( pd_17_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1136 = ( pd_19_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1137 = ( (~ pencrypt_0_)  &  pinreg_36_  &  n_n1327  &  wire7712 ) ;
 assign wire1138 = ( pencrypt_0_  &  pinreg_28_  &  n_n1327  &  wire7712 ) ;
 assign wire1140 = ( pc_15_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1141 = ( pc_19_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1142 = ( pc_16_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1143 = ( pc_18_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1144 = ( pinreg_42_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1145 = ( pencrypt_0_  &  pinreg_34_  &  n_n1327  &  wire7712 ) ;
 assign wire1152 = ( (~ n_n1690)  &  n_n1693  &  wire286  &  wire308 ) ;
 assign wire1156 = ( (~ n_n1691)  &  n_n1692  &  wire309  &  wire285 ) ;
 assign wire1180 = ( pcount_3_  &  pcount_new_0_ ) | ( pcount_3_  &  wire1182 ) | ( pcount_3_  &  wire1519 ) ;
 assign wire1181 = ( (~ preset_0_)  &  (~ pload_key_0_)  &  wire392 ) | ( (~ preset_0_)  &  (~ n_n1327)  &  wire392 ) ;
 assign wire1182 = ( (~ pcount_2_)  &  (~ preset_0_)  &  (~ pload_key_0_) ) | ( (~ pcount_2_)  &  (~ preset_0_)  &  (~ n_n1327) ) ;
 assign wire1184 = ( pd_13_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1185 = ( pd_17_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1186 = ( pd_14_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1187 = ( pd_16_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1188 = ( pdata_in_5_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1189 = ( pinreg_52_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1191 = ( pc_23_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1192 = ( pc_27_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1193 = ( pc_24_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1194 = ( pc_26_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1195 = ( pinreg_43_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1196 = ( pencrypt_0_  &  pinreg_35_  &  n_n1327  &  wire7712 ) ;
 assign wire1198 = ( pc_14_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1199 = ( pc_18_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1200 = ( pc_15_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1201 = ( pc_17_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1202 = ( pinreg_50_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1203 = ( pinreg_42_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1211 = ( (~ pdata_20_)  &  n_n1327  &  wire8264 ) | ( (~ pdata_20_)  &  n_n1327  &  wire8265 ) | ( pdata_20_  &  n_n1327  &  (~ wire8264)  &  (~ wire8265) ) ;
 assign wire1216 = ( (~ n_n1726)  &  (~ n_n1729)  &  wire531  &  wire7856 ) ;
 assign wire1220 = ( wire265  &  wire295  &  wire7844 ) ;
 assign wire1221 = ( n_n1725  &  n_n1729  &  wire265  &  wire7853 ) ;
 assign wire1222 = ( (~ n_n1726)  &  n_n1729  &  wire531  &  wire506 ) ;
 assign wire1229 = ( (~ pdata_23_)  &  n_n1327  &  wire323 ) | ( (~ pdata_23_)  &  n_n1327  &  wire8210 ) | ( pdata_23_  &  n_n1327  &  (~ wire323)  &  (~ wire8210) ) ;
 assign wire1238 = ( (~ pdata_17_)  &  (~ n_n1327)  &  wire322 ) | ( (~ pdata_17_)  &  (~ n_n1327)  &  wire8253 ) | ( pdata_17_  &  (~ n_n1327)  &  (~ wire322)  &  (~ wire8253) ) ;
 assign wire1242 = ( n_n1686  &  (~ n_n1685)  &  wire523  &  wire320 ) ;
 assign wire1243 = ( (~ n_n1686)  &  (~ n_n1685)  &  wire533  &  wire604 ) ;
 assign wire1244 = ( (~ pdata_36_)  &  pc_27_  &  wire1249 ) | ( pdata_36_  &  (~ pc_27_)  &  wire1249 ) | ( (~ pdata_36_)  &  pc_27_  &  wire1250 ) | ( pdata_36_  &  (~ pc_27_)  &  wire1250 ) ;
 assign wire1245 = ( n_n1687  &  wire1253 ) | ( n_n1687  &  wire1254 ) | ( n_n1687  &  wire8247 ) ;
 assign wire1246 = ( pdata_35_  &  pc_2_  &  wire321  &  wire320 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  wire321  &  wire320 ) ;
 assign wire1249 = ( (~ pdata_35_)  &  pc_2_  &  (~ n_n1683)  &  wire320 ) | ( pdata_35_  &  (~ pc_2_)  &  (~ n_n1683)  &  wire320 ) ;
 assign wire1250 = ( wire307  &  wire533 ) ;
 assign wire1253 = ( pdata_36_  &  pc_27_  &  wire307  &  wire268 ) | ( (~ pdata_36_)  &  (~ pc_27_)  &  wire307  &  wire268 ) ;
 assign wire1254 = ( (~ n_n1684)  &  n_n1686  &  (~ n_n1685)  &  wire523 ) ;
 assign wire1257 = ( pd_25_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1258 = ( pd_1_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1259 = ( pd_26_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1260 = ( pd_0_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1261 = ( pdata_in_3_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1262 = ( pencrypt_0_  &  pinreg_54_  &  n_n1327  &  wire7712 ) ;
 assign wire1264 = ( pd_14_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1265 = ( pd_18_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1266 = ( pd_15_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1267 = ( pd_17_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1268 = ( pinreg_52_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1269 = ( pencrypt_0_  &  pinreg_44_  &  n_n1327  &  wire7712 ) ;
 assign wire1271 = ( pc_24_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1272 = ( pc_0_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1273 = ( pc_25_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1274 = ( pc_27_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1275 = ( (~ pencrypt_0_)  &  pinreg_35_  &  n_n1327  &  wire7712 ) ;
 assign wire1276 = ( pencrypt_0_  &  pinreg_27_  &  n_n1327  &  wire7712 ) ;
 assign wire1278 = ( pc_13_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1279 = ( pc_17_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1280 = ( pc_14_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1281 = ( pc_16_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1282 = ( (~ pencrypt_0_)  &  pdata_in_1_  &  n_n1327  &  wire7712 ) ;
 assign wire1283 = ( pinreg_50_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1291 = ( wire246  &  (~ wire271)  &  wire585 ) ;
 assign wire1301 = ( n_n1719  &  n_n1721  &  wire7731 ) | ( n_n1719  &  n_n1721  &  wire8215 ) ;
 assign wire1319 = ( (~ pdata_23_)  &  (~ n_n1327)  &  wire323 ) | ( (~ pdata_23_)  &  (~ n_n1327)  &  wire8210 ) | ( pdata_23_  &  (~ n_n1327)  &  (~ wire323)  &  (~ wire8210) ) ;
 assign wire1324 = ( wire270  &  wire525  &  wire537 ) ;
 assign wire1325 = ( pdata_44_  &  pc_7_  &  wire426 ) | ( (~ pdata_44_)  &  (~ pc_7_)  &  wire426 ) | ( pdata_44_  &  pc_7_  &  wire1331 ) | ( (~ pdata_44_)  &  (~ pc_7_)  &  wire1331 ) ;
 assign wire1326 = ( (~ pdata_43_)  &  pc_25_  &  wire507  &  wire302 ) | ( pdata_43_  &  (~ pc_25_)  &  wire507  &  wire302 ) ;
 assign wire1327 = ( (~ pdata_44_)  &  pc_7_  &  wire526  &  wire7948 ) | ( pdata_44_  &  (~ pc_7_)  &  wire526  &  wire7948 ) ;
 assign wire1331 = ( wire302  &  wire8204 ) ;
 assign wire1341 = ( pd_20_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1342 = ( pd_24_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1343 = ( pd_21_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1344 = ( pd_23_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1345 = ( pinreg_4_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1346 = ( pdata_in_4_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1348 = ( pd_11_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1349 = ( pd_15_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1350 = ( pd_12_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1351 = ( pd_14_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1352 = ( (~ pencrypt_0_)  &  pinreg_13_  &  n_n1327  &  wire7712 ) ;
 assign wire1353 = ( pinreg_5_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1355 = ( pc_21_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1356 = ( pc_25_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1357 = ( pc_22_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1358 = ( pc_24_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1359 = ( (~ pencrypt_0_)  &  pdata_in_2_  &  n_n1327  &  wire7712 ) ;
 assign wire1360 = ( pinreg_51_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1362 = ( pc_12_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1363 = ( pc_16_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1364 = ( pc_13_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1365 = ( pc_15_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1366 = ( pinreg_1_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1367 = ( pencrypt_0_  &  pdata_in_1_  &  n_n1327  &  wire7712 ) ;
 assign wire1380 = ( (~ pdata_36_)  &  pc_27_  &  wire1390 ) | ( pdata_36_  &  (~ pc_27_)  &  wire1390 ) | ( (~ pdata_36_)  &  pc_27_  &  wire8175 ) | ( pdata_36_  &  (~ pc_27_)  &  wire8175 ) ;
 assign wire1383 = ( (~ n_n1688)  &  (~ n_n1683)  &  wire598 ) | ( n_n1687  &  n_n1688  &  n_n1683  &  wire598 ) ;
 assign wire1384 = ( (~ pdata_40_)  &  pc_9_  &  wire604  &  wire8144 ) | ( pdata_40_  &  (~ pc_9_)  &  wire604  &  wire8144 ) ;
 assign wire1385 = ( pdata_35_  &  pc_2_  &  (~ n_n1688)  &  wire320 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  (~ n_n1688)  &  wire320 ) ;
 assign wire1386 = ( pdata_35_  &  pc_2_  &  wire307  &  wire569 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  wire307  &  wire569 ) ;
 assign wire1389 = ( (~ pdata_35_)  &  pc_2_  &  wire604  &  wire623 ) | ( pdata_35_  &  (~ pc_2_)  &  wire604  &  wire623 ) ;
 assign wire1390 = ( pdata_40_  &  pc_9_  &  wire624 ) | ( (~ pdata_40_)  &  (~ pc_9_)  &  wire624 ) ;
 assign wire1391 = ( (~ n_n1684)  &  (~ n_n1686)  &  n_n1687  &  wire523 ) ;
 assign wire1392 = ( (~ pdata_40_)  &  pc_9_  &  wire307  &  wire8144 ) | ( pdata_40_  &  (~ pc_9_)  &  wire307  &  wire8144 ) ;
 assign wire1397 = ( (~ n_n1684)  &  (~ n_n1686)  &  wire523  &  wire8170 ) ;
 assign wire1399 = ( n_n1686  &  n_n1685  &  wire321  &  wire569 ) ;
 assign wire1411 = ( (~ pdata_36_)  &  pc_27_  &  wire8162 ) | ( pdata_36_  &  (~ pc_27_)  &  wire8162 ) | ( (~ pdata_36_)  &  pc_27_  &  wire8163 ) | ( pdata_36_  &  (~ pc_27_)  &  wire8163 ) ;
 assign wire1412 = ( (~ pdata_35_)  &  pc_2_  &  wire307  &  wire320 ) | ( pdata_35_  &  (~ pc_2_)  &  wire307  &  wire320 ) ;
 assign wire1413 = ( n_n1687  &  (~ n_n1685)  &  wire321  &  wire8144 ) ;
 assign wire1418 = ( pdata_35_  &  pc_2_  &  wire307  &  wire638 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  wire307  &  wire638 ) ;
 assign wire1420 = ( (~ pdata_40_)  &  pc_9_  &  wire604  &  wire8144 ) | ( pdata_40_  &  (~ pc_9_)  &  wire604  &  wire8144 ) ;
 assign wire1421 = ( (~ pdata_35_)  &  pc_2_  &  wire533  &  wire604 ) | ( pdata_35_  &  (~ pc_2_)  &  wire533  &  wire604 ) ;
 assign wire1425 = ( (~ n_n1684)  &  (~ n_n1686)  &  wire523  &  wire8155 ) ;
 assign wire1426 = ( (~ n_n1686)  &  (~ n_n1685)  &  wire604  &  wire569 ) ;
 assign wire1427 = ( n_n1686  &  (~ n_n1685)  &  wire307  &  wire569 ) ;
 assign wire1428 = ( n_n1686  &  (~ n_n1685)  &  wire321  &  wire320 ) ;
 assign wire1429 = ( (~ n_n1686)  &  n_n1685  &  wire523  &  wire320 ) ;
 assign wire1430 = ( n_n1686  &  (~ n_n1685)  &  wire321  &  wire569 ) ;
 assign wire1434 = ( n_n1686  &  n_n1685  &  wire523  &  wire320 ) ;
 assign wire1435 = ( pdata_36_  &  pc_27_  &  wire1437 ) | ( (~ pdata_36_)  &  (~ pc_27_)  &  wire1437 ) | ( pdata_36_  &  pc_27_  &  wire1438 ) | ( (~ pdata_36_)  &  (~ pc_27_)  &  wire1438 ) ;
 assign wire1436 = ( n_n1687  &  (~ n_n1685)  &  wire307  &  wire8144 ) ;
 assign wire1437 = ( n_n1684  &  n_n1686  &  n_n1687  &  wire604 ) ;
 assign wire1438 = ( pdata_35_  &  pc_2_  &  wire307  &  wire533 ) | ( (~ pdata_35_)  &  (~ pc_2_)  &  wire307  &  wire533 ) ;
 assign wire1439 = ( n_n1687  &  n_n1685  &  wire321  &  wire598 ) ;
 assign wire1440 = ( (~ n_n1685)  &  wire1441 ) | ( (~ n_n1685)  &  wire1442 ) | ( (~ n_n1685)  &  wire1443 ) ;
 assign wire1441 = ( (~ n_n1684)  &  (~ n_n1686)  &  (~ n_n1687)  &  wire523 ) ;
 assign wire1442 = ( (~ pdata_35_)  &  pc_2_  &  wire533  &  wire604 ) | ( pdata_35_  &  (~ pc_2_)  &  wire533  &  wire604 ) ;
 assign wire1443 = ( (~ pdata_40_)  &  pc_9_  &  wire523  &  wire8144 ) | ( pdata_40_  &  (~ pc_9_)  &  wire523  &  wire8144 ) ;
 assign wire1444 = ( n_n1686  &  n_n1685  &  wire307  &  wire569 ) ;
 assign wire1445 = ( (~ n_n1684)  &  n_n1686  &  wire523  &  wire8143 ) ;
 assign wire1446 = ( (~ n_n1686)  &  (~ n_n1685)  &  wire320  &  wire604 ) ;
 assign wire1447 = ( n_n1687  &  n_n1685  &  wire321  &  wire8144 ) ;
 assign wire1474 = ( pd_2_  &  pdata_49_  &  wire1483 ) | ( (~ pd_2_)  &  (~ pdata_49_)  &  wire1483 ) | ( pd_2_  &  pdata_49_  &  wire1484 ) | ( (~ pd_2_)  &  (~ pdata_49_)  &  wire1484 ) ;
 assign wire1475 = ( n_n1698  &  wire8134 ) | ( n_n1700  &  n_n1698  &  wire650 ) ;
 assign wire1476 = ( wire552  &  wire579  &  wire7772 ) ;
 assign wire1477 = ( pdata_47_  &  pd_12_  &  wire289  &  wire303 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire289  &  wire303 ) ;
 assign wire1478 = ( (~ pdata_47_)  &  pd_12_  &  wire289  &  wire283 ) | ( pdata_47_  &  (~ pd_12_)  &  wire289  &  wire283 ) ;
 assign wire1483 = ( pd_8_  &  pdata_50_  &  (~ wire262)  &  wire527 ) | ( (~ pd_8_)  &  (~ pdata_50_)  &  (~ wire262)  &  wire527 ) ;
 assign wire1484 = ( pdata_47_  &  pd_12_  &  wire552  &  wire261 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire552  &  wire261 ) ;
 assign wire1494 = ( n_n1710  &  n_n1708  &  (~ wire247)  &  wire302 ) ;
 assign wire1495 = ( (~ n_n1712)  &  n_n1711  &  wire508  &  wire7943 ) ;
 assign wire1496 = ( pdata_43_  &  pc_25_  &  wire431 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire431 ) | ( pdata_43_  &  pc_25_  &  wire1501 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire1501 ) ;
 assign wire1498 = ( pdata_43_  &  pc_25_  &  wire525  &  wire267 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire525  &  wire267 ) ;
 assign wire1501 = ( (~ pdata_42_)  &  pc_3_  &  (~ n_n1712)  &  wire503 ) | ( pdata_42_  &  (~ pc_3_)  &  (~ n_n1712)  &  wire503 ) ;
 assign wire1503 = ( pdata_41_  &  pc_11_  &  wire536  &  wire8125 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  wire536  &  wire8125 ) ;
 assign wire1505 = ( (~ pdata_44_)  &  pc_7_  &  n_n1711  &  wire7943 ) | ( pdata_44_  &  (~ pc_7_)  &  n_n1711  &  wire7943 ) ;
 assign wire1508 = ( wire549  &  wire536  &  wire515 ) ;
 assign wire1509 = ( (~ n_n1712)  &  n_n1708  &  wire507  &  wire503 ) | ( n_n1712  &  (~ n_n1708)  &  wire507  &  wire503 ) ;
 assign wire1510 = ( (~ n_n1710)  &  n_n1708  &  wire302  &  wire536 ) ;
 assign wire1519 = ( (~ pcount_1_)  &  (~ preset_0_)  &  (~ pload_key_0_) ) | ( (~ pcount_1_)  &  (~ preset_0_)  &  (~ n_n1327) ) ;
 assign wire1521 = ( pd_19_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1522 = ( pd_23_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1523 = ( pd_20_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1524 = ( pd_22_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1525 = ( pinreg_12_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1526 = ( pinreg_4_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1528 = ( pd_12_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1529 = ( pd_16_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1530 = ( pd_13_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1531 = ( pd_15_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1532 = ( pinreg_5_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1533 = ( pdata_in_5_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1535 = ( pc_22_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1536 = ( pc_26_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1537 = ( pc_23_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1538 = ( pc_25_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1539 = ( pinreg_51_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1540 = ( pinreg_43_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1542 = ( pc_11_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1543 = ( pc_15_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1544 = ( pc_12_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1545 = ( pc_14_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1546 = ( pinreg_9_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1547 = ( pinreg_1_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1556 = ( (~ n_n1690)  &  (~ n_n1694)  &  wire308  &  wire8084 ) ;
 assign wire1559 = ( n_n1691  &  wire433 ) | ( n_n1691  &  (~ n_n1692)  &  wire676 ) ;
 assign wire1560 = ( (~ n_n1694)  &  n_n1689  &  wire310  &  wire301 ) ;
 assign wire1561 = ( n_n1690  &  (~ n_n1693)  &  wire286  &  wire8088 ) ;
 assign wire1562 = ( (~ n_n1691)  &  n_n1692  &  (~ n_n1689)  &  wire285 ) ;
 assign wire1574 = ( (~ n_n1694)  &  (~ n_n1689)  &  wire301  &  wire524 ) ;
 assign wire1576 = ( (~ n_n1690)  &  n_n1694  &  wire310  &  wire308 ) ;
 assign wire1597 = ( pdata_44_  &  pc_6_  &  wire286  &  wire8067 ) | ( (~ pdata_44_)  &  (~ pc_6_)  &  wire286  &  wire8067 ) ;
 assign wire1598 = ( (~ n_n1691)  &  n_n1689  &  wire285  &  wire524 ) ;
 assign wire1599 = ( pdata_43_  &  pc_15_  &  wire310  &  wire308 ) | ( (~ pdata_43_)  &  (~ pc_15_)  &  wire310  &  wire308 ) ;
 assign wire1600 = ( (~ pdata_43_)  &  pc_15_  &  wire309  &  wire301 ) | ( pdata_43_  &  (~ pc_15_)  &  wire309  &  wire301 ) ;
 assign wire1601 = ( (~ pdata_44_)  &  pc_6_  &  wire380 ) | ( pdata_44_  &  (~ pc_6_)  &  wire380 ) | ( (~ pdata_44_)  &  pc_6_  &  wire1607 ) | ( pdata_44_  &  (~ pc_6_)  &  wire1607 ) ;
 assign wire1602 = ( (~ pdata_46_)  &  pc_19_  &  wire309  &  wire285 ) | ( pdata_46_  &  (~ pc_19_)  &  wire309  &  wire285 ) ;
 assign wire1607 = ( pdata_47_  &  pc_12_  &  wire263  &  wire308 ) | ( (~ pdata_47_)  &  (~ pc_12_)  &  wire263  &  wire308 ) ;
 assign wire1617 = ( n_n1690  &  n_n1691  &  wire309  &  wire286 ) ;
 assign wire1618 = ( n_n1694  &  (~ n_n1689)  &  wire310  &  wire534 ) ;
 assign wire1619 = ( pdata_43_  &  pc_15_  &  wire1620 ) | ( (~ pdata_43_)  &  (~ pc_15_)  &  wire1620 ) | ( pdata_43_  &  pc_15_  &  wire1621 ) | ( (~ pdata_43_)  &  (~ pc_15_)  &  wire1621 ) ;
 assign wire1620 = ( (~ pdata_48_)  &  pc_1_  &  wire524  &  wire8063 ) | ( pdata_48_  &  (~ pc_1_)  &  wire524  &  wire8063 ) ;
 assign wire1621 = ( (~ pdata_45_)  &  pc_26_  &  wire301  &  wire8057 ) | ( pdata_45_  &  (~ pc_26_)  &  wire301  &  wire8057 ) ;
 assign wire1625 = ( wire286  &  wire308  &  wire8060 ) ;
 assign wire1626 = ( (~ n_n1690)  &  (~ n_n1694)  &  wire308  &  wire524 ) ;
 assign wire1630 = ( wire285  &  wire308  &  wire8055 ) ;
 assign wire1631 = ( (~ pdata_48_)  &  pc_1_  &  wire1633 ) | ( pdata_48_  &  (~ pc_1_)  &  wire1633 ) | ( (~ pdata_48_)  &  pc_1_  &  wire1634 ) | ( pdata_48_  &  (~ pc_1_)  &  wire1634 ) ;
 assign wire1632 = ( wire286  &  wire301  &  wire8057 ) ;
 assign wire1633 = ( pdata_44_  &  pc_6_  &  wire286  &  wire534 ) | ( (~ pdata_44_)  &  (~ pc_6_)  &  wire286  &  wire534 ) ;
 assign wire1634 = ( pdata_46_  &  pc_19_  &  wire285  &  wire310 ) | ( (~ pdata_46_)  &  (~ pc_19_)  &  wire285  &  wire310 ) ;
 assign wire1647 = ( (~ pdata_14_)  &  (~ n_n1327)  &  wire8053 ) | ( (~ pdata_14_)  &  (~ n_n1327)  &  wire8054 ) | ( pdata_14_  &  (~ n_n1327)  &  (~ wire8053)  &  (~ wire8054) ) ;
 assign wire1651 = ( (~ n_n1725)  &  (~ n_n1730)  &  wire543  &  wire295 ) ;
 assign wire1652 = ( n_n1726  &  n_n1729  &  wire506  &  wire562 ) ;
 assign wire1653 = ( wire543  &  wire588  &  wire7857 ) ;
 assign wire1654 = ( (~ n_n1726)  &  n_n1725  &  n_n1729  &  wire7846 ) ;
 assign wire1655 = ( pd_7_  &  pdata_62_  &  wire506  &  wire7850 ) | ( (~ pd_7_)  &  (~ pdata_62_)  &  wire506  &  wire7850 ) ;
 assign wire1656 = ( n_n1726  &  (~ n_n1729)  &  wire297  &  wire7856 ) ;
 assign wire1657 = ( pd_21_  &  pdata_61_  &  wire297  &  wire7996 ) | ( (~ pd_21_)  &  (~ pdata_61_)  &  wire297  &  wire7996 ) ;
 assign wire1659 = ( pdata_32_  &  pd_3_  &  wire280 ) | ( (~ pdata_32_)  &  (~ pd_3_)  &  wire280 ) | ( pdata_32_  &  pd_3_  &  wire1756 ) | ( (~ pdata_32_)  &  (~ pd_3_)  &  wire1756 ) ;
 assign wire1660 = ( (~ n_n1726)  &  (~ n_n1730)  &  n_n1727  &  wire511 ) ;
 assign wire1666 = ( pd_22_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1667 = ( pd_26_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1668 = ( pd_23_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1669 = ( pd_25_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1670 = ( (~ pencrypt_0_)  &  pinreg_19_  &  n_n1327  &  wire7712 ) ;
 assign wire1671 = ( pencrypt_0_  &  pinreg_11_  &  n_n1327  &  wire7712 ) ;
 assign wire1673 = ( pd_9_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1674 = ( pd_13_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1675 = ( pd_10_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1676 = ( pd_12_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1677 = ( (~ pencrypt_0_)  &  pinreg_29_  &  n_n1327  &  wire7712 ) ;
 assign wire1678 = ( pencrypt_0_  &  pinreg_21_  &  n_n1327  &  wire7712 ) ;
 assign wire1680 = ( pc_19_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1681 = ( pc_23_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1682 = ( pc_20_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1683 = ( pc_22_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1684 = ( (~ pencrypt_0_)  &  pinreg_10_  &  n_n1327  &  wire7712 ) ;
 assign wire1685 = ( pinreg_2_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1687 = ( pc_10_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1688 = ( pc_14_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1689 = ( pc_11_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1690 = ( pc_13_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1691 = ( (~ pencrypt_0_)  &  pinreg_17_  &  n_n1327  &  wire7712 ) ;
 assign wire1692 = ( pinreg_9_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1695 = ( (~ pcount_0_)  &  poutreg_61_ ) ;
 assign wire1698 = ( n_n1704  &  wire1704 ) | ( n_n1704  &  wire1705 ) | ( n_n1704  &  wire1706 ) ;
 assign wire1699 = ( (~ n_n1704)  &  wire1707 ) | ( (~ n_n1704)  &  wire1708 ) | ( (~ n_n1704)  &  wire1709 ) ;
 assign wire1704 = ( pdata_32_  &  pc_16_  &  wire264  &  wire519 ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  wire264  &  wire519 ) ;
 assign wire1705 = ( pdata_34_  &  pc_23_  &  wire592  &  wire319 ) | ( (~ pdata_34_)  &  (~ pc_23_)  &  wire592  &  wire319 ) ;
 assign wire1706 = ( (~ pdata_32_)  &  pc_16_  &  n_n1703  &  wire7912 ) | ( pdata_32_  &  (~ pc_16_)  &  n_n1703  &  wire7912 ) ;
 assign wire1707 = ( (~ pdata_34_)  &  pc_23_  &  wire496  &  wire319 ) | ( pdata_34_  &  (~ pc_23_)  &  wire496  &  wire319 ) ;
 assign wire1708 = ( (~ n_n1706)  &  n_n1701  &  n_n1703  &  wire591 ) | ( n_n1706  &  n_n1701  &  (~ n_n1703)  &  wire591 ) | ( (~ n_n1706)  &  (~ n_n1701)  &  (~ n_n1703)  &  wire591 ) ;
 assign wire1709 = ( (~ n_n1702)  &  n_n1705  &  n_n1701  &  wire519 ) | ( n_n1702  &  n_n1705  &  (~ n_n1701)  &  wire519 ) | ( (~ n_n1702)  &  (~ n_n1705)  &  (~ n_n1701)  &  wire519 ) ;
 assign wire1714 = ( (~ wire496)  &  wire513  &  wire595 ) ;
 assign wire1716 = ( wire512  &  wire594  &  wire520 ) ;
 assign wire1723 = ( (~ pdata_4_)  &  n_n1327  &  wire7871 ) | ( (~ pdata_4_)  &  n_n1327  &  wire7872 ) | ( pdata_4_  &  n_n1327  &  (~ wire7871)  &  (~ wire7872) ) ;
 assign wire1741 = ( n_n1726  &  (~ n_n1730)  &  wire297  &  wire543 ) ;
 assign wire1742 = ( (~ pd_21_)  &  pdata_61_  &  wire424 ) | ( pd_21_  &  (~ pdata_61_)  &  wire424 ) | ( (~ pd_21_)  &  pdata_61_  &  wire439 ) | ( pd_21_  &  (~ pdata_61_)  &  wire439 ) ;
 assign wire1744 = ( (~ pdata_59_)  &  pd_17_  &  wire295  &  wire511 ) | ( pdata_59_  &  (~ pd_17_)  &  wire295  &  wire511 ) ;
 assign wire1745 = ( wire297  &  wire543  &  wire7857 ) ;
 assign wire1746 = ( (~ n_n1725)  &  (~ n_n1729)  &  wire295  &  wire7856 ) ;
 assign wire1747 = ( (~ n_n1726)  &  n_n1727  &  n_n1729  &  wire7846 ) ;
 assign wire1753 = ( (~ n_n1726)  &  (~ n_n1727)  &  (~ n_n1729)  &  wire7856 ) ;
 assign wire1754 = ( wire295  &  wire511 ) ;
 assign wire1756 = ( (~ pdata_59_)  &  pd_17_  &  n_n1729  &  wire295 ) | ( pdata_59_  &  (~ pd_17_)  &  n_n1729  &  wire295 ) ;
 assign wire1758 = ( n_n1726  &  n_n1730  &  wire543  &  wire562 ) ;
 assign wire1759 = ( n_n1726  &  n_n1729  &  wire297  &  wire506 ) ;
 assign wire1760 = ( wire531  &  wire543  &  wire7857 ) ;
 assign wire1761 = ( wire506  &  wire562  &  wire7850 ) ;
 assign wire1766 = ( pd_21_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1767 = ( pd_25_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1768 = ( pd_22_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1769 = ( pd_24_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1770 = ( pdata_in_4_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1771 = ( pencrypt_0_  &  pinreg_19_  &  n_n1327  &  wire7712 ) ;
 assign wire1773 = ( pd_10_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1774 = ( pd_14_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1775 = ( pd_11_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1776 = ( pd_13_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1777 = ( (~ pencrypt_0_)  &  pinreg_21_  &  n_n1327  &  wire7712 ) ;
 assign wire1778 = ( pencrypt_0_  &  pinreg_13_  &  n_n1327  &  wire7712 ) ;
 assign wire1780 = ( pc_20_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1781 = ( pc_24_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1782 = ( pc_21_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1783 = ( pc_23_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1784 = ( pinreg_2_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1785 = ( pencrypt_0_  &  pdata_in_2_  &  n_n1327  &  wire7712 ) ;
 assign wire1787 = ( pc_9_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1788 = ( pc_13_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1789 = ( pc_10_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1790 = ( pc_12_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1791 = ( (~ pencrypt_0_)  &  pinreg_25_  &  n_n1327  &  wire7712 ) ;
 assign wire1792 = ( pencrypt_0_  &  pinreg_17_  &  n_n1327  &  wire7712 ) ;
 assign wire1805 = ( wire270  &  wire526  &  wire536 ) ;
 assign wire1806 = ( wire247  &  wire328  &  wire503 ) ;
 assign wire1807 = ( (~ n_n1710)  &  (~ n_n1708)  &  wire302  &  wire536 ) ;
 assign wire1808 = ( pdata_41_  &  pc_11_  &  wire1813 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  wire1813 ) | ( pdata_41_  &  pc_11_  &  wire1814 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  wire1814 ) ;
 assign wire1809 = ( n_n1710  &  wire1815 ) | ( n_n1710  &  wire1816 ) | ( n_n1710  &  wire1817 ) ;
 assign wire1810 = ( n_n1707  &  n_n1711  &  wire7943  &  wire7962 ) ;
 assign wire1813 = ( (~ pdata_43_)  &  pc_25_  &  wire507  &  wire302 ) | ( pdata_43_  &  (~ pc_25_)  &  wire507  &  wire302 ) ;
 assign wire1814 = ( pdata_43_  &  pc_25_  &  wire525  &  wire526 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire525  &  wire526 ) ;
 assign wire1815 = ( wire525  &  wire7960 ) ;
 assign wire1816 = ( (~ pdata_43_)  &  pc_25_  &  (~ n_n1707)  &  wire302 ) | ( pdata_43_  &  (~ pc_25_)  &  (~ n_n1707)  &  wire302 ) ;
 assign wire1817 = ( pdata_43_  &  pc_25_  &  wire525  &  wire302 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire525  &  wire302 ) ;
 assign wire1818 = ( n_n1710  &  (~ n_n1708)  &  wire525  &  wire549 ) ;
 assign wire1819 = ( (~ n_n1712)  &  n_n1711  &  wire525  &  wire7943 ) ;
 assign wire1829 = ( n_n1712  &  n_n1708  &  wire525  &  wire503 ) ;
 assign wire1830 = ( wire526  &  wire7948  &  wire7949 ) ;
 assign wire1834 = ( (~ n_n1710)  &  n_n1708  &  wire525  &  wire302 ) ;
 assign wire1835 = ( n_n1712  &  n_n1711  &  wire536  &  wire7943 ) ;
 assign wire1836 = ( (~ pdata_43_)  &  pc_25_  &  wire1837 ) | ( pdata_43_  &  (~ pc_25_)  &  wire1837 ) | ( (~ pdata_43_)  &  pc_25_  &  wire1838 ) | ( pdata_43_  &  (~ pc_25_)  &  wire1838 ) ;
 assign wire1837 = ( (~ pdata_41_)  &  pc_11_  &  wire507  &  wire526 ) | ( pdata_41_  &  (~ pc_11_)  &  wire507  &  wire526 ) ;
 assign wire1838 = ( pdata_41_  &  pc_11_  &  wire537  &  wire536 ) | ( (~ pdata_41_)  &  (~ pc_11_)  &  wire537  &  wire536 ) ;
 assign wire1839 = ( (~ n_n1712)  &  n_n1708  &  wire508  &  wire503 ) ;
 assign wire1841 = ( pdata_43_  &  pc_25_  &  wire526  &  wire724 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire526  &  wire724 ) ;
 assign wire1842 = ( pdata_43_  &  pc_25_  &  wire525  &  wire302 ) | ( (~ pdata_43_)  &  (~ pc_25_)  &  wire525  &  wire302 ) ;
 assign wire1857 = ( pd_26_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1858 = ( pd_2_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1859 = ( pd_27_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1860 = ( pd_1_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1861 = ( (~ pencrypt_0_)  &  pinreg_54_  &  n_n1327  &  wire7712 ) ;
 assign wire1862 = ( pencrypt_0_  &  pinreg_46_  &  n_n1327  &  wire7712 ) ;
 assign wire1864 = ( pc_27_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1865 = ( pc_3_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1866 = ( pc_0_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1867 = ( pc_2_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1868 = ( pinreg_40_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire1869 = ( pinreg_32_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1882 = ( pc_26_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1883 = ( pc_2_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1884 = ( pc_27_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1885 = ( pc_1_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire1886 = ( (~ pencrypt_0_)  &  pinreg_48_  &  n_n1327  &  wire7712 ) ;
 assign wire1887 = ( pinreg_40_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire1894 = ( pdata_33_  &  pc_10_  &  wire1902 ) | ( (~ pdata_33_)  &  (~ pc_10_)  &  wire1902 ) | ( pdata_33_  &  pc_10_  &  wire1903 ) | ( (~ pdata_33_)  &  (~ pc_10_)  &  wire1903 ) ;
 assign wire1895 = ( (~ pdata_33_)  &  pc_10_  &  wire626 ) | ( pdata_33_  &  (~ pc_10_)  &  wire626 ) ;
 assign wire1896 = ( pdata_34_  &  pc_23_  &  wire592  &  wire319 ) | ( (~ pdata_34_)  &  (~ pc_23_)  &  wire592  &  wire319 ) ;
 assign wire1897 = ( (~ pdata_32_)  &  pc_16_  &  wire568  &  wire7912 ) | ( pdata_32_  &  (~ pc_16_)  &  wire568  &  wire7912 ) ;
 assign wire1902 = ( pdata_36_  &  pc_4_  &  wire269  &  wire591 ) | ( (~ pdata_36_)  &  (~ pc_4_)  &  wire269  &  wire591 ) ;
 assign wire1903 = ( (~ pdata_32_)  &  pc_16_  &  n_n1701  &  wire7912 ) | ( pdata_32_  &  (~ pc_16_)  &  n_n1701  &  wire7912 ) ;
 assign wire1904 = ( (~ pdata_36_)  &  pc_4_  &  wire269  &  wire591 ) | ( pdata_36_  &  (~ pc_4_)  &  wire269  &  wire591 ) ;
 assign wire1905 = ( (~ n_n1706)  &  n_n1705  &  wire512 ) | ( n_n1706  &  (~ n_n1705)  &  wire512  &  n_n1703 ) ;
 assign wire1906 = ( (~ pdata_32_)  &  pc_16_  &  (~ n_n1701)  &  wire7912 ) | ( pdata_32_  &  (~ pc_16_)  &  (~ n_n1701)  &  wire7912 ) ;
 assign wire1913 = ( (~ n_n1706)  &  (~ n_n1705)  &  wire592  &  wire567 ) ;
 assign wire1914 = ( wire532  &  wire513  &  wire7908 ) ;
 assign wire1917 = ( (~ pdata_33_)  &  pc_10_  &  wire1920 ) | ( pdata_33_  &  (~ pc_10_)  &  wire1920 ) | ( (~ pdata_33_)  &  pc_10_  &  wire1921 ) | ( pdata_33_  &  (~ pc_10_)  &  wire1921 ) ;
 assign wire1918 = ( wire512  &  wire520  &  wire567 ) ;
 assign wire1919 = ( (~ n_n1706)  &  (~ n_n1705)  &  wire568  &  wire592 ) ;
 assign wire1920 = ( (~ pdata_32_)  &  pc_16_  &  (~ wire496)  &  wire513 ) | ( pdata_32_  &  (~ pc_16_)  &  (~ wire496)  &  wire513 ) ;
 assign wire1921 = ( pdata_32_  &  pc_16_  &  wire592  &  wire519 ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  wire592  &  wire519 ) ;
 assign wire1922 = ( wire594  &  wire532  &  wire520 ) ;
 assign wire1923 = ( (~ n_n1704)  &  wire1925 ) | ( (~ n_n1704)  &  (~ n_n1703)  &  wire722 ) ;
 assign wire1925 = ( pdata_32_  &  pc_16_  &  wire512  &  wire519 ) | ( (~ pdata_32_)  &  (~ pc_16_)  &  wire512  &  wire519 ) ;
 assign wire1929 = ( wire512  &  wire568  &  wire520 ) ;
 assign wire1930 = ( (~ wire496)  &  wire513  &  wire7908 ) ;
 assign wire1949 = ( (~ pdata_3_)  &  (~ n_n1327)  &  wire324 ) | ( (~ pdata_3_)  &  (~ n_n1327)  &  wire7905 ) | ( pdata_3_  &  (~ n_n1327)  &  (~ wire324)  &  (~ wire7905) ) ;
 assign wire1953 = ( wire245  &  wire313  &  wire7894 ) ;
 assign wire1955 = ( (~ n_n1717)  &  wire1962 ) | ( (~ n_n1717)  &  wire1964 ) | ( (~ n_n1717)  &  wire7898 ) ;
 assign wire1956 = ( n_n1715  &  n_n1717  &  wire517  &  wire528 ) ;
 assign wire1962 = ( (~ pd_22_)  &  pdata_53_  &  wire245  &  wire274 ) | ( pd_22_  &  (~ pdata_53_)  &  wire245  &  wire274 ) ;
 assign wire1964 = ( (~ pd_16_)  &  pdata_54_  &  n_n1713  &  wire528 ) | ( pd_16_  &  (~ pdata_54_)  &  n_n1713  &  wire528 ) ;
 assign wire1969 = ( n_n1715  &  n_n1717  &  wire505  &  wire558 ) ;
 assign wire1970 = ( (~ n_n1715)  &  n_n1717  &  wire284  &  wire7884 ) ;
 assign wire1973 = ( wire540  &  wire509  &  wire751 ) ;
 assign wire1977 = ( wire517  &  wire505  &  wire555 ) ;
 assign wire1978 = ( n_n1715  &  n_n1717  &  wire313  &  wire528 ) ;
 assign wire1979 = ( n_n1715  &  n_n1717  &  wire284  &  wire558 ) ;
 assign wire1980 = ( (~ n_n1715)  &  n_n1717  &  wire528  &  wire7884 ) ;
 assign wire1981 = ( n_n1715  &  n_n1717  &  wire737  &  wire7884 ) ;
 assign wire1982 = ( wire313  &  wire505  &  wire555 ) ;
 assign wire1983 = ( (~ n_n1715)  &  n_n1717  &  wire558  &  wire509 ) ;
 assign wire1996 = ( pd_0_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire1997 = ( pd_4_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire1998 = ( pd_1_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire1999 = ( pd_3_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2000 = ( (~ pencrypt_0_)  &  pinreg_38_  &  n_n1327  &  wire7712 ) ;
 assign wire2001 = ( pinreg_30_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2003 = ( pc_1_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2004 = ( pc_5_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2005 = ( pc_2_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2006 = ( pc_4_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2007 = ( (~ pencrypt_0_)  &  pinreg_24_  &  n_n1327  &  wire7712 ) ;
 assign wire2008 = ( pencrypt_0_  &  pinreg_16_  &  n_n1327  &  wire7712 ) ;
 assign wire2017 = ( (~ pdata_4_)  &  (~ n_n1327)  &  wire7871 ) | ( (~ pdata_4_)  &  (~ n_n1327)  &  wire7872 ) | ( pdata_4_  &  (~ n_n1327)  &  (~ wire7871)  &  (~ wire7872) ) ;
 assign wire2021 = ( (~ n_n1729)  &  wire531  &  wire7856 ) | ( (~ n_n1729)  &  wire295  &  wire7856 ) ;
 assign wire2022 = ( n_n1725  &  wire2032 ) | ( n_n1725  &  wire2033 ) | ( n_n1725  &  wire2034 ) ;
 assign wire2023 = ( pdata_59_  &  pd_17_  &  wire531  &  wire511 ) | ( (~ pdata_59_)  &  (~ pd_17_)  &  wire531  &  wire511 ) ;
 assign wire2025 = ( n_n1726  &  n_n1729  &  wire297  &  wire7846 ) ;
 assign wire2026 = ( n_n1726  &  (~ n_n1728)  &  wire562  &  wire7863 ) ;
 assign wire2027 = ( (~ n_n1726)  &  (~ n_n1730)  &  (~ n_n1727)  &  wire511 ) ;
 assign wire2032 = ( (~ pdata_59_)  &  pd_17_  &  wire295  &  wire511 ) | ( pdata_59_  &  (~ pd_17_)  &  wire295  &  wire511 ) ;
 assign wire2033 = ( (~ n_n1726)  &  n_n1727  &  (~ n_n1729)  &  wire7856 ) ;
 assign wire2034 = ( pd_7_  &  pdata_62_  &  wire506  &  wire7850 ) | ( (~ pd_7_)  &  (~ pdata_62_)  &  wire506  &  wire7850 ) ;
 assign wire2035 = ( wire543  &  wire743  &  wire7860 ) ;
 assign wire2036 = ( n_n1726  &  n_n1730  &  wire297  &  wire511 ) ;
 assign wire2037 = ( n_n1726  &  (~ n_n1729)  &  wire562  &  wire7856 ) ;
 assign wire2038 = ( n_n1725  &  n_n1729  &  wire506  &  wire295 ) ;
 assign wire2039 = ( (~ n_n1726)  &  (~ n_n1729)  &  wire297  &  wire7856 ) ;
 assign wire2040 = ( n_n1726  &  (~ n_n1730)  &  wire297  &  wire511 ) ;
 assign wire2041 = ( wire543  &  wire562  &  wire7857 ) ;
 assign wire2044 = ( (~ n_n1725)  &  n_n1730  &  wire543  &  wire295 ) ;
 assign wire2046 = ( wire297  &  wire506  &  wire7850 ) ;
 assign wire2048 = ( (~ n_n1726)  &  n_n1730  &  wire588  &  wire511 ) ;
 assign wire2049 = ( (~ n_n1725)  &  (~ n_n1729)  &  wire506  &  wire295 ) ;
 assign wire2050 = ( wire295  &  wire7844  &  wire7845 ) ;
 assign wire2051 = ( (~ n_n1726)  &  n_n1729  &  wire531  &  wire7846 ) ;
 assign wire2066 = ( pd_27_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2067 = ( pd_3_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2068 = ( pd_0_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2069 = ( pd_2_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2070 = ( (~ pencrypt_0_)  &  pinreg_46_  &  n_n1327  &  wire7712 ) ;
 assign wire2071 = ( pencrypt_0_  &  pinreg_38_  &  n_n1327  &  wire7712 ) ;
 assign wire2073 = ( pc_0_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2074 = ( pc_4_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2075 = ( pc_1_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2076 = ( pc_3_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2077 = ( pinreg_32_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire2078 = ( pencrypt_0_  &  pinreg_24_  &  n_n1327  &  wire7712 ) ;
 assign wire2091 = ( pd_2_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2092 = ( pd_6_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2093 = ( pd_3_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2094 = ( pd_5_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2095 = ( (~ pencrypt_0_)  &  pinreg_22_  &  n_n1327  &  wire7712 ) ;
 assign wire2096 = ( pencrypt_0_  &  pinreg_14_  &  n_n1327  &  wire7712 ) ;
 assign wire2098 = ( pc_3_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2099 = ( pc_7_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2100 = ( pc_4_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2101 = ( pc_6_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2102 = ( pinreg_8_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire2103 = ( pinreg_0_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2110 = ( pdata_59_  &  pd_5_  &  wire306  &  wire518 ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  wire306  &  wire518 ) ;
 assign wire2111 = ( n_n1723  &  n_n1721  &  wire315  &  wire586 ) | ( (~ n_n1723)  &  (~ n_n1721)  &  wire315  &  wire586 ) ;
 assign wire2112 = ( n_n1720  &  wire428 ) | ( n_n1720  &  n_n1719  &  wire643 ) ;
 assign wire2113 = ( n_n1721  &  wire2123 ) | ( n_n1721  &  wire2124 ) | ( n_n1721  &  wire2125 ) ;
 assign wire2123 = ( (~ pd_20_)  &  pdata_56_  &  wire246  &  (~ wire271) ) | ( pd_20_  &  (~ pdata_56_)  &  wire246  &  (~ wire271) ) ;
 assign wire2124 = ( pd_20_  &  pdata_56_  &  wire529  &  wire586 ) | ( (~ pd_20_)  &  (~ pdata_56_)  &  wire529  &  wire586 ) ;
 assign wire2125 = ( pd_20_  &  pdata_56_  &  wire315  &  (~ wire417) ) | ( (~ pd_20_)  &  (~ pdata_56_)  &  wire315  &  (~ wire417) ) ;
 assign wire2127 = ( wire306  &  wire715 ) ;
 assign wire2143 = ( pd_1_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2144 = ( pd_5_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2145 = ( pd_2_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2146 = ( pd_4_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2147 = ( pinreg_30_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire2148 = ( pencrypt_0_  &  pinreg_22_  &  n_n1327  &  wire7712 ) ;
 assign wire2150 = ( pc_2_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2151 = ( pc_6_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2152 = ( pc_3_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2153 = ( pc_5_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2154 = ( (~ pencrypt_0_)  &  pinreg_16_  &  n_n1327  &  wire7712 ) ;
 assign wire2155 = ( pinreg_8_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2162 = ( (~ pd_2_)  &  pdata_49_  &  wire666 ) | ( pd_2_  &  (~ pdata_49_)  &  wire666 ) ;
 assign wire2167 = ( n_n1696  &  (~ n_n1695)  &  n_n1697  &  wire7791 ) | ( (~ n_n1696)  &  n_n1695  &  (~ n_n1697)  &  wire7791 ) ;
 assign wire2169 = ( (~ pd_8_)  &  pdata_50_  &  wire289  &  wire262 ) | ( pd_8_  &  (~ pdata_50_)  &  wire289  &  wire262 ) ;
 assign wire2175 = ( wire304  &  wire7794 ) ;
 assign wire2182 = ( wire516  &  wire303  &  wire539 ) ;
 assign wire2184 = ( wire552  &  wire579  &  wire7771 ) ;
 assign wire2195 = ( wire631  &  wire579  &  wire7771 ) ;
 assign wire2198 = ( pd_8_  &  pdata_50_  &  wire527  &  wire7783 ) | ( (~ pd_8_)  &  (~ pdata_50_)  &  wire527  &  wire7783 ) ;
 assign wire2202 = ( (~ n_n1696)  &  (~ n_n1700)  &  n_n1697  &  wire289 ) | ( (~ n_n1696)  &  n_n1700  &  (~ n_n1697)  &  wire289 ) | ( n_n1696  &  (~ n_n1700)  &  (~ n_n1697)  &  wire289 ) ;
 assign wire2208 = ( (~ pdata_47_)  &  pd_12_  &  wire261  &  wire635 ) | ( pdata_47_  &  (~ pd_12_)  &  wire261  &  wire635 ) ;
 assign wire2209 = ( pdata_47_  &  pd_12_  &  wire283  &  wire304 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire283  &  wire304 ) ;
 assign wire2210 = ( pdata_47_  &  pd_12_  &  n_n1695  &  wire303 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  n_n1695  &  wire303 ) ;
 assign wire2211 = ( wire289  &  wire303 ) ;
 assign wire2212 = ( wire283  &  wire516  &  wire539 ) ;
 assign wire2214 = ( wire504  &  wire516  &  wire7776 ) ;
 assign wire2218 = ( wire283  &  wire516  &  wire7776 ) ;
 assign wire2219 = ( wire504  &  wire579  &  wire7772 ) ;
 assign wire2222 = ( (~ n_n1700)  &  n_n1698  &  wire552  &  wire516 ) ;
 assign wire2223 = ( wire504  &  wire579  &  wire7771 ) ;
 assign wire2224 = ( wire283  &  wire304  &  (~ wire420) ) ;
 assign wire2225 = ( wire579  &  wire303  &  wire7772 ) ;
 assign wire2227 = ( wire539  &  wire726 ) ;
 assign wire2228 = ( pd_2_  &  pdata_49_  &  wire2231 ) | ( (~ pd_2_)  &  (~ pdata_49_)  &  wire2231 ) | ( pd_2_  &  pdata_49_  &  wire2232 ) | ( (~ pd_2_)  &  (~ pdata_49_)  &  wire2232 ) ;
 assign wire2231 = ( pdata_47_  &  pd_12_  &  wire304  &  wire303 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire304  &  wire303 ) ;
 assign wire2232 = ( pdata_47_  &  pd_12_  &  wire289  &  wire552 ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  wire289  &  wire552 ) ;
 assign wire2249 = ( pd_17_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2250 = ( pd_21_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2251 = ( pd_18_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2252 = ( pd_20_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2253 = ( (~ pencrypt_0_)  &  pinreg_28_  &  n_n1327  &  wire7712 ) ;
 assign wire2254 = ( pencrypt_0_  &  pinreg_20_  &  n_n1327  &  wire7712 ) ;
 assign wire2256 = ( pd_4_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2257 = ( pd_8_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2258 = ( pd_5_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2259 = ( pd_7_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2260 = ( pinreg_6_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire2261 = ( pdata_in_6_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2263 = ( pc_5_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2264 = ( pc_9_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2265 = ( pc_6_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2266 = ( pc_8_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2267 = ( (~ pencrypt_0_)  &  pdata_in_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2268 = ( pencrypt_0_  &  pinreg_49_  &  n_n1327  &  wire7712 ) ;
 assign wire2275 = ( pd_20_  &  pdata_56_  &  wire529  &  wire646 ) | ( (~ pd_20_)  &  (~ pdata_56_)  &  wire529  &  wire646 ) ;
 assign wire2276 = ( (~ n_n1723)  &  (~ n_n1721)  &  wire586  &  wire7741 ) ;
 assign wire2277 = ( (~ n_n1724)  &  n_n1721  &  wire315  &  wire584 ) ;
 assign wire2278 = ( wire306  &  wire417  &  wire541 ) ;
 assign wire2293 = ( (~ pdata_60_)  &  pd_24_  &  wire2294 ) | ( pdata_60_  &  (~ pd_24_)  &  wire2294 ) | ( (~ pdata_60_)  &  pd_24_  &  wire2295 ) | ( pdata_60_  &  (~ pd_24_)  &  wire2295 ) ;
 assign wire2294 = ( pd_27_  &  pdata_58_  &  wire518  &  wire510 ) | ( (~ pd_27_)  &  (~ pdata_58_)  &  wire518  &  wire510 ) ;
 assign wire2295 = ( (~ pd_27_)  &  pdata_58_  &  wire7731  &  wire7732 ) | ( pd_27_  &  (~ pdata_58_)  &  wire7731  &  wire7732 ) ;
 assign wire2304 = ( n_n1719  &  n_n1721  &  wire518  &  wire584 ) ;
 assign wire2306 = ( wire315  &  (~ wire417)  &  wire585 ) ;
 assign wire2309 = ( wire529  &  wire510  &  wire7733 ) ;
 assign wire2311 = ( (~ n_n1723)  &  n_n1721  &  wire315  &  wire586 ) ;
 assign wire2334 = ( pd_3_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2335 = ( pd_7_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2336 = ( pd_4_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2337 = ( pd_6_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2338 = ( (~ pencrypt_0_)  &  pinreg_14_  &  n_n1327  &  wire7712 ) ;
 assign wire2339 = ( pinreg_6_  &  pencrypt_0_  &  n_n1327  &  wire7712 ) ;
 assign wire2341 = ( pc_17_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2342 = ( pc_21_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2343 = ( pc_18_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2344 = ( pc_20_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2345 = ( (~ pencrypt_0_)  &  pinreg_26_  &  n_n1327  &  wire7712 ) ;
 assign wire2346 = ( pencrypt_0_  &  pinreg_18_  &  n_n1327  &  wire7712 ) ;
 assign wire2348 = ( pc_4_  &  wire514  &  (~ n_n1329)  &  wire7710 ) ;
 assign wire2349 = ( pc_8_  &  wire514  &  (~ n_n1329)  &  wire7711 ) ;
 assign wire2350 = ( pc_5_  &  wire514  &  n_n1329  &  wire7710 ) ;
 assign wire2351 = ( pc_7_  &  wire514  &  n_n1329  &  wire7711 ) ;
 assign wire2352 = ( pinreg_0_  &  (~ pencrypt_0_)  &  n_n1327  &  wire7712 ) ;
 assign wire2353 = ( pencrypt_0_  &  pdata_in_0_  &  n_n1327  &  wire7712 ) ;
 assign wire7710 = ( (~ pencrypt_0_)  &  (~ pencrypt_mode_0_) ) | ( (~ pencrypt_mode_0_)  &  (~ n_n1327) ) ;
 assign wire7711 = ( pencrypt_0_  &  pencrypt_mode_0_ ) | ( pencrypt_mode_0_  &  (~ n_n1327) ) ;
 assign wire7712 = ( pload_key_0_  &  (~ preset_0_) ) ;
 assign wire7714 = ( wire2352 ) | ( wire2353 ) | ( pc_6_  &  wire254 ) ;
 assign wire7717 = ( wire2348 ) | ( wire2349 ) | ( wire7714 ) ;
 assign wire7719 = ( wire2345 ) | ( wire2346 ) | ( pc_19_  &  wire254 ) ;
 assign wire7722 = ( wire2341 ) | ( wire2342 ) | ( wire7719 ) ;
 assign wire7724 = ( wire2338 ) | ( wire2339 ) | ( pd_5_  &  wire254 ) ;
 assign wire7727 = ( wire2334 ) | ( wire2335 ) | ( wire7724 ) ;
 assign wire7729 = ( pd_10_  &  pdata_60_  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  (~ pdata_60_)  &  (~ pd_24_)  &  pdata_57_ ) | ( (~ pd_10_)  &  pdata_60_  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire7731 = ( pd_10_  &  pd_15_  &  pdata_57_  &  pdata_55_ ) | ( (~ pd_10_)  &  pd_15_  &  (~ pdata_57_)  &  pdata_55_ ) | ( pd_10_  &  (~ pd_15_)  &  pdata_57_  &  (~ pdata_55_) ) | ( (~ pd_10_)  &  (~ pd_15_)  &  (~ pdata_57_)  &  (~ pdata_55_) ) ;
 assign wire7732 = ( pdata_59_  &  pd_20_  &  pd_5_  &  pdata_56_ ) | ( (~ pdata_59_)  &  pd_20_  &  (~ pd_5_)  &  pdata_56_ ) | ( pdata_59_  &  (~ pd_20_)  &  pd_5_  &  (~ pdata_56_) ) | ( (~ pdata_59_)  &  (~ pd_20_)  &  (~ pd_5_)  &  (~ pdata_56_) ) ;
 assign wire7733 = ( (~ pd_27_)  &  (~ pd_15_)  &  pdata_58_  &  pdata_55_ ) | ( pd_27_  &  (~ pd_15_)  &  (~ pdata_58_)  &  pdata_55_ ) | ( (~ pd_27_)  &  pd_15_  &  pdata_58_  &  (~ pdata_55_) ) | ( pd_27_  &  pd_15_  &  (~ pdata_58_)  &  (~ pdata_55_) ) ;
 assign wire7738 = ( (~ pdata_59_)  &  pd_5_  &  (~ pd_15_)  &  pdata_55_ ) | ( pdata_59_  &  (~ pd_5_)  &  (~ pd_15_)  &  pdata_55_ ) | ( (~ pdata_59_)  &  pd_5_  &  pd_15_  &  (~ pdata_55_) ) | ( pdata_59_  &  (~ pd_5_)  &  pd_15_  &  (~ pdata_55_) ) ;
 assign wire7741 = ( pd_10_  &  pdata_60_  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  (~ pdata_60_)  &  (~ pd_24_)  &  pdata_57_ ) | ( (~ pd_10_)  &  pdata_60_  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire7744 = ( pdata_60_  &  pd_24_  &  pd_15_  &  pdata_55_ ) | ( (~ pdata_60_)  &  (~ pd_24_)  &  pd_15_  &  pdata_55_ ) | ( pdata_60_  &  pd_24_  &  (~ pd_15_)  &  (~ pdata_55_) ) | ( (~ pdata_60_)  &  (~ pd_24_)  &  (~ pd_15_)  &  (~ pdata_55_) ) ;
 assign wire7745 = ( (~ pd_20_)  &  (~ pd_27_)  &  pdata_58_  &  pdata_56_ ) | ( (~ pd_20_)  &  pd_27_  &  (~ pdata_58_)  &  pdata_56_ ) | ( pd_20_  &  (~ pd_27_)  &  pdata_58_  &  (~ pdata_56_) ) | ( pd_20_  &  pd_27_  &  (~ pdata_58_)  &  (~ pdata_56_) ) ;
 assign wire7747 = ( wire2278 ) | ( n_n1722  &  wire586  &  wire7745 ) ;
 assign wire7748 = ( wire402 ) | ( wire2276 ) | ( wire2277 ) ;
 assign wire7751 = ( wire7748 ) | ( pdata_59_  &  pd_5_  &  wire645 ) | ( (~ pdata_59_)  &  (~ pd_5_)  &  wire645 ) ;
 assign wire7752 = ( wire472 ) | ( wire2293 ) | ( wire747  &  wire7729 ) ;
 assign wire7753 = ( wire335 ) | ( wire401 ) | ( wire2275 ) | ( wire7747 ) ;
 assign wire7755 = ( (~ pcount_0_)  &  poutreg_9_ ) | ( pcount_0_  &  poutreg_17_  &  (~ wire577) ) ;
 assign wire7757 = ( wire2267 ) | ( wire2268 ) | ( pc_7_  &  wire254 ) ;
 assign wire7760 = ( wire2263 ) | ( wire2264 ) | ( wire7757 ) ;
 assign wire7762 = ( wire2260 ) | ( wire2261 ) | ( pd_6_  &  wire254 ) ;
 assign wire7765 = ( wire2256 ) | ( wire2257 ) | ( wire7762 ) ;
 assign wire7767 = ( wire2253 ) | ( wire2254 ) | ( pd_19_  &  wire254 ) ;
 assign wire7770 = ( wire2249 ) | ( wire2250 ) | ( wire7767 ) ;
 assign wire7771 = ( pdata_48_  &  pd_23_  &  pd_26_  &  pdata_52_ ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  pd_26_  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  (~ pd_26_)  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  (~ pd_26_)  &  (~ pdata_52_) ) ;
 assign wire7772 = ( pdata_48_  &  pd_23_  &  (~ pd_26_)  &  pdata_52_ ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  (~ pd_26_)  &  pdata_52_ ) | ( pdata_48_  &  pd_23_  &  pd_26_  &  (~ pdata_52_) ) | ( (~ pdata_48_)  &  (~ pd_23_)  &  pd_26_  &  (~ pdata_52_) ) ;
 assign wire7775 = ( wire2222 ) | ( wire2223 ) | ( wire2224 ) | ( wire2225 ) ;
 assign wire7776 = ( pdata_47_  &  pd_12_  &  pd_2_  &  pdata_49_ ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  pd_2_  &  pdata_49_ ) | ( pdata_47_  &  pd_12_  &  (~ pd_2_)  &  (~ pdata_49_) ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  (~ pd_2_)  &  (~ pdata_49_) ) ;
 assign wire7783 = ( pdata_47_  &  pd_12_  &  (~ pd_18_)  &  pdata_51_ ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  (~ pd_18_)  &  pdata_51_ ) | ( pdata_47_  &  pd_12_  &  pd_18_  &  (~ pdata_51_) ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  pd_18_  &  (~ pdata_51_) ) ;
 assign wire7785 = ( wire467 ) | ( wire2195 ) | ( wire2198 ) ;
 assign wire7786 = ( wire471 ) | ( wire2227 ) | ( wire2228 ) | ( wire7775 ) ;
 assign wire7787 = ( pd_2_  &  pdata_49_  &  wire634 ) | ( (~ pd_2_)  &  (~ pdata_49_)  &  wire634 ) | ( (~ pd_2_)  &  pdata_49_  &  wire632 ) | ( pd_2_  &  (~ pdata_49_)  &  wire632 ) ;
 assign wire7791 = ( pdata_48_  &  pdata_47_  &  pd_12_  &  pd_23_ ) | ( pdata_48_  &  (~ pdata_47_)  &  (~ pd_12_)  &  pd_23_ ) | ( (~ pdata_48_)  &  pdata_47_  &  pd_12_  &  (~ pd_23_) ) | ( (~ pdata_48_)  &  (~ pdata_47_)  &  (~ pd_12_)  &  (~ pd_23_) ) ;
 assign wire7793 = ( pdata_47_  &  pd_12_  &  pd_26_  &  pdata_52_ ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  pd_26_  &  pdata_52_ ) | ( pdata_47_  &  pd_12_  &  (~ pd_26_)  &  (~ pdata_52_) ) | ( (~ pdata_47_)  &  (~ pd_12_)  &  (~ pd_26_)  &  (~ pdata_52_) ) ;
 assign wire7794 = ( (~ pdata_47_)  &  pd_12_  &  (~ pd_8_)  &  pdata_50_ ) | ( pdata_47_  &  (~ pd_12_)  &  (~ pd_8_)  &  pdata_50_ ) | ( (~ pdata_47_)  &  pd_12_  &  pd_8_  &  (~ pdata_50_) ) | ( pdata_47_  &  (~ pd_12_)  &  pd_8_  &  (~ pdata_50_) ) ;
 assign wire7795 = ( (~ n_n1696)  &  (~ n_n1697)  &  wire289 ) | ( n_n1696  &  (~ n_n1697)  &  wire7793 ) ;
 assign wire7799 = ( wire467 ) | ( wire336 ) | ( (~ n_n1698)  &  wire669 ) ;
 assign wire7800 = ( (~ pcount_0_)  &  poutreg_19_ ) | ( pcount_0_  &  poutreg_27_  &  (~ wire577) ) ;
 assign wire7802 = ( wire2154 ) | ( wire2155 ) | ( pc_4_  &  wire254 ) ;
 assign wire7805 = ( wire2150 ) | ( wire2151 ) | ( wire7802 ) ;
 assign wire7807 = ( wire2147 ) | ( wire2148 ) | ( pd_3_  &  wire254 ) ;
 assign wire7810 = ( wire2143 ) | ( wire2144 ) | ( wire7807 ) ;
 assign wire7816 = ( wire472 ) | ( wire2293 ) | ( wire747  &  wire7729 ) ;
 assign wire7819 = ( wire2110 ) | ( wire2111 ) | ( wire2112 ) | ( wire2113 ) ;
 assign wire7820 = ( (~ pcount_0_)  &  poutreg_7_ ) | ( pcount_0_  &  poutreg_15_  &  (~ wire577) ) ;
 assign wire7822 = ( wire2102 ) | ( wire2103 ) | ( pc_5_  &  wire254 ) ;
 assign wire7825 = ( wire2098 ) | ( wire2099 ) | ( wire7822 ) ;
 assign wire7827 = ( wire2095 ) | ( wire2096 ) | ( pd_4_  &  wire254 ) ;
 assign wire7830 = ( wire2091 ) | ( wire2092 ) | ( wire7827 ) ;
 assign wire7831 = ( pcount_0_  &  pdata_38_  &  wire577 ) | ( pcount_0_  &  poutreg_16_  &  (~ wire577) ) ;
 assign wire7833 = ( wire2077 ) | ( wire2078 ) | ( pc_2_  &  wire254 ) ;
 assign wire7836 = ( wire2073 ) | ( wire2074 ) | ( wire7833 ) ;
 assign wire7838 = ( wire2070 ) | ( wire2071 ) | ( pd_1_  &  wire254 ) ;
 assign wire7841 = ( wire2066 ) | ( wire2067 ) | ( wire7838 ) ;
 assign wire7844 = ( (~ pdata_32_)  &  pdata_60_  &  pd_13_  &  pd_3_ ) | ( (~ pdata_32_)  &  (~ pdata_60_)  &  (~ pd_13_)  &  pd_3_ ) | ( pdata_32_  &  pdata_60_  &  pd_13_  &  (~ pd_3_) ) | ( pdata_32_  &  (~ pdata_60_)  &  (~ pd_13_)  &  (~ pd_3_) ) ;
 assign wire7845 = ( pdata_59_  &  pd_21_  &  pd_17_  &  pdata_61_ ) | ( (~ pdata_59_)  &  pd_21_  &  (~ pd_17_)  &  pdata_61_ ) | ( pdata_59_  &  (~ pd_21_)  &  pd_17_  &  (~ pdata_61_) ) | ( (~ pdata_59_)  &  (~ pd_21_)  &  (~ pd_17_)  &  (~ pdata_61_) ) ;
 assign wire7846 = ( (~ pdata_59_)  &  (~ pd_21_)  &  pd_17_  &  pdata_61_ ) | ( pdata_59_  &  (~ pd_21_)  &  (~ pd_17_)  &  pdata_61_ ) | ( (~ pdata_59_)  &  pd_21_  &  pd_17_  &  (~ pdata_61_) ) | ( pdata_59_  &  pd_21_  &  (~ pd_17_)  &  (~ pdata_61_) ) ;
 assign wire7850 = ( pdata_60_  &  pd_13_  &  pd_0_  &  pdata_63_ ) | ( (~ pdata_60_)  &  (~ pd_13_)  &  pd_0_  &  pdata_63_ ) | ( pdata_60_  &  pd_13_  &  (~ pd_0_)  &  (~ pdata_63_) ) | ( (~ pdata_60_)  &  (~ pd_13_)  &  (~ pd_0_)  &  (~ pdata_63_) ) ;
 assign wire7852 = ( wire2044 ) | ( wire2046 ) | ( wire316  &  wire713 ) ;
 assign wire7853 = ( (~ pd_7_)  &  pd_0_  &  pdata_62_  &  pdata_63_ ) | ( pd_7_  &  pd_0_  &  (~ pdata_62_)  &  pdata_63_ ) | ( (~ pd_7_)  &  (~ pd_0_)  &  pdata_62_  &  (~ pdata_63_) ) | ( pd_7_  &  (~ pd_0_)  &  (~ pdata_62_)  &  (~ pdata_63_) ) ;
 assign wire7856 = ( (~ pdata_59_)  &  (~ pd_21_)  &  pd_17_  &  pdata_61_ ) | ( pdata_59_  &  (~ pd_21_)  &  (~ pd_17_)  &  pdata_61_ ) | ( (~ pdata_59_)  &  pd_21_  &  pd_17_  &  (~ pdata_61_) ) | ( pdata_59_  &  pd_21_  &  (~ pd_17_)  &  (~ pdata_61_) ) ;
 assign wire7857 = ( (~ pdata_59_)  &  pd_17_  &  pd_0_  &  pdata_63_ ) | ( pdata_59_  &  (~ pd_17_)  &  pd_0_  &  pdata_63_ ) | ( (~ pdata_59_)  &  pd_17_  &  (~ pd_0_)  &  (~ pdata_63_) ) | ( pdata_59_  &  (~ pd_17_)  &  (~ pd_0_)  &  (~ pdata_63_) ) ;
 assign wire7860 = ( pdata_59_  &  pd_17_  &  pd_0_  &  pdata_63_ ) | ( (~ pdata_59_)  &  (~ pd_17_)  &  pd_0_  &  pdata_63_ ) | ( pdata_59_  &  pd_17_  &  (~ pd_0_)  &  (~ pdata_63_) ) | ( (~ pdata_59_)  &  (~ pd_17_)  &  (~ pd_0_)  &  (~ pdata_63_) ) ;
 assign wire7863 = ( pdata_59_  &  pd_17_  &  pdata_60_  &  pd_13_ ) | ( (~ pdata_59_)  &  (~ pd_17_)  &  pdata_60_  &  pd_13_ ) | ( pdata_59_  &  pd_17_  &  (~ pdata_60_)  &  (~ pd_13_) ) | ( (~ pdata_59_)  &  (~ pd_17_)  &  (~ pdata_60_)  &  (~ pd_13_) ) ;
 assign wire7865 = ( wire2023 ) | ( wire297  &  wire543  &  wire7860 ) ;
 assign wire7866 = ( wire2026 ) | ( wire2025 ) ;
 assign wire7867 = ( wire396 ) | ( wire2021 ) | ( wire2027 ) ;
 assign wire7871 = ( wire475 ) | ( wire7865 ) | ( wire7866 ) | ( wire7867 ) ;
 assign wire7872 = ( wire470 ) | ( wire413 ) | ( wire2022 ) | ( wire7852 ) ;
 assign wire7873 = ( pdata_37_  &  pcount_0_  &  wire577 ) | ( pcount_0_  &  poutreg_24_  &  (~ wire577) ) ;
 assign wire7875 = ( wire2007 ) | ( wire2008 ) | ( pc_3_  &  wire254 ) ;
 assign wire7878 = ( wire2003 ) | ( wire2004 ) | ( wire7875 ) ;
 assign wire7880 = ( wire2000 ) | ( wire2001 ) | ( pd_2_  &  wire254 ) ;
 assign wire7883 = ( wire1996 ) | ( wire1997 ) | ( wire7880 ) ;
 assign wire7884 = ( (~ pd_22_)  &  pd_19_  &  pdata_53_  &  pdata_56_ ) | ( pd_22_  &  pd_19_  &  (~ pdata_53_)  &  pdata_56_ ) | ( (~ pd_22_)  &  (~ pd_19_)  &  pdata_53_  &  (~ pdata_56_) ) | ( pd_22_  &  (~ pd_19_)  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire7894 = ( (~ pd_11_)  &  (~ pd_16_)  &  pdata_54_  &  pdata_52_ ) | ( (~ pd_11_)  &  pd_16_  &  (~ pdata_54_)  &  pdata_52_ ) | ( pd_11_  &  (~ pd_16_)  &  pdata_54_  &  (~ pdata_52_) ) | ( pd_11_  &  pd_16_  &  (~ pdata_54_)  &  (~ pdata_52_) ) ;
 assign wire7898 = ( (~ n_n1716)  &  (~ n_n1713)  &  wire284 ) | ( n_n1715  &  n_n1716  &  n_n1713  &  wire284 ) ;
 assign wire7900 = ( (~ pd_22_)  &  pd_19_  &  pdata_53_  &  pdata_56_ ) | ( pd_22_  &  pd_19_  &  (~ pdata_53_)  &  pdata_56_ ) | ( (~ pd_22_)  &  (~ pd_19_)  &  pdata_53_  &  (~ pdata_56_) ) | ( pd_22_  &  (~ pd_19_)  &  (~ pdata_53_)  &  (~ pdata_56_) ) ;
 assign wire7901 = ( wire1953 ) | ( wire305  &  wire528  &  wire7900 ) ;
 assign wire7902 = ( wire1956 ) | ( wire305  &  wire655 ) ;
 assign wire7905 = ( wire407 ) | ( wire1955 ) | ( wire7901 ) | ( wire7902 ) ;
 assign wire7908 = ( pdata_32_  &  (~ pdata_33_)  &  pc_10_  &  pc_16_ ) | ( pdata_32_  &  pdata_33_  &  (~ pc_10_)  &  pc_16_ ) | ( (~ pdata_32_)  &  (~ pdata_33_)  &  pc_10_  &  (~ pc_16_) ) | ( (~ pdata_32_)  &  pdata_33_  &  (~ pc_10_)  &  (~ pc_16_) ) ;
 assign wire7912 = ( pdata_35_  &  (~ pc_13_)  &  pc_0_  &  pdata_63_ ) | ( (~ pdata_35_)  &  (~ pc_13_)  &  (~ pc_0_)  &  pdata_63_ ) | ( pdata_35_  &  pc_13_  &  pc_0_  &  (~ pdata_63_) ) | ( (~ pdata_35_)  &  pc_13_  &  (~ pc_0_)  &  (~ pdata_63_) ) ;
 assign wire7919 = ( wire1894 ) | ( wire1917 ) | ( wire1918 ) | ( wire1919 ) ;
 assign wire7920 = ( wire465 ) | ( wire333 ) | ( wire1896 ) | ( wire1897 ) ;
 assign wire7923 = ( (~ pcount_0_)  &  poutreg_15_ ) | ( pcount_0_  &  poutreg_23_  &  (~ wire577) ) ;
 assign wire7925 = ( wire1886 ) | ( wire1887 ) | ( pc_0_  &  wire254 ) ;
 assign wire7928 = ( wire1882 ) | ( wire1883 ) | ( wire7925 ) ;
 assign wire7929 = ( pcount_0_  &  pdata_45_  &  wire577 ) | ( pcount_0_  &  poutreg_26_  &  (~ wire577) ) ;
 assign wire7931 = ( wire1868 ) | ( wire1869 ) | ( pc_1_  &  wire254 ) ;
 assign wire7934 = ( wire1864 ) | ( wire1865 ) | ( wire7931 ) ;
 assign wire7936 = ( wire1861 ) | ( wire1862 ) | ( pd_0_  &  wire254 ) ;
 assign wire7939 = ( wire1857 ) | ( wire1858 ) | ( wire7936 ) ;
 assign wire7943 = ( (~ pdata_43_)  &  (~ pdata_41_)  &  pc_11_  &  pc_25_ ) | ( (~ pdata_43_)  &  pdata_41_  &  (~ pc_11_)  &  pc_25_ ) | ( pdata_43_  &  (~ pdata_41_)  &  pc_11_  &  (~ pc_25_) ) | ( pdata_43_  &  pdata_41_  &  (~ pc_11_)  &  (~ pc_25_) ) ;
 assign wire7946 = ( wire1835 ) | ( wire1834 ) ;
 assign wire7948 = ( (~ pdata_43_)  &  pdata_42_  &  pc_25_  &  pc_3_ ) | ( pdata_43_  &  pdata_42_  &  (~ pc_25_)  &  pc_3_ ) | ( (~ pdata_43_)  &  (~ pdata_42_)  &  pc_25_  &  (~ pc_3_) ) | ( pdata_43_  &  (~ pdata_42_)  &  (~ pc_25_)  &  (~ pc_3_) ) ;
 assign wire7949 = ( pdata_44_  &  (~ pdata_41_)  &  pc_11_  &  pc_7_ ) | ( pdata_44_  &  pdata_41_  &  (~ pc_11_)  &  pc_7_ ) | ( (~ pdata_44_)  &  (~ pdata_41_)  &  pc_11_  &  (~ pc_7_) ) | ( (~ pdata_44_)  &  pdata_41_  &  (~ pc_11_)  &  (~ pc_7_) ) ;
 assign wire7952 = ( wire480 ) | ( wire508  &  wire549  &  wire515 ) ;
 assign wire7953 = ( wire398 ) | ( wire1834 ) | ( wire1835 ) | ( wire1836 ) ;
 assign wire7960 = ( (~ pdata_43_)  &  (~ pc_22_)  &  pc_25_  &  pdata_39_ ) | ( pdata_43_  &  (~ pc_22_)  &  (~ pc_25_)  &  pdata_39_ ) | ( (~ pdata_43_)  &  pc_22_  &  pc_25_  &  (~ pdata_39_) ) | ( pdata_43_  &  pc_22_  &  (~ pc_25_)  &  (~ pdata_39_) ) ;
 assign wire7962 = ( (~ pdata_42_)  &  pc_22_  &  pc_3_  &  pdata_39_ ) | ( pdata_42_  &  pc_22_  &  (~ pc_3_)  &  pdata_39_ ) | ( (~ pdata_42_)  &  (~ pc_22_)  &  pc_3_  &  (~ pdata_39_) ) | ( pdata_42_  &  (~ pc_22_)  &  (~ pc_3_)  &  (~ pdata_39_) ) ;
 assign wire7966 = ( wire474 ) | ( wire1806 ) | ( wire1810 ) ;
 assign wire7967 = ( wire1805 ) | ( wire1807 ) | ( wire1808 ) | ( wire1809 ) ;
 assign wire7969 = ( (~ pcount_0_)  &  poutreg_17_ ) | ( pcount_0_  &  poutreg_25_  &  (~ wire577) ) ;
 assign wire7971 = ( wire1791 ) | ( wire1792 ) | ( pc_11_  &  wire254 ) ;
 assign wire7974 = ( wire1787 ) | ( wire1788 ) | ( wire7971 ) ;
 assign wire7976 = ( wire1784 ) | ( wire1785 ) | ( pc_22_  &  wire254 ) ;
 assign wire7979 = ( wire1780 ) | ( wire1781 ) | ( wire7976 ) ;
 assign wire7981 = ( wire1777 ) | ( wire1778 ) | ( pd_12_  &  wire254 ) ;
 assign wire7984 = ( wire1773 ) | ( wire1774 ) | ( wire7981 ) ;
 assign wire7986 = ( wire1770 ) | ( wire1771 ) | ( pd_23_  &  wire254 ) ;
 assign wire7989 = ( wire1766 ) | ( wire1767 ) | ( wire7986 ) ;
 assign wire7996 = ( (~ pdata_60_)  &  pd_13_  &  pd_0_  &  pdata_63_ ) | ( pdata_60_  &  (~ pd_13_)  &  pd_0_  &  pdata_63_ ) | ( (~ pdata_60_)  &  pd_13_  &  (~ pd_0_)  &  (~ pdata_63_) ) | ( pdata_60_  &  (~ pd_13_)  &  (~ pd_0_)  &  (~ pdata_63_) ) ;
 assign wire8000 = ( wire1747 ) | ( wire1746 ) ;
 assign wire8001 = ( wire381 ) | ( wire1741 ) | ( wire1744 ) | ( wire1745 ) ;
 assign wire8004 = ( wire470 ) | ( wire8001 ) ;
 assign wire8005 = ( wire475 ) | ( wire338 ) | ( wire413 ) ;
 assign wire8006 = ( wire1742 ) | ( wire8000 ) | ( n_n1725  &  wire708 ) ;
 assign wire8008 = ( (~ pcount_0_)  &  poutreg_1_ ) | ( pcount_0_  &  poutreg_9_  &  (~ wire577) ) ;
 assign wire8009 = ( (~ pcount_0_)  &  poutreg_25_ ) | ( pcount_0_  &  poutreg_33_  &  (~ wire577) ) ;
 assign wire8010 = ( pdata_59_  &  pcount_0_  &  wire577 ) | ( pcount_0_  &  poutreg_46_  &  (~ wire577) ) ;
 assign wire8013 = ( wire1714 ) | ( wire1716 ) | ( (~ n_n1704)  &  wire712 ) ;
 assign wire8018 = ( wire333 ) | ( (~ n_n1703)  &  (~ wire496)  &  wire319 ) ;
 assign wire8019 = ( wire1698 ) | ( wire1917 ) | ( wire1918 ) | ( wire1919 ) ;
 assign wire8023 = ( wire1691 ) | ( wire1692 ) | ( pc_12_  &  wire254 ) ;
 assign wire8026 = ( wire1687 ) | ( wire1688 ) | ( wire8023 ) ;
 assign wire8028 = ( wire1684 ) | ( wire1685 ) | ( pc_21_  &  wire254 ) ;
 assign wire8031 = ( wire1680 ) | ( wire1681 ) | ( wire8028 ) ;
 assign wire8033 = ( wire1677 ) | ( wire1678 ) | ( pd_11_  &  wire254 ) ;
 assign wire8036 = ( wire1673 ) | ( wire1674 ) | ( wire8033 ) ;
 assign wire8038 = ( wire1670 ) | ( wire1671 ) | ( pd_24_  &  wire254 ) ;
 assign wire8041 = ( wire1666 ) | ( wire1667 ) | ( wire8038 ) ;
 assign wire8047 = ( wire1654 ) | ( n_n1728  &  wire295  &  wire7844 ) ;
 assign wire8048 = ( wire1651 ) | ( wire1652 ) | ( wire1660 ) ;
 assign wire8049 = ( wire1653 ) | ( wire1655 ) | ( wire1656 ) | ( wire1657 ) ;
 assign wire8053 = ( wire338 ) | ( wire1659 ) | ( wire8047 ) | ( wire8048 ) ;
 assign wire8054 = ( wire470 ) | ( wire413 ) | ( wire7852 ) | ( wire8049 ) ;
 assign wire8055 = ( (~ pdata_45_)  &  (~ pdata_44_)  &  pc_6_  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_44_  &  (~ pc_6_)  &  pc_26_ ) | ( pdata_45_  &  (~ pdata_44_)  &  pc_6_  &  (~ pc_26_) ) | ( pdata_45_  &  pdata_44_  &  (~ pc_6_)  &  (~ pc_26_) ) ;
 assign wire8057 = ( pdata_48_  &  (~ pdata_44_)  &  pc_6_  &  pc_1_ ) | ( pdata_48_  &  pdata_44_  &  (~ pc_6_)  &  pc_1_ ) | ( (~ pdata_48_)  &  (~ pdata_44_)  &  pc_6_  &  (~ pc_1_) ) | ( (~ pdata_48_)  &  pdata_44_  &  (~ pc_6_)  &  (~ pc_1_) ) ;
 assign wire8058 = ( wire1630 ) | ( wire286  &  wire301  &  wire8057 ) ;
 assign wire8060 = ( (~ pdata_47_)  &  (~ pdata_44_)  &  pc_12_  &  pc_6_ ) | ( pdata_47_  &  (~ pdata_44_)  &  (~ pc_12_)  &  pc_6_ ) | ( (~ pdata_47_)  &  pdata_44_  &  pc_12_  &  (~ pc_6_) ) | ( pdata_47_  &  pdata_44_  &  (~ pc_12_)  &  (~ pc_6_) ) ;
 assign wire8062 = ( wire1625 ) | ( wire1626 ) | ( wire546  &  wire716 ) ;
 assign wire8063 = ( pdata_47_  &  (~ pdata_46_)  &  pc_12_  &  pc_19_ ) | ( (~ pdata_47_)  &  (~ pdata_46_)  &  (~ pc_12_)  &  pc_19_ ) | ( pdata_47_  &  pdata_46_  &  pc_12_  &  (~ pc_19_) ) | ( (~ pdata_47_)  &  pdata_46_  &  (~ pc_12_)  &  (~ pc_19_) ) ;
 assign wire8066 = ( wire1618 ) | ( wire1617 ) ;
 assign wire8067 = ( pdata_48_  &  pdata_47_  &  pc_12_  &  pc_1_ ) | ( pdata_48_  &  (~ pdata_47_)  &  (~ pc_12_)  &  pc_1_ ) | ( (~ pdata_48_)  &  pdata_47_  &  pc_12_  &  (~ pc_1_) ) | ( (~ pdata_48_)  &  (~ pdata_47_)  &  (~ pc_12_)  &  (~ pc_1_) ) ;
 assign wire8074 = ( wire1602 ) | ( n_n1694  &  wire331  &  wire310 ) ;
 assign wire8075 = ( wire1597 ) | ( wire1598 ) | ( wire1599 ) | ( wire1600 ) ;
 assign wire8077 = ( wire476 ) | ( wire8075 ) ;
 assign wire8078 = ( wire1601 ) | ( wire1619 ) | ( wire8066 ) | ( wire8074 ) ;
 assign wire8080 = ( pdata_47_  &  pcount_0_  &  wire577 ) | ( pcount_0_  &  poutreg_10_  &  (~ wire577) ) ;
 assign wire8081 = ( pcount_0_  &  pdata_44_  &  wire577 ) | ( pcount_0_  &  poutreg_34_  &  (~ wire577) ) ;
 assign wire8084 = ( (~ pdata_45_)  &  (~ pdata_44_)  &  pc_6_  &  pc_26_ ) | ( (~ pdata_45_)  &  pdata_44_  &  (~ pc_6_)  &  pc_26_ ) | ( pdata_45_  &  (~ pdata_44_)  &  pc_6_  &  (~ pc_26_) ) | ( pdata_45_  &  pdata_44_  &  (~ pc_6_)  &  (~ pc_26_) ) ;
 assign wire8088 = ( pdata_48_  &  pdata_46_  &  pc_19_  &  pc_1_ ) | ( pdata_48_  &  (~ pdata_46_)  &  (~ pc_19_)  &  pc_1_ ) | ( (~ pdata_48_)  &  pdata_46_  &  pc_19_  &  (~ pc_1_) ) | ( (~ pdata_48_)  &  (~ pdata_46_)  &  (~ pc_19_)  &  (~ pc_1_) ) ;
 assign wire8089 = ( wire1556 ) | ( wire574  &  wire672 ) ;
 assign wire8091 = ( wire1562 ) | ( wire309  &  wire673 ) ;
 assign wire8092 = ( wire1560 ) | ( wire1561 ) | ( wire8089 ) ;
 assign wire8096 = ( wire468 ) | ( wire476 ) | ( wire1559 ) | ( wire8091 ) ;
 assign wire8097 = ( (~ pcount_0_)  &  poutreg_37_ ) | ( pcount_0_  &  poutreg_45_  &  (~ wire577) ) ;
 assign wire8099 = ( wire1546 ) | ( wire1547 ) | ( pc_13_  &  wire254 ) ;
 assign wire8102 = ( wire1542 ) | ( wire1543 ) | ( wire8099 ) ;
 assign wire8104 = ( wire1539 ) | ( wire1540 ) | ( pc_24_  &  wire254 ) ;
 assign wire8107 = ( wire1535 ) | ( wire1536 ) | ( wire8104 ) ;
 assign wire8109 = ( wire1532 ) | ( wire1533 ) | ( pd_14_  &  wire254 ) ;
 assign wire8112 = ( wire1528 ) | ( wire1529 ) | ( wire8109 ) ;
 assign wire8114 = ( wire1525 ) | ( wire1526 ) | ( pd_21_  &  wire254 ) ;
 assign wire8117 = ( wire1521 ) | ( wire1522 ) | ( wire8114 ) ;
 assign wire8125 = ( pdata_43_  &  pdata_40_  &  pc_18_  &  pc_25_ ) | ( pdata_43_  &  (~ pdata_40_)  &  (~ pc_18_)  &  pc_25_ ) | ( (~ pdata_43_)  &  pdata_40_  &  pc_18_  &  (~ pc_25_) ) | ( (~ pdata_43_)  &  (~ pdata_40_)  &  (~ pc_18_)  &  (~ pc_25_) ) ;
 assign wire8130 = ( wire473 ) | ( wire1494 ) | ( wire1495 ) ;
 assign wire8131 = ( wire1496 ) | ( wire1498 ) | ( n_n1712  &  wire696 ) ;
 assign wire8134 = ( n_n1699  &  n_n1695  &  wire649 ) | ( (~ n_n1699)  &  (~ n_n1695)  &  wire7783 ) ;
 assign wire8138 = ( wire467 ) | ( wire1476 ) | ( wire1477 ) | ( wire1478 ) ;
 assign wire8139 = ( wire471 ) | ( wire2228 ) | ( wire539  &  wire726 ) ;
 assign wire8140 = ( wire336 ) | ( wire1474 ) | ( wire1475 ) ;
 assign wire8143 = ( pdata_36_  &  pdata_40_  &  pc_9_  &  pc_27_ ) | ( pdata_36_  &  (~ pdata_40_)  &  (~ pc_9_)  &  pc_27_ ) | ( (~ pdata_36_)  &  pdata_40_  &  pc_9_  &  (~ pc_27_) ) | ( (~ pdata_36_)  &  (~ pdata_40_)  &  (~ pc_9_)  &  (~ pc_27_) ) ;
 assign wire8144 = ( pdata_35_  &  (~ pdata_37_)  &  pc_14_  &  pc_2_ ) | ( pdata_35_  &  pdata_37_  &  (~ pc_14_)  &  pc_2_ ) | ( (~ pdata_35_)  &  (~ pdata_37_)  &  pc_14_  &  (~ pc_2_) ) | ( (~ pdata_35_)  &  pdata_37_  &  (~ pc_14_)  &  (~ pc_2_) ) ;
 assign wire8150 = ( wire1436 ) | ( wire1434 ) ;
 assign wire8153 = ( wire405 ) | ( wire1429 ) | ( wire1430 ) ;
 assign wire8154 = ( wire1435 ) | ( wire1439 ) | ( wire1440 ) | ( wire8150 ) ;
 assign wire8155 = ( (~ pdata_36_)  &  pdata_40_  &  pc_9_  &  pc_27_ ) | ( (~ pdata_36_)  &  (~ pdata_40_)  &  (~ pc_9_)  &  pc_27_ ) | ( pdata_36_  &  pdata_40_  &  pc_9_  &  (~ pc_27_) ) | ( pdata_36_  &  (~ pdata_40_)  &  (~ pc_9_)  &  (~ pc_27_) ) ;
 assign wire8160 = ( pdata_36_  &  pdata_37_  &  pc_27_  &  pc_14_ ) | ( (~ pdata_36_)  &  pdata_37_  &  (~ pc_27_)  &  pc_14_ ) | ( pdata_36_  &  (~ pdata_37_)  &  pc_27_  &  (~ pc_14_) ) | ( (~ pdata_36_)  &  (~ pdata_37_)  &  (~ pc_27_)  &  (~ pc_14_) ) ;
 assign wire8162 = ( wire1421 ) | ( (~ n_n1684)  &  n_n1687  &  wire523 ) ;
 assign wire8163 = ( wire1418 ) | ( wire1420 ) | ( n_n1686  &  wire639 ) ;
 assign wire8165 = ( wire1412 ) | ( wire1413 ) | ( wire636  &  wire8160 ) ;
 assign wire8166 = ( wire8165 ) | ( wire463 ) ;
 assign wire8168 = ( (~ pcount_0_)  &  poutreg_27_ ) | ( pcount_0_  &  poutreg_35_  &  (~ wire577) ) ;
 assign wire8169 = ( pcount_0_  &  pdata_51_  &  wire577 ) | ( pcount_0_  &  poutreg_44_  &  (~ wire577) ) ;
 assign wire8170 = ( pdata_36_  &  (~ pdata_40_)  &  pc_9_  &  pc_27_ ) | ( pdata_36_  &  pdata_40_  &  (~ pc_9_)  &  pc_27_ ) | ( (~ pdata_36_)  &  (~ pdata_40_)  &  pc_9_  &  (~ pc_27_) ) | ( (~ pdata_36_)  &  pdata_40_  &  (~ pc_9_)  &  (~ pc_27_) ) ;
 assign wire8175 = ( wire1389 ) | ( wire1391 ) | ( wire1392 ) ;
 assign wire8176 = ( wire462 ) | ( pdata_36_  &  pc_27_  &  wire620 ) | ( (~ pdata_36_)  &  (~ pc_27_)  &  wire620 ) ;
 assign wire8178 = ( (~ pcount_0_)  &  poutreg_49_ ) | ( pcount_0_  &  poutreg_57_  &  (~ wire577) ) ;
 assign wire8179 = ( pcount_0_  &  pdata_41_  &  wire577 ) | ( pcount_0_  &  poutreg_58_  &  (~ wire577) ) ;
 assign wire8181 = ( wire1366 ) | ( wire1367 ) | ( pc_14_  &  wire254 ) ;
 assign wire8184 = ( wire1362 ) | ( wire1363 ) | ( wire8181 ) ;
 assign wire8186 = ( wire1359 ) | ( wire1360 ) | ( pc_23_  &  wire254 ) ;
 assign wire8189 = ( wire1355 ) | ( wire1356 ) | ( wire8186 ) ;
 assign wire8191 = ( wire1352 ) | ( wire1353 ) | ( pd_13_  &  wire254 ) ;
 assign wire8194 = ( wire1348 ) | ( wire1349 ) | ( wire8191 ) ;
 assign wire8196 = ( wire1345 ) | ( wire1346 ) | ( pd_22_  &  wire254 ) ;
 assign wire8199 = ( wire1341 ) | ( wire1342 ) | ( wire8196 ) ;
 assign wire8202 = ( (~ pc_22_)  &  pdata_39_  &  wire247 ) | ( pc_22_  &  (~ pdata_39_)  &  wire247 ) ;
 assign wire8204 = ( pdata_43_  &  pdata_41_  &  pc_11_  &  pc_25_ ) | ( pdata_43_  &  (~ pdata_41_)  &  (~ pc_11_)  &  pc_25_ ) | ( (~ pdata_43_)  &  pdata_41_  &  pc_11_  &  (~ pc_25_) ) | ( (~ pdata_43_)  &  (~ pdata_41_)  &  (~ pc_11_)  &  (~ pc_25_) ) ;
 assign wire8206 = ( wire1327 ) | ( (~ n_n1710)  &  wire328  &  wire536 ) ;
 assign wire8207 = ( wire1324 ) | ( wire1326 ) | ( wire630  &  wire8202 ) ;
 assign wire8210 = ( wire398 ) | ( wire1325 ) | ( wire8206 ) | ( wire8207 ) ;
 assign wire8211 = ( pcount_0_  &  pdata_39_  &  wire577 ) | ( pcount_0_  &  poutreg_8_  &  (~ wire577) ) ;
 assign wire8212 = ( pcount_0_  &  pdata_52_  &  wire577 ) | ( pcount_0_  &  poutreg_36_  &  (~ wire577) ) ;
 assign wire8215 = ( (~ pdata_59_)  &  (~ pd_10_)  &  pd_5_  &  pdata_57_ ) | ( pdata_59_  &  (~ pd_10_)  &  (~ pd_5_)  &  pdata_57_ ) | ( (~ pdata_59_)  &  pd_10_  &  pd_5_  &  (~ pdata_57_) ) | ( pdata_59_  &  pd_10_  &  (~ pd_5_)  &  (~ pdata_57_) ) ;
 assign wire8217 = ( (~ n_n1719)  &  (~ n_n1722)  &  wire692 ) | ( (~ n_n1719)  &  n_n1722  &  wire691 ) | ( n_n1719  &  (~ n_n1722)  &  wire691 ) ;
 assign wire8218 = ( wire472 ) | ( n_n1723  &  wire427 ) | ( n_n1723  &  wire1301 ) ;
 assign wire8219 = ( wire335 ) | ( wire1291 ) | ( wire8217 ) ;
 assign wire8221 = ( (~ pcount_0_)  &  poutreg_35_ ) | ( pcount_0_  &  poutreg_43_  &  (~ wire577) ) ;
 assign wire8223 = ( wire1282 ) | ( wire1283 ) | ( pc_15_  &  wire254 ) ;
 assign wire8226 = ( wire1278 ) | ( wire1279 ) | ( wire8223 ) ;
 assign wire8228 = ( wire1275 ) | ( wire1276 ) | ( pc_26_  &  wire254 ) ;
 assign wire8231 = ( wire1271 ) | ( wire1272 ) | ( wire8228 ) ;
 assign wire8233 = ( wire1268 ) | ( wire1269 ) | ( pd_16_  &  wire254 ) ;
 assign wire8236 = ( wire1264 ) | ( wire1265 ) | ( wire8233 ) ;
 assign wire8238 = ( wire1261 ) | ( wire1262 ) | ( pd_27_  &  wire254 ) ;
 assign wire8241 = ( wire1257 ) | ( wire1258 ) | ( wire8238 ) ;
 assign wire8245 = ( pdata_35_  &  pdata_37_  &  pc_14_  &  pc_2_ ) | ( pdata_35_  &  (~ pdata_37_)  &  (~ pc_14_)  &  pc_2_ ) | ( (~ pdata_35_)  &  pdata_37_  &  pc_14_  &  (~ pc_2_) ) | ( (~ pdata_35_)  &  (~ pdata_37_)  &  (~ pc_14_)  &  (~ pc_2_) ) ;
 assign wire8246 = ( (~ pdata_37_)  &  (~ pc_20_)  &  pc_14_  &  pdata_39_ ) | ( pdata_37_  &  (~ pc_20_)  &  (~ pc_14_)  &  pdata_39_ ) | ( (~ pdata_37_)  &  pc_20_  &  pc_14_  &  (~ pdata_39_) ) | ( pdata_37_  &  pc_20_  &  (~ pc_14_)  &  (~ pdata_39_) ) ;
 assign wire8247 = ( n_n1685  &  wire8246 ) | ( n_n1685  &  wire321  &  wire8245 ) ;
 assign wire8250 = ( wire1242 ) | ( wire1243 ) | ( wire1246 ) ;
 assign wire8253 = ( wire405 ) | ( wire1244 ) | ( wire1245 ) | ( wire8250 ) ;
 assign wire8254 = ( (~ pcount_0_)  &  poutreg_5_ ) | ( pcount_0_  &  poutreg_13_  &  (~ wire577) ) ;
 assign wire8258 = ( wire1216 ) | ( n_n1729  &  (~ wire265)  &  wire295 ) ;
 assign wire8259 = ( wire1220 ) | ( wire588  &  wire700 ) ;
 assign wire8263 = ( wire1221 ) | ( wire1222 ) | ( wire297  &  wire701 ) ;
 assign wire8264 = ( wire475 ) | ( wire338 ) | ( wire8258 ) | ( wire8259 ) ;
 assign wire8265 = ( wire413 ) | ( wire7852 ) | ( wire8263 ) ;
 assign wire8266 = ( (~ pcount_0_)  &  poutreg_29_ ) | ( pcount_0_  &  poutreg_37_  &  (~ wire577) ) ;
 assign wire8267 = ( (~ pcount_0_)  &  poutreg_47_ ) | ( pcount_0_  &  poutreg_55_  &  (~ wire577) ) ;
 assign wire8268 = ( pcount_0_  &  pdata_49_  &  wire577 ) | ( pcount_0_  &  poutreg_60_  &  (~ wire577) ) ;
 assign wire8270 = ( wire1202 ) | ( wire1203 ) | ( pc_16_  &  wire254 ) ;
 assign wire8273 = ( wire1198 ) | ( wire1199 ) | ( wire8270 ) ;
 assign wire8275 = ( wire1195 ) | ( wire1196 ) | ( pc_25_  &  wire254 ) ;
 assign wire8278 = ( wire1191 ) | ( wire1192 ) | ( wire8275 ) ;
 assign wire8280 = ( wire1188 ) | ( wire1189 ) | ( pd_15_  &  wire254 ) ;
 assign wire8283 = ( wire1184 ) | ( wire1185 ) | ( wire8280 ) ;
 assign wire8284 = ( pcount_0_  &  pdata_63_  &  wire577 ) | ( pcount_0_  &  poutreg_14_  &  (~ wire577) ) ;
 assign wire8285 = ( pcount_0_  &  pdata_33_  &  wire577 ) | ( pcount_0_  &  poutreg_56_  &  (~ wire577) ) ;
 assign wire8289 = ( wire1152 ) | ( wire285  &  wire678 ) ;
 assign wire8290 = ( wire1156 ) | ( (~ n_n1693)  &  wire286  &  wire331 ) ;
 assign wire8291 = ( wire409 ) | ( wire432 ) | ( wire263  &  wire677 ) ;
 assign wire8293 = ( wire468 ) | ( wire1617 ) | ( wire1618 ) | ( wire1619 ) ;
 assign wire8294 = ( wire8289 ) | ( wire8290 ) | ( wire8291 ) ;
 assign wire8296 = ( poutreg_51_  &  (~ pcount_0_) ) | ( pcount_0_  &  poutreg_59_  &  (~ wire577) ) ;
 assign wire8298 = ( wire1144 ) | ( wire1145 ) | ( pc_17_  &  wire254 ) ;
 assign wire8301 = ( wire1140 ) | ( wire1141 ) | ( wire8298 ) ;
 assign wire8303 = ( wire1137 ) | ( wire1138 ) | ( pd_18_  &  wire254 ) ;
 assign wire8306 = ( wire1133 ) | ( wire1134 ) | ( wire8303 ) ;
 assign wire8308 = ( wire1130 ) | ( wire1131 ) | ( pd_25_  &  wire254 ) ;
 assign wire8311 = ( wire1126 ) | ( wire1127 ) | ( wire8308 ) ;
 assign wire8312 = ( (~ pcount_0_)  &  poutreg_3_ ) | ( pcount_0_  &  poutreg_11_  &  (~ wire577) ) ;
 assign wire8319 = ( pd_11_  &  (~ pd_4_)  &  pdata_52_  &  pdata_55_ ) | ( (~ pd_11_)  &  (~ pd_4_)  &  (~ pdata_52_)  &  pdata_55_ ) | ( pd_11_  &  pd_4_  &  pdata_52_  &  (~ pdata_55_) ) | ( (~ pd_11_)  &  pd_4_  &  (~ pdata_52_)  &  (~ pdata_55_) ) ;
 assign wire8320 = ( wire305  &  wire313 ) | ( wire274  &  wire8319 ) ;
 assign wire8322 = ( wire1099 ) | ( wire284  &  wire680 ) ;
 assign wire8323 = ( wire379 ) | ( wire1098 ) | ( wire1102 ) ;
 assign wire8326 = ( wire411 ) | ( wire1101 ) | ( wire8322 ) | ( wire8323 ) ;
 assign wire8327 = ( (~ pcount_0_)  &  poutreg_45_ ) | ( poutreg_53_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8328 = ( pcount_0_  &  pdata_57_  &  wire577 ) | ( poutreg_62_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8330 = ( wire1087 ) | ( wire1088 ) | ( pc_18_  &  wire254 ) ;
 assign wire8333 = ( wire1083 ) | ( wire1084 ) | ( wire8330 ) ;
 assign wire8335 = ( wire1080 ) | ( wire1081 ) | ( pc_27_  &  wire254 ) ;
 assign wire8338 = ( wire1076 ) | ( wire1077 ) | ( wire8335 ) ;
 assign wire8340 = ( wire1073 ) | ( wire1074 ) | ( pd_17_  &  wire254 ) ;
 assign wire8343 = ( wire1069 ) | ( wire1070 ) | ( wire8340 ) ;
 assign wire8345 = ( wire1066 ) | ( wire1067 ) | ( pd_26_  &  wire254 ) ;
 assign wire8348 = ( wire1062 ) | ( wire1063 ) | ( wire8345 ) ;
 assign wire8350 = ( pdata_40_  &  pc_20_  &  pc_9_  &  pdata_39_ ) | ( (~ pdata_40_)  &  pc_20_  &  (~ pc_9_)  &  pdata_39_ ) | ( pdata_40_  &  (~ pc_20_)  &  pc_9_  &  (~ pdata_39_) ) | ( (~ pdata_40_)  &  (~ pc_20_)  &  (~ pc_9_)  &  (~ pdata_39_) ) ;
 assign wire8352 = ( wire1056 ) | ( (~ wire268)  &  wire8350 ) ;
 assign wire8353 = ( wire484 ) | ( wire603 ) | ( wire1057 ) ;
 assign wire8355 = ( wire1047 ) | ( wire1050 ) | ( wire606  &  wire664 ) ;
 assign wire8356 = ( wire1439 ) | ( wire1440 ) | ( wire8355 ) ;
 assign wire8358 = ( pcount_0_  &  pdata_55_  &  wire577 ) | ( pcount_0_  &  poutreg_12_  &  (~ wire577) ) ;
 assign wire8359 = ( (~ pcount_0_)  &  poutreg_39_ ) | ( pcount_0_  &  poutreg_47_  &  (~ wire577) ) ;
 assign wire8360 = ( pcount_0_  &  pdata_58_  &  wire577 ) | ( pcount_0_  &  poutreg_54_  &  (~ wire577) ) ;
 assign wire8361 = ( poutreg_53_  &  (~ pcount_0_) ) | ( pcount_0_  &  poutreg_61_  &  (~ wire577) ) ;
 assign wire8362 = ( pcount_0_  &  pdata_60_  &  wire577 ) | ( pcount_0_  &  poutreg_38_  &  (~ wire577) ) ;
 assign wire8364 = ( wire1012 ) | ( wire1973 ) | ( wire505  &  wire750 ) ;
 assign wire8367 = ( pd_11_  &  (~ pd_22_)  &  pdata_53_  &  pdata_52_ ) | ( pd_11_  &  pd_22_  &  (~ pdata_53_)  &  pdata_52_ ) | ( (~ pd_11_)  &  (~ pd_22_)  &  pdata_53_  &  (~ pdata_52_) ) | ( (~ pd_11_)  &  pd_22_  &  (~ pdata_53_)  &  (~ pdata_52_) ) ;
 assign wire8370 = ( wire1002 ) | ( wire245  &  wire683 ) ;
 assign wire8371 = ( wire1000 ) | ( wire1001 ) | ( wire1005 ) ;
 assign wire8374 = ( wire469 ) | ( wire1004 ) | ( wire8370 ) | ( wire8371 ) ;
 assign wire8375 = ( (~ pcount_0_)  &  poutreg_43_ ) | ( poutreg_51_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8376 = ( pcount_0_  &  pdata_50_  &  wire577 ) | ( poutreg_52_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8377 = ( (~ pcount_0_)  &  poutreg_55_ ) | ( poutreg_63_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8378 = ( pdata_44_  &  pdata_43_  &  pc_7_  &  pc_25_ ) | ( (~ pdata_44_)  &  pdata_43_  &  (~ pc_7_)  &  pc_25_ ) | ( pdata_44_  &  (~ pdata_43_)  &  pc_7_  &  (~ pc_25_) ) | ( (~ pdata_44_)  &  (~ pdata_43_)  &  (~ pc_7_)  &  (~ pc_25_) ) ;
 assign wire8382 = ( wire977 ) | ( (~ n_n1710)  &  wire526  &  wire7948 ) ;
 assign wire8383 = ( wire431 ) | ( wire976 ) | ( wire312  &  wire653 ) ;
 assign wire8385 = ( wire1836 ) | ( wire7946 ) | ( wire8382 ) | ( wire8383 ) ;
 assign wire8389 = ( (~ pdata_48_)  &  (~ pdata_47_)  &  pd_12_  &  pd_23_ ) | ( (~ pdata_48_)  &  pdata_47_  &  (~ pd_12_)  &  pd_23_ ) | ( pdata_48_  &  (~ pdata_47_)  &  pd_12_  &  (~ pd_23_) ) | ( pdata_48_  &  pdata_47_  &  (~ pd_12_)  &  (~ pd_23_) ) ;
 assign wire8393 = ( wire336 ) | ( wire954 ) | ( wire955 ) | ( wire958 ) ;
 assign wire8396 = ( wire471 ) | ( wire956 ) | ( wire957 ) ;
 assign wire8397 = ( (~ pcount_0_)  &  poutreg_41_ ) | ( pcount_0_  &  poutreg_49_  &  (~ wire577) ) ;
 assign wire8400 = ( pdata_33_  &  pc_10_  &  wire264 ) | ( (~ pdata_33_)  &  (~ pc_10_)  &  wire264 ) ;
 assign wire8402 = ( wire934 ) | ( wire935 ) | ( wire325  &  wire8400 ) ;
 assign wire8403 = ( wire1917 ) | ( wire1918 ) | ( wire1919 ) | ( wire8402 ) ;
 assign wire8404 = ( wire937 ) | ( wire465 ) ;
 assign wire8406 = ( pcount_0_  &  pdata_53_  &  wire577 ) | ( pcount_0_  &  poutreg_28_  &  (~ wire577) ) ;
 assign wire8407 = ( pcount_0_  &  pdata_42_  &  wire577 ) | ( pcount_0_  &  poutreg_50_  &  (~ wire577) ) ;
 assign wire8413 = ( wire433 ) | ( wire904 ) | ( wire909 ) ;
 assign wire8414 = ( wire905 ) | ( wire908 ) | ( wire285  &  wire688 ) ;
 assign wire8416 = ( wire476 ) | ( wire468 ) ;
 assign wire8417 = ( wire1619 ) | ( wire1631 ) | ( wire8058 ) | ( wire8066 ) ;
 assign wire8418 = ( wire8413 ) | ( wire8414 ) | ( wire286  &  wire689 ) ;
 assign wire8420 = ( (~ pdata_36_)  &  (~ pdata_34_)  &  pc_23_  &  pc_4_ ) | ( (~ pdata_36_)  &  pdata_34_  &  (~ pc_23_)  &  pc_4_ ) | ( pdata_36_  &  (~ pdata_34_)  &  pc_23_  &  (~ pc_4_) ) | ( pdata_36_  &  pdata_34_  &  (~ pc_23_)  &  (~ pc_4_) ) ;
 assign wire8421 = ( (~ pdata_36_)  &  (~ pc_13_)  &  pc_4_  &  pdata_63_ ) | ( pdata_36_  &  (~ pc_13_)  &  (~ pc_4_)  &  pdata_63_ ) | ( (~ pdata_36_)  &  pc_13_  &  pc_4_  &  (~ pdata_63_) ) | ( pdata_36_  &  pc_13_  &  (~ pc_4_)  &  (~ pdata_63_) ) ;
 assign wire8423 = ( wire592  &  wire319 ) | ( pdata_34_  &  pc_23_  &  wire319 ) | ( (~ pdata_34_)  &  (~ pc_23_)  &  wire319 ) ;
 assign wire8424 = ( (~ pdata_32_)  &  (~ pdata_34_)  &  pc_16_  &  pc_23_ ) | ( pdata_32_  &  (~ pdata_34_)  &  (~ pc_16_)  &  pc_23_ ) | ( (~ pdata_32_)  &  pdata_34_  &  pc_16_  &  (~ pc_23_) ) | ( pdata_32_  &  pdata_34_  &  (~ pc_16_)  &  (~ pc_23_) ) ;
 assign wire8428 = ( wire465 ) | ( (~ n_n1704)  &  wire889 ) | ( (~ n_n1704)  &  wire8423 ) ;
 assign wire8429 = ( wire333 ) | ( wire883 ) | ( n_n1704  &  wire662 ) ;
 assign wire8432 = ( pdata_59_  &  pdata_60_  &  pd_24_  &  pd_5_ ) | ( pdata_59_  &  (~ pdata_60_)  &  (~ pd_24_)  &  pd_5_ ) | ( (~ pdata_59_)  &  pdata_60_  &  pd_24_  &  (~ pd_5_) ) | ( (~ pdata_59_)  &  (~ pdata_60_)  &  (~ pd_24_)  &  (~ pd_5_) ) ;
 assign wire8433 = ( pd_10_  &  (~ pdata_60_)  &  pd_24_  &  pdata_57_ ) | ( pd_10_  &  pdata_60_  &  (~ pd_24_)  &  pdata_57_ ) | ( (~ pd_10_)  &  (~ pdata_60_)  &  pd_24_  &  (~ pdata_57_) ) | ( (~ pd_10_)  &  pdata_60_  &  (~ pd_24_)  &  (~ pdata_57_) ) ;
 assign wire8435 = ( (~ pd_27_)  &  pdata_58_  &  wire529 ) | ( pd_27_  &  (~ pdata_58_)  &  wire529 ) ;
 assign wire8437 = ( wire866 ) | ( wire863 ) ;
 assign wire8439 = ( wire862 ) | ( wire246  &  wire709 ) | ( (~ wire246)  &  wire8435 ) ;
 assign wire8440 = ( wire2293 ) | ( wire8437 ) | ( wire747  &  wire7729 ) ;
 assign wire8441 = ( wire335 ) | ( wire8439 ) | ( wire710  &  wire8432 ) ;
 assign wire8443 = ( (~ pcount_0_)  &  poutreg_21_ ) | ( pcount_0_  &  poutreg_29_  &  (~ wire577) ) ;
 assign wire8444 = ( pcount_0_  &  pdata_43_  &  wire577 ) | ( pcount_0_  &  poutreg_42_  &  (~ wire577) ) ;
 assign wire8446 = ( wire850 ) | ( wire851 ) | ( pd_20_  &  wire254 ) ;
 assign wire8449 = ( wire846 ) | ( wire847 ) | ( wire8446 ) ;
 assign wire8457 = ( wire824 ) | ( wire825 ) | ( wire827 ) | ( wire828 ) ;
 assign wire8459 = ( wire477 ) | ( wire8457 ) | ( (~ n_n1716)  &  wire705 ) ;
 assign wire8460 = ( pcount_0_  &  pdata_61_  &  wire577 ) | ( pcount_0_  &  poutreg_30_  &  (~ wire577) ) ;
 assign wire8461 = ( (~ pcount_0_)  &  poutreg_33_ ) | ( pcount_0_  &  poutreg_41_  &  (~ wire577) ) ;
 assign wire8462 = ( pcount_0_  &  pdata_34_  &  wire577 ) | ( pcount_0_  &  poutreg_48_  &  (~ wire577) ) ;
 assign wire8464 = ( wire802 ) | ( wire803 ) | ( pc_20_  &  wire254 ) ;
 assign wire8467 = ( wire798 ) | ( wire799 ) | ( wire8464 ) ;
 assign wire8469 = ( wire795 ) | ( wire796 ) | ( pd_10_  &  wire254 ) ;
 assign wire8472 = ( wire791 ) | ( wire792 ) | ( wire8469 ) ;
 assign wire8473 = ( (~ pcount_0_)  &  poutreg_23_ ) | ( pcount_0_  &  poutreg_31_  &  (~ wire577) ) ;
 assign wire8474 = ( pdata_35_  &  pcount_0_  &  wire577 ) | ( poutreg_40_  &  pcount_0_  &  (~ wire577) ) ;
 assign wire8476 = ( wire774 ) | ( wire775 ) | ( pc_10_  &  wire254 ) ;
 assign wire8479 = ( wire770 ) | ( wire771 ) | ( wire8476 ) ;
 assign wire8480 = ( pdata_36_  &  pcount_0_  &  wire577 ) | ( pcount_0_  &  poutreg_32_  &  (~ wire577) ) ;
 assign wire8481 = ( (~ pcount_0_)  &  poutreg_31_ ) | ( pcount_0_  &  poutreg_39_  &  (~ wire577) ) ;
 assign wire8482 = ( pcount_0_  &  pdata_54_  &  wire577 ) | ( pcount_0_  &  poutreg_20_  &  (~ wire577) ) ;
 assign wire8483 = ( (~ pcount_0_)  &  poutreg_11_ ) | ( pcount_0_  &  poutreg_19_  &  (~ wire577) ) ;
 assign wire8484 = ( pcount_0_  &  pdata_62_  &  wire577 ) | ( pcount_0_  &  poutreg_22_  &  (~ wire577) ) ;
 assign wire8485 = ( (~ pcount_0_)  &  poutreg_13_ ) | ( pcount_0_  &  poutreg_21_  &  (~ wire577) ) ;
 assign wire8487 = ( wire455 ) | ( wire456 ) | ( pd_9_  &  wire254 ) ;
 assign wire8490 = ( wire451 ) | ( wire452 ) | ( wire8487 ) ;
 assign wire8492 = ( wire435 ) | ( wire436 ) | ( pc_8_  &  wire254 ) ;
 assign wire8495 = ( wire422 ) | ( wire425 ) | ( wire8492 ) ;
 assign wire8497 = ( wire418 ) | ( wire419 ) | ( pd_7_  &  wire254 ) ;
 assign wire8500 = ( wire404 ) | ( wire414 ) | ( wire8497 ) ;
 assign wire8501 = ( pdata_46_  &  pcount_0_  &  wire577 ) | ( pcount_0_  &  poutreg_18_  &  (~ wire577) ) ;
 assign wire8503 = ( wire383 ) | ( wire384 ) | ( pc_9_  &  wire254 ) ;
 assign wire8506 = ( wire376 ) | ( wire377 ) | ( wire8503 ) ;
 assign wire8508 = ( wire339 ) | ( wire374 ) | ( pd_8_  &  wire254 ) ;
 assign wire8511 = ( wire327 ) | ( wire329 ) | ( wire8508 ) ;


endmodule

