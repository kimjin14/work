module s38417 (
	pg1943, pg1249, pg3219, pg3229, pg3217, pg3228, pg3218, pg3227, 
	pg2637, pg3222, pg3233, pg3212, pg3221, pg3234, pclk, pg3220, pg3215, pg3226, 
	pg3216, pg3225, pg3230, pg3213, pg3224, pg3231, pg3214, pg3223, pg3232, pg51, 
	pg563, pg8012, pg8023, pg8265, pg16297, pg8167, pg8266, pg8275, pg4090, pg7161, 
	pg7194, pg8021, pg8175, pg8263, pg8274, pg7052, pg8264, pg8273, pg7390, pg8261, 
	pg8272, pg8262, pg8271, pg16355, pg24734, pg6573, pg7084, pg7264, pg7334, pg8007, 
	pg8106, pg8270, pg8251, pg8260, pg4590, pg6642, pg6750, pg7302, pg4450, pg6225, 
	pg26135, pg4088, pg5472, pg6442, pg8030, pg16437, pg25435, pg5511, pg7014, pg16399, 
	pg16496, pg27380, pg6313, pg5612, pg6231, pg26149, pg5437, pg5657, pg6979, pg25420, 
	pg25442, pg3993, pg6911, pg6944, pg4323, pg6712, pg6837, pg7519, pg25489, pg5686, 
	pg5738, pg6447, pg26104, pg4200, pg4321, pg5388, pg5555, pg7229, pg5549, pg5637, 
	pg5648, pg5747, pg5629, pg6518, pg7425, pg5595, pg8082, pg5695, pg6368, pg6485, 
	pg6782, pg7961, pg7357, pg5796, pg7909, pg7956, pg8096, pg8258, pg8269, pg6677, 
	pg8087, pg8249, pg8267, pg6895, pg7487, pg8259, pg8268);

input pg1943;
input pg1249;
input pg3219;
input pg3229;
input pg3217;
input pg3228;
input pg3218;
input pg3227;
input pg2637;
input pg3222;
input pg3233;
input pg3212;
input pg3221;
input pg3234;
input pclk;
input pg3220;
input pg3215;
input pg3226;
input pg3216;
input pg3225;
input pg3230;
input pg3213;
input pg3224;
input pg3231;
input pg3214;
input pg3223;
input pg3232;
input pg51;
input pg563;
output pg8012;
output pg8023;
output pg8265;
output pg16297;
output pg8167;
output pg8266;
output pg8275;
output pg4090;
output pg7161;
output pg7194;
output pg8021;
output pg8175;
output pg8263;
output pg8274;
output pg7052;
output pg8264;
output pg8273;
output pg7390;
output pg8261;
output pg8272;
output pg8262;
output pg8271;
output pg16355;
output pg24734;
output pg6573;
output pg7084;
output pg7264;
output pg7334;
output pg8007;
output pg8106;
output pg8270;
output pg8251;
output pg8260;
output pg4590;
output pg6642;
output pg6750;
output pg7302;
output pg4450;
output pg6225;
output pg26135;
output pg4088;
output pg5472;
output pg6442;
output pg8030;
output pg16437;
output pg25435;
output pg5511;
output pg7014;
output pg16399;
output pg16496;
output pg27380;
output pg6313;
output pg5612;
output pg6231;
output pg26149;
output pg5437;
output pg5657;
output pg6979;
output pg25420;
output pg25442;
output pg3993;
output pg6911;
output pg6944;
output pg4323;
output pg6712;
output pg6837;
output pg7519;
output pg25489;
output pg5686;
output pg5738;
output pg6447;
output pg26104;
output pg4200;
output pg4321;
output pg5388;
output pg5555;
output pg7229;
output pg5549;
output pg5637;
output pg5648;
output pg5747;
output pg5629;
output pg6518;
output pg7425;
output pg5595;
output pg8082;
output pg5695;
output pg6368;
output pg6485;
output pg6782;
output pg7961;
output pg7357;
output pg5796;
output pg7909;
output pg7956;
output pg8096;
output pg8258;
output pg8269;
output pg6677;
output pg8087;
output pg8249;
output pg8267;
output pg6895;
output pg7487;
output pg8259;
output pg8268;
wire ng25450;
wire ng30801;
wire ng17341;
wire ng22030;
wire ng22064;
wire ng30258;
wire ng26529;
wire ng27256;
wire ng28744;
wire ng26808;
wire ng30455;
wire ng11510;
wire ng18678;
wire ng24174;
wire ng27279;
wire ng24498;
wire ng26541;
wire ng24426;
wire ng20892;
wire ng20946;
wire ng21051;
wire ng25262;
wire ng22146;
wire ng22066;
wire ng22128;
wire ng25223;
wire ng30654;
wire ng30264;
wire ng30670;
wire ng29354;
wire ng27284;
wire ng28767;
wire ng29612;
wire ng26661;
wire ng11519;
wire ng26183;
wire ng23081;
wire ng23039;
wire ng27328;
wire ng28355;
wire ng26781;
wire ng20926;
wire ng20995;
wire ng20913;
wire ng22247;
wire ng22044;
wire ng22130;
wire ng25224;
wire ng30281;
wire ng27129;
wire ng27288;
wire ng29205;
wire ng26824;
wire ng30503;
wire ng18794;
wire ng24208;
wire ng27306;
wire ng24534;
wire ng28361;
wire ng13445;
wire ng23339;
wire ng20916;
wire ng21019;
wire ng21072;
wire ng22172;
wire ng25247;
wire ng30672;
wire ng30282;
wire ng30686;
wire ng29357;
wire ng27322;
wire ng29221;
wire ng27767;
wire ng18780;
wire ng24209;
wire ng27336;
wire ng20962;
wire ng21026;
wire ng21075;
wire ng21063;
wire ng29454;
wire ng25451;
wire ng30798;
wire ng17429;
wire ng22028;
wire ng22049;
wire ng30263;
wire ng25932;
wire ng27259;
wire ng28735;
wire ng26812;
wire ng30702;
wire ng11494;
wire ng21842;
wire ng23399;
wire ng27268;
wire ng24507;
wire ng28348;
wire ng25185;
wire ng20880;
wire ng20967;
wire ng21032;
wire ng25266;
wire ng22162;
wire ng22056;
wire ng22106;
wire ng30648;
wire ng30676;
wire ng30259;
wire ng30677;
wire ng29110;
wire ng27298;
wire ng28759;
wire ng29616;
wire ng29179;
wire ng19024;
wire ng26120;
wire ng23111;
wire ng23014;
wire ng13171;
wire ng27315;
wire ng28360;
wire ng26272;
wire ng27678;
wire ng20912;
wire ng21016;
wire ng20898;
wire ng22263;
wire ng22057;
wire ng22114;
wire ng25217;
wire ng30295;
wire ng27612;
wire ng27275;
wire ng29212;
wire ng26821;
wire ng30338;
wire ng11564;
wire ng12524;
wire ng24219;
wire ng27320;
wire ng24524;
wire ng26559;
wire ng13444;
wire ng24434;
wire ng20934;
wire ng21001;
wire ng21056;
wire ng22184;
wire ng25251;
wire ng30690;
wire ng30274;
wire ng30691;
wire ng29112;
wire ng27309;
wire ng29213;
wire ng30341;
wire ng11576;
wire ng21847;
wire ng23418;
wire ng27325;
wire ng23348;
wire ng21043;
wire ng21081;
wire ng25272;
wire ng29453;
wire ng25452;
wire ng17247;
wire ng17383;
wire ng22125;
wire ng25220;
wire ng30268;
wire ng27594;
wire ng27255;
wire ng28732;
wire ng27759;
wire ng11509;
wire ng12487;
wire ng23385;
wire ng13149;
wire ng27280;
wire ng27327;
wire ng28344;
wire ng26660;
wire ng20893;
wire ng20945;
wire ng21011;
wire ng22218;
wire ng22177;
wire ng22042;
wire ng22127;
wire ng30681;
wire ng30247;
wire ng30642;
wire ng28635;
wire ng27313;
wire ng26809;
wire ng27765;
wire ng29173;
wire ng23126;
wire ng24222;
wire ng26534;
wire ng27301;
wire ng28346;
wire ng13427;
wire ng21033;
wire ng20975;
wire ng25270;
wire ng22043;
wire ng22131;
wire ng25225;
wire ng30294;
wire ng28147;
wire ng27289;
wire ng28760;
wire ng26816;
wire ng29178;
wire ng23413;
wire ng12482;
wire ng27331;
wire ng24535;
wire ng26573;
wire ng13447;
wire ng20752;
wire ng20915;
wire ng21023;
wire ng22183;
wire ng22173;
wire ng25256;
wire ng30660;
wire ng30304;
wire ng30694;
wire ng13110;
wire ng27292;
wire ng28782;
wire ng30356;
wire ng11592;
wire ng12539;
wire ng23407;
wire ng13175;
wire ng27337;
wire ng24438;
wire ng20963;
wire ng21074;
wire ng25280;
wire ng29456;
wire ng28420;
wire ng17229;
wire ng17271;
wire ng22143;
wire ng25228;
wire ng30635;
wire ng27120;
wire ng27258;
wire ng27293;
wire ng30468;
wire ng11493;
wire ng18726;
wire ng23117;
wire ng27269;
wire ng24491;
wire ng28342;
wire ng26776;
wire ng20901;
wire ng20966;
wire ng21031;
wire ng22231;
wire ng22163;
wire ng22055;
wire ng22105;
wire ng30687;
wire ng30270;
wire ng30647;
wire ng28146;
wire ng28738;
wire ng26806;
wire ng29609;
wire ng29170;
wire ng23392;
wire ng24212;
wire ng13124;
wire ng27314;
wire ng13426;
wire ng13428;
wire ng21017;
wire ng20952;
wire ng22234;
wire ng22035;
wire ng22150;
wire ng25233;
wire ng25234;
wire ng28636;
wire ng27302;
wire ng28771;
wire ng26820;
wire ng29181;
wire ng11565;
wire ng24182;
wire ng24243;
wire ng27321;
wire ng24525;
wire ng26592;
wire ng13446;
wire ng21972;
wire ng20899;
wire ng21042;
wire ng22192;
wire ng22185;
wire ng25252;
wire ng30666;
wire ng30303;
wire ng25067;
wire ng29582;
wire ng27308;
wire ng28773;
wire ng29182;
wire ng18820;
wire ng21970;
wire ng27326;
wire ng25197;
wire ng20940;
wire ng21006;
wire ng25288;
wire ng29455;
wire ng26037;
wire ng17246;
wire ng29939;
wire ng17248;
wire ng28313;
wire ng30668;
wire ng30262;
wire ng30669;
wire ng29579;
wire ng27278;
wire ng26106;
wire ng23093;
wire ng13410;
wire ng20314;
wire ng21010;
wire ng22242;
wire ng25221;
wire ng30277;
wire ng28746;
wire ng26810;
wire ng11538;
wire ng23406;
wire ng12467;
wire ng27285;
wire ng24511;
wire ng26569;
wire ng21034;
wire ng20976;
wire ng22178;
wire ng22074;
wire ng22091;
wire ng22152;
wire ng29111;
wire ng27317;
wire ng28772;
wire ng29613;
wire ng30704;
wire ng26675;
wire ng23030;
wire ng13135;
wire ng27341;
wire ng13449;
wire ng20978;
wire ng21041;
wire ng21022;
wire ng22182;
wire ng22194;
wire ng25257;
wire ng30667;
wire ng30260;
wire ng30297;
wire ng27621;
wire ng27291;
wire ng28763;
wire ng29185;
wire ng11572;
wire ng23133;
wire ng24538;
wire ng26616;
wire ng13464;
wire ng22269;
wire ng29458;
wire ng17226;
wire ng29936;
wire ng17303;
wire ng30674;
wire ng30257;
wire ng30245;
wire ng27253;
wire ng27267;
wire ng23067;
wire ng13411;
wire ng16654;
wire ng20923;
wire ng22029;
wire ng25215;
wire ng30269;
wire ng28758;
wire ng26813;
wire ng11522;
wire ng24179;
wire ng24235;
wire ng27339;
wire ng24522;
wire ng26557;
wire ng21052;
wire ng20996;
wire ng22167;
wire ng22059;
wire ng22112;
wire ng22168;
wire ng29355;
wire ng27303;
wire ng28778;
wire ng27768;
wire ng30706;
wire ng26670;
wire ng23058;
wire ng29113;
wire ng27290;
wire ng27333;
wire ng22651;
wire ng13448;
wire ng20999;
wire ng21054;
wire ng21003;
wire ng22170;
wire ng25227;
wire ng25253;
wire ng30673;
wire ng30256;
wire ng30652;
wire ng27131;
wire ng27307;
wire ng27342;
wire ng29187;
wire ng19048;
wire ng23114;
wire ng27343;
wire ng13463;
wire ng22284;
wire ng29457;
wire ng17235;
wire ng30796;
wire ng17270;
wire ng28696;
wire ng30246;
wire ng25027;
wire ng27277;
wire ng13412;
wire ng23136;
wire ng20891;
wire ng22067;
wire ng25222;
wire ng30643;
wire ng30701;
wire ng26669;
wire ng11518;
wire ng24181;
wire ng27329;
wire ng24532;
wire ng22615;
wire ng21035;
wire ng21018;
wire ng22149;
wire ng22073;
wire ng22092;
wire ng22180;
wire ng29581;
wire ng27318;
wire ng29218;
wire ng27766;
wire ng30708;
wire ng23124;
wire ng24231;
wire ng27305;
wire ng24513;
wire ng25194;
wire ng20953;
wire ng20979;
wire ng21071;
wire ng20980;
wire ng22280;
wire ng25236;
wire ng30289;
wire ng30693;
wire ng30253;
wire ng30659;
wire ng28637;
wire ng27335;
wire ng26672;
wire ng11573;
wire ng27338;
wire ng24557;
wire ng13462;
wire ng22299;
wire ng17269;
wire ng29941;
wire ng17340;
wire ng30248;
wire ng30675;
wire ng29353;
wire ng13413;
wire ng20682;
wire ng23324;
wire ng22147;
wire ng25230;
wire ng30285;
wire ng30703;
wire ng26665;
wire ng27273;
wire ng27316;
wire ng28351;
wire ng21053;
wire ng20997;
wire ng22166;
wire ng22058;
wire ng22113;
wire ng22169;
wire ng27264;
wire ng27304;
wire ng28761;
wire ng27764;
wire ng30487;
wire ng11563;
wire ng23097;
wire ng23123;
wire ng13164;
wire ng27319;
wire ng27346;
wire ng26671;
wire ng20935;
wire ng21000;
wire ng21055;
wire ng21002;
wire ng22267;
wire ng25245;
wire ng25259;
wire ng30695;
wire ng30290;
wire ng30665;
wire ng28148;
wire ng27276;
wire ng27324;
wire ng26676;
wire ng27344;
wire ng24548;
wire ng26596;
wire ng29459;
wire ng22026;
wire ng22100;
wire ng22037;
wire ng22080;
wire ng25207;
wire ng30275;
wire ng30284;
wire ng27760;
wire ng29167;
wire ng27294;
wire ng24508;
wire ng13417;
wire ng20879;
wire ng22087;
wire ng22148;
wire ng25232;
wire ng30293;
wire ng30638;
wire ng11536;
wire ng28350;
wire ng13433;
wire ng24430;
wire ng20911;
wire ng20974;
wire ng25244;
wire ng30692;
wire ng30252;
wire ng25056;
wire ng22076;
wire ng22139;
wire ng25237;
wire ng28783;
wire ng29618;
wire ng26025;
wire ng11574;
wire ng27347;
wire ng28368;
wire ng16718;
wire ng28328;
wire ng21005;
wire ng21062;
wire ng29460;
wire ng30908;
wire ng30982;
wire ng25191;
wire ng16844;
wire ng16854;
wire ng23358;
wire ng22122;
wire ng22031;
wire ng22101;
wire ng25211;
wire ng30637;
wire ng30276;
wire ng28736;
wire ng29169;
wire ng11511;
wire ng27281;
wire ng24499;
wire ng22578;
wire ng13416;
wire ng20944;
wire ng22033;
wire ng22164;
wire ng25240;
wire ng30298;
wire ng30278;
wire ng11520;
wire ng24501;
wire ng24072;
wire ng23329;
wire ng20925;
wire ng20993;
wire ng25250;
wire ng30688;
wire ng30255;
wire ng30689;
wire ng11548;
wire ng22061;
wire ng22117;
wire ng30296;
wire ng28788;
wire ng27771;
wire ng11590;
wire ng27345;
wire ng28364;
wire ng13458;
wire ng13466;
wire ng20918;
wire ng20983;
wire ng21028;
wire ng29655;
wire ng30119;
wire ng30983;
wire ng24445;
wire ng16853;
wire ng16845;
wire ng24473;
wire ng22141;
wire ng22038;
wire ng22079;
wire ng25206;
wire ng30640;
wire ng30254;
wire ng28745;
wire ng29606;
wire ng19012;
wire ng23000;
wire ng13111;
wire ng21435;
wire ng13418;
wire ng20991;
wire ng25209;
wire ng25248;
wire ng27123;
wire ng27271;
wire ng11537;
wire ng18763;
wire ng24510;
wire ng26547;
wire ng13434;
wire ng26666;
wire ng20910;
wire ng20973;
wire ng22090;
wire ng22151;
wire ng25255;
wire ng30664;
wire ng30280;
wire ng30684;
wire ng26667;
wire ng22077;
wire ng22140;
wire ng30679;
wire ng26817;
wire ng29623;
wire ng11575;
wire ng30055;
wire ng23047;
wire ng13143;
wire ng27348;
wire ng28358;
wire ng22687;
wire ng24092;
wire ng20939;
wire ng21061;
wire ng21007;
wire ng29972;
wire ng30910;
wire ng30980;
wire ng23330;
wire ng16860;
wire ng16880;
wire ng18542;
wire ng25201;
wire ng22123;
wire ng22032;
wire ng22065;
wire ng25204;
wire ng30645;
wire ng30292;
wire ng28754;
wire ng27762;
wire ng30482;
wire ng21346;
wire ng23022;
wire ng21851;
wire ng24059;
wire ng20947;
wire ng20969;
wire ng25214;
wire ng25241;
wire ng27603;
wire ng27263;
wire ng11521;
wire ng12507;
wire ng24521;
wire ng28354;
wire ng25189;
wire ng20897;
wire ng20951;
wire ng22075;
wire ng22132;
wire ng30279;
wire ng30658;
wire ng30250;
wire ng30678;
wire ng29620;
wire ng11549;
wire ng22097;
wire ng22153;
wire ng30283;
wire ng26822;
wire ng29621;
wire ng11591;
wire ng26144;
wire ng23076;
wire ng30072;
wire ng27354;
wire ng28371;
wire ng30061;
wire ng13465;
wire ng21025;
wire ng21073;
wire ng20965;
wire ng29973;
wire ng30909;
wire ng30981;
wire ng26048;
wire ng16803;
wire ng16861;
wire ng16802;
wire ng28421;
wire ng17236;
wire ng22142;
wire ng22039;
wire ng22124;
wire ng25219;
wire ng25229;
wire ng30641;
wire ng30636;
wire ng28634;
wire ng27266;
wire ng26803;
wire ng29611;
wire ng26659;
wire ng23092;
wire ng24206;
wire ng13160;
wire ng27296;
wire ng28353;
wire ng27672;
wire ng20921;
wire ng20990;
wire ng20924;
wire ng20948;
wire ng22041;
wire ng22089;
wire ng30649;
wire ng30251;
wire ng25935;
wire ng27270;
wire ng27282;
wire ng29204;
wire ng27761;
wire ng30500;
wire ng21843;
wire ng24213;
wire ng13155;
wire ng27300;
wire ng13429;
wire ng20333;
wire ng20882;
wire ng20972;
wire ng25263;
wire ng22191;
wire ng25242;
wire ng30657;
wire ng30266;
wire ng30656;
wire ng26815;
wire ng19036;
wire ng22078;
wire ng22171;
wire ng25940;
wire ng26825;
wire ng30709;
wire ng23132;
wire ng24225;
wire ng13194;
wire ng24527;
wire ng28367;
wire ng13461;
wire ng26677;
wire ng20964;
wire ng21060;
wire ng20941;
wire ng20877;
wire ng29974;
wire ng30912;
wire ng30986;
wire ng23359;
wire ng16866;
wire ng18907;
wire ng16823;
wire ng28425;
wire ng17302;
wire ng22161;
wire ng22047;
wire ng22103;
wire ng25213;
wire ng25239;
wire ng30680;
wire ng30639;
wire ng28145;
wire ng29201;
wire ng26804;
wire ng29608;
wire ng26664;
wire ng11492;
wire ng24216;
wire ng24215;
wire ng27312;
wire ng28349;
wire ng28199;
wire ng20902;
wire ng21009;
wire ng20894;
wire ng20970;
wire ng22054;
wire ng22104;
wire ng30655;
wire ng30249;
wire ng26530;
wire ng27262;
wire ng27272;
wire ng29198;
wire ng27763;
wire ng30485;
wire ng18707;
wire ng27286;
wire ng13430;
wire ng16671;
wire ng20896;
wire ng20950;
wire ng25267;
wire ng22179;
wire ng25235;
wire ng30651;
wire ng30272;
wire ng30650;
wire ng28749;
wire ng11546;
wire ng22098;
wire ng22154;
wire ng26823;
wire ng30707;
wire ng24238;
wire ng24237;
wire ng24537;
wire ng28363;
wire ng21974;
wire ng26795;
wire ng20981;
wire ng21045;
wire ng20919;
wire ng21046;
wire ng29975;
wire ng30911;
wire ng30987;
wire ng22002;
wire ng16857;
wire ng21964;
wire ng19152;
wire ng29656;
wire ng22025;
wire ng22063;
wire ng22081;
wire ng25218;
wire ng30261;
wire ng30653;
wire ng30661;
wire ng27265;
wire ng29197;
wire ng26807;
wire ng30700;
wire ng29172;
wire ng11495;
wire ng24207;
wire ng24228;
wire ng27261;
wire ng27295;
wire ng28345;
wire ng26545;
wire ng13415;
wire ng28668;
wire ng20922;
wire ng20989;
wire ng20881;
wire ng20992;
wire ng22145;
wire ng22040;
wire ng22088;
wire ng25231;
wire ng30662;
wire ng30271;
wire ng30682;
wire ng27257;
wire ng27283;
wire ng28747;
wire ng26814;
wire ng30470;
wire ng23110;
wire ng27299;
wire ng13431;
wire ng21969;
wire ng27718;
wire ng20927;
wire ng20994;
wire ng20883;
wire ng25243;
wire ng30683;
wire ng30299;
wire ng30644;
wire ng27287;
wire ng26130;
wire ng27323;
wire ng26826;
wire ng30505;
wire ng24226;
wire ng24250;
wire ng27310;
wire ng24547;
wire ng13459;
wire ng20789;
wire ng27243;
wire ng21004;
wire ng21027;
wire ng21094;
wire ng21029;
wire ng20497;
wire ng29976;
wire ng30914;
wire ng30984;
wire ng26786;
wire ng21966;
wire ng18837;
wire ng20825;
wire ng29166;
wire ng22027;
wire ng22048;
wire ng22102;
wire ng25212;
wire ng30267;
wire ng30646;
wire ng29109;
wire ng27260;
wire ng29194;
wire ng26805;
wire ng30699;
wire ng26655;
wire ng11491;
wire ng24178;
wire ng12457;
wire ng27311;
wire ng24519;
wire ng26553;
wire ng13414;
wire ng20875;
wire ng20903;
wire ng20968;
wire ng20876;
wire ng25260;
wire ng22126;
wire ng22034;
wire ng22068;
wire ng22129;
wire ng30286;
wire ng30265;
wire ng25042;
wire ng29580;
wire ng27297;
wire ng29209;
wire ng26818;
wire ng30705;
wire ng24223;
wire ng13432;
wire ng20717;
wire ng28321;
wire ng20949;
wire ng21015;
wire ng21070;
wire ng25249;
wire ng30663;
wire ng30302;
wire ng30288;
wire ng26531;
wire ng11547;
wire ng28903;
wire ng29226;
wire ng26827;
wire ng30566;
wire ng24214;
wire ng12499;
wire ng26575;
wire ng13460;
wire ng20375;
wire ng27724;
wire ng20982;
wire ng21044;
wire ng21082;
wire ng21047;
wire ng20884;
wire ng29977;
wire ng30913;
wire ng30985;
wire ng26031;
wire ng16824;
wire ng16566;
wire ng18868;
wire ng20417;
wire ng18885;
wire ng18782;
wire ng29978;
wire ng30940;
wire ng19173;
wire ng19149;
wire ng17222;
wire ng29979;
wire ng30915;
wire ng21878;
wire ng20874;
wire ng17225;
wire ng30989;
wire ng25202;
wire ng19184;
wire ng19144;
wire ng17234;
wire ng25265;
wire ng24446;
wire ng26798;
wire ng18852;
wire ng17224;
wire ng30287;
wire ng22193;
wire ng22099;
wire ng16835;
wire ng18804;
wire ng21989;
wire ng18835;
wire ng17228;
wire ng30671;
wire ng22200;
wire ng22115;
wire ng16851;
wire ng18755;
wire ng23357;
wire ng18821;
wire ng30273;
wire ng18743;
wire ng22045;
wire ng22138;
wire ng27769;
wire ng24476;
wire ng18803;
wire ng25938;
wire ng21845;
wire ng22060;
wire ng22116;
wire ng28774;
wire ng25199;
wire ng19154;
wire ng19172;
wire ng27274;
wire ng23400;
wire ng20936;
wire ng21039;
wire ng20917;
wire ng22249;
wire ng27334;
wire ng16181;
wire ng21880;
wire ng20376;
wire ng27330;
wire ng23137;
wire ng20954;
wire ng21020;
wire ng20937;
wire ng25279;
wire ng16132;
wire ng18883;
wire ng18836;
wire ng26811;
wire ng24218;
wire ng13182;
wire ng20977;
wire ng21040;
wire ng21080;
wire ng25271;
wire ng26532;
wire ng18866;
wire ng19178;
wire ng18867;
wire ng29617;
wire ng24230;
wire ng20955;
wire ng21021;
wire ng20900;
wire ng25268;
wire ng30291;
wire ng19153;
wire ng18906;
wire ng18957;
wire ng29184;
wire ng27332;
wire ng28357;
wire ng28362;
wire ng16692;
wire ng28325;
wire ng30301;
wire ng12433;
wire ng20310;
wire ng19167;
wire ng18942;
wire ng21882;
wire ng11545;
wire ng27340;
wire ng24545;
wire ng28366;
wire ng28990;
wire ng20353;
wire ng27722;
wire ng30300;
wire ng18754;
wire ng19163;
wire ng19162;
wire ng18968;
wire ng18669;
wire ng28352;
wire ng13443;
wire ng24083;
wire ng27682;
wire ng25246;
wire ng18781;
wire ng20343;
wire ng19157;
wire ng18975;
wire ng18719;
wire ng28356;
wire ng13442;
wire ng13450;
wire ng26789;
wire ng22155;
wire wire3193;
wire wire3281;
wire wire3282;
wire ng26137;
wire wire3138;
wire wire3224;
wire wire3425;
wire wire3049;
wire wire3142;
wire ng13002;
wire ng12866;
wire ng12959;
wire ng12978;
wire ng12933;
wire ng12836;
wire ng12899;
wire ng13022;
wire ng12994;
wire ng11730;
wire ng13123;
wire ng12324;
wire wire3199;
wire ng12288;
wire wire3200;
wire wire3201;
wire ng13134;
wire ng12233;
wire ng12271;
wire ng12124;
wire ng12008;
wire ng12306;
wire ng12329;
wire ng12184;
wire ng12234;
wire ng11965;
wire ng12068;
wire ng11964;
wire ng12231;
wire ng12305;
wire ng10839;
wire ng12269;
wire ng10822;
wire wire3351;
wire wire3352;
wire wire3926;
wire wire3945;
wire ng12180;
wire ng12108;
wire ng15970;
wire ng13165;
wire ng15950;
wire wire3283;
wire ng23979;
wire ng18079;
wire ng18183;
wire ng18346;
wire wire3054;
wire wire3065;
wire wire3326;
wire wire3368;
wire ng23486;
wire ng18319;
wire ng18395;
wire ng18478;
wire ng18578;
wire ng18606;
wire ng18053;
wire ng18231;
wire wire3055;
wire wire3066;
wire wire3105;
wire wire3369;
wire ng23537;
wire ng22157;
wire ng10747;
wire wire3370;
wire ng24038;
wire ng27566;
wire ng27576;
wire ng17031;
wire wire3371;
wire wire3372;
wire ng24695;
wire ng11663;
wire ng28529;
wire ng12820;
wire ng25958;
wire ng26327;
wire ng12968;
wire ng29677;
wire ng30033;
wire ng30015;
wire ng30016;
wire ng11600;
wire ng11647;
wire ng17086;
wire ng24712;
wire ng22399;
wire ng24683;
wire ng12876;
wire ng22381;
wire ng17051;
wire ng11644;
wire ng13378;
wire ng27834;
wire ng11687;
wire ng17151;
wire ng22400;
wire ng11653;
wire ng27892;
wire ng11955;
wire ng29713;
wire ng11330;
wire ng12250;
wire ng27824;
wire ng30622;
wire ng30926;
wire ng21711;
wire ng21796;
wire ng10706;
wire ng10238;
wire ng17124;
wire ng11678;
wire ng10677;
wire ng11952;
wire ng12005;
wire ng11733;
wire ng13146;
wire ng13113;
wire ng13137;
wire ng17973;
wire ng12945;
wire wire3046;
wire ng18218;
wire ng11624;
wire ng13142;
wire ng11800;
wire ng12352;
wire ng12195;
wire ng12991;
wire ng12107;
wire ng12941;
wire ng11902;
wire ng26126;
wire wire3252;
wire wire3204;
wire ng12245;
wire wire3205;
wire ng12249;
wire wire3206;
wire ng12292;
wire ng13126;
wire ng11875;
wire wire3296;
wire ng24009;
wire wire3139;
wire wire3310;
wire wire3221;
wire ng27551;
wire ng11870;
wire wire3197;
wire ng27550;
wire wire3374;
wire ng12755;
wire ng26915;
wire ng11675;
wire ng28501;
wire ng27563;
wire wire3175;
wire wire3359;
wire ng28556;
wire ng12971;
wire wire3180;
wire wire3190;
wire wire3361;
wire ng29680;
wire ng29670;
wire ng30030;
wire ng30032;
wire ng18419;
wire ng17887;
wire ng17807;
wire ng17729;
wire wire3106;
wire wire3284;
wire ng23478;
wire ng22396;
wire ng12916;
wire ng11621;
wire ng26145;
wire ng26151;
wire ng11873;
wire ng27811;
wire ng29728;
wire ng30034;
wire ng11781;
wire ng12970;
wire ng18561;
wire ng25853;
wire ng27751;
wire ng11860;
wire ng12121;
wire ng17197;
wire ng23539;
wire ng18363;
wire ng18441;
wire ng18195;
wire ng18290;
wire wire3067;
wire wire3285;
wire wire3375;
wire ng23502;
wire wire3286;
wire wire3287;
wire wire3333;
wire ng13145;
wire ng11721;
wire wire3246;
wire wire3247;
wire wire3248;
wire ng12145;
wire ng13001;
wire ng12100;
wire ng12044;
wire ng12698;
wire ng10793;
wire ng11915;
wire ng11726;
wire ng11833;
wire ng23495;
wire wire3377;
wire ng16655;
wire wire3748;
wire ng26374;
wire ng12992;
wire ng29672;
wire ng30021;
wire ng11630;
wire ng11666;
wire ng12248;
wire ng12097;
wire ng10814;
wire ng12152;
wire ng10801;
wire wire3288;
wire ng23071;
wire ng12974;
wire ng27875;
wire ng12999;
wire ng25099;
wire wire3194;
wire ng27577;
wire ng21746;
wire ng25874;
wire ng27756;
wire ng23349;
wire ng12920;
wire ng12890;
wire ng12852;
wire ng12789;
wire ng25818;
wire wire3210;
wire ng12216;
wire ng8430;
wire ng11889;
wire ng11975;
wire ng11882;
wire wire3304;
wire ng24043;
wire ng23335;
wire ng11828;
wire ng27529;
wire ng25078;
wire wire3353;
wire ng27528;
wire wire3380;
wire ng12949;
wire ng16672;
wire ng12930;
wire ng12797;
wire ng12858;
wire ng12828;
wire ng25964;
wire wire3234;
wire wire3935;
wire ng24676;
wire ng29912;
wire ng28584;
wire wire3426;
wire ng29671;
wire ng12207;
wire ng23107;
wire ng18598;
wire ng24723;
wire ng24700;
wire ng11946;
wire ng27802;
wire ng17942;
wire wire3196;
wire ng11263;
wire ng27883;
wire ng28842;
wire ng23377;
wire ng23368;
wire wire3327;
wire ng23533;
wire ng18096;
wire ng17998;
wire ng18492;
wire wire3056;
wire wire3107;
wire ng23511;
wire ng12194;
wire ng12172;
wire ng12112;
wire ng12035;
wire ng26087;
wire wire3944;
wire wire3253;
wire ng12060;
wire ng12293;
wire ng11999;
wire ng12263;
wire ng12171;
wire ng11914;
wire ng21770;
wire ng12169;
wire ng10851;
wire ng12291;
wire ng12214;
wire wire3233;
wire wire3354;
wire wire3364;
wire wire3437;
wire wire3440;
wire ng23340;
wire wire3530;
wire ng26869;
wire ng11917;
wire ng26931;
wire ng29681;
wire ng29920;
wire ng12033;
wire ng10789;
wire ng12080;
wire ng10784;
wire wire3344;
wire wire3345;
wire wire3929;
wire wire3949;
wire ng18548;
wire ng18639;
wire wire3289;
wire ng23521;
wire ng29741;
wire wire3183;
wire wire3341;
wire ng30594;
wire ng16643;
wire ng22016;
wire ng21991;
wire ng16693;
wire ng17985;
wire ng12146;
wire ng12967;
wire ng12000;
wire ng26154;
wire ng12849;
wire ng11916;
wire ng12880;
wire ng12781;
wire ng12939;
wire ng12747;
wire ng12912;
wire ng12328;
wire wire3328;
wire ng23489;
wire wire3290;
wire wire3220;
wire ng24004;
wire ng27850;
wire wire3235;
wire wire3930;
wire ng27743;
wire ng26878;
wire ng12043;
wire wire3117;
wire ng29732;
wire ng29705;
wire ng29751;
wire ng30035;
wire ng25082;
wire ng11962;
wire ng23372;
wire ng21976;
wire ng27585;
wire ng26947;
wire wire3908;
wire ng18458;
wire ng18514;
wire ng18383;
wire wire3068;
wire wire3291;
wire wire3386;
wire ng23518;
wire wire3444;
wire ng18325;
wire ng15830;
wire wire3259;
wire ng12208;
wire ng11784;
wire ng11896;
wire ng12162;
wire wire3292;
wire wire3293;
wire ng11912;
wire ng27567;
wire wire3570;
wire ng26887;
wire ng26925;
wire ng26283;
wire ng18630;
wire ng29748;
wire ng27729;
wire wire3150;
wire ng30610;
wire ng30614;
wire wire3925;
wire ng11807;
wire ng29684;
wire ng21996;
wire ng26938;
wire ng26928;
wire ng25969;
wire wire3909;
wire ng23513;
wire wire3439;
wire ng18102;
wire ng12179;
wire ng12099;
wire ng11991;
wire ng11935;
wire ng11773;
wire ng26096;
wire ng26099;
wire wire3140;
wire ng22005;
wire wire3595;
wire wire3236;
wire ng25954;
wire ng25764;
wire wire3237;
wire wire3936;
wire ng27738;
wire ng26897;
wire ng27482;
wire wire3118;
wire ng13399;
wire ng30588;
wire ng30632;
wire wire3189;
wire wire3338;
wire ng30602;
wire ng25091;
wire ng27814;
wire ng27827;
wire ng11988;
wire ng22083;
wire ng22050;
wire ng23528;
wire ng10711;
wire ng26107;
wire ng26110;
wire wire3141;
wire wire3229;
wire wire3833;
wire wire3137;
wire wire3230;
wire ng13055;
wire ng11831;
wire ng11872;
wire ng13004;
wire ng23353;
wire wire3389;
wire ng26941;
wire wire3119;
wire ng22093;
wire ng27855;
wire ng29721;
wire ng22108;
wire ng23331;
wire ng23325;
wire wire3151;
wire ng18556;
wire ng18212;
wire ng18115;
wire wire3108;
wire wire3297;
wire ng23505;
wire ng11839;
wire wire3216;
wire ng11863;
wire ng30597;
wire wire3198;
wire ng27382;
wire ng27379;
wire ng28845;
wire ng27113;
wire wire3143;
wire ng30629;
wire wire3427;
wire ng11744;
wire ng11905;
wire ng12154;
wire ng12048;
wire ng22134;
wire ng26902;
wire ng26892;
wire wire3302;
wire ng26906;
wire ng27462;
wire ng27900;
wire ng27730;
wire ng30605;
wire ng30927;
wire wire3303;
wire ng23320;
wire wire3395;
wire ng11987;
wire wire3277;
wire wire3227;
wire wire3835;
wire wire3834;
wire wire3442;
wire ng22118;
wire ng27157;
wire ng26911;
wire wire3120;
wire ng27897;
wire ng17194;
wire ng17177;
wire ng11992;
wire ng11938;
wire wire3278;
wire ng27865;
wire wire3836;
wire ng11830;
wire wire3217;
wire ng15757;
wire ng15719;
wire ng15841;
wire wire3397;
wire ng27582;
wire ng30031;
wire ng23388;
wire wire3307;
wire wire3308;
wire ng12057;
wire ng23360;
wire ng23950;
wire ng17183;
wire wire3400;
wire ng26417;
wire wire3323;
wire wire3403;
wire wire3921;
wire ng23497;
wire ng17162;
wire ng30305;
wire ng11981;
wire wire3174;
wire wire3339;
wire wire3942;
wire wire3313;
wire ng23526;
wire ng8381;
wire ng12082;
wire ng29710;
wire wire3280;
wire ng11974;
wire wire3314;
wire ng11188;
wire ng12988;
wire wire3188;
wire wire3336;
wire wire3697;
wire wire3156;
wire wire3435;
wire wire3315;
wire wire3316;
wire wire3317;
wire wire3195;
wire ng11262;
wire wire3309;
wire ng11979;
wire ng12036;
wire wire3279;
wire ng29718;
wire wire3319;
wire wire3157;
wire ng12026;
wire wire3121;
wire wire3122;
wire ng12090;
wire ng12224;
wire ng22009;
wire wire3123;
wire wire3124;
wire ng23395;
wire wire3324;
wire ng23381;
wire ng21983;
wire ng22069;
wire wire3320;
wire wire3321;
wire ng22021;
wire wire3159;
wire ng12213;
wire ng23364;
wire wire3325;
wire wire3073;
wire ng17139;
wire ng23344;
wire wire3784;
wire wire3788;
wire ng26918;
wire wire3074;
wire wire3075;
wire wire3076;
wire wire3116;
wire wire3034;
wire wire3035;
wire wire3036;
wire wire3037;
wire wire3050;
wire wire3079;
wire wire3097;
wire wire3101;
wire wire3167;
wire wire3168;
wire wire3213;
wire wire3322;
wire wire3388;
wire wire3390;
wire wire3391;
wire wire3392;
wire wire3393;
wire wire3394;
wire wire3396;
wire wire3404;
wire wire3422;
wire wire3423;
wire wire3424;
wire wire3441;
wire wire3448;
wire wire3449;
wire wire3450;
wire wire3451;
wire wire3488;
wire wire3512;
wire wire3515;
wire wire3527;
wire wire3528;
wire wire3529;
wire wire3545;
wire wire3564;
wire wire3594;
wire wire3621;
wire wire3639;
wire wire3660;
wire wire3661;
wire wire3672;
wire wire3673;
wire wire3714;
wire wire3715;
wire wire3721;
wire wire3727;
wire wire3808;
wire wire3815;
wire wire3845;
wire wire3846;
wire wire3850;
wire wire3851;
wire wire3852;
wire wire3854;
wire wire3855;
wire wire3856;
wire wire3857;
wire wire3858;
wire wire3885;
wire wire3886;
wire wire3893;
wire wire3894;
wire wire3902;
wire wire3931;
wire wire4030;
wire wire4076;
wire wire4080;
wire wire4104;
wire wire4105;
wire wire4115;
wire wire4121;
wire wire4133;
wire wire4135;
wire wire4155;
wire wire4214;
wire wire4215;
wire wire4217;
wire wire4239;
wire wire4250;
wire wire4254;
wire wire4255;
wire wire4265;
wire wire4271;
wire wire4282;
wire wire4284;
wire wire4286;
wire wire4287;
wire wire4288;
wire wire4291;
wire wire4292;
wire wire4302;
wire wire4305;
wire wire4306;
wire wire4309;
wire wire4315;
wire wire4319;
wire wire4320;
wire wire4321;
wire wire4323;
wire wire4345;
wire wire4346;
wire wire4347;
wire wire4348;
wire wire4349;
wire wire4350;
wire wire4351;
wire wire4359;
wire wire4360;
wire wire4376;
wire wire4379;
wire wire4380;
wire wire4381;
wire wire4382;
wire wire4383;
wire wire4384;
wire wire4385;
wire wire4386;
wire wire4397;
wire wire4415;
wire wire4416;
wire wire4420;
wire wire4425;
wire wire4426;
wire wire4432;
wire wire4434;
wire wire4436;
wire wire4467;
wire wire4476;
wire wire4477;
wire wire4478;
wire wire4479;
wire wire4487;
wire wire4493;
wire wire4506;
wire wire4560;
wire wire4568;
wire wire4571;
wire wire4588;
wire wire4610;
wire wire4647;
wire wire4648;
wire wire4654;
wire wire4662;
wire wire4673;
wire wire4683;
wire wire4685;
wire wire4686;
wire wire4687;
wire wire4690;
wire wire4691;
wire wire4692;
wire wire4695;
wire wire4696;
wire wire4703;
wire wire4708;
wire wire4721;
wire wire4722;
wire wire4748;
wire wire4757;
wire wire4770;
wire wire4771;
wire wire4772;
wire wire4775;
wire wire4776;
wire wire4780;
wire wire4784;
wire wire4807;
wire wire4808;
wire wire4809;
wire wire4810;
wire wire4869;
wire wire4872;
wire wire4873;
wire wire4874;
wire wire4875;
wire wire4888;
wire wire4889;
wire wire4918;
wire wire4928;
wire wire4932;
wire wire4947;
wire wire4955;
wire wire4961;
wire wire4964;
wire wire4975;
wire wire4983;
wire wire4985;
wire wire5013;
wire wire5021;
wire wire5029;
wire wire5030;
wire wire5031;
wire wire5034;
wire wire5035;
wire wire5049;
wire wire5060;
wire wire5069;
wire wire5070;
wire wire5071;
wire wire5072;
wire wire5073;
wire wire5074;
wire wire5075;
wire wire5088;
wire wire5091;
wire wire5092;
wire wire5093;
wire wire5094;
wire wire5096;
wire wire5101;
wire wire5102;
wire wire5104;
wire wire5109;
wire wire5110;
wire wire5112;
wire wire5113;
wire wire5114;
wire wire5117;
wire wire5118;
wire wire5120;
wire wire5125;
wire wire5126;
wire wire5128;
wire wire5129;
wire wire5130;
wire wire5131;
wire wire5132;
wire wire5133;
wire wire5134;
wire wire5136;
wire wire5141;
wire wire5142;
wire wire5144;
wire wire5145;
wire wire5146;
wire wire5147;
wire wire5148;
wire wire5149;
wire wire5150;
wire wire5152;
wire wire5153;
wire wire5154;
wire wire5155;
wire wire5156;
wire wire5157;
wire wire5158;
wire wire5160;
wire wire5161;
wire wire5162;
wire wire5165;
wire wire5166;
wire wire5168;
wire wire5169;
wire wire5170;
wire wire5173;
wire wire5174;
wire wire5176;
wire wire5177;
wire wire5199;
wire wire5200;
wire wire5202;
wire wire5203;
wire wire5204;
wire wire5205;
wire wire5206;
wire wire5210;
wire wire5211;
wire wire5212;
wire wire5213;
wire wire5214;
wire wire5216;
wire wire5217;
wire wire5219;
wire wire5220;
wire wire5222;
wire wire5223;
wire wire5224;
wire wire5225;
wire wire5226;
wire wire5227;
wire wire5228;
wire wire5229;
wire wire5230;
wire wire5231;
wire wire5232;
wire wire5237;
wire wire5238;
wire wire5239;
wire wire5244;
wire wire5245;
wire wire5248;
wire wire5251;
wire wire5252;
wire wire5253;
wire wire5254;
wire wire5256;
wire wire5257;
wire wire5258;
wire wire5261;
wire wire5262;
wire wire5264;
wire wire5267;
wire wire5268;
wire wire5269;
wire wire5270;
wire wire5272;
wire wire5273;
wire wire5274;
wire wire5275;
wire wire5276;
wire wire5277;
wire wire5278;
wire wire5286;
wire wire5287;
wire wire5288;
wire wire5303;
wire wire5326;
wire wire5335;
wire wire5341;
wire wire5351;
wire wire5356;
wire wire5370;
wire wire5371;
wire wire5382;
wire wire5419;
wire wire5422;
wire wire5423;
wire wire5424;
wire wire5425;
wire wire5435;
wire wire5442;
wire wire5443;
wire wire5445;
wire wire5464;
wire wire5469;
wire wire5475;
wire wire5492;
wire wire5512;
wire wire5525;
wire wire5526;
wire wire5527;
wire wire5557;
wire wire5564;
wire wire5571;
wire wire5572;
wire wire5573;
wire wire5577;
wire wire5605;
wire wire5606;
wire wire5619;
wire wire5626;
wire wire5673;
wire wire5694;
wire wire5702;
wire wire5707;
wire wire5726;
wire wire5739;
wire wire5740;
wire wire5749;
wire wire5751;
wire wire5752;
wire wire5753;
wire wire5754;
wire wire5755;
wire wire5759;
wire wire5760;
wire wire5761;
wire wire5762;
wire wire5763;
wire wire5765;
wire wire5766;
wire wire5768;
wire wire5769;
wire wire5771;
wire wire5772;
wire wire5774;
wire wire5775;
wire wire5780;
wire wire5781;
wire wire5787;
wire wire5793;
wire wire5794;
wire wire5795;
wire wire5804;
wire wire5805;
wire wire5810;
wire wire5831;
wire wire5832;
wire wire5833;
wire wire5836;
wire wire5837;
wire wire5849;
wire wire5850;
wire wire5851;
wire wire5854;
wire wire5858;
wire wire5879;
wire wire5883;
wire wire5886;
wire wire5893;
wire wire5894;
wire wire5895;
wire wire5899;
wire wire5902;
wire wire5903;
wire wire5963;
wire wire5964;
wire wire5965;
wire wire5973;
wire wire5976;
wire wire5993;
wire wire5994;
wire wire6005;
wire wire6006;
wire wire6015;
wire wire6043;
wire wire6055;
wire wire6057;
wire wire6089;
wire wire6094;
wire wire6095;
wire wire6103;
wire wire6105;
wire wire6107;
wire wire6114;
wire wire6138;
wire wire6140;
wire wire6155;
wire wire6170;
wire wire6171;
wire wire6175;
wire wire6176;
wire wire6177;
wire wire6178;
wire wire6179;
wire wire6180;
wire wire6188;
wire wire6190;
wire wire6207;
wire wire6208;
wire wire6209;
wire wire6212;
wire wire6213;
wire wire6217;
wire wire6218;
wire wire6219;
wire wire6220;
wire wire6221;
wire wire6222;
wire wire6223;
wire wire6240;
wire wire6255;
wire wire6263;
wire wire6278;
wire wire6281;
wire wire6282;
wire wire6283;
wire wire6284;
wire wire6292;
wire wire6301;
wire wire6302;
wire wire6303;
wire wire6304;
wire wire6305;
wire wire6306;
wire wire6307;
wire wire6308;
wire wire6329;
wire wire6330;
wire wire6331;
wire wire6332;
wire wire6333;
wire wire6334;
wire wire6335;
wire wire6337;
wire wire6342;
wire wire6343;
wire wire6345;
wire wire6346;
wire wire6347;
wire wire6348;
wire wire6349;
wire wire6350;
wire wire6351;
wire wire6353;
wire wire6358;
wire wire6359;
wire wire6361;
wire wire6362;
wire wire6363;
wire wire6366;
wire wire6367;
wire wire6369;
wire wire6370;
wire wire6371;
wire wire6374;
wire wire6375;
wire wire6377;
wire wire6380;
wire wire6381;
wire wire6382;
wire wire6383;
wire wire6385;
wire wire6386;
wire wire6387;
wire wire6388;
wire wire6389;
wire wire6390;
wire wire6391;
wire wire6393;
wire wire6394;
wire wire6395;
wire wire6398;
wire wire6399;
wire wire6401;
wire wire6402;
wire wire6403;
wire wire6406;
wire wire6407;
wire wire6409;
wire wire6410;
wire wire6411;
wire wire6414;
wire wire6415;
wire wire6424;
wire wire6425;
wire wire6434;
wire wire6441;
wire wire6442;
wire wire6443;
wire wire6444;
wire wire6445;
wire wire6446;
wire wire6447;
wire wire6448;
wire wire6452;
wire wire6459;
wire wire6464;
wire wire6465;
wire wire6468;
wire wire6473;
wire wire6474;
wire wire6488;
wire wire6508;
wire wire6514;
wire wire6515;
wire wire6516;
wire wire6519;
wire wire6520;
wire wire6532;
wire wire6533;
wire wire6534;
wire wire6535;
wire wire6536;
wire wire6537;
wire wire6538;
wire wire6539;
wire wire6544;
wire wire6545;
wire wire6546;
wire wire6547;
wire wire6552;
wire wire6553;
wire wire6564;
wire wire6572;
wire wire6581;
wire wire6582;
wire wire6583;
wire wire6584;
wire wire6585;
wire wire6586;
wire wire6587;
wire wire6588;
wire wire6609;
wire wire6614;
wire wire6615;
wire wire6617;
wire wire6618;
wire wire6619;
wire wire6622;
wire wire6623;
wire wire6625;
wire wire6626;
wire wire6627;
wire wire6628;
wire wire6629;
wire wire6630;
wire wire6631;
wire wire6633;
wire wire6638;
wire wire6639;
wire wire6641;
wire wire6644;
wire wire6645;
wire wire6646;
wire wire6647;
wire wire6649;
wire wire6654;
wire wire6655;
wire wire6657;
wire wire6660;
wire wire6661;
wire wire6662;
wire wire6663;
wire wire6665;
wire wire6666;
wire wire6667;
wire wire6670;
wire wire6671;
wire wire6673;
wire wire6674;
wire wire6675;
wire wire6678;
wire wire6679;
wire wire6681;
wire wire6682;
wire wire6683;
wire wire6684;
wire wire6685;
wire wire6686;
wire wire6687;
wire wire6689;
wire wire6690;
wire wire6691;
wire wire6694;
wire wire6695;
wire wire6702;
wire wire6720;
wire wire6732;
wire wire6737;
wire wire6738;
wire wire6771;
wire wire6791;
wire wire6818;
wire wire6819;
wire wire6820;
wire wire6821;
wire wire6822;
wire wire6823;
wire wire6824;
wire wire6875;
wire wire6881;
wire wire6883;
wire wire6921;
wire wire6922;
wire wire6923;
wire wire6925;
wire wire6926;
wire wire6927;
wire wire6928;
wire wire6929;
wire wire6930;
wire wire6931;
wire wire6932;
wire wire6933;
wire wire6934;
wire wire6939;
wire wire6940;
wire wire6941;
wire wire6946;
wire wire6947;
wire wire6950;
wire wire6951;
wire wire6952;
wire wire6955;
wire wire6956;
wire wire6958;
wire wire6959;
wire wire6960;
wire wire6963;
wire wire6964;
wire wire6966;
wire wire6969;
wire wire6970;
wire wire6971;
wire wire6972;
wire wire6974;
wire wire6975;
wire wire6976;
wire wire6977;
wire wire6978;
wire wire6979;
wire wire6980;
wire wire6982;
wire wire6983;
wire wire6984;
wire wire6985;
wire wire6988;
wire wire6989;
wire wire6990;
wire wire6991;
wire wire6993;
wire wire6994;
wire wire6996;
wire wire6997;
wire wire6999;
wire wire7000;
wire wire7002;
wire wire7003;
wire wire7005;
wire wire7006;
wire wire7011;
wire wire7012;
wire wire7014;
wire wire7026;
wire wire7029;
wire wire7030;
wire wire7045;
wire wire7046;
wire wire7048;
wire wire7057;
wire wire7058;
wire wire7069;
wire wire7070;
wire wire7078;
wire wire7083;
wire wire7084;
wire wire7111;
wire wire7114;
wire wire7119;
wire wire7120;
wire wire7121;
wire wire7124;
wire wire7125;
wire wire7127;
wire wire7128;
wire wire7129;
wire wire7132;
wire wire7133;
wire wire7135;
wire wire7138;
wire wire7139;
wire wire7140;
wire wire7141;
wire wire7143;
wire wire7144;
wire wire7145;
wire wire7148;
wire wire7149;
wire wire7152;
wire wire7153;
wire wire7154;
wire wire7159;
wire wire7160;
wire wire7162;
wire wire7163;
wire wire7164;
wire wire7165;
wire wire7166;
wire wire7167;
wire wire7168;
wire wire7170;
wire wire7175;
wire wire7176;
wire wire7190;
wire wire7191;
wire wire7192;
wire wire7196;
wire wire7201;
wire wire7202;
wire wire7204;
wire wire7209;
wire wire7210;
wire wire7213;
wire wire7218;
wire wire7219;
wire wire7225;
wire wire7227;
wire wire7228;
wire wire7229;
wire wire7230;
wire wire7231;
wire wire7232;
wire wire7233;
wire wire7234;
wire wire7235;
wire wire7240;
wire wire7241;
wire wire7246;
wire wire7249;
wire wire7250;
wire wire7251;
wire wire7252;
wire wire7262;
wire wire7267;
wire wire7268;
wire wire7270;
wire wire7273;
wire wire7274;
wire wire7275;
wire wire7276;
wire wire7278;
wire wire7283;
wire wire7284;
wire wire7307;
wire wire7308;
wire wire7327;
wire wire7331;
wire wire7336;
wire wire7337;
wire wire7342;
wire wire7343;
wire wire7344;
wire wire7359;
wire wire7364;
wire wire7365;
wire wire7366;
wire wire7383;
wire wire7384;
wire wire7385;
wire wire7386;
wire wire7387;
wire wire7388;
wire wire7389;
wire wire7390;
wire wire7391;
wire wire7392;
wire wire7393;
wire wire7394;
wire wire7395;
wire wire7396;
wire wire7397;
wire wire7398;
wire wire7399;
wire wire7400;
wire wire7409;
wire wire7414;
wire wire7415;
wire wire7417;
wire wire7422;
wire wire7423;
wire wire7425;
wire wire7430;
wire wire7431;
wire wire7435;
wire wire7436;
wire wire7437;
wire wire7438;
wire wire7439;
wire wire7440;
wire wire7441;
wire wire7442;
wire wire7443;
wire wire7444;
wire wire7445;
wire wire7446;
wire wire7447;
wire wire7448;
wire wire7449;
wire wire7450;
wire wire7451;
wire wire7452;
wire wire7455;
wire wire7456;
wire wire7459;
wire wire7464;
wire wire7465;
wire wire7467;
wire wire7472;
wire wire7473;
wire wire7475;
wire wire7480;
wire wire7481;
wire wire7483;
wire wire7488;
wire wire7489;
wire wire7491;
wire wire7496;
wire wire7497;
wire wire7500;
wire wire7504;
wire wire7509;
wire wire7510;
wire wire7512;
wire wire7517;
wire wire7518;
wire wire7520;
wire wire7521;
wire wire7522;
wire wire7523;
wire wire7524;
wire wire7525;
wire wire7526;
wire wire7528;
wire wire7531;
wire wire7532;
wire wire7533;
wire wire7534;
wire wire7536;
wire wire7541;
wire wire7542;
wire wire7544;
wire wire7549;
wire wire7550;
wire wire7552;
wire wire7553;
wire wire7554;
wire wire7555;
wire wire7556;
wire wire7557;
wire wire7558;
wire wire7560;
wire wire7565;
wire wire7566;
wire wire7568;
wire wire7573;
wire wire7574;
wire wire7576;
wire wire7577;
wire wire7578;
wire wire7579;
wire wire7580;
wire wire7581;
wire wire7582;
wire wire7584;
wire wire7585;
wire wire7586;
wire wire7587;
wire wire7588;
wire wire7589;
wire wire7590;
wire wire7592;
wire wire7597;
wire wire7598;
wire wire7600;
wire wire7601;
wire wire7602;
wire wire7603;
wire wire7604;
wire wire7605;
wire wire7606;
wire wire7612;
wire wire7617;
wire wire7618;
wire wire7627;
wire wire7633;
wire wire7635;
wire wire7636;
wire wire7637;
wire wire7638;
wire wire7639;
wire wire7640;
wire wire7641;
wire wire7644;
wire wire7649;
wire wire7650;
wire wire7651;
wire wire7652;
wire wire7653;
wire wire7660;
wire wire7661;
wire wire7662;
wire wire7665;
wire wire7666;
wire wire7668;
wire wire7669;
wire wire7670;
wire wire7671;
wire wire7672;
wire wire7673;
wire wire7674;
wire wire7676;
wire wire7677;
wire wire7678;
wire wire7681;
wire wire7682;
wire wire7684;
wire wire7685;
wire wire7686;
wire wire7687;
wire wire7688;
wire wire7689;
wire wire7690;
wire wire7692;
wire wire7693;
wire wire7694;
wire wire7697;
wire wire7698;
wire wire7700;
wire wire7701;
wire wire7702;
wire wire7703;
wire wire7704;
wire wire7708;
wire wire7709;
wire wire7710;
wire wire7711;
wire wire7712;
wire wire7714;
wire wire7715;
wire wire7717;
wire wire7718;
wire wire7720;
wire wire7721;
wire wire7723;
wire wire7724;
wire wire7729;
wire wire7730;
wire wire7732;
wire wire7734;
wire wire7735;
wire wire7736;
wire wire7737;
wire wire7738;
wire wire7741;
wire wire7742;
wire wire7743;
wire wire7745;
wire wire7746;
wire wire7748;
wire wire7749;
wire wire7751;
wire wire7752;
wire wire7754;
wire wire7755;
wire wire7756;
wire wire7757;
wire wire7758;
wire wire7759;
wire wire7760;
wire wire7763;
wire wire7764;
wire wire7769;
wire wire7770;
wire wire7771;
wire wire7776;
wire wire7777;
wire wire7779;
wire wire7784;
wire wire7785;
wire wire7787;
wire wire7792;
wire wire7793;
wire wire7797;
wire wire7802;
wire wire7803;
wire wire7807;
wire wire7808;
wire wire7809;
wire wire7812;
wire wire7813;
wire wire7815;
wire wire7816;
wire wire7817;
wire wire7820;
wire wire7821;
wire wire7829;
wire wire7830;
wire wire7837;
wire wire7844;
wire wire7845;
wire wire7846;
wire wire7850;
wire wire7855;
wire wire7856;
wire wire7858;
wire wire7863;
wire wire7864;
wire wire7867;
wire wire7868;
wire wire7869;
wire wire7870;
wire wire7871;
wire wire7872;
wire wire7873;
wire wire7879;
wire wire7881;
wire wire7882;
wire wire7883;
wire wire7884;
wire wire7885;
wire wire7886;
wire wire7887;
wire wire7888;
wire wire7892;
wire wire7897;
wire wire7898;
wire wire7900;
wire wire7901;
wire wire7902;
wire wire7903;
wire wire7904;
wire wire7905;
wire wire7906;
wire wire7914;
wire wire7919;
wire wire7920;
wire wire7922;
wire wire7927;
wire wire7928;
wire wire7930;
wire wire7931;
wire wire7932;
wire wire7933;
wire wire7934;
wire wire7935;
wire wire7936;
wire wire7941;
wire wire7954;
wire wire7955;
wire wire7972;
wire wire7976;
wire wire7977;
wire wire7978;
wire wire7979;
wire wire7981;
wire wire7982;
wire wire7987;
wire wire7988;
wire wire7989;
wire wire8004;
wire wire8009;
wire wire8010;
wire wire8011;
wire wire8026;
wire wire8027;
wire wire8028;
wire wire8029;
wire wire8030;
wire wire8035;
wire wire8036;
wire wire8041;
wire wire8042;
wire wire8043;
wire wire8044;
wire wire8046;
wire wire8047;
wire wire8050;
wire wire8051;
wire wire8054;
wire wire8055;
wire wire8056;
wire wire8057;
wire wire8058;
wire wire8059;
wire wire8060;
wire wire8062;
wire wire8067;
wire wire8068;
wire wire8070;
wire wire8075;
wire wire8076;
wire wire8086;
wire wire8087;
wire wire8088;
wire wire8089;
wire wire8090;
wire wire8094;
wire wire8095;
wire wire8098;
wire wire8103;
wire wire8104;
wire wire8106;
wire wire8111;
wire wire8112;
wire wire8114;
wire wire8119;
wire wire8120;
wire wire8122;
wire wire8127;
wire wire8128;
wire wire8130;
wire wire8131;
wire wire8132;
wire wire8133;
wire wire8134;
wire wire8135;
wire wire8136;
wire wire8138;
wire wire8141;
wire wire8142;
wire wire8143;
wire wire8144;
wire wire8146;
wire wire8147;
wire wire8151;
wire wire8156;
wire wire8157;
wire wire8159;
wire wire8164;
wire wire8165;
wire wire8167;
wire wire8168;
wire wire8169;
wire wire8170;
wire wire8171;
wire wire8172;
wire wire8173;
wire wire8175;
wire wire8180;
wire wire8181;
wire wire8183;
wire wire8188;
wire wire8189;
wire wire8191;
wire wire8196;
wire wire8197;
wire wire8199;
wire wire8202;
wire wire8203;
wire wire8204;
wire wire8205;
wire wire8207;
wire wire8212;
wire wire8213;
wire wire8215;
wire wire8220;
wire wire8221;
wire wire8223;
wire wire8228;
wire wire8229;
wire wire8231;
wire wire8236;
wire wire8237;
wire wire8239;
wire wire8244;
wire wire8245;
wire wire8247;
wire wire8252;
wire wire8253;
wire wire8274;
wire wire8275;
wire wire8280;
wire wire8281;
wire wire8282;
wire wire8283;
wire wire8284;
wire wire8285;
wire wire8287;
wire wire8288;
wire wire8290;
wire wire8292;
wire wire8293;
wire wire8295;
wire wire8296;
wire wire8298;
wire wire8299;
wire wire8301;
wire wire8302;
wire wire8304;
wire wire8305;
wire wire8310;
wire wire8311;
wire wire8314;
wire wire8315;
wire wire8316;
wire wire8317;
wire wire8318;
wire wire8323;
wire wire8324;
wire wire8326;
wire wire8327;
wire wire8329;
wire wire8330;
wire wire8332;
wire wire8334;
wire wire8335;
wire wire8336;
wire wire8337;
wire wire8338;
wire wire8339;
wire wire8340;
wire wire8341;
wire wire8342;
wire wire8344;
wire wire8347;
wire wire8348;
wire wire8349;
wire wire8350;
wire wire8352;
wire wire8357;
wire wire8358;
wire wire8360;
wire wire8361;
wire wire8362;
wire wire8365;
wire wire8366;
wire wire8368;
wire wire8373;
wire wire8374;
wire wire8376;
wire wire8380;
wire wire8381;
wire wire8382;
wire wire8383;
wire wire8384;
wire wire8385;
wire wire8386;
wire wire8387;
wire wire8389;
wire wire8390;
wire wire8392;
wire wire8393;
wire wire8395;
wire wire8396;
wire wire8397;
wire wire8398;
wire wire8399;
wire wire8400;
wire wire8401;
wire wire8402;
wire wire8405;
wire wire8406;
wire wire8414;
wire wire8415;
wire wire8416;
wire wire8419;
wire wire8420;
wire wire8422;
wire wire8423;
wire wire8424;
wire wire8425;
wire wire8426;
wire wire8427;
wire wire8428;
wire wire8430;
wire wire8431;
wire wire8432;
wire wire8433;
wire wire8434;
wire wire8435;
wire wire8436;
wire wire8439;
wire wire8440;
wire wire8441;
wire wire8446;
wire wire8447;
wire wire8449;
wire wire8450;
wire wire8451;
wire wire8452;
wire wire8453;
wire wire8454;
wire wire8455;
wire wire8457;
wire wire8460;
wire wire8461;
wire wire8462;
wire wire8463;
wire wire8469;
wire wire8474;
wire wire8475;
wire wire8482;
wire wire8484;
wire wire8487;
wire wire8488;
wire wire8491;
wire wire8492;
wire wire8493;
wire wire8494;
wire wire8495;
wire wire8496;
wire wire8497;
wire wire8498;
wire wire8502;
wire wire8503;
wire wire8504;
wire wire8505;
wire wire8506;
wire wire8507;
wire wire8508;
wire wire8510;
wire wire8515;
wire wire8516;
wire wire8524;
wire wire8529;
wire wire8530;
wire wire8532;
wire wire8533;
wire wire8534;
wire wire8535;
wire wire8536;
wire wire8537;
wire wire8538;
wire wire8540;
wire wire8543;
wire wire8544;
wire wire8545;
wire wire8546;
wire wire8556;
wire wire8557;
wire wire8566;
wire wire8569;
wire wire8591;
wire wire8594;
wire wire8596;
wire wire8597;
wire wire8602;
wire wire8603;
wire wire8604;
wire wire8619;
wire wire8624;
wire wire8625;
wire wire8626;
wire wire8641;
wire wire8649;
wire wire8650;
wire wire8663;
wire wire8668;
wire wire8669;
wire wire8671;
wire wire8676;
wire wire8677;
wire wire8679;
wire wire8684;
wire wire8685;
wire wire8689;
wire wire8690;
wire wire8691;
wire wire8692;
wire wire8693;
wire wire8694;
wire wire8695;
wire wire8696;
wire wire8697;
wire wire8698;
wire wire8699;
wire wire8700;
wire wire8701;
wire wire8702;
wire wire8703;
wire wire8704;
wire wire8705;
wire wire8706;
wire wire8709;
wire wire8710;
wire wire8713;
wire wire8718;
wire wire8719;
wire wire8721;
wire wire8726;
wire wire8727;
wire wire8729;
wire wire8734;
wire wire8735;
wire wire8737;
wire wire8738;
wire wire8739;
wire wire8740;
wire wire8741;
wire wire8742;
wire wire8743;
wire wire8745;
wire wire8750;
wire wire8751;
wire wire8754;
wire wire8757;
wire wire8762;
wire wire8763;
wire wire8765;
wire wire8770;
wire wire8771;
wire wire8773;
wire wire8774;
wire wire8775;
wire wire8776;
wire wire8777;
wire wire8778;
wire wire8779;
wire wire8781;
wire wire8786;
wire wire8787;
wire wire8789;
wire wire8790;
wire wire8791;
wire wire8792;
wire wire8793;
wire wire8794;
wire wire8795;
wire wire8797;
wire wire8802;
wire wire8803;
wire wire8805;
wire wire8806;
wire wire8807;
wire wire8808;
wire wire8809;
wire wire8810;
wire wire8811;
wire wire8813;
wire wire8818;
wire wire8819;
wire wire8821;
wire wire8822;
wire wire8823;
wire wire8824;
wire wire8825;
wire wire8826;
wire wire8827;
wire wire8829;
wire wire8830;
wire wire8831;
wire wire8834;
wire wire8835;
wire wire8837;
wire wire8840;
wire wire8841;
wire wire8842;
wire wire8843;
wire wire8845;
wire wire8846;
wire wire8847;
wire wire8848;
wire wire8849;
wire wire8850;
wire wire8851;
wire wire8853;
wire wire8858;
wire wire8859;
wire wire8865;
wire wire8870;
wire wire8871;
wire wire8879;
wire wire8880;
wire wire8881;
wire wire8882;
wire wire8883;
wire wire8884;
wire wire8885;
wire wire8886;
wire wire8907;
wire wire8908;
wire wire8909;
wire wire8912;
wire wire8913;
wire wire8915;
wire wire8918;
wire wire8919;
wire wire8920;
wire wire8921;
wire wire8923;
wire wire8924;
wire wire8925;
wire wire8926;
wire wire8927;
wire wire8928;
wire wire8929;
wire wire8931;
wire wire8932;
wire wire8933;
wire wire8934;
wire wire8935;
wire wire8936;
wire wire8937;
wire wire8939;
wire wire8940;
wire wire8941;
wire wire8942;
wire wire8943;
wire wire8944;
wire wire8945;
wire wire8947;
wire wire8952;
wire wire8953;
wire wire8955;
wire wire8956;
wire wire8957;
wire wire8958;
wire wire8959;
wire wire8960;
wire wire8961;
wire wire8963;
wire wire8968;
wire wire8969;
wire wire8971;
wire wire8972;
wire wire8973;
wire wire8974;
wire wire8975;
wire wire8976;
wire wire8977;
wire wire8979;
wire wire8984;
wire wire8985;
wire wire8987;
wire wire8988;
wire wire8989;
wire wire8990;
wire wire8991;
wire wire8992;
wire wire8993;
wire wire9005;
wire wire9007;
wire wire9008;
wire wire9009;
wire wire9010;
wire wire9011;
wire wire9012;
wire wire9013;
wire wire9014;
wire wire9015;
wire wire9019;
wire wire9020;
wire wire9022;
wire wire9023;
wire wire9025;
wire wire9026;
wire wire9028;
wire wire9029;
wire wire9030;
wire wire9031;
wire wire9032;
wire wire9033;
wire wire9034;
wire wire9035;
wire wire9036;
wire wire9037;
wire wire9041;
wire wire9044;
wire wire9049;
wire wire9054;
wire wire9055;
wire wire9057;
wire wire9060;
wire wire9061;
wire wire9062;
wire wire9063;
wire wire9065;
wire wire9070;
wire wire9071;
wire wire9073;
wire wire9074;
wire wire9075;
wire wire9078;
wire wire9079;
wire wire9082;
wire wire9083;
wire wire9084;
wire wire9085;
wire wire9086;
wire wire9087;
wire wire9088;
wire wire9089;
wire wire9090;
wire wire9092;
wire wire9097;
wire wire9098;
wire wire9100;
wire wire9101;
wire wire9102;
wire wire9103;
wire wire9104;
wire wire9105;
wire wire9106;
wire wire9118;
wire wire9128;
wire wire9129;
wire wire9130;
wire wire9134;
wire wire9139;
wire wire9140;
wire wire9142;
wire wire9143;
wire wire9144;
wire wire9145;
wire wire9146;
wire wire9147;
wire wire9148;
wire wire9150;
wire wire9153;
wire wire9154;
wire wire9155;
wire wire9156;
wire wire9165;
wire wire9167;
wire wire9168;
wire wire9169;
wire wire9170;
wire wire9171;
wire wire9172;
wire wire9173;
wire wire9174;
wire wire9178;
wire wire9179;
wire wire9180;
wire wire9183;
wire wire9184;
wire wire9186;
wire wire9187;
wire wire9188;
wire wire9189;
wire wire9190;
wire wire9191;
wire wire9192;
wire wire9202;
wire wire9207;
wire wire9208;
wire wire9210;
wire wire9215;
wire wire9216;
wire wire9218;
wire wire9221;
wire wire9222;
wire wire9223;
wire wire9224;
wire wire9238;
wire wire9239;
wire wire9260;
wire wire9263;
wire wire9265;
wire wire9266;
wire wire9271;
wire wire9272;
wire wire9273;
wire wire9288;
wire wire9293;
wire wire9294;
wire wire9295;
wire wire9313;
wire wire9318;
wire wire9319;
wire wire9332;
wire wire9337;
wire wire9338;
wire wire9340;
wire wire9345;
wire wire9346;
wire wire9356;
wire wire9357;
wire wire9358;
wire wire9359;
wire wire9360;
wire wire9364;
wire wire9365;
wire wire9368;
wire wire9373;
wire wire9374;
wire wire9376;
wire wire9381;
wire wire9382;
wire wire9384;
wire wire9389;
wire wire9390;
wire wire9392;
wire wire9393;
wire wire9394;
wire wire9395;
wire wire9396;
wire wire9397;
wire wire9398;
wire wire9400;
wire wire9405;
wire wire9406;
wire wire9408;
wire wire9413;
wire wire9414;
wire wire9416;
wire wire9421;
wire wire9422;
wire wire9425;
wire wire9429;
wire wire9434;
wire wire9435;
wire wire9437;
wire wire9442;
wire wire9443;
wire wire9445;
wire wire9450;
wire wire9451;
wire wire9453;
wire wire9458;
wire wire9459;
wire wire9461;
wire wire9464;
wire wire9465;
wire wire9466;
wire wire9467;
wire wire9469;
wire wire9472;
wire wire9473;
wire wire9474;
wire wire9475;
wire wire9477;
wire wire9482;
wire wire9483;
wire wire9485;
wire wire9490;
wire wire9491;
wire wire9493;
wire wire9498;
wire wire9499;
wire wire9501;
wire wire9506;
wire wire9507;
wire wire9509;
wire wire9514;
wire wire9515;
wire wire9517;
wire wire9518;
wire wire9519;
wire wire9520;
wire wire9521;
wire wire9522;
wire wire9523;
wire wire9525;
wire wire9530;
wire wire9531;
wire wire9538;
wire wire9542;
wire wire9543;
wire wire9544;
wire wire9547;
wire wire9548;
wire wire9549;
wire wire9550;
wire wire9559;
wire wire30881;
wire wire30883;
wire wire30884;
wire wire30886;
wire wire30887;
wire wire30889;
wire wire30892;
wire wire30893;
wire wire30896;
wire wire30897;
wire wire30898;
wire wire30899;
wire wire30900;
wire wire30902;
wire wire30903;
wire wire30904;
wire wire30905;
wire wire30906;
wire wire30911;
wire wire30912;
wire wire30913;
wire wire30914;
wire wire30915;
wire wire30918;
wire wire30924;
wire wire30925;
wire wire30927;
wire wire30928;
wire wire30934;
wire wire30935;
wire wire30937;
wire wire30938;
wire wire30944;
wire wire30945;
wire wire30947;
wire wire30948;
wire wire30954;
wire wire30955;
wire wire30957;
wire wire30958;
wire wire30964;
wire wire30965;
wire wire30967;
wire wire30968;
wire wire30974;
wire wire30975;
wire wire30977;
wire wire30978;
wire wire30979;
wire wire30985;
wire wire30986;
wire wire30988;
wire wire30989;
wire wire30995;
wire wire30996;
wire wire30998;
wire wire30999;
wire wire31008;
wire wire31009;
wire wire31015;
wire wire31016;
wire wire31018;
wire wire31019;
wire wire31025;
wire wire31028;
wire wire31029;
wire wire31035;
wire wire31038;
wire wire31039;
wire wire31045;
wire wire31046;
wire wire31048;
wire wire31049;
wire wire31050;
wire wire31051;
wire wire31052;
wire wire31053;
wire wire31054;
wire wire31057;
wire wire31058;
wire wire31059;
wire wire31060;
wire wire31061;
wire wire31062;
wire wire31063;
wire wire31065;
wire wire31066;
wire wire31067;
wire wire31074;
wire wire31075;
wire wire31077;
wire wire31078;
wire wire31079;
wire wire31081;
wire wire31083;
wire wire31084;
wire wire31085;
wire wire31086;
wire wire31087;
wire wire31089;
wire wire31091;
wire wire31092;
wire wire31102;
wire wire31103;
wire wire31106;
wire wire31112;
wire wire31113;
wire wire31115;
wire wire31116;
wire wire31122;
wire wire31123;
wire wire31126;
wire wire31129;
wire wire31130;
wire wire31131;
wire wire31132;
wire wire31133;
wire wire31134;
wire wire31137;
wire wire31138;
wire wire31143;
wire wire31144;
wire wire31145;
wire wire31147;
wire wire31149;
wire wire31156;
wire wire31157;
wire wire31159;
wire wire31160;
wire wire31162;
wire wire31164;
wire wire31166;
wire wire31167;
wire wire31168;
wire wire31171;
wire wire31172;
wire wire31178;
wire wire31179;
wire wire31181;
wire wire31182;
wire wire31191;
wire wire31192;
wire wire31198;
wire wire31199;
wire wire31201;
wire wire31202;
wire wire31208;
wire wire31209;
wire wire31211;
wire wire31212;
wire wire31214;
wire wire31215;
wire wire31216;
wire wire31218;
wire wire31220;
wire wire31221;
wire wire31222;
wire wire31223;
wire wire31224;
wire wire31225;
wire wire31226;
wire wire31227;
wire wire31231;
wire wire31232;
wire wire31233;
wire wire31234;
wire wire31235;
wire wire31236;
wire wire31245;
wire wire31248;
wire wire31249;
wire wire31250;
wire wire31251;
wire wire31261;
wire wire31264;
wire wire31265;
wire wire31266;
wire wire31267;
wire wire31269;
wire wire31270;
wire wire31271;
wire wire31272;
wire wire31273;
wire wire31274;
wire wire31279;
wire wire31281;
wire wire31283;
wire wire31284;
wire wire31285;
wire wire31287;
wire wire31289;
wire wire31292;
wire wire31293;
wire wire31297;
wire wire31298;
wire wire31311;
wire wire31312;
wire wire31314;
wire wire31315;
wire wire31321;
wire wire31322;
wire wire31324;
wire wire31325;
wire wire31331;
wire wire31334;
wire wire31335;
wire wire31336;
wire wire31345;
wire wire31346;
wire wire31353;
wire wire31355;
wire wire31356;
wire wire31360;
wire wire31361;
wire wire31362;
wire wire31365;
wire wire31368;
wire wire31370;
wire wire31372;
wire wire31374;
wire wire31375;
wire wire31376;
wire wire31377;
wire wire31382;
wire wire31383;
wire wire31391;
wire wire31392;
wire wire31394;
wire wire31395;
wire wire31404;
wire wire31405;
wire wire31411;
wire wire31414;
wire wire31415;
wire wire31418;
wire wire31419;
wire wire31420;
wire wire31426;
wire wire31427;
wire wire31428;
wire wire31431;
wire wire31432;
wire wire31436;
wire wire31437;
wire wire31438;
wire wire31449;
wire wire31450;
wire wire31456;
wire wire31457;
wire wire31459;
wire wire31460;
wire wire31469;
wire wire31470;
wire wire31471;
wire wire31472;
wire wire31479;
wire wire31480;
wire wire31482;
wire wire31483;
wire wire31489;
wire wire31492;
wire wire31493;
wire wire31500;
wire wire31502;
wire wire31503;
wire wire31509;
wire wire31510;
wire wire31512;
wire wire31513;
wire wire31514;
wire wire31518;
wire wire31522;
wire wire31523;
wire wire31524;
wire wire31550;
wire wire31551;
wire wire31553;
wire wire31555;
wire wire31557;
wire wire31559;
wire wire31562;
wire wire31565;
wire wire31568;
wire wire31577;
wire wire31578;
wire wire31579;
wire wire31580;
wire wire31582;
wire wire31584;
wire wire31585;
wire wire31586;
wire wire31587;
wire wire31588;
wire wire31589;
wire wire31591;
wire wire31592;
wire wire31602;
wire wire31605;
wire wire31606;
wire wire31613;
wire wire31615;
wire wire31616;
wire wire31627;
wire wire31628;
wire wire31639;
wire wire31640;
wire wire31651;
wire wire31652;
wire wire31663;
wire wire31664;
wire wire31672;
wire wire31673;
wire wire31675;
wire wire31676;
wire wire31684;
wire wire31685;
wire wire31687;
wire wire31688;
wire wire31699;
wire wire31700;
wire wire31708;
wire wire31709;
wire wire31711;
wire wire31712;
wire wire31723;
wire wire31724;
wire wire31727;
wire wire31728;
wire wire31729;
wire wire31730;
wire wire31731;
wire wire31732;
wire wire31733;
wire wire31734;
wire wire31735;
wire wire31741;
wire wire31742;
wire wire31743;
wire wire31746;
wire wire31748;
wire wire31750;
wire wire31752;
wire wire31753;
wire wire31754;
wire wire31755;
wire wire31760;
wire wire31761;
wire wire31767;
wire wire31768;
wire wire31770;
wire wire31771;
wire wire31774;
wire wire31775;
wire wire31785;
wire wire31786;
wire wire31793;
wire wire31795;
wire wire31796;
wire wire31805;
wire wire31806;
wire wire31812;
wire wire31815;
wire wire31816;
wire wire31817;
wire wire31823;
wire wire31824;
wire wire31826;
wire wire31827;
wire wire31828;
wire wire31834;
wire wire31835;
wire wire31837;
wire wire31838;
wire wire31844;
wire wire31845;
wire wire31847;
wire wire31848;
wire wire31854;
wire wire31855;
wire wire31857;
wire wire31858;
wire wire31867;
wire wire31868;
wire wire31874;
wire wire31875;
wire wire31877;
wire wire31878;
wire wire31887;
wire wire31888;
wire wire31897;
wire wire31898;
wire wire31904;
wire wire31905;
wire wire31907;
wire wire31908;
wire wire31909;
wire wire31910;
wire wire31911;
wire wire31912;
wire wire31915;
wire wire31916;
wire wire31918;
wire wire31919;
wire wire31920;
wire wire31921;
wire wire31922;
wire wire31924;
wire wire31925;
wire wire31931;
wire wire31932;
wire wire31934;
wire wire31935;
wire wire31936;
wire wire31937;
wire wire31938;
wire wire31939;
wire wire31963;
wire wire31964;
wire wire31967;
wire wire31973;
wire wire31974;
wire wire31976;
wire wire31977;
wire wire31983;
wire wire31984;
wire wire31987;
wire wire31996;
wire wire31997;
wire wire31998;
wire wire31999;
wire wire32000;
wire wire32001;
wire wire32004;
wire wire32005;
wire wire32010;
wire wire32011;
wire wire32017;
wire wire32018;
wire wire32020;
wire wire32021;
wire wire32023;
wire wire32025;
wire wire32027;
wire wire32028;
wire wire32030;
wire wire32032;
wire wire32034;
wire wire32035;
wire wire32038;
wire wire32039;
wire wire32045;
wire wire32046;
wire wire32048;
wire wire32049;
wire wire32058;
wire wire32059;
wire wire32065;
wire wire32066;
wire wire32068;
wire wire32069;
wire wire32071;
wire wire32072;
wire wire32073;
wire wire32075;
wire wire32077;
wire wire32078;
wire wire32079;
wire wire32080;
wire wire32081;
wire wire32082;
wire wire32083;
wire wire32084;
wire wire32088;
wire wire32089;
wire wire32090;
wire wire32091;
wire wire32092;
wire wire32093;
wire wire32102;
wire wire32105;
wire wire32106;
wire wire32107;
wire wire32108;
wire wire32118;
wire wire32121;
wire wire32122;
wire wire32123;
wire wire32124;
wire wire32126;
wire wire32127;
wire wire32128;
wire wire32129;
wire wire32130;
wire wire32131;
wire wire32135;
wire wire32136;
wire wire32140;
wire wire32142;
wire wire32144;
wire wire32145;
wire wire32146;
wire wire32147;
wire wire32148;
wire wire32149;
wire wire32150;
wire wire32151;
wire wire32155;
wire wire32156;
wire wire32157;
wire wire32160;
wire wire32161;
wire wire32164;
wire wire32166;
wire wire32174;
wire wire32177;
wire wire32178;
wire wire32184;
wire wire32185;
wire wire32187;
wire wire32188;
wire wire32197;
wire wire32198;
wire wire32199;
wire wire32200;
wire wire32206;
wire wire32207;
wire wire32209;
wire wire32210;
wire wire32219;
wire wire32220;
wire wire32224;
wire wire32225;
wire wire32226;
wire wire32229;
wire wire32231;
wire wire32233;
wire wire32235;
wire wire32236;
wire wire32237;
wire wire32238;
wire wire32243;
wire wire32244;
wire wire32245;
wire wire32246;
wire wire32247;
wire wire32248;
wire wire32249;
wire wire32252;
wire wire32253;
wire wire32259;
wire wire32260;
wire wire32262;
wire wire32263;
wire wire32269;
wire wire32272;
wire wire32273;
wire wire32282;
wire wire32283;
wire wire32289;
wire wire32290;
wire wire32292;
wire wire32293;
wire wire32303;
wire wire32304;
wire wire32313;
wire wire32314;
wire wire32321;
wire wire32323;
wire wire32324;
wire wire32332;
wire wire32334;
wire wire32335;
wire wire32337;
wire wire32339;
wire wire32341;
wire wire32343;
wire wire32360;
wire wire32363;
wire wire32366;
wire wire32377;
wire wire32378;
wire wire32379;
wire wire32380;
wire wire32384;
wire wire32385;
wire wire32386;
wire wire32387;
wire wire32388;
wire wire32389;
wire wire32396;
wire wire32397;
wire wire32399;
wire wire32400;
wire wire32407;
wire wire32409;
wire wire32410;
wire wire32416;
wire wire32419;
wire wire32420;
wire wire32429;
wire wire32430;
wire wire32431;
wire wire32432;
wire wire32434;
wire wire32440;
wire wire32441;
wire wire32443;
wire wire32444;
wire wire32445;
wire wire32446;
wire wire32448;
wire wire32449;
wire wire32451;
wire wire32452;
wire wire32456;
wire wire32458;
wire wire32459;
wire wire32460;
wire wire32461;
wire wire32462;
wire wire32463;
wire wire32464;
wire wire32465;
wire wire32466;
wire wire32469;
wire wire32470;
wire wire32471;
wire wire32486;
wire wire32487;
wire wire32489;
wire wire32490;
wire wire32492;
wire wire32494;
wire wire32500;
wire wire32504;
wire wire32508;
wire wire32511;
wire wire32514;
wire wire32524;
wire wire32525;
wire wire32526;
wire wire32527;
wire wire32529;
wire wire32531;
wire wire32532;
wire wire32533;
wire wire32534;
wire wire32535;
wire wire32536;
wire wire32538;
wire wire32539;
wire wire32540;
wire wire32541;
wire wire32543;
wire wire32545;
wire wire32546;
wire wire32547;
wire wire32549;
wire wire32552;
wire wire32553;
wire wire32554;
wire wire32556;
wire wire32559;
wire wire32560;
wire wire32561;
wire wire32563;
wire wire32564;
wire wire32566;
wire wire32567;
wire wire32568;
wire wire32569;
wire wire32575;
wire wire32576;
wire wire32578;
wire wire32587;
wire wire32588;
wire wire32590;
wire wire32591;
wire wire32597;
wire wire32598;
wire wire32600;
wire wire32601;
wire wire32607;
wire wire32608;
wire wire32610;
wire wire32611;
wire wire32617;
wire wire32618;
wire wire32620;
wire wire32621;
wire wire32630;
wire wire32631;
wire wire32637;
wire wire32638;
wire wire32640;
wire wire32641;
wire wire32647;
wire wire32648;
wire wire32650;
wire wire32651;
wire wire32652;
wire wire32658;
wire wire32659;
wire wire32661;
wire wire32662;
wire wire32668;
wire wire32671;
wire wire32672;
wire wire32678;
wire wire32679;
wire wire32681;
wire wire32682;
wire wire32688;
wire wire32689;
wire wire32691;
wire wire32692;
wire wire32698;
wire wire32699;
wire wire32701;
wire wire32702;
wire wire32703;
wire wire32709;
wire wire32710;
wire wire32712;
wire wire32713;
wire wire32715;
wire wire32716;
wire wire32717;
wire wire32718;
wire wire32721;
wire wire32722;
wire wire32724;
wire wire32725;
wire wire32726;
wire wire32727;
wire wire32728;
wire wire32730;
wire wire32731;
wire wire32740;
wire wire32741;
wire wire32742;
wire wire32744;
wire wire32746;
wire wire32747;
wire wire32748;
wire wire32749;
wire wire32750;
wire wire32752;
wire wire32754;
wire wire32755;
wire wire32765;
wire wire32766;
wire wire32769;
wire wire32775;
wire wire32776;
wire wire32778;
wire wire32779;
wire wire32785;
wire wire32786;
wire wire32789;
wire wire32792;
wire wire32793;
wire wire32794;
wire wire32795;
wire wire32796;
wire wire32797;
wire wire32800;
wire wire32801;
wire wire32806;
wire wire32807;
wire wire32816;
wire wire32817;
wire wire32819;
wire wire32825;
wire wire32828;
wire wire32829;
wire wire32831;
wire wire32833;
wire wire32835;
wire wire32837;
wire wire32839;
wire wire32840;
wire wire32841;
wire wire32842;
wire wire32843;
wire wire32844;
wire wire32845;
wire wire32846;
wire wire32847;
wire wire32848;
wire wire32855;
wire wire32856;
wire wire32858;
wire wire32859;
wire wire32865;
wire wire32866;
wire wire32869;
wire wire32875;
wire wire32876;
wire wire32878;
wire wire32879;
wire wire32883;
wire wire32884;
wire wire32886;
wire wire32887;
wire wire32893;
wire wire32894;
wire wire32895;
wire wire32896;
wire wire32897;
wire wire32898;
wire wire32899;
wire wire32902;
wire wire32903;
wire wire32904;
wire wire32906;
wire wire32907;
wire wire32908;
wire wire32918;
wire wire32921;
wire wire32922;
wire wire32923;
wire wire32924;
wire wire32934;
wire wire32937;
wire wire32938;
wire wire32939;
wire wire32940;
wire wire32942;
wire wire32943;
wire wire32944;
wire wire32945;
wire wire32946;
wire wire32947;
wire wire32952;
wire wire32954;
wire wire32956;
wire wire32957;
wire wire32958;
wire wire32959;
wire wire32960;
wire wire32961;
wire wire32962;
wire wire32963;
wire wire32975;
wire wire32977;
wire wire32979;
wire wire32985;
wire wire32986;
wire wire32988;
wire wire32989;
wire wire32995;
wire wire32996;
wire wire32998;
wire wire32999;
wire wire33008;
wire wire33009;
wire wire33018;
wire wire33019;
wire wire33023;
wire wire33024;
wire wire33025;
wire wire33033;
wire wire33034;
wire wire33036;
wire wire33037;
wire wire33039;
wire wire33041;
wire wire33043;
wire wire33045;
wire wire33046;
wire wire33047;
wire wire33048;
wire wire33053;
wire wire33054;
wire wire33063;
wire wire33064;
wire wire33070;
wire wire33071;
wire wire33074;
wire wire33080;
wire wire33081;
wire wire33083;
wire wire33084;
wire wire33087;
wire wire33088;
wire wire33089;
wire wire33091;
wire wire33097;
wire wire33098;
wire wire33099;
wire wire33101;
wire wire33102;
wire wire33103;
wire wire33105;
wire wire33106;
wire wire33107;
wire wire33108;
wire wire33115;
wire wire33117;
wire wire33118;
wire wire33124;
wire wire33125;
wire wire33127;
wire wire33128;
wire wire33135;
wire wire33137;
wire wire33138;
wire wire33144;
wire wire33145;
wire wire33147;
wire wire33148;
wire wire33154;
wire wire33155;
wire wire33157;
wire wire33158;
wire wire33164;
wire wire33165;
wire wire33167;
wire wire33168;
wire wire33184;
wire wire33186;
wire wire33187;
wire wire33189;
wire wire33191;
wire wire33193;
wire wire33201;
wire wire33205;
wire wire33208;
wire wire33211;
wire wire33221;
wire wire33222;
wire wire33223;
wire wire33224;
wire wire33226;
wire wire33228;
wire wire33229;
wire wire33230;
wire wire33231;
wire wire33232;
wire wire33233;
wire wire33248;
wire wire33249;
wire wire33251;
wire wire33252;
wire wire33254;
wire wire33256;
wire wire33258;
wire wire33260;
wire wire33270;
wire wire33273;
wire wire33276;
wire wire33286;
wire wire33287;
wire wire33288;
wire wire33289;
wire wire33293;
wire wire33294;
wire wire33295;
wire wire33296;
wire wire33297;
wire wire33298;
wire wire33306;
wire wire33308;
wire wire33309;
wire wire33318;
wire wire33319;
wire wire33326;
wire wire33328;
wire wire33329;
wire wire33336;
wire wire33338;
wire wire33339;
wire wire33340;
wire wire33341;
wire wire33343;
wire wire33353;
wire wire33354;
wire wire33355;
wire wire33357;
wire wire33359;
wire wire33361;
wire wire33363;
wire wire33364;
wire wire33365;
wire wire33366;
wire wire33367;
wire wire33368;
wire wire33369;
wire wire33370;
wire wire33371;
wire wire33372;
wire wire33376;
wire wire33377;
wire wire33378;
wire wire33380;
wire wire33382;
wire wire33383;
wire wire33384;
wire wire33385;
wire wire33387;
wire wire33388;
wire wire33390;
wire wire33391;
wire wire33392;
wire wire33393;
wire wire33398;
wire wire33399;
wire wire33401;
wire wire33402;
wire wire33403;
wire wire33404;
wire wire33405;
wire wire33413;
wire wire33414;
wire wire33415;
wire wire33416;
wire wire33417;
wire wire33425;
wire wire33426;
wire wire33428;
wire wire33429;
wire wire33438;
wire wire33439;
wire wire33445;
wire wire33446;
wire wire33448;
wire wire33449;
wire wire33458;
wire wire33459;
wire wire33468;
wire wire33469;
wire wire33475;
wire wire33476;
wire wire33478;
wire wire33479;
wire wire33485;
wire wire33486;
wire wire33488;
wire wire33489;
wire wire33498;
wire wire33499;
wire wire33505;
wire wire33506;
wire wire33508;
wire wire33509;
wire wire33515;
wire wire33516;
wire wire33518;
wire wire33519;
wire wire33528;
wire wire33529;
wire wire33535;
wire wire33536;
wire wire33538;
wire wire33539;
wire wire33545;
wire wire33546;
wire wire33548;
wire wire33549;
wire wire33550;
wire wire33551;
wire wire33557;
wire wire33560;
wire wire33561;
wire wire33563;
wire wire33564;
wire wire33565;
wire wire33566;
wire wire33569;
wire wire33570;
wire wire33572;
wire wire33573;
wire wire33574;
wire wire33575;
wire wire33576;
wire wire33578;
wire wire33579;
wire wire33585;
wire wire33586;
wire wire33588;
wire wire33589;
wire wire33590;
wire wire33591;
wire wire33592;
wire wire33593;
wire wire33617;
wire wire33618;
wire wire33621;
wire wire33627;
wire wire33628;
wire wire33630;
wire wire33631;
wire wire33637;
wire wire33638;
wire wire33640;
wire wire33641;
wire wire33647;
wire wire33648;
wire wire33651;
wire wire33660;
wire wire33661;
wire wire33662;
wire wire33663;
wire wire33664;
wire wire33665;
wire wire33668;
wire wire33669;
wire wire33674;
wire wire33675;
wire wire33676;
wire wire33677;
wire wire33678;
wire wire33679;
wire wire33703;
wire wire33704;
wire wire33706;
wire wire33707;
wire wire33713;
wire wire33714;
wire wire33716;
wire wire33717;
wire wire33723;
wire wire33724;
wire wire33726;
wire wire33727;
wire wire33736;
wire wire33737;
wire wire33738;
wire wire33739;
wire wire33740;
wire wire33741;
wire wire33744;
wire wire33745;
wire wire33747;
wire wire33749;
wire wire33751;
wire wire33752;
wire wire33754;
wire wire33755;
wire wire33756;
wire wire33766;
wire wire33769;
wire wire33770;
wire wire33771;
wire wire33772;
wire wire33782;
wire wire33785;
wire wire33786;
wire wire33787;
wire wire33788;
wire wire33790;
wire wire33791;
wire wire33792;
wire wire33793;
wire wire33794;
wire wire33795;
wire wire33799;
wire wire33800;
wire wire33805;
wire wire33807;
wire wire33808;
wire wire33809;
wire wire33811;
wire wire33812;
wire wire33813;
wire wire33814;
wire wire33815;
wire wire33819;
wire wire33823;
wire wire33824;
wire wire33827;
wire wire33829;
wire wire33837;
wire wire33838;
wire wire33840;
wire wire33841;
wire wire33847;
wire wire33850;
wire wire33851;
wire wire33857;
wire wire33858;
wire wire33860;
wire wire33861;
wire wire33862;
wire wire33868;
wire wire33871;
wire wire33872;
wire wire33876;
wire wire33877;
wire wire33878;
wire wire33886;
wire wire33887;
wire wire33889;
wire wire33890;
wire wire33892;
wire wire33894;
wire wire33896;
wire wire33898;
wire wire33899;
wire wire33900;
wire wire33901;
wire wire33906;
wire wire33907;
wire wire33913;
wire wire33914;
wire wire33917;
wire wire33923;
wire wire33924;
wire wire33926;
wire wire33927;
wire wire33934;
wire wire33935;
wire wire33937;
wire wire33938;
wire wire33940;
wire wire33941;
wire wire33942;
wire wire33944;
wire wire33948;
wire wire33954;
wire wire33955;
wire wire33957;
wire wire33958;
wire wire33967;
wire wire33968;
wire wire33974;
wire wire33975;
wire wire33977;
wire wire33978;
wire wire33986;
wire wire33988;
wire wire33989;
wire wire33995;
wire wire33998;
wire wire33999;
wire wire34006;
wire wire34008;
wire wire34009;
wire wire34016;
wire wire34018;
wire wire34019;
wire wire34020;
wire wire34024;
wire wire34028;
wire wire34034;
wire wire34035;
wire wire34037;
wire wire34038;
wire wire34040;
wire wire34041;
wire wire34042;
wire wire34043;
wire wire34044;
wire wire34045;
wire wire34048;
wire wire34049;
wire wire34051;
wire wire34052;
wire wire34054;
wire wire34055;
wire wire34057;
wire wire34058;
wire wire34060;
wire wire34061;
wire wire34062;
wire wire34063;
wire wire34064;
wire wire34065;
wire wire34066;
wire wire34067;
wire wire34068;
wire wire34069;
wire wire34070;
wire wire34071;
wire wire34072;
wire wire34074;
wire wire34075;
wire wire34076;
wire wire34079;
wire wire34081;
wire wire34082;
wire wire34083;
wire wire34084;
wire wire34087;
wire wire34088;
wire wire34089;
wire wire34091;
wire wire34093;
wire wire34094;
wire wire34095;
wire wire34096;
wire wire34097;
wire wire34099;
wire wire34100;
wire wire34114;
wire wire34115;
wire wire34117;
wire wire34118;
wire wire34120;
wire wire34122;
wire wire34124;
wire wire34134;
wire wire34138;
wire wire34141;
wire wire34144;
wire wire34154;
wire wire34155;
wire wire34156;
wire wire34157;
wire wire34161;
wire wire34162;
wire wire34163;
wire wire34164;
wire wire34165;
wire wire34166;
wire wire34176;
wire wire34177;
wire wire34183;
wire wire34186;
wire wire34187;
wire wire34194;
wire wire34196;
wire wire34197;
wire wire34198;
wire wire34199;
wire wire34201;
wire wire34202;
wire wire34204;
wire wire34205;
wire wire34213;
wire wire34215;
wire wire34216;
wire wire34217;
wire wire34219;
wire wire34221;
wire wire34223;
wire wire34225;
wire wire34226;
wire wire34227;
wire wire34228;
wire wire34229;
wire wire34230;
wire wire34231;
wire wire34232;
wire wire34235;
wire wire34236;
wire wire34237;
wire wire34238;
wire wire34239;
wire wire34243;
wire wire34244;
wire wire34245;
wire wire34247;
wire wire34249;
wire wire34250;
wire wire34251;
wire wire34252;
wire wire34253;
wire wire34254;
wire wire34255;
wire wire34260;
wire wire34261;
wire wire34262;
wire wire34264;
wire wire34265;
wire wire34266;
wire wire34267;
wire wire34269;
wire wire34270;
wire wire34273;
wire wire34274;
wire wire34281;
wire wire34283;
wire wire34284;
wire wire34289;
wire wire34290;
wire wire34291;
wire wire34293;
wire wire34294;
wire wire34295;
wire wire34296;
wire wire34297;
wire wire34298;
wire wire34299;
wire wire34300;
wire wire34301;
wire wire34302;
wire wire34303;
wire wire34304;
wire wire34305;
wire wire34306;
wire wire34307;
wire wire34308;
wire wire34309;
wire wire34310;
wire wire34311;
wire wire34312;
wire wire34313;
wire wire34314;
wire wire34315;
wire wire34316;
wire wire34317;
wire wire34318;
wire wire34319;
wire wire34320;
wire wire34321;
wire wire34322;
wire wire34323;
wire wire34324;
wire wire34325;
wire wire34326;
wire wire34327;
wire wire34328;
wire wire34329;
wire wire34330;
wire wire34331;
wire wire34332;
wire wire34333;
wire wire34334;
wire wire34335;
wire wire34336;
wire wire34337;
wire wire34338;
wire wire34339;
wire wire34340;
wire wire34341;
wire wire34342;
wire wire34343;
wire wire34344;
wire wire34345;
wire wire34346;
wire wire34351;
wire wire34352;
wire wire34353;
wire wire34354;
wire wire34355;
wire wire34356;
wire wire34357;
wire wire34358;
wire wire34359;
wire wire34360;
wire wire34361;
wire wire34362;
wire wire34363;
wire wire34364;
wire wire34371;
wire wire34372;
wire wire34373;
wire wire34374;
wire wire34385;
wire wire34386;
wire wire34389;
wire wire34390;
wire wire34395;
wire wire34402;
wire wire34403;
wire wire34410;
wire wire34412;
wire wire34418;
wire wire34419;
wire wire34421;
wire wire34422;
wire wire34428;
wire wire34429;
wire wire34430;
wire wire34432;
wire wire34434;
wire wire34435;
wire wire34438;
wire wire34439;
wire wire34440;
wire wire34449;
wire wire34450;
wire wire34451;
wire wire34452;
wire wire34453;
wire wire34459;
wire wire34460;
wire wire34462;
wire wire34463;
wire wire34469;
wire wire34470;
wire wire34472;
wire wire34473;
wire wire34482;
wire wire34484;
wire wire34485;
wire wire34496;
wire wire34497;
wire wire34505;
wire wire34508;
wire wire34509;
wire wire34517;
wire wire34518;
wire wire34520;
wire wire34521;
wire wire34530;
wire wire34532;
wire wire34533;
wire wire34544;
wire wire34545;
wire wire34553;
wire wire34556;
wire wire34557;
wire wire34566;
wire wire34568;
wire wire34569;
wire wire34578;
wire wire34580;
wire wire34581;
wire wire34584;
wire wire34585;
wire wire34586;
wire wire34587;
wire wire34588;
wire wire34589;
wire wire34590;
wire wire34591;
wire wire34592;
wire wire34598;
wire wire34599;
wire wire34600;
wire wire34603;
wire wire34605;
wire wire34607;
wire wire34609;
wire wire34610;
wire wire34611;
wire wire34612;
wire wire34617;
wire wire34618;
wire wire34619;
wire wire34620;
wire wire34622;
wire wire34625;
wire wire34633;
wire wire34634;
wire wire34636;
wire wire34637;
wire wire34638;
wire wire34642;
wire wire34645;
wire wire34648;
wire wire34651;
wire wire34653;
wire wire34655;
wire wire34657;
wire wire34658;
wire wire34663;
wire wire34664;
wire wire34668;
wire wire34675;
wire wire34677;
wire wire34679;
wire wire34686;
wire wire34689;
wire wire34690;
wire wire34696;
wire wire34697;
wire wire34700;
wire wire34706;
wire wire34707;
wire wire34709;
wire wire34710;
wire wire34716;
wire wire34719;
wire wire34722;
wire wire34725;
wire wire34727;
wire wire34729;
wire wire34731;
wire wire34732;
wire wire34737;
wire wire34738;
wire wire34741;
wire wire34742;
wire wire34743;
wire wire34744;
wire wire34746;
wire wire34747;
wire wire34748;
wire wire34755;
wire wire34757;
wire wire34758;
wire wire34767;
wire wire34768;
wire wire34776;
wire wire34777;
wire wire34779;
wire wire34780;
wire wire34791;
wire wire34792;
wire wire34800;
wire wire34801;
wire wire34803;
wire wire34804;
wire wire34813;
wire wire34815;
wire wire34816;
wire wire34825;
wire wire34827;
wire wire34828;
wire wire34836;
wire wire34839;
wire wire34840;
wire wire34851;
wire wire34852;
wire wire34861;
wire wire34863;
wire wire34864;
wire wire34873;
wire wire34875;
wire wire34876;
wire wire34879;
wire wire34880;
wire wire34881;
wire wire34882;
wire wire34883;
wire wire34884;
wire wire34885;
wire wire34886;
wire wire34887;
wire wire34893;
wire wire34894;
wire wire34895;
wire wire34898;
wire wire34900;
wire wire34902;
wire wire34904;
wire wire34905;
wire wire34906;
wire wire34907;
wire wire34912;
wire wire34913;
wire wire34916;
wire wire34924;
wire wire34927;
wire wire34928;
wire wire34932;
wire wire34933;
wire wire34934;
wire wire34937;
wire wire34948;
wire wire34949;
wire wire34956;
wire wire34958;
wire wire34962;
wire wire34963;
wire wire34965;
wire wire34969;
wire wire34970;
wire wire34971;
wire wire34972;
wire wire34973;
wire wire34974;
wire wire34978;
wire wire34982;
wire wire34983;
wire wire34985;
wire wire34987;
wire wire34989;
wire wire34990;
wire wire34992;
wire wire34996;
wire wire34997;
wire wire35003;
wire wire35004;
wire wire35007;
wire wire35013;
wire wire35014;
wire wire35018;
wire wire35019;
wire wire35020;
wire wire35021;
wire wire35022;
wire wire35023;
wire wire35029;
wire wire35030;
wire wire35032;
wire wire35033;
wire wire35038;
wire wire35039;
wire wire35040;
wire wire35041;
wire wire35042;
wire wire35043;
wire wire35044;
wire wire35045;
wire wire35046;
wire wire35047;
wire wire35057;
wire wire35060;
wire wire35061;
wire wire35062;
wire wire35063;
wire wire35064;
wire wire35065;
wire wire35066;
wire wire35067;
wire wire35068;
wire wire35069;
wire wire35070;
wire wire35071;
wire wire35072;
wire wire35073;
wire wire35074;
wire wire35075;
wire wire35076;
wire wire35077;
wire wire35078;
wire wire35079;
wire wire35080;
wire wire35081;
wire wire35082;
wire wire35083;
wire wire35084;
wire wire35085;
wire wire35086;
wire wire35087;
wire wire35088;
wire wire35089;
wire wire35090;
wire wire35091;
wire wire35092;
wire wire35093;
wire wire35094;
wire wire35095;
wire wire35096;
wire wire35097;
wire wire35098;
wire wire35099;
wire wire35100;
wire wire35101;
wire wire35102;
wire wire35103;
wire wire35104;
wire wire35105;
wire wire35106;
wire wire35107;
wire wire35108;
wire wire35109;
wire wire35110;
wire wire35115;
wire wire35116;
wire wire35117;
wire wire35118;
wire wire35119;
wire wire35120;
wire wire35121;
wire wire35122;
wire wire35123;
wire wire35124;
wire wire35125;
wire wire35126;
wire wire35127;
wire wire35128;
wire wire35135;
wire wire35136;
wire wire35137;
wire wire35138;
wire wire35143;
wire wire35144;
wire wire35146;
wire wire35147;
wire wire35148;
wire wire35150;
wire wire35154;
wire wire35156;
wire wire35157;
wire wire35159;
wire wire35160;
wire wire35161;
wire wire35162;
wire wire35163;
wire wire35164;
wire wire35165;
wire wire35167;
wire wire35169;
wire wire35170;
wire wire35171;
wire wire35172;
wire wire35174;
wire wire35175;
wire wire35184;
wire wire35186;
wire wire35190;
wire wire35191;
wire wire35193;
wire wire35194;
wire wire35195;
wire wire35197;
wire wire35199;
wire wire35200;
wire wire35202;
wire wire35203;
wire wire35208;
wire wire35210;
wire wire35211;
wire wire35225;
wire wire35226;
wire wire35228;
wire wire35229;
wire wire35231;
wire wire35233;
wire wire35235;
wire wire35237;
wire wire35247;
wire wire35250;
wire wire35253;
wire wire35263;
wire wire35264;
wire wire35265;
wire wire35266;
wire wire35270;
wire wire35271;
wire wire35272;
wire wire35273;
wire wire35274;
wire wire35275;
wire wire35277;
wire wire35278;
wire wire35280;
wire wire35281;
wire wire35284;
wire wire35285;
wire wire35288;
wire wire35294;
wire wire35295;
wire wire35304;
wire wire35306;
wire wire35307;
wire wire35308;
wire wire35309;
wire wire35310;
wire wire35318;
wire wire35319;
wire wire35320;
wire wire35321;
wire wire35323;
wire wire35325;
wire wire35326;
wire wire35327;
wire wire35328;
wire wire35330;
wire wire35331;
wire wire35336;
wire wire35337;
wire wire35338;
wire wire35341;
wire wire35345;
wire wire35346;
wire wire35347;
wire wire35349;
wire wire35350;
wire wire35352;
wire wire35358;
wire wire35362;
wire wire35367;
wire wire35368;
wire wire35369;
wire wire35371;
wire wire35375;
wire wire35378;
wire wire35379;
wire wire35380;
wire wire35381;
wire wire35384;
wire wire35390;
wire wire35391;
wire wire35394;
wire wire35395;
wire wire35396;
wire wire35397;
wire wire35405;
wire wire35408;
wire wire35409;
wire wire35418;
wire wire35419;
wire wire35426;
wire wire35428;
wire wire35429;
wire wire35430;
wire wire35437;
wire wire35440;
wire wire35441;
wire wire35442;
wire wire35444;
wire wire35445;
wire wire35446;
wire wire35447;
wire wire35448;
wire wire35449;
wire wire35450;
wire wire35451;
wire wire35454;
wire wire35455;
wire wire35456;
wire wire35457;
wire wire35458;
wire wire35462;
wire wire35463;
wire wire35473;
wire wire35475;
wire wire35477;
wire wire35479;
wire wire35489;
wire wire35492;
wire wire35495;
wire wire35505;
wire wire35506;
wire wire35507;
wire wire35508;
wire wire35510;
wire wire35512;
wire wire35513;
wire wire35514;
wire wire35515;
wire wire35516;
wire wire35517;
wire wire35519;
wire wire35521;
wire wire35522;
wire wire35524;
wire wire35525;
wire wire35527;
wire wire35528;
wire wire35530;
wire wire35532;
wire wire35534;
wire wire35536;
wire wire35538;
wire wire35539;
wire wire35540;
wire wire35541;
wire wire35542;
wire wire35543;
wire wire35544;
wire wire35549;
wire wire35550;
wire wire35551;
wire wire35553;
wire wire35554;
wire wire35555;
wire wire35557;
wire wire35564;
wire wire35565;
wire wire35566;
wire wire35568;
wire wire35574;
wire wire35575;
wire wire35577;
wire wire35578;
wire wire35585;
wire wire35587;
wire wire35588;
wire wire35597;
wire wire35598;
wire wire35607;
wire wire35608;
wire wire35614;
wire wire35615;
wire wire35617;
wire wire35618;
wire wire35627;
wire wire35628;
wire wire35634;
wire wire35635;
wire wire35637;
wire wire35638;
wire wire35645;
wire wire35647;
wire wire35648;
wire wire35655;
wire wire35657;
wire wire35658;
wire wire35664;
wire wire35665;
wire wire35667;
wire wire35668;
wire wire35674;
wire wire35677;
wire wire35678;
wire wire35687;
wire wire35688;
wire wire35690;
wire wire35691;
wire wire35692;
wire wire35693;
wire wire35694;
wire wire35695;
wire wire35698;
wire wire35699;
wire wire35701;
wire wire35703;
wire wire35705;
wire wire35707;
wire wire35708;
wire wire35709;
wire wire35710;
wire wire35711;
wire wire35712;
wire wire35713;
wire wire35714;
wire wire35716;
wire wire35717;
wire wire35721;
wire wire35723;
wire wire35725;
wire wire35732;
wire wire35734;
wire wire35735;
wire wire35737;
wire wire35738;
wire wire35739;
wire wire35740;
wire wire35741;
wire wire35742;
wire wire35745;
wire wire35746;
wire wire35747;
wire wire35748;
wire wire35750;
wire wire35751;
wire wire35752;
wire wire35753;
wire wire35755;
wire wire35758;
wire wire35759;
wire wire35768;
wire wire35769;
wire wire35770;
wire wire35771;
wire wire35772;
wire wire35774;
wire wire35775;
wire wire35776;
wire wire35777;
wire wire35778;
wire wire35779;
wire wire35780;
wire wire35781;
wire wire35790;
wire wire35791;
wire wire35792;
wire wire35794;
wire wire35795;
wire wire35796;
wire wire35798;
wire wire35799;
wire wire35802;
wire wire35806;
wire wire35812;
wire wire35814;
wire wire35816;
wire wire35819;
wire wire35823;
wire wire35830;
wire wire35833;
wire wire35834;
wire wire35836;
wire wire35837;
wire wire35838;
wire wire35839;
wire wire35840;
wire wire35841;
wire wire35844;
wire wire35845;
wire wire35860;
wire wire35862;
wire wire35864;
wire wire35866;
wire wire35867;
wire wire35872;
wire wire35873;
wire wire35874;
wire wire35875;
wire wire35876;
wire wire35877;
wire wire35884;
wire wire35886;
wire wire35895;
wire wire35900;
wire wire35901;
wire wire35902;
wire wire35903;
wire wire35904;
wire wire35905;
wire wire35906;
wire wire35907;
wire wire35908;
wire wire35909;
wire wire35910;
wire wire35911;
wire wire35912;
wire wire35913;
wire wire35915;
wire wire35917;
wire wire35918;
wire wire35920;
wire wire35927;
wire wire35929;
wire wire35931;
wire wire35932;
wire wire35933;
wire wire35934;
wire wire35937;
wire wire35939;
wire wire35941;
wire wire35943;
wire wire35944;
wire wire35945;
wire wire35946;
wire wire35947;
wire wire35948;
wire wire35949;
wire wire35950;
wire wire35952;
wire wire35953;
wire wire35957;
wire wire35961;
wire wire35964;
wire wire35965;
wire wire35966;
wire wire35967;
wire wire35968;
wire wire35969;
wire wire35970;
wire wire35971;
wire wire35972;
wire wire35973;
wire wire35974;
wire wire35975;
wire wire35976;
wire wire35977;
wire wire35978;
wire wire35979;
wire wire35980;
wire wire35981;
wire wire35982;
wire wire35983;
wire wire35984;
wire wire35985;
wire wire35986;
wire wire35987;
wire wire35988;
wire wire35989;
wire wire35990;
wire wire35991;
wire wire35992;
wire wire35993;
wire wire35994;
wire wire35995;
wire wire35996;
wire wire35997;
wire wire35998;
wire wire35999;
wire wire36000;
wire wire36001;
wire wire36002;
wire wire36003;
wire wire36004;
wire wire36005;
wire wire36006;
wire wire36007;
wire wire36008;
wire wire36009;
wire wire36010;
wire wire36011;
wire wire36012;
wire wire36013;
wire wire36014;
wire wire36019;
wire wire36020;
wire wire36021;
wire wire36022;
wire wire36023;
wire wire36024;
wire wire36025;
wire wire36026;
wire wire36027;
wire wire36028;
wire wire36029;
wire wire36030;
wire wire36031;
wire wire36032;
wire wire36039;
wire wire36040;
wire wire36041;
wire wire36042;
wire wire36045;
wire wire36047;
wire wire36048;
wire wire36050;
wire wire36054;
wire wire36055;
wire wire36057;
wire wire36058;
wire wire36064;
wire wire36065;
wire wire36077;
wire wire36078;
wire wire36081;
wire wire36082;
wire wire36083;
wire wire36084;
wire wire36086;
wire wire36089;
wire wire36090;
wire wire36091;
wire wire36093;
wire wire36095;
wire wire36096;
wire wire36097;
wire wire36098;
wire wire36109;
wire wire36110;
wire wire36111;
wire wire36115;
wire wire36116;
wire wire36119;
wire wire36120;
wire wire36121;
wire wire36122;
wire wire36131;
wire wire36132;
wire wire36135;
wire wire36136;
wire wire36139;
wire wire36140;
wire wire36142;
wire wire36144;
wire wire36145;
wire wire36146;
wire wire36147;
wire wire36148;
wire wire36150;
wire wire36151;
wire wire36160;
wire wire36162;
wire wire36170;
wire wire36171;
wire wire36172;
wire wire36173;
wire wire36175;
wire wire36176;
wire wire36177;
wire wire36183;
wire wire36184;
wire wire36188;
wire wire36189;
wire wire36190;
wire wire36192;
wire wire36193;
wire wire36198;
wire wire36201;
wire wire36202;
wire wire36203;
wire wire36204;
wire wire36205;
wire wire36206;
wire wire36207;
wire wire36208;
wire wire36209;
wire wire36210;
wire wire36211;
wire wire36212;
wire wire36213;
wire wire36214;
wire wire36215;
wire wire36216;
wire wire36217;
wire wire36218;
wire wire36219;
wire wire36220;
wire wire36221;
wire wire36222;
wire wire36223;
wire wire36224;
wire wire36225;
wire wire36226;
wire wire36227;
wire wire36228;
wire wire36229;
wire wire36230;
wire wire36231;
wire wire36232;
wire wire36233;
wire wire36234;
wire wire36235;
wire wire36236;
wire wire36237;
wire wire36238;
wire wire36239;
wire wire36240;
wire wire36241;
wire wire36242;
wire wire36243;
wire wire36244;
wire wire36245;
wire wire36246;
wire wire36247;
wire wire36248;
wire wire36249;
wire wire36250;
wire wire36251;
wire wire36256;
wire wire36257;
wire wire36258;
wire wire36259;
wire wire36260;
wire wire36261;
wire wire36262;
wire wire36263;
wire wire36264;
wire wire36265;
wire wire36266;
wire wire36267;
wire wire36268;
wire wire36269;
wire wire36276;
wire wire36277;
wire wire36278;
wire wire36279;
wire wire36284;
wire wire36287;
wire wire36288;
wire wire36289;
wire wire36290;
wire wire36297;
wire wire36302;
wire wire36303;
wire wire36304;
wire wire36305;
wire wire36306;
wire wire36307;
wire wire36311;
wire wire36312;
wire wire36314;
wire wire36321;
wire wire36323;
wire wire36324;
wire wire36325;
wire wire36326;
wire wire36327;
wire wire36330;
wire wire36331;
wire wire36334;
wire wire36335;
wire wire36342;
wire wire36344;
wire wire36346;
wire wire36347;
wire wire36348;
wire wire36349;
wire wire36352;
wire wire36353;
wire wire36356;
wire wire36357;
wire wire36362;
wire wire36364;
wire wire36369;
wire wire36370;
wire wire36377;
wire wire36378;
wire wire36379;
wire wire36380;
wire wire36381;
wire wire36382;
wire wire36383;
wire wire36385;
wire wire36386;
wire wire36387;
wire wire36388;
wire wire36389;
wire wire36390;
wire wire36391;
wire wire36412;
wire wire36413;
wire wire36414;
wire wire36415;
wire wire36416;
wire wire36417;
wire wire36418;
wire wire36419;
wire wire36420;
wire wire36426;
wire wire36427;
wire wire36428;
wire wire36431;
wire wire36433;
wire wire36435;
wire wire36437;
wire wire36438;
wire wire36439;
wire wire36440;
wire wire36445;
wire wire36446;
wire wire36455;
wire wire36456;
wire wire36457;
wire wire36458;
wire wire36459;
wire wire36461;
wire wire36462;
wire wire36463;
wire wire36465;
wire wire36474;
wire wire36476;
reg ng3097;

reg ng3108;

reg ng3185;

reg ng3135;

reg ng141;

reg ng155;

reg ng258;

reg ng83;

reg ng369;

reg ng414;

reg ng441;

reg ng318;

reg ng452;

reg ng380;

reg ng557;

reg ng574;

reg ng461;

reg ng535;

reg ng575;

reg ng590;

reg ng490;

reg ng646;

reg ng703;

reg ng714;

reg ng722;

reg ng736;

reg ng821;

reg ng835;

reg ng849;

reg ng863;

reg ng924;

reg ng939;

reg ng954;

reg ng744;

reg ng1085;

reg ng1113;

reg ng1000;

reg ng1090;

reg ng969;

reg ng992;

reg ng1053;

reg ng1082;

reg ng1255;

reg ng1173;

reg ng1151;

reg ng1186;

reg ng1267;

reg ng1303;

reg ng1211;

reg ng1352;

reg ng1392;

reg ng1403;

reg ng1411;

reg ng1425;

reg ng1527;

reg ng1535;

reg ng1552;

reg ng1642;

reg ng1453;

reg ng1739;

reg ng1798;

reg ng1825;

reg ng1700;

reg ng1834;

reg ng1890;

reg ng1945;

reg ng1858;

reg ng1922;

reg ng1959;

reg ng1973;

reg ng1991;

reg ng1912;

reg ng2033;

reg ng2082;

reg ng2090;

reg ng2104;

reg ng2237;

reg ng2251;

reg ng2312;

reg ng2327;

reg ng2342;

reg ng2124;

reg ng2436;

reg ng2495;

reg ng2523;

reg ng2362;

reg ng2426;

reg ng2455;

reg ng2631;

reg ng2648;

reg ng2536;

reg ng2609;

reg ng2649;

reg ng2772;

reg ng2786;

reg ng2797;

reg ng2805;

reg ng3044;

reg ng3098;

reg ng3107;

reg ng3088;

reg ng3139;

reg ng145;

reg ng154;

reg ng261;

reg ng88;

reg ng358;

reg ng411;

reg ng444;

reg ng317;

reg ng286;

reg ng381;

reg ng554;

reg ng565;

reg ng458;

reg ng542;

reg ng577;

reg ng593;

reg ng611;

reg ng660;

reg ng702;

reg ng715;

reg ng724;

reg ng734;

reg ng817;

reg ng839;

reg ng848;

reg ng921;

reg ng882;

reg ng936;

reg ng957;

reg ng749;

reg ng1075;

reg ng1115;

reg ng1001;

reg ng1008;

reg ng970;

reg ng986;

reg ng985;

reg ng1083;

reg ng1250;

reg ng1174;

reg ng1171;

reg ng1244;

reg ng1269;

reg ng1306;

reg pg16355;

reg ng1365;

reg ng1391;

reg ng1404;

reg ng1413;

reg ng1423;

reg ng1523;

reg ng1539;

reg ng1551;

reg ng1585;

reg ng1448;

reg ng1750;

reg ng1801;

reg ng1822;

reg ng1701;

reg ng1833;

reg ng1893;

reg ng1954;

reg ng1859;

reg ng1915;

reg ng1960;

reg ng1970;

reg ng1871;

reg ng1911;

reg ng2026;

reg ng2078;

reg ng2094;

reg ng2103;

reg ng2235;

reg ng2247;

reg ng2270;

reg ng2324;

reg ng2345;

reg ng2129;

reg ng2459;

reg ng2492;

reg ng2394;

reg ng2363;

reg ng2425;

reg ng2456;

reg ng2628;

reg ng2639;

reg ng2533;

reg ng2616;

reg ng2651;

reg ng2727;

reg ng2784;

reg ng2793;

reg ng2809;

reg ng3043;

reg ng3099;

reg ng3158;

reg ng3179;

reg ng3110;

reg ng164;

reg ng178;

reg ng264;

reg ng74;

reg ng343;

reg ng408;

reg ng448;

reg ng450;

reg ng285;

reg ng382;

reg ng513;

reg ng572;

reg ng455;

reg ng543;

reg ng580;

reg ng584;

reg ng608;

reg ng672;

reg ng705;

reg ng712;

reg ng723;

reg ng738;

reg ng820;

reg ng836;

reg ng844;

reg ng885;

reg ng900;

reg ng912;

reg ng753;

reg ng1078;

reg ng1119;

reg ng1134;

reg ng1010;

reg ng1029;

reg ng1055;

reg ng1210;

reg ng1175;

reg ng1155;

reg ng1234;

reg ng1268;

reg ng1291;

reg ng1216;

reg ng1315;

reg ng1402;

reg ng1416;

reg ng1420;

reg ng1525;

reg ng1540;

reg ng1554;

reg ng1573;

reg ng1444;

reg ng1765;

reg ng1792;

reg ng1819;

reg ng1703;

reg ng1660;

reg ng1903;

reg ng1947;

reg ng1839;

reg ng1908;

reg ng1958;

reg ng1979;

reg ng1874;

reg ng1914;

reg ng2020;

reg ng2080;

reg ng2113;

reg ng2209;

reg ng2239;

reg ng2250;

reg ng2306;

reg ng2285;

reg ng2348;

reg ng2256;

reg ng2444;

reg ng2489;

reg ng2395;

reg ng2529;

reg ng2457;

reg ng2587;

reg ng2646;

reg ng2530;

reg ng2617;

reg ng2654;

reg ng2720;

reg ng2777;

reg ng2795;

reg ng2810;

reg ng3046;

reg ng3100;

reg ng3155;

reg ng3182;

reg ng3120;

reg ng162;

reg ng174;

reg ng222;

reg ng79;

reg ng346;

reg ng391;

reg ng319;

reg ng451;

reg ng284;

reg ng383;

reg ng510;

reg ng573;

reg ng488;

reg ng544;

reg ng579;

reg ng587;

reg ng605;

reg ng666;

reg ng701;

reg ng710;

reg ng719;

reg ng739;

reg ng822;

reg ng837;

reg ng846;

reg ng888;

reg ng942;

reg ng915;

reg ng758;

reg ng1095;

reg ng1116;

reg ng999;

reg ng1009;

reg ng1036;

reg ng1054;

reg ng1081;

reg ng1142;

reg ng1152;

reg ng1235;

reg ng1264;

reg ng1215;

reg ng1217;

reg ng1312;

reg ng1406;

reg ng1415;

reg ng1424;

reg ng1524;

reg ng1538;

reg ng1550;

reg ng1555;

reg ng1439;

reg ng1742;

reg ng1795;

reg ng1816;

reg ng1704;

reg ng1835;

reg ng1904;

reg ng1946;

reg ng1842;

reg ng1852;

reg ng1962;

reg ng1976;

reg ng1877;

reg ng1913;

reg ng2013;

reg ng2079;

reg ng2111;

reg ng2205;

reg ng2240;

reg ng2252;

reg ng2309;

reg ng2282;

reg ng2160;

reg ng2120;

reg ng2433;

reg ng2486;

reg ng2397;

reg ng2528;

reg ng2458;

reg ng2584;

reg ng2647;

reg ng2563;

reg ng2618;

reg ng2653;

reg ng2734;

reg ng2776;

reg ng2785;

reg ng2808;

reg ng3045;

reg ng2900;

reg ng3093;

reg ng3104;

reg ng3173;

reg ng3123;

reg ng195;

reg ng255;

reg ng270;

reg ng52;

reg ng388;

reg ng298;

reg ng367;

reg ng570;

reg ng487;

reg ng529;

reg ng659;

reg ng721;

reg ng737;

reg ng856;

reg ng876;

reg ng1098;

reg ng1125;

reg ng1141;

reg ng976;

reg ng1145;

reg ng1214;

reg ng1263;

reg ng1282;

reg ng1183;

reg ng1407;

reg ng1418;

reg ng1511;

reg ng1531;

reg ng1534;

reg ng1545;

reg ng1435;

reg ng1757;

reg ng1809;

reg ng1693;

reg ng1696;

reg ng1783;

reg ng1944;

reg ng1870;

reg ng1865;

reg ng1929;

reg ng1939;

reg ng1966;

reg ng1886;

reg ng1917;

reg ng2089;

reg ng2100;

reg ng2108;

reg ng2207;

reg ng2238;

reg ng2255;

reg ng2315;

reg ng2294;

reg ng2339;

reg ng2142;

reg ng2418;

reg ng2483;

reg ng2398;

reg ng2355;

reg ng2366;

reg ng2439;

reg ng2644;

reg ng2562;

reg ng2670;

reg ng2571;

reg ng2610;

reg ng2812;

reg ng3048;

reg ng3094;

reg ng3103;

reg ng3176;

reg ng3124;

reg ng198;

reg ng252;

reg ng213;

reg ng354;

reg ng398;

reg ng342;

reg ng366;

reg ng571;

reg ng486;

reg ng530;

reg ng630;

reg ng711;

reg ng830;

reg ng860;

reg ng873;

reg ng1101;

reg ng1122;

reg ng966;

reg ng975;

reg ng1148;

reg ng1158;

reg ng1270;

reg ng1285;

reg ng1180;

reg ng1405;

reg ng1414;

reg ng1515;

reg ng1530;

reg ng1532;

reg ng1541;

reg ng1430;

reg ng1754;

reg ng1807;

reg ng1828;

reg ng1697;

reg ng1785;

reg ng1949;

reg ng1948;

reg ng1845;

reg ng1928;

reg ng1956;

reg ng1965;

reg ng1887;

reg ng1916;

reg ng2087;

reg ng2096;

reg ng2112;

reg ng2206;

reg ng2245;

reg ng2254;

reg ng2318;

reg ng2291;

reg ng2297;

reg ng2147;

reg ng2421;

reg ng2466;

reg ng2396;

reg ng2354;

reg ng2374;

reg ng2432;

reg ng2645;

reg ng2561;

reg ng2652;

reg ng2580;

reg ng2608;

reg ng2813;

reg ng3047;

reg ng3095;

reg ng3106;

reg ng3167;

reg ng3125;

reg ng216;

reg ng92;

reg ng376;

reg ng349;

reg ng372;

reg ng324;

reg ng531;

reg ng633;

reg ng698;

reg ng840;

reg ng861;

reg ng918;

reg ng1002;

reg ng1089;

reg ng967;

reg ng978;

reg ng1164;

reg ng1245;

reg ng1272;

reg ng1288;

reg ng1193;

reg ng1409;

reg ng1417;

reg ng1512;

reg ng1526;

reg ng1536;

reg ng1544;

reg ng1426;

reg ng1769;

reg ng1804;

reg ng1830;

reg ng1698;

reg ng1832;

reg ng1950;

reg ng1868;

reg ng1860;

reg ng1924;

reg ng1957;

reg ng1967;

reg ng2040;

reg ng2081;

reg ng2091;

reg ng2099;

reg ng2109;

reg ng2117;

reg ng2246;

reg ng2261;

reg ng2273;

reg ng2288;

reg ng2300;

reg ng2133;

reg ng2463;

reg ng2478;

reg ng2357;

reg ng2364;

reg ng2428;

reg ng2447;

reg ng2399;

reg ng2656;

reg ng2676;

reg ng2607;

reg ng2811;

reg ng3096;

reg ng3105;

reg ng3170;

reg ng3126;

reg ng219;

reg ng273;

reg ng56;

reg ng368;

reg ng379;

reg ng397;

reg ng532;

reg ng640;

reg ng653;

reg ng847;

reg ng859;

reg ng879;

reg ng1003;

reg ng1091;

reg ng968;

reg ng977;

reg ng1221;

reg ng1262;

reg ng1271;

reg ng1300;

reg ng1192;

reg ng1410;

reg ng1419;

reg ng1513;

reg ng1528;

reg ng1537;

reg ng1546;

reg ng1735;

reg ng1779;

reg ng1808;

reg ng1829;

reg ng1699;

reg ng1831;

reg ng1951;

reg ng1867;

reg ng1861;

reg ng1923;

reg ng1955;

reg ng1964;

reg ng2052;

reg ng2083;

reg ng2092;

reg ng2101;

reg ng2110;

reg ng2119;

reg ng2244;

reg ng2253;

reg ng2276;

reg ng2330;

reg ng2303;

reg ng2138;

reg ng2429;

reg ng2473;

reg ng2479;

reg ng2356;

reg ng2365;

reg ng2427;

reg ng2454;

reg ng2472;

reg ng2657;

reg ng2673;

reg ng2568;

reg ng3049;

reg ng2888;

reg ng130;

reg ng144;

reg ng158;

reg ng172;

reg ng192;

reg ng207;

reg ng449;

reg ng322;

reg ng279;

reg ng290;

reg ng357;

reg ng578;

reg ng599;

reg ng506;

reg ng537;

reg ng700;

reg ng838;

reg ng852;

reg ng866;

reg ng894;

reg ng909;

reg ng1137;

reg ng972;

reg ng1044;

reg ng1070;

reg ng1209;

reg ng1294;

reg ng1223;

reg ng1332;

reg ng1389;

reg ng1400;

reg ng1560;

reg ng1582;

reg ng1597;

reg ng1466;

reg ng1666;

reg ng1730;

reg ng1753;

reg ng1705;

reg ng2217;

reg ng2231;

reg ng2248;

reg ng2503;

reg ng2387;

reg ng2477;

reg ng2359;

reg ng2417;

reg ng2443;

reg ng2655;

reg ng2691;

reg ng2599;

reg ng2704;

reg ng2766;

reg ng2783;

reg ng2794;

reg ng3050;

reg ng3062;

reg ng3073;

reg ng3013;

reg pg8274;

reg pg8265;

reg ng2896;

reg ng131;

reg ng146;

reg ng156;

reg ng168;

reg ng231;

reg ng204;

reg ng427;

reg ng323;

reg ng454;

reg ng291;

reg ng353;

reg ng582;

reg ng596;

reg ng507;

reg ng536;

reg ng707;

reg ng831;

reg ng850;

reg ng862;

reg ng897;

reg ng951;

reg ng1138;

reg ng971;

reg ng1051;

reg ng1069;

reg ng1252;

reg ng1273;

reg ng1224;

reg ng1339;

reg ng1387;

reg ng1396;

reg ng1561;

reg ng1579;

reg ng1600;

reg ng1654;

reg ng1667;

reg ng1723;

reg ng1760;

reg ng1778;

reg ng2221;

reg ng2230;

reg ng2264;

reg ng2501;

reg ng2522;

reg ng2525;

reg ng2358;

reg ng2424;

reg ng2442;

reg ng2659;

reg ng2688;

reg ng2603;

reg ng2615;

reg ng2773;

reg ng2782;

reg ng2804;

reg ng3051;

reg ng3061;

reg ng3074;

reg ng3002;

reg pg8273;

reg pg8266;

reg ng2892;

reg ng129;

reg ng149;

reg ng153;

reg ng170;

reg ng234;

reg ng249;

reg ng428;

reg ng312;

reg ng453;

reg ng299;

reg ng365;

reg ng484;

reg ng549;

reg pg16297;

reg ng541;

reg ng720;

reg ng826;

reg ng857;

reg ng865;

reg ng767;

reg ng1045;

reg ng1139;

reg ng974;

reg ng1052;

reg ng1196;

reg ng1251;

reg ng1276;

reg ng1177;

reg ng1227;

reg ng1358;

reg ng1384;

reg ng1398;

reg ng1529;

reg ng1543;

reg ng1559;

reg ng1624;

reg ng1636;

reg ng1651;

reg ng1784;

reg ng1668;

reg ng1732;

reg ng1748;

reg ng1777;

reg ng2222;

reg ng2233;

reg ng2321;

reg ng2504;

reg ng2389;

reg ng2526;

reg ng2361;

reg ng2380;

reg ng2441;

reg ng2559;

reg ng2623;

reg ng2660;

reg ng2679;

reg ng2581;

reg ng2612;

reg ng2774;

reg ng2792;

reg ng2803;

reg ng3052;

reg ng3064;

reg ng3071;

reg ng3006;

reg pg8272;

reg pg8262;

reg pg8258;

reg ng2903;

reg ng133;

reg ng148;

reg ng157;

reg ng169;

reg ng237;

reg ng210;

reg ng426;

reg ng447;

reg ng320;

reg ng305;

reg ng364;

reg ng464;

reg ng548;

reg ng525;

reg ng538;

reg ng730;

reg ng728;

reg ng858;

reg ng867;

reg ng762;

reg ng1056;

reg ng1140;

reg ng973;

reg ng1074;

reg ng1199;

reg ng1260;

reg ng1279;

reg ng1297;

reg ng1309;

reg ng1346;

reg ng1388;

reg ng1397;

reg ng1533;

reg ng1542;

reg ng1567;

reg ng1621;

reg ng1594;

reg ng1648;

reg ng1695;

reg ng1669;

reg ng1731;

reg ng1749;

reg ng1776;

reg ng2220;

reg ng2229;

reg ng2333;

reg ng2507;

reg ng2388;

reg ng2527;

reg ng2360;

reg ng2373;

reg ng2440;

reg ng2539;

reg ng2622;

reg ng2658;

reg ng2694;

reg pg16437;

reg ng2611;

reg ng2781;

reg ng2790;

reg ng2799;

reg ng3053;

reg ng3063;

reg ng3072;

reg ng2998;

reg pg8268;

reg pg8264;

reg ng2817;

reg ng3101;

reg ng3164;

reg ng134;

reg ng151;

reg ng159;

reg ng176;

reg ng179;

reg ng240;

reg ng225;

reg ng65;

reg ng373;

reg ng429;

reg ng314;

reg ng404;

reg ng283;

reg ng350;

reg ng387;

reg ng524;

reg ng568;

reg ng480;

reg ng465;

reg ng558;

reg ng585;

reg ng620;

reg ng679;

reg ng704;

reg ng718;

reg ng729;

reg ng732;

reg ng853;

reg ng834;

reg ng845;

reg ng927;

reg ng906;

reg ng776;

reg ng1033;

reg ng1048;

reg ng1107;

reg ng1135;

reg ng1007;

reg ng1037;

reg ng1066;

reg ng1240;

reg ng1259;

reg ng1165;

reg ng1229;

reg ng1266;

reg ng1218;

reg ng1345;

reg ng1385;

reg ng1393;

reg ng1421;

reg ng1514;

reg ng1553;

reg ng1615;

reg ng1630;

reg ng1609;

reg ng1813;

reg ng1662;

reg ng1680;

reg ng1746;

reg ng1775;

reg ng2224;

reg ng2232;

reg ng2156;

reg ng2510;

reg ng2391;

reg ng2462;

reg ng2598;

reg ng2642;

reg ng2555;

reg ng2540;

reg ng2632;

reg ng2661;

reg ng2685;

reg ng2606;

reg ng2746;

reg ng2779;

reg ng2787;

reg ng2801;

reg ng3054;

reg ng3055;

reg ng3066;

reg ng3077;

reg ng3028;

reg pg5388;

reg ng3083;

reg ng2990;

reg ng2933;

reg ng3102;

reg ng3161;

reg ng132;

reg ng147;

reg ng163;

reg ng175;

reg ng177;

reg ng201;

reg ng228;

reg ng70;

reg ng423;

reg ng432;

reg ng313;

reg ng402;

reg ng282;

reg ng287;

reg ng394;

reg ng523;

reg ng489;

reg ng479;

reg ng468;

reg ng499;

reg ng586;

reg ng617;

reg ng686;

reg ng706;

reg ng716;

reg ng725;

reg ng733;

reg ng823;

reg ng832;

reg ng841;

reg ng930;

reg ng903;

reg ng771;

reg ng1030;

reg ng1071;

reg ng1104;

reg ng1136;

reg ng1006;

reg ng1038;

reg ng1059;

reg ng1243;

reg ng1258;

reg ng1253;

reg ng1230;

reg ng1265;

reg ng1219;

reg ng1316;

reg ng1386;

reg ng1395;

reg ng1422;

reg ng1516;

reg ng1557;

reg ng1612;

reg ng1633;

reg ng1606;

reg ng1789;

reg ng1663;

reg ng1672;

reg ng1747;

reg ng1768;

reg ng2225;

reg ng2234;

reg ng2258;

reg ng2513;

reg ng2390;

reg ng2469;

reg ng2597;

reg ng2564;

reg ng2554;

reg ng2543;

reg ng2574;

reg ng2664;

reg ng2682;

reg ng2707;

reg ng2740;

reg ng2775;

reg ng2791;

reg ng2800;

reg ng2802;

reg ng3056;

reg ng3065;

reg ng3078;

reg ng3018;

reg ng2986;

reg pg8271;

reg ng2991;

reg ng2950;

reg ng3191;

reg ng185;

reg ng142;

reg ng150;

reg ng160;

reg ng171;

reg ng186;

reg ng246;

reg ng267;

reg ng361;

reg ng420;

reg ng435;

reg ng316;

reg ng321;

reg ng281;

reg ng288;

reg ng352;

reg ng395;

reg ng569;

reg ng566;

reg ng478;

reg ng471;

reg ng576;

reg ng583;

reg ng614;

reg ng493;

reg ng534;

reg ng692;

reg ng709;

reg ng713;

reg ng727;

reg ng731;

reg ng819;

reg ng829;

reg ng843;

reg ng864;

reg ng933;

reg ng948;

reg ng960;

reg ng1041;

reg ng1060;

reg ng1114;

reg ng1128;

reg ng1005;

reg ng1039;

reg ng1068;

reg ng1084;

reg ng1257;

reg ng1254;

reg ng1167;

reg ng1261;

reg ng1220;

reg ng1319;

reg ng1372;

reg ng1394;

reg ng1401;

reg ng1412;

reg ng1558;

reg ng1576;

reg ng1588;

reg ng1603;

reg ng1727;

reg ng1664;

reg ng1679;

reg ng1738;

reg ng1764;

reg ng2448;

reg ng2516;

reg ng2393;

reg ng2470;

reg ng2643;

reg ng2640;

reg ng2553;

reg ng2546;

reg ng2650;

reg ng2667;

reg ng2604;

reg ng2714;

reg ng2753;

reg ng2778;

reg ng2788;

reg ng2796;

reg ng2806;

reg ng3080;

reg ng3057;

reg ng3068;

reg ng3075;

reg ng3024;

reg ng2987;

reg ng2992;

reg pg8261;

reg ng2883;

reg ng3128;

reg ng3147;

reg ng143;

reg ng152;

reg ng161;

reg ng173;

reg ng189;

reg ng243;

reg ng61;

reg ng384;

reg ng417;

reg ng438;

reg ng315;

reg ng403;

reg ng280;

reg ng289;

reg ng351;

reg ng396;

reg ng564;

reg ng567;

reg ng477;

reg ng528;

reg ng559;

reg ng581;

reg ng602;

reg ng496;

reg ng533;

reg ng699;

reg ng708;

reg ng717;

reg ng726;

reg ng735;

reg ng818;

reg ng833;

reg ng842;

reg ng851;

reg ng891;

reg ng945;

reg ng780;

reg ng740;

reg ng1063;

reg ng1110;

reg ng1131;

reg ng1004;

reg ng1040;

reg ng1067;

reg ng1011;

reg ng1256;

reg ng1176;

reg ng1166;

reg ng1228;

reg ng1222;

reg ng1326;

reg ng1378;

reg ng1390;

reg ng1399;

reg ng1408;

reg ng1556;

reg ng1618;

reg ng1591;

reg ng1645;

reg ng1457;

reg ng1665;

reg ng1686;

reg ng1745;

reg ng1763;

reg ng2498;

reg ng2519;

reg ng2392;

reg ng2471;

reg ng2638;

reg ng2641;

reg ng2552;

reg ng2602;

reg ng2633;

reg ng2565;

reg ng2605;

reg ng2733;

reg ng2760;

reg ng2780;

reg ng2789;

reg ng2798;

reg ng2807;

reg ng3079;

reg ng3058;

reg ng3067;

reg ng3076;

reg ng3010;

reg pg8275;

reg pg8267;

reg pg8259;

reg ng809;

reg pg7334;

reg ng113;

reg ng2200;

reg ng3084;

reg ng3059;

reg ng3070;

reg pg4323;

reg ng789;

reg pg8175;

reg ng2857;

reg ng3085;

reg ng3060;

reg ng3069;

reg ng805;

reg pg7519;

reg ng117;

reg pg8096;

reg ng3086;

reg ng2997;

reg ng3032;

reg pg8021;

reg pg4590;

reg ng785;

reg pg8023;

reg ng97;

reg ng3087;

reg ng2993;

reg ng3036;

reg ng2908;

reg ng2935;

reg ng2969;

reg ng1481;

reg ng3091;

reg ng1570;

reg ng1670;

reg ng1734;

reg ng2210;

reg ng2227;

reg pg8269;

reg pg8260;

reg ng2912;

reg ng2934;

reg ng2972;

reg ng1486;

reg ng3092;

reg ng1627;

reg ng1671;

reg ng1733;

reg ng2208;

reg ng2223;

reg pg8270;

reg pg8263;

reg ng2917;

reg ng2941;

reg ng2963;

reg ng1491;

reg ng1639;

reg ng1761;

reg ng1937;

reg ng2218;

reg ng2226;

reg ng2524;

reg ng2924;

reg ng2938;

reg ng2966;

reg ng1496;

reg ng1462;

reg ng1762;

reg ng1934;

reg ng2219;

reg ng2228;

reg ng2502;

reg ng2920;

reg ng2947;

reg ng2981;

reg pg8251;

reg ng793;

reg pg4321;

reg ng1724;

reg ng1952;

reg ng1836;

reg ng2085;

reg ng2093;

reg ng2107;

reg ng2118;

reg ng2451;

reg ng2984;

reg ng2944;

reg ng2874;

reg ng2877;

reg pg6895;

reg ng121;

reg ng1772;

reg ng1953;

reg ng1869;

reg ng2086;

reg ng2095;

reg ng2105;

reg ng2114;

reg ng2257;

reg ng2985;

reg ng2956;

reg ng2975;

reg ng1471;

reg ng101;

reg ng2170;

reg ng1810;

reg ng1846;

reg ng1938;

reg ng2084;

reg ng2098;

reg ng2102;

reg ng2116;

reg ng2151;

reg ng2953;

reg ng2978;

reg ng1476;

reg pg4450;

reg ng2175;

reg ng1694;

reg ng1849;

reg ng1880;

reg ng2088;

reg ng2097;

reg ng2106;

reg ng2115;

reg ng2336;

reg ng2929;

reg ng2962;

reg ng801;

reg pg8249;

reg ng105;

reg ng2180;

reg ng2165;

reg ng1702;

reg ng1963;

reg ng1994;

reg ng1997;

reg ng1905;

reg ng2010;

reg ng2072;

reg ng2279;

reg ng2879;

reg ng2959;

reg pg6225;

reg ng2873;

reg pg4200;

reg ng2185;

reg ng2878;

reg ng1661;

reg ng1961;

reg ng1982;

reg ng2000;

reg pg16399;

reg ng2039;

reg ng2066;

reg ng2267;

reg ng1506;

reg pg4090;

reg ng797;

reg pg4088;

reg ng109;

reg ng2190;

reg ng3210;

reg ng1985;

reg ng1910;

reg ng1918;

reg ng2059;

reg ng2249;

reg ng1501;

reg ng813;

reg pg6442;

reg ng125;

reg pg3993;

reg ng2195;

reg ng3211;

reg ng1988;

reg ng1909;

reg ng1921;

reg ng2046;

reg ng2236;

always  @(posedge pclk)
	ng3097<=ng25450;

 always  @(posedge pclk)
	ng3108<=ng30801;

 always  @(posedge pclk)
	ng3185<=ng17341;

 always  @(posedge pclk)
	ng3135<=pg26149;

 always  @(posedge pclk)
	ng141<=ng22030;

 always  @(posedge pclk)
	ng155<=ng22064;

 always  @(posedge pclk)
	ng258<=ng30258;

 always  @(posedge pclk)
	ng83<=ng26529;

 always  @(posedge pclk)
	ng369<=ng27256;

 always  @(posedge pclk)
	ng414<=ng28744;

 always  @(posedge pclk)
	ng441<=ng26808;

 always  @(posedge pclk)
	ng318<=ng30455;

 always  @(posedge pclk)
	ng452<=ng11510;

 always  @(posedge pclk)
	ng380<=ng373;

 always  @(posedge pclk)
	ng557<=ng18678;

 always  @(posedge pclk)
	ng574<=ng465;

 always  @(posedge pclk)
	ng461<=ng24174;

 always  @(posedge pclk)
	ng535<=ng528;

 always  @(posedge pclk)
	ng575<=ng27279;

 always  @(posedge pclk)
	ng590<=ng24498;

 always  @(posedge pclk)
	ng490<=ng26541;

 always  @(posedge pclk)
	ng646<=ng24426;

 always  @(posedge pclk)
	ng703<=ng20892;

 always  @(posedge pclk)
	ng714<=ng20946;

 always  @(posedge pclk)
	ng722<=ng21051;

 always  @(posedge pclk)
	ng736<=ng25262;

 always  @(posedge pclk)
	ng821<=ng22146;

 always  @(posedge pclk)
	ng835<=ng22066;

 always  @(posedge pclk)
	ng849<=ng22128;

 always  @(posedge pclk)
	ng863<=ng25223;

 always  @(posedge pclk)
	ng924<=ng30654;

 always  @(posedge pclk)
	ng939<=ng30264;

 always  @(posedge pclk)
	ng954<=ng30670;

 always  @(posedge pclk)
	ng744<=ng29354;

 always  @(posedge pclk)
	ng1085<=ng27284;

 always  @(posedge pclk)
	ng1113<=ng28767;

 always  @(posedge pclk)
	ng1000<=ng29612;

 always  @(posedge pclk)
	ng1090<=ng26661;

 always  @(posedge pclk)
	ng969<=ng11519;

 always  @(posedge pclk)
	ng992<=ng26183;

 always  @(posedge pclk)
	ng1053<=ng1052;

 always  @(posedge pclk)
	ng1082<=ng1075;

 always  @(posedge pclk)
	ng1255<=ng1250;

 always  @(posedge pclk)
	ng1173<=ng23081;

 always  @(posedge pclk)
	ng1151<=ng23039;

 always  @(posedge pclk)
	ng1186<=ng1235;

 always  @(posedge pclk)
	ng1267<=ng27328;

 always  @(posedge pclk)
	ng1303<=ng28355;

 always  @(posedge pclk)
	ng1211<=pg16355;

 always  @(posedge pclk)
	ng1352<=ng26781;

 always  @(posedge pclk)
	ng1392<=ng20926;

 always  @(posedge pclk)
	ng1403<=ng20995;

 always  @(posedge pclk)
	ng1411<=ng20913;

 always  @(posedge pclk)
	ng1425<=ng22247;

 always  @(posedge pclk)
	ng1527<=ng22044;

 always  @(posedge pclk)
	ng1535<=ng22130;

 always  @(posedge pclk)
	ng1552<=ng25224;

 always  @(posedge pclk)
	ng1642<=ng30281;

 always  @(posedge pclk)
	ng1453<=ng27129;

 always  @(posedge pclk)
	ng1739<=ng27288;

 always  @(posedge pclk)
	ng1798<=ng29205;

 always  @(posedge pclk)
	ng1825<=ng26824;

 always  @(posedge pclk)
	ng1700<=ng30503;

 always  @(posedge pclk)
	ng1834<=ng1833;

 always  @(posedge pclk)
	ng1890<=ng18794;

 always  @(posedge pclk)
	ng1945<=ng1954;

 always  @(posedge pclk)
	ng1858<=ng24208;

 always  @(posedge pclk)
	ng1922<=ng1915;

 always  @(posedge pclk)
	ng1959<=ng27306;

 always  @(posedge pclk)
	ng1973<=ng24534;

 always  @(posedge pclk)
	ng1991<=ng28361;

 always  @(posedge pclk)
	ng1912<=ng13445;

 always  @(posedge pclk)
	ng2033<=ng23339;

 always  @(posedge pclk)
	ng2082<=ng20916;

 always  @(posedge pclk)
	ng2090<=ng21019;

 always  @(posedge pclk)
	ng2104<=ng21072;

 always  @(posedge pclk)
	ng2237<=ng22172;

 always  @(posedge pclk)
	ng2251<=ng25247;

 always  @(posedge pclk)
	ng2312<=ng30672;

 always  @(posedge pclk)
	ng2327<=ng30282;

 always  @(posedge pclk)
	ng2342<=ng30686;

 always  @(posedge pclk)
	ng2124<=ng29357;

 always  @(posedge pclk)
	ng2436<=ng27322;

 always  @(posedge pclk)
	ng2495<=ng29221;

 always  @(posedge pclk)
	ng2523<=ng27767;

 always  @(posedge pclk)
	ng2362<=ng2361;

 always  @(posedge pclk)
	ng2426<=ng2425;

 always  @(posedge pclk)
	ng2455<=ng2448;

 always  @(posedge pclk)
	ng2631<=ng18780;

 always  @(posedge pclk)
	ng2648<=ng2540;

 always  @(posedge pclk)
	ng2536<=ng24209;

 always  @(posedge pclk)
	ng2609<=ng2602;

 always  @(posedge pclk)
	ng2649<=ng27336;

 always  @(posedge pclk)
	ng2772<=ng20962;

 always  @(posedge pclk)
	ng2786<=ng21026;

 always  @(posedge pclk)
	ng2797<=ng21075;

 always  @(posedge pclk)
	ng2805<=ng21063;

 always  @(posedge pclk)
	ng3044<=ng29454;

 always  @(posedge pclk)
	ng3098<=ng25451;

 always  @(posedge pclk)
	ng3107<=ng30798;

 always  @(posedge pclk)
	ng3088<=ng17429;

 always  @(posedge pclk)
	ng3139<=pg27380;

 always  @(posedge pclk)
	ng145<=ng22028;

 always  @(posedge pclk)
	ng154<=ng22049;

 always  @(posedge pclk)
	ng261<=ng30263;

 always  @(posedge pclk)
	ng88<=ng25932;

 always  @(posedge pclk)
	ng358<=ng27259;

 always  @(posedge pclk)
	ng411<=ng28735;

 always  @(posedge pclk)
	ng444<=ng26812;

 always  @(posedge pclk)
	ng317<=ng30702;

 always  @(posedge pclk)
	ng286<=ng11494;

 always  @(posedge pclk)
	ng381<=ng380;

 always  @(posedge pclk)
	ng554<=ng21842;

 always  @(posedge pclk)
	ng565<=ng574;

 always  @(posedge pclk)
	ng458<=ng23399;

 always  @(posedge pclk)
	ng542<=ng535;

 always  @(posedge pclk)
	ng577<=ng27268;

 always  @(posedge pclk)
	ng593<=ng24507;

 always  @(posedge pclk)
	ng611<=ng28348;

 always  @(posedge pclk)
	ng660<=ng25185;

 always  @(posedge pclk)
	ng702<=ng20880;

 always  @(posedge pclk)
	ng715<=ng20967;

 always  @(posedge pclk)
	ng724<=ng21032;

 always  @(posedge pclk)
	ng734<=ng25266;

 always  @(posedge pclk)
	ng817<=ng22162;

 always  @(posedge pclk)
	ng839<=ng22056;

 always  @(posedge pclk)
	ng848<=ng22106;

 always  @(posedge pclk)
	ng921<=ng30648;

 always  @(posedge pclk)
	ng882<=ng30676;

 always  @(posedge pclk)
	ng936<=ng30259;

 always  @(posedge pclk)
	ng957<=ng30677;

 always  @(posedge pclk)
	ng749<=ng29110;

 always  @(posedge pclk)
	ng1075<=ng27298;

 always  @(posedge pclk)
	ng1115<=ng28759;

 always  @(posedge pclk)
	ng1001<=ng29616;

 always  @(posedge pclk)
	ng1008<=ng29179;

 always  @(posedge pclk)
	ng970<=ng969;

 always  @(posedge pclk)
	ng986<=ng19024;

 always  @(posedge pclk)
	ng985<=ng26120;

 always  @(posedge pclk)
	ng1083<=ng1082;

 always  @(posedge pclk)
	ng1250<=ng1142;

 always  @(posedge pclk)
	ng1174<=ng23111;

 always  @(posedge pclk)
	ng1171<=ng23014;

 always  @(posedge pclk)
	ng1244<=ng13171;

 always  @(posedge pclk)
	ng1269<=ng27315;

 always  @(posedge pclk)
	ng1306<=ng28360;

 always  @(posedge pclk)
	pg16355<=ng26272;

 always  @(posedge pclk)
	ng1365<=ng27678;

 always  @(posedge pclk)
	ng1391<=ng20912;

 always  @(posedge pclk)
	ng1404<=ng21016;

 always  @(posedge pclk)
	ng1413<=ng20898;

 always  @(posedge pclk)
	ng1423<=ng22263;

 always  @(posedge pclk)
	ng1523<=ng22057;

 always  @(posedge pclk)
	ng1539<=ng22114;

 always  @(posedge pclk)
	ng1551<=ng25217;

 always  @(posedge pclk)
	ng1585<=ng30295;

 always  @(posedge pclk)
	ng1448<=ng27612;

 always  @(posedge pclk)
	ng1750<=ng27275;

 always  @(posedge pclk)
	ng1801<=ng29212;

 always  @(posedge pclk)
	ng1822<=ng26821;

 always  @(posedge pclk)
	ng1701<=ng30338;

 always  @(posedge pclk)
	ng1833<=ng11564;

 always  @(posedge pclk)
	ng1893<=ng12524;

 always  @(posedge pclk)
	ng1954<=ng1846;

 always  @(posedge pclk)
	ng1859<=ng24219;

 always  @(posedge pclk)
	ng1915<=ng1908;

 always  @(posedge pclk)
	ng1960<=ng27320;

 always  @(posedge pclk)
	ng1970<=ng24524;

 always  @(posedge pclk)
	ng1871<=ng26559;

 always  @(posedge pclk)
	ng1911<=ng13444;

 always  @(posedge pclk)
	ng2026<=ng24434;

 always  @(posedge pclk)
	ng2078<=ng20934;

 always  @(posedge pclk)
	ng2094<=ng21001;

 always  @(posedge pclk)
	ng2103<=ng21056;

 always  @(posedge pclk)
	ng2235<=ng22184;

 always  @(posedge pclk)
	ng2247<=ng25251;

 always  @(posedge pclk)
	ng2270<=ng30690;

 always  @(posedge pclk)
	ng2324<=ng30274;

 always  @(posedge pclk)
	ng2345<=ng30691;

 always  @(posedge pclk)
	ng2129<=ng29112;

 always  @(posedge pclk)
	ng2459<=ng27309;

 always  @(posedge pclk)
	ng2492<=ng29213;

 always  @(posedge pclk)
	ng2394<=ng30341;

 always  @(posedge pclk)
	ng2363<=ng11576;

 always  @(posedge pclk)
	ng2425<=ng2418;

 always  @(posedge pclk)
	ng2456<=ng2455;

 always  @(posedge pclk)
	ng2628<=ng21847;

 always  @(posedge pclk)
	ng2639<=ng2648;

 always  @(posedge pclk)
	ng2533<=ng23418;

 always  @(posedge pclk)
	ng2616<=ng2609;

 always  @(posedge pclk)
	ng2651<=ng27325;

 always  @(posedge pclk)
	ng2727<=ng23348;

 always  @(posedge pclk)
	ng2784<=ng21043;

 always  @(posedge pclk)
	ng2793<=ng21081;

 always  @(posedge pclk)
	ng2809<=ng25272;

 always  @(posedge pclk)
	ng3043<=ng29453;

 always  @(posedge pclk)
	ng3099<=ng25452;

 always  @(posedge pclk)
	ng3158<=ng17247;

 always  @(posedge pclk)
	ng3179<=ng17383;

 always  @(posedge pclk)
	ng3110<=pg25435;

 always  @(posedge pclk)
	ng164<=ng22125;

 always  @(posedge pclk)
	ng178<=ng25220;

 always  @(posedge pclk)
	ng264<=ng30268;

 always  @(posedge pclk)
	ng74<=ng27594;

 always  @(posedge pclk)
	ng343<=ng27255;

 always  @(posedge pclk)
	ng408<=ng28732;

 always  @(posedge pclk)
	ng448<=ng27759;

 always  @(posedge pclk)
	ng450<=ng11509;

 always  @(posedge pclk)
	ng285<=ng284;

 always  @(posedge pclk)
	ng382<=ng376;

 always  @(posedge pclk)
	ng513<=ng12487;

 always  @(posedge pclk)
	ng572<=ng461;

 always  @(posedge pclk)
	ng455<=ng23385;

 always  @(posedge pclk)
	ng543<=ng13149;

 always  @(posedge pclk)
	ng580<=ng27280;

 always  @(posedge pclk)
	ng584<=ng27327;

 always  @(posedge pclk)
	ng608<=ng28344;

 always  @(posedge pclk)
	ng672<=ng26660;

 always  @(posedge pclk)
	ng705<=ng20893;

 always  @(posedge pclk)
	ng712<=ng20945;

 always  @(posedge pclk)
	ng723<=ng21011;

 always  @(posedge pclk)
	ng738<=ng22218;

 always  @(posedge pclk)
	ng820<=ng22177;

 always  @(posedge pclk)
	ng836<=ng22042;

 always  @(posedge pclk)
	ng844<=ng22127;

 always  @(posedge pclk)
	ng885<=ng30681;

 always  @(posedge pclk)
	ng900<=ng30247;

 always  @(posedge pclk)
	ng912<=ng30642;

 always  @(posedge pclk)
	ng753<=ng28635;

 always  @(posedge pclk)
	ng1078<=ng27313;

 always  @(posedge pclk)
	ng1119<=ng26809;

 always  @(posedge pclk)
	ng1134<=ng27765;

 always  @(posedge pclk)
	ng1010<=ng29173;

 always  @(posedge pclk)
	ng1029<=ng1041;

 always  @(posedge pclk)
	ng1055<=ng1054;

 always  @(posedge pclk)
	ng1210<=ng1209;

 always  @(posedge pclk)
	ng1175<=ng23126;

 always  @(posedge pclk)
	ng1155<=ng24222;

 always  @(posedge pclk)
	ng1234<=ng26534;

 always  @(posedge pclk)
	ng1268<=ng27301;

 always  @(posedge pclk)
	ng1291<=ng28346;

 always  @(posedge pclk)
	ng1216<=ng13427;

 always  @(posedge pclk)
	ng1315<=ng1312;

 always  @(posedge pclk)
	ng1402<=ng21033;

 always  @(posedge pclk)
	ng1416<=ng20975;

 always  @(posedge pclk)
	ng1420<=ng25270;

 always  @(posedge pclk)
	ng1525<=ng22043;

 always  @(posedge pclk)
	ng1540<=ng22131;

 always  @(posedge pclk)
	ng1554<=ng25225;

 always  @(posedge pclk)
	ng1573<=ng30294;

 always  @(posedge pclk)
	ng1444<=ng28147;

 always  @(posedge pclk)
	ng1765<=ng27289;

 always  @(posedge pclk)
	ng1792<=ng28760;

 always  @(posedge pclk)
	ng1819<=ng26816;

 always  @(posedge pclk)
	ng1703<=ng29178;

 always  @(posedge pclk)
	ng1660<=ng1835;

 always  @(posedge pclk)
	ng1903<=ng1893;

 always  @(posedge pclk)
	ng1947<=ng1946;

 always  @(posedge pclk)
	ng1839<=ng23413;

 always  @(posedge pclk)
	ng1908<=ng12482;

 always  @(posedge pclk)
	ng1958<=ng27331;

 always  @(posedge pclk)
	ng1979<=ng24535;

 always  @(posedge pclk)
	ng1874<=ng26573;

 always  @(posedge pclk)
	ng1914<=ng13447;

 always  @(posedge pclk)
	ng2020<=ng20752;

 always  @(posedge pclk)
	ng2080<=ng20915;

 always  @(posedge pclk)
	ng2113<=ng21023;

 always  @(posedge pclk)
	ng2209<=ng22183;

 always  @(posedge pclk)
	ng2239<=ng22173;

 always  @(posedge pclk)
	ng2250<=ng25256;

 always  @(posedge pclk)
	ng2306<=ng30660;

 always  @(posedge pclk)
	ng2285<=ng30304;

 always  @(posedge pclk)
	ng2348<=ng30694;

 always  @(posedge pclk)
	ng2256<=ng13110;

 always  @(posedge pclk)
	ng2444<=ng27292;

 always  @(posedge pclk)
	ng2489<=ng28782;

 always  @(posedge pclk)
	ng2395<=ng30356;

 always  @(posedge pclk)
	ng2529<=ng11592;

 always  @(posedge pclk)
	ng2457<=ng2451;

 always  @(posedge pclk)
	ng2587<=ng12539;

 always  @(posedge pclk)
	ng2646<=ng2536;

 always  @(posedge pclk)
	ng2530<=ng23407;

 always  @(posedge pclk)
	ng2617<=ng13175;

 always  @(posedge pclk)
	ng2654<=ng27337;

 always  @(posedge pclk)
	ng2720<=ng24438;

 always  @(posedge pclk)
	ng2777<=ng20963;

 always  @(posedge pclk)
	ng2795<=ng21074;

 always  @(posedge pclk)
	ng2810<=ng25280;

 always  @(posedge pclk)
	ng3046<=ng29456;

 always  @(posedge pclk)
	ng3100<=ng28420;

 always  @(posedge pclk)
	ng3155<=ng17229;

 always  @(posedge pclk)
	ng3182<=ng17271;

 always  @(posedge pclk)
	ng3120<=pg26104;

 always  @(posedge pclk)
	ng162<=ng22143;

 always  @(posedge pclk)
	ng174<=ng25228;

 always  @(posedge pclk)
	ng222<=ng30635;

 always  @(posedge pclk)
	ng79<=ng27120;

 always  @(posedge pclk)
	ng346<=ng27258;

 always  @(posedge pclk)
	ng391<=ng27293;

 always  @(posedge pclk)
	ng319<=ng30468;

 always  @(posedge pclk)
	ng451<=ng450;

 always  @(posedge pclk)
	ng284<=ng11493;

 always  @(posedge pclk)
	ng383<=ng382;

 always  @(posedge pclk)
	ng510<=ng18726;

 always  @(posedge pclk)
	ng573<=ng572;

 always  @(posedge pclk)
	ng488<=ng23117;

 always  @(posedge pclk)
	ng544<=ng543;

 always  @(posedge pclk)
	ng579<=ng27269;

 always  @(posedge pclk)
	ng587<=ng24491;

 always  @(posedge pclk)
	ng605<=ng28342;

 always  @(posedge pclk)
	ng666<=ng26776;

 always  @(posedge pclk)
	ng701<=ng20901;

 always  @(posedge pclk)
	ng710<=ng20966;

 always  @(posedge pclk)
	ng719<=ng21031;

 always  @(posedge pclk)
	ng739<=ng22231;

 always  @(posedge pclk)
	ng822<=ng22163;

 always  @(posedge pclk)
	ng837<=ng22055;

 always  @(posedge pclk)
	ng846<=ng22105;

 always  @(posedge pclk)
	ng888<=ng30687;

 always  @(posedge pclk)
	ng942<=ng30270;

 always  @(posedge pclk)
	ng915<=ng30647;

 always  @(posedge pclk)
	ng758<=ng28146;

 always  @(posedge pclk)
	ng1095<=ng28738;

 always  @(posedge pclk)
	ng1116<=ng26806;

 always  @(posedge pclk)
	ng999<=ng29609;

 always  @(posedge pclk)
	ng1009<=ng29170;

 always  @(posedge pclk)
	ng1036<=ng1029;

 always  @(posedge pclk)
	ng1054<=ng1048;

 always  @(posedge pclk)
	ng1081<=ng1074;

 always  @(posedge pclk)
	ng1142<=ng23392;

 always  @(posedge pclk)
	ng1152<=ng24212;

 always  @(posedge pclk)
	ng1235<=ng13124;

 always  @(posedge pclk)
	ng1264<=ng27314;

 always  @(posedge pclk)
	ng1215<=ng13426;

 always  @(posedge pclk)
	ng1217<=ng13428;

 always  @(posedge pclk)
	ng1312<=ng1309;

 always  @(posedge pclk)
	ng1406<=ng21017;

 always  @(posedge pclk)
	ng1415<=ng20952;

 always  @(posedge pclk)
	ng1424<=ng22234;

 always  @(posedge pclk)
	ng1524<=ng22035;

 always  @(posedge pclk)
	ng1538<=ng22150;

 always  @(posedge pclk)
	ng1550<=ng25233;

 always  @(posedge pclk)
	ng1555<=ng25234;

 always  @(posedge pclk)
	ng1439<=ng28636;

 always  @(posedge pclk)
	ng1742<=ng27302;

 always  @(posedge pclk)
	ng1795<=ng28771;

 always  @(posedge pclk)
	ng1816<=ng26820;

 always  @(posedge pclk)
	ng1704<=ng29181;

 always  @(posedge pclk)
	ng1835<=ng11565;

 always  @(posedge pclk)
	ng1904<=ng1903;

 always  @(posedge pclk)
	ng1946<=ng1849;

 always  @(posedge pclk)
	ng1842<=ng24182;

 always  @(posedge pclk)
	ng1852<=ng24243;

 always  @(posedge pclk)
	ng1962<=ng27321;

 always  @(posedge pclk)
	ng1976<=ng24525;

 always  @(posedge pclk)
	ng1877<=ng26592;

 always  @(posedge pclk)
	ng1913<=ng13446;

 always  @(posedge pclk)
	ng2013<=ng21972;

 always  @(posedge pclk)
	ng2079<=ng20899;

 always  @(posedge pclk)
	ng2111<=ng21042;

 always  @(posedge pclk)
	ng2205<=ng22192;

 always  @(posedge pclk)
	ng2240<=ng22185;

 always  @(posedge pclk)
	ng2252<=ng25252;

 always  @(posedge pclk)
	ng2309<=ng30666;

 always  @(posedge pclk)
	ng2282<=ng30303;

 always  @(posedge pclk)
	ng2160<=ng25067;

 always  @(posedge pclk)
	ng2120<=ng29582;

 always  @(posedge pclk)
	ng2433<=ng27308;

 always  @(posedge pclk)
	ng2486<=ng28773;

 always  @(posedge pclk)
	ng2397<=ng29182;

 always  @(posedge pclk)
	ng2528<=ng2527;

 always  @(posedge pclk)
	ng2458<=ng2457;

 always  @(posedge pclk)
	ng2584<=ng18820;

 always  @(posedge pclk)
	ng2647<=ng2646;

 always  @(posedge pclk)
	ng2563<=ng21970;

 always  @(posedge pclk)
	ng2618<=ng2617;

 always  @(posedge pclk)
	ng2653<=ng27326;

 always  @(posedge pclk)
	ng2734<=ng25197;

 always  @(posedge pclk)
	ng2776<=ng20940;

 always  @(posedge pclk)
	ng2785<=ng21006;

 always  @(posedge pclk)
	ng2808<=ng25288;

 always  @(posedge pclk)
	ng3045<=ng29455;

 always  @(posedge pclk)
	ng2900<=ng26037;

 always  @(posedge pclk)
	ng3093<=ng17246;

 always  @(posedge pclk)
	ng3104<=ng29939;

 always  @(posedge pclk)
	ng3173<=ng17248;

 always  @(posedge pclk)
	ng3123<=ng28313;

 always  @(posedge pclk)
	ng195<=ng30668;

 always  @(posedge pclk)
	ng255<=ng30262;

 always  @(posedge pclk)
	ng270<=ng30669;

 always  @(posedge pclk)
	ng52<=ng29579;

 always  @(posedge pclk)
	ng388<=ng27278;

 always  @(posedge pclk)
	ng298<=ng26106;

 always  @(posedge pclk)
	ng367<=ng361;

 always  @(posedge pclk)
	ng570<=ng458;

 always  @(posedge pclk)
	ng487<=ng23093;

 always  @(posedge pclk)
	ng529<=ng13410;

 always  @(posedge pclk)
	ng659<=ng20314;

 always  @(posedge pclk)
	ng721<=ng21010;

 always  @(posedge pclk)
	ng737<=ng22242;

 always  @(posedge pclk)
	ng856<=ng25221;

 always  @(posedge pclk)
	ng876<=ng30277;

 always  @(posedge pclk)
	ng1098<=ng28746;

 always  @(posedge pclk)
	ng1125<=ng26810;

 always  @(posedge pclk)
	ng1141<=ng11538;

 always  @(posedge pclk)
	ng976<=ng975;

 always  @(posedge pclk)
	ng1145<=ng23406;

 always  @(posedge pclk)
	ng1214<=ng12467;

 always  @(posedge pclk)
	ng1263<=ng27285;

 always  @(posedge pclk)
	ng1282<=ng24511;

 always  @(posedge pclk)
	ng1183<=ng26569;

 always  @(posedge pclk)
	ng1407<=ng21034;

 always  @(posedge pclk)
	ng1418<=ng20976;

 always  @(posedge pclk)
	ng1511<=ng22178;

 always  @(posedge pclk)
	ng1531<=ng22074;

 always  @(posedge pclk)
	ng1534<=ng22091;

 always  @(posedge pclk)
	ng1545<=ng22152;

 always  @(posedge pclk)
	ng1435<=ng29111;

 always  @(posedge pclk)
	ng1757<=ng27317;

 always  @(posedge pclk)
	ng1809<=ng28772;

 always  @(posedge pclk)
	ng1693<=ng29613;

 always  @(posedge pclk)
	ng1696<=ng30704;

 always  @(posedge pclk)
	ng1783<=ng26675;

 always  @(posedge pclk)
	ng1944<=ng1836;

 always  @(posedge pclk)
	ng1870<=ng1948;

 always  @(posedge pclk)
	ng1865<=ng23030;

 always  @(posedge pclk)
	ng1929<=ng13135;

 always  @(posedge pclk)
	ng1939<=ng1938;

 always  @(posedge pclk)
	ng1966<=ng27341;

 always  @(posedge pclk)
	ng1886<=ng1880;

 always  @(posedge pclk)
	ng1917<=ng13449;

 always  @(posedge pclk)
	ng2089<=ng20978;

 always  @(posedge pclk)
	ng2100<=ng21041;

 always  @(posedge pclk)
	ng2108<=ng21022;

 always  @(posedge pclk)
	ng2207<=ng22182;

 always  @(posedge pclk)
	ng2238<=ng22194;

 always  @(posedge pclk)
	ng2255<=ng25257;

 always  @(posedge pclk)
	ng2315<=ng30667;

 always  @(posedge pclk)
	ng2294<=ng30260;

 always  @(posedge pclk)
	ng2339<=ng30297;

 always  @(posedge pclk)
	ng2142<=ng27621;

 always  @(posedge pclk)
	ng2418<=ng27291;

 always  @(posedge pclk)
	ng2483<=ng28763;

 always  @(posedge pclk)
	ng2398<=ng29185;

 always  @(posedge pclk)
	ng2355<=ng11572;

 always  @(posedge pclk)
	ng2366<=ng2365;

 always  @(posedge pclk)
	ng2439<=ng2432;

 always  @(posedge pclk)
	ng2644<=ng2533;

 always  @(posedge pclk)
	ng2562<=ng23133;

 always  @(posedge pclk)
	ng2670<=ng24538;

 always  @(posedge pclk)
	ng2571<=ng26616;

 always  @(posedge pclk)
	ng2610<=ng13464;

 always  @(posedge pclk)
	ng2812<=ng22269;

 always  @(posedge pclk)
	ng3048<=ng29458;

 always  @(posedge pclk)
	ng3094<=ng17226;

 always  @(posedge pclk)
	ng3103<=ng29936;

 always  @(posedge pclk)
	ng3176<=ng17303;

 always  @(posedge pclk)
	ng3124<=pg25442;

 always  @(posedge pclk)
	ng198<=ng30674;

 always  @(posedge pclk)
	ng252<=ng30257;

 always  @(posedge pclk)
	ng213<=ng30245;

 always  @(posedge pclk)
	ng354<=ng27253;

 always  @(posedge pclk)
	ng398<=ng27267;

 always  @(posedge pclk)
	ng342<=ng354;

 always  @(posedge pclk)
	ng366<=ng365;

 always  @(posedge pclk)
	ng571<=ng570;

 always  @(posedge pclk)
	ng486<=ng23067;

 always  @(posedge pclk)
	ng530<=ng13411;

 always  @(posedge pclk)
	ng630<=ng16654;

 always  @(posedge pclk)
	ng711<=ng20923;

 always  @(posedge pclk)
	ng830<=ng22029;

 always  @(posedge pclk)
	ng860<=ng25215;

 always  @(posedge pclk)
	ng873<=ng30269;

 always  @(posedge pclk)
	ng1101<=ng28758;

 always  @(posedge pclk)
	ng1122<=ng26813;

 always  @(posedge pclk)
	ng966<=ng1141;

 always  @(posedge pclk)
	ng975<=ng11522;

 always  @(posedge pclk)
	ng1148<=ng24179;

 always  @(posedge pclk)
	ng1158<=ng24235;

 always  @(posedge pclk)
	ng1270<=ng27339;

 always  @(posedge pclk)
	ng1285<=ng24522;

 always  @(posedge pclk)
	ng1180<=ng26557;

 always  @(posedge pclk)
	ng1405<=ng21052;

 always  @(posedge pclk)
	ng1414<=ng20996;

 always  @(posedge pclk)
	ng1515<=ng22167;

 always  @(posedge pclk)
	ng1530<=ng22059;

 always  @(posedge pclk)
	ng1532<=ng22112;

 always  @(posedge pclk)
	ng1541<=ng22168;

 always  @(posedge pclk)
	ng1430<=ng29355;

 always  @(posedge pclk)
	ng1754<=ng27303;

 always  @(posedge pclk)
	ng1807<=ng28778;

 always  @(posedge pclk)
	ng1828<=ng27768;

 always  @(posedge pclk)
	ng1697<=ng30706;

 always  @(posedge pclk)
	ng1785<=ng26670;

 always  @(posedge pclk)
	ng1949<=ng1944;

 always  @(posedge pclk)
	ng1948<=ng1852;

 always  @(posedge pclk)
	ng1845<=ng23058;

 always  @(posedge pclk)
	ng1928<=ng29113;

 always  @(posedge pclk)
	ng1956<=ng27290;

 always  @(posedge pclk)
	ng1965<=ng27333;

 always  @(posedge pclk)
	ng1887<=ng22651;

 always  @(posedge pclk)
	ng1916<=ng13448;

 always  @(posedge pclk)
	ng2087<=ng20999;

 always  @(posedge pclk)
	ng2096<=ng21054;

 always  @(posedge pclk)
	ng2112<=ng21003;

 always  @(posedge pclk)
	ng2206<=ng22170;

 always  @(posedge pclk)
	ng2245<=ng25227;

 always  @(posedge pclk)
	ng2254<=ng25253;

 always  @(posedge pclk)
	ng2318<=ng30673;

 always  @(posedge pclk)
	ng2291<=ng30256;

 always  @(posedge pclk)
	ng2297<=ng30652;

 always  @(posedge pclk)
	ng2147<=ng27131;

 always  @(posedge pclk)
	ng2421<=ng27307;

 always  @(posedge pclk)
	ng2466<=ng27342;

 always  @(posedge pclk)
	ng2396<=ng29187;

 always  @(posedge pclk)
	ng2354<=ng2529;

 always  @(posedge pclk)
	ng2374<=ng19048;

 always  @(posedge pclk)
	ng2432<=ng2444;

 always  @(posedge pclk)
	ng2645<=ng2644;

 always  @(posedge pclk)
	ng2561<=ng23114;

 always  @(posedge pclk)
	ng2652<=ng27343;

 always  @(posedge pclk)
	ng2580<=ng2574;

 always  @(posedge pclk)
	ng2608<=ng13463;

 always  @(posedge pclk)
	ng2813<=ng22284;

 always  @(posedge pclk)
	ng3047<=ng29457;

 always  @(posedge pclk)
	ng3095<=ng17235;

 always  @(posedge pclk)
	ng3106<=ng30796;

 always  @(posedge pclk)
	ng3167<=ng17270;

 always  @(posedge pclk)
	ng3125<=ng28696;

 always  @(posedge pclk)
	ng216<=ng30246;

 always  @(posedge pclk)
	ng92<=ng25027;

 always  @(posedge pclk)
	ng376<=ng27277;

 always  @(posedge pclk)
	ng349<=ng342;

 always  @(posedge pclk)
	ng372<=ng384;

 always  @(posedge pclk)
	ng324<=ng397;

 always  @(posedge pclk)
	ng531<=ng13412;

 always  @(posedge pclk)
	ng633<=ng23136;

 always  @(posedge pclk)
	ng698<=ng20891;

 always  @(posedge pclk)
	ng840<=ng22067;

 always  @(posedge pclk)
	ng861<=ng25222;

 always  @(posedge pclk)
	ng918<=ng30643;

 always  @(posedge pclk)
	ng1002<=ng30701;

 always  @(posedge pclk)
	ng1089<=ng26669;

 always  @(posedge pclk)
	ng967<=ng11518;

 always  @(posedge pclk)
	ng978<=ng977;

 always  @(posedge pclk)
	ng1164<=ng24181;

 always  @(posedge pclk)
	ng1245<=ng1244;

 always  @(posedge pclk)
	ng1272<=ng27329;

 always  @(posedge pclk)
	ng1288<=ng24532;

 always  @(posedge pclk)
	ng1193<=ng22615;

 always  @(posedge pclk)
	ng1409<=ng21035;

 always  @(posedge pclk)
	ng1417<=ng21018;

 always  @(posedge pclk)
	ng1512<=ng22149;

 always  @(posedge pclk)
	ng1526<=ng22073;

 always  @(posedge pclk)
	ng1536<=ng22092;

 always  @(posedge pclk)
	ng1544<=ng22180;

 always  @(posedge pclk)
	ng1426<=ng29581;

 always  @(posedge pclk)
	ng1769<=ng27318;

 always  @(posedge pclk)
	ng1804<=ng29218;

 always  @(posedge pclk)
	ng1830<=ng27766;

 always  @(posedge pclk)
	ng1698<=ng30708;

 always  @(posedge pclk)
	ng1832<=ng1831;

 always  @(posedge pclk)
	ng1950<=ng1839;

 always  @(posedge pclk)
	ng1868<=ng23124;

 always  @(posedge pclk)
	ng1860<=ng24231;

 always  @(posedge pclk)
	ng1924<=ng1923;

 always  @(posedge pclk)
	ng1957<=ng27305;

 always  @(posedge pclk)
	ng1967<=ng24513;

 always  @(posedge pclk)
	ng2040<=ng25194;

 always  @(posedge pclk)
	ng2081<=ng20953;

 always  @(posedge pclk)
	ng2091<=ng20979;

 always  @(posedge pclk)
	ng2099<=ng21071;

 always  @(posedge pclk)
	ng2109<=ng20980;

 always  @(posedge pclk)
	ng2117<=ng22280;

 always  @(posedge pclk)
	ng2246<=ng25236;

 always  @(posedge pclk)
	ng2261<=ng30289;

 always  @(posedge pclk)
	ng2273<=ng30693;

 always  @(posedge pclk)
	ng2288<=ng30253;

 always  @(posedge pclk)
	ng2300<=ng30659;

 always  @(posedge pclk)
	ng2133<=ng28637;

 always  @(posedge pclk)
	ng2463<=ng27335;

 always  @(posedge pclk)
	ng2478<=ng26672;

 always  @(posedge pclk)
	ng2357<=ng11573;

 always  @(posedge pclk)
	ng2364<=ng2363;

 always  @(posedge pclk)
	ng2428<=ng2427;

 always  @(posedge pclk)
	ng2447<=ng2459;

 always  @(posedge pclk)
	ng2399<=ng2472;

 always  @(posedge pclk)
	ng2656<=ng27338;

 always  @(posedge pclk)
	ng2676<=ng24557;

 always  @(posedge pclk)
	ng2607<=ng13462;

 always  @(posedge pclk)
	ng2811<=ng22299;

 always  @(posedge pclk)
	ng3096<=ng17269;

 always  @(posedge pclk)
	ng3105<=ng29941;

 always  @(posedge pclk)
	ng3170<=ng17340;

 always  @(posedge pclk)
	ng3126<=pg25420;

 always  @(posedge pclk)
	ng219<=ng30248;

 always  @(posedge pclk)
	ng273<=ng30675;

 always  @(posedge pclk)
	ng56<=ng29353;

 always  @(posedge pclk)
	ng368<=ng367;

 always  @(posedge pclk)
	ng379<=ng372;

 always  @(posedge pclk)
	ng397<=ng391;

 always  @(posedge pclk)
	ng532<=ng13413;

 always  @(posedge pclk)
	ng640<=ng20682;

 always  @(posedge pclk)
	ng653<=ng23324;

 always  @(posedge pclk)
	ng847<=ng22147;

 always  @(posedge pclk)
	ng859<=ng25230;

 always  @(posedge pclk)
	ng879<=ng30285;

 always  @(posedge pclk)
	ng1003<=ng30703;

 always  @(posedge pclk)
	ng1091<=ng26665;

 always  @(posedge pclk)
	ng968<=ng967;

 always  @(posedge pclk)
	ng977<=ng2873;

 always  @(posedge pclk)
	ng1221<=ng1214;

 always  @(posedge pclk)
	ng1262<=ng27273;

 always  @(posedge pclk)
	ng1271<=ng27316;

 always  @(posedge pclk)
	ng1300<=ng28351;

 always  @(posedge pclk)
	ng1192<=ng1186;

 always  @(posedge pclk)
	ng1410<=ng21053;

 always  @(posedge pclk)
	ng1419<=ng20997;

 always  @(posedge pclk)
	ng1513<=ng22166;

 always  @(posedge pclk)
	ng1528<=ng22058;

 always  @(posedge pclk)
	ng1537<=ng22113;

 always  @(posedge pclk)
	ng1546<=ng22169;

 always  @(posedge pclk)
	ng1735<=ng27264;

 always  @(posedge pclk)
	ng1779<=ng27304;

 always  @(posedge pclk)
	ng1808<=ng28761;

 always  @(posedge pclk)
	ng1829<=ng27764;

 always  @(posedge pclk)
	ng1699<=ng30487;

 always  @(posedge pclk)
	ng1831<=ng11563;

 always  @(posedge pclk)
	ng1951<=ng1950;

 always  @(posedge pclk)
	ng1867<=ng23097;

 always  @(posedge pclk)
	ng1861<=ng23123;

 always  @(posedge pclk)
	ng1923<=ng13164;

 always  @(posedge pclk)
	ng1955<=ng27319;

 always  @(posedge pclk)
	ng1964<=ng27346;

 always  @(posedge pclk)
	ng2052<=ng26671;

 always  @(posedge pclk)
	ng2083<=ng20935;

 always  @(posedge pclk)
	ng2092<=ng21000;

 always  @(posedge pclk)
	ng2101<=ng21055;

 always  @(posedge pclk)
	ng2110<=ng21002;

 always  @(posedge pclk)
	ng2119<=ng22267;

 always  @(posedge pclk)
	ng2244<=ng25245;

 always  @(posedge pclk)
	ng2253<=ng25259;

 always  @(posedge pclk)
	ng2276<=ng30695;

 always  @(posedge pclk)
	ng2330<=ng30290;

 always  @(posedge pclk)
	ng2303<=ng30665;

 always  @(posedge pclk)
	ng2138<=ng28148;

 always  @(posedge pclk)
	ng2429<=ng27276;

 always  @(posedge pclk)
	ng2473<=ng27324;

 always  @(posedge pclk)
	ng2479<=ng26676;

 always  @(posedge pclk)
	ng2356<=ng2355;

 always  @(posedge pclk)
	ng2365<=ng2878;

 always  @(posedge pclk)
	ng2427<=ng2421;

 always  @(posedge pclk)
	ng2454<=ng2447;

 always  @(posedge pclk)
	ng2472<=ng2466;

 always  @(posedge pclk)
	ng2657<=ng27344;

 always  @(posedge pclk)
	ng2673<=ng24548;

 always  @(posedge pclk)
	ng2568<=ng26596;

 always  @(posedge pclk)
	ng3049<=ng29459;

 always  @(posedge pclk)
	ng2888<=ng22026;

 always  @(posedge pclk)
	ng130<=ng22100;

 always  @(posedge pclk)
	ng144<=ng22037;

 always  @(posedge pclk)
	ng158<=ng22080;

 always  @(posedge pclk)
	ng172<=ng25207;

 always  @(posedge pclk)
	ng192<=ng30275;

 always  @(posedge pclk)
	ng207<=ng30284;

 always  @(posedge pclk)
	ng449<=ng27760;

 always  @(posedge pclk)
	ng322<=ng29167;

 always  @(posedge pclk)
	ng279<=ng454;

 always  @(posedge pclk)
	ng290<=ng2857;

 always  @(posedge pclk)
	ng357<=ng369;

 always  @(posedge pclk)
	ng578<=ng27294;

 always  @(posedge pclk)
	ng599<=ng24508;

 always  @(posedge pclk)
	ng506<=ng499;

 always  @(posedge pclk)
	ng537<=ng13417;

 always  @(posedge pclk)
	ng700<=ng20879;

 always  @(posedge pclk)
	ng838<=ng22087;

 always  @(posedge pclk)
	ng852<=ng22148;

 always  @(posedge pclk)
	ng866<=ng25232;

 always  @(posedge pclk)
	ng894<=ng30293;

 always  @(posedge pclk)
	ng909<=ng30638;

 always  @(posedge pclk)
	ng1137<=ng11536;

 always  @(posedge pclk)
	ng972<=ng971;

 always  @(posedge pclk)
	ng1044<=ng1056;

 always  @(posedge pclk)
	ng1070<=ng1069;

 always  @(posedge pclk)
	ng1209<=ng1199;

 always  @(posedge pclk)
	ng1294<=ng28350;

 always  @(posedge pclk)
	ng1223<=ng13433;

 always  @(posedge pclk)
	ng1332<=ng24430;

 always  @(posedge pclk)
	ng1389<=ng20911;

 always  @(posedge pclk)
	ng1400<=ng20974;

 always  @(posedge pclk)
	ng1560<=ng25244;

 always  @(posedge pclk)
	ng1582<=ng30692;

 always  @(posedge pclk)
	ng1597<=ng30252;

 always  @(posedge pclk)
	ng1466<=ng25056;

 always  @(posedge pclk)
	ng1666<=ng1665;

 always  @(posedge pclk)
	ng1730<=ng1723;

 always  @(posedge pclk)
	ng1753<=ng1765;

 always  @(posedge pclk)
	ng1705<=ng1778;

 always  @(posedge pclk)
	ng2217<=ng22076;

 always  @(posedge pclk)
	ng2231<=ng22139;

 always  @(posedge pclk)
	ng2248<=ng25237;

 always  @(posedge pclk)
	ng2503<=ng28783;

 always  @(posedge pclk)
	ng2387<=ng29618;

 always  @(posedge pclk)
	ng2477<=ng26025;

 always  @(posedge pclk)
	ng2359<=ng11574;

 always  @(posedge pclk)
	ng2417<=ng2429;

 always  @(posedge pclk)
	ng2443<=ng2442;

 always  @(posedge pclk)
	ng2655<=ng27347;

 always  @(posedge pclk)
	ng2691<=ng28368;

 always  @(posedge pclk)
	ng2599<=pg16437;

 always  @(posedge pclk)
	ng2704<=ng16718;

 always  @(posedge pclk)
	ng2766<=ng28328;

 always  @(posedge pclk)
	ng2783<=ng21005;

 always  @(posedge pclk)
	ng2794<=ng21062;

 always  @(posedge pclk)
	ng3050<=ng29460;

 always  @(posedge pclk)
	ng3062<=ng30908;

 always  @(posedge pclk)
	ng3073<=ng30982;

 always  @(posedge pclk)
	ng3013<=ng25191;

 always  @(posedge pclk)
	pg8274<=ng16844;

 always  @(posedge pclk)
	pg8265<=ng16854;

 always  @(posedge pclk)
	ng2896<=ng23358;

 always  @(posedge pclk)
	ng131<=ng22122;

 always  @(posedge pclk)
	ng146<=ng22031;

 always  @(posedge pclk)
	ng156<=ng22101;

 always  @(posedge pclk)
	ng168<=ng25211;

 always  @(posedge pclk)
	ng231<=ng30637;

 always  @(posedge pclk)
	ng204<=ng30276;

 always  @(posedge pclk)
	ng427<=ng28736;

 always  @(posedge pclk)
	ng323<=ng29169;

 always  @(posedge pclk)
	ng454<=ng11511;

 always  @(posedge pclk)
	ng291<=ng290;

 always  @(posedge pclk)
	ng353<=ng352;

 always  @(posedge pclk)
	ng582<=ng27281;

 always  @(posedge pclk)
	ng596<=ng24499;

 always  @(posedge pclk)
	ng507<=ng22578;

 always  @(posedge pclk)
	ng536<=ng13416;

 always  @(posedge pclk)
	ng707<=ng20944;

 always  @(posedge pclk)
	ng831<=ng22033;

 always  @(posedge pclk)
	ng850<=ng22164;

 always  @(posedge pclk)
	ng862<=ng25240;

 always  @(posedge pclk)
	ng897<=ng30298;

 always  @(posedge pclk)
	ng951<=ng30278;

 always  @(posedge pclk)
	ng1138<=ng1137;

 always  @(posedge pclk)
	ng971<=ng11520;

 always  @(posedge pclk)
	ng1051<=ng1044;

 always  @(posedge pclk)
	ng1069<=ng1063;

 always  @(posedge pclk)
	ng1252<=ng1155;

 always  @(posedge pclk)
	ng1273<=ng24501;

 always  @(posedge pclk)
	ng1224<=ng24072;

 always  @(posedge pclk)
	ng1339<=ng23329;

 always  @(posedge pclk)
	ng1387<=ng20925;

 always  @(posedge pclk)
	ng1396<=ng20993;

 always  @(posedge pclk)
	ng1561<=ng25250;

 always  @(posedge pclk)
	ng1579<=ng30688;

 always  @(posedge pclk)
	ng1600<=ng30255;

 always  @(posedge pclk)
	ng1654<=ng30689;

 always  @(posedge pclk)
	ng1667<=ng11548;

 always  @(posedge pclk)
	ng1723<=ng1735;

 always  @(posedge pclk)
	ng1760<=ng1753;

 always  @(posedge pclk)
	ng1778<=ng1772;

 always  @(posedge pclk)
	ng2221<=ng22061;

 always  @(posedge pclk)
	ng2230<=ng22117;

 always  @(posedge pclk)
	ng2264<=ng30296;

 always  @(posedge pclk)
	ng2501<=ng28788;

 always  @(posedge pclk)
	ng2522<=ng27771;

 always  @(posedge pclk)
	ng2525<=ng11590;

 always  @(posedge pclk)
	ng2358<=ng2357;

 always  @(posedge pclk)
	ng2424<=ng2417;

 always  @(posedge pclk)
	ng2442<=ng2436;

 always  @(posedge pclk)
	ng2659<=ng27345;

 always  @(posedge pclk)
	ng2688<=ng28364;

 always  @(posedge pclk)
	ng2603<=ng13458;

 always  @(posedge pclk)
	ng2615<=ng13466;

 always  @(posedge pclk)
	ng2773<=ng20918;

 always  @(posedge pclk)
	ng2782<=ng20983;

 always  @(posedge pclk)
	ng2804<=ng21028;

 always  @(posedge pclk)
	ng3051<=ng29655;

 always  @(posedge pclk)
	ng3061<=ng30119;

 always  @(posedge pclk)
	ng3074<=ng30983;

 always  @(posedge pclk)
	ng3002<=ng24445;

 always  @(posedge pclk)
	pg8273<=ng16853;

 always  @(posedge pclk)
	pg8266<=ng16845;

 always  @(posedge pclk)
	ng2892<=ng24473;

 always  @(posedge pclk)
	ng129<=ng22141;

 always  @(posedge pclk)
	ng149<=ng22038;

 always  @(posedge pclk)
	ng153<=ng22079;

 always  @(posedge pclk)
	ng170<=ng25206;

 always  @(posedge pclk)
	ng234<=ng30640;

 always  @(posedge pclk)
	ng249<=ng30254;

 always  @(posedge pclk)
	ng428<=ng28745;

 always  @(posedge pclk)
	ng312<=ng29606;

 always  @(posedge pclk)
	ng453<=ng452;

 always  @(posedge pclk)
	ng299<=ng19012;

 always  @(posedge pclk)
	ng365<=ng358;

 always  @(posedge pclk)
	ng484<=ng23000;

 always  @(posedge pclk)
	ng549<=ng13111;

 always  @(posedge pclk)
	pg16297<=ng21435;

 always  @(posedge pclk)
	ng541<=ng13418;

 always  @(posedge pclk)
	ng720<=ng20991;

 always  @(posedge pclk)
	ng826<=ng2950;

 always  @(posedge pclk)
	ng857<=ng25209;

 always  @(posedge pclk)
	ng865<=ng25248;

 always  @(posedge pclk)
	ng767<=ng27123;

 always  @(posedge pclk)
	ng1045<=ng27271;

 always  @(posedge pclk)
	ng1139<=ng11537;

 always  @(posedge pclk)
	ng974<=ng973;

 always  @(posedge pclk)
	ng1052<=ng1045;

 always  @(posedge pclk)
	ng1196<=ng18763;

 always  @(posedge pclk)
	ng1251<=ng1260;

 always  @(posedge pclk)
	ng1276<=ng24510;

 always  @(posedge pclk)
	ng1177<=ng26547;

 always  @(posedge pclk)
	ng1227<=ng13434;

 always  @(posedge pclk)
	ng1358<=ng26666;

 always  @(posedge pclk)
	ng1384<=ng20910;

 always  @(posedge pclk)
	ng1398<=ng20973;

 always  @(posedge pclk)
	ng1529<=ng22090;

 always  @(posedge pclk)
	ng1543<=ng22151;

 always  @(posedge pclk)
	ng1559<=ng25255;

 always  @(posedge pclk)
	ng1624<=ng30664;

 always  @(posedge pclk)
	ng1636<=ng30280;

 always  @(posedge pclk)
	ng1651<=ng30684;

 always  @(posedge pclk)
	ng1784<=ng26667;

 always  @(posedge pclk)
	ng1668<=ng1667;

 always  @(posedge pclk)
	ng1732<=ng1731;

 always  @(posedge pclk)
	ng1748<=ng1742;

 always  @(posedge pclk)
	ng1777<=ng1776;

 always  @(posedge pclk)
	ng2222<=ng22077;

 always  @(posedge pclk)
	ng2233<=ng22140;

 always  @(posedge pclk)
	ng2321<=ng30679;

 always  @(posedge pclk)
	ng2504<=ng26817;

 always  @(posedge pclk)
	ng2389<=ng29623;

 always  @(posedge pclk)
	ng2526<=ng2525;

 always  @(posedge pclk)
	ng2361<=ng11575;

 always  @(posedge pclk)
	ng2380<=ng30055;

 always  @(posedge pclk)
	ng2441<=ng2440;

 always  @(posedge pclk)
	ng2559<=ng23047;

 always  @(posedge pclk)
	ng2623<=ng13143;

 always  @(posedge pclk)
	ng2660<=ng27348;

 always  @(posedge pclk)
	ng2679<=ng28358;

 always  @(posedge pclk)
	ng2581<=ng22687;

 always  @(posedge pclk)
	ng2612<=ng24092;

 always  @(posedge pclk)
	ng2774<=ng20939;

 always  @(posedge pclk)
	ng2792<=ng21061;

 always  @(posedge pclk)
	ng2803<=ng21007;

 always  @(posedge pclk)
	ng3052<=ng29972;

 always  @(posedge pclk)
	ng3064<=ng30910;

 always  @(posedge pclk)
	ng3071<=ng30980;

 always  @(posedge pclk)
	ng3006<=ng23330;

 always  @(posedge pclk)
	pg8272<=ng16860;

 always  @(posedge pclk)
	pg8262<=ng16880;

 always  @(posedge pclk)
	pg8258<=ng18542;

 always  @(posedge pclk)
	ng2903<=ng25201;

 always  @(posedge pclk)
	ng133<=ng22123;

 always  @(posedge pclk)
	ng148<=ng22032;

 always  @(posedge pclk)
	ng157<=ng22065;

 always  @(posedge pclk)
	ng169<=ng25204;

 always  @(posedge pclk)
	ng237<=ng30645;

 always  @(posedge pclk)
	ng210<=ng30292;

 always  @(posedge pclk)
	ng426<=ng28754;

 always  @(posedge pclk)
	ng447<=ng27762;

 always  @(posedge pclk)
	ng320<=ng30482;

 always  @(posedge pclk)
	ng305<=ng21346;

 always  @(posedge pclk)
	ng364<=ng357;

 always  @(posedge pclk)
	ng464<=ng23022;

 always  @(posedge pclk)
	ng548<=ng21851;

 always  @(posedge pclk)
	ng525<=pg16297;

 always  @(posedge pclk)
	ng538<=ng24059;

 always  @(posedge pclk)
	ng730<=ng20947;

 always  @(posedge pclk)
	ng728<=ng20969;

 always  @(posedge pclk)
	ng858<=ng25214;

 always  @(posedge pclk)
	ng867<=ng25241;

 always  @(posedge pclk)
	ng762<=ng27603;

 always  @(posedge pclk)
	ng1056<=ng27263;

 always  @(posedge pclk)
	ng1140<=ng1139;

 always  @(posedge pclk)
	ng973<=ng11521;

 always  @(posedge pclk)
	ng1074<=ng1085;

 always  @(posedge pclk)
	ng1199<=ng12507;

 always  @(posedge pclk)
	ng1260<=ng1152;

 always  @(posedge pclk)
	ng1279<=ng24521;

 always  @(posedge pclk)
	ng1297<=ng28354;

 always  @(posedge pclk)
	ng1309<=ng3080;

 always  @(posedge pclk)
	ng1346<=ng25189;

 always  @(posedge pclk)
	ng1388<=ng20897;

 always  @(posedge pclk)
	ng1397<=ng20951;

 always  @(posedge pclk)
	ng1533<=ng22075;

 always  @(posedge pclk)
	ng1542<=ng22132;

 always  @(posedge pclk)
	ng1567<=ng30279;

 always  @(posedge pclk)
	ng1621<=ng30658;

 always  @(posedge pclk)
	ng1594<=ng30250;

 always  @(posedge pclk)
	ng1648<=ng30678;

 always  @(posedge pclk)
	ng1695<=ng29620;

 always  @(posedge pclk)
	ng1669<=ng11549;

 always  @(posedge pclk)
	ng1731<=ng1724;

 always  @(posedge pclk)
	ng1749<=ng1748;

 always  @(posedge pclk)
	ng1776<=ng1769;

 always  @(posedge pclk)
	ng2220<=ng22097;

 always  @(posedge pclk)
	ng2229<=ng22153;

 always  @(posedge pclk)
	ng2333<=ng30283;

 always  @(posedge pclk)
	ng2507<=ng26822;

 always  @(posedge pclk)
	ng2388<=ng29621;

 always  @(posedge pclk)
	ng2527<=ng11591;

 always  @(posedge pclk)
	ng2360<=ng2359;

 always  @(posedge pclk)
	ng2373<=ng26144;

 always  @(posedge pclk)
	ng2440<=ng2433;

 always  @(posedge pclk)
	ng2539<=ng23076;

 always  @(posedge pclk)
	ng2622<=ng30072;

 always  @(posedge pclk)
	ng2658<=ng27354;

 always  @(posedge pclk)
	ng2694<=ng28371;

 always  @(posedge pclk)
	pg16437<=ng30061;

 always  @(posedge pclk)
	ng2611<=ng13465;

 always  @(posedge pclk)
	ng2781<=ng21025;

 always  @(posedge pclk)
	ng2790<=ng21073;

 always  @(posedge pclk)
	ng2799<=ng20965;

 always  @(posedge pclk)
	ng3053<=ng29973;

 always  @(posedge pclk)
	ng3063<=ng30909;

 always  @(posedge pclk)
	ng3072<=ng30981;

 always  @(posedge pclk)
	ng2998<=ng26048;

 always  @(posedge pclk)
	pg8268<=ng16803;

 always  @(posedge pclk)
	pg8264<=ng16861;

 always  @(posedge pclk)
	ng2817<=ng16802;

 always  @(posedge pclk)
	ng3101<=ng28421;

 always  @(posedge pclk)
	ng3164<=ng17236;

 always  @(posedge pclk)
	ng134<=ng22142;

 always  @(posedge pclk)
	ng151<=ng22039;

 always  @(posedge pclk)
	ng159<=ng22124;

 always  @(posedge pclk)
	ng176<=ng25219;

 always  @(posedge pclk)
	ng179<=ng25229;

 always  @(posedge pclk)
	ng240<=ng30641;

 always  @(posedge pclk)
	ng225<=ng30636;

 always  @(posedge pclk)
	ng65<=ng28634;

 always  @(posedge pclk)
	ng373<=ng27266;

 always  @(posedge pclk)
	ng429<=ng26803;

 always  @(posedge pclk)
	ng314<=ng29611;

 always  @(posedge pclk)
	ng404<=ng26659;

 always  @(posedge pclk)
	ng283<=ng282;

 always  @(posedge pclk)
	ng350<=ng343;

 always  @(posedge pclk)
	ng387<=ng398;

 always  @(posedge pclk)
	ng524<=ng523;

 always  @(posedge pclk)
	ng568<=ng471;

 always  @(posedge pclk)
	ng480<=ng23092;

 always  @(posedge pclk)
	ng465<=ng24206;

 always  @(posedge pclk)
	ng558<=ng13160;

 always  @(posedge pclk)
	ng585<=ng27296;

 always  @(posedge pclk)
	ng620<=ng28353;

 always  @(posedge pclk)
	ng679<=ng27672;

 always  @(posedge pclk)
	ng704<=ng20921;

 always  @(posedge pclk)
	ng718<=ng20990;

 always  @(posedge pclk)
	ng729<=ng20924;

 always  @(posedge pclk)
	ng732<=ng20948;

 always  @(posedge pclk)
	ng853<=ng823;

 always  @(posedge pclk)
	ng834<=ng22041;

 always  @(posedge pclk)
	ng845<=ng22089;

 always  @(posedge pclk)
	ng927<=ng30649;

 always  @(posedge pclk)
	ng906<=ng30251;

 always  @(posedge pclk)
	ng776<=ng25935;

 always  @(posedge pclk)
	ng1033<=ng27270;

 always  @(posedge pclk)
	ng1048<=ng27282;

 always  @(posedge pclk)
	ng1107<=ng29204;

 always  @(posedge pclk)
	ng1135<=ng27761;

 always  @(posedge pclk)
	ng1007<=ng30500;

 always  @(posedge pclk)
	ng1037<=ng1030;

 always  @(posedge pclk)
	ng1066<=ng1059;

 always  @(posedge pclk)
	ng1240<=ng21843;

 always  @(posedge pclk)
	ng1259<=ng1258;

 always  @(posedge pclk)
	ng1165<=ng24213;

 always  @(posedge pclk)
	ng1229<=ng13155;

 always  @(posedge pclk)
	ng1266<=ng27300;

 always  @(posedge pclk)
	ng1218<=ng13429;

 always  @(posedge pclk)
	ng1345<=ng20333;

 always  @(posedge pclk)
	ng1385<=ng20882;

 always  @(posedge pclk)
	ng1393<=ng20972;

 always  @(posedge pclk)
	ng1421<=ng25263;

 always  @(posedge pclk)
	ng1514<=ng22191;

 always  @(posedge pclk)
	ng1553<=ng25242;

 always  @(posedge pclk)
	ng1615<=ng30657;

 always  @(posedge pclk)
	ng1630<=ng30266;

 always  @(posedge pclk)
	ng1609<=ng30656;

 always  @(posedge pclk)
	ng1813<=ng26815;

 always  @(posedge pclk)
	ng1662<=ng1661;

 always  @(posedge pclk)
	ng1680<=ng19036;

 always  @(posedge pclk)
	ng1746<=ng1739;

 always  @(posedge pclk)
	ng1775<=ng1768;

 always  @(posedge pclk)
	ng2224<=ng22078;

 always  @(posedge pclk)
	ng2232<=ng22171;

 always  @(posedge pclk)
	ng2156<=ng25940;

 always  @(posedge pclk)
	ng2510<=ng26825;

 always  @(posedge pclk)
	ng2391<=ng30709;

 always  @(posedge pclk)
	ng2462<=ng2473;

 always  @(posedge pclk)
	ng2598<=ng2597;

 always  @(posedge pclk)
	ng2642<=ng2546;

 always  @(posedge pclk)
	ng2555<=ng23132;

 always  @(posedge pclk)
	ng2540<=ng24225;

 always  @(posedge pclk)
	ng2632<=ng13194;

 always  @(posedge pclk)
	ng2661<=ng24527;

 always  @(posedge pclk)
	ng2685<=ng28367;

 always  @(posedge pclk)
	ng2606<=ng13461;

 always  @(posedge pclk)
	ng2746<=ng26677;

 always  @(posedge pclk)
	ng2779<=ng20964;

 always  @(posedge pclk)
	ng2787<=ng21060;

 always  @(posedge pclk)
	ng2801<=ng20941;

 always  @(posedge pclk)
	ng3054<=ng20877;

 always  @(posedge pclk)
	ng3055<=ng29974;

 always  @(posedge pclk)
	ng3066<=ng30912;

 always  @(posedge pclk)
	ng3077<=ng30986;

 always  @(posedge pclk)
	ng3028<=ng23359;

 always  @(posedge pclk)
	pg5388<=pg3234;

 always  @(posedge pclk)
	ng3083<=ng16866;

 always  @(posedge pclk)
	ng2990<=ng18907;

 always  @(posedge pclk)
	ng2933<=ng16823;

 always  @(posedge pclk)
	ng3102<=ng28425;

 always  @(posedge pclk)
	ng3161<=ng17302;

 always  @(posedge pclk)
	ng132<=ng22161;

 always  @(posedge pclk)
	ng147<=ng22047;

 always  @(posedge pclk)
	ng163<=ng22103;

 always  @(posedge pclk)
	ng175<=ng25213;

 always  @(posedge pclk)
	ng177<=ng25239;

 always  @(posedge pclk)
	ng201<=ng30680;

 always  @(posedge pclk)
	ng228<=ng30639;

 always  @(posedge pclk)
	ng70<=ng28145;

 always  @(posedge pclk)
	ng423<=ng29201;

 always  @(posedge pclk)
	ng432<=ng26804;

 always  @(posedge pclk)
	ng313<=ng29608;

 always  @(posedge pclk)
	ng402<=ng26664;

 always  @(posedge pclk)
	ng282<=ng11492;

 always  @(posedge pclk)
	ng287<=ng286;

 always  @(posedge pclk)
	ng394<=ng387;

 always  @(posedge pclk)
	ng523<=ng513;

 always  @(posedge pclk)
	ng489<=ng568;

 always  @(posedge pclk)
	ng479<=ng24216;

 always  @(posedge pclk)
	ng468<=ng24215;

 always  @(posedge pclk)
	ng499<=ng549;

 always  @(posedge pclk)
	ng586<=ng27312;

 always  @(posedge pclk)
	ng617<=ng28349;

 always  @(posedge pclk)
	ng686<=ng28199;

 always  @(posedge pclk)
	ng706<=ng20902;

 always  @(posedge pclk)
	ng716<=ng21009;

 always  @(posedge pclk)
	ng725<=ng20894;

 always  @(posedge pclk)
	ng733<=ng20970;

 always  @(posedge pclk)
	ng823<=ng826;

 always  @(posedge pclk)
	ng832<=ng22054;

 always  @(posedge pclk)
	ng841<=ng22104;

 always  @(posedge pclk)
	ng930<=ng30655;

 always  @(posedge pclk)
	ng903<=ng30249;

 always  @(posedge pclk)
	ng771<=ng26530;

 always  @(posedge pclk)
	ng1030<=ng27262;

 always  @(posedge pclk)
	ng1071<=ng27272;

 always  @(posedge pclk)
	ng1104<=ng29198;

 always  @(posedge pclk)
	ng1136<=ng27763;

 always  @(posedge pclk)
	ng1006<=ng30485;

 always  @(posedge pclk)
	ng1038<=ng1037;

 always  @(posedge pclk)
	ng1059<=ng1071;

 always  @(posedge pclk)
	ng1243<=ng18707;

 always  @(posedge pclk)
	ng1258<=ng1148;

 always  @(posedge pclk)
	ng1253<=ng1252;

 always  @(posedge pclk)
	ng1230<=ng1229;

 always  @(posedge pclk)
	ng1265<=ng27286;

 always  @(posedge pclk)
	ng1219<=ng13430;

 always  @(posedge pclk)
	ng1316<=ng16671;

 always  @(posedge pclk)
	ng1386<=ng20896;

 always  @(posedge pclk)
	ng1395<=ng20950;

 always  @(posedge pclk)
	ng1422<=ng25267;

 always  @(posedge pclk)
	ng1516<=ng22179;

 always  @(posedge pclk)
	ng1557<=ng25235;

 always  @(posedge pclk)
	ng1612<=ng30651;

 always  @(posedge pclk)
	ng1633<=ng30272;

 always  @(posedge pclk)
	ng1606<=ng30650;

 always  @(posedge pclk)
	ng1789<=ng28749;

 always  @(posedge pclk)
	ng1663<=ng11546;

 always  @(posedge pclk)
	ng1672<=ng1671;

 always  @(posedge pclk)
	ng1747<=ng1746;

 always  @(posedge pclk)
	ng1768<=ng1779;

 always  @(posedge pclk)
	ng2225<=ng22098;

 always  @(posedge pclk)
	ng2234<=ng22154;

 always  @(posedge pclk)
	ng2258<=ng2256;

 always  @(posedge pclk)
	ng2513<=ng26823;

 always  @(posedge pclk)
	ng2390<=ng30707;

 always  @(posedge pclk)
	ng2469<=ng2462;

 always  @(posedge pclk)
	ng2597<=ng2587;

 always  @(posedge pclk)
	ng2564<=ng2642;

 always  @(posedge pclk)
	ng2554<=ng24238;

 always  @(posedge pclk)
	ng2543<=ng24237;

 always  @(posedge pclk)
	ng2574<=ng2623;

 always  @(posedge pclk)
	ng2664<=ng24537;

 always  @(posedge pclk)
	ng2682<=ng28363;

 always  @(posedge pclk)
	ng2707<=ng21974;

 always  @(posedge pclk)
	ng2740<=ng26795;

 always  @(posedge pclk)
	ng2775<=ng20981;

 always  @(posedge pclk)
	ng2791<=ng21045;

 always  @(posedge pclk)
	ng2800<=ng20919;

 always  @(posedge pclk)
	ng2802<=ng21046;

 always  @(posedge pclk)
	ng3056<=ng29975;

 always  @(posedge pclk)
	ng3065<=ng30911;

 always  @(posedge pclk)
	ng3078<=ng30987;

 always  @(posedge pclk)
	ng3018<=ng22002;

 always  @(posedge pclk)
	ng2986<=pg5388;

 always  @(posedge pclk)
	pg8271<=ng16857;

 always  @(posedge pclk)
	ng2991<=ng21964;

 always  @(posedge pclk)
	ng2950<=ng19152;

 always  @(posedge pclk)
	ng3191<=pg24734;

 always  @(posedge pclk)
	ng185<=ng29656;

 always  @(posedge pclk)
	ng142<=ng22025;

 always  @(posedge pclk)
	ng150<=ng22063;

 always  @(posedge pclk)
	ng160<=ng22081;

 always  @(posedge pclk)
	ng171<=ng25218;

 always  @(posedge pclk)
	ng186<=ng30261;

 always  @(posedge pclk)
	ng246<=ng30653;

 always  @(posedge pclk)
	ng267<=ng30661;

 always  @(posedge pclk)
	ng361<=ng27265;

 always  @(posedge pclk)
	ng420<=ng29197;

 always  @(posedge pclk)
	ng435<=ng26807;

 always  @(posedge pclk)
	ng316<=ng30700;

 always  @(posedge pclk)
	ng321<=ng29172;

 always  @(posedge pclk)
	ng281<=ng280;

 always  @(posedge pclk)
	ng288<=ng11495;

 always  @(posedge pclk)
	ng352<=ng346;

 always  @(posedge pclk)
	ng395<=ng388;

 always  @(posedge pclk)
	ng569<=ng564;

 always  @(posedge pclk)
	ng566<=ng468;

 always  @(posedge pclk)
	ng478<=ng24207;

 always  @(posedge pclk)
	ng471<=ng24228;

 always  @(posedge pclk)
	ng576<=ng27261;

 always  @(posedge pclk)
	ng583<=ng27295;

 always  @(posedge pclk)
	ng614<=ng28345;

 always  @(posedge pclk)
	ng493<=ng26545;

 always  @(posedge pclk)
	ng534<=ng13415;

 always  @(posedge pclk)
	ng692<=ng28668;

 always  @(posedge pclk)
	ng709<=ng20922;

 always  @(posedge pclk)
	ng713<=ng20989;

 always  @(posedge pclk)
	ng727<=ng20881;

 always  @(posedge pclk)
	ng731<=ng20992;

 always  @(posedge pclk)
	ng819<=ng22145;

 always  @(posedge pclk)
	ng829<=ng22040;

 always  @(posedge pclk)
	ng843<=ng22088;

 always  @(posedge pclk)
	ng864<=ng25231;

 always  @(posedge pclk)
	ng933<=ng30662;

 always  @(posedge pclk)
	ng948<=ng30271;

 always  @(posedge pclk)
	ng960<=ng30682;

 always  @(posedge pclk)
	ng1041<=ng27257;

 always  @(posedge pclk)
	ng1060<=ng27283;

 always  @(posedge pclk)
	ng1114<=ng28747;

 always  @(posedge pclk)
	ng1128<=ng26814;

 always  @(posedge pclk)
	ng1005<=ng30470;

 always  @(posedge pclk)
	ng1039<=ng1033;

 always  @(posedge pclk)
	ng1068<=ng1067;

 always  @(posedge pclk)
	ng1084<=ng1078;

 always  @(posedge pclk)
	ng1257<=ng1256;

 always  @(posedge pclk)
	ng1254<=ng1158;

 always  @(posedge pclk)
	ng1167<=ng23110;

 always  @(posedge pclk)
	ng1261<=ng27299;

 always  @(posedge pclk)
	ng1220<=ng13431;

 always  @(posedge pclk)
	ng1319<=ng21969;

 always  @(posedge pclk)
	ng1372<=ng27718;

 always  @(posedge pclk)
	ng1394<=ng20927;

 always  @(posedge pclk)
	ng1401<=ng20994;

 always  @(posedge pclk)
	ng1412<=ng20883;

 always  @(posedge pclk)
	ng1558<=ng25243;

 always  @(posedge pclk)
	ng1576<=ng30683;

 always  @(posedge pclk)
	ng1588<=ng30299;

 always  @(posedge pclk)
	ng1603<=ng30644;

 always  @(posedge pclk)
	ng1727<=ng27287;

 always  @(posedge pclk)
	ng1664<=ng1663;

 always  @(posedge pclk)
	ng1679<=ng26130;

 always  @(posedge pclk)
	ng1738<=ng1750;

 always  @(posedge pclk)
	ng1764<=ng1763;

 always  @(posedge pclk)
	ng2448<=ng27323;

 always  @(posedge pclk)
	ng2516<=ng26826;

 always  @(posedge pclk)
	ng2393<=ng30505;

 always  @(posedge pclk)
	ng2470<=ng2463;

 always  @(posedge pclk)
	ng2643<=ng2638;

 always  @(posedge pclk)
	ng2640<=ng2543;

 always  @(posedge pclk)
	ng2553<=ng24226;

 always  @(posedge pclk)
	ng2546<=ng24250;

 always  @(posedge pclk)
	ng2650<=ng27310;

 always  @(posedge pclk)
	ng2667<=ng24547;

 always  @(posedge pclk)
	ng2604<=ng13459;

 always  @(posedge pclk)
	ng2714<=ng20789;

 always  @(posedge pclk)
	ng2753<=ng27243;

 always  @(posedge pclk)
	ng2778<=ng21004;

 always  @(posedge pclk)
	ng2788<=ng21027;

 always  @(posedge pclk)
	ng2796<=ng21094;

 always  @(posedge pclk)
	ng2806<=ng21029;

 always  @(posedge pclk)
	ng3080<=ng20497;

 always  @(posedge pclk)
	ng3057<=ng29976;

 always  @(posedge pclk)
	ng3068<=ng30914;

 always  @(posedge pclk)
	ng3075<=ng30984;

 always  @(posedge pclk)
	ng3024<=ng26786;

 always  @(posedge pclk)
	ng2987<=pg16496;

 always  @(posedge pclk)
	ng2992<=ng21966;

 always  @(posedge pclk)
	pg8261<=ng18837;

 always  @(posedge pclk)
	ng2883<=ng20825;

 always  @(posedge pclk)
	ng3128<=ng29166;

 always  @(posedge pclk)
	ng3147<=pg26135;

 always  @(posedge pclk)
	ng143<=ng22027;

 always  @(posedge pclk)
	ng152<=ng22048;

 always  @(posedge pclk)
	ng161<=ng22102;

 always  @(posedge pclk)
	ng173<=ng25212;

 always  @(posedge pclk)
	ng189<=ng30267;

 always  @(posedge pclk)
	ng243<=ng30646;

 always  @(posedge pclk)
	ng61<=ng29109;

 always  @(posedge pclk)
	ng384<=ng27260;

 always  @(posedge pclk)
	ng417<=ng29194;

 always  @(posedge pclk)
	ng438<=ng26805;

 always  @(posedge pclk)
	ng315<=ng30699;

 always  @(posedge pclk)
	ng403<=ng26655;

 always  @(posedge pclk)
	ng280<=ng11491;

 always  @(posedge pclk)
	ng289<=ng288;

 always  @(posedge pclk)
	ng351<=ng350;

 always  @(posedge pclk)
	ng396<=ng395;

 always  @(posedge pclk)
	ng564<=ng455;

 always  @(posedge pclk)
	ng567<=ng566;

 always  @(posedge pclk)
	ng477<=ng24178;

 always  @(posedge pclk)
	ng528<=ng12457;

 always  @(posedge pclk)
	ng559<=ng558;

 always  @(posedge pclk)
	ng581<=ng27311;

 always  @(posedge pclk)
	ng602<=ng24519;

 always  @(posedge pclk)
	ng496<=ng26553;

 always  @(posedge pclk)
	ng533<=ng13414;

 always  @(posedge pclk)
	ng699<=ng20875;

 always  @(posedge pclk)
	ng708<=ng20903;

 always  @(posedge pclk)
	ng717<=ng20968;

 always  @(posedge pclk)
	ng726<=ng20876;

 always  @(posedge pclk)
	ng735<=ng25260;

 always  @(posedge pclk)
	ng818<=ng22126;

 always  @(posedge pclk)
	ng833<=ng22034;

 always  @(posedge pclk)
	ng842<=ng22068;

 always  @(posedge pclk)
	ng851<=ng22129;

 always  @(posedge pclk)
	ng891<=ng30286;

 always  @(posedge pclk)
	ng945<=ng30265;

 always  @(posedge pclk)
	ng780<=ng25042;

 always  @(posedge pclk)
	ng740<=ng29580;

 always  @(posedge pclk)
	ng1063<=ng27297;

 always  @(posedge pclk)
	ng1110<=ng29209;

 always  @(posedge pclk)
	ng1131<=ng26818;

 always  @(posedge pclk)
	ng1004<=ng30705;

 always  @(posedge pclk)
	ng1040<=ng1039;

 always  @(posedge pclk)
	ng1067<=ng1060;

 always  @(posedge pclk)
	ng1011<=ng1084;

 always  @(posedge pclk)
	ng1256<=ng1145;

 always  @(posedge pclk)
	ng1176<=ng1254;

 always  @(posedge pclk)
	ng1166<=ng24223;

 always  @(posedge pclk)
	ng1228<=ng1221;

 always  @(posedge pclk)
	ng1222<=ng13432;

 always  @(posedge pclk)
	ng1326<=ng20717;

 always  @(posedge pclk)
	ng1378<=ng28321;

 always  @(posedge pclk)
	ng1390<=ng20949;

 always  @(posedge pclk)
	ng1399<=ng21015;

 always  @(posedge pclk)
	ng1408<=ng21070;

 always  @(posedge pclk)
	ng1556<=ng25249;

 always  @(posedge pclk)
	ng1618<=ng30663;

 always  @(posedge pclk)
	ng1591<=ng30302;

 always  @(posedge pclk)
	ng1645<=ng30288;

 always  @(posedge pclk)
	ng1457<=ng26531;

 always  @(posedge pclk)
	ng1665<=ng11547;

 always  @(posedge pclk)
	ng1686<=ng28903;

 always  @(posedge pclk)
	ng1745<=ng1738;

 always  @(posedge pclk)
	ng1763<=ng1757;

 always  @(posedge pclk)
	ng2498<=ng29226;

 always  @(posedge pclk)
	ng2519<=ng26827;

 always  @(posedge pclk)
	ng2392<=ng30566;

 always  @(posedge pclk)
	ng2471<=ng2470;

 always  @(posedge pclk)
	ng2638<=ng2530;

 always  @(posedge pclk)
	ng2641<=ng2640;

 always  @(posedge pclk)
	ng2552<=ng24214;

 always  @(posedge pclk)
	ng2602<=ng12499;

 always  @(posedge pclk)
	ng2633<=ng2632;

 always  @(posedge pclk)
	ng2565<=ng26575;

 always  @(posedge pclk)
	ng2605<=ng13460;

 always  @(posedge pclk)
	ng2733<=ng20375;

 always  @(posedge pclk)
	ng2760<=ng27724;

 always  @(posedge pclk)
	ng2780<=ng20982;

 always  @(posedge pclk)
	ng2789<=ng21044;

 always  @(posedge pclk)
	ng2798<=ng21082;

 always  @(posedge pclk)
	ng2807<=ng21047;

 always  @(posedge pclk)
	ng3079<=ng20884;

 always  @(posedge pclk)
	ng3058<=ng29977;

 always  @(posedge pclk)
	ng3067<=ng30913;

 always  @(posedge pclk)
	ng3076<=ng30985;

 always  @(posedge pclk)
	ng3010<=ng26031;

 always  @(posedge pclk)
	pg8275<=ng16824;

 always  @(posedge pclk)
	pg8267<=ng16566;

 always  @(posedge pclk)
	pg8259<=ng18868;

 always  @(posedge pclk)
	ng809<=pg4090;

 always  @(posedge pclk)
	pg7334<=ng20417;

 always  @(posedge pclk)
	ng113<=pg8023;

 always  @(posedge pclk)
	ng2200<=ng18885;

 always  @(posedge pclk)
	ng3084<=ng18782;

 always  @(posedge pclk)
	ng3059<=ng29978;

 always  @(posedge pclk)
	ng3070<=ng30940;

 always  @(posedge pclk)
	pg4323<=ng19173;

 always  @(posedge pclk)
	ng789<=pg6895;

 always  @(posedge pclk)
	pg8175<=ng19149;

 always  @(posedge pclk)
	ng2857<=pg8096;

 always  @(posedge pclk)
	ng3085<=ng17222;

 always  @(posedge pclk)
	ng3060<=ng29979;

 always  @(posedge pclk)
	ng3069<=ng30915;

 always  @(posedge pclk)
	ng805<=pg4323;

 always  @(posedge pclk)
	pg7519<=ng21878;

 always  @(posedge pclk)
	ng117<=pg4321;

 always  @(posedge pclk)
	pg8096<=ng20874;

 always  @(posedge pclk)
	ng3086<=ng17225;

 always  @(posedge pclk)
	ng2997<=ng30989;

 always  @(posedge pclk)
	ng3032<=ng25202;

 always  @(posedge pclk)
	pg8021<=pg51;

 always  @(posedge pclk)
	pg4590<=ng19184;

 always  @(posedge pclk)
	ng785<=pg7334;

 always  @(posedge pclk)
	pg8023<=ng19144;

 always  @(posedge pclk)
	ng97<=pg4450;

 always  @(posedge pclk)
	ng3087<=ng17234;

 always  @(posedge pclk)
	ng2993<=ng25265;

 always  @(posedge pclk)
	ng3036<=ng24446;

 always  @(posedge pclk)
	ng2908<=ng26798;

 always  @(posedge pclk)
	ng2935<=pg3228;

 always  @(posedge pclk)
	ng2969<=pg3218;

 always  @(posedge pclk)
	ng1481<=ng18852;

 always  @(posedge pclk)
	ng3091<=ng17224;

 always  @(posedge pclk)
	ng1570<=ng30287;

 always  @(posedge pclk)
	ng1670<=ng1669;

 always  @(posedge pclk)
	ng1734<=ng1733;

 always  @(posedge pclk)
	ng2210<=ng22193;

 always  @(posedge pclk)
	ng2227<=ng22099;

 always  @(posedge pclk)
	pg8269<=ng16835;

 always  @(posedge pclk)
	pg8260<=ng18804;

 always  @(posedge pclk)
	ng2912<=ng21989;

 always  @(posedge pclk)
	ng2934<=pg3212;

 always  @(posedge pclk)
	ng2972<=pg3217;

 always  @(posedge pclk)
	ng1486<=ng18835;

 always  @(posedge pclk)
	ng3092<=ng17228;

 always  @(posedge pclk)
	ng1627<=ng30671;

 always  @(posedge pclk)
	ng1671<=ng2877;

 always  @(posedge pclk)
	ng1733<=ng1727;

 always  @(posedge pclk)
	ng2208<=ng22200;

 always  @(posedge pclk)
	ng2223<=ng22115;

 always  @(posedge pclk)
	pg8270<=ng16851;

 always  @(posedge pclk)
	pg8263<=ng18755;

 always  @(posedge pclk)
	ng2917<=ng23357;

 always  @(posedge pclk)
	ng2941<=pg3226;

 always  @(posedge pclk)
	ng2963<=pg3220;

 always  @(posedge pclk)
	ng1491<=ng18821;

 always  @(posedge pclk)
	ng1639<=ng30273;

 always  @(posedge pclk)
	ng1761<=ng1754;

 always  @(posedge pclk)
	ng1937<=ng18743;

 always  @(posedge pclk)
	ng2218<=ng22045;

 always  @(posedge pclk)
	ng2226<=ng22138;

 always  @(posedge pclk)
	ng2524<=ng27769;

 always  @(posedge pclk)
	ng2924<=ng24476;

 always  @(posedge pclk)
	ng2938<=pg3227;

 always  @(posedge pclk)
	ng2966<=pg3219;

 always  @(posedge pclk)
	ng1496<=ng18803;

 always  @(posedge pclk)
	ng1462<=ng25938;

 always  @(posedge pclk)
	ng1762<=ng1761;

 always  @(posedge pclk)
	ng1934<=ng21845;

 always  @(posedge pclk)
	ng2219<=ng22060;

 always  @(posedge pclk)
	ng2228<=ng22116;

 always  @(posedge pclk)
	ng2502<=ng28774;

 always  @(posedge pclk)
	ng2920<=ng25199;

 always  @(posedge pclk)
	ng2947<=pg3224;

 always  @(posedge pclk)
	ng2981<=pg3214;

 always  @(posedge pclk)
	pg8251<=ng19154;

 always  @(posedge pclk)
	ng793<=pg6442;

 always  @(posedge pclk)
	pg4321<=ng19172;

 always  @(posedge pclk)
	ng1724<=ng27274;

 always  @(posedge pclk)
	ng1952<=ng1842;

 always  @(posedge pclk)
	ng1836<=ng23400;

 always  @(posedge pclk)
	ng2085<=ng20936;

 always  @(posedge pclk)
	ng2093<=ng21039;

 always  @(posedge pclk)
	ng2107<=ng20917;

 always  @(posedge pclk)
	ng2118<=ng22249;

 always  @(posedge pclk)
	ng2451<=ng27334;

 always  @(posedge pclk)
	ng2984<=ng16181;

 always  @(posedge pclk)
	ng2944<=pg3225;

 always  @(posedge pclk)
	ng2874<=pg3213;

 always  @(posedge pclk)
	ng2877<=ng21880;

 always  @(posedge pclk)
	pg6895<=ng20376;

 always  @(posedge pclk)
	ng121<=pg4088;

 always  @(posedge pclk)
	ng1772<=ng27330;

 always  @(posedge pclk)
	ng1953<=ng1952;

 always  @(posedge pclk)
	ng1869<=ng23137;

 always  @(posedge pclk)
	ng2086<=ng20954;

 always  @(posedge pclk)
	ng2095<=ng21020;

 always  @(posedge pclk)
	ng2105<=ng20937;

 always  @(posedge pclk)
	ng2114<=ng25279;

 always  @(posedge pclk)
	ng2257<=ng2258;

 always  @(posedge pclk)
	ng2985<=ng16132;

 always  @(posedge pclk)
	ng2956<=pg3222;

 always  @(posedge pclk)
	ng2975<=pg3216;

 always  @(posedge pclk)
	ng1471<=ng18883;

 always  @(posedge pclk)
	ng101<=pg4200;

 always  @(posedge pclk)
	ng2170<=ng18836;

 always  @(posedge pclk)
	ng1810<=ng26811;

 always  @(posedge pclk)
	ng1846<=ng24218;

 always  @(posedge pclk)
	ng1938<=ng13182;

 always  @(posedge pclk)
	ng2084<=ng20977;

 always  @(posedge pclk)
	ng2098<=ng21040;

 always  @(posedge pclk)
	ng2102<=ng21080;

 always  @(posedge pclk)
	ng2116<=ng25271;

 always  @(posedge pclk)
	ng2151<=ng26532;

 always  @(posedge pclk)
	ng2953<=pg3223;

 always  @(posedge pclk)
	ng2978<=pg3215;

 always  @(posedge pclk)
	ng1476<=ng18866;

 always  @(posedge pclk)
	pg4450<=ng19178;

 always  @(posedge pclk)
	ng2175<=ng18867;

 always  @(posedge pclk)
	ng1694<=ng29617;

 always  @(posedge pclk)
	ng1849<=ng24230;

 always  @(posedge pclk)
	ng1880<=ng1929;

 always  @(posedge pclk)
	ng2088<=ng20955;

 always  @(posedge pclk)
	ng2097<=ng21021;

 always  @(posedge pclk)
	ng2106<=ng20900;

 always  @(posedge pclk)
	ng2115<=ng25268;

 always  @(posedge pclk)
	ng2336<=ng30291;

 always  @(posedge pclk)
	ng2929<=pg8021;

 always  @(posedge pclk)
	ng2962<=pg3232;

 always  @(posedge pclk)
	ng801<=pg4590;

 always  @(posedge pclk)
	pg8249<=ng19153;

 always  @(posedge pclk)
	ng105<=pg3993;

 always  @(posedge pclk)
	ng2180<=ng18906;

 always  @(posedge pclk)
	ng2165<=ng18957;

 always  @(posedge pclk)
	ng1702<=ng29184;

 always  @(posedge pclk)
	ng1963<=ng27332;

 always  @(posedge pclk)
	ng1994<=ng28357;

 always  @(posedge pclk)
	ng1997<=ng28362;

 always  @(posedge pclk)
	ng1905<=pg16399;

 always  @(posedge pclk)
	ng2010<=ng16692;

 always  @(posedge pclk)
	ng2072<=ng28325;

 always  @(posedge pclk)
	ng2279<=ng30301;

 always  @(posedge pclk)
	ng2879<=ng12433;

 always  @(posedge pclk)
	ng2959<=pg3221;

 always  @(posedge pclk)
	pg6225<=ng20310;

 always  @(posedge pclk)
	ng2873<=pg7519;

 always  @(posedge pclk)
	pg4200<=ng19167;

 always  @(posedge pclk)
	ng2185<=ng18942;

 always  @(posedge pclk)
	ng2878<=ng21882;

 always  @(posedge pclk)
	ng1661<=ng11545;

 always  @(posedge pclk)
	ng1961<=ng27340;

 always  @(posedge pclk)
	ng1982<=ng24545;

 always  @(posedge pclk)
	ng2000<=ng28366;

 always  @(posedge pclk)
	pg16399<=ng28990;

 always  @(posedge pclk)
	ng2039<=ng20353;

 always  @(posedge pclk)
	ng2066<=ng27722;

 always  @(posedge pclk)
	ng2267<=ng30300;

 always  @(posedge pclk)
	ng1506<=ng18754;

 always  @(posedge pclk)
	pg4090<=ng19163;

 always  @(posedge pclk)
	ng797<=pg6225;

 always  @(posedge pclk)
	pg4088<=ng19162;

 always  @(posedge pclk)
	ng109<=pg8175;

 always  @(posedge pclk)
	ng2190<=ng18968;

 always  @(posedge pclk)
	ng3210<=ng18669;

 always  @(posedge pclk)
	ng1985<=ng28352;

 always  @(posedge pclk)
	ng1910<=ng13443;

 always  @(posedge pclk)
	ng1918<=ng24083;

 always  @(posedge pclk)
	ng2059<=ng27682;

 always  @(posedge pclk)
	ng2249<=ng25246;

 always  @(posedge pclk)
	ng1501<=ng18781;

 always  @(posedge pclk)
	ng813<=pg8251;

 always  @(posedge pclk)
	pg6442<=ng20343;

 always  @(posedge pclk)
	ng125<=pg8249;

 always  @(posedge pclk)
	pg3993<=ng19157;

 always  @(posedge pclk)
	ng2195<=ng18975;

 always  @(posedge pclk)
	ng3211<=ng18719;

 always  @(posedge pclk)
	ng1988<=ng28356;

 always  @(posedge pclk)
	ng1909<=ng13442;

 always  @(posedge pclk)
	ng1921<=ng13450;

 always  @(posedge pclk)
	ng2046<=ng26789;

 always  @(posedge pclk)
	ng2236<=ng22155;

 assign pg24734 = ( ng17973 ) | ( (~ ng3123)  &  (~ ng8381)  &  (~ wire30893) ) ;
 assign pg26135 = ( wire36306 ) | ( wire36307 ) | ( wire36311 ) ;
 assign pg25435 = ( wire6564 ) | ( wire34622 ) ;
 assign pg16496 = ( (~ ng2987) ) | ( pg5388  &  (~ ng2986) ) ;
 assign pg27380 = ( wire7046 ) | ( wire7048 ) | ( wire34087 ) ;
 assign pg26149 = ( wire30913 ) | ( wire30914 ) | ( wire30918 ) ;
 assign pg25420 = ( (~ pg3233) ) | ( pg3230 ) | ( ng3126  &  wire3217 ) ;
 assign pg25442 = ( (~ pg3233) ) | ( pg3230 ) | ( ng3124  &  wire3217 ) ;
 assign pg25489 = ( wire3034 ) | ( wire3035 ) | ( wire3036 ) | ( wire3037 ) ;
 assign pg26104 = ( wire34973 ) | ( wire34974 ) | ( wire34978 ) ;
 assign ng25450 = ( ng3097  &  (~ ng1309) ) | ( ng544  &  ng1309  &  ng499 ) ;
 assign ng30801 = ( ng3108  &  (~ ng1315) ) | ( ng1315  &  ng30072 ) ;
 assign ng17341 = ( ng3185  &  (~ ng1312) ) | ( ng1312  &  ng2574 ) ;
 assign ng22030 = ( ng141  &  (~ ng853) ) | ( ng141  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng105) ) ;
 assign ng22064 = ( ng155  &  (~ ng823) ) | ( ng155  &  (~ ng2257) ) | ( ng823  &  (~ ng121)  &  ng2257 ) ;
 assign ng30258 = ( ng258  &  (~ ng826) ) | ( ng826  &  ng29671 ) ;
 assign ng26529 = ( ng83  &  ng25932 ) | ( ng83  &  (~ ng88)  &  (~ ng17031) ) | ( (~ ng83)  &  (~ ng25932)  &  ng88  &  (~ ng17031) ) ;
 assign ng27256 = ( ng369  &  (~ ng826) ) | ( ng369  &  wire3290 ) | ( ng826  &  (~ wire3290)  &  (~ ng21976) ) ;
 assign ng28744 = ( ng414  &  (~ ng853) ) | ( ng853  &  ng27528 ) ;
 assign ng26808 = ( ng441  &  (~ ng823) ) | ( ng823  &  wire3156 ) ;
 assign ng30455 = ( ng318  &  (~ ng826) ) | ( ng826  &  ng29912 ) ;
 assign ng11510 = ( (~ ng121) ) ;
 assign ng18678 = ( (~ ng554)  &  ng1315 ) | ( ng557  &  (~ ng1315) ) ;
 assign ng24174 = ( ng461  &  (~ ng853) ) | ( ng853  &  (~ ng11624)  &  wire31336 ) ;
 assign ng27279 = ( ng575  &  (~ ng1315) ) | ( ng575  &  (~ ng22578) ) | ( ng1315  &  ng22578  &  (~ ng23360) ) ;
 assign ng24498 = ( wire9005 ) | ( ng590  &  (~ ng1312) ) ;
 assign ng26541 = ( ng490  &  (~ ng1309) ) | ( ng1309  &  ng12245  &  wire3444 ) ;
 assign ng24426 = ( ng646  &  ng10677  &  (~ wire31591) ) | ( ng646  &  ng10677  &  (~ wire31592) ) | ( (~ ng646)  &  ng10677  &  wire31591  &  wire31592 ) ;
 assign ng20892 = ( ng703  &  ng13113 ) | ( (~ ng633)  &  (~ ng13113) ) ;
 assign ng20946 = ( ng714  &  ng13123 ) | ( (~ ng672)  &  (~ ng13123) ) ;
 assign ng21051 = ( ng722  &  ng11721 ) | ( (~ ng686)  &  (~ ng11721) ) ;
 assign ng25262 = ( ng736  &  ng13113 ) | ( (~ ng13113)  &  wire31760 ) | ( (~ ng13113)  &  wire31761 ) ;
 assign ng22146 = ( ng821  &  (~ ng826) ) | ( ng821  &  (~ ng2257) ) | ( ng826  &  (~ ng789)  &  ng2257 ) ;
 assign ng22066 = ( ng835  &  (~ ng853) ) | ( ng835  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng801) ) ;
 assign ng22128 = ( ng849  &  ng15950 ) | ( (~ ng15950)  &  wire31770 ) | ( (~ ng15950)  &  wire31771 ) ;
 assign ng25223 = ( ng863  &  (~ ng13110) ) | ( ng863  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng785) ) ;
 assign ng30654 = ( ng924  &  (~ ng853) ) | ( ng853  &  wire32135 ) | ( ng853  &  wire32136 ) ;
 assign ng30264 = ( ng939  &  (~ ng823) ) | ( ng823  &  ng29672 ) ;
 assign ng30670 = ( ng954  &  (~ ng826) ) | ( ng826  &  wire32160 ) | ( ng826  &  wire32161 ) ;
 assign ng29354 = ( (~ ng744)  &  (~ ng17031)  &  ng26878 ) | ( ng744  &  (~ ng17031)  &  (~ ng26878) ) ;
 assign ng27284 = ( ng1085  &  (~ ng826) ) | ( ng1085  &  wire3293 ) | ( ng826  &  (~ wire3293)  &  (~ ng22005) ) ;
 assign ng28767 = ( wire8488 ) | ( wire32246 ) ;
 assign ng29612 = ( wire8484 ) | ( ng1000  &  (~ ng823) ) ;
 assign ng26661 = ( wire8482 ) | ( ng1090  &  (~ ng826) ) | ( ng1090  &  (~ ng2257) ) ;
 assign ng11519 = ( (~ ng797) ) ;
 assign ng26183 = ( wire32253 ) | ( ng986  &  ng21346  &  ng823 ) ;
 assign ng23081 = ( ng1173  &  (~ ng826) ) | ( ng826  &  (~ wire32262)  &  (~ wire32263) ) ;
 assign ng23039 = ( ng1151  &  (~ ng853) ) | ( ng853  &  wire32219 ) | ( ng853  &  wire32220 ) ;
 assign ng27328 = ( ng1267  &  (~ ng1315) ) | ( ng1267  &  (~ ng22615) ) | ( ng1315  &  ng22615  &  (~ ng23377) ) ;
 assign ng28355 = ( ng1303  &  (~ ng1312) ) | ( ng1312  &  ng27157 ) ;
 assign ng26781 = ( (~ ng23979)  &  wire32578 ) | ( (~ ng26666)  &  (~ ng23979)  &  wire32576 ) ;
 assign ng20926 = ( ng1392  &  ng13126 ) | ( (~ ng1339)  &  (~ ng13126) ) ;
 assign ng20995 = ( ng1403  &  ng13134 ) | ( (~ ng1352)  &  (~ ng13134) ) ;
 assign ng20913 = ( ng1411  &  ng11726 ) | ( (~ ng1378)  &  (~ ng11726) ) ;
 assign ng22247 = ( ng1425  &  (~ ng1312) ) | ( ng1425  &  (~ ng1316) ) | ( (~ ng1316)  &  (~ ng13126) ) ;
 assign ng22044 = ( ng1527  &  (~ ng826) ) | ( ng1527  &  (~ ng2257) ) | ( ng826  &  (~ ng1486)  &  ng2257 ) ;
 assign ng22130 = ( ng1535  &  (~ ng853) ) | ( ng1535  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng1501) ) ;
 assign ng25224 = ( ng1552  &  (~ ng13110) ) | ( ng1552  &  (~ ng823) ) | ( ng13110  &  ng823  &  wire3921 ) ;
 assign ng30281 = ( ng1642  &  (~ ng823) ) | ( ng823  &  ng29680 ) ;
 assign ng27129 = ( wire7941 ) | ( (~ ng26531)  &  wire32977 ) ;
 assign ng27288 = ( ng1739  &  (~ ng823) ) | ( ng1739  &  wire3309 ) | ( ng823  &  (~ ng21996)  &  (~ wire3309) ) ;
 assign ng29205 = ( ng1798  &  (~ ng826) ) | ( ng826  &  ng11952  &  ng27567 ) | ( ng826  &  (~ ng11952)  &  (~ ng27567) ) ;
 assign ng26824 = ( ng1825  &  (~ ng853) ) | ( ng853  &  wire3159 ) ;
 assign ng30503 = ( ng1700  &  (~ ng823) ) | ( ng823  &  wire7829 ) | ( ng823  &  wire7830 ) ;
 assign ng18794 = ( ng1890  &  (~ ng1315) ) | ( ng1315  &  ng1937 ) ;
 assign ng24208 = ( ng1858  &  (~ ng826) ) | ( ng826  &  ng11666  &  wire32944 ) ;
 assign ng27306 = ( ng1959  &  (~ ng1309) ) | ( ng1959  &  (~ ng22651) ) | ( ng1309  &  ng22651  &  (~ ng22093) ) ;
 assign ng24534 = ( wire7732 ) | ( ng1973  &  (~ ng1315) ) ;
 assign ng28361 = ( wire7633 ) | ( ng1991  &  (~ ng1315) ) ;
 assign ng13445 = ( (~ ng1662) ) ;
 assign ng23339 = ( wire7627 ) | ( (~ ng21972)  &  wire33416 ) ;
 assign ng20916 = ( ng2082  &  ng13142 ) | ( (~ ng2013)  &  (~ ng13142) ) ;
 assign ng21019 = ( ng2090  &  ng11730 ) | ( (~ ng2040)  &  (~ ng11730) ) ;
 assign ng21072 = ( ng2104  &  ng13137 ) | ( (~ ng2066)  &  (~ ng13137) ) ;
 assign ng22172 = ( ng2237  &  ng15950 ) | ( (~ ng15950)  &  wire33428 ) | ( (~ ng15950)  &  wire33429 ) ;
 assign ng25247 = ( ng2251  &  (~ ng13110) ) | ( ng2251  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng2165) ) ;
 assign ng30672 = ( ng2312  &  (~ ng853) ) | ( ng853  &  wire33799 ) | ( ng853  &  wire33800 ) ;
 assign ng30282 = ( ng2327  &  (~ ng823) ) | ( ng823  &  ng29681 ) ;
 assign ng30686 = ( ng2342  &  (~ ng826) ) | ( ng826  &  wire33823 ) | ( ng826  &  wire33824 ) ;
 assign ng29357 = ( (~ ng2124)  &  (~ ng17031)  &  ng26897 ) | ( ng2124  &  (~ ng17031)  &  (~ ng26897) ) ;
 assign ng27322 = ( ng2436  &  (~ ng853) ) | ( ng2436  &  wire3313 ) | ( ng853  &  (~ wire3313)  &  (~ ng22009) ) ;
 assign ng29221 = ( ng2495  &  (~ ng823) ) | ( ng823  &  ng12005  &  ng27577 ) | ( ng823  &  (~ ng12005)  &  (~ ng27577) ) ;
 assign ng27767 = ( ng2523  &  (~ ng826) ) | ( ng826  &  (~ ng24038)  &  wire33948 ) | ( ng2523  &  (~ ng24038)  &  (~ wire33948) ) ;
 assign ng18780 = ( (~ ng2628)  &  ng1315 ) | ( ng2631  &  (~ ng1315) ) ;
 assign ng24209 = ( ng2536  &  (~ ng853) ) | ( ng853  &  (~ ng11678)  &  wire33862 ) ;
 assign ng27336 = ( ng2649  &  (~ ng1315) ) | ( ng2649  &  (~ ng22687) ) | ( ng1315  &  ng22687  &  (~ ng23381) ) ;
 assign ng20962 = ( ng2772  &  ng11733 ) | ( (~ ng2714)  &  (~ ng11733) ) ;
 assign ng21026 = ( ng2786  &  ng13145 ) | ( (~ ng2734)  &  (~ ng13145) ) ;
 assign ng21075 = ( ng2797  &  ng13146 ) | ( (~ ng2760)  &  (~ ng13146) ) ;
 assign ng21063 = ( ng2805  &  wire3216 ) | ( (~ wire3216)  &  wire33977 ) | ( (~ wire3216)  &  wire33978 ) ;
 assign ng29454 = ( wire3425 ) | ( wire7057 ) | ( wire7058 ) ;
 assign ng25451 = ( ng3098  &  (~ ng1312) ) | ( ng1312  &  ng21851 ) ;
 assign ng30798 = ( ng3107  &  (~ ng1312) ) | ( ng1312  &  ng30072 ) ;
 assign ng17429 = ( ng3088  &  (~ ng1315) ) | ( ng1315  &  ng2574 ) ;
 assign ng22028 = ( ng145  &  (~ ng826) ) | ( ng145  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng109) ) ;
 assign ng22049 = ( ng154  &  (~ ng826) ) | ( ng154  &  (~ ng2257) ) | ( ng826  &  (~ ng121)  &  ng2257 ) ;
 assign ng30263 = ( ng261  &  (~ ng823) ) | ( ng823  &  ng29671 ) ;
 assign ng25932 = ( ng88  &  (~ ng92)  &  ng13165 ) | ( (~ ng88)  &  ng92  &  ng17197 ) | ( ng88  &  (~ ng92)  &  ng17197 ) | ( ng88  &  ng13165  &  (~ ng17197) ) ;
 assign ng27259 = ( ng358  &  (~ ng823) ) | ( ng358  &  wire3290 ) | ( ng823  &  (~ wire3290)  &  (~ ng21976) ) ;
 assign ng28735 = ( ng411  &  (~ ng823) ) | ( ng823  &  ng27528 ) ;
 assign ng26812 = ( ng444  &  (~ ng853) ) | ( ng853  &  wire3156 ) ;
 assign ng30702 = ( ng317  &  (~ ng853) ) | ( ng853  &  ng30030 ) ;
 assign ng11494 = ( (~ ng101) ) ;
 assign ng21842 = ( wire3142 ) | ( ng554  &  (~ ng1315) ) ;
 assign ng23399 = ( ng458  &  (~ ng823) ) | ( ng823  &  (~ ng11624)  &  wire31336 ) ;
 assign ng27268 = ( ng577  &  (~ ng1312) ) | ( ng577  &  (~ ng22578) ) | ( ng1312  &  ng22578  &  (~ ng23360) ) ;
 assign ng24507 = ( wire7014 ) | ( ng593  &  (~ ng1315) ) ;
 assign ng28348 = ( wire6923 ) | ( ng611  &  (~ ng1315) ) ;
 assign ng25185 = ( wire6921 ) | ( wire6922 ) ;
 assign ng20880 = ( ng702  &  ng13123 ) | ( (~ ng633)  &  (~ ng13123) ) ;
 assign ng20967 = ( ng715  &  ng13113 ) | ( (~ ng672)  &  (~ ng13113) ) ;
 assign ng21032 = ( ng724  &  ng13113 ) | ( (~ ng686)  &  (~ ng13113) ) ;
 assign ng25266 = ( ng734  &  ng11721 ) | ( (~ ng11721)  &  wire31760 ) | ( (~ ng11721)  &  wire31761 ) ;
 assign ng22162 = ( ng817  &  (~ ng853) ) | ( ng817  &  (~ ng2257) ) | ( ng853  &  (~ ng785)  &  ng2257 ) ;
 assign ng22056 = ( ng839  &  (~ ng826) ) | ( ng839  &  (~ ng2257) ) | ( ng826  &  (~ ng805)  &  ng2257 ) ;
 assign ng22106 = ( ng848  &  ng15970 ) | ( (~ ng15970)  &  wire31770 ) | ( (~ ng15970)  &  wire31771 ) ;
 assign ng30648 = ( ng921  &  (~ ng823) ) | ( ng823  &  wire32135 ) | ( ng823  &  wire32136 ) ;
 assign ng30676 = ( ng882  &  (~ ng826) ) | ( ng826  &  wire34273 ) | ( ng826  &  wire34274 ) ;
 assign ng30259 = ( ng936  &  (~ ng826) ) | ( ng826  &  ng29672 ) ;
 assign ng30677 = ( ng957  &  (~ ng823) ) | ( ng823  &  wire32160 ) | ( ng823  &  wire32161 ) ;
 assign ng29110 = ( (~ ng26878)  &  wire34283 ) | ( (~ ng28635)  &  (~ ng26878)  &  wire34281 ) ;
 assign ng27298 = ( ng1075  &  (~ ng823) ) | ( ng1075  &  wire3293 ) | ( ng823  &  (~ wire3293)  &  (~ ng22005) ) ;
 assign ng28759 = ( wire6883 ) | ( wire34284 ) ;
 assign ng29616 = ( wire6881 ) | ( ng1001  &  (~ ng853) ) ;
 assign ng29179 = ( wire34295 ) | ( ng853  &  (~ ng27850)  &  wire34293 ) ;
 assign ng19024 = ( (~ wire32219)  &  (~ wire32220) ) ;
 assign ng26120 = ( wire34371 ) | ( wire34372 ) | ( wire34373 ) | ( wire34374 ) ;
 assign ng23111 = ( ng1174  &  (~ ng823) ) | ( ng823  &  (~ wire32262)  &  (~ wire32263) ) ;
 assign ng23014 = ( ng1171  &  (~ ng823) ) | ( ng823  &  wire32219 ) | ( ng823  &  wire32220 ) ;
 assign ng13171 = ( wire34385 ) | ( wire34386 ) ;
 assign ng27315 = ( ng1269  &  (~ ng1312) ) | ( ng1269  &  (~ ng22615) ) | ( ng1312  &  ng22615  &  (~ ng23377) ) ;
 assign ng28360 = ( ng1306  &  (~ ng1315) ) | ( ng1315  &  ng27157 ) ;
 assign ng26272 = ( wire34390 ) | ( ng1312  &  (~ ng1192)  &  ng21435 ) ;
 assign ng27678 = ( (~ ng1365)  &  (~ ng1312)  &  ng23979 ) | ( (~ ng1365)  &  (~ ng1316)  &  ng23979 ) | ( ng1365  &  (~ ng1312)  &  (~ ng23979) ) | ( ng1365  &  (~ ng1316)  &  (~ ng23979) ) ;
 assign ng20912 = ( ng1391  &  ng13134 ) | ( (~ ng1339)  &  (~ ng13134) ) ;
 assign ng21016 = ( ng1404  &  ng13126 ) | ( (~ ng1352)  &  (~ ng13126) ) ;
 assign ng20898 = ( ng1413  &  ng13126 ) | ( (~ ng1378)  &  (~ ng13126) ) ;
 assign ng22263 = ( ng1423  &  (~ ng1315) ) | ( ng1423  &  (~ ng1316) ) | ( (~ ng1316)  &  (~ ng11726) ) ;
 assign ng22057 = ( ng1523  &  (~ ng853) ) | ( ng1523  &  (~ ng2257) ) | ( ng853  &  (~ ng1481)  &  ng2257 ) ;
 assign ng22114 = ( ng1539  &  (~ ng826) ) | ( ng1539  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng1506) ) ;
 assign ng25217 = ( ng1551  &  (~ ng13110) ) | ( ng1551  &  (~ ng826) ) | ( ng13110  &  ng826  &  wire3921 ) ;
 assign ng30295 = ( ng1585  &  (~ ng826) ) | ( ng826  &  wire6791 ) | ( ng826  &  wire34395 ) ;
 assign ng27612 = ( (~ ng1448)  &  (~ ng17031)  &  ng23528 ) | ( ng1448  &  (~ ng17031)  &  (~ ng23528) ) ;
 assign ng27275 = ( ng1750  &  (~ ng826) ) | ( ng1750  &  wire3309 ) | ( ng826  &  (~ ng21996)  &  (~ wire3309) ) ;
 assign ng29212 = ( ng1801  &  (~ ng823) ) | ( ng823  &  ng11952  &  ng27567 ) | ( ng823  &  (~ ng11952)  &  (~ ng27567) ) ;
 assign ng26821 = ( ng1822  &  (~ ng823) ) | ( ng823  &  wire3159 ) ;
 assign ng30338 = ( ng1701  &  (~ ng853) ) | ( ng853  &  wire7829 ) | ( ng853  &  wire7830 ) ;
 assign ng11564 = ( (~ ng1501) ) ;
 assign ng12524 = ( wire7763 ) | ( wire7764 ) | ( wire33184 ) | ( wire33186 ) ;
 assign ng24219 = ( ng1859  &  (~ ng823) ) | ( ng823  &  ng11666  &  wire32944 ) ;
 assign ng27320 = ( ng1960  &  (~ ng1312) ) | ( ng1960  &  (~ ng22651) ) | ( ng1312  &  ng22651  &  (~ ng22093) ) ;
 assign ng24524 = ( wire6771 ) | ( ng1970  &  (~ ng1312) ) ;
 assign ng26559 = ( ng1871  &  (~ ng1309) ) | ( ng1309  &  ng12324  &  wire3442 ) ;
 assign ng13444 = ( (~ ng1660) ) ;
 assign ng24434 = ( ng2026  &  (~ ng10238)  &  (~ wire33413) ) | ( ng2026  &  (~ ng10238)  &  (~ wire33414) ) | ( (~ ng2026)  &  (~ ng10238)  &  wire33413  &  wire33414 ) ;
 assign ng20934 = ( ng2078  &  ng11730 ) | ( (~ ng2020)  &  (~ ng11730) ) ;
 assign ng21001 = ( ng2094  &  ng13142 ) | ( (~ ng2052)  &  (~ ng13142) ) ;
 assign ng21056 = ( ng2103  &  ng13142 ) | ( (~ ng2066)  &  (~ ng13142) ) ;
 assign ng22184 = ( ng2235  &  ng13165 ) | ( (~ ng13165)  &  wire33428 ) | ( (~ ng13165)  &  wire33429 ) ;
 assign ng25251 = ( ng2247  &  (~ ng13110) ) | ( ng2247  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng2170) ) ;
 assign ng30690 = ( ng2270  &  (~ ng826) ) | ( ng826  &  wire34402 ) | ( ng826  &  wire34403 ) ;
 assign ng30274 = ( ng2324  &  (~ ng826) ) | ( ng826  &  ng29681 ) ;
 assign ng30691 = ( ng2345  &  (~ ng823) ) | ( ng823  &  wire33823 ) | ( ng823  &  wire33824 ) ;
 assign ng29112 = ( (~ ng26897)  &  wire34412 ) | ( (~ ng28637)  &  (~ ng26897)  &  wire34410 ) ;
 assign ng27309 = ( ng2459  &  (~ ng826) ) | ( ng2459  &  wire3313 ) | ( ng826  &  (~ ng23353)  &  (~ wire3313) ) ;
 assign ng29213 = ( ng2492  &  (~ ng826) ) | ( ng826  &  ng12005  &  ng27577 ) | ( ng826  &  (~ ng12005)  &  (~ ng27577) ) ;
 assign ng30341 = ( ng2394  &  (~ ng823) ) | ( ng823  &  ng29920 ) ;
 assign ng11576 = ( (~ ng2165) ) ;
 assign ng21847 = ( wire3142 ) | ( ng2628  &  (~ ng1315) ) ;
 assign ng23418 = ( ng2533  &  (~ ng823) ) | ( ng823  &  (~ ng11678)  &  wire33862 ) ;
 assign ng27325 = ( ng2651  &  (~ ng1312) ) | ( ng2651  &  (~ ng22687) ) | ( ng1312  &  ng22687  &  (~ ng23381) ) ;
 assign ng23348 = ( wire6702 ) | ( (~ ng21974)  &  wire34452 ) ;
 assign ng21043 = ( ng2784  &  ng11733 ) | ( (~ ng2734)  &  (~ ng11733) ) ;
 assign ng21081 = ( ng2793  &  ng11733 ) | ( (~ ng2753)  &  (~ ng11733) ) ;
 assign ng25272 = ( ng2809  &  ng13146 ) | ( (~ ng13146)  &  wire34617 ) | ( (~ ng13146)  &  wire34618 ) ;
 assign ng29453 = ( wire6572 ) | ( wire34074 ) | ( wire34075 ) | ( wire34620 ) ;
 assign ng25452 = ( ng3099  &  (~ ng1315) ) | ( ng1315  &  ng21851 ) ;
 assign ng17247 = ( ng3158  &  (~ ng1312) ) | ( ng1312  &  ng499 ) ;
 assign ng17383 = ( ng3179  &  (~ ng1315) ) | ( ng1315  &  ng1880 ) ;
 assign ng22125 = ( ng164  &  ng15950 ) | ( (~ ng15950)  &  wire31201 ) | ( (~ ng15950)  &  wire31202 ) ;
 assign ng25220 = ( ng178  &  (~ ng13110) ) | ( ng178  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng12876) ) ;
 assign ng30268 = ( ng264  &  (~ ng853) ) | ( ng853  &  ng29671 ) ;
 assign ng27594 = ( (~ ng74)  &  (~ ng17031)  &  ng23497 ) | ( ng74  &  (~ ng17031)  &  (~ ng23497) ) ;
 assign ng27255 = ( ng343  &  (~ ng823) ) | ( ng343  &  wire3290 ) | ( ng823  &  (~ wire3290)  &  (~ ng23320) ) ;
 assign ng28732 = ( ng408  &  (~ ng826) ) | ( ng826  &  ng27528 ) ;
 assign ng27759 = ( ng448  &  wire3595 ) | ( (~ wire3595)  &  (~ wire34663)  &  (~ wire34664) ) ;
 assign ng11509 = ( (~ ng125) ) ;
 assign ng12487 = ( wire31550 ) | ( wire31551 ) ;
 assign ng23385 = ( ng455  &  (~ ng826) ) | ( ng826  &  (~ ng11624)  &  wire31336 ) ;
 assign ng13149 = ( wire6519 ) | ( wire6520 ) | ( wire34675 ) | ( wire34677 ) ;
 assign ng27280 = ( ng580  &  (~ ng1312) ) | ( ng580  &  (~ ng22578) ) | ( ng1312  &  ng22578  &  (~ ng22050) ) ;
 assign ng27327 = ( ng584  &  (~ ng1315) ) | ( ng584  &  (~ ng22578) ) | ( ng1315  &  ng22578  &  (~ ng22083) ) ;
 assign ng28344 = ( wire6508 ) | ( ng608  &  (~ ng1312) ) ;
 assign ng26660 = ( (~ ng660)  &  ng672  &  ng10677 ) | ( ng660  &  ng672  &  ng10677  &  wire3319 ) | ( ng660  &  (~ ng672)  &  ng10677  &  (~ wire3319) ) ;
 assign ng20893 = ( ng705  &  ng13123 ) | ( (~ ng653)  &  (~ ng13123) ) ;
 assign ng20945 = ( ng712  &  ng13113 ) | ( (~ ng660)  &  (~ ng13113) ) ;
 assign ng21011 = ( ng723  &  ng13123 ) | ( (~ ng686)  &  (~ ng13123) ) ;
 assign ng22218 = ( ng738  &  (~ ng1309) ) | ( ng738  &  (~ ng630) ) | ( (~ ng630)  &  (~ ng13123) ) ;
 assign ng22177 = ( ng820  &  (~ ng853) ) | ( ng820  &  (~ ng2257) ) | ( ng853  &  (~ ng789)  &  ng2257 ) ;
 assign ng22042 = ( ng836  &  (~ ng826) ) | ( ng836  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng801) ) ;
 assign ng22127 = ( ng844  &  (~ ng853) ) | ( ng844  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng813) ) ;
 assign ng30681 = ( ng885  &  (~ ng823) ) | ( ng823  &  wire34273 ) | ( ng823  &  wire34274 ) ;
 assign ng30247 = ( ng900  &  (~ ng826) ) | ( ng826  &  wire6488 ) | ( ng826  &  wire34686 ) ;
 assign ng30642 = ( ng912  &  (~ ng823) ) | ( ng823  &  wire34689 ) | ( ng823  &  wire34690 ) ;
 assign ng28635 = ( ng753  &  (~ ng758)  &  (~ ng17031) ) | ( ng753  &  ng758  &  (~ ng17031)  &  wire3303 ) | ( (~ ng753)  &  ng758  &  (~ ng17031)  &  (~ wire3303) ) ;
 assign ng27313 = ( ng1078  &  (~ ng853) ) | ( ng1078  &  wire3293 ) | ( ng853  &  (~ wire3293)  &  (~ ng22005) ) ;
 assign ng26809 = ( wire6452 ) | ( ng1119  &  (~ ng823) ) ;
 assign ng27765 = ( ng1134  &  wire3530 ) | ( (~ wire3530)  &  (~ wire34737)  &  (~ wire34738) ) ;
 assign ng29173 = ( wire34743 ) | ( ng823  &  (~ ng27850)  &  wire34293 ) ;
 assign ng23126 = ( ng1175  &  (~ ng853) ) | ( ng853  &  (~ wire32262)  &  (~ wire32263) ) ;
 assign ng24222 = ( ng1155  &  (~ ng823) ) | ( ng823  &  ng11647  &  wire31828 ) ;
 assign ng26534 = ( wire30883 ) | ( (~ ng1186)  &  ng1309  &  ng21851 ) ;
 assign ng27301 = ( ng1268  &  (~ ng1309) ) | ( ng1268  &  (~ ng22615) ) | ( ng1309  &  ng22615  &  (~ ng23377) ) ;
 assign ng28346 = ( ng1291  &  (~ ng1309) ) | ( ng1309  &  wire6424 ) | ( ng1309  &  wire34748 ) ;
 assign ng13427 = ( (~ ng1140) ) ;
 assign ng21033 = ( ng1402  &  ng11726 ) | ( (~ ng1352)  &  (~ ng11726) ) ;
 assign ng20975 = ( ng1416  &  ng10706 ) | ( (~ ng10706)  &  wire32272 ) | ( (~ ng10706)  &  wire32273 ) ;
 assign ng25270 = ( ng1420  &  ng11726 ) | ( (~ ng11726)  &  wire34912 ) | ( (~ ng11726)  &  wire34913 ) ;
 assign ng22043 = ( ng1525  &  (~ ng823) ) | ( ng1525  &  (~ ng2257) ) | ( ng823  &  (~ ng1481)  &  ng2257 ) ;
 assign ng22131 = ( ng1540  &  (~ ng823) ) | ( ng1540  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng1506) ) ;
 assign ng25225 = ( ng1554  &  (~ ng13110) ) | ( ng1554  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng1476) ) ;
 assign ng30294 = ( ng1573  &  (~ ng853) ) | ( ng853  &  wire6292 ) | ( ng853  &  wire34916 ) ;
 assign ng28147 = ( (~ ng1448)  &  ng1444  &  (~ ng17031) ) | ( ng1444  &  (~ ng17031)  &  (~ ng23528) ) | ( ng1448  &  (~ ng1444)  &  (~ ng17031)  &  ng23528 ) ;
 assign ng27289 = ( ng1765  &  (~ ng826) ) | ( ng1765  &  wire3309 ) | ( ng826  &  (~ ng23349)  &  (~ wire3309) ) ;
 assign ng28760 = ( ng1792  &  (~ ng823) ) | ( ng823  &  ng27566 ) ;
 assign ng26816 = ( ng1819  &  (~ ng826) ) | ( ng826  &  wire3159 ) ;
 assign ng29178 = ( wire34934 ) | ( ng826  &  (~ ng27875)  &  wire34932 ) ;
 assign ng23413 = ( ng1839  &  (~ ng823) ) | ( ng823  &  (~ ng11666)  &  wire32979 ) ;
 assign ng12482 = ( wire3049 ) | ( wire7724 ) | ( wire33248 ) | ( wire33252 ) ;
 assign ng27331 = ( (~ ng1315)  &  ng1958 ) | ( ng1958  &  (~ ng22651) ) | ( ng1315  &  ng22651  &  (~ ng22093) ) ;
 assign ng24535 = ( wire6255 ) | ( (~ ng1312)  &  ng1979 ) ;
 assign ng26573 = ( (~ ng1312)  &  ng1874 ) | ( ng1312  &  ng12324  &  wire3442 ) ;
 assign ng13447 = ( (~ ng1666) ) ;
 assign ng20752 = ( (~ ng1312)  &  ng2020  &  wire3259 ) | ( ng2020  &  (~ ng2010)  &  wire3259 ) | ( (~ ng1312)  &  (~ ng2020)  &  (~ wire3259) ) | ( (~ ng2020)  &  (~ ng2010)  &  (~ wire3259) ) ;
 assign ng20915 = ( ng2080  &  ng13137 ) | ( (~ ng2020)  &  (~ ng13137) ) ;
 assign ng21023 = ( ng2113  &  (~ ng10238) ) | ( ng10238  &  wire33167 ) | ( ng10238  &  wire33168 ) ;
 assign ng22183 = ( ng2209  &  (~ ng826) ) | ( ng2209  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2170) ) ;
 assign ng22173 = ( ng2239  &  ng15970 ) | ( (~ ng15970)  &  wire33630 ) | ( (~ ng15970)  &  wire33631 ) ;
 assign ng25256 = ( ng2250  &  (~ ng13110) ) | ( ng2250  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng2165) ) ;
 assign ng30660 = ( ng2306  &  (~ ng826) ) | ( ng826  &  wire33799 ) | ( ng826  &  wire33800 ) ;
 assign ng30304 = ( ng2285  &  (~ ng853) ) | ( ng853  &  wire6240 ) | ( ng853  &  wire34937 ) ;
 assign ng30694 = ( ng2348  &  (~ ng853) ) | ( ng853  &  wire33823 ) | ( ng853  &  wire33824 ) ;
 assign ng13110 = ( wire31297  &  wire31298  &  wire31774  &  wire31775 ) ;
 assign ng27292 = ( ng2444  &  (~ ng826) ) | ( ng2444  &  wire3313 ) | ( ng826  &  (~ wire3313)  &  (~ ng22009) ) ;
 assign ng28782 = ( ng2489  &  (~ ng853) ) | ( ng853  &  ng27576 ) ;
 assign ng30356 = ( ng2395  &  (~ ng853) ) | ( ng853  &  ng29920 ) ;
 assign ng11592 = ( (~ ng2190) ) ;
 assign ng12539 = ( wire34948 ) | ( wire34949 ) ;
 assign ng23407 = ( ng2530  &  (~ ng826) ) | ( ng826  &  (~ ng11678)  &  wire33862 ) ;
 assign ng13175 = ( wire6212 ) | ( wire6213 ) | ( wire34956 ) | ( wire34958 ) ;
 assign ng27337 = ( (~ ng1312)  &  ng2654 ) | ( ng2654  &  (~ ng22687) ) | ( ng1312  &  ng22687  &  (~ ng22118) ) ;
 assign ng24438 = ( ng2720  &  ng10747  &  (~ wire34449) ) | ( ng2720  &  ng10747  &  (~ wire34450) ) | ( (~ ng2720)  &  ng10747  &  wire34449  &  wire34450 ) ;
 assign ng20963 = ( ng2777  &  ng13145 ) | ( (~ ng2707)  &  (~ ng13145) ) ;
 assign ng21074 = ( ng2795  &  ng13145 ) | ( (~ ng2753)  &  (~ ng13145) ) ;
 assign ng25280 = ( ng2810  &  ng13145 ) | ( (~ ng13145)  &  wire34617 ) | ( (~ ng13145)  &  wire34618 ) ;
 assign ng29456 = ( wire6190 ) | ( wire34074 ) | ( wire34075 ) | ( wire34963 ) ;
 assign ng28420 = ( wire6188 ) | ( ng3100  &  (~ ng1309) ) ;
 assign ng17229 = ( ng3155  &  (~ ng1309) ) | ( ng1309  &  ng499 ) ;
 assign ng17271 = ( ng3182  &  (~ ng1309) ) | ( ng1309  &  ng2574 ) ;
 assign ng22143 = ( ng162  &  ng13165 ) | ( (~ ng13165)  &  wire31201 ) | ( (~ ng13165)  &  wire31202 ) ;
 assign ng25228 = ( (~ ng13110)  &  ng174 ) | ( ng174  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng97) ) ;
 assign ng30635 = ( ng222  &  (~ ng826) ) | ( ng826  &  wire34982 ) | ( ng826  &  wire34983 ) ;
 assign ng27120 = ( wire6155 ) | ( (~ ng26529)  &  wire34985 ) ;
 assign ng27258 = ( ng346  &  (~ ng853) ) | ( ng346  &  wire3290 ) | ( ng853  &  (~ wire3290)  &  (~ ng23320) ) ;
 assign ng27293 = ( ng391  &  (~ ng853) ) | ( ng391  &  wire3290 ) | ( ng853  &  (~ ng21991)  &  (~ wire3290) ) ;
 assign ng30468 = ( ng319  &  (~ ng823) ) | ( ng823  &  ng29912 ) ;
 assign ng11493 = ( (~ ng105) ) ;
 assign ng18726 = ( ng557  &  ng1315 ) | ( (~ ng1315)  &  ng510 ) ;
 assign ng23117 = ( ng488  &  (~ ng853) ) | ( ng853  &  (~ wire31394)  &  (~ wire31395) ) ;
 assign ng27269 = ( ng579  &  (~ ng1309) ) | ( ng579  &  (~ ng22578) ) | ( ng1309  &  ng22578  &  (~ ng22050) ) ;
 assign ng24491 = ( wire6140 ) | ( ng587  &  (~ ng1309) ) ;
 assign ng28342 = ( wire6138 ) | ( ng605  &  (~ ng1309) ) ;
 assign ng26776 = ( (~ ng23950)  &  wire34992 ) | ( (~ ng26660)  &  (~ ng23950)  &  wire34990 ) ;
 assign ng20901 = ( ng701  &  ng11721 ) | ( (~ ng633)  &  (~ ng11721) ) ;
 assign ng20966 = ( ng710  &  ng11721 ) | ( (~ ng660)  &  (~ ng11721) ) ;
 assign ng21031 = ( ng719  &  ng11721 ) | ( (~ ng679)  &  (~ ng11721) ) ;
 assign ng22231 = ( (~ ng1312)  &  ng739 ) | ( ng739  &  (~ ng630) ) | ( (~ ng630)  &  (~ ng13113) ) ;
 assign ng22163 = ( ng822  &  (~ ng823) ) | ( ng822  &  (~ ng2257) ) | ( ng823  &  (~ ng789)  &  ng2257 ) ;
 assign ng22055 = ( ng837  &  (~ ng823) ) | ( ng837  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng801) ) ;
 assign ng22105 = ( ng846  &  (~ ng823) ) | ( ng846  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng813) ) ;
 assign ng30687 = ( ng888  &  (~ ng853) ) | ( ng853  &  wire34273 ) | ( ng853  &  wire34274 ) ;
 assign ng30270 = ( ng942  &  (~ ng853) ) | ( ng853  &  ng29672 ) ;
 assign ng30647 = ( ng915  &  (~ ng853) ) | ( ng853  &  wire34689 ) | ( ng853  &  wire34690 ) ;
 assign ng28146 = ( ng758  &  (~ ng762)  &  (~ ng17031) ) | ( ng758  &  (~ ng17031)  &  (~ ng23513) ) | ( (~ ng758)  &  ng762  &  (~ ng17031)  &  ng23513 ) ;
 assign ng28738 = ( ng1095  &  (~ ng826) ) | ( ng826  &  ng27550 ) ;
 assign ng26806 = ( wire6107 ) | ( ng1116  &  (~ ng826) ) ;
 assign ng29609 = ( wire6105 ) | ( ng999  &  (~ ng826) ) ;
 assign ng29170 = ( wire34997 ) | ( ng826  &  (~ ng27850)  &  wire34293 ) ;
 assign ng23392 = ( ng1142  &  (~ ng826) ) | ( ng826  &  (~ ng11647)  &  wire32200 ) ;
 assign ng24212 = ( ng1152  &  (~ ng826) ) | ( ng826  &  ng11647  &  wire31828 ) ;
 assign ng13124 = ( wire3049 ) | ( wire6089 ) | ( wire35003 ) | ( wire35007 ) ;
 assign ng27314 = ( (~ ng1315)  &  ng1264 ) | ( ng1264  &  (~ ng22615) ) | ( ng1315  &  ng22615  &  (~ ng22069) ) ;
 assign ng13426 = ( (~ ng1138) ) ;
 assign ng13428 = ( (~ ng966) ) ;
 assign ng21017 = ( ng1406  &  ng13134 ) | ( (~ ng1365)  &  (~ ng13134) ) ;
 assign ng20952 = ( ng1415  &  wire3204 ) | ( (~ wire3204)  &  wire32272 ) | ( (~ wire3204)  &  wire32273 ) ;
 assign ng22234 = ( (~ ng1309)  &  ng1424 ) | ( ng1424  &  (~ ng1316) ) | ( (~ ng1316)  &  (~ ng13134) ) ;
 assign ng22035 = ( ng1524  &  (~ ng826) ) | ( ng1524  &  (~ ng2257) ) | ( ng826  &  (~ ng1481)  &  ng2257 ) ;
 assign ng22150 = ( ng1538  &  (~ ng853) ) | ( ng1538  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng1506) ) ;
 assign ng25233 = ( (~ ng13110)  &  ng1550 ) | ( ng1550  &  (~ ng853) ) | ( ng13110  &  ng853  &  wire3921 ) ;
 assign ng25234 = ( (~ ng13110)  &  ng1555 ) | ( ng1555  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng1476) ) ;
 assign ng28636 = ( (~ ng1444)  &  ng1439  &  (~ ng17031) ) | ( ng1444  &  ng1439  &  (~ ng17031)  &  wire3325 ) | ( ng1444  &  (~ ng1439)  &  (~ ng17031)  &  (~ wire3325) ) ;
 assign ng27302 = ( ng1742  &  (~ ng853) ) | ( ng1742  &  wire3309 ) | ( ng853  &  (~ ng21996)  &  (~ wire3309) ) ;
 assign ng28771 = ( ng1795  &  (~ ng853) ) | ( ng853  &  ng27566 ) ;
 assign ng26820 = ( wire6057 ) | ( ng1816  &  (~ ng853) ) ;
 assign ng29181 = ( wire35014 ) | ( ng823  &  (~ ng27875)  &  wire34932 ) ;
 assign ng11565 = ( (~ ng1496) ) ;
 assign ng24182 = ( ng1842  &  (~ ng853) ) | ( ng853  &  (~ ng11666)  &  wire32979 ) ;
 assign ng24243 = ( ng1852  &  (~ ng853) ) | ( ng853  &  ng11666  &  wire32703 ) ;
 assign ng27321 = ( (~ ng1309)  &  ng1962 ) | ( ng1962  &  (~ ng22651) ) | ( ng1309  &  ng22651  &  (~ ng23388) ) ;
 assign ng24525 = ( wire6043 ) | ( (~ ng1309)  &  ng1976 ) ;
 assign ng26592 = ( (~ ng1315)  &  ng1877 ) | ( ng1315  &  ng12324  &  wire3442 ) ;
 assign ng13446 = ( (~ ng1664) ) ;
 assign ng21972 = ( (~ ng2020)  &  ng2013  &  (~ ng10238) ) | ( ng2020  &  ng2013  &  (~ ng10238)  &  wire3259 ) | ( ng2020  &  (~ ng2013)  &  (~ ng10238)  &  (~ wire3259) ) ;
 assign ng20899 = ( ng2079  &  ng13142 ) | ( (~ ng2020)  &  (~ ng13142) ) ;
 assign ng21042 = ( ng2111  &  wire3201 ) | ( (~ wire3201)  &  wire33167 ) | ( (~ wire3201)  &  wire33168 ) ;
 assign ng22192 = ( ng2205  &  (~ ng853) ) | ( ng2205  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2165) ) ;
 assign ng22185 = ( ng2240  &  ng15950 ) | ( (~ ng15950)  &  wire33630 ) | ( (~ ng15950)  &  wire33631 ) ;
 assign ng25252 = ( (~ ng13110)  &  ng2252 ) | ( ng2252  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng2165) ) ;
 assign ng30666 = ( ng2309  &  (~ ng823) ) | ( ng823  &  wire33799 ) | ( ng823  &  wire33800 ) ;
 assign ng30303 = ( ng2282  &  (~ ng823) ) | ( ng823  &  wire6240 ) | ( ng823  &  wire34937 ) ;
 assign ng25067 = ( (~ ng2160)  &  ng17197 ) | ( ng2160  &  (~ ng853)  &  (~ ng17197) ) | ( ng2160  &  (~ ng2257)  &  (~ ng17197) ) ;
 assign ng29582 = ( ng2120  &  (~ ng17031)  &  wire3372 ) | ( (~ ng2120)  &  (~ ng17031)  &  (~ wire3372) ) ;
 assign ng27308 = ( ng2433  &  (~ ng823) ) | ( ng2433  &  wire3313 ) | ( ng823  &  (~ wire3313)  &  (~ ng22009) ) ;
 assign ng28773 = ( ng2486  &  (~ ng823) ) | ( ng823  &  ng27576 ) ;
 assign ng29182 = ( wire35020 ) | ( ng826  &  (~ ng27892)  &  wire35018 ) ;
 assign ng18820 = ( ng2631  &  ng1315 ) | ( (~ ng1315)  &  ng2584 ) ;
 assign ng21970 = ( ng2563  &  (~ ng853) ) | ( ng853  &  (~ wire33937)  &  (~ wire33938) ) ;
 assign ng27326 = ( (~ ng1309)  &  ng2653 ) | ( ng2653  &  (~ ng22687) ) | ( ng1309  &  ng22687  &  (~ ng22118) ) ;
 assign ng25197 = ( wire6005 ) | ( wire6006 ) ;
 assign ng20940 = ( ng2776  &  ng13146 ) | ( (~ ng2707)  &  (~ ng13146) ) ;
 assign ng21006 = ( ng2785  &  ng13146 ) | ( (~ ng2734)  &  (~ ng13146) ) ;
 assign ng25288 = ( ng2808  &  ng11733 ) | ( (~ ng11733)  &  wire34617 ) | ( (~ ng11733)  &  wire34618 ) ;
 assign ng29455 = ( wire3425 ) | ( wire5993 ) | ( wire5994 ) ;
 assign ng26037 = ( ng2900  &  (~ wire3139)  &  wire3395 ) | ( (~ ng2900)  &  (~ wire3139)  &  (~ wire3395) ) ;
 assign ng17246 = ( (~ ng1315)  &  ng3093 ) | ( ng1315  &  ng1939 ) ;
 assign ng29939 = ( (~ ng1312)  &  ng3104 ) | ( ng1312  &  wire9559 ) | ( ng1312  &  wire30886 ) ;
 assign ng17248 = ( (~ ng1309)  &  ng3173 ) | ( ng1309  &  ng1880 ) ;
 assign ng28313 = ( ng3123  &  (~ ng17973) ) | ( (~ ng17973)  &  ng8381 ) | ( (~ ng17973)  &  wire30893 ) ;
 assign ng30668 = ( ng195  &  (~ ng826) ) | ( ng826  &  wire35038 ) | ( ng826  &  wire35039 ) ;
 assign ng30262 = ( ng255  &  (~ ng853) ) | ( ng853  &  ng29670 ) ;
 assign ng30669 = ( ng270  &  (~ ng823) ) | ( ng823  &  ng30021 ) ;
 assign ng29579 = ( ng52  &  (~ ng17031)  &  wire3371 ) | ( (~ ng52)  &  (~ ng17031)  &  (~ wire3371) ) ;
 assign ng27278 = ( ng388  &  (~ ng823) ) | ( ng388  &  wire3290 ) | ( ng823  &  (~ ng21991)  &  (~ wire3290) ) ;
 assign ng26106 = ( wire35135 ) | ( wire35136 ) | ( wire35137 ) | ( wire35138 ) ;
 assign ng23093 = ( ng487  &  (~ ng823) ) | ( ng823  &  (~ wire31394)  &  (~ wire31395) ) ;
 assign ng13410 = ( (~ ng451) ) ;
 assign ng20314 = ( (~ ng1315)  &  ng659 ) | ( ng1315  &  wire31471  &  wire31472 ) ;
 assign ng21010 = ( ng721  &  ng13113 ) | ( (~ ng679)  &  (~ ng13113) ) ;
 assign ng22242 = ( (~ ng1315)  &  ng737 ) | ( ng737  &  (~ ng630) ) | ( (~ ng630)  &  (~ ng11721) ) ;
 assign ng25221 = ( (~ ng13110)  &  ng856 ) | ( ng856  &  (~ ng853) ) | ( ng13110  &  ng853  &  wire3909 ) ;
 assign ng30277 = ( wire5899 ) | ( ng876  &  (~ ng823) ) ;
 assign ng28746 = ( ng1098  &  (~ ng823) ) | ( ng823  &  ng27550 ) ;
 assign ng26810 = ( ng1125  &  (~ ng826) ) | ( ng826  &  wire3157 ) ;
 assign ng11538 = ( (~ ng805) ) ;
 assign ng23406 = ( ng1145  &  (~ ng823) ) | ( ng823  &  (~ ng11647)  &  wire32200 ) ;
 assign ng12467 = ( wire8405 ) | ( wire8406 ) | ( wire32332 ) | ( wire32334 ) ;
 assign ng27285 = ( (~ ng1312)  &  ng1263 ) | ( ng1263  &  (~ ng22615) ) | ( ng1312  &  ng22615  &  (~ ng23364) ) ;
 assign ng24511 = ( wire5879 ) | ( (~ ng1309)  &  ng1282 ) ;
 assign ng26569 = ( (~ ng1315)  &  ng1183 ) | ( ng1315  &  ng12288  &  wire3439 ) ;
 assign ng21034 = ( ng1407  &  ng13126 ) | ( (~ ng1365)  &  (~ ng13126) ) ;
 assign ng20976 = ( ng1418  &  wire3204 ) | ( (~ wire3204)  &  wire32292 ) | ( (~ wire3204)  &  wire32293 ) ;
 assign ng22178 = ( ng1511  &  (~ ng853) ) | ( ng1511  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng1471) ) ;
 assign ng22074 = ( ng1531  &  (~ ng823) ) | ( ng1531  &  (~ ng2257) ) | ( ng823  &  (~ ng1491)  &  ng2257 ) ;
 assign ng22091 = ( ng1534  &  (~ ng823) ) | ( ng1534  &  (~ ng2257) ) | ( ng823  &  (~ ng1496)  &  ng2257 ) ;
 assign ng22152 = ( ng1545  &  ng15970 ) | ( (~ ng15970)  &  wire32828 ) | ( (~ ng15970)  &  wire32829 ) ;
 assign ng29111 = ( (~ ng26887)  &  wire35159 ) | ( (~ ng28636)  &  (~ ng26887)  &  wire35157 ) ;
 assign ng27317 = ( ng1757  &  (~ ng853) ) | ( ng1757  &  wire3309 ) | ( ng853  &  (~ ng23349)  &  (~ wire3309) ) ;
 assign ng28772 = ( wire5858 ) | ( wire35161 ) ;
 assign ng29613 = ( wire5854 ) | ( ng1693  &  (~ ng826) ) ;
 assign ng30704 = ( ng1696  &  (~ ng826) ) | ( ng826  &  ng30032 ) ;
 assign ng26675 = ( ng1783  &  (~ ng853) ) | ( ng1783  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng24683) ) ;
 assign ng23030 = ( ng1865  &  (~ ng823) ) | ( ng823  &  wire33018 ) | ( ng823  &  wire33019 ) ;
 assign ng13135 = ( wire5836 ) | ( wire5837 ) | ( wire35184 ) | ( wire35186 ) ;
 assign ng27341 = ( (~ ng1312)  &  ng1966 ) | ( ng1966  &  (~ ng22651) ) | ( ng1312  &  ng22651  &  (~ ng22134) ) ;
 assign ng13449 = ( (~ ng1670) ) ;
 assign ng20978 = ( ng2089  &  ng13137 ) | ( (~ ng2026)  &  (~ ng13137) ) ;
 assign ng21041 = ( ng2100  &  ng13142 ) | ( (~ ng2059)  &  (~ ng13142) ) ;
 assign ng21022 = ( ng2108  &  wire3201 ) | ( (~ wire3201)  &  wire33147 ) | ( (~ wire3201)  &  wire33148 ) ;
 assign ng22182 = ( ng2207  &  (~ ng823) ) | ( ng2207  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2165) ) ;
 assign ng22194 = ( ng2238  &  ng13165 ) | ( (~ ng13165)  &  wire33630 ) | ( (~ ng13165)  &  wire33631 ) ;
 assign ng25257 = ( (~ ng13110)  &  ng2255 ) | ( ng2255  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng12974) ) ;
 assign ng30667 = ( ng2315  &  (~ ng826) ) | ( ng826  &  wire35190 ) | ( ng826  &  wire35191 ) ;
 assign ng30260 = ( ng2294  &  (~ ng853) ) | ( ng853  &  wire5810 ) | ( ng853  &  wire35193 ) ;
 assign ng30297 = ( ng2339  &  (~ ng853) ) | ( ng853  &  ng29684 ) ;
 assign ng27621 = ( (~ ng2142)  &  (~ ng17031)  &  ng23539 ) | ( ng2142  &  (~ ng17031)  &  (~ ng23539) ) ;
 assign ng27291 = ( ng2418  &  (~ ng823) ) | ( ng2418  &  wire3313 ) | ( ng823  &  (~ wire3313)  &  (~ ng23344) ) ;
 assign ng28763 = ( ng2483  &  (~ ng826) ) | ( ng826  &  ng27576 ) ;
 assign ng29185 = ( wire35211 ) | ( ng823  &  (~ ng27892)  &  wire35018 ) ;
 assign ng11572 = ( (~ ng2185) ) ;
 assign ng23133 = ( ng2562  &  (~ ng823) ) | ( ng823  &  (~ wire33937)  &  (~ wire33938) ) ;
 assign ng24538 = ( wire5749 ) | ( (~ ng1309)  &  ng2670 ) ;
 assign ng26616 = ( (~ ng1315)  &  ng2571 ) | ( ng1315  &  ng12352  &  wire3435 ) ;
 assign ng13464 = ( (~ ng2362) ) ;
 assign ng22269 = ( (~ ng1309)  &  ng2812 ) | ( ng2812  &  (~ ng2704) ) | ( (~ ng2704)  &  (~ ng13146) ) ;
 assign ng29458 = ( wire5739 ) | ( wire35278 ) ;
 assign ng17226 = ( (~ ng1309)  &  ng3094 ) | ( ng1309  &  ng2633 ) ;
 assign ng29936 = ( (~ ng1309)  &  ng3103 ) | ( ng1309  &  wire9559 ) | ( ng1309  &  wire30886 ) ;
 assign ng17303 = ( ng1312  &  ng1880 ) | ( (~ ng1312)  &  ng3176 ) ;
 assign ng30674 = ( ng198  &  (~ ng823) ) | ( ng823  &  wire35038 ) | ( ng823  &  wire35039 ) ;
 assign ng30257 = ( ng252  &  (~ ng823) ) | ( ng823  &  ng29670 ) ;
 assign ng30245 = ( ng213  &  (~ ng826) ) | ( ng826  &  wire5726 ) | ( ng826  &  wire35280 ) ;
 assign ng27253 = ( ng354  &  (~ ng826) ) | ( ng354  &  wire3290 ) | ( ng826  &  (~ wire3290)  &  (~ ng23320) ) ;
 assign ng27267 = ( ng398  &  (~ ng826) ) | ( ng398  &  wire3290 ) | ( ng826  &  (~ ng21991)  &  (~ wire3290) ) ;
 assign ng23067 = ( ng486  &  (~ ng826) ) | ( ng826  &  (~ wire31394)  &  (~ wire31395) ) ;
 assign ng13411 = ( (~ ng453) ) ;
 assign ng16654 = ( ng1315  &  ng510 ) | ( (~ ng1315)  &  ng630 ) ;
 assign ng20923 = ( ng711  &  ng13123 ) | ( (~ ng660)  &  (~ ng13123) ) ;
 assign ng22029 = ( ng830  &  (~ ng826) ) | ( ng830  &  (~ ng2257) ) | ( ng826  &  (~ ng793)  &  ng2257 ) ;
 assign ng25215 = ( (~ ng13110)  &  ng860 ) | ( ng860  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng789) ) ;
 assign ng30269 = ( wire5707 ) | ( ng873  &  (~ ng826) ) ;
 assign ng28758 = ( ng1101  &  (~ ng853) ) | ( ng853  &  ng27550 ) ;
 assign ng26813 = ( wire5702 ) | ( ng1122  &  (~ ng853) ) ;
 assign ng11522 = ( (~ ng785) ) ;
 assign ng24179 = ( ng1148  &  (~ ng853) ) | ( ng853  &  (~ ng11647)  &  wire32200 ) ;
 assign ng24235 = ( ng1158  &  (~ ng853) ) | ( ng853  &  ng11647  &  wire31828 ) ;
 assign ng27339 = ( (~ ng1315)  &  ng1270 ) | ( ng1270  &  (~ ng22615) ) | ( ng1315  &  ng22615  &  (~ ng22108) ) ;
 assign ng24522 = ( wire5694 ) | ( (~ ng1312)  &  ng1285 ) ;
 assign ng26557 = ( (~ ng1312)  &  ng1180 ) | ( ng1312  &  ng12288  &  wire3439 ) ;
 assign ng21052 = ( ng1405  &  ng11726 ) | ( (~ ng1365)  &  (~ ng11726) ) ;
 assign ng20996 = ( ng1414  &  wire3200 ) | ( (~ wire3200)  &  wire32272 ) | ( (~ wire3200)  &  wire32273 ) ;
 assign ng22167 = ( ng1515  &  (~ ng826) ) | ( ng1515  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng1476) ) ;
 assign ng22059 = ( ng1530  &  (~ ng826) ) | ( ng1530  &  (~ ng2257) ) | ( ng826  &  (~ ng1491)  &  ng2257 ) ;
 assign ng22112 = ( ng1532  &  (~ ng853) ) | ( ng1532  &  (~ ng2257) ) | ( ng853  &  (~ ng1496)  &  ng2257 ) ;
 assign ng22168 = ( ng1541  &  ng13165 ) | ( (~ ng13165)  &  wire32816 ) | ( (~ ng13165)  &  wire32817 ) ;
 assign ng29355 = ( (~ ng1430)  &  (~ ng17031)  &  ng26887 ) | ( ng1430  &  (~ ng17031)  &  (~ ng26887) ) ;
 assign ng27303 = ( ng1754  &  (~ ng823) ) | ( ng1754  &  wire3309 ) | ( ng823  &  (~ ng23349)  &  (~ wire3309) ) ;
 assign ng28778 = ( wire5673 ) | ( wire35284 ) ;
 assign ng27768 = ( ng1828  &  (~ ng853) ) | ( ng853  &  (~ ng24004)  &  wire35288 ) | ( ng1828  &  (~ ng24004)  &  (~ wire35288) ) ;
 assign ng30706 = ( ng1697  &  (~ ng823) ) | ( ng823  &  ng30032 ) ;
 assign ng26670 = ( ng1785  &  (~ ng823) ) | ( ng1785  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng24683) ) ;
 assign ng23058 = ( ng1845  &  (~ ng853) ) | ( ng853  &  wire33018 ) | ( ng853  &  wire33019 ) ;
 assign ng29113 = ( wire9559 ) | ( wire30886 ) ;
 assign ng27290 = ( (~ ng1309)  &  ng1956 ) | ( ng1956  &  (~ ng22651) ) | ( ng1309  &  ng22651  &  (~ ng23372) ) ;
 assign ng27333 = ( (~ ng1309)  &  ng1965 ) | ( ng1965  &  (~ ng22651) ) | ( ng1309  &  ng22651  &  (~ ng22134) ) ;
 assign ng22651 = ( wire7769 ) | ( wire7770 ) | ( (~ ng12324)  &  wire3442 ) ;
 assign ng13448 = ( (~ ng1668) ) ;
 assign ng20999 = ( ng2087  &  ng11730 ) | ( (~ ng2026)  &  (~ ng11730) ) ;
 assign ng21054 = ( ng2096  &  ng11730 ) | ( (~ ng2046)  &  (~ ng11730) ) ;
 assign ng21003 = ( ng2112  &  wire3199 ) | ( (~ wire3199)  &  wire33167 ) | ( (~ wire3199)  &  wire33168 ) ;
 assign ng22170 = ( ng2206  &  (~ ng826) ) | ( ng2206  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2165) ) ;
 assign ng25227 = ( (~ ng13110)  &  ng2245 ) | ( ng2245  &  (~ ng826) ) | ( ng13110  &  ng826  &  wire3908 ) ;
 assign ng25253 = ( (~ ng13110)  &  ng2254 ) | ( ng2254  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng12974) ) ;
 assign ng30673 = ( ng2318  &  (~ ng823) ) | ( ng823  &  wire35190 ) | ( ng823  &  wire35191 ) ;
 assign ng30256 = ( ng2291  &  (~ ng823) ) | ( ng823  &  wire5810 ) | ( ng823  &  wire35193 ) ;
 assign ng30652 = ( ng2297  &  (~ ng826) ) | ( ng826  &  wire35294 ) | ( ng826  &  wire35295 ) ;
 assign ng27131 = ( wire5626 ) | ( (~ ng26532)  &  wire35304 ) ;
 assign ng27307 = ( ng2421  &  (~ ng853) ) | ( ng2421  &  wire3313 ) | ( ng853  &  (~ wire3313)  &  (~ ng23344) ) ;
 assign ng27342 = ( ng2466  &  (~ ng853) ) | ( ng2466  &  wire3313 ) | ( ng853  &  (~ wire3313)  &  (~ ng22021) ) ;
 assign ng29187 = ( wire35308 ) | ( ng853  &  (~ ng27892)  &  wire35018 ) ;
 assign ng19048 = ( (~ wire3046)  &  (~ wire7246)  &  (~ wire33868)  &  (~ wire33872) ) ;
 assign ng23114 = ( ng2561  &  (~ ng826) ) | ( ng826  &  (~ wire33937)  &  (~ wire33938) ) ;
 assign ng27343 = ( (~ ng1315)  &  ng2652 ) | ( ng2652  &  (~ ng22687) ) | ( ng1315  &  ng22687  &  (~ ng22118) ) ;
 assign ng13463 = ( (~ ng2360) ) ;
 assign ng22284 = ( (~ ng1312)  &  ng2813 ) | ( ng2813  &  (~ ng2704) ) | ( (~ ng1312)  &  (~ ng13145) ) | ( (~ ng2704)  &  (~ ng13145) ) ;
 assign ng29457 = ( wire5605 ) | ( wire35310 ) ;
 assign ng17235 = ( (~ ng1312)  &  ng3095 ) | ( ng1312  &  ng2633 ) ;
 assign ng30796 = ( (~ ng1309)  &  ng3106 ) | ( ng1309  &  ng30072 ) ;
 assign ng17270 = ( ng1186  &  ng1312 ) | ( (~ ng1312)  &  ng3167 ) ;
 assign ng28696 = ( (~ wire6564)  &  (~ wire34622) ) ;
 assign ng30246 = ( ng216  &  (~ ng823) ) | ( ng823  &  wire5726 ) | ( ng823  &  wire35280 ) ;
 assign ng25027 = ( (~ ng92)  &  ng17197 ) | ( ng92  &  (~ ng853)  &  (~ ng17197) ) | ( ng92  &  (~ ng2257)  &  (~ ng17197) ) ;
 assign ng27277 = ( ng376  &  (~ ng853) ) | ( ng376  &  wire3290 ) | ( ng853  &  (~ wire3290)  &  (~ ng23331) ) ;
 assign ng13412 = ( (~ ng279) ) ;
 assign ng23136 = ( ng633  &  (~ ng640)  &  ng10677 ) | ( ng633  &  ng640  &  ng10677  &  wire3252 ) | ( (~ ng633)  &  ng640  &  ng10677  &  (~ wire3252) ) ;
 assign ng20891 = ( ng698  &  ng11721 ) | ( (~ ng640)  &  (~ ng11721) ) ;
 assign ng22067 = ( ng840  &  (~ ng823) ) | ( ng840  &  (~ ng2257) ) | ( ng823  &  (~ ng805)  &  ng2257 ) ;
 assign ng25222 = ( (~ ng13110)  &  ng861 ) | ( ng861  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng789) ) ;
 assign ng30643 = ( ng918  &  (~ ng826) ) | ( ng826  &  wire32135 ) | ( ng826  &  wire32136 ) ;
 assign ng30701 = ( ng1002  &  (~ ng826) ) | ( ng826  &  ng30031 ) ;
 assign ng26669 = ( wire5564 ) | ( ng1089  &  (~ ng853) ) | ( ng1089  &  (~ ng2257) ) ;
 assign ng11518 = ( (~ ng801) ) ;
 assign ng24181 = ( ng1164  &  (~ ng826) ) | ( ng826  &  ng11647  &  wire32128 ) ;
 assign ng27329 = ( (~ ng1312)  &  ng1272 ) | ( ng1272  &  (~ ng22615) ) | ( ng1312  &  ng22615  &  (~ ng22108) ) ;
 assign ng24532 = ( wire5557 ) | ( (~ ng1315)  &  ng1288 ) ;
 assign ng22615 = ( wire8439 ) | ( wire8440 ) | ( (~ ng12288)  &  wire3439 ) ;
 assign ng21035 = ( ng1409  &  ng13134 ) | ( (~ ng1372)  &  (~ ng13134) ) ;
 assign ng21018 = ( ng1417  &  wire3200 ) | ( (~ wire3200)  &  wire32292 ) | ( (~ wire3200)  &  wire32293 ) ;
 assign ng22149 = ( ng1512  &  (~ ng826) ) | ( ng1512  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng1471) ) ;
 assign ng22073 = ( ng1526  &  (~ ng853) ) | ( ng1526  &  (~ ng2257) ) | ( ng853  &  (~ ng1486)  &  ng2257 ) ;
 assign ng22092 = ( ng1536  &  (~ ng826) ) | ( ng1536  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng1501) ) ;
 assign ng22180 = ( ng1544  &  ng13165 ) | ( (~ ng13165)  &  wire32828 ) | ( (~ ng13165)  &  wire32829 ) ;
 assign ng29581 = ( ng1426  &  (~ ng17031)  &  wire3400 ) | ( (~ ng1426)  &  (~ ng17031)  &  (~ wire3400) ) ;
 assign ng27318 = ( ng1769  &  (~ ng823) ) | ( ng1769  &  wire3309 ) | ( ng823  &  (~ ng22016)  &  (~ wire3309) ) ;
 assign ng29218 = ( ng1804  &  (~ ng853) ) | ( ng853  &  ng11952  &  ng27567 ) | ( ng853  &  (~ ng11952)  &  (~ ng27567) ) ;
 assign ng27766 = ( ng1830  &  (~ ng823) ) | ( ng823  &  (~ ng24004)  &  wire35288 ) | ( ng1830  &  (~ ng24004)  &  (~ wire35288) ) ;
 assign ng30708 = ( ng1698  &  (~ ng853) ) | ( ng853  &  ng30032 ) ;
 assign ng23124 = ( ng1868  &  (~ ng823) ) | ( ng823  &  (~ wire33063)  &  (~ wire33064) ) ;
 assign ng24231 = ( ng1860  &  (~ ng853) ) | ( ng853  &  ng11666  &  wire32944 ) ;
 assign ng27305 = ( (~ ng1312)  &  ng1957 ) | ( (~ ng22651)  &  ng1957 ) | ( ng1312  &  ng22651  &  (~ ng23372) ) ;
 assign ng24513 = ( wire5527 ) | ( (~ ng1309)  &  ng1967 ) ;
 assign ng25194 = ( wire5525 ) | ( wire5526 ) ;
 assign ng20953 = ( ng2081  &  ng11730 ) | ( (~ ng2013)  &  (~ ng11730) ) ;
 assign ng20979 = ( ng2091  &  ng13142 ) | ( (~ ng2040)  &  (~ ng13142) ) ;
 assign ng21071 = ( ng2099  &  ng11730 ) | ( (~ ng2059)  &  (~ ng11730) ) ;
 assign ng20980 = ( ng2109  &  wire3199 ) | ( (~ wire3199)  &  wire33147 ) | ( (~ wire3199)  &  wire33148 ) ;
 assign ng22280 = ( (~ ng1315)  &  ng2117 ) | ( ng2117  &  (~ ng2010) ) | ( (~ ng2010)  &  (~ ng11730) ) ;
 assign ng25236 = ( (~ ng13110)  &  ng2246 ) | ( ng2246  &  (~ ng823) ) | ( ng13110  &  ng823  &  wire3908 ) ;
 assign ng30289 = ( ng2261  &  (~ ng826) ) | ( ng826  &  wire5512 ) | ( ng826  &  wire35341 ) ;
 assign ng30693 = ( ng2273  &  (~ ng823) ) | ( ng823  &  wire34402 ) | ( ng823  &  wire34403 ) ;
 assign ng30253 = ( ng2288  &  (~ ng826) ) | ( ng826  &  wire5810 ) | ( ng826  &  wire35193 ) ;
 assign ng30659 = ( ng2300  &  (~ ng823) ) | ( ng823  &  wire35294 ) | ( ng823  &  wire35295 ) ;
 assign ng28637 = ( ng2133  &  (~ ng2138)  &  (~ ng17031) ) | ( ng2133  &  ng2138  &  (~ ng17031)  &  wire3323 ) | ( (~ ng2133)  &  ng2138  &  (~ ng17031)  &  (~ wire3323) ) ;
 assign ng27335 = ( ng2463  &  (~ ng823) ) | ( ng2463  &  wire3313 ) | ( ng823  &  (~ wire3313)  &  (~ ng22021) ) ;
 assign ng26672 = ( ng2478  &  (~ ng826) ) | ( ng2478  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng24700) ) ;
 assign ng11573 = ( (~ ng2180) ) ;
 assign ng27338 = ( (~ ng1309)  &  ng2656 ) | ( ng2656  &  (~ ng22687) ) | ( ng1309  &  ng22687  &  (~ ng23395) ) ;
 assign ng24557 = ( wire5492 ) | ( (~ ng1315)  &  ng2676 ) ;
 assign ng13462 = ( (~ ng2358) ) ;
 assign ng22299 = ( (~ ng1315)  &  ng2811 ) | ( ng2811  &  (~ ng2704) ) | ( (~ ng2704)  &  (~ ng11733) ) ;
 assign ng17269 = ( (~ ng1315)  &  ng3096 ) | ( ng1315  &  ng2633 ) ;
 assign ng29941 = ( (~ ng1315)  &  ng3105 ) | ( ng1315  &  wire9559 ) | ( ng1315  &  wire30886 ) ;
 assign ng17340 = ( ng1186  &  ng1315 ) | ( (~ ng1315)  &  ng3170 ) ;
 assign ng30248 = ( ng219  &  (~ ng853) ) | ( ng853  &  wire5726 ) | ( ng853  &  wire35280 ) ;
 assign ng30675 = ( ng273  &  (~ ng853) ) | ( ng853  &  ng30021 ) ;
 assign ng29353 = ( (~ ng56)  &  (~ ng17031)  &  ng26869 ) | ( ng56  &  (~ ng17031)  &  (~ ng26869) ) ;
 assign ng13413 = ( (~ ng281) ) ;
 assign ng20682 = ( (~ ng1312)  &  ng640  &  wire3252 ) | ( (~ ng630)  &  ng640  &  wire3252 ) | ( (~ ng1312)  &  (~ ng640)  &  (~ wire3252) ) | ( (~ ng630)  &  (~ ng640)  &  (~ wire3252) ) ;
 assign ng23324 = ( wire5475 ) | ( (~ ng23136)  &  wire35345 ) ;
 assign ng22147 = ( ng847  &  ng13165 ) | ( (~ ng13165)  &  wire31770 ) | ( (~ ng13165)  &  wire31771 ) ;
 assign ng25230 = ( (~ ng13110)  &  ng859 ) | ( ng859  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng789) ) ;
 assign ng30285 = ( wire5469 ) | ( ng879  &  (~ ng853) ) ;
 assign ng30703 = ( ng1003  &  (~ ng823) ) | ( ng823  &  ng30031 ) ;
 assign ng26665 = ( wire5464 ) | ( ng1091  &  (~ ng823) ) | ( ng1091  &  (~ ng2257) ) ;
 assign ng27273 = ( (~ ng1309)  &  ng1262 ) | ( (~ ng22615)  &  ng1262 ) | ( ng1309  &  ng22615  &  (~ ng23364) ) ;
 assign ng27316 = ( (~ ng1309)  &  ng1271 ) | ( (~ ng22615)  &  ng1271 ) | ( ng1309  &  ng22615  &  (~ ng22108) ) ;
 assign ng28351 = ( (~ ng1309)  &  ng1300 ) | ( ng1309  &  ng27157 ) ;
 assign ng21053 = ( ng1410  &  ng13126 ) | ( (~ ng1372)  &  (~ ng13126) ) ;
 assign ng20997 = ( ng1419  &  ng10706 ) | ( (~ ng10706)  &  wire32292 ) | ( (~ ng10706)  &  wire32293 ) ;
 assign ng22166 = ( ng1513  &  (~ ng823) ) | ( ng1513  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng1471) ) ;
 assign ng22058 = ( ng1528  &  (~ ng823) ) | ( ng1528  &  (~ ng2257) ) | ( ng823  &  (~ ng1486)  &  ng2257 ) ;
 assign ng22113 = ( ng1537  &  (~ ng823) ) | ( ng1537  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng1501) ) ;
 assign ng22169 = ( ng1546  &  ng15950 ) | ( (~ ng15950)  &  wire32828 ) | ( (~ ng15950)  &  wire32829 ) ;
 assign ng27264 = ( ng1735  &  (~ ng826) ) | ( ng1735  &  wire3309 ) | ( ng826  &  (~ ng23335)  &  (~ wire3309) ) ;
 assign ng27304 = ( ng1779  &  (~ ng826) ) | ( ng1779  &  wire3309 ) | ( ng826  &  (~ ng22016)  &  (~ wire3309) ) ;
 assign ng28761 = ( wire5435 ) | ( wire35352 ) ;
 assign ng27764 = ( ng1829  &  (~ ng826) ) | ( ng826  &  (~ ng24004)  &  wire35288 ) | ( ng1829  &  (~ ng24004)  &  (~ wire35288) ) ;
 assign ng30487 = ( ng1699  &  (~ ng826) ) | ( ng826  &  wire7829 ) | ( ng826  &  wire7830 ) ;
 assign ng11563 = ( (~ ng1506) ) ;
 assign ng23097 = ( ng1867  &  (~ ng826) ) | ( ng826  &  (~ wire33063)  &  (~ wire33064) ) ;
 assign ng23123 = ( ng1861  &  (~ ng826) ) | ( ng826  &  wire33018 ) | ( ng826  &  wire33019 ) ;
 assign ng13164 = ( wire3049 ) | ( wire5419 ) | ( wire35358 ) | ( wire35362 ) ;
 assign ng27319 = ( (~ ng1315)  &  ng1955 ) | ( (~ ng22651)  &  ng1955 ) | ( ng1315  &  ng22651  &  (~ ng23372) ) ;
 assign ng27346 = ( (~ ng1315)  &  ng1964 ) | ( (~ ng22651)  &  ng1964 ) | ( ng1315  &  ng22651  &  (~ ng22134) ) ;
 assign ng26671 = ( (~ ng2040)  &  ng2052  &  (~ ng10238) ) | ( ng2040  &  ng2052  &  (~ ng10238)  &  wire3296 ) | ( ng2040  &  (~ ng2052)  &  (~ ng10238)  &  (~ wire3296) ) ;
 assign ng20935 = ( ng2083  &  ng13137 ) | ( (~ ng2013)  &  (~ ng13137) ) ;
 assign ng21000 = ( ng2092  &  ng13137 ) | ( (~ ng2040)  &  (~ ng13137) ) ;
 assign ng21055 = ( ng2101  &  ng13137 ) | ( (~ ng2059)  &  (~ ng13137) ) ;
 assign ng21002 = ( ng2110  &  (~ ng10238) ) | ( ng10238  &  wire33147 ) | ( ng10238  &  wire33148 ) ;
 assign ng22267 = ( (~ ng1312)  &  ng2119 ) | ( ng2119  &  (~ ng2010) ) | ( (~ ng2010)  &  (~ ng13137) ) ;
 assign ng25245 = ( (~ ng13110)  &  ng2244 ) | ( ng2244  &  (~ ng853) ) | ( ng13110  &  ng853  &  wire3908 ) ;
 assign ng25259 = ( (~ ng13110)  &  ng2253 ) | ( ng2253  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng12974) ) ;
 assign ng30695 = ( ng2276  &  (~ ng853) ) | ( ng853  &  wire34402 ) | ( ng853  &  wire34403 ) ;
 assign ng30290 = ( ng2330  &  (~ ng853) ) | ( ng853  &  ng29681 ) ;
 assign ng30665 = ( ng2303  &  (~ ng853) ) | ( ng853  &  wire35294 ) | ( ng853  &  wire35295 ) ;
 assign ng28148 = ( (~ ng2142)  &  ng2138  &  (~ ng17031) ) | ( ng2138  &  (~ ng17031)  &  (~ ng23539) ) | ( ng2142  &  (~ ng2138)  &  (~ ng17031)  &  ng23539 ) ;
 assign ng27276 = ( ng2429  &  (~ ng826) ) | ( ng2429  &  wire3313 ) | ( ng826  &  (~ wire3313)  &  (~ ng23344) ) ;
 assign ng27324 = ( ng2473  &  (~ ng826) ) | ( ng2473  &  wire3313 ) | ( ng826  &  (~ wire3313)  &  (~ ng22021) ) ;
 assign ng26676 = ( ng2479  &  (~ ng823) ) | ( ng2479  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng24700) ) ;
 assign ng27344 = ( (~ ng1312)  &  ng2657 ) | ( ng2657  &  (~ ng22687) ) | ( ng1312  &  ng22687  &  (~ ng23395) ) ;
 assign ng24548 = ( wire5382 ) | ( (~ ng1312)  &  ng2673 ) ;
 assign ng26596 = ( (~ ng1312)  &  ng2568 ) | ( ng1312  &  ng12352  &  wire3435 ) ;
 assign ng29459 = ( wire5370 ) | ( wire5371 ) | ( wire35369 ) ;
 assign ng22026 = ( ng2888  &  (~ ng2950)  &  (~ wire3139) ) | ( (~ ng2888)  &  ng2950  &  ng2883  &  (~ wire3139) ) | ( ng2888  &  ng2950  &  (~ ng2883)  &  (~ wire3139) ) ;
 assign ng22100 = ( ng130  &  (~ ng826) ) | ( ng130  &  (~ ng2257) ) | ( ng826  &  (~ ng97)  &  ng2257 ) ;
 assign ng22037 = ( ng144  &  (~ ng853) ) | ( ng144  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng109) ) ;
 assign ng22080 = ( ng158  &  (~ ng823) ) | ( ng158  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng125) ) ;
 assign ng25207 = ( (~ ng13110)  &  ng172 ) | ( ng172  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng101) ) ;
 assign ng30275 = ( ng192  &  (~ ng853) ) | ( ng853  &  wire5356 ) | ( ng853  &  wire35375 ) ;
 assign ng30284 = ( ng207  &  (~ ng823) ) | ( ng823  &  wire5351 ) | ( ng823  &  wire35378 ) ;
 assign ng27760 = ( ng449  &  wire3570 ) | ( (~ wire3570)  &  (~ wire34663)  &  (~ wire34664) ) ;
 assign ng29167 = ( wire35381 ) | ( (~ ng15970)  &  ng17051  &  (~ ng27834) ) ;
 assign ng27294 = ( (~ ng1315)  &  ng578 ) | ( ng578  &  (~ ng22578) ) | ( ng1315  &  ng22578  &  (~ ng22050) ) ;
 assign ng24508 = ( wire5335 ) | ( (~ ng1312)  &  ng599 ) ;
 assign ng13417 = ( (~ ng289) ) ;
 assign ng20879 = ( ng700  &  ng13113 ) | ( (~ ng640)  &  (~ ng13113) ) ;
 assign ng22087 = ( ng838  &  (~ ng853) ) | ( ng838  &  (~ ng2257) ) | ( ng853  &  (~ ng805)  &  ng2257 ) ;
 assign ng22148 = ( ng852  &  ng15950 ) | ( (~ ng15950)  &  wire32020 ) | ( (~ ng15950)  &  wire32021 ) ;
 assign ng25232 = ( (~ ng13110)  &  ng866 ) | ( ng866  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng12916) ) ;
 assign ng30293 = ( ng894  &  (~ ng823) ) | ( ng823  &  wire5326 ) | ( ng823  &  wire35384 ) ;
 assign ng30638 = ( ng909  &  (~ ng826) ) | ( ng826  &  wire34689 ) | ( ng826  &  wire34690 ) ;
 assign ng11536 = ( (~ ng813) ) ;
 assign ng28350 = ( (~ ng1312)  &  ng1294 ) | ( ng1312  &  wire6424 ) | ( ng1312  &  wire34748 ) ;
 assign ng13433 = ( (~ ng976) ) ;
 assign ng24430 = ( ng1332  &  ng10706  &  (~ wire32566) ) | ( ng1332  &  ng10706  &  (~ wire32567) ) | ( (~ ng1332)  &  ng10706  &  wire32566  &  wire32567 ) ;
 assign ng20911 = ( ng1389  &  ng13126 ) | ( (~ ng1319)  &  (~ ng13126) ) ;
 assign ng20974 = ( ng1400  &  ng13134 ) | ( (~ ng1358)  &  (~ ng13134) ) ;
 assign ng25244 = ( (~ ng13110)  &  ng1560 ) | ( ng1560  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng12945) ) ;
 assign ng30692 = ( ng1582  &  (~ ng853) ) | ( ng853  &  wire35390 ) | ( ng853  &  wire35391 ) ;
 assign ng30252 = ( ng1597  &  (~ ng823) ) | ( ng823  &  wire5303 ) | ( ng823  &  wire35394 ) ;
 assign ng25056 = ( (~ ng1466)  &  ng17197 ) | ( ng1466  &  (~ ng853)  &  (~ ng17197) ) | ( ng1466  &  (~ ng2257)  &  (~ ng17197) ) ;
 assign ng22076 = ( ng2217  &  (~ ng853) ) | ( ng2217  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2175) ) ;
 assign ng22139 = ( ng2231  &  (~ ng823) ) | ( ng2231  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2195) ) ;
 assign ng25237 = ( (~ ng13110)  &  ng2248 ) | ( ng2248  &  (~ ng826) ) | ( ng13110  &  ng826  &  (~ ng2170) ) ;
 assign ng28783 = ( wire5288 ) | ( wire35396 ) ;
 assign ng29618 = ( ng2387  &  (~ ng826) ) | ( ng826  &  wire5286 ) | ( ng826  &  wire5287 ) ;
 assign ng26025 = ( ng2477  &  (~ ng853) ) | ( ng2477  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng24700) ) ;
 assign ng11574 = ( (~ ng2175) ) ;
 assign ng27347 = ( (~ ng1315)  &  ng2655 ) | ( ng2655  &  (~ ng22687) ) | ( ng1315  &  ng22687  &  (~ ng23395) ) ;
 assign ng28368 = ( (~ ng1312)  &  ng2691 ) | ( ng1312  &  wire5200 ) | ( ng1312  &  wire35555 ) ;
 assign ng16718 = ( ng1315  &  ng2584 ) | ( (~ ng1315)  &  ng2704 ) ;
 assign ng28328 = ( ng2766  &  (~ ng2760)  &  ng10747 ) | ( ng2766  &  ng2760  &  ng10747  &  wire3370 ) | ( (~ ng2766)  &  ng2760  &  ng10747  &  (~ wire3370) ) ;
 assign ng21005 = ( ng2783  &  ng13145 ) | ( (~ ng2720)  &  (~ ng13145) ) ;
 assign ng21062 = ( ng2794  &  ng13146 ) | ( (~ ng2753)  &  (~ ng13146) ) ;
 assign ng29460 = ( wire5176 ) | ( wire5177 ) | ( wire35566 ) ;
 assign ng30908 = ( wire3833 ) | ( wire5049 ) | ( (~ ng29728)  &  wire3229 ) ;
 assign ng30982 = ( wire5013 ) | ( wire5021 ) | ( wire35751 ) | ( wire35753 ) ;
 assign ng25191 = ( ng3013  &  ng21796  &  wire3333 ) | ( ng3013  &  ng21796  &  (~ wire35755) ) | ( (~ ng3013)  &  ng21796  &  (~ wire3333)  &  wire35755 ) ;
 assign ng16844 = ( ng3063  &  ng2987 ) | ( ng3044  &  (~ ng2987) ) ;
 assign ng16854 = ( ng3072  &  ng2987 ) | ( ng3053  &  (~ ng2987) ) ;
 assign ng23358 = ( (~ ng2888)  &  ng2896  &  (~ wire3139) ) | ( (~ ng2888)  &  ng2896  &  (~ wire3310) ) | ( ng2888  &  (~ ng2896)  &  (~ wire3310) ) | ( ng2888  &  ng2896  &  (~ wire3139)  &  wire3310 ) ;
 assign ng22122 = ( ng131  &  (~ ng823) ) | ( ng131  &  (~ ng2257) ) | ( ng823  &  (~ ng97)  &  ng2257 ) ;
 assign ng22031 = ( ng146  &  (~ ng823) ) | ( ng146  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng109) ) ;
 assign ng22101 = ( ng156  &  (~ ng853) ) | ( ng156  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng125) ) ;
 assign ng25211 = ( (~ ng13110)  &  ng168 ) | ( ng168  &  (~ ng853) ) | ( ng13110  &  ng853  &  wire3942 ) ;
 assign ng30637 = ( ng231  &  (~ ng826) ) | ( ng826  &  wire35768 ) | ( ng826  &  wire35769 ) ;
 assign ng30276 = ( ng204  &  (~ ng826) ) | ( ng826  &  wire5351 ) | ( ng826  &  wire35378 ) ;
 assign ng28736 = ( wire4985 ) | ( wire35770 ) ;
 assign ng29169 = ( wire35772 ) | ( (~ ng15950)  &  ng17051  &  (~ ng27834) ) ;
 assign ng11511 = ( (~ ng117) ) ;
 assign ng27281 = ( (~ ng1309)  &  ng582 ) | ( ng582  &  (~ ng22578) ) | ( ng1309  &  ng22578  &  (~ ng23368) ) ;
 assign ng24499 = ( wire4975 ) | ( (~ ng1309)  &  ng596 ) ;
 assign ng22578 = ( wire9082 ) | ( wire9083 ) | ( (~ ng12245)  &  wire3444 ) ;
 assign ng13416 = ( (~ ng287) ) ;
 assign ng20944 = ( ng707  &  ng11721 ) | ( (~ ng646)  &  (~ ng11721) ) ;
 assign ng22033 = ( ng831  &  (~ ng823) ) | ( ng831  &  (~ ng2257) ) | ( ng823  &  (~ ng793)  &  ng2257 ) ;
 assign ng22164 = ( ng850  &  ng13165 ) | ( (~ ng13165)  &  wire32020 ) | ( (~ ng13165)  &  wire32021 ) ;
 assign ng25240 = ( (~ ng13110)  &  ng862 ) | ( ng862  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng785) ) ;
 assign ng30298 = ( ng897  &  (~ ng853) ) | ( ng853  &  wire5326 ) | ( ng853  &  wire35384 ) ;
 assign ng30278 = ( ng951  &  (~ ng853) ) | ( ng853  &  ng29677 ) ;
 assign ng11520 = ( (~ ng793) ) ;
 assign ng24501 = ( wire4955 ) | ( (~ ng1309)  &  ng1273 ) ;
 assign ng24072 = ( (~ pg3229)  &  ng992 ) | ( pg3229  &  (~ ng978) ) ;
 assign ng23329 = ( wire4947 ) | ( (~ ng21969)  &  wire35791 ) ;
 assign ng20925 = ( ng1387  &  ng11726 ) | ( (~ ng1319)  &  (~ ng11726) ) ;
 assign ng20993 = ( ng1396  &  ng11726 ) | ( (~ ng1346)  &  (~ ng11726) ) ;
 assign ng25250 = ( (~ ng13110)  &  ng1561 ) | ( ng1561  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng12945) ) ;
 assign ng30688 = ( ng1579  &  (~ ng823) ) | ( ng823  &  wire35390 ) | ( ng823  &  wire35391 ) ;
 assign ng30255 = ( ng1600  &  (~ ng853) ) | ( ng853  &  wire5303 ) | ( ng853  &  wire35394 ) ;
 assign ng30689 = ( wire4928 ) | ( ng1654  &  (~ ng853) ) ;
 assign ng11548 = ( (~ ng1476) ) ;
 assign ng22061 = ( ng2221  &  (~ ng826) ) | ( ng2221  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2180) ) ;
 assign ng22117 = ( ng2230  &  (~ ng826) ) | ( ng2230  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2195) ) ;
 assign ng30296 = ( ng2264  &  (~ ng823) ) | ( ng823  &  wire5512 ) | ( ng823  &  wire35341 ) ;
 assign ng28788 = ( wire4918 ) | ( wire35798 ) ;
 assign ng27771 = ( ng2522  &  (~ ng853) ) | ( ng853  &  (~ ng24038)  &  wire33948 ) | ( ng2522  &  (~ ng24038)  &  (~ wire33948) ) ;
 assign ng11590 = ( (~ ng2200) ) ;
 assign ng27345 = ( (~ ng1309)  &  ng2659 ) | ( ng2659  &  (~ ng22687) ) | ( ng1309  &  ng22687  &  (~ ng22157) ) ;
 assign ng28364 = ( (~ ng1309)  &  ng2688 ) | ( ng1309  &  wire5200 ) | ( ng1309  &  wire35555 ) ;
 assign ng13458 = ( (~ ng2526) ) ;
 assign ng13466 = ( (~ ng2366) ) ;
 assign ng20918 = ( ng2773  &  ng13146 ) | ( (~ ng2714)  &  (~ ng13146) ) ;
 assign ng20983 = ( ng2782  &  ng13146 ) | ( (~ ng2720)  &  (~ ng13146) ) ;
 assign ng21028 = ( ng2804  &  ng10747 ) | ( (~ ng10747)  &  wire33957 ) | ( (~ ng10747)  &  wire33958 ) ;
 assign ng29655 = ( wire35814 ) | ( ng510  &  (~ ng27382)  &  ng27379 ) | ( ng510  &  ng27382  &  (~ ng27379) ) ;
 assign ng30119 = ( wire35862 ) | ( ng1196  &  (~ ng28842)  &  ng28845 ) | ( ng1196  &  ng28842  &  (~ ng28845) ) ;
 assign ng30983 = ( wire3427 ) | ( wire4809 ) | ( wire4810 ) ;
 assign ng24445 = ( ng3002  &  (~ ng3006)  &  ng21796 ) | ( ng3002  &  ng21796  &  wire3333 ) | ( (~ ng3002)  &  ng3006  &  ng21796  &  (~ wire3333) ) ;
 assign ng16853 = ( ng3064  &  ng2987 ) | ( ng3045  &  (~ ng2987) ) ;
 assign ng16845 = ( ng3071  &  ng2987 ) | ( ng3052  &  (~ ng2987) ) ;
 assign ng24473 = ( (~ ng23358)  &  wire35872 ) | ( (~ wire3139)  &  wire35873 ) ;
 assign ng22141 = ( ng129  &  (~ ng853) ) | ( ng129  &  (~ ng2257) ) | ( ng853  &  (~ ng97)  &  ng2257 ) ;
 assign ng22038 = ( ng149  &  (~ ng823) ) | ( ng149  &  (~ ng2257) ) | ( ng823  &  (~ ng113)  &  ng2257 ) ;
 assign ng22079 = ( ng153  &  (~ ng853) ) | ( ng153  &  (~ ng2257) ) | ( ng853  &  (~ ng121)  &  ng2257 ) ;
 assign ng25206 = ( (~ ng13110)  &  ng170 ) | ( ng170  &  (~ ng823) ) | ( ng13110  &  ng823  &  wire3942 ) ;
 assign ng30640 = ( ng234  &  (~ ng823) ) | ( ng823  &  wire35768 ) | ( ng823  &  wire35769 ) ;
 assign ng30254 = ( ng249  &  (~ ng826) ) | ( ng826  &  ng29670 ) ;
 assign ng28745 = ( wire4784 ) | ( wire35874 ) ;
 assign ng29606 = ( wire4780 ) | ( ng312  &  (~ ng826) ) ;
 assign ng19012 = ( (~ wire9183)  &  (~ wire9184)  &  (~ wire31353)  &  (~ wire31355) ) ;
 assign ng23000 = ( ng484  &  (~ ng823) ) | ( ng823  &  wire31355 ) | ( ng823  &  wire31356 ) ;
 assign ng13111 = ( wire4775 ) | ( wire4776 ) | ( wire35884 ) | ( wire35886 ) ;
 assign ng21435 = ( pg16297  &  (~ ng506) ) | ( ng1312  &  (~ ng506) ) | ( ng506  &  ng507 ) ;
 assign ng13418 = ( (~ ng291) ) ;
 assign ng20991 = ( ng720  &  ng13123 ) | ( (~ ng679)  &  (~ ng13123) ) ;
 assign ng25209 = ( (~ ng13110)  &  ng857 ) | ( (~ ng826)  &  ng857 ) | ( ng13110  &  ng826  &  wire3909 ) ;
 assign ng25248 = ( (~ ng13110)  &  ng865 ) | ( ng865  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng12916) ) ;
 assign ng27123 = ( wire4757 ) | ( (~ ng26530)  &  (~ ng17031)  &  wire35895 ) ;
 assign ng27271 = ( ng1045  &  (~ ng823) ) | ( ng1045  &  wire3293 ) | ( ng823  &  (~ wire3293)  &  (~ ng21983) ) ;
 assign ng11537 = ( (~ ng809) ) ;
 assign ng18763 = ( (~ ng1315)  &  ng1196 ) | ( ng1315  &  ng1243 ) ;
 assign ng24510 = ( wire4748 ) | ( (~ ng1312)  &  ng1276 ) ;
 assign ng26547 = ( (~ ng1309)  &  ng1177 ) | ( ng1309  &  ng12288  &  wire3439 ) ;
 assign ng13434 = ( (~ ng978) ) ;
 assign ng26666 = ( ng1358  &  (~ ng1346)  &  ng10706 ) | ( ng1358  &  ng1346  &  wire3283  &  ng10706 ) | ( (~ ng1358)  &  ng1346  &  (~ wire3283)  &  ng10706 ) ;
 assign ng20910 = ( ng1384  &  ng11726 ) | ( (~ ng1326)  &  (~ ng11726) ) ;
 assign ng20973 = ( ng1398  &  ng13126 ) | ( (~ ng1346)  &  (~ ng13126) ) ;
 assign ng22090 = ( ng1529  &  (~ ng853) ) | ( ng1529  &  (~ ng2257) ) | ( ng853  &  (~ ng1491)  &  ng2257 ) ;
 assign ng22151 = ( ng1543  &  ng15950 ) | ( (~ ng15950)  &  wire32816 ) | ( (~ ng15950)  &  wire32817 ) ;
 assign ng25255 = ( (~ ng13110)  &  ng1559 ) | ( ng1559  &  (~ ng853) ) | ( ng13110  &  ng853  &  (~ ng12945) ) ;
 assign ng30664 = ( ng1624  &  (~ ng823) ) | ( ng823  &  wire35900 ) | ( ng823  &  wire35901 ) ;
 assign ng30280 = ( wire4722 ) | ( ng1636  &  (~ ng853) ) ;
 assign ng30684 = ( wire4721 ) | ( ng1651  &  (~ ng823) ) ;
 assign ng26667 = ( (~ ng826)  &  ng1784 ) | ( ng1784  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng24683) ) ;
 assign ng22077 = ( ng2222  &  (~ ng823) ) | ( ng2222  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2180) ) ;
 assign ng22140 = ( (~ ng826)  &  ng2233 ) | ( ng2233  &  (~ ng2257) ) | ( ng826  &  (~ ng2200)  &  ng2257 ) ;
 assign ng30679 = ( ng2321  &  (~ ng853) ) | ( ng853  &  wire35190 ) | ( ng853  &  wire35191 ) ;
 assign ng26817 = ( wire4708 ) | ( (~ ng826)  &  ng2504 ) ;
 assign ng29623 = ( ng2389  &  (~ ng853) ) | ( ng853  &  wire5286 ) | ( ng853  &  wire5287 ) ;
 assign ng11575 = ( (~ ng2170) ) ;
 assign ng30055 = ( wire35920 ) | ( wire4703  &  wire35918 ) | ( wire35917  &  wire35918 ) ;
 assign ng23047 = ( ng2559  &  (~ ng823) ) | ( ng823  &  wire33871 ) | ( ng823  &  wire33872 ) ;
 assign ng13143 = ( wire4695 ) | ( wire4696 ) | ( wire35927 ) | ( wire35929 ) ;
 assign ng27348 = ( (~ ng1312)  &  ng2660 ) | ( ng2660  &  (~ ng22687) ) | ( ng1312  &  ng22687  &  (~ ng22157) ) ;
 assign ng28358 = ( wire4683 ) | ( (~ ng1309)  &  ng2679 ) ;
 assign ng22687 = ( wire7152 ) | ( wire7153 ) | ( (~ ng12352)  &  wire3435 ) ;
 assign ng24092 = ( pg3229  &  (~ ng2366) ) | ( (~ pg3229)  &  ng2380 ) ;
 assign ng20939 = ( ng2774  &  ng13145 ) | ( (~ ng2714)  &  (~ ng13145) ) ;
 assign ng21061 = ( ng2792  &  ng13145 ) | ( (~ ng2740)  &  (~ ng13145) ) ;
 assign ng21007 = ( ng2803  &  wire3206 ) | ( (~ wire3206)  &  wire33957 ) | ( (~ wire3206)  &  wire33958 ) ;
 assign ng29972 = ( wire3835 ) | ( wire4662 ) | ( (~ ng27855)  &  wire3227 ) ;
 assign ng30910 = ( wire3834 ) | ( wire4654 ) | ( (~ ng29741)  &  wire3229 ) ;
 assign ng30980 = ( wire3427 ) | ( wire4647 ) | ( wire4648 ) ;
 assign ng23330 = ( wire4807 ) | ( wire4808 ) ;
 assign ng16860 = ( ng3065  &  ng2987 ) | ( ng3046  &  (~ ng2987) ) ;
 assign ng16880 = ( ng3074  &  ng2987 ) | ( ng3056  &  (~ ng2987) ) ;
 assign ng18542 = ( pg3231  &  (~ ng12999)  &  ng12988 ) | ( (~ ng3120)  &  (~ ng12999)  &  ng12988 ) | ( pg3231  &  ng12999  &  (~ ng12988) ) | ( (~ ng3120)  &  ng12999  &  (~ ng12988) ) | ( (~ pg3231)  &  ng3120  &  ng12999  &  ng12988 ) | ( (~ pg3231)  &  ng3120  &  (~ ng12999)  &  (~ ng12988) ) ;
 assign ng25201 = ( ng2903  &  (~ wire3139)  &  (~ wire35032) ) | ( ng2903  &  (~ wire3139)  &  (~ wire35033) ) | ( (~ ng2903)  &  (~ wire3139)  &  wire35032  &  wire35033 ) ;
 assign ng22123 = ( (~ ng826)  &  ng133 ) | ( ng133  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng101) ) ;
 assign ng22032 = ( (~ ng826)  &  ng148 ) | ( ng148  &  (~ ng2257) ) | ( ng826  &  (~ ng113)  &  ng2257 ) ;
 assign ng22065 = ( (~ ng826)  &  ng157 ) | ( ng157  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng125) ) ;
 assign ng25204 = ( (~ ng13110)  &  ng169 ) | ( (~ ng826)  &  ng169 ) | ( ng13110  &  ng826  &  wire3942 ) ;
 assign ng30645 = ( ng237  &  (~ ng853) ) | ( ng853  &  wire35768 ) | ( ng853  &  wire35769 ) ;
 assign ng30292 = ( ng210  &  (~ ng853) ) | ( ng853  &  wire5351 ) | ( ng853  &  wire35378 ) ;
 assign ng28754 = ( wire4610 ) | ( wire35961 ) ;
 assign ng27762 = ( ng447  &  wire3788 ) | ( (~ wire3788)  &  (~ wire34663)  &  (~ wire34664) ) ;
 assign ng30482 = ( ng320  &  (~ ng853) ) | ( ng853  &  ng29912 ) ;
 assign ng21346 = ( (~ ng298)  &  (~ ng299) ) | ( ng299  &  ng305  &  (~ ng823) ) ;
 assign ng23022 = ( ng464  &  (~ ng853) ) | ( ng853  &  wire31355 ) | ( ng853  &  wire31356 ) ;
 assign ng21851 = ( ng544  &  ng499 ) | ( (~ ng1309)  &  (~ ng499)  &  ng548 ) ;
 assign ng24059 = ( pg3229  &  (~ ng291) ) | ( (~ pg3229)  &  ng305 ) ;
 assign ng20947 = ( ng730  &  ng10677 ) | ( (~ ng10677)  &  wire31449 ) | ( (~ ng10677)  &  wire31450 ) ;
 assign ng20969 = ( ng728  &  wire3205 ) | ( (~ wire3205)  &  wire31449 ) | ( (~ wire3205)  &  wire31450 ) ;
 assign ng25214 = ( (~ ng13110)  &  ng858 ) | ( ng858  &  (~ ng823) ) | ( ng13110  &  ng823  &  wire3909 ) ;
 assign ng25241 = ( (~ ng13110)  &  ng867 ) | ( ng867  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng12916) ) ;
 assign ng27603 = ( (~ ng762)  &  (~ ng17031)  &  ng23513 ) | ( ng762  &  (~ ng17031)  &  (~ ng23513) ) ;
 assign ng27263 = ( ng1056  &  (~ ng826) ) | ( ng1056  &  wire3293 ) | ( ng826  &  (~ wire3293)  &  (~ ng21983) ) ;
 assign ng11521 = ( (~ ng789) ) ;
 assign ng12507 = ( wire3049 ) | ( wire8305 ) | ( wire32486 ) | ( wire32490 ) ;
 assign ng24521 = ( wire4588 ) | ( (~ ng1315)  &  ng1279 ) ;
 assign ng28354 = ( (~ ng1315)  &  ng1297 ) | ( ng1315  &  wire6424 ) | ( ng1315  &  wire34748 ) ;
 assign ng25189 = ( wire8274 ) | ( wire8275 ) ;
 assign ng20897 = ( ng1388  &  ng13134 ) | ( (~ ng1319)  &  (~ ng13134) ) ;
 assign ng20951 = ( ng1397  &  ng13134 ) | ( (~ ng1346)  &  (~ ng13134) ) ;
 assign ng22075 = ( (~ ng826)  &  ng1533 ) | ( ng1533  &  (~ ng2257) ) | ( ng826  &  (~ ng1496)  &  ng2257 ) ;
 assign ng22132 = ( ng1542  &  ng15970 ) | ( (~ ng15970)  &  wire32816 ) | ( (~ ng15970)  &  wire32817 ) ;
 assign ng30279 = ( (~ ng826)  &  ng1567 ) | ( ng826  &  wire6292 ) | ( ng826  &  wire34916 ) ;
 assign ng30658 = ( (~ ng826)  &  ng1621 ) | ( ng826  &  wire35900 ) | ( ng826  &  wire35901 ) ;
 assign ng30250 = ( (~ ng826)  &  ng1594 ) | ( ng826  &  wire5303 ) | ( ng826  &  wire35394 ) ;
 assign ng30678 = ( wire4571 ) | ( (~ ng826)  &  ng1648 ) ;
 assign ng29620 = ( wire4568 ) | ( ng1695  &  (~ ng853) ) ;
 assign ng11549 = ( (~ ng1471) ) ;
 assign ng22097 = ( ng2220  &  (~ ng853) ) | ( ng2220  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2180) ) ;
 assign ng22153 = ( ng2229  &  (~ ng853) ) | ( ng2229  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2195) ) ;
 assign ng30283 = ( (~ ng826)  &  ng2333 ) | ( ng826  &  ng29684 ) ;
 assign ng26822 = ( wire4560 ) | ( ng2507  &  (~ ng823) ) ;
 assign ng29621 = ( ng2388  &  (~ ng823) ) | ( ng823  &  wire5286 ) | ( ng823  &  wire5287 ) ;
 assign ng11591 = ( (~ ng2195) ) ;
 assign ng26144 = ( wire36039 ) | ( wire36040 ) | ( wire36041 ) | ( wire36042 ) ;
 assign ng23076 = ( ng2539  &  (~ ng853) ) | ( ng853  &  wire33871 ) | ( ng853  &  wire33872 ) ;
 assign ng30072 = ( wire30889 ) | ( wire9559  &  wire30887 ) | ( wire30886  &  wire30887 ) ;
 assign ng27354 = ( (~ ng1315)  &  ng2658 ) | ( (~ ng22687)  &  ng2658 ) | ( ng1315  &  ng22687  &  (~ ng22157) ) ;
 assign ng28371 = ( (~ ng1315)  &  ng2694 ) | ( ng1315  &  wire5200 ) | ( ng1315  &  wire35555 ) ;
 assign ng30061 = ( wire36050 ) | ( wire4506  &  wire36048 ) | ( wire36047  &  wire36048 ) ;
 assign ng13465 = ( (~ ng2364) ) ;
 assign ng21025 = ( ng2781  &  ng11733 ) | ( (~ ng2720)  &  (~ ng11733) ) ;
 assign ng21073 = ( ng2790  &  ng11733 ) | ( (~ ng2740)  &  (~ ng11733) ) ;
 assign ng20965 = ( ng2799  &  ng11733 ) | ( (~ ng2766)  &  (~ ng11733) ) ;
 assign ng29973 = ( wire3836 ) | ( wire4493 ) | ( wire3227  &  (~ ng27865) ) ;
 assign ng30909 = ( wire3834 ) | ( wire4487 ) | ( (~ ng29732)  &  wire3229 ) ;
 assign ng30981 = ( wire4479 ) | ( wire5021 ) | ( wire35751 ) | ( wire36055 ) ;
 assign ng26048 = ( (~ ng25265)  &  (~ ng21796) ) | ( (~ ng2998)  &  (~ ng25265)  &  ng2993 ) | ( ng2998  &  ng25265  &  ng21796 ) | ( ng2998  &  (~ ng2993)  &  ng21796 ) ;
 assign ng16803 = ( ng3066  &  ng2987 ) | ( ng3047  &  (~ ng2987) ) ;
 assign ng16861 = ( ng3073  &  ng2987 ) | ( ng3055  &  (~ ng2987) ) ;
 assign ng16802 = ( (~ pg51)  &  ng2950 ) ;
 assign ng28421 = ( wire4467 ) | ( (~ ng1312)  &  ng3101 ) ;
 assign ng17236 = ( ng1186  &  ng1309 ) | ( (~ ng1309)  &  ng3164 ) ;
 assign ng22142 = ( ng134  &  (~ ng823) ) | ( ng134  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng101) ) ;
 assign ng22039 = ( (~ ng826)  &  ng151 ) | ( ng151  &  (~ ng2257) ) | ( ng826  &  (~ ng117)  &  ng2257 ) ;
 assign ng22124 = ( ng159  &  ng13165 ) | ( (~ ng13165)  &  wire31159 ) | ( (~ ng13165)  &  wire31160 ) ;
 assign ng25219 = ( (~ ng13110)  &  ng176 ) | ( ng176  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng97) ) ;
 assign ng25229 = ( (~ ng13110)  &  ng179 ) | ( ng179  &  (~ ng823) ) | ( ng13110  &  ng823  &  (~ ng12876) ) ;
 assign ng30641 = ( (~ ng826)  &  ng240 ) | ( ng826  &  wire36064 ) | ( ng826  &  wire36065 ) ;
 assign ng30636 = ( ng225  &  (~ ng823) ) | ( ng823  &  wire34982 ) | ( ng823  &  wire34983 ) ;
 assign ng28634 = ( ng65  &  (~ ng70)  &  (~ ng17031) ) | ( ng65  &  ng70  &  (~ ng17031)  &  wire3324 ) | ( (~ ng65)  &  ng70  &  (~ ng17031)  &  (~ wire3324) ) ;
 assign ng27266 = ( ng373  &  (~ ng823) ) | ( ng373  &  wire3290 ) | ( ng823  &  (~ wire3290)  &  (~ ng23331) ) ;
 assign ng26803 = ( wire4436 ) | ( (~ ng826)  &  ng429 ) ;
 assign ng29611 = ( wire4434 ) | ( ng314  &  (~ ng853) ) ;
 assign ng26659 = ( wire4432 ) | ( ng404  &  (~ ng823) ) | ( ng404  &  (~ ng2257) ) ;
 assign ng23092 = ( (~ ng826)  &  ng480 ) | ( ng826  &  wire31355 ) | ( ng826  &  wire31356 ) ;
 assign ng24206 = ( ng465  &  (~ ng826) ) | ( ng826  &  ng11624  &  wire31067 ) ;
 assign ng13160 = ( wire3049 ) | ( wire4420 ) | ( wire36077 ) | ( wire36081 ) ;
 assign ng27296 = ( (~ ng1309)  &  ng585 ) | ( (~ ng22578)  &  ng585 ) | ( ng1309  &  ng22578  &  (~ ng22083) ) ;
 assign ng28353 = ( (~ ng1315)  &  ng620 ) | ( ng1315  &  wire4415 ) | ( ng1315  &  wire36086 ) ;
 assign ng27672 = ( (~ ng1312)  &  (~ ng679)  &  ng23950 ) | ( (~ ng630)  &  (~ ng679)  &  ng23950 ) | ( (~ ng1312)  &  ng679  &  (~ ng23950) ) | ( (~ ng630)  &  ng679  &  (~ ng23950) ) ;
 assign ng20921 = ( ng704  &  ng11721 ) | ( (~ ng653)  &  (~ ng11721) ) ;
 assign ng20990 = ( ng718  &  ng13113 ) | ( (~ ng666)  &  (~ ng13113) ) ;
 assign ng20924 = ( ng729  &  wire3210 ) | ( (~ wire3210)  &  wire31449 ) | ( (~ wire3210)  &  wire31450 ) ;
 assign ng20948 = ( ng732  &  wire3210 ) | ( (~ wire3210)  &  wire31469 ) | ( (~ wire3210)  &  wire31470 ) ;
 assign ng22041 = ( (~ ng823)  &  ng834 ) | ( ng834  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng797) ) ;
 assign ng22089 = ( (~ ng826)  &  ng845 ) | ( ng845  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng813) ) ;
 assign ng30649 = ( (~ ng826)  &  ng927 ) | ( ng826  &  ng30016 ) ;
 assign ng30251 = ( (~ ng853)  &  ng906 ) | ( ng853  &  wire6488 ) | ( ng853  &  wire34686 ) ;
 assign ng25935 = ( ng776  &  (~ ng780)  &  ng13165 ) | ( (~ ng776)  &  ng780  &  ng17197 ) | ( ng776  &  (~ ng780)  &  ng17197 ) | ( ng776  &  ng13165  &  (~ ng17197) ) ;
 assign ng27270 = ( (~ ng853)  &  ng1033 ) | ( ng1033  &  wire3293 ) | ( ng853  &  (~ wire3293)  &  (~ ng23325) ) ;
 assign ng27282 = ( ng1048  &  (~ ng853) ) | ( ng1048  &  wire3293 ) | ( ng853  &  (~ wire3293)  &  (~ ng21983) ) ;
 assign ng29204 = ( (~ ng823)  &  ng1107 ) | ( ng823  &  ng11902  &  ng27551 ) | ( ng823  &  (~ ng11902)  &  (~ ng27551) ) ;
 assign ng27761 = ( ng1135  &  wire3784 ) | ( (~ wire3784)  &  (~ wire34737)  &  (~ wire34738) ) ;
 assign ng30500 = ( (~ ng853)  &  ng1007 ) | ( ng853  &  wire4359 ) | ( ng853  &  wire4360 ) ;
 assign ng21843 = ( wire3142 ) | ( (~ ng1315)  &  ng1240 ) ;
 assign ng24213 = ( (~ ng823)  &  ng1165 ) | ( ng823  &  ng11647  &  wire32128 ) ;
 assign ng13155 = ( wire36131 ) | ( wire36132 ) ;
 assign ng27300 = ( (~ ng1312)  &  ng1266 ) | ( (~ ng22615)  &  ng1266 ) | ( ng1312  &  ng22615  &  (~ ng22069) ) ;
 assign ng13429 = ( (~ ng968) ) ;
 assign ng20333 = ( (~ ng1315)  &  ng1345 ) | ( ng1315  &  wire31471  &  wire31472 ) ;
 assign ng20882 = ( ng1385  &  ng13134 ) | ( (~ ng1326)  &  (~ ng13134) ) ;
 assign ng20972 = ( ng1393  &  ng11726 ) | ( (~ ng1332)  &  (~ ng11726) ) ;
 assign ng25263 = ( ng1421  &  ng13134 ) | ( (~ ng13134)  &  wire34912 ) | ( (~ ng13134)  &  wire34913 ) ;
 assign ng22191 = ( (~ ng853)  &  ng1514 ) | ( ng1514  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng1476) ) ;
 assign ng25242 = ( (~ ng13110)  &  ng1553 ) | ( (~ ng853)  &  ng1553 ) | ( ng13110  &  ng853  &  (~ ng1476) ) ;
 assign ng30657 = ( (~ ng823)  &  ng1615 ) | ( ng823  &  wire36135 ) | ( ng823  &  wire36136 ) ;
 assign ng30266 = ( wire4323 ) | ( (~ ng826)  &  ng1630 ) ;
 assign ng30656 = ( (~ ng853)  &  ng1609 ) | ( ng853  &  ng30015 ) ;
 assign ng26815 = ( wire4315 ) | ( (~ ng823)  &  ng1813 ) ;
 assign ng19036 = ( (~ wire33018)  &  (~ wire33019) ) ;
 assign ng22078 = ( (~ ng826)  &  ng2224 ) | ( ng2224  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2185) ) ;
 assign ng22171 = ( (~ ng853)  &  ng2232 ) | ( ng2232  &  (~ ng2257) ) | ( ng853  &  (~ ng2200)  &  ng2257 ) ;
 assign ng25940 = ( (~ ng2160)  &  ng2156  &  ng13165 ) | ( (~ ng2160)  &  ng2156  &  ng17197 ) | ( ng2160  &  (~ ng2156)  &  ng17197 ) | ( ng2156  &  ng13165  &  (~ ng17197) ) ;
 assign ng26825 = ( wire4309 ) | ( (~ ng853)  &  ng2510 ) ;
 assign ng30709 = ( (~ ng823)  &  ng2391 ) | ( ng823  &  ng30033 ) ;
 assign ng23132 = ( (~ ng826)  &  ng2555 ) | ( ng826  &  wire33871 ) | ( ng826  &  wire33872 ) ;
 assign ng24225 = ( ng2540  &  (~ ng826) ) | ( ng826  &  ng11678  &  wire33551 ) ;
 assign ng13194 = ( wire4291 ) | ( wire4292 ) | ( wire36160 ) | ( wire36162 ) ;
 assign ng24527 = ( wire4284 ) | ( (~ ng1309)  &  ng2661 ) ;
 assign ng28367 = ( wire4282 ) | ( (~ ng1315)  &  ng2685 ) ;
 assign ng13461 = ( (~ ng2356) ) ;
 assign ng26677 = ( (~ ng2734)  &  ng2746  &  ng10747 ) | ( ng2734  &  ng2746  &  ng10747  &  wire3304 ) | ( ng2734  &  (~ ng2746)  &  ng10747  &  (~ wire3304) ) ;
 assign ng20964 = ( ng2779  &  ng13146 ) | ( (~ ng2727)  &  (~ ng13146) ) ;
 assign ng21060 = ( ng2787  &  ng11733 ) | ( (~ ng2746)  &  (~ ng11733) ) ;
 assign ng20941 = ( ng2801  &  ng13145 ) | ( (~ ng2766)  &  (~ ng13145) ) ;
 assign ng20877 = ( (~ pg3234)  &  ng3080 ) ;
 assign ng29974 = ( wire3836 ) | ( wire4271 ) | ( (~ ng27883)  &  wire3227 ) ;
 assign ng30912 = ( wire36170 ) | ( ng1890  &  (~ ng1937)  &  (~ ng29751) ) ;
 assign ng30986 = ( wire4254 ) | ( wire4255 ) | ( wire36173 ) ;
 assign ng23359 = ( (~ ng3028)  &  (~ wire3292) ) | ( ng3028  &  ng21796  &  wire3292 ) | ( ng3028  &  wire3292  &  wire36176 ) ;
 assign ng16866 = ( ng3051  &  (~ ng2987) ) | ( ng2987  &  ng3070 ) ;
 assign ng18907 = ( ng3061  &  (~ ng2987) ) | ( ng2987  &  ng2997 ) ;
 assign ng16823 = ( (~ pg51)  &  ng2817 ) ;
 assign ng28425 = ( wire4239 ) | ( (~ ng1315)  &  ng3102 ) ;
 assign ng17302 = ( ng1315  &  ng499 ) | ( (~ ng1315)  &  ng3161 ) ;
 assign ng22161 = ( (~ ng853)  &  ng132 ) | ( ng132  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng101) ) ;
 assign ng22047 = ( (~ ng853)  &  ng147 ) | ( ng147  &  (~ ng2257) ) | ( ng853  &  (~ ng113)  &  ng2257 ) ;
 assign ng22103 = ( ng163  &  ng15970 ) | ( (~ ng15970)  &  wire31201 ) | ( (~ ng15970)  &  wire31202 ) ;
 assign ng25213 = ( (~ ng13110)  &  ng175 ) | ( (~ ng826)  &  ng175 ) | ( ng13110  &  ng826  &  (~ ng97) ) ;
 assign ng25239 = ( (~ ng13110)  &  ng177 ) | ( (~ ng853)  &  ng177 ) | ( ng13110  &  ng853  &  (~ ng12876) ) ;
 assign ng30680 = ( (~ ng853)  &  ng201 ) | ( ng853  &  wire35038 ) | ( ng853  &  wire35039 ) ;
 assign ng30639 = ( (~ ng853)  &  ng228 ) | ( ng853  &  wire34982 ) | ( ng853  &  wire34983 ) ;
 assign ng28145 = ( (~ ng74)  &  ng70  &  (~ ng17031) ) | ( ng70  &  (~ ng17031)  &  (~ ng23497) ) | ( ng74  &  (~ ng70)  &  (~ ng17031)  &  ng23497 ) ;
 assign ng29201 = ( (~ ng853)  &  ng423 ) | ( ng853  &  ng11860  &  ng27529 ) | ( ng853  &  (~ ng11860)  &  (~ ng27529) ) ;
 assign ng26804 = ( wire4217 ) | ( (~ ng823)  &  ng432 ) ;
 assign ng29608 = ( wire4215 ) | ( (~ ng823)  &  ng313 ) ;
 assign ng26664 = ( wire4214 ) | ( (~ ng853)  &  ng402 ) | ( ng402  &  (~ ng2257) ) ;
 assign ng11492 = ( (~ ng109) ) ;
 assign ng24216 = ( (~ ng853)  &  ng479 ) | ( ng853  &  ng11624  &  wire31271 ) ;
 assign ng24215 = ( (~ ng823)  &  ng468 ) | ( ng823  &  ng11624  &  wire31067 ) ;
 assign ng27312 = ( (~ ng1312)  &  ng586 ) | ( (~ ng22578)  &  ng586 ) | ( ng1312  &  ng22578  &  (~ ng22083) ) ;
 assign ng28349 = ( (~ ng1312)  &  ng617 ) | ( ng1312  &  wire4415 ) | ( ng1312  &  wire36086 ) ;
 assign ng28199 = ( (~ ng679)  &  ng686  &  ng10677 ) | ( ng686  &  ng10677  &  (~ ng23950) ) | ( ng679  &  (~ ng686)  &  ng10677  &  ng23950 ) ;
 assign ng20902 = ( ng706  &  ng13113 ) | ( (~ ng653)  &  (~ ng13113) ) ;
 assign ng21009 = ( ng716  &  ng11721 ) | ( (~ ng666)  &  (~ ng11721) ) ;
 assign ng20894 = ( ng725  &  ng11721 ) | ( (~ ng692)  &  (~ ng11721) ) ;
 assign ng20970 = ( ng733  &  ng10677 ) | ( (~ ng10677)  &  wire31469 ) | ( (~ ng10677)  &  wire31470 ) ;
 assign ng22054 = ( (~ ng853)  &  ng832 ) | ( ng832  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng797) ) ;
 assign ng22104 = ( (~ ng853)  &  ng841 ) | ( ng841  &  (~ ng2257) ) | ( ng853  &  (~ ng809)  &  ng2257 ) ;
 assign ng30655 = ( (~ ng823)  &  ng930 ) | ( ng823  &  ng30016 ) ;
 assign ng30249 = ( (~ ng823)  &  ng903 ) | ( ng823  &  wire6488 ) | ( ng823  &  wire34686 ) ;
 assign ng26530 = ( ng25935  &  ng771 ) | ( (~ ng776)  &  ng771  &  (~ ng17031) ) | ( (~ ng25935)  &  ng776  &  (~ ng771)  &  (~ ng17031) ) ;
 assign ng27262 = ( (~ ng823)  &  ng1030 ) | ( ng1030  &  wire3293 ) | ( ng823  &  (~ wire3293)  &  (~ ng23325) ) ;
 assign ng27272 = ( (~ ng826)  &  ng1071 ) | ( ng1071  &  wire3293 ) | ( ng826  &  (~ ng23340)  &  (~ wire3293) ) ;
 assign ng29198 = ( (~ ng826)  &  ng1104 ) | ( ng826  &  ng11902  &  ng27551 ) | ( ng826  &  (~ ng11902)  &  (~ ng27551) ) ;
 assign ng27763 = ( ng1136  &  wire3697 ) | ( (~ wire3697)  &  (~ wire34737)  &  (~ wire34738) ) ;
 assign ng30485 = ( (~ ng823)  &  ng1006 ) | ( ng823  &  wire4359 ) | ( ng823  &  wire4360 ) ;
 assign ng18707 = ( ng1315  &  (~ ng1240) ) | ( (~ ng1315)  &  ng1243 ) ;
 assign ng27286 = ( (~ ng1309)  &  ng1265 ) | ( (~ ng22615)  &  ng1265 ) | ( ng1309  &  ng22615  &  (~ ng22069) ) ;
 assign ng13430 = ( (~ ng970) ) ;
 assign ng16671 = ( ng1315  &  ng1196 ) | ( (~ ng1315)  &  ng1316 ) ;
 assign ng20896 = ( ng1386  &  ng13126 ) | ( (~ ng1326)  &  (~ ng13126) ) ;
 assign ng20950 = ( ng1395  &  ng13126 ) | ( (~ ng1332)  &  (~ ng13126) ) ;
 assign ng25267 = ( ng1422  &  ng13126 ) | ( (~ ng13126)  &  wire34912 ) | ( (~ ng13126)  &  wire34913 ) ;
 assign ng22179 = ( (~ ng823)  &  ng1516 ) | ( ng1516  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng1476) ) ;
 assign ng25235 = ( (~ ng13110)  &  ng1557 ) | ( (~ ng826)  &  ng1557 ) | ( ng13110  &  ng826  &  (~ ng1471) ) ;
 assign ng30651 = ( (~ ng826)  &  ng1612 ) | ( ng826  &  wire36135 ) | ( ng826  &  wire36136 ) ;
 assign ng30272 = ( wire4155 ) | ( (~ ng823)  &  ng1633 ) ;
 assign ng30650 = ( (~ ng823)  &  ng1606 ) | ( ng823  &  ng30015 ) ;
 assign ng28749 = ( (~ ng826)  &  ng1789 ) | ( ng826  &  ng27566 ) ;
 assign ng11546 = ( (~ ng1486) ) ;
 assign ng22098 = ( (~ ng823)  &  ng2225 ) | ( ng2225  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2185) ) ;
 assign ng22154 = ( (~ ng823)  &  ng2234 ) | ( ng2234  &  (~ ng2257) ) | ( ng823  &  (~ ng2200)  &  ng2257 ) ;
 assign ng26823 = ( (~ ng826)  &  ng2513 ) | ( ng826  &  wire3151 ) ;
 assign ng30707 = ( (~ ng826)  &  ng2390 ) | ( ng826  &  ng30033 ) ;
 assign ng24238 = ( (~ ng853)  &  ng2554 ) | ( ng853  &  ng11678  &  wire33792 ) ;
 assign ng24237 = ( (~ ng823)  &  ng2543 ) | ( ng823  &  ng11678  &  wire33551 ) ;
 assign ng24537 = ( wire4135 ) | ( (~ ng1312)  &  ng2664 ) ;
 assign ng28363 = ( wire4133 ) | ( (~ ng1312)  &  ng2682 ) ;
 assign ng21974 = ( ng2707  &  (~ ng2714)  &  ng10747 ) | ( ng2707  &  ng2714  &  ng10747  &  wire3248 ) | ( (~ ng2707)  &  ng2714  &  ng10747  &  (~ wire3248) ) ;
 assign ng26795 = ( (~ ng26677)  &  wire36183 ) | ( (~ ng24043)  &  wire36184 ) ;
 assign ng20981 = ( ng2775  &  ng11733 ) | ( (~ ng2707)  &  (~ ng11733) ) ;
 assign ng21045 = ( ng2791  &  ng13146 ) | ( (~ ng2740)  &  (~ ng13146) ) ;
 assign ng20919 = ( ng2800  &  ng13146 ) | ( (~ ng2766)  &  (~ ng13146) ) ;
 assign ng21046 = ( ng2802  &  wire3216 ) | ( (~ wire3216)  &  wire33957 ) | ( (~ wire3216)  &  wire33958 ) ;
 assign ng29975 = ( wire3835 ) | ( wire4121 ) | ( wire3227  &  (~ ng27897) ) ;
 assign ng30911 = ( wire3833 ) | ( wire4115 ) | ( (~ ng29748)  &  wire3229 ) ;
 assign ng30987 = ( wire4104 ) | ( wire4105 ) | ( wire36190 ) ;
 assign ng22002 = ( wire36177 ) | ( (~ ng21796)  &  (~ wire4250)  &  (~ wire36175) ) ;
 assign ng16857 = ( ng3050  &  (~ ng2987) ) | ( ng2987  &  ng3069 ) ;
 assign ng21964 = ( ng2990  &  ng12999  &  ng12988 ) | ( (~ ng2990)  &  (~ ng12999)  &  ng12988 ) | ( (~ ng2990)  &  ng12999  &  (~ ng12988) ) | ( ng2990  &  (~ ng12999)  &  (~ ng12988) ) ;
 assign ng19152 = ( pg51 ) | ( ng2933 ) ;
 assign ng29656 = ( (~ wire7046)  &  (~ wire7048)  &  (~ wire34087) ) ;
 assign ng22025 = ( (~ ng826)  &  ng142 ) | ( ng142  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng105) ) ;
 assign ng22063 = ( (~ ng853)  &  ng150 ) | ( ng150  &  (~ ng2257) ) | ( ng853  &  (~ ng117)  &  ng2257 ) ;
 assign ng22081 = ( ng160  &  ng15970 ) | ( (~ ng15970)  &  wire31159 ) | ( (~ ng15970)  &  wire31160 ) ;
 assign ng25218 = ( (~ ng13110)  &  ng171 ) | ( (~ ng853)  &  ng171 ) | ( ng13110  &  ng853  &  (~ ng101) ) ;
 assign ng30261 = ( (~ ng826)  &  ng186 ) | ( ng826  &  wire5356 ) | ( ng826  &  wire35375 ) ;
 assign ng30653 = ( (~ ng853)  &  ng246 ) | ( ng853  &  wire36064 ) | ( ng853  &  wire36065 ) ;
 assign ng30661 = ( (~ ng826)  &  ng267 ) | ( ng826  &  ng30021 ) ;
 assign ng27265 = ( ng361  &  (~ ng853) ) | ( ng361  &  wire3290 ) | ( ng853  &  (~ wire3290)  &  (~ ng21976) ) ;
 assign ng29197 = ( (~ ng823)  &  ng420 ) | ( ng823  &  ng11860  &  ng27529 ) | ( ng823  &  (~ ng11860)  &  (~ ng27529) ) ;
 assign ng26807 = ( wire4080 ) | ( (~ ng853)  &  ng435 ) ;
 assign ng30700 = ( (~ ng823)  &  ng316 ) | ( ng823  &  ng30030 ) ;
 assign ng29172 = ( wire36193 ) | ( (~ ng13165)  &  ng17051  &  (~ ng27834) ) ;
 assign ng11495 = ( (~ ng97) ) ;
 assign ng24207 = ( (~ ng823)  &  ng478 ) | ( ng823  &  ng11624  &  wire31271 ) ;
 assign ng24228 = ( ng471  &  (~ ng853) ) | ( ng853  &  ng11624  &  wire31067 ) ;
 assign ng27261 = ( (~ ng1309)  &  ng576 ) | ( (~ ng22578)  &  ng576 ) | ( ng1309  &  ng22578  &  (~ ng23360) ) ;
 assign ng27295 = ( (~ ng1312)  &  ng583 ) | ( (~ ng22578)  &  ng583 ) | ( ng1312  &  ng22578  &  (~ ng23368) ) ;
 assign ng28345 = ( (~ ng1309)  &  ng614 ) | ( ng1309  &  wire4415 ) | ( ng1309  &  wire36086 ) ;
 assign ng26545 = ( (~ ng1312)  &  ng493 ) | ( ng1312  &  ng12245  &  wire3444 ) ;
 assign ng13415 = ( (~ ng285) ) ;
 assign ng28668 = ( (~ ng686)  &  ng692  &  ng10677 ) | ( ng686  &  ng692  &  ng10677  &  wire3380 ) | ( ng686  &  (~ ng692)  &  ng10677  &  (~ wire3380) ) ;
 assign ng20922 = ( ng709  &  ng13113 ) | ( (~ ng646)  &  (~ ng13113) ) ;
 assign ng20989 = ( ng713  &  ng11721 ) | ( (~ ng672)  &  (~ ng11721) ) ;
 assign ng20881 = ( ng727  &  ng13113 ) | ( (~ ng692)  &  (~ ng13113) ) ;
 assign ng20992 = ( ng731  &  wire3205 ) | ( (~ wire3205)  &  wire31469 ) | ( (~ wire3205)  &  wire31470 ) ;
 assign ng22145 = ( (~ ng823)  &  ng819 ) | ( ng819  &  (~ ng2257) ) | ( ng823  &  (~ ng785)  &  ng2257 ) ;
 assign ng22040 = ( (~ ng853)  &  ng829 ) | ( ng829  &  (~ ng2257) ) | ( ng853  &  (~ ng793)  &  ng2257 ) ;
 assign ng22088 = ( (~ ng823)  &  ng843 ) | ( ng843  &  (~ ng2257) ) | ( ng823  &  (~ ng809)  &  ng2257 ) ;
 assign ng25231 = ( (~ ng13110)  &  ng864 ) | ( (~ ng823)  &  ng864 ) | ( ng13110  &  ng823  &  (~ ng785) ) ;
 assign ng30662 = ( (~ ng853)  &  ng933 ) | ( ng853  &  ng30016 ) ;
 assign ng30271 = ( (~ ng823)  &  ng948 ) | ( ng823  &  ng29677 ) ;
 assign ng30682 = ( (~ ng853)  &  ng960 ) | ( ng853  &  wire32160 ) | ( ng853  &  wire32161 ) ;
 assign ng27257 = ( ng1041  &  (~ ng826) ) | ( ng1041  &  wire3293 ) | ( ng826  &  (~ wire3293)  &  (~ ng23325) ) ;
 assign ng27283 = ( (~ ng823)  &  ng1060 ) | ( ng1060  &  wire3293 ) | ( ng823  &  (~ ng23340)  &  (~ wire3293) ) ;
 assign ng28747 = ( wire4030 ) | ( wire36198 ) ;
 assign ng26814 = ( (~ ng823)  &  ng1128 ) | ( ng823  &  wire3157 ) ;
 assign ng30470 = ( (~ ng826)  &  ng1005 ) | ( ng826  &  wire4359 ) | ( ng826  &  wire4360 ) ;
 assign ng23110 = ( (~ ng826)  &  ng1167 ) | ( ng826  &  wire32219 ) | ( ng826  &  wire32220 ) ;
 assign ng27299 = ( (~ ng1315)  &  ng1261 ) | ( (~ ng22615)  &  ng1261 ) | ( ng1315  &  ng22615  &  (~ ng23364) ) ;
 assign ng13431 = ( (~ ng972) ) ;
 assign ng21969 = ( ng1319  &  (~ ng1326)  &  ng10706 ) | ( ng1319  &  ng1326  &  ng10706  &  wire3253 ) | ( (~ ng1319)  &  ng1326  &  ng10706  &  (~ wire3253) ) ;
 assign ng27718 = ( (~ ng1365)  &  ng1372  &  ng10706 ) | ( ng1372  &  (~ ng23979)  &  ng10706 ) | ( ng1365  &  (~ ng1372)  &  ng23979  &  ng10706 ) ;
 assign ng20927 = ( ng1394  &  ng13134 ) | ( (~ ng1332)  &  (~ ng13134) ) ;
 assign ng20994 = ( ng1401  &  ng13126 ) | ( (~ ng1358)  &  (~ ng13126) ) ;
 assign ng20883 = ( ng1412  &  ng13134 ) | ( (~ ng1378)  &  (~ ng13134) ) ;
 assign ng25243 = ( (~ ng13110)  &  ng1558 ) | ( (~ ng823)  &  ng1558 ) | ( ng13110  &  ng823  &  (~ ng1471) ) ;
 assign ng30683 = ( (~ ng826)  &  ng1576 ) | ( ng826  &  wire35390 ) | ( ng826  &  wire35391 ) ;
 assign ng30299 = ( (~ ng823)  &  ng1588 ) | ( ng823  &  wire6791 ) | ( ng823  &  wire34395 ) ;
 assign ng30644 = ( (~ ng826)  &  ng1603 ) | ( ng826  &  ng30015 ) ;
 assign ng27287 = ( (~ ng853)  &  ng1727 ) | ( ng1727  &  wire3309 ) | ( ng853  &  (~ ng23335)  &  (~ wire3309) ) ;
 assign ng26130 = ( wire36276 ) | ( wire36277 ) | ( wire36278 ) | ( wire36279 ) ;
 assign ng27323 = ( ng2448  &  (~ ng823) ) | ( ng2448  &  wire3313 ) | ( ng823  &  (~ ng23353)  &  (~ wire3313) ) ;
 assign ng26826 = ( (~ ng823)  &  ng2516 ) | ( ng823  &  wire3151 ) ;
 assign ng30505 = ( (~ ng826)  &  ng2393 ) | ( ng826  &  ng29920 ) ;
 assign ng24226 = ( (~ ng823)  &  ng2553 ) | ( ng823  &  ng11678  &  wire33792 ) ;
 assign ng24250 = ( (~ ng853)  &  ng2546 ) | ( ng853  &  ng11678  &  wire33551 ) ;
 assign ng27310 = ( (~ ng1309)  &  ng2650 ) | ( (~ ng22687)  &  ng2650 ) | ( ng1309  &  ng22687  &  (~ ng23381) ) ;
 assign ng24547 = ( wire3931 ) | ( (~ ng1315)  &  ng2667 ) ;
 assign ng13459 = ( (~ ng2528) ) ;
 assign ng20789 = ( (~ ng1312)  &  ng2714  &  wire3248 ) | ( (~ ng2704)  &  ng2714  &  wire3248 ) | ( (~ ng1312)  &  (~ ng2714)  &  (~ wire3248) ) | ( (~ ng2704)  &  (~ ng2714)  &  (~ wire3248) ) ;
 assign ng27243 = ( (~ ng1312)  &  (~ ng2753)  &  ng24043 ) | ( (~ ng2704)  &  (~ ng2753)  &  ng24043 ) | ( (~ ng1312)  &  ng2753  &  (~ ng24043) ) | ( (~ ng2704)  &  ng2753  &  (~ ng24043) ) ;
 assign ng21004 = ( ng2778  &  ng11733 ) | ( (~ ng2727)  &  (~ ng11733) ) ;
 assign ng21027 = ( ng2788  &  ng13146 ) | ( (~ ng2746)  &  (~ ng13146) ) ;
 assign ng21094 = ( ng2796  &  ng11733 ) | ( (~ ng2760)  &  (~ ng11733) ) ;
 assign ng21029 = ( ng2806  &  wire3206 ) | ( (~ wire3206)  &  wire33977 ) | ( (~ wire3206)  &  wire33978 ) ;
 assign ng20497 = ( pg3234 ) | ( ng3079 ) ;
 assign ng29976 = ( wire36284 ) | ( ng1196  &  (~ ng1243)  &  (~ ng27900) ) ;
 assign ng30914 = ( wire36288 ) | ( ng1890  &  (~ ng1937)  &  (~ ng29713) ) ;
 assign ng30984 = ( wire3885 ) | ( wire36290 ) ;
 assign ng26786 = ( ng3024  &  (~ ng3010)  &  ng21796 ) | ( ng3024  &  ng3010  &  ng21796  &  wire3403 ) | ( (~ ng3024)  &  ng3010  &  ng21796  &  (~ wire3403) ) ;
 assign ng21966 = ( ng3083  &  ng11621  &  ng13399 ) | ( (~ ng3083)  &  (~ ng11621)  &  ng13399 ) | ( (~ ng3083)  &  ng11621  &  (~ ng13399) ) | ( ng3083  &  (~ ng11621)  &  (~ ng13399) ) ;
 assign ng18837 = ( ng3077  &  ng2987 ) | ( (~ ng2987)  &  ng3059 ) ;
 assign ng20825 = ( pg8021 ) | ( wire35371 ) | ( wire35029  &  wire35030 ) ;
 assign ng29166 = ( (~ wire36306)  &  (~ wire36307)  &  (~ wire36311) ) ;
 assign ng22027 = ( (~ ng823)  &  ng143 ) | ( ng143  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng105) ) ;
 assign ng22048 = ( (~ ng823)  &  ng152 ) | ( ng152  &  (~ ng2257) ) | ( ng823  &  (~ ng117)  &  ng2257 ) ;
 assign ng22102 = ( ng161  &  ng15950 ) | ( (~ ng15950)  &  wire31159 ) | ( (~ ng15950)  &  wire31160 ) ;
 assign ng25212 = ( (~ ng13110)  &  ng173 ) | ( (~ ng823)  &  ng173 ) | ( ng13110  &  ng823  &  (~ ng101) ) ;
 assign ng30267 = ( (~ ng823)  &  ng189 ) | ( ng823  &  wire5356 ) | ( ng823  &  wire35375 ) ;
 assign ng30646 = ( (~ ng823)  &  ng243 ) | ( ng823  &  wire36064 ) | ( ng823  &  wire36065 ) ;
 assign ng29109 = ( (~ ng26869)  &  wire36314 ) | ( (~ ng28634)  &  (~ ng26869)  &  wire36312 ) ;
 assign ng27260 = ( ng384  &  (~ ng826) ) | ( ng384  &  wire3290 ) | ( ng826  &  (~ wire3290)  &  (~ ng23331) ) ;
 assign ng29194 = ( (~ ng826)  &  ng417 ) | ( ng826  &  ng11860  &  ng27529 ) | ( ng826  &  (~ ng11860)  &  (~ ng27529) ) ;
 assign ng26805 = ( (~ ng826)  &  ng438 ) | ( ng826  &  wire3156 ) ;
 assign ng30699 = ( (~ ng826)  &  ng315 ) | ( ng826  &  ng30030 ) ;
 assign ng26655 = ( wire3815 ) | ( (~ ng826)  &  ng403 ) | ( ng403  &  (~ ng2257) ) ;
 assign ng11491 = ( (~ ng113) ) ;
 assign ng24178 = ( (~ ng826)  &  ng477 ) | ( ng826  &  ng11624  &  wire31271 ) ;
 assign ng12457 = ( wire3049 ) | ( wire7006 ) | ( wire34114 ) | ( wire34118 ) ;
 assign ng27311 = ( (~ ng1315)  &  ng581 ) | ( (~ ng22578)  &  ng581 ) | ( ng1315  &  ng22578  &  (~ ng23368) ) ;
 assign ng24519 = ( wire3808 ) | ( (~ ng1315)  &  ng602 ) ;
 assign ng26553 = ( (~ ng1315)  &  ng496 ) | ( ng1315  &  ng12245  &  wire3444 ) ;
 assign ng13414 = ( (~ ng283) ) ;
 assign ng20875 = ( ng699  &  ng13123 ) | ( (~ ng640)  &  (~ ng13123) ) ;
 assign ng20903 = ( ng708  &  ng13123 ) | ( (~ ng646)  &  (~ ng13123) ) ;
 assign ng20968 = ( ng717  &  ng13123 ) | ( (~ ng666)  &  (~ ng13123) ) ;
 assign ng20876 = ( ng726  &  ng13123 ) | ( (~ ng692)  &  (~ ng13123) ) ;
 assign ng25260 = ( ng735  &  ng13123 ) | ( (~ ng13123)  &  wire31760 ) | ( (~ ng13123)  &  wire31761 ) ;
 assign ng22126 = ( (~ ng826)  &  ng818 ) | ( ng818  &  (~ ng2257) ) | ( ng826  &  (~ ng785)  &  ng2257 ) ;
 assign ng22034 = ( (~ ng826)  &  ng833 ) | ( ng833  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng797) ) ;
 assign ng22068 = ( (~ ng826)  &  ng842 ) | ( ng842  &  (~ ng2257) ) | ( ng826  &  (~ ng809)  &  ng2257 ) ;
 assign ng22129 = ( ng851  &  ng15970 ) | ( (~ ng15970)  &  wire32020 ) | ( (~ ng15970)  &  wire32021 ) ;
 assign ng30286 = ( (~ ng826)  &  ng891 ) | ( ng826  &  wire5326 ) | ( ng826  &  wire35384 ) ;
 assign ng30265 = ( (~ ng826)  &  ng945 ) | ( ng826  &  ng29677 ) ;
 assign ng25042 = ( (~ ng780)  &  ng17197 ) | ( (~ ng853)  &  ng780  &  (~ ng17197) ) | ( ng780  &  (~ ng2257)  &  (~ ng17197) ) ;
 assign ng29580 = ( ng740  &  (~ ng17031)  &  wire3389 ) | ( (~ ng740)  &  (~ ng17031)  &  (~ wire3389) ) ;
 assign ng27297 = ( ng1063  &  (~ ng853) ) | ( ng1063  &  wire3293 ) | ( ng853  &  (~ ng23340)  &  (~ wire3293) ) ;
 assign ng29209 = ( (~ ng853)  &  ng1110 ) | ( ng853  &  ng11902  &  ng27551 ) | ( ng853  &  (~ ng11902)  &  (~ ng27551) ) ;
 assign ng26818 = ( (~ ng853)  &  ng1131 ) | ( ng853  &  wire3157 ) ;
 assign ng30705 = ( (~ ng853)  &  ng1004 ) | ( ng853  &  ng30031 ) ;
 assign ng24223 = ( (~ ng853)  &  ng1166 ) | ( ng853  &  ng11647  &  wire32128 ) ;
 assign ng13432 = ( (~ ng974) ) ;
 assign ng20717 = ( (~ ng1312)  &  ng1326  &  wire3253 ) | ( (~ ng1316)  &  ng1326  &  wire3253 ) | ( (~ ng1312)  &  (~ ng1326)  &  (~ wire3253) ) | ( (~ ng1316)  &  (~ ng1326)  &  (~ wire3253) ) ;
 assign ng28321 = ( (~ ng1372)  &  ng1378  &  ng10706 ) | ( ng1372  &  ng1378  &  ng10706  &  wire3377 ) | ( ng1372  &  (~ ng1378)  &  ng10706  &  (~ wire3377) ) ;
 assign ng20949 = ( ng1390  &  ng11726 ) | ( (~ ng1339)  &  (~ ng11726) ) ;
 assign ng21015 = ( ng1399  &  ng11726 ) | ( (~ ng1358)  &  (~ ng11726) ) ;
 assign ng21070 = ( ng1408  &  ng11726 ) | ( (~ ng1372)  &  (~ ng11726) ) ;
 assign ng25249 = ( (~ ng13110)  &  ng1556 ) | ( (~ ng853)  &  ng1556 ) | ( ng13110  &  ng853  &  (~ ng1471) ) ;
 assign ng30663 = ( (~ ng853)  &  ng1618 ) | ( ng853  &  wire36135 ) | ( ng853  &  wire36136 ) ;
 assign ng30302 = ( (~ ng853)  &  ng1591 ) | ( ng853  &  wire6791 ) | ( ng853  &  wire34395 ) ;
 assign ng30288 = ( (~ ng853)  &  ng1645 ) | ( ng853  &  ng29680 ) ;
 assign ng26531 = ( ng1457  &  ng25938 ) | ( ng1457  &  (~ ng1462)  &  (~ ng17031) ) | ( (~ ng1457)  &  (~ ng25938)  &  ng1462  &  (~ ng17031) ) ;
 assign ng11547 = ( (~ ng1481) ) ;
 assign ng28903 = ( wire4703 ) | ( wire35917 ) ;
 assign ng29226 = ( (~ ng853)  &  ng2498 ) | ( ng853  &  ng12005  &  ng27577 ) | ( ng853  &  (~ ng12005)  &  (~ ng27577) ) ;
 assign ng26827 = ( (~ ng853)  &  ng2519 ) | ( ng853  &  wire3151 ) ;
 assign ng30566 = ( (~ ng853)  &  ng2392 ) | ( ng853  &  ng30033 ) ;
 assign ng24214 = ( (~ ng826)  &  ng2552 ) | ( ng826  &  ng11678  &  wire33792 ) ;
 assign ng12499 = ( wire3049 ) | ( wire5775 ) | ( wire35225 ) | ( wire35229 ) ;
 assign ng26575 = ( (~ ng1309)  &  ng2565 ) | ( ng1309  &  ng12352  &  wire3435 ) ;
 assign ng13460 = ( (~ ng2354) ) ;
 assign ng20375 = ( (~ ng1315)  &  ng2733 ) | ( ng1315  &  wire31471  &  wire31472 ) ;
 assign ng27724 = ( (~ ng2753)  &  ng2760  &  ng10747 ) | ( ng2760  &  ng10747  &  (~ ng24043) ) | ( ng2753  &  (~ ng2760)  &  ng10747  &  ng24043 ) ;
 assign ng20982 = ( ng2780  &  ng13145 ) | ( (~ ng2727)  &  (~ ng13145) ) ;
 assign ng21044 = ( ng2789  &  ng13145 ) | ( (~ ng2746)  &  (~ ng13145) ) ;
 assign ng21082 = ( ng2798  &  ng13145 ) | ( (~ ng2760)  &  (~ ng13145) ) ;
 assign ng21047 = ( ng2807  &  ng10747 ) | ( (~ ng10747)  &  wire33977 ) | ( (~ ng10747)  &  wire33978 ) ;
 assign ng20884 = ( (~ pg3234)  &  ng3054 ) ;
 assign ng29977 = ( wire36321 ) | ( ng1196  &  (~ ng1243)  &  (~ ng27802) ) ;
 assign ng30913 = ( wire36323 ) | ( ng1890  &  (~ ng1937)  &  (~ ng29705) ) ;
 assign ng30985 = ( wire3714 ) | ( wire36325 ) ;
 assign ng26031 = ( ng3010  &  ng21796  &  wire3403 ) | ( (~ ng3010)  &  ng21796  &  (~ wire3403) ) ;
 assign ng16824 = ( ng3062  &  ng2987 ) | ( ng3043  &  (~ ng2987) ) ;
 assign ng16566 = ( pg3231  &  (~ ng11621)  &  ng13399 ) | ( (~ ng3120)  &  (~ ng11621)  &  ng13399 ) | ( pg3231  &  ng11621  &  (~ ng13399) ) | ( (~ ng3120)  &  ng11621  &  (~ ng13399) ) | ( (~ pg3231)  &  ng3120  &  ng11621  &  ng13399 ) | ( (~ pg3231)  &  ng3120  &  (~ ng11621)  &  (~ ng13399) ) ;
 assign ng18868 = ( ng3078  &  ng2987 ) | ( (~ ng2987)  &  ng3060 ) ;
 assign ng20417 = ( pg7334  &  ng2879 ) | ( ng2963  &  (~ ng2879) ) ;
 assign ng18885 = ( ng2874  &  ng2879 ) | ( ng2200  &  (~ ng2879) ) ;
 assign ng18782 = ( ng1315  &  ng559 ) | ( (~ ng1315)  &  ng3084 ) ;
 assign ng29978 = ( wire36327 ) | ( ng1196  &  (~ ng1243)  &  (~ ng27814) ) ;
 assign ng30940 = ( wire36344 ) | ( ng1890  &  (~ ng30034)  &  ng30035 ) | ( ng1890  &  ng30034  &  (~ ng30035) ) ;
 assign ng19173 = ( pg4323  &  ng2879 ) | ( ng2978  &  (~ ng2879) ) ;
 assign ng19149 = ( pg8175  &  ng2879 ) | ( ng2944  &  (~ ng2879) ) ;
 assign ng17222 = ( ng1309  &  ng1245 ) | ( (~ ng1309)  &  ng3085 ) ;
 assign ng29979 = ( wire36347 ) | ( ng1196  &  (~ ng1243)  &  (~ ng27827) ) ;
 assign ng30915 = ( wire36349 ) | ( ng1890  &  (~ ng1937)  &  (~ ng29721) ) ;
 assign ng21878 = ( wire3639 ) | ( pg7519  &  ng2879 ) ;
 assign ng20874 = ( wire3621 ) | ( pg8096  &  ng2879 ) ;
 assign ng17225 = ( ng1312  &  ng1245 ) | ( (~ ng1312)  &  ng3086 ) ;
 assign ng30989 = ( wire36364 ) | ( ng2584  &  (~ ng30926)  &  ng30927 ) | ( ng2584  &  ng30926  &  (~ ng30927) ) ;
 assign ng25202 = ( wire3594 ) | ( ng3032  &  ng24446 ) | ( (~ ng24446)  &  wire36370 ) ;
 assign ng19184 = ( pg4590  &  ng2879 ) | ( ng2975  &  (~ ng2879) ) ;
 assign ng19144 = ( pg8023  &  ng2879 ) | ( ng2947  &  (~ ng2879) ) ;
 assign ng17234 = ( ng1315  &  ng1245 ) | ( (~ ng1315)  &  ng3087 ) ;
 assign ng25265 = ( wire4476 ) | ( wire4477 ) | ( wire4478 ) ;
 assign ng24446 = ( (~ ng3028)  &  ng3036  &  ng21711 ) | ( (~ ng3028)  &  ng3036  &  (~ wire3292) ) | ( ng3028  &  (~ ng3036)  &  (~ wire3292) ) | ( ng3028  &  ng3036  &  ng21711  &  wire3292 ) ;
 assign ng26798 = ( (~ ng2900)  &  ng2908  &  (~ wire3139) ) | ( ng2900  &  ng2908  &  (~ wire3139)  &  wire3395 ) | ( ng2900  &  (~ ng2908)  &  (~ wire3139)  &  (~ wire3395) ) ;
 assign ng18852 = ( ng2941  &  ng2879 ) | ( ng1481  &  (~ ng2879) ) ;
 assign ng17224 = ( ng1309  &  ng1939 ) | ( (~ ng1309)  &  ng3091 ) ;
 assign ng30287 = ( (~ ng823)  &  ng1570 ) | ( ng823  &  wire6292 ) | ( ng823  &  wire34916 ) ;
 assign ng22193 = ( (~ ng823)  &  ng2210 ) | ( ng2210  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2170) ) ;
 assign ng22099 = ( (~ ng826)  &  ng2227 ) | ( ng2227  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2190) ) ;
 assign ng16835 = ( ng3048  &  (~ ng2987) ) | ( ng2987  &  ng3067 ) ;
 assign ng18804 = ( (~ ng2987)  &  ng3058 ) | ( ng2987  &  ng3076 ) ;
 assign ng21989 = ( wire36379 ) | ( wire3139  &  (~ wire3564)  &  (~ wire36377) ) ;
 assign ng18835 = ( ng2944  &  ng2879 ) | ( ng1486  &  (~ ng2879) ) ;
 assign ng17228 = ( ng1312  &  ng1939 ) | ( (~ ng1312)  &  ng3092 ) ;
 assign ng30671 = ( (~ ng853)  &  ng1627 ) | ( ng853  &  wire35900 ) | ( ng853  &  wire35901 ) ;
 assign ng22200 = ( (~ ng853)  &  ng2208 ) | ( ng2208  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2170) ) ;
 assign ng22115 = ( (~ ng853)  &  ng2223 ) | ( ng2223  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2185) ) ;
 assign ng16851 = ( ng3068  &  ng2987 ) | ( ng3049  &  (~ ng2987) ) ;
 assign ng18755 = ( ng3075  &  ng2987 ) | ( ng3057  &  (~ ng2987) ) ;
 assign ng23357 = ( wire3545 ) | ( wire36383 ) ;
 assign ng18821 = ( ng2947  &  ng2879 ) | ( ng1491  &  (~ ng2879) ) ;
 assign ng30273 = ( (~ ng826)  &  ng1639 ) | ( ng826  &  ng29680 ) ;
 assign ng18743 = ( (~ ng1315)  &  ng1937 ) | ( ng1315  &  (~ ng1934) ) ;
 assign ng22045 = ( (~ ng826)  &  ng2218 ) | ( ng2218  &  (~ ng2257) ) | ( ng826  &  ng2257  &  (~ ng2175) ) ;
 assign ng22138 = ( (~ ng853)  &  ng2226 ) | ( ng2226  &  (~ ng2257) ) | ( ng853  &  ng2257  &  (~ ng2190) ) ;
 assign ng27769 = ( (~ ng823)  &  ng2524 ) | ( ng823  &  (~ ng24038)  &  wire33948 ) | ( ng2524  &  (~ ng24038)  &  (~ wire33948) ) ;
 assign ng24476 = ( wire3527 ) | ( wire3528 ) | ( wire3529 ) ;
 assign ng18803 = ( ng2953  &  ng2879 ) | ( ng1496  &  (~ ng2879) ) ;
 assign ng25938 = ( (~ ng1466)  &  ng1462  &  ng13165 ) | ( (~ ng1466)  &  ng1462  &  ng17197 ) | ( ng1466  &  (~ ng1462)  &  ng17197 ) | ( ng1462  &  ng13165  &  (~ ng17197) ) ;
 assign ng21845 = ( wire3142 ) | ( (~ ng1315)  &  ng1934 ) ;
 assign ng22060 = ( (~ ng823)  &  ng2219 ) | ( ng2219  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2175) ) ;
 assign ng22116 = ( (~ ng823)  &  ng2228 ) | ( ng2228  &  (~ ng2257) ) | ( ng823  &  ng2257  &  (~ ng2190) ) ;
 assign ng28774 = ( wire3515 ) | ( wire36388 ) ;
 assign ng25199 = ( wire36391 ) | ( ng2920  &  wire3529 ) | ( ng2920  &  wire36387 ) ;
 assign ng19154 = ( pg8251  &  ng2879 ) | ( ng2874  &  (~ ng2879) ) ;
 assign ng19172 = ( pg4321  &  ng2879 ) | ( ng2953  &  (~ ng2879) ) ;
 assign ng27274 = ( ng1724  &  (~ ng823) ) | ( ng1724  &  wire3309 ) | ( ng823  &  (~ ng23335)  &  (~ wire3309) ) ;
 assign ng23400 = ( ng1836  &  (~ ng826) ) | ( ng826  &  (~ ng11666)  &  wire32979 ) ;
 assign ng20936 = ( ng2085  &  ng13142 ) | ( (~ ng2033)  &  (~ ng13142) ) ;
 assign ng21039 = ( ng2093  &  ng11730 ) | ( (~ ng2052)  &  (~ ng11730) ) ;
 assign ng20917 = ( ng2107  &  ng13137 ) | ( (~ ng2072)  &  (~ ng13137) ) ;
 assign ng22249 = ( (~ ng1309)  &  ng2118 ) | ( ng2118  &  (~ ng2010) ) | ( (~ ng2010)  &  (~ ng13142) ) ;
 assign ng27334 = ( ng2451  &  (~ ng853) ) | ( ng2451  &  wire3313 ) | ( ng853  &  (~ ng23353)  &  (~ wire3313) ) ;
 assign ng16181 = ( ng2934  &  ng11330  &  ng11263 ) | ( (~ ng2934)  &  (~ ng11330)  &  ng11263 ) | ( (~ ng2934)  &  ng11330  &  (~ ng11263) ) | ( ng2934  &  (~ ng11330)  &  (~ ng11263) ) ;
 assign ng21880 = ( wire3488 ) | ( ng2877  &  (~ ng2879) ) ;
 assign ng20376 = ( pg6895  &  ng2879 ) | ( ng2966  &  (~ ng2879) ) ;
 assign ng27330 = ( ng1772  &  (~ ng853) ) | ( ng1772  &  wire3309 ) | ( ng853  &  (~ ng22016)  &  (~ wire3309) ) ;
 assign ng23137 = ( (~ ng853)  &  ng1869 ) | ( ng853  &  (~ wire33063)  &  (~ wire33064) ) ;
 assign ng20954 = ( ng2086  &  ng13137 ) | ( (~ ng2033)  &  (~ ng13137) ) ;
 assign ng21020 = ( ng2095  &  ng13137 ) | ( (~ ng2052)  &  (~ ng13137) ) ;
 assign ng20937 = ( ng2105  &  ng11730 ) | ( (~ ng2072)  &  (~ ng11730) ) ;
 assign ng25279 = ( ng2114  &  ng11730 ) | ( (~ ng11730)  &  wire36445 ) | ( (~ ng11730)  &  wire36446 ) ;
 assign ng16132 = ( ng2962  &  ng11188  &  ng11262 ) | ( (~ ng2962)  &  (~ ng11188)  &  ng11262 ) | ( (~ ng2962)  &  ng11188  &  (~ ng11262) ) | ( ng2962  &  (~ ng11188)  &  (~ ng11262) ) ;
 assign ng18883 = ( ng2935  &  ng2879 ) | ( ng1471  &  (~ ng2879) ) ;
 assign ng18836 = ( ng2966  &  ng2879 ) | ( ng2170  &  (~ ng2879) ) ;
 assign ng26811 = ( wire3404 ) | ( (~ ng826)  &  ng1810 ) ;
 assign ng24218 = ( ng1846  &  (~ ng826) ) | ( ng826  &  ng11666  &  wire32703 ) ;
 assign ng13182 = ( wire36455 ) | ( wire36456 ) ;
 assign ng20977 = ( ng2084  &  ng11730 ) | ( (~ ng2033)  &  (~ ng11730) ) ;
 assign ng21040 = ( ng2098  &  ng13137 ) | ( (~ ng2046)  &  (~ ng13137) ) ;
 assign ng21080 = ( ng2102  &  ng11730 ) | ( (~ ng2066)  &  (~ ng11730) ) ;
 assign ng25271 = ( ng2116  &  ng13137 ) | ( (~ ng13137)  &  wire36445 ) | ( (~ ng13137)  &  wire36446 ) ;
 assign ng26532 = ( ng25940  &  ng2151 ) | ( (~ ng2156)  &  ng2151  &  (~ ng17031) ) | ( (~ ng25940)  &  ng2156  &  (~ ng2151)  &  (~ ng17031) ) ;
 assign ng18866 = ( ng2938  &  ng2879 ) | ( ng1476  &  (~ ng2879) ) ;
 assign ng19178 = ( pg4450  &  ng2879 ) | ( ng2935  &  (~ ng2879) ) ;
 assign ng18867 = ( ng2969  &  ng2879 ) | ( ng2175  &  (~ ng2879) ) ;
 assign ng29617 = ( wire3322 ) | ( (~ ng823)  &  ng1694 ) ;
 assign ng24230 = ( ng1849  &  (~ ng823) ) | ( ng823  &  ng11666  &  wire32703 ) ;
 assign ng20955 = ( ng2088  &  ng13142 ) | ( (~ ng2026)  &  (~ ng13142) ) ;
 assign ng21021 = ( ng2097  &  ng13142 ) | ( (~ ng2046)  &  (~ ng13142) ) ;
 assign ng20900 = ( ng2106  &  ng13142 ) | ( (~ ng2072)  &  (~ ng13142) ) ;
 assign ng25268 = ( ng2115  &  ng13142 ) | ( (~ ng13142)  &  wire36445 ) | ( (~ ng13142)  &  wire36446 ) ;
 assign ng30291 = ( (~ ng823)  &  ng2336 ) | ( ng823  &  ng29684 ) ;
 assign ng19153 = ( pg8249  &  ng2879 ) | ( (~ ng2879)  &  ng2959 ) ;
 assign ng18906 = ( ng2972  &  ng2879 ) | ( ng2180  &  (~ ng2879) ) ;
 assign ng18957 = ( ng2963  &  ng2879 ) | ( ng2165  &  (~ ng2879) ) ;
 assign ng29184 = ( wire36458 ) | ( ng853  &  (~ ng27875)  &  wire34932 ) ;
 assign ng27332 = ( (~ ng1312)  &  ng1963 ) | ( (~ ng22651)  &  ng1963 ) | ( ng1312  &  ng22651  &  (~ ng23388) ) ;
 assign ng28357 = ( (~ ng1309)  &  ng1994 ) | ( ng1309  &  wire3168 ) | ( ng1309  &  wire36463 ) ;
 assign ng28362 = ( (~ ng1312)  &  ng1997 ) | ( ng1312  &  wire3168 ) | ( ng1312  &  wire36463 ) ;
 assign ng16692 = ( ng1890  &  ng1315 ) | ( (~ ng1315)  &  ng2010 ) ;
 assign ng28325 = ( ng2072  &  (~ ng2066)  &  (~ ng10238) ) | ( ng2072  &  ng2066  &  (~ ng10238)  &  wire3374 ) | ( (~ ng2072)  &  ng2066  &  (~ ng10238)  &  (~ wire3374) ) ;
 assign ng30301 = ( (~ ng826)  &  ng2279 ) | ( ng826  &  wire6240 ) | ( ng826  &  wire34937 ) ;
 assign ng12433 = ( (~ ng2879) ) | ( pg8021  &  (~ ng2929) ) ;
 assign ng20310 = ( pg6225  &  ng2879 ) | ( ng2972  &  (~ ng2879) ) ;
 assign ng19167 = ( pg4200  &  ng2879 ) | ( ng2938  &  (~ ng2879) ) ;
 assign ng18942 = ( ng2975  &  ng2879 ) | ( (~ ng2879)  &  ng2185 ) ;
 assign ng21882 = ( wire3101 ) | ( ng2878  &  (~ ng2879) ) ;
 assign ng11545 = ( (~ ng1491) ) ;
 assign ng27340 = ( (~ ng1315)  &  ng1961 ) | ( (~ ng22651)  &  ng1961 ) | ( ng1315  &  ng22651  &  (~ ng23388) ) ;
 assign ng24545 = ( wire3097 ) | ( (~ ng1315)  &  ng1982 ) ;
 assign ng28366 = ( (~ ng1315)  &  ng2000 ) | ( ng1315  &  wire3168 ) | ( ng1315  &  wire36463 ) ;
 assign ng28990 = ( wire4506 ) | ( wire36047 ) ;
 assign ng20353 = ( (~ ng1315)  &  ng2039 ) | ( ng1315  &  wire31471  &  wire31472 ) ;
 assign ng27722 = ( ng2066  &  (~ ng2059)  &  (~ ng10238) ) | ( ng2066  &  (~ ng10238)  &  (~ ng24009) ) | ( (~ ng2066)  &  ng2059  &  (~ ng10238)  &  ng24009 ) ;
 assign ng30300 = ( (~ ng853)  &  ng2267 ) | ( ng853  &  wire5512 ) | ( ng853  &  wire35341 ) ;
 assign ng18754 = ( ng2879  &  ng2959 ) | ( (~ ng2879)  &  ng1506 ) ;
 assign ng19163 = ( pg4090  &  ng2879 ) | ( ng2981  &  (~ ng2879) ) ;
 assign ng19162 = ( pg4088  &  ng2879 ) | ( ng2956  &  (~ ng2879) ) ;
 assign ng18968 = ( ng2978  &  ng2879 ) | ( (~ ng2879)  &  ng2190 ) ;
 assign ng18669 = ( ng1309  &  ng559 ) | ( (~ ng1309)  &  ng3210 ) ;
 assign ng28352 = ( wire3079 ) | ( (~ ng1309)  &  ng1985 ) ;
 assign ng13443 = ( (~ ng1834) ) ;
 assign ng24083 = ( pg3229  &  (~ ng1672) ) | ( (~ pg3229)  &  ng1686 ) ;
 assign ng27682 = ( (~ ng1312)  &  (~ ng2059)  &  ng24009 ) | ( (~ ng2010)  &  (~ ng2059)  &  ng24009 ) | ( (~ ng1312)  &  ng2059  &  (~ ng24009) ) | ( (~ ng2010)  &  ng2059  &  (~ ng24009) ) ;
 assign ng25246 = ( (~ ng13110)  &  ng2249 ) | ( (~ ng823)  &  ng2249 ) | ( ng13110  &  ng823  &  (~ ng2170) ) ;
 assign ng18781 = ( ng2956  &  ng2879 ) | ( (~ ng2879)  &  ng1501 ) ;
 assign ng20343 = ( pg6442  &  ng2879 ) | ( ng2969  &  (~ ng2879) ) ;
 assign ng19157 = ( pg3993  &  ng2879 ) | ( ng2941  &  (~ ng2879) ) ;
 assign ng18975 = ( ng2981  &  ng2879 ) | ( (~ ng2879)  &  ng2195 ) ;
 assign ng18719 = ( ng1312  &  ng559 ) | ( (~ ng1312)  &  ng3211 ) ;
 assign ng28356 = ( wire3050 ) | ( (~ ng1312)  &  ng1988 ) ;
 assign ng13442 = ( (~ ng1832) ) ;
 assign ng13450 = ( (~ ng1672) ) ;
 assign ng26789 = ( (~ ng24009)  &  wire36476 ) | ( (~ ng26671)  &  (~ ng24009)  &  wire36474 ) ;
 assign ng22155 = ( ng2236  &  ng15970 ) | ( (~ ng15970)  &  wire33428 ) | ( (~ ng15970)  &  wire33429 ) ;
 assign wire3193 = ( ng3139 ) | ( ng3147 ) ;
 assign wire3281 = ( ng2991 ) | ( ng2992 ) ;
 assign wire3282 = ( ng2984 ) | ( ng2985 ) ;
 assign ng26137 = ( wire34076 ) | ( wire3336  &  (~ wire31627)  &  (~ wire31628) ) ;
 assign wire3138 = ( (~ ng557)  &  (~ ng510)  &  ng525 ) ;
 assign wire3224 = ( (~ ng557)  &  ng510 ) ;
 assign wire3425 = ( wire3944 ) | ( wire3140  &  (~ wire34074)  &  (~ wire34075) ) ;
 assign wire3049 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire3142 = ( ng1315  &  (~ wire31522) ) | ( ng1315  &  (~ wire31523) ) | ( ng1315  &  (~ wire31524) ) ;
 assign ng13002 = ( wire3046 ) | ( wire7592 ) | ( wire33445 ) | ( wire33449 ) ;
 assign ng12866 = ( wire33458 ) | ( wire33459 ) ;
 assign ng12959 = ( wire33468 ) | ( wire33469 ) ;
 assign ng12978 = ( wire3046 ) | ( wire7568 ) | ( wire33475 ) | ( wire33479 ) ;
 assign ng12933 = ( wire3046 ) | ( wire7560 ) | ( wire33485 ) | ( wire33489 ) ;
 assign ng12836 = ( wire33498 ) | ( wire33499 ) ;
 assign ng12899 = ( wire3046 ) | ( wire7544 ) | ( wire33505 ) | ( wire33509 ) ;
 assign ng13022 = ( wire3046 ) | ( wire7536 ) | ( wire33515 ) | ( wire33519 ) ;
 assign ng12994 = ( wire3046 ) | ( wire7528 ) | ( wire33557 ) | ( wire33561 ) ;
 assign ng11730 = ( (~ ng1315) ) | ( (~ ng1905) ) | ( ng2039 ) | ( (~ ng1918) ) ;
 assign ng13123 = ( (~ ng1309) ) | ( ng659 ) | ( (~ ng525) ) | ( (~ ng538) ) ;
 assign ng12324 = ( wire3049 ) | ( wire7779 ) | ( wire33144 ) | ( wire33148 ) ;
 assign wire3199 = ( (~ ng1309) ) | ( (~ ng2010) ) ;
 assign ng12288 = ( wire3049 ) | ( wire8457 ) | ( wire32269 ) | ( wire32273 ) ;
 assign wire3200 = ( (~ ng1315) ) | ( (~ ng1316) ) ;
 assign wire3201 = ( (~ ng1315) ) | ( (~ ng2010) ) ;
 assign ng13134 = ( (~ ng1211) ) | ( (~ ng1309) ) | ( (~ ng1224) ) | ( ng1345 ) ;
 assign ng12233 = ( wire6694 ) | ( wire6695 ) | ( wire34530 ) | ( wire34532 ) ;
 assign ng12271 = ( wire34544 ) | ( wire34545 ) ;
 assign ng12124 = ( wire6678 ) | ( wire6679 ) | ( wire34578 ) | ( wire34580 ) ;
 assign ng12008 = ( wire6670 ) | ( wire6671 ) | ( wire34566 ) | ( wire34568 ) ;
 assign ng12306 = ( wire3049 ) | ( wire6657 ) | ( wire34553 ) | ( wire34557 ) ;
 assign ng12329 = ( wire3049 ) | ( wire6649 ) | ( wire34517 ) | ( wire34521 ) ;
 assign ng12184 = ( wire3049 ) | ( wire6641 ) | ( wire34505 ) | ( wire34509 ) ;
 assign ng12234 = ( wire3049 ) | ( wire6633 ) | ( wire34459 ) | ( wire34463 ) ;
 assign ng11965 = ( wire34496 ) | ( wire34497 ) ;
 assign ng12068 = ( wire6622 ) | ( wire6623 ) | ( wire34482 ) | ( wire34484 ) ;
 assign ng11964 = ( wire3049 ) | ( wire6609 ) | ( wire34469 ) | ( wire34473 ) ;
 assign ng12231 = ( wire3049 ) | ( wire7135 ) | ( wire33995 ) | ( wire33999 ) ;
 assign ng12305 = ( wire7132 ) | ( wire7133 ) | ( wire34006 ) | ( wire34008 ) ;
 assign ng10839 = ( wire5261 ) | ( wire5262 ) | ( wire35426 ) | ( wire35428 ) ;
 assign ng12269 = ( wire7124 ) | ( wire7125 ) | ( wire34016 ) | ( wire34018 ) ;
 assign ng10822 = ( wire3049 ) | ( wire5248 ) | ( wire35405 ) | ( wire35409 ) ;
 assign wire3351 = ( wire33998  &  (~ wire35408)  &  (~ wire35409) ) | ( wire33999  &  (~ wire35408)  &  (~ wire35409) ) ;
 assign wire3352 = ( (~ wire33998)  &  (~ wire33999)  &  wire35408 ) | ( (~ wire33998)  &  (~ wire33999)  &  wire35409 ) ;
 assign wire3926 = ( wire33988  &  wire34018 ) | ( wire33989  &  wire34018 ) | ( wire33988  &  wire34019 ) | ( wire33989  &  wire34019 ) ;
 assign wire3945 = ( (~ wire35418)  &  (~ wire35419)  &  (~ wire35428)  &  (~ wire35429) ) ;
 assign ng12180 = ( wire3046 ) | ( wire7213 ) | ( wire33934 ) | ( wire33938 ) ;
 assign ng12108 = ( wire33063 ) | ( wire33064 ) ;
 assign ng15970 = ( (~ ng826) ) | ( (~ ng2257) ) ;
 assign ng13165 = ( (~ ng853) ) | ( (~ ng2257) ) ;
 assign ng15950 = ( (~ ng823) ) | ( (~ ng2257) ) ;
 assign wire3283 = ( (~ ng1332) ) | ( (~ ng1339) ) | ( (~ ng1319) ) | ( (~ wire32567) ) ;
 assign ng23979 = ( ng1332  &  wire32566  &  wire32567  &  wire32575 ) ;
 assign ng18079 = ( (~ wire31038)  &  (~ wire31039)  &  wire31159 ) | ( (~ wire31038)  &  (~ wire31039)  &  wire31160 ) | ( wire31038  &  (~ wire31159)  &  (~ wire31160) ) | ( wire31039  &  (~ wire31159)  &  (~ wire31160) ) ;
 assign ng18183 = ( ng121  &  wire30947 ) | ( ng121  &  wire30948 ) | ( (~ ng121)  &  (~ wire30947)  &  (~ wire30948) ) ;
 assign ng18346 = ( ng105  &  wire31028 ) | ( ng105  &  wire31029 ) | ( (~ ng105)  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire3054 = ( (~ ng113)  &  wire30988 ) | ( (~ ng113)  &  wire30989 ) | ( ng113  &  (~ wire30988)  &  (~ wire30989) ) ;
 assign wire3065 = ( (~ ng97)  &  wire31048 ) | ( (~ ng97)  &  wire31049 ) | ( ng97  &  (~ wire31048)  &  (~ wire31049) ) ;
 assign wire3326 = ( (~ ng18079)  &  (~ ng18183) ) | ( (~ ng18346)  &  wire3054 ) ;
 assign wire3368 = ( (~ ng2257) ) | ( wire31077 ) | ( wire31078 ) ;
 assign ng23486 = ( wire31249 ) | ( wire31250 ) | ( wire31251 ) ;
 assign ng18319 = ( ng2170  &  wire33508 ) | ( ng2170  &  wire33509 ) | ( (~ ng2170)  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign ng18395 = ( (~ wire33428)  &  (~ wire33429)  &  wire33458 ) | ( (~ wire33428)  &  (~ wire33429)  &  wire33459 ) | ( wire33428  &  (~ wire33458)  &  (~ wire33459) ) | ( wire33429  &  (~ wire33458)  &  (~ wire33459) ) ;
 assign ng18478 = ( ng2195  &  wire33498 ) | ( ng2195  &  wire33499 ) | ( (~ ng2195)  &  (~ wire33498)  &  (~ wire33499) ) ;
 assign ng18578 = ( ng2175  &  wire33448 ) | ( ng2175  &  wire33449 ) | ( (~ ng2175)  &  (~ wire33448)  &  (~ wire33449) ) ;
 assign ng18606 = ( (~ wire33438)  &  (~ wire33439)  &  wire33630 ) | ( (~ wire33438)  &  (~ wire33439)  &  wire33631 ) | ( wire33438  &  (~ wire33630)  &  (~ wire33631) ) | ( wire33439  &  (~ wire33630)  &  (~ wire33631) ) ;
 assign ng18053 = ( ng2200  &  wire33478 ) | ( ng2200  &  wire33479 ) | ( (~ ng2200)  &  (~ wire33478)  &  (~ wire33479) ) ;
 assign ng18231 = ( ng2180  &  wire33488 ) | ( ng2180  &  wire33489 ) | ( (~ ng2180)  &  (~ wire33488)  &  (~ wire33489) ) ;
 assign wire3055 = ( (~ ng2165)  &  wire33560 ) | ( (~ ng2165)  &  wire33561 ) | ( ng2165  &  (~ wire33560)  &  (~ wire33561) ) ;
 assign wire3066 = ( (~ ng2190)  &  wire33468 ) | ( (~ ng2190)  &  wire33469 ) | ( ng2190  &  (~ wire33468)  &  (~ wire33469) ) ;
 assign wire3105 = ( (~ ng2185)  &  wire33518 ) | ( (~ ng2185)  &  wire33519 ) | ( ng2185  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire3369 = ( (~ ng2257) ) | ( wire33588 ) | ( wire33589 ) ;
 assign ng23537 = ( wire3369 ) | ( wire34428  &  wire34429  &  wire34430 ) ;
 assign ng22157 = ( pg3229  &  wire33998  &  wire35799 ) | ( pg3229  &  wire33999  &  wire35799 ) | ( (~ pg3229)  &  (~ wire33998)  &  (~ wire33999)  &  wire35799 ) ;
 assign ng10747 = ( (~ ng1312) ) | ( (~ ng2704) ) ;
 assign wire3370 = ( (~ ng2753) ) | ( (~ ng24043) ) ;
 assign ng24038 = ( (~ wire7190)  &  (~ wire7191)  &  (~ wire7192)  &  wire33944 ) ;
 assign ng27566 = ( (~ ng2257)  &  (~ ng11912)  &  (~ ng27567) ) | ( ng2257  &  ng11912  &  (~ ng25091) ) | ( ng2257  &  (~ ng11912)  &  (~ ng27567)  &  (~ ng25091) ) ;
 assign ng27576 = ( ng2257  &  (~ ng25099)  &  ng11962 ) | ( (~ ng2257)  &  (~ ng27577)  &  (~ ng11962) ) | ( ng2257  &  (~ ng25099)  &  (~ ng27577)  &  (~ ng11962) ) ;
 assign ng17031 = ( ng853  &  ng2257  &  wire31297  &  wire31298 ) ;
 assign wire3371 = ( (~ ng74) ) | ( (~ ng56) ) | ( (~ ng23497) ) | ( (~ wire35057) ) ;
 assign wire3372 = ( (~ ng2124) ) | ( (~ ng2142) ) | ( (~ ng23539) ) | ( (~ wire33829) ) ;
 assign ng24695 = ( wire32093 ) | ( (~ wire32088)  &  (~ wire32089)  &  wire32092 ) ;
 assign ng11663 = ( wire8834 ) | ( wire8835 ) | ( wire31793 ) | ( wire31795 ) ;
 assign ng28529 = ( ng25818 ) | ( wire32131 ) | ( ng27850  &  wire32130 ) ;
 assign ng12820 = ( wire31785 ) | ( wire31786 ) ;
 assign ng25958 = ( (~ ng11663) ) | ( (~ ng11600) ) | ( ng11647  &  (~ ng12941) ) | ( ng11663  &  ng11600  &  (~ ng11647)  &  ng12941 ) ;
 assign ng26327 = ( (~ ng25958)  &  (~ ng16655)  &  wire31785 ) | ( (~ ng25958)  &  (~ ng16655)  &  wire31786 ) | ( (~ ng25958)  &  ng16655  &  (~ wire31785)  &  (~ wire31786) ) ;
 assign ng12968 = ( wire3046 ) | ( wire8757 ) | ( wire31834 ) | ( wire31838 ) ;
 assign ng29677 = ( wire4961 ) | ( wire4964 ) | ( wire35780 ) | ( wire35781 ) ;
 assign ng30033 = ( (~ ng11678)  &  (~ ng24723)  &  wire4302 ) | ( (~ ng11678)  &  (~ ng24723)  &  wire36151 ) | ( ng11678  &  (~ ng24723)  &  (~ wire4302)  &  (~ wire36151) ) ;
 assign ng30015 = ( wire3361 ) | ( wire4319 ) | ( wire4320 ) | ( wire4321 ) ;
 assign ng30016 = ( wire4397 ) | ( wire36096 ) | ( wire36097 ) | ( wire36098 ) ;
 assign ng11600 = ( wire31805 ) | ( wire31806 ) ;
 assign ng11647 = ( wire3046 ) | ( wire8837 ) | ( wire31812 ) | ( wire31816 ) ;
 assign ng17086 = ( wire31815  &  wire32128 ) | ( wire31816  &  wire32128 ) ;
 assign ng24712 = ( wire7977 ) | ( wire7978 ) | ( wire7979 ) ;
 assign ng22399 = ( wire32897 ) | ( wire32898 ) | ( wire32903 ) | ( wire32904 ) ;
 assign ng24683 = ( (~ ng22399)  &  (~ wire32906)  &  (~ wire32907)  &  (~ wire32908) ) ;
 assign ng12876 = ( wire31360  &  wire31361 ) ;
 assign ng22381 = ( wire31231 ) | ( wire31232 ) ;
 assign ng17051 = ( wire30977  &  wire31271 ) | ( wire30978  &  wire31271 ) ;
 assign ng11644 = ( wire3046 ) | ( wire9437 ) | ( wire30954 ) | ( wire30958 ) ;
 assign ng13378 = ( wire3046 ) | ( wire9429 ) | ( wire30964 ) | ( wire30968 ) ;
 assign ng27834 = ( wire9265 ) | ( ng23486  &  ng23478  &  wire31270 ) ;
 assign ng11687 = ( wire33528 ) | ( wire33529 ) ;
 assign ng17151 = ( wire33548  &  wire33792 ) | ( wire33549  &  wire33792 ) ;
 assign ng22400 = ( wire33674 ) | ( wire33675 ) | ( wire33751 ) | ( wire33752 ) ;
 assign ng11653 = ( wire3046 ) | ( wire7504 ) | ( wire33535 ) | ( wire33539 ) ;
 assign ng27892 = ( wire7336 ) | ( ng23533  &  ng23521  &  wire33791 ) ;
 assign ng11955 = ( wire3049 ) | ( wire5104 ) | ( wire35574 ) | ( wire35578 ) ;
 assign ng29713 = ( ng11955  &  ng12292  &  wire3074 ) | ( ng12292  &  (~ ng21770)  &  wire3074 ) | ( (~ ng11955)  &  (~ ng12292)  &  ng21770  &  wire3074 ) ;
 assign ng11330 = ( (~ ng2935)  &  ng2941  &  ng2938  &  ng2944 ) | ( ng2935  &  (~ ng2941)  &  ng2938  &  ng2944 ) | ( ng2935  &  ng2941  &  (~ ng2938)  &  ng2944 ) | ( (~ ng2935)  &  (~ ng2941)  &  (~ ng2938)  &  ng2944 ) | ( ng2935  &  ng2941  &  ng2938  &  (~ ng2944) ) | ( (~ ng2935)  &  (~ ng2941)  &  ng2938  &  (~ ng2944) ) | ( (~ ng2935)  &  ng2941  &  (~ ng2938)  &  (~ ng2944) ) | ( ng2935  &  (~ ng2941)  &  (~ ng2938)  &  (~ ng2944) ) ;
 assign ng12250 = ( wire6366 ) | ( wire6367 ) | ( wire34813 ) | ( wire34815 ) ;
 assign ng27824 = ( ng12288  &  ng12250  &  wire3076 ) | ( ng12288  &  (~ ng21746)  &  wire3076 ) | ( (~ ng12288)  &  (~ ng12250)  &  ng21746  &  wire3076 ) ;
 assign ng30622 = ( wire35752 ) | ( wire3341  &  (~ wire34532)  &  (~ wire34533) ) ;
 assign ng30926 = ( (~ ng30622)  &  ng30610  &  ng30614  &  ng30629 ) | ( ng30622  &  (~ ng30610)  &  ng30614  &  ng30629 ) | ( ng30622  &  ng30610  &  (~ ng30614)  &  ng30629 ) | ( (~ ng30622)  &  (~ ng30610)  &  (~ ng30614)  &  ng30629 ) | ( ng30622  &  ng30610  &  ng30614  &  (~ ng30629) ) | ( (~ ng30622)  &  (~ ng30610)  &  ng30614  &  (~ ng30629) ) | ( (~ ng30622)  &  ng30610  &  (~ ng30614)  &  (~ ng30629) ) | ( ng30622  &  (~ ng30610)  &  (~ ng30614)  &  (~ ng30629) ) ;
 assign ng21711 = ( ng21796 ) | ( wire4250 ) | ( wire36175 ) ;
 assign ng21796 = ( (~ pg3234)  &  (~ wire35758) ) | ( (~ pg3234)  &  (~ wire35759) ) ;
 assign ng10706 = ( (~ ng1312) ) | ( (~ ng1316) ) ;
 assign ng10238 = ( ng1312  &  ng2010 ) ;
 assign ng17124 = ( wire32650  &  wire32944 ) | ( wire32651  &  wire32944 ) ;
 assign ng11678 = ( wire3046 ) | ( wire7512 ) | ( wire33545 ) | ( wire33549 ) ;
 assign ng10677 = ( (~ ng1312) ) | ( (~ ng630) ) ;
 assign ng11952 = ( wire33018 ) | ( wire33019 ) ;
 assign ng12005 = ( wire3046 ) | ( wire7246 ) | ( wire33868 ) | ( wire33872 ) ;
 assign ng11733 = ( (~ ng1315) ) | ( (~ ng2599) ) | ( (~ ng2612) ) | ( ng2733 ) ;
 assign ng13146 = ( (~ ng1309) ) | ( (~ ng2599) ) | ( (~ ng2612) ) | ( ng2733 ) ;
 assign ng13113 = ( (~ ng1312) ) | ( ng659 ) | ( (~ ng525) ) | ( (~ ng538) ) ;
 assign ng13137 = ( (~ ng1312) ) | ( (~ ng1905) ) | ( ng2039 ) | ( (~ ng1918) ) ;
 assign ng17973 = ( (~ pg3233) ) | ( pg3230 ) ;
 assign ng12945 = ( wire33023  &  wire33024 ) ;
 assign wire3046 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853) ) ;
 assign ng18218 = ( wire7863 ) | ( wire7864 ) | ( wire33083 ) | ( wire33084 ) ;
 assign ng11624 = ( wire3046 ) | ( wire9445 ) | ( wire30974 ) | ( wire30978 ) ;
 assign ng13142 = ( (~ ng1309) ) | ( (~ ng1905) ) | ( ng2039 ) | ( (~ ng1918) ) ;
 assign ng11800 = ( wire3046 ) | ( wire9416 ) | ( wire31156 ) | ( wire31160 ) ;
 assign ng12352 = ( wire3049 ) | ( wire7170 ) | ( wire33954 ) | ( wire33958 ) ;
 assign ng12195 = ( wire31723 ) | ( wire31724 ) ;
 assign ng12991 = ( wire3046 ) | ( wire8853 ) | ( wire31844 ) | ( wire31848 ) ;
 assign ng12107 = ( wire33008 ) | ( wire33009 ) ;
 assign ng12941 = ( wire3046 ) | ( wire8797 ) | ( wire31823 ) | ( wire31827 ) ;
 assign ng11902 = ( wire32219 ) | ( wire32220 ) ;
 assign ng26126 = ( wire34619 ) | ( wire3339  &  (~ wire31699)  &  (~ wire31700) ) ;
 assign wire3252 = ( (~ ng1315) ) | ( ng659 ) ;
 assign wire3204 = ( (~ ng1309) ) | ( (~ ng1316) ) ;
 assign ng12245 = ( wire31449 ) | ( wire31450 ) ;
 assign wire3205 = ( (~ ng1315) ) | ( (~ ng630) ) ;
 assign ng12249 = ( wire3049 ) | ( wire8441 ) | ( wire32289 ) | ( wire32293 ) ;
 assign wire3206 = ( (~ ng1309) ) | ( (~ ng2704) ) ;
 assign ng12292 = ( wire3049 ) | ( wire7787 ) | ( wire33164 ) | ( wire33168 ) ;
 assign ng13126 = ( (~ ng1211) ) | ( (~ ng1312) ) | ( (~ ng1224) ) | ( ng1345 ) ;
 assign ng11875 = ( wire32816 ) | ( wire32817 ) ;
 assign wire3296 = ( (~ ng2033) ) | ( (~ ng2026) ) | ( (~ ng2020) ) | ( (~ wire33414) ) ;
 assign ng24009 = ( ng2026  &  wire33413  &  wire33414  &  wire36465 ) ;
 assign wire3139 = ( pg8021 ) | ( wire35029  &  wire35030 ) ;
 assign wire3310 = ( (~ ng2950) ) | ( ng20825 ) ;
 assign wire3221 = ( ng1312  &  (~ wire31522) ) | ( ng1312  &  (~ wire31523) ) | ( ng1312  &  (~ wire31524) ) ;
 assign ng27551 = ( wire6114 ) | ( wire3197  &  (~ wire32243)  &  (~ wire32244) ) ;
 assign ng11870 = ( wire3046 ) | ( wire8510 ) | ( wire32206 ) | ( wire32210 ) ;
 assign wire3197 = ( ng2257  &  (~ ng25082)  &  (~ wire32209)  &  (~ wire32210) ) ;
 assign ng27550 = ( (~ ng2257)  &  (~ ng27551)  &  (~ ng11870) ) | ( ng2257  &  ng11870  &  (~ ng25082) ) | ( ng2257  &  (~ ng27551)  &  (~ ng11870)  &  (~ ng25082) ) ;
 assign wire3374 = ( (~ ng2059) ) | ( (~ ng24009) ) ;
 assign ng12755 = ( wire3046 ) | ( wire8781 ) | ( wire31854 ) | ( wire31858 ) ;
 assign ng26915 = ( ng26925 ) | ( wire32142 ) ;
 assign ng11675 = ( wire32630 ) | ( wire32631 ) ;
 assign ng28501 = ( ng25764 ) | ( wire31274 ) | ( ng27834  &  wire31273 ) ;
 assign ng27563 = ( (~ ng16643)  &  ng12781  &  ng12939  &  (~ ng25954) ) | ( ng16643  &  (~ ng12781)  &  (~ ng12939)  &  (~ ng25954) ) ;
 assign wire3175 = ( wire31274 ) | ( ng27834  &  wire31273 ) ;
 assign wire3359 = ( ng11624  &  ng25764  &  (~ ng27738) ) | ( ng25764  &  (~ ng27738)  &  (~ wire30979) ) ;
 assign ng28556 = ( ng25853 ) | ( wire32947 ) | ( ng27875  &  wire32946 ) ;
 assign ng12971 = ( wire3046 ) | ( wire8231 ) | ( wire32587 ) | ( wire32591 ) ;
 assign wire3180 = ( wire32947 ) | ( ng27875  &  wire32946 ) ;
 assign wire3190 = ( (~ ng12828)  &  wire32650 ) | ( (~ ng12828)  &  wire32651 ) | ( (~ ng12828)  &  (~ wire32652) ) | ( ng12828  &  (~ wire32650)  &  (~ wire32651)  &  wire32652 ) ;
 assign wire3361 = ( (~ ng27751)  &  (~ ng16672)  &  wire8146 ) | ( (~ ng27751)  &  (~ ng16672)  &  wire8147 ) ;
 assign ng29680 = ( wire7954 ) | ( wire7955 ) | ( wire32962 ) | ( wire32963 ) ;
 assign ng29670 = ( wire5973 ) | ( wire5976 ) | ( wire35046 ) | ( wire35047 ) ;
 assign ng30030 = ( (~ ng11624)  &  (~ ng24676)  &  wire7026 ) | ( (~ ng11624)  &  (~ ng24676)  &  wire34100 ) | ( ng11624  &  (~ ng24676)  &  (~ wire7026)  &  (~ wire34100) ) ;
 assign ng30032 = ( (~ ng24712)  &  (~ ng11666)  &  wire5849 ) | ( (~ ng24712)  &  (~ ng11666)  &  wire35175 ) | ( (~ ng24712)  &  ng11666  &  (~ wire5849)  &  (~ wire35175) ) ;
 assign ng18419 = ( (~ wire30937)  &  (~ wire30938)  &  wire31201 ) | ( (~ wire30937)  &  (~ wire30938)  &  wire31202 ) | ( wire30937  &  (~ wire31201)  &  (~ wire31202) ) | ( wire30938  &  (~ wire31201)  &  (~ wire31202) ) ;
 assign ng17887 = ( ng109  &  wire30927 ) | ( ng109  &  wire30928 ) | ( (~ ng109)  &  (~ wire30927)  &  (~ wire30928) ) ;
 assign ng17807 = ( ng117  &  wire30998 ) | ( ng117  &  wire30999 ) | ( (~ ng117)  &  (~ wire30998)  &  (~ wire30999) ) ;
 assign ng17729 = ( ng125  &  wire31008 ) | ( ng125  &  wire31009 ) | ( (~ ng125)  &  (~ wire31008)  &  (~ wire31009) ) ;
 assign wire3106 = ( (~ ng101)  &  wire31018 ) | ( (~ ng101)  &  wire31019 ) | ( ng101  &  (~ wire31018)  &  (~ wire31019) ) ;
 assign wire3284 = ( (~ ng17887)  &  (~ ng17807) ) | ( (~ ng18419)  &  (~ ng17729) ) ;
 assign ng23478 = ( wire31265 ) | ( wire31266 ) | ( wire31267 ) ;
 assign ng22396 = ( wire32088 ) | ( wire32089 ) ;
 assign ng12916 = ( wire32224  &  wire32225 ) ;
 assign ng11621 = ( (~ pg8271)  &  pg8270  &  pg8269  &  pg8268 ) | ( pg8271  &  (~ pg8270)  &  pg8269  &  pg8268 ) | ( pg8271  &  pg8270  &  (~ pg8269)  &  pg8268 ) | ( (~ pg8271)  &  (~ pg8270)  &  (~ pg8269)  &  pg8268 ) | ( pg8271  &  pg8270  &  pg8269  &  (~ pg8268) ) | ( (~ pg8271)  &  (~ pg8270)  &  pg8269  &  (~ pg8268) ) | ( (~ pg8271)  &  pg8270  &  (~ pg8269)  &  (~ pg8268) ) | ( pg8271  &  (~ pg8270)  &  (~ pg8269)  &  (~ pg8268) ) ;
 assign ng26145 = ( wire35023 ) | ( wire3339  &  (~ wire31711)  &  (~ wire31712) ) ;
 assign ng26151 = ( wire34962 ) | ( wire3336  &  (~ wire31605)  &  (~ wire31606) ) ;
 assign ng11873 = ( wire3049 ) | ( wire6377 ) | ( wire34836 ) | ( wire34840 ) ;
 assign ng27811 = ( ng12249  &  ng11873  &  wire3076 ) | ( ng12249  &  (~ ng21746)  &  wire3076 ) | ( (~ ng12249)  &  (~ ng11873)  &  ng21746  &  wire3076 ) ;
 assign ng29728 = ( ng12292  &  ng12263  &  wire3074 ) | ( ng12292  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12292)  &  (~ ng12263)  &  ng21770  &  wire3074 ) ;
 assign ng30034 = ( (~ ng29728)  &  ng29741  &  ng29732  &  ng29748 ) | ( ng29728  &  (~ ng29741)  &  ng29732  &  ng29748 ) | ( ng29728  &  ng29741  &  (~ ng29732)  &  ng29748 ) | ( (~ ng29728)  &  (~ ng29741)  &  (~ ng29732)  &  ng29748 ) | ( ng29728  &  ng29741  &  ng29732  &  (~ ng29748) ) | ( (~ ng29728)  &  (~ ng29741)  &  ng29732  &  (~ ng29748) ) | ( (~ ng29728)  &  ng29741  &  (~ ng29732)  &  (~ ng29748) ) | ( ng29728  &  (~ ng29741)  &  (~ ng29732)  &  (~ ng29748) ) ;
 assign ng11781 = ( wire3046 ) | ( wire9400 ) | ( wire31198 ) | ( wire31202 ) ;
 assign ng12970 = ( wire3046 ) | ( wire8239 ) | ( wire32709 ) | ( wire32713 ) ;
 assign ng18561 = ( ng1471  &  wire32712 ) | ( ng1471  &  wire32713 ) | ( (~ ng1471)  &  (~ wire32712)  &  (~ wire32713) ) ;
 assign ng25853 = ( wire8147 ) | ( ng25964  &  wire32721  &  wire32722 ) ;
 assign ng27751 = ( wire32947 ) | ( ng27875  &  wire32946 ) ;
 assign ng11860 = ( wire9183 ) | ( wire9184 ) | ( wire31353 ) | ( wire31355 ) ;
 assign ng12121 = ( wire3046 ) | ( wire7196 ) | ( wire33913 ) | ( wire33917 ) ;
 assign ng17197 = ( ng2892  &  ng853 ) | ( ng2903  &  ng853 ) | ( ng853  &  (~ wire31298) ) ;
 assign ng23539 = ( ng853  &  (~ wire31297)  &  wire33827 ) | ( ng853  &  (~ wire31298)  &  wire33827 ) ;
 assign ng18363 = ( ng801  &  wire31847 ) | ( ng801  &  wire31848 ) | ( (~ ng801)  &  (~ wire31847)  &  (~ wire31848) ) ;
 assign ng18441 = ( ng793  &  wire31837 ) | ( ng793  &  wire31838 ) | ( (~ ng793)  &  (~ wire31837)  &  (~ wire31838) ) ;
 assign ng18195 = ( (~ wire31770)  &  (~ wire31771)  &  wire31907 ) | ( (~ wire31770)  &  (~ wire31771)  &  wire31908 ) | ( wire31770  &  (~ wire31907)  &  (~ wire31908) ) | ( wire31771  &  (~ wire31907)  &  (~ wire31908) ) ;
 assign ng18290 = ( ng809  &  wire31857 ) | ( ng809  &  wire31858 ) | ( (~ ng809)  &  (~ wire31857)  &  (~ wire31858) ) ;
 assign wire3067 = ( (~ ng785)  &  wire31826 ) | ( (~ ng785)  &  wire31827 ) | ( ng785  &  (~ wire31826)  &  (~ wire31827) ) ;
 assign wire3285 = ( (~ ng18363)  &  (~ ng18441) ) | ( (~ ng18195)  &  (~ ng18290) ) ;
 assign wire3375 = ( (~ ng2257) ) | ( wire31934 ) | ( wire31935 ) ;
 assign ng23502 = ( wire32106 ) | ( wire32107 ) | ( wire32108 ) ;
 assign wire3286 = ( ng159 ) | ( (~ ng853) ) ;
 assign wire3287 = ( (~ ng826) ) | ( ng151 ) ;
 assign wire3333 = ( (~ ng3080) ) | ( (~ ng2998) ) | ( (~ ng2993) ) ;
 assign ng13145 = ( (~ ng1312) ) | ( (~ ng2599) ) | ( (~ ng2612) ) | ( ng2733 ) ;
 assign ng11721 = ( (~ ng1315) ) | ( ng659 ) | ( (~ ng525) ) | ( (~ ng538) ) ;
 assign wire3246 = ( ng3139 ) | ( (~ ng3147) ) ;
 assign wire3247 = ( (~ ng3135) ) | ( ng3120 ) ;
 assign wire3248 = ( (~ ng1315) ) | ( ng2733 ) ;
 assign ng12145 = ( wire9078 ) | ( wire9079 ) | ( wire31500 ) | ( wire31502 ) ;
 assign ng13001 = ( wire3046 ) | ( wire8247 ) | ( wire32597 ) | ( wire32601 ) ;
 assign ng12100 = ( wire6414 ) | ( wire6415 ) | ( wire34755 ) | ( wire34757 ) ;
 assign ng12044 = ( wire3046 ) | ( wire8469 ) | ( wire32259 ) | ( wire32263 ) ;
 assign ng12698 = ( wire3046 ) | ( wire9525 ) | ( wire30944 ) | ( wire30948 ) ;
 assign ng10793 = ( wire3049 ) | ( wire8368 ) | ( wire32396 ) | ( wire32400 ) ;
 assign ng11915 = ( wire5165 ) | ( wire5166 ) | ( wire35585 ) | ( wire35587 ) ;
 assign ng11726 = ( (~ ng1211) ) | ( (~ ng1315) ) | ( (~ ng1224) ) | ( ng1345 ) ;
 assign ng11833 = ( wire3046 ) | ( wire8865 ) | ( wire31767 ) | ( wire31771 ) ;
 assign ng23495 = ( wire3368 ) | ( wire31426  &  wire31427  &  wire31428 ) ;
 assign wire3377 = ( (~ ng1365) ) | ( (~ ng23979) ) ;
 assign ng16655 = ( (~ wire31815)  &  (~ wire31816)  &  wire31817 ) ;
 assign wire3748 = ( (~ ng12941) ) | ( (~ wire31828) ) | ( (~ wire31815)  &  (~ wire31816) ) ;
 assign ng26374 = ( ng11666  &  ng12858  &  (~ ng25964) ) | ( ng12858  &  (~ ng25964)  &  (~ wire32652) ) | ( (~ ng11666)  &  (~ ng12858)  &  (~ ng25964)  &  wire32652 ) ;
 assign ng12992 = ( wire3046 ) | ( wire8207 ) | ( wire32607 ) | ( wire32611 ) ;
 assign ng29672 = ( wire8566 ) | ( wire8569 ) | ( wire32150 ) | ( wire32151 ) ;
 assign ng30021 = ( wire3359 ) | ( wire5963 ) | ( wire5964 ) | ( wire5965 ) ;
 assign ng11630 = ( wire3046 ) | ( wire8159 ) | ( wire32637 ) | ( wire32641 ) ;
 assign ng11666 = ( wire3046 ) | ( wire8151 ) | ( wire32647 ) | ( wire32651 ) ;
 assign ng12248 = ( wire32303 ) | ( wire32304 ) ;
 assign ng12097 = ( wire8419 ) | ( wire8420 ) | ( wire32321 ) | ( wire32323 ) ;
 assign ng10814 = ( wire8365 ) | ( wire8366 ) | ( wire32407 ) | ( wire32409 ) ;
 assign ng12152 = ( wire32313 ) | ( wire32314 ) ;
 assign ng10801 = ( wire3049 ) | ( wire8344 ) | ( wire32416 ) | ( wire32420 ) ;
 assign wire3288 = ( wire32429 ) | ( wire32430 ) | ( (~ wire32419)  &  (~ wire32420) ) ;
 assign ng23071 = ( wire8329 ) | ( wire8330 ) | ( wire32560 ) | ( wire32561 ) ;
 assign ng12974 = ( wire33876  &  wire33877 ) ;
 assign ng27875 = ( wire7981 ) | ( ng23518  &  ng23505  &  wire32943 ) ;
 assign ng12999 = ( (~ pg8263)  &  pg8261  &  pg8260  &  pg8259 ) | ( pg8263  &  (~ pg8261)  &  pg8260  &  pg8259 ) | ( pg8263  &  pg8261  &  (~ pg8260)  &  pg8259 ) | ( (~ pg8263)  &  (~ pg8261)  &  (~ pg8260)  &  pg8259 ) | ( pg8263  &  pg8261  &  pg8260  &  (~ pg8259) ) | ( (~ pg8263)  &  (~ pg8261)  &  pg8260  &  (~ pg8259) ) | ( (~ pg8263)  &  pg8261  &  (~ pg8260)  &  (~ pg8259) ) | ( pg8263  &  (~ pg8261)  &  (~ pg8260)  &  (~ pg8259) ) ;
 assign ng25099 = ( ng12005  &  ng11917 ) | ( ng12005  &  wire3925 ) | ( ng12005  &  wire33878 ) | ( (~ ng12005)  &  (~ ng11917)  &  (~ wire33878) ) ;
 assign wire3194 = ( ng2257  &  (~ ng25099)  &  (~ wire33889)  &  (~ wire33890) ) ;
 assign ng27577 = ( wire7225 ) | ( wire3194  &  (~ wire33906)  &  (~ wire33907) ) ;
 assign ng21746 = ( wire35840 ) | ( wire35841 ) | ( wire35845 ) ;
 assign ng25874 = ( wire7500 ) | ( ng25969  &  wire33569  &  wire33570 ) ;
 assign ng27756 = ( ng24723 ) | ( wire7327 ) | ( ng27892  &  wire33794 ) ;
 assign ng23349 = ( wire3122  &  ng12213  &  wire33008 ) | ( wire3122  &  ng12213  &  wire33009 ) | ( (~ wire3122)  &  (~ wire33008)  &  (~ wire33009) ) ;
 assign ng12920 = ( wire3046 ) | ( wire8813 ) | ( wire31874 ) | ( wire31878 ) ;
 assign ng12890 = ( wire31887 ) | ( wire31888 ) ;
 assign ng12852 = ( wire31897 ) | ( wire31898 ) ;
 assign ng12789 = ( wire3046 ) | ( wire8765 ) | ( wire31904 ) | ( wire31908 ) ;
 assign ng25818 = ( wire8754 ) | ( ng25958  &  wire31915  &  wire31916 ) ;
 assign wire3210 = ( (~ ng1309) ) | ( (~ ng630) ) ;
 assign ng12216 = ( wire35597 ) | ( wire35598 ) ;
 assign ng8430 = ( ng3110  &  (~ ng3124)  &  (~ ng3126)  &  (~ ng3191) ) ;
 assign ng11889 = ( wire3046 ) | ( wire9384 ) | ( wire31122 ) | ( wire31126 ) ;
 assign ng11975 = ( wire3046 ) | ( wire9134 ) | ( wire31391 ) | ( wire31395 ) ;
 assign ng11882 = ( wire3046 ) | ( wire7467 ) | ( wire33627 ) | ( wire33631 ) ;
 assign wire3304 = ( (~ ng2727) ) | ( (~ ng2720) ) | ( (~ ng2707) ) | ( (~ wire34450) ) ;
 assign ng24043 = ( ng2720  &  wire34449  &  wire34450  &  wire35557 ) ;
 assign ng23335 = ( wire5442 ) | ( wire5443 ) | ( wire35350 ) ;
 assign ng11828 = ( wire31345 ) | ( wire31346 ) ;
 assign ng27529 = ( wire9165 ) | ( wire3195  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign ng25078 = ( ng11781  &  ng11860 ) | ( ng11860  &  wire3936 ) | ( ng11860  &  wire31362 ) | ( (~ ng11781)  &  (~ ng11860)  &  (~ wire31362) ) ;
 assign wire3353 = ( (~ ng25078)  &  wire31345 ) | ( (~ ng25078)  &  wire31346 ) ;
 assign ng27528 = ( (~ ng2257)  &  (~ ng11828)  &  ng25078 ) | ( ng2257  &  ng11828  &  (~ ng25078) ) | ( ng11828  &  ng27529  &  (~ ng25078) ) | ( (~ ng11828)  &  (~ ng27529)  &  (~ ng25078) ) ;
 assign wire3380 = ( (~ ng679) ) | ( (~ ng23950) ) ;
 assign ng12949 = ( wire3046 ) | ( wire8223 ) | ( wire32617 ) | ( wire32621 ) ;
 assign ng16672 = ( (~ wire32650)  &  (~ wire32651)  &  wire32652 ) ;
 assign ng12930 = ( wire3046 ) | ( wire8215 ) | ( wire32658 ) | ( wire32662 ) ;
 assign ng12797 = ( wire3046 ) | ( wire8191 ) | ( wire32678 ) | ( wire32682 ) ;
 assign ng12858 = ( wire3046 ) | ( wire8183 ) | ( wire32688 ) | ( wire32692 ) ;
 assign ng12828 = ( wire3046 ) | ( wire8175 ) | ( wire32698 ) | ( wire32702 ) ;
 assign ng25964 = ( (~ ng11675) ) | ( (~ ng11630) ) | ( (~ ng12970)  &  ng11666 ) | ( ng11675  &  ng12970  &  ng11630  &  (~ ng11666) ) ;
 assign wire3234 = ( wire32945 ) | ( (~ ng1704)  &  ng823 ) ;
 assign wire3935 = ( ng2257  &  wire32740 ) | ( ng2257  &  wire32741 ) ;
 assign ng24676 = ( wire31236 ) | ( (~ wire31231)  &  (~ wire31232)  &  wire31235 ) ;
 assign ng29912 = ( ng11644  &  (~ ng24676)  &  wire9118 ) | ( ng11644  &  (~ ng24676)  &  wire31438 ) | ( (~ ng11644)  &  (~ ng24676)  &  (~ wire9118)  &  (~ wire31438) ) ;
 assign ng28584 = ( ng25874 ) | ( wire33795 ) | ( ng27892  &  wire33794 ) ;
 assign wire3426 = ( ng26931 ) | ( (~ ng12866)  &  ng11678 ) | ( (~ ng12866)  &  (~ wire33550) ) | ( ng12866  &  (~ ng11678)  &  wire33550 ) ;
 assign ng29671 = ( wire9238 ) | ( wire9239 ) | ( wire31292 ) | ( wire31293 ) ;
 assign ng12207 = ( wire32429 ) | ( wire32430 ) ;
 assign ng23107 = ( wire8318 ) | ( wire32465 ) | ( wire32470 ) | ( wire32471 ) ;
 assign ng18598 = ( wire3049 ) | ( wire32529 ) | ( wire32535 ) | ( wire32536 ) ;
 assign ng24723 = ( (~ ng22400)  &  wire33754 ) | ( (~ ng22400)  &  wire33755 ) | ( (~ ng22400)  &  wire33756 ) ;
 assign ng24700 = ( (~ ng22400)  &  (~ wire33754)  &  (~ wire33755)  &  (~ wire33756) ) ;
 assign ng11946 = ( wire3049 ) | ( wire6353 ) | ( wire34800 ) | ( wire34804 ) ;
 assign ng27802 = ( ng12288  &  (~ ng21746)  &  wire3076 ) | ( ng12288  &  ng11946  &  wire3076 ) | ( (~ ng12288)  &  ng21746  &  (~ ng11946)  &  wire3076 ) ;
 assign ng17942 = ( ng1506  &  wire32620 ) | ( ng1506  &  wire32621 ) | ( (~ ng1506)  &  (~ wire32620)  &  (~ wire32621) ) ;
 assign wire3196 = ( ng2257  &  (~ ng25091)  &  (~ wire33036)  &  (~ wire33037) ) ;
 assign ng11263 = ( (~ ng2947)  &  ng2956  &  ng2953  &  ng2959 ) | ( ng2947  &  (~ ng2956)  &  ng2953  &  ng2959 ) | ( ng2947  &  ng2956  &  (~ ng2953)  &  ng2959 ) | ( (~ ng2947)  &  (~ ng2956)  &  (~ ng2953)  &  ng2959 ) | ( ng2947  &  ng2956  &  ng2953  &  (~ ng2959) ) | ( (~ ng2947)  &  (~ ng2956)  &  ng2953  &  (~ ng2959) ) | ( (~ ng2947)  &  ng2956  &  (~ ng2953)  &  (~ ng2959) ) | ( ng2947  &  (~ ng2956)  &  (~ ng2953)  &  (~ ng2959) ) ;
 assign ng27883 = ( ng12249  &  (~ ng21746)  &  wire3076 ) | ( ng12249  &  ng12099  &  wire3076 ) | ( (~ ng12249)  &  ng21746  &  (~ ng12099)  &  wire3076 ) ;
 assign ng28842 = ( (~ ng27883)  &  ng27855  &  ng27897  &  ng27865 ) | ( ng27883  &  (~ ng27855)  &  ng27897  &  ng27865 ) | ( ng27883  &  ng27855  &  (~ ng27897)  &  ng27865 ) | ( (~ ng27883)  &  (~ ng27855)  &  (~ ng27897)  &  ng27865 ) | ( ng27883  &  ng27855  &  ng27897  &  (~ ng27865) ) | ( (~ ng27883)  &  (~ ng27855)  &  ng27897  &  (~ ng27865) ) | ( (~ ng27883)  &  ng27855  &  (~ ng27897)  &  (~ ng27865) ) | ( ng27883  &  (~ ng27855)  &  (~ ng27897)  &  (~ ng27865) ) ;
 assign ng23377 = ( (~ ng12152)  &  wire3123 ) | ( ng12152  &  (~ wire3123)  &  wire32303 ) | ( ng12152  &  (~ wire3123)  &  wire32304 ) ;
 assign ng23368 = ( (~ ng12080)  &  wire3118 ) | ( ng12080  &  (~ wire3118)  &  wire31482 ) | ( ng12080  &  (~ wire3118)  &  wire31483 ) ;
 assign wire3327 = ( (~ ng18395)  &  (~ ng18578) ) | ( (~ ng18478)  &  wire3055 ) ;
 assign ng23533 = ( wire33770 ) | ( wire33771 ) | ( wire33772 ) ;
 assign ng18096 = ( ng789  &  wire31785 ) | ( ng789  &  wire31786 ) | ( (~ ng789)  &  (~ wire31785)  &  (~ wire31786) ) ;
 assign ng17998 = ( ng797  &  wire31897 ) | ( ng797  &  wire31898 ) | ( (~ ng797)  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign ng18492 = ( (~ wire31867)  &  (~ wire31868)  &  wire32020 ) | ( (~ wire31867)  &  (~ wire31868)  &  wire32021 ) | ( wire31867  &  (~ wire32020)  &  (~ wire32021) ) | ( wire31868  &  (~ wire32020)  &  (~ wire32021) ) ;
 assign wire3056 = ( (~ ng813)  &  wire31877 ) | ( (~ ng813)  &  wire31878 ) | ( ng813  &  (~ wire31877)  &  (~ wire31878) ) ;
 assign wire3107 = ( (~ ng805)  &  wire31887 ) | ( (~ ng805)  &  wire31888 ) | ( ng805  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign ng23511 = ( wire3375 ) | ( wire34289  &  wire34290  &  wire34291 ) ;
 assign ng12194 = ( wire31469 ) | ( wire31470 ) ;
 assign ng12172 = ( wire35607 ) | ( wire35608 ) ;
 assign ng12112 = ( wire3049 ) | ( wire5136 ) | ( wire35614 ) | ( wire35618 ) ;
 assign ng12035 = ( wire3049 ) | ( wire8979 ) | ( wire31708 ) | ( wire31712 ) ;
 assign ng26087 = ( wire35277 ) | ( wire3336  &  (~ wire31687)  &  (~ wire31688) ) ;
 assign wire3944 = ( ng21851  &  ng17139 ) | ( ng17139  &  wire34028 ) ;
 assign wire3253 = ( (~ ng1315) ) | ( ng1345 ) ;
 assign ng12060 = ( wire35627 ) | ( wire35628 ) ;
 assign ng12293 = ( wire3049 ) | ( wire5120 ) | ( wire35634 ) | ( wire35638 ) ;
 assign ng11999 = ( wire5117 ) | ( wire5118 ) | ( wire35645 ) | ( wire35647 ) ;
 assign ng12263 = ( wire5173 ) | ( wire5174 ) | ( wire35655 ) | ( wire35657 ) ;
 assign ng12171 = ( wire3049 ) | ( wire5096 ) | ( wire35664 ) | ( wire35668 ) ;
 assign ng11914 = ( wire3049 ) | ( wire5088 ) | ( wire35674 ) | ( wire35678 ) ;
 assign ng21770 = ( wire35694 ) | ( wire35695 ) | ( wire35699 ) ;
 assign ng12169 = ( wire7812 ) | ( wire7813 ) | ( wire33135 ) | ( wire33137 ) ;
 assign ng10851 = ( wire33353 ) | ( wire33354 ) ;
 assign ng12291 = ( wire7665 ) | ( wire7666 ) | ( wire33336 ) | ( wire33338 ) ;
 assign ng12214 = ( wire3049 ) | ( wire7797 ) | ( wire33124 ) | ( wire33128 ) ;
 assign wire3233 = ( wire33127 ) | ( wire33128 ) | ( (~ wire33117)  &  (~ wire33118) ) ;
 assign wire3354 = ( wire33137  &  (~ wire33328)  &  (~ wire33329) ) | ( wire33138  &  (~ wire33328)  &  (~ wire33329) ) ;
 assign wire3364 = ( (~ wire33137)  &  (~ wire33138)  &  wire33328 ) | ( (~ wire33137)  &  (~ wire33138)  &  wire33329 ) ;
 assign wire3437 = ( (~ wire33308)  &  (~ wire33309)  &  (~ wire33318)  &  (~ wire33319) ) ;
 assign wire3440 = ( wire33117  &  wire33127 ) | ( wire33118  &  wire33127 ) | ( wire33117  &  wire33128 ) | ( wire33118  &  wire33128 ) ;
 assign ng23340 = ( (~ ng12043)  &  wire3117 ) | ( ng12043  &  (~ wire3117)  &  wire36109 ) | ( ng12043  &  (~ wire3117)  &  wire36110 ) ;
 assign wire3530 = ( (~ ng853) ) | ( (~ wire34737)  &  (~ wire34738)  &  (~ wire34741) ) ;
 assign ng26869 = ( ng74  &  ng23497  &  wire35057 ) ;
 assign ng11917 = ( wire3046 ) | ( wire7612 ) | ( wire33425 ) | ( wire33429 ) ;
 assign ng26931 = ( (~ ng27585) ) | ( wire33805 ) | ( wire33807 ) | ( wire33819 ) ;
 assign ng29681 = ( wire7307 ) | ( wire7308 ) | ( wire33814 ) | ( wire33815 ) ;
 assign ng29920 = ( ng11687  &  (~ ng24723)  &  wire6720 ) | ( ng11687  &  (~ ng24723)  &  wire34440 ) | ( (~ ng11687)  &  (~ ng24723)  &  (~ wire6720)  &  (~ wire34440) ) ;
 assign ng12033 = ( wire3049 ) | ( wire9057 ) | ( wire31489 ) | ( wire31493 ) ;
 assign ng10789 = ( wire34176 ) | ( wire34177 ) ;
 assign ng12080 = ( wire3049 ) | ( wire9049 ) | ( wire31509 ) | ( wire31513 ) ;
 assign ng10784 = ( wire6955 ) | ( wire6956 ) | ( wire34194 ) | ( wire34196 ) ;
 assign wire3344 = ( wire31492  &  (~ wire34196)  &  (~ wire34197) ) | ( wire31493  &  (~ wire34196)  &  (~ wire34197) ) ;
 assign wire3345 = ( (~ wire31492)  &  (~ wire31493)  &  wire34196 ) | ( (~ wire31492)  &  (~ wire31493)  &  wire34197 ) ;
 assign wire3929 = ( wire31482  &  wire31512 ) | ( wire31483  &  wire31512 ) | ( wire31482  &  wire31513 ) | ( wire31483  &  wire31513 ) ;
 assign wire3949 = ( (~ wire34176)  &  (~ wire34177)  &  (~ wire34215)  &  (~ wire34216) ) ;
 assign ng18548 = ( wire9030 ) | ( wire31582 ) | ( wire31588 ) | ( wire31589 ) ;
 assign ng18639 = ( wire5224 ) | ( wire35510 ) | ( wire35516 ) | ( wire35517 ) ;
 assign wire3289 = ( (~ ng18319)  &  (~ ng18053) ) | ( (~ ng18606)  &  (~ ng18231) ) ;
 assign ng23521 = ( wire33786 ) | ( wire33787 ) | ( wire33788 ) ;
 assign ng29741 = ( ng12292  &  ng12171  &  wire3074 ) | ( ng12292  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12292)  &  (~ ng12171)  &  ng21770  &  wire3074 ) ;
 assign wire3183 = ( ng2574  &  (~ ng30072)  &  ng12328  &  (~ wire35748) ) ;
 assign wire3341 = ( (~ ng12328)  &  wire3075  &  wire35745 ) | ( (~ ng12328)  &  wire3075  &  wire35746 ) ;
 assign ng30594 = ( wire36172 ) | ( wire3341  &  (~ wire34496)  &  (~ wire34497) ) ;
 assign ng16643 = ( (~ wire30977)  &  (~ wire30978)  &  wire30979 ) ;
 assign ng22016 = ( pg3229  &  wire32998  &  wire35336 ) | ( pg3229  &  wire32999  &  wire35336 ) | ( (~ pg3229)  &  (~ wire32998)  &  (~ wire32999)  &  wire35336 ) ;
 assign ng21991 = ( pg3229  &  wire31324  &  wire34987 ) | ( pg3229  &  wire31325  &  wire34987 ) | ( (~ pg3229)  &  (~ wire31324)  &  (~ wire31325)  &  wire34987 ) ;
 assign ng16693 = ( (~ wire33548)  &  (~ wire33549)  &  wire33550 ) ;
 assign ng17985 = ( wire9155 ) | ( wire9156 ) | ( wire31414 ) | ( wire31415 ) ;
 assign ng12146 = ( wire31699 ) | ( wire31700 ) ;
 assign ng12967 = ( wire3046 ) | ( wire9501 ) | ( wire30985 ) | ( wire30989 ) ;
 assign ng12000 = ( wire3046 ) | ( wire7483 ) | ( wire33647 ) | ( wire33651 ) ;
 assign ng26154 = ( wire35309 ) | ( wire3339  &  (~ wire31651)  &  (~ wire31652) ) ;
 assign ng12849 = ( wire3046 ) | ( wire9493 ) | ( wire30995 ) | ( wire30999 ) ;
 assign ng11916 = ( wire3046 ) | ( wire7475 ) | ( wire33617 ) | ( wire33621 ) ;
 assign ng12880 = ( wire31008 ) | ( wire31009 ) ;
 assign ng12781 = ( wire3046 ) | ( wire9485 ) | ( wire31015 ) | ( wire31019 ) ;
 assign ng12939 = ( wire3046 ) | ( wire9469 ) | ( wire31025 ) | ( wire31029 ) ;
 assign ng12747 = ( wire3046 ) | ( wire9461 ) | ( wire31035 ) | ( wire31039 ) ;
 assign ng12912 = ( wire3046 ) | ( wire9453 ) | ( wire31045 ) | ( wire31049 ) ;
 assign ng12328 = ( wire3049 ) | ( wire7154 ) | ( wire33974 ) | ( wire33978 ) ;
 assign wire3328 = ( (~ ng17998)  &  (~ ng18492) ) | ( (~ ng18096)  &  wire3056 ) ;
 assign ng23489 = ( wire32122 ) | ( wire32123 ) | ( wire32124 ) ;
 assign wire3290 = ( (~ ng11644)  &  ng10711 ) | ( (~ ng13378)  &  ng10711 ) | ( (~ ng11624)  &  ng10711 ) | ( (~ ng11644)  &  ng13378  &  (~ ng11624) ) ;
 assign wire3220 = ( ng1309  &  (~ wire31522) ) | ( ng1309  &  (~ wire31523) ) | ( ng1309  &  (~ wire31524) ) ;
 assign ng24004 = ( (~ wire7844)  &  (~ wire7845)  &  (~ wire7846)  &  wire35285 ) ;
 assign ng27850 = ( wire8596 ) | ( ng23502  &  ng23489  &  wire32127 ) ;
 assign wire3235 = ( wire32129 ) | ( (~ ng1010)  &  ng823 ) ;
 assign wire3930 = ( ng2257  &  wire31934 ) | ( ng2257  &  wire31935 ) ;
 assign ng27743 = ( wire32131 ) | ( ng27850  &  wire32130 ) ;
 assign ng26878 = ( ng762  &  ng23513  &  wire32166 ) ;
 assign ng12043 = ( wire3046 ) | ( wire8540 ) | ( wire32174 ) | ( wire32178 ) ;
 assign wire3117 = ( pg3229  &  wire32187 ) | ( pg3229  &  wire32188 ) | ( (~ pg3229)  &  (~ wire32187)  &  (~ wire32188) ) ;
 assign ng29732 = ( ng12324  &  ng12216  &  wire3074 ) | ( ng12324  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12324)  &  (~ ng12216)  &  ng21770  &  wire3074 ) ;
 assign ng29705 = ( ng12324  &  ng11999  &  wire3074 ) | ( ng12324  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12324)  &  (~ ng11999)  &  ng21770  &  wire3074 ) ;
 assign ng29751 = ( ng12292  &  ng12060  &  wire3074 ) | ( ng12292  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12292)  &  (~ ng12060)  &  ng21770  &  wire3074 ) ;
 assign ng30035 = ( (~ ng29713)  &  ng29705  &  ng29751  &  ng29721 ) | ( ng29713  &  (~ ng29705)  &  ng29751  &  ng29721 ) | ( ng29713  &  ng29705  &  (~ ng29751)  &  ng29721 ) | ( (~ ng29713)  &  (~ ng29705)  &  (~ ng29751)  &  ng29721 ) | ( ng29713  &  ng29705  &  ng29751  &  (~ ng29721) ) | ( (~ ng29713)  &  (~ ng29705)  &  ng29751  &  (~ ng29721) ) | ( (~ ng29713)  &  ng29705  &  (~ ng29751)  &  (~ ng29721) ) | ( ng29713  &  (~ ng29705)  &  (~ ng29751)  &  (~ ng29721) ) ;
 assign ng25082 = ( ng11902  &  wire3930 ) | ( ng11902  &  ng11807 ) | ( ng11902  &  wire32226 ) | ( (~ ng11902)  &  (~ ng11807)  &  (~ wire32226) ) ;
 assign ng11962 = ( wire3046 ) | ( wire7235 ) | ( wire33886 ) | ( wire33890 ) ;
 assign ng23372 = ( pg3229  &  (~ ng12291) ) | ( (~ pg3229)  &  (~ wire3233) ) | ( (~ ng12169)  &  ng12291  &  wire3233 ) ;
 assign ng21976 = ( (~ ng12026)  &  wire3121 ) | ( ng12026  &  (~ wire31334)  &  (~ wire31335) ) ;
 assign ng27585 = ( (~ ng13002)  &  (~ ng12899)  &  ng16693  &  (~ ng25969) ) | ( ng13002  &  ng12899  &  (~ ng16693)  &  (~ ng25969) ) ;
 assign ng26947 = ( (~ ng27585) ) | ( (~ ng12933)  &  ng11678 ) | ( (~ ng12933)  &  (~ wire33550) ) | ( ng12933  &  (~ ng11678)  &  wire33550 ) ;
 assign wire3908 = ( ng2200  &  ng2185  &  (~ ng2190)  &  (~ ng2195) ) ;
 assign ng18458 = ( ng1491  &  wire32600 ) | ( ng1491  &  wire32601 ) | ( (~ ng1491)  &  (~ wire32600)  &  (~ wire32601) ) ;
 assign ng18514 = ( ng1481  &  wire32610 ) | ( ng1481  &  wire32611 ) | ( (~ ng1481)  &  (~ wire32610)  &  (~ wire32611) ) ;
 assign ng18383 = ( ng1501  &  wire32681 ) | ( ng1501  &  wire32682 ) | ( (~ ng1501)  &  (~ wire32681)  &  (~ wire32682) ) ;
 assign wire3068 = ( wire32701  &  wire32816 ) | ( wire32702  &  wire32816 ) | ( wire32701  &  wire32817 ) | ( wire32702  &  wire32817 ) | ( (~ wire32701)  &  (~ wire32702)  &  (~ wire32816)  &  (~ wire32817) ) ;
 assign wire3291 = ( (~ ng18561)  &  (~ ng18514) ) | ( (~ ng18458)  &  (~ ng18383) ) ;
 assign wire3386 = ( (~ ng2257) ) | ( wire32740 ) | ( wire32741 ) ;
 assign ng23518 = ( wire32922 ) | ( wire32923 ) | ( wire32924 ) ;
 assign wire3444 = ( ng510  &  wire31459 ) | ( ng510  &  wire31460 ) ;
 assign ng18325 = ( wire7209 ) | ( wire7210 ) | ( wire33926 ) | ( wire33927 ) ;
 assign ng15830 = ( ng3135 ) | ( ng3120 ) | ( wire3193 ) | ( (~ ng8430) ) ;
 assign wire3259 = ( (~ ng1315) ) | ( ng2039 ) ;
 assign ng12208 = ( wire6406 ) | ( wire6407 ) | ( wire34873 ) | ( wire34875 ) ;
 assign ng11784 = ( wire3046 ) | ( wire8729 ) | ( wire31963 ) | ( wire31967 ) ;
 assign ng11896 = ( wire3049 ) | ( wire8963 ) | ( wire31684 ) | ( wire31688 ) ;
 assign ng12162 = ( wire3046 ) | ( wire7922 ) | ( wire32985 ) | ( wire32989 ) ;
 assign wire3292 = ( (~ ng13004) ) | ( (~ ng3018)  &  ng13004 ) | ( pg3234  &  (~ wire36176) ) | ( ng13004  &  (~ wire36176) ) ;
 assign wire3293 = ( (~ ng11663)  &  ng10711 ) | ( (~ ng11600)  &  ng10711 ) | ( (~ ng11647)  &  ng10711 ) | ( (~ ng11663)  &  ng11600  &  (~ ng11647) ) ;
 assign ng11912 = ( wire3046 ) | ( wire7892 ) | ( wire33033 ) | ( wire33037 ) ;
 assign ng27567 = ( wire7879 ) | ( wire3196  &  (~ wire33053)  &  (~ wire33054) ) ;
 assign wire3570 = ( (~ ng823) ) | ( (~ wire34663)  &  (~ wire34664)  &  (~ wire34668) ) ;
 assign ng26887 = ( ng1448  &  ng23528  &  wire35156 ) ;
 assign ng26925 = ( ng25958 ) | ( wire32140 ) | ( ng12820  &  ng16655 ) | ( (~ ng12820)  &  (~ ng16655) ) ;
 assign ng26283 = ( ng11624  &  ng12781  &  (~ ng25954) ) | ( ng12781  &  (~ ng25954)  &  (~ wire30979) ) | ( (~ ng11624)  &  (~ ng12781)  &  (~ ng25954)  &  wire30979 ) ;
 assign ng18630 = ( wire7756 ) | ( wire33226 ) | ( wire33232 ) | ( wire33233 ) ;
 assign ng29748 = ( ng12324  &  ng12112  &  wire3074 ) | ( ng12324  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12324)  &  (~ ng12112)  &  ng21770  &  wire3074 ) ;
 assign ng27729 = ( wire5577 ) | ( ng23502  &  ng23489  &  wire35319 ) ;
 assign wire3150 = ( (~ ng23489) ) | ( (~ wire32106)  &  (~ wire32107)  &  (~ wire32108) ) ;
 assign ng30610 = ( wire35957 ) | ( wire3341  &  (~ wire34556)  &  (~ wire34557) ) ;
 assign ng30614 = ( wire36054 ) | ( wire3338  &  (~ wire34544)  &  (~ wire34545) ) ;
 assign wire3925 = ( ng2257  &  wire33588 ) | ( ng2257  &  wire33589 ) ;
 assign ng11807 = ( wire3046 ) | ( wire8679 ) | ( wire32017 ) | ( wire32021 ) ;
 assign ng29684 = ( wire5804 ) | ( wire5805 ) | ( wire35202 ) | ( wire35203 ) ;
 assign ng21996 = ( (~ ng12162)  &  wire3122 ) | ( ng12162  &  (~ wire33008)  &  (~ wire33009) ) ;
 assign ng26938 = ( (~ ng27582) ) | ( wire32952 ) ;
 assign ng26928 = ( (~ ng27582) ) | ( wire32952 ) | ( wire32954 ) ;
 assign ng25969 = ( (~ ng11687) ) | ( (~ ng11653) ) | ( (~ ng12994)  &  ng11678 ) | ( ng12994  &  ng11687  &  ng11653  &  (~ ng11678) ) ;
 assign wire3909 = ( (~ ng809)  &  (~ ng805)  &  ng801  &  ng813 ) ;
 assign ng23513 = ( ng853  &  (~ wire31297)  &  wire32164 ) | ( ng853  &  (~ wire31298)  &  wire32164 ) ;
 assign wire3439 = ( ng1196  &  wire32282 ) | ( ng1196  &  wire32283 ) ;
 assign ng18102 = ( wire6464 ) | ( wire6465 ) | ( wire34709 ) | ( wire34710 ) ;
 assign ng12179 = ( wire3046 ) | ( wire7278 ) | ( wire33857 ) | ( wire33861 ) ;
 assign ng12099 = ( wire6398 ) | ( wire6399 ) | ( wire34861 ) | ( wire34863 ) ;
 assign ng11991 = ( wire34851 ) | ( wire34852 ) ;
 assign ng11935 = ( wire31404 ) | ( wire31405 ) ;
 assign ng11773 = ( wire3046 ) | ( wire8114 ) | ( wire32785 ) | ( wire32789 ) ;
 assign ng26096 = ( wire35368 ) | ( wire3339  &  (~ wire31663)  &  (~ wire31664) ) ;
 assign ng26099 = ( wire35367 ) | ( wire3339  &  (~ wire31675)  &  (~ wire31676) ) ;
 assign wire3140 = ( ng557  &  (~ ng510) ) ;
 assign ng22005 = ( pg3229  &  wire32187  &  wire32199 ) | ( pg3229  &  wire32188  &  wire32199 ) | ( (~ pg3229)  &  (~ wire32187)  &  (~ wire32188)  &  wire32199 ) ;
 assign wire3595 = ( (~ ng826) ) | ( (~ wire34663)  &  (~ wire34664)  &  (~ wire34668) ) ;
 assign wire3236 = ( wire33793 ) | ( (~ ng2398)  &  ng823 ) ;
 assign ng25954 = ( (~ ng11644) ) | ( (~ ng13378) ) | ( ng11624  &  (~ ng12912) ) | ( ng11644  &  ng13378  &  (~ ng11624)  &  ng12912 ) ;
 assign ng25764 = ( wire9425 ) | ( wire31057  &  wire31058 ) ;
 assign wire3237 = ( wire31272 ) | ( (~ ng323)  &  ng823 ) ;
 assign wire3936 = ( ng2257  &  wire31077 ) | ( ng2257  &  wire31078 ) ;
 assign ng27738 = ( wire31274 ) | ( ng27834  &  wire31273 ) ;
 assign ng26897 = ( ng2142  &  ng23539  &  wire33829 ) ;
 assign ng27482 = ( wire8556 ) | ( wire8557 ) ;
 assign wire3118 = ( pg3229  &  wire31492 ) | ( pg3229  &  wire31493 ) | ( (~ pg3229)  &  (~ wire31492)  &  (~ wire31493) ) ;
 assign ng13399 = ( (~ pg8275)  &  pg8274  &  pg8273  &  pg8272 ) | ( pg8275  &  (~ pg8274)  &  pg8273  &  pg8272 ) | ( pg8275  &  pg8274  &  (~ pg8273)  &  pg8272 ) | ( (~ pg8275)  &  (~ pg8274)  &  (~ pg8273)  &  pg8272 ) | ( pg8275  &  pg8274  &  pg8273  &  (~ pg8272) ) | ( (~ pg8275)  &  (~ pg8274)  &  pg8273  &  (~ pg8272) ) | ( (~ pg8275)  &  pg8274  &  (~ pg8273)  &  (~ pg8272) ) | ( pg8275  &  (~ pg8274)  &  (~ pg8273)  &  (~ pg8272) ) ;
 assign ng30588 = ( wire36324 ) | ( wire3338  &  (~ wire34484)  &  (~ wire34485) ) ;
 assign ng30632 = ( wire36289 ) | ( wire3341  &  (~ wire34580)  &  (~ wire34581) ) ;
 assign wire3189 = ( ng2574  &  (~ ng30072)  &  ng12352  &  (~ wire35748) ) ;
 assign wire3338 = ( (~ ng12352)  &  wire3075  &  wire35745 ) | ( (~ ng12352)  &  wire3075  &  wire35746 ) ;
 assign ng30602 = ( wire36189 ) | ( wire3338  &  (~ wire34520)  &  (~ wire34521) ) ;
 assign ng25091 = ( ng11952  &  ng11875 ) | ( ng11952  &  wire3935 ) | ( ng11952  &  wire33025 ) | ( (~ ng11952)  &  (~ ng11875)  &  (~ wire33025) ) ;
 assign ng27814 = ( ng12249  &  (~ ng21746)  &  wire3076 ) | ( ng12249  &  ng11905  &  wire3076 ) | ( (~ ng12249)  &  ng21746  &  (~ ng11905)  &  wire3076 ) ;
 assign ng27827 = ( ng12288  &  (~ ng21746)  &  wire3076 ) | ( ng12288  &  ng11872  &  wire3076 ) | ( (~ ng12288)  &  ng21746  &  (~ ng11872)  &  wire3076 ) ;
 assign ng11988 = ( wire3046 ) | ( wire6468 ) | ( wire34696 ) | ( wire34700 ) ;
 assign ng22083 = ( pg3229  &  wire31492  &  wire34679 ) | ( pg3229  &  wire31493  &  wire34679 ) | ( (~ pg3229)  &  (~ wire31492)  &  (~ wire31493)  &  wire34679 ) ;
 assign ng22050 = ( (~ ng12080)  &  wire31502 ) | ( (~ ng12080)  &  wire31503 ) | ( (~ wire3118)  &  (~ wire31502)  &  (~ wire31503) ) ;
 assign ng23528 = ( ng853  &  (~ wire31297)  &  wire32975 ) | ( ng853  &  (~ wire31298)  &  wire32975 ) ;
 assign ng10711 = ( (~ ng2892)  &  (~ ng2903)  &  wire31298 ) ;
 assign ng26107 = ( wire35565 ) | ( wire3336  &  (~ wire31723)  &  (~ wire31724) ) ;
 assign ng26110 = ( wire35564 ) | ( wire3336  &  (~ wire31639)  &  (~ wire31640) ) ;
 assign wire3141 = ( (~ ng1890)  &  (~ ng1937)  &  ng1905 ) ;
 assign wire3229 = ( ng1890  &  (~ ng1937) ) ;
 assign wire3833 = ( wire3277 ) | ( wire3280  &  wire35716 ) | ( wire3280  &  wire35717 ) ;
 assign wire3137 = ( (~ ng2631)  &  (~ ng2584)  &  ng2599 ) ;
 assign wire3230 = ( (~ ng2631)  &  ng2584 ) ;
 assign ng13055 = ( wire31522  &  wire31523  &  wire31524 ) ;
 assign ng11831 = ( wire31663 ) | ( wire31664 ) ;
 assign ng11872 = ( wire6374 ) | ( wire6375 ) | ( wire34825 ) | ( wire34827 ) ;
 assign ng13004 = ( wire35758  &  wire35759 ) ;
 assign ng23353 = ( (~ ng12179)  &  wire3120 ) | ( ng12179  &  (~ wire3120)  &  wire34421 ) | ( ng12179  &  (~ wire3120)  &  wire34422 ) ;
 assign wire3389 = ( (~ ng744) ) | ( (~ ng762) ) | ( (~ ng23513) ) | ( (~ wire32166) ) ;
 assign ng26941 = ( (~ ng27585) ) | ( wire33805 ) | ( wire33807 ) ;
 assign wire3119 = ( (~ pg3229)  &  wire33137 ) | ( (~ pg3229)  &  wire33138 ) | ( pg3229  &  (~ wire33137)  &  (~ wire33138) ) ;
 assign ng22093 = ( (~ ng12214)  &  wire33117 ) | ( (~ ng12214)  &  wire33118 ) | ( wire3119  &  (~ wire33117)  &  (~ wire33118) ) ;
 assign ng27855 = ( ng12249  &  (~ ng21746)  &  wire3076 ) | ( ng12249  &  ng12208  &  wire3076 ) | ( (~ ng12249)  &  ng21746  &  (~ ng12208)  &  wire3076 ) ;
 assign ng29721 = ( ng12324  &  ng11914  &  wire3074 ) | ( ng12324  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12324)  &  (~ ng11914)  &  ng21770  &  wire3074 ) ;
 assign ng22108 = ( pg3229  &  wire32323  &  wire35281 ) | ( pg3229  &  wire32324  &  wire35281 ) | ( (~ pg3229)  &  (~ wire32323)  &  (~ wire32324)  &  wire35281 ) ;
 assign ng23331 = ( (~ ng11974)  &  (~ wire3121) ) | ( ng11974  &  wire3121  &  wire34636 ) | ( ng11974  &  wire3121  &  wire34637 ) ;
 assign ng23325 = ( wire4376 ) | ( wire4379 ) | ( wire36115 ) ;
 assign wire3151 = ( ng12180  &  wire7190 ) | ( ng12180  &  wire7191 ) | ( ng12180  &  wire7192 ) | ( (~ ng12180)  &  (~ wire7190)  &  (~ wire7191)  &  (~ wire7192) ) ;
 assign ng18556 = ( (~ wire32590)  &  (~ wire32591)  &  wire32828 ) | ( (~ wire32590)  &  (~ wire32591)  &  wire32829 ) | ( wire32590  &  (~ wire32828)  &  (~ wire32829) ) | ( wire32591  &  (~ wire32828)  &  (~ wire32829) ) ;
 assign ng18212 = ( ng1476  &  wire32691 ) | ( ng1476  &  wire32692 ) | ( (~ ng1476)  &  (~ wire32691)  &  (~ wire32692) ) ;
 assign ng18115 = ( ng1486  &  wire32671 ) | ( ng1486  &  wire32672 ) | ( (~ ng1486)  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire3108 = ( (~ ng1496)  &  wire32661 ) | ( (~ ng1496)  &  wire32662 ) | ( ng1496  &  (~ wire32661)  &  (~ wire32662) ) ;
 assign wire3297 = ( (~ ng17942)  &  (~ ng18212) ) | ( (~ ng18556)  &  (~ ng18115) ) ;
 assign ng23505 = ( wire32938 ) | ( wire32939 ) | ( wire32940 ) ;
 assign ng11839 = ( wire3046 ) | ( wire8070 ) | ( wire32865 ) | ( wire32869 ) ;
 assign wire3216 = ( (~ ng1315) ) | ( (~ ng2704) ) ;
 assign ng11863 = ( wire3049 ) | ( wire8947 ) | ( wire31672 ) | ( wire31676 ) ;
 assign ng30597 = ( wire36171 ) | ( wire3341  &  (~ wire34568)  &  (~ wire34569) ) ;
 assign wire3198 = ( ng2631  &  (~ ng2584) ) ;
 assign ng27382 = ( (~ ng26087)  &  ng26154  &  ng26099  &  ng26110 ) | ( ng26087  &  (~ ng26154)  &  ng26099  &  ng26110 ) | ( ng26087  &  ng26154  &  (~ ng26099)  &  ng26110 ) | ( (~ ng26087)  &  (~ ng26154)  &  (~ ng26099)  &  ng26110 ) | ( ng26087  &  ng26154  &  ng26099  &  (~ ng26110) ) | ( (~ ng26087)  &  (~ ng26154)  &  ng26099  &  (~ ng26110) ) | ( (~ ng26087)  &  ng26154  &  (~ ng26099)  &  (~ ng26110) ) | ( ng26087  &  (~ ng26154)  &  (~ ng26099)  &  (~ ng26110) ) ;
 assign ng27379 = ( (~ ng26137)  &  ng26126  &  ng26145  &  ng26151 ) | ( ng26137  &  (~ ng26126)  &  ng26145  &  ng26151 ) | ( ng26137  &  ng26126  &  (~ ng26145)  &  ng26151 ) | ( (~ ng26137)  &  (~ ng26126)  &  (~ ng26145)  &  ng26151 ) | ( ng26137  &  ng26126  &  ng26145  &  (~ ng26151) ) | ( (~ ng26137)  &  (~ ng26126)  &  ng26145  &  (~ ng26151) ) | ( (~ ng26137)  &  ng26126  &  (~ ng26145)  &  (~ ng26151) ) | ( ng26137  &  (~ ng26126)  &  (~ ng26145)  &  (~ ng26151) ) ;
 assign ng28845 = ( (~ ng27802)  &  ng27814  &  ng27827  &  ng27900 ) | ( ng27802  &  (~ ng27814)  &  ng27827  &  ng27900 ) | ( ng27802  &  ng27814  &  (~ ng27827)  &  ng27900 ) | ( (~ ng27802)  &  (~ ng27814)  &  (~ ng27827)  &  ng27900 ) | ( ng27802  &  ng27814  &  ng27827  &  (~ ng27900) ) | ( (~ ng27802)  &  (~ ng27814)  &  ng27827  &  (~ ng27900) ) | ( (~ ng27802)  &  ng27814  &  (~ ng27827)  &  (~ ng27900) ) | ( ng27802  &  (~ ng27814)  &  (~ ng27827)  &  (~ ng27900) ) ;
 assign ng27113 = ( wire30883 ) | ( wire35816 ) | ( ng21851  &  wire30881 ) ;
 assign wire3143 = ( ng1211  &  (~ ng1196)  &  (~ ng1243) ) ;
 assign ng30629 = ( wire35864 ) | ( wire3338  &  (~ wire34508)  &  (~ wire34509) ) ;
 assign wire3427 = ( ng17194  &  ng30305 ) | ( ng17194  &  (~ ng17183)  &  (~ ng30305)  &  (~ wire35751) ) ;
 assign ng11744 = ( wire3046 ) | ( wire9368 ) | ( wire31102 ) | ( wire31106 ) ;
 assign ng11905 = ( wire34791 ) | ( wire34792 ) ;
 assign ng12154 = ( wire3049 ) | ( wire6337 ) | ( wire34776 ) | ( wire34780 ) ;
 assign ng12048 = ( wire34767 ) | ( wire34768 ) ;
 assign ng22134 = ( pg3229  &  wire3440  &  wire33137 ) | ( pg3229  &  wire3440  &  wire33138 ) | ( (~ pg3229)  &  wire3440  &  (~ wire33137)  &  (~ wire33138) ) ;
 assign ng26902 = ( (~ ng27563) ) | ( wire31279 ) | ( wire31281 ) ;
 assign ng26892 = ( (~ ng27563) ) | ( wire31279 ) | ( wire31281 ) | ( wire31283 ) ;
 assign wire3302 = ( ng11630  &  ng11666  &  wire32630 ) | ( ng11630  &  (~ ng11666)  &  wire32630 ) | ( ng11630  &  ng11666  &  wire32631 ) | ( ng11630  &  (~ ng11666)  &  wire32631 ) ;
 assign ng26906 = ( ng26925 ) | ( wire32142 ) | ( wire32155 ) ;
 assign ng27462 = ( ng11624  &  ng12747  &  (~ ng26892) ) | ( ng12747  &  (~ ng26892)  &  (~ wire30979) ) | ( (~ ng11624)  &  (~ ng12747)  &  (~ ng26892)  &  wire30979 ) ;
 assign ng27900 = ( ng12249  &  (~ ng21746)  &  wire3076 ) | ( ng12249  &  ng11991  &  wire3076 ) | ( (~ ng12249)  &  ng21746  &  (~ ng11991)  &  wire3076 ) ;
 assign ng27730 = ( wire7837 ) | ( ng23518  &  ng23505  &  wire33102 ) ;
 assign ng30605 = ( wire36188 ) | ( wire3338  &  (~ wire34472)  &  (~ wire34473) ) ;
 assign ng30927 = ( (~ ng30588)  &  ng30632  &  ng30597  &  ng30605 ) | ( ng30588  &  (~ ng30632)  &  ng30597  &  ng30605 ) | ( ng30588  &  ng30632  &  (~ ng30597)  &  ng30605 ) | ( (~ ng30588)  &  (~ ng30632)  &  (~ ng30597)  &  ng30605 ) | ( ng30588  &  ng30632  &  ng30597  &  (~ ng30605) ) | ( (~ ng30588)  &  (~ ng30632)  &  ng30597  &  (~ ng30605) ) | ( (~ ng30588)  &  ng30632  &  (~ ng30597)  &  (~ ng30605) ) | ( ng30588  &  (~ ng30632)  &  (~ ng30597)  &  (~ ng30605) ) ;
 assign wire3303 = ( (~ ng762) ) | ( (~ ng23513) ) ;
 assign ng23320 = ( wire6544 ) | ( wire6545 ) | ( wire6546 ) ;
 assign wire3395 = ( (~ ng2892) ) | ( (~ ng2950) ) | ( (~ ng2903) ) | ( (~ wire35033) ) ;
 assign ng11987 = ( wire3046 ) | ( wire8524 ) | ( wire32184 ) | ( wire32188 ) ;
 assign wire3277 = ( ng17177  &  wire9559 ) | ( ng17177  &  wire30886 ) | ( ng17177  &  wire35568 ) ;
 assign wire3227 = ( ng1196  &  (~ ng1243) ) ;
 assign wire3835 = ( wire3278 ) | ( wire3279  &  wire35952 ) | ( wire3279  &  wire35953 ) ;
 assign wire3834 = ( wire3277 ) | ( wire3280  &  (~ wire35716)  &  (~ wire35717) ) ;
 assign wire3442 = ( ng1890  &  wire33157 ) | ( ng1890  &  wire33158 ) ;
 assign ng22118 = ( (~ ng12269)  &  wire34008 ) | ( (~ ng12269)  &  wire34009 ) | ( (~ wire3124)  &  (~ wire34008)  &  (~ wire34009) ) ;
 assign ng27157 = ( wire8280 ) | ( (~ ng23107)  &  wire32539 ) | ( (~ ng23107)  &  wire32564 ) ;
 assign ng26911 = ( (~ ng27563) ) | ( wire31279 ) ;
 assign wire3120 = ( pg3229  &  wire33840 ) | ( pg3229  &  wire33841 ) | ( (~ pg3229)  &  (~ wire33840)  &  (~ wire33841) ) ;
 assign ng27897 = ( ng12288  &  (~ ng21746)  &  wire3076 ) | ( ng12288  &  ng12048  &  wire3076 ) | ( (~ ng12288)  &  ng21746  &  (~ ng12048)  &  wire3076 ) ;
 assign ng17194 = ( ng2631  &  (~ ng2584) ) | ( (~ ng2584)  &  ng2599 ) ;
 assign ng17177 = ( (~ ng1890)  &  ng1937 ) | ( (~ ng1890)  &  ng1905 ) ;
 assign ng11992 = ( wire3046 ) | ( wire8098 ) | ( wire32765 ) | ( wire32769 ) ;
 assign ng11938 = ( wire31651 ) | ( wire31652 ) ;
 assign wire3278 = ( ng1211  &  (~ ng1196)  &  ng27113 ) | ( (~ ng1196)  &  ng1243  &  ng27113 ) ;
 assign ng27865 = ( ng12288  &  (~ ng21746)  &  wire3076 ) | ( ng12288  &  ng12154  &  wire3076 ) | ( (~ ng12288)  &  ng21746  &  (~ ng12154)  &  wire3076 ) ;
 assign wire3836 = ( wire3278 ) | ( wire3279  &  (~ wire35952)  &  (~ wire35953) ) ;
 assign ng11830 = ( wire31639 ) | ( wire31640 ) ;
 assign wire3217 = ( (~ ng8381)  &  (~ wire30893) ) | ( (~ wire3246)  &  (~ ng8381)  &  (~ wire30892) ) ;
 assign ng15757 = ( ng3135 ) | ( ng3120 ) | ( (~ ng8430) ) | ( wire30897 ) ;
 assign ng15719 = ( ng3135 ) | ( ng3120 ) | ( wire3246 ) | ( (~ ng8430) ) ;
 assign ng15841 = ( ng3135 ) | ( ng3120 ) | ( (~ ng8430) ) | ( wire30896 ) ;
 assign wire3397 = ( ng3135  &  ng3120  &  (~ wire3246)  &  (~ ng8381) ) | ( ng3135  &  (~ ng3120)  &  (~ wire3246)  &  (~ ng8381) ) ;
 assign ng27582 = ( ng12992  &  (~ ng16672)  &  ng12858  &  (~ ng25964) ) | ( (~ ng12992)  &  ng16672  &  (~ ng12858)  &  (~ ng25964) ) ;
 assign ng30031 = ( (~ ng24695)  &  (~ ng11647)  &  wire5571 ) | ( (~ ng24695)  &  (~ ng11647)  &  wire35331 ) | ( (~ ng24695)  &  ng11647  &  (~ wire5571)  &  (~ wire35331) ) ;
 assign ng23388 = ( (~ ng12214)  &  (~ wire3119) ) | ( ng12214  &  wire3119  &  wire33338 ) | ( ng12214  &  wire3119  &  wire33339 ) ;
 assign wire3307 = ( (~ ng826) ) | ( ng133 ) ;
 assign wire3308 = ( ng149 ) | ( (~ ng823) ) ;
 assign ng12057 = ( wire3046 ) | ( wire7850 ) | ( wire33070 ) | ( wire33074 ) ;
 assign ng23360 = ( wire9041 ) | ( wire9044 ) | ( wire31518 ) ;
 assign ng23950 = ( ng646  &  wire31591  &  wire31592  &  wire34989 ) ;
 assign ng17183 = ( (~ ng2631)  &  ng2584 ) | ( (~ ng2631)  &  ng2599 ) ;
 assign wire3400 = ( (~ ng1448) ) | ( (~ ng1430) ) | ( (~ ng23528) ) | ( (~ wire35156) ) ;
 assign ng26417 = ( (~ ng16693)  &  (~ ng25969)  &  wire33508 ) | ( (~ ng16693)  &  (~ ng25969)  &  wire33509 ) | ( ng16693  &  (~ ng25969)  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign wire3323 = ( (~ ng2142) ) | ( (~ ng23539) ) ;
 assign wire3403 = ( (~ ng3013) ) | ( (~ ng3002) ) | ( (~ ng3006) ) | ( wire3333 ) ;
 assign wire3921 = ( ng1491  &  (~ ng1496)  &  ng1506  &  (~ ng1501) ) ;
 assign ng23497 = ( ng853  &  (~ wire31297)  &  wire34625 ) | ( ng853  &  (~ wire31298)  &  wire34625 ) ;
 assign ng17162 = ( ng1211  &  (~ ng1196) ) | ( (~ ng1196)  &  ng1243 ) ;
 assign ng30305 = ( pg2637 ) | ( ng30072 ) | ( ng2633 ) ;
 assign ng11981 = ( wire3046 ) | ( wire8713 ) | ( wire31983 ) | ( wire31987 ) ;
 assign wire3174 = ( (~ wire3073)  &  wire31469 ) | ( (~ wire3073)  &  wire31470 ) ;
 assign wire3339 = ( (~ ng12194)  &  (~ wire3073)  &  wire34048 ) | ( (~ ng12194)  &  (~ wire3073)  &  wire34049 ) ;
 assign wire3942 = ( ng113  &  (~ ng117)  &  (~ ng121)  &  ng125 ) ;
 assign wire3313 = ( (~ ng11687)  &  ng10711 ) | ( (~ ng11653)  &  ng10711 ) | ( (~ ng11678)  &  ng10711 ) | ( (~ ng11687)  &  ng11653  &  (~ ng11678) ) ;
 assign ng23526 = ( wire3386 ) | ( wire33097  &  wire33098  &  wire33099 ) ;
 assign ng8381 = ( ng3110 ) | ( ng3124 ) | ( ng3126 ) | ( ng3191 ) ;
 assign ng12082 = ( wire31627 ) | ( wire31628 ) ;
 assign ng29710 = ( ng12292  &  ng11915  &  wire3074 ) | ( ng12292  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12292)  &  (~ ng11915)  &  ng21770  &  wire3074 ) ;
 assign wire3280 = ( (~ ng1890)  &  ng1937 ) ;
 assign ng11974 = ( wire3046 ) | ( wire9218 ) | ( wire31331 ) | ( wire31335 ) ;
 assign wire3314 = ( ng11653  &  ng11678  &  wire33528 ) | ( ng11653  &  (~ ng11678)  &  wire33528 ) | ( ng11653  &  ng11678  &  wire33529 ) | ( ng11653  &  (~ ng11678)  &  wire33529 ) ;
 assign ng11188 = ( (~ ng2981)  &  ng2874  &  ng2975  &  ng2978 ) | ( ng2981  &  (~ ng2874)  &  ng2975  &  ng2978 ) | ( ng2981  &  ng2874  &  (~ ng2975)  &  ng2978 ) | ( (~ ng2981)  &  (~ ng2874)  &  (~ ng2975)  &  ng2978 ) | ( ng2981  &  ng2874  &  ng2975  &  (~ ng2978) ) | ( (~ ng2981)  &  (~ ng2874)  &  ng2975  &  (~ ng2978) ) | ( (~ ng2981)  &  ng2874  &  (~ ng2975)  &  (~ ng2978) ) | ( ng2981  &  (~ ng2874)  &  (~ ng2975)  &  (~ ng2978) ) ;
 assign ng12988 = ( (~ pg8265)  &  pg8266  &  pg8264  &  pg8262 ) | ( pg8265  &  (~ pg8266)  &  pg8264  &  pg8262 ) | ( pg8265  &  pg8266  &  (~ pg8264)  &  pg8262 ) | ( (~ pg8265)  &  (~ pg8266)  &  (~ pg8264)  &  pg8262 ) | ( pg8265  &  pg8266  &  pg8264  &  (~ pg8262) ) | ( (~ pg8265)  &  (~ pg8266)  &  pg8264  &  (~ pg8262) ) | ( (~ pg8265)  &  pg8266  &  (~ pg8264)  &  (~ pg8262) ) | ( pg8265  &  (~ pg8266)  &  (~ pg8264)  &  (~ pg8262) ) ;
 assign wire3188 = ( (~ wire3073)  &  wire31449 ) | ( (~ wire3073)  &  wire31450 ) ;
 assign wire3336 = ( (~ ng12245)  &  (~ wire3073)  &  wire34048 ) | ( (~ ng12245)  &  (~ wire3073)  &  wire34049 ) ;
 assign wire3697 = ( (~ ng823) ) | ( (~ wire34737)  &  (~ wire34738)  &  (~ wire34741) ) ;
 assign wire3156 = ( ng11975  &  wire9128 ) | ( ng11975  &  wire9129 ) | ( ng11975  &  wire9130 ) | ( (~ ng11975)  &  (~ wire9128)  &  (~ wire9129)  &  (~ wire9130) ) ;
 assign wire3435 = ( ng2584  &  wire33967 ) | ( ng2584  &  wire33968 ) ;
 assign wire3315 = ( (~ ng853) ) | ( ng841 ) ;
 assign wire3316 = ( ng852 ) | ( (~ ng823) ) ;
 assign wire3317 = ( ng13378  &  ng11624  &  wire30957 ) | ( ng13378  &  (~ ng11624)  &  wire30957 ) | ( ng13378  &  ng11624  &  wire30958 ) | ( ng13378  &  (~ ng11624)  &  wire30958 ) ;
 assign wire3195 = ( ng2257  &  (~ ng25078)  &  (~ wire31345)  &  (~ wire31346) ) ;
 assign ng11262 = ( (~ ng2969)  &  ng2972  &  ng2963  &  ng2966 ) | ( ng2969  &  (~ ng2972)  &  ng2963  &  ng2966 ) | ( ng2969  &  ng2972  &  (~ ng2963)  &  ng2966 ) | ( (~ ng2969)  &  (~ ng2972)  &  (~ ng2963)  &  ng2966 ) | ( ng2969  &  ng2972  &  ng2963  &  (~ ng2966) ) | ( (~ ng2969)  &  (~ ng2972)  &  ng2963  &  (~ ng2966) ) | ( (~ ng2969)  &  ng2972  &  (~ ng2963)  &  (~ ng2966) ) | ( ng2969  &  (~ ng2972)  &  (~ ng2963)  &  (~ ng2966) ) ;
 assign wire3309 = ( (~ ng11675)  &  ng10711 ) | ( (~ ng11630)  &  ng10711 ) | ( (~ ng11666)  &  ng10711 ) | ( (~ ng11675)  &  ng11630  &  (~ ng11666) ) ;
 assign ng11979 = ( wire3049 ) | ( wire8915 ) | ( wire31602 ) | ( wire31606 ) ;
 assign ng12036 = ( wire8912 ) | ( wire8913 ) | ( wire31613 ) | ( wire31615 ) ;
 assign wire3279 = ( (~ ng1196)  &  ng1243 ) ;
 assign ng29718 = ( ng12324  &  ng12293  &  wire3074 ) | ( ng12324  &  (~ ng21770)  &  wire3074 ) | ( (~ ng12324)  &  (~ ng12293)  &  ng21770  &  wire3074 ) ;
 assign wire3319 = ( (~ ng646) ) | ( (~ ng633) ) | ( (~ ng640) ) | ( (~ wire31592) ) ;
 assign wire3157 = ( ng12044  &  wire5893 ) | ( ng12044  &  wire5894 ) | ( ng12044  &  wire5895 ) | ( (~ ng12044)  &  (~ wire5893)  &  (~ wire5894)  &  (~ wire5895) ) ;
 assign ng12026 = ( wire3046 ) | ( wire9210 ) | ( wire31311 ) | ( wire31315 ) ;
 assign wire3121 = ( (~ pg3229)  &  wire31324 ) | ( (~ pg3229)  &  wire31325 ) | ( pg3229  &  (~ wire31324)  &  (~ wire31325) ) ;
 assign wire3122 = ( (~ pg3229)  &  wire32998 ) | ( (~ pg3229)  &  wire32999 ) | ( pg3229  &  (~ wire32998)  &  (~ wire32999) ) ;
 assign ng12090 = ( wire32197 ) | ( wire32198 ) ;
 assign ng12224 = ( wire3046 ) | ( wire7270 ) | ( wire33847 ) | ( wire33851 ) ;
 assign ng22009 = ( (~ wire3120)  &  (~ ng12224) ) | ( ng12224  &  (~ wire33860)  &  (~ wire33861) ) ;
 assign wire3123 = ( pg3229  &  wire32323 ) | ( pg3229  &  wire32324 ) | ( (~ pg3229)  &  (~ wire32323)  &  (~ wire32324) ) ;
 assign wire3124 = ( pg3229  &  wire33998 ) | ( pg3229  &  wire33999 ) | ( (~ pg3229)  &  (~ wire33998)  &  (~ wire33999) ) ;
 assign ng23395 = ( (~ ng12269)  &  wire3124 ) | ( ng12269  &  (~ wire3124)  &  wire33988 ) | ( ng12269  &  (~ wire3124)  &  wire33989 ) ;
 assign wire3324 = ( (~ ng74) ) | ( (~ ng23497) ) ;
 assign ng23381 = ( wire7111 ) | ( wire7114 ) | ( wire34024 ) ;
 assign ng21983 = ( (~ wire3117)  &  (~ ng12090) ) | ( ng12090  &  (~ wire32177)  &  (~ wire32178) ) ;
 assign ng22069 = ( (~ ng12207)  &  (~ wire3123) ) | ( ng12207  &  (~ wire32313)  &  (~ wire32314) ) ;
 assign wire3320 = ( ng1515 ) | ( (~ ng826) ) ;
 assign wire3321 = ( ng1531 ) | ( (~ ng823) ) ;
 assign ng22021 = ( pg3229  &  wire33840  &  wire35306 ) | ( pg3229  &  wire33841  &  wire35306 ) | ( (~ pg3229)  &  (~ wire33840)  &  (~ wire33841)  &  wire35306 ) ;
 assign wire3159 = ( ng12108  &  wire7844 ) | ( ng12108  &  wire7845 ) | ( ng12108  &  wire7846 ) | ( (~ ng12108)  &  (~ wire7844)  &  (~ wire7845)  &  (~ wire7846) ) ;
 assign ng12213 = ( wire3046 ) | ( wire6278 ) | ( wire34924 ) | ( wire34928 ) ;
 assign ng23364 = ( wire5883 ) | ( wire5886 ) | ( wire35154 ) ;
 assign wire3325 = ( (~ ng1448) ) | ( (~ ng23528) ) ;
 assign wire3073 = ( (~ ng499) ) | ( ng21851 ) | ( wire34028 ) ;
 assign ng17139 = ( ng557  &  (~ ng510) ) | ( (~ ng510)  &  ng525 ) ;
 assign ng23344 = ( wire5793 ) | ( wire5794 ) | ( wire5795 ) ;
 assign wire3784 = ( (~ ng826) ) | ( (~ wire34737)  &  (~ wire34738)  &  (~ wire34741) ) ;
 assign wire3788 = ( (~ ng853) ) | ( (~ wire34663)  &  (~ wire34664)  &  (~ wire34668) ) ;
 assign ng26918 = ( (~ ng27582) ) | ( wire32952 ) | ( wire32954 ) | ( wire32956 ) ;
 assign wire3074 = ( ng1880  &  (~ wire9559)  &  (~ wire30886)  &  (~ wire35568) ) ;
 assign wire3075 = ( (~ pg2637)  &  ng2574  &  (~ ng30072)  &  (~ ng2633) ) ;
 assign wire3076 = ( ng1186  &  (~ ng27113) ) ;
 assign wire3116 = ( pg3231 ) | ( (~ ng3139) ) ;
 assign pg8012 = ( ng826 ) ;
 assign pg8167 = ( ng823 ) ;
 assign pg7161 = ( ng1312 ) ;
 assign pg7194 = ( ng1312 ) ;
 assign pg7052 = ( ng1309 ) ;
 assign pg7390 = ( ng1312 ) ;
 assign pg6573 = ( ng826 ) ;
 assign pg7084 = ( ng823 ) ;
 assign pg7264 = ( ng823 ) ;
 assign pg8007 = ( ng823 ) ;
 assign pg8106 = ( ng1309 ) ;
 assign pg6642 = ( ng1312 ) ;
 assign pg6750 = ( ng1309 ) ;
 assign pg7302 = ( ng1309 ) ;
 assign pg5472 = ( ng826 ) ;
 assign pg8030 = ( ng1312 ) ;
 assign pg5511 = ( ng826 ) ;
 assign pg7014 = ( ng823 ) ;
 assign pg6313 = ( ng823 ) ;
 assign pg5612 = ( ng2258 ) ;
 assign pg6231 = ( ng826 ) ;
 assign pg5437 = ( ng826 ) ;
 assign pg5657 = ( ng1309 ) ;
 assign pg6979 = ( ng1309 ) ;
 assign pg6911 = ( ng1312 ) ;
 assign pg6944 = ( ng1312 ) ;
 assign pg6712 = ( ng823 ) ;
 assign pg6837 = ( ng826 ) ;
 assign pg5686 = ( ng1312 ) ;
 assign pg5738 = ( ng1312 ) ;
 assign pg6447 = ( ng823 ) ;
 assign pg5555 = ( ng826 ) ;
 assign pg7229 = ( ng1309 ) ;
 assign pg5549 = ( ng2258 ) ;
 assign pg5637 = ( ng2258 ) ;
 assign pg5648 = ( ng1312 ) ;
 assign pg5747 = ( ng1309 ) ;
 assign pg5629 = ( ng1309 ) ;
 assign pg6518 = ( ng823 ) ;
 assign pg7425 = ( ng1309 ) ;
 assign pg5595 = ( ng2258 ) ;
 assign pg8082 = ( ng823 ) ;
 assign pg5695 = ( ng1309 ) ;
 assign pg6368 = ( ng826 ) ;
 assign pg6485 = ( ng1309 ) ;
 assign pg6782 = ( ng823 ) ;
 assign pg7961 = ( ng826 ) ;
 assign pg7357 = ( ng1312 ) ;
 assign pg5796 = ( ng1312 ) ;
 assign pg7909 = ( ng826 ) ;
 assign pg7956 = ( ng823 ) ;
 assign pg6677 = ( ng1309 ) ;
 assign pg8087 = ( ng826 ) ;
 assign pg7487 = ( ng1312 ) ;
 assign wire3034 = ( ng3097  &  ng3139  &  ng3120  &  ng3147 ) ;
 assign wire3035 = ( (~ ng3120)  &  (~ ng3147)  &  ng2984 ) | ( (~ ng3120)  &  (~ ng3147)  &  ng2985 ) ;
 assign wire3036 = ( (~ ng3139)  &  ng2991  &  (~ ng3147) ) | ( (~ ng3139)  &  ng2992  &  (~ ng3147) ) ;
 assign wire3037 = ( (~ ng3139)  &  (~ ng3120)  &  (~ ng3147) ) ;
 assign wire3050 = ( ng1312  &  wire7635 ) | ( ng1312  &  wire7636 ) | ( ng1312  &  wire7637 ) ;
 assign wire3079 = ( ng1309  &  wire7635 ) | ( ng1309  &  wire7636 ) | ( ng1309  &  wire7637 ) ;
 assign wire3097 = ( wire3142  &  (~ wire33296)  &  (~ wire33297)  &  (~ wire33298) ) ;
 assign wire3101 = ( ng2879  &  ng11188  &  ng11262  &  wire3116 ) | ( ng2879  &  (~ ng11188)  &  (~ ng11262)  &  wire3116 ) | ( ng2879  &  (~ ng11188)  &  ng11262  &  (~ wire3116) ) | ( ng2879  &  ng11188  &  (~ ng11262)  &  (~ wire3116) ) ;
 assign wire3167 = ( ng18630  &  (~ wire33376)  &  (~ wire33377)  &  wire36459 ) ;
 assign wire3168 = ( wire7640  &  wire36462 ) | ( wire33399  &  wire36462 ) | ( wire33401  &  wire36462 ) ;
 assign wire3213 = ( (~ ng2257)  &  ng1702  &  ng17124 ) | ( ng1702  &  (~ ng17124)  &  ng23526 ) ;
 assign wire3322 = ( ng823  &  (~ ng24712)  &  wire35163 ) | ( ng823  &  (~ ng24712)  &  wire35164 ) ;
 assign wire3388 = ( ng1868  &  ng1867  &  ng1869 ) ;
 assign wire3390 = ( (~ ng1315)  &  ng1867  &  ng1869 ) ;
 assign wire3391 = ( (~ ng1312)  &  ng1868  &  ng1869 ) ;
 assign wire3392 = ( (~ ng1309)  &  ng1868  &  ng1867 ) ;
 assign wire3393 = ( (~ ng1312)  &  (~ ng1315)  &  ng1869 ) ;
 assign wire3394 = ( (~ ng1312)  &  (~ ng1309)  &  ng1868 ) ;
 assign wire3396 = ( (~ ng1315)  &  (~ ng1309)  &  ng1867 ) ;
 assign wire3404 = ( ng826  &  (~ ng2257)  &  (~ ng12057) ) | ( ng826  &  (~ ng18218)  &  (~ ng12057) ) | ( ng826  &  ng2257  &  (~ ng18218)  &  ng12057 ) ;
 assign wire3422 = ( wire36426  &  wire36431 ) | ( wire36427  &  wire36431 ) | ( wire36428  &  wire36431 ) ;
 assign wire3423 = ( wire36426  &  wire36433 ) | ( wire36427  &  wire36433 ) | ( wire36428  &  wire36433 ) ;
 assign wire3424 = ( wire36426  &  wire36435 ) | ( wire36427  &  wire36435 ) | ( wire36428  &  wire36435 ) ;
 assign wire3441 = ( wire36426  &  wire36437 ) | ( wire36427  &  wire36437 ) | ( wire36428  &  wire36437 ) ;
 assign wire3448 = ( wire36426  &  wire36438 ) | ( wire36427  &  wire36438 ) | ( wire36428  &  wire36438 ) ;
 assign wire3449 = ( wire36426  &  wire36439 ) | ( wire36427  &  wire36439 ) | ( wire36428  &  wire36439 ) ;
 assign wire3450 = ( wire36426  &  wire36440 ) | ( wire36427  &  wire36440 ) | ( wire36428  &  wire36440 ) ;
 assign wire3451 = ( wire3049  &  wire36426 ) | ( wire3049  &  wire36427 ) | ( wire3049  &  wire36428 ) ;
 assign wire3488 = ( ng2879  &  ng11330  &  ng11263  &  wire3116 ) | ( ng2879  &  (~ ng11330)  &  (~ ng11263)  &  wire3116 ) | ( ng2879  &  (~ ng11330)  &  ng11263  &  (~ wire3116) ) | ( ng2879  &  ng11330  &  (~ ng11263)  &  (~ wire3116) ) ;
 assign wire3512 = ( (~ ng2924)  &  ng2920  &  (~ wire3139) ) | ( (~ ng2924)  &  ng2920  &  wire36378 ) ;
 assign wire3515 = ( (~ ng15970)  &  (~ wire33906)  &  (~ wire33907)  &  wire35395 ) ;
 assign wire3527 = ( (~ wire3139)  &  (~ wire36379)  &  wire36385 ) | ( wire36378  &  (~ wire36379)  &  wire36385 ) ;
 assign wire3528 = ( (~ ng2917)  &  ng2924  &  (~ wire3139) ) | ( (~ ng2917)  &  ng2924  &  wire36378 ) ;
 assign wire3529 = ( ng2924  &  wire3545 ) | ( ng2924  &  wire36383 ) ;
 assign wire3545 = ( (~ wire3139)  &  (~ wire36379)  &  wire36382 ) | ( wire36378  &  (~ wire36379)  &  wire36382 ) ;
 assign wire3564 = ( (~ pg8021)  &  ng2924 ) | ( (~ pg8021)  &  (~ ng2920) ) ;
 assign wire3594 = ( ng3032  &  (~ ng3036)  &  ng21796 ) | ( ng3032  &  (~ ng3036)  &  wire36176 ) ;
 assign wire3621 = ( (~ ng2879)  &  ng11330  &  ng11263  &  wire3116 ) | ( (~ ng2879)  &  (~ ng11330)  &  (~ ng11263)  &  wire3116 ) | ( (~ ng2879)  &  (~ ng11330)  &  ng11263  &  (~ wire3116) ) | ( (~ ng2879)  &  ng11330  &  (~ ng11263)  &  (~ wire3116) ) ;
 assign wire3639 = ( (~ ng2879)  &  ng11188  &  ng11262  &  wire3116 ) | ( (~ ng2879)  &  (~ ng11188)  &  (~ ng11262)  &  wire3116 ) | ( (~ ng2879)  &  (~ ng11188)  &  ng11262  &  (~ wire3116) ) | ( (~ ng2879)  &  ng11188  &  (~ ng11262)  &  (~ wire3116) ) ;
 assign wire3660 = ( wire3141  &  wire9559 ) | ( wire3141  &  wire30886 ) | ( wire3141  &  wire35568 ) ;
 assign wire3661 = ( (~ ng1890)  &  ng1917  &  (~ ng1937)  &  ng1905 ) ;
 assign wire3672 = ( (~ wire9559)  &  (~ wire30886)  &  (~ wire35568)  &  wire36331 ) ;
 assign wire3673 = ( (~ wire9559)  &  (~ wire30886)  &  (~ wire35568)  &  wire36335 ) ;
 assign wire3714 = ( ng12068  &  wire3230  &  (~ wire36324) ) | ( (~ wire3338)  &  wire3230  &  (~ wire36324) ) ;
 assign wire3715 = ( (~ ng2631)  &  (~ ng2584)  &  ng2608  &  ng2599 ) ;
 assign wire3721 = ( (~ ng1890)  &  ng1914  &  (~ ng1937)  &  ng1905 ) ;
 assign wire3727 = ( ng1211  &  (~ ng1196)  &  (~ ng1243)  &  ng1220 ) ;
 assign wire3808 = ( wire3142  &  (~ wire34164)  &  (~ wire34165)  &  (~ wire34166) ) ;
 assign wire3815 = ( (~ ng15970)  &  ng22381 ) | ( (~ ng15970)  &  wire31236 ) | ( (~ ng15970)  &  (~ ng22381)  &  wire31235 ) ;
 assign wire3845 = ( ng3105  &  (~ wire3193)  &  (~ wire3247)  &  ng8430 ) ;
 assign wire3846 = ( (~ ng3128)  &  (~ ng8381)  &  (~ wire30893) ) ;
 assign wire3850 = ( (~ ng3135)  &  ng3099  &  ng8430  &  (~ wire30898) ) ;
 assign wire3851 = ( ng3106  &  (~ wire3247)  &  ng8430  &  (~ wire30899) ) ;
 assign wire3852 = ( ng3108  &  ng8430  &  (~ wire30902) ) ;
 assign wire3854 = ( (~ ng3135)  &  ng3103  &  ng8430  &  (~ wire30904) ) ;
 assign wire3855 = ( (~ ng3135)  &  ng3104  &  ng8430  &  (~ wire30903) ) ;
 assign wire3856 = ( ng3107  &  ng8430  &  (~ wire30905) ) ;
 assign wire3857 = ( (~ ng3139)  &  ng3147  &  (~ ng8381)  &  (~ wire30892) ) ;
 assign wire3858 = ( (~ ng3135)  &  ng3100  &  ng8430  &  (~ wire30900) ) ;
 assign wire3885 = ( ng12124  &  wire3230  &  (~ wire36289) ) | ( (~ wire3341)  &  wire3230  &  (~ wire36289) ) ;
 assign wire3886 = ( (~ ng2631)  &  (~ ng2584)  &  ng2607  &  ng2599 ) ;
 assign wire3893 = ( wire3141  &  wire9559 ) | ( wire3141  &  wire30886 ) | ( wire3141  &  wire35568 ) ;
 assign wire3894 = ( (~ ng1890)  &  ng1916  &  (~ ng1937)  &  ng1905 ) ;
 assign wire3902 = ( ng1211  &  (~ ng1196)  &  (~ ng1243)  &  ng1219 ) ;
 assign wire3931 = ( wire3142  &  (~ wire35515)  &  (~ wire35516)  &  (~ wire35517) ) ;
 assign wire4030 = ( (~ ng15970)  &  (~ wire32243)  &  (~ wire32244)  &  wire32245 ) ;
 assign wire4076 = ( ng321  &  (~ ng2257)  &  ng17051 ) | ( ng321  &  (~ ng17051)  &  ng23495 ) ;
 assign wire4080 = ( ng853  &  (~ ng2257)  &  (~ ng11935) ) | ( ng853  &  (~ ng17985)  &  (~ ng11935) ) | ( ng853  &  ng2257  &  (~ ng17985)  &  ng11935 ) ;
 assign wire4104 = ( ng11964  &  wire3230  &  (~ wire36188) ) | ( (~ wire3338)  &  wire3230  &  (~ wire36188) ) ;
 assign wire4105 = ( ng12329  &  wire3198  &  (~ wire36189) ) | ( (~ wire3338)  &  wire3198  &  (~ wire36189) ) ;
 assign wire4115 = ( (~ ng1890)  &  ng1912  &  (~ ng1937)  &  ng1905 ) ;
 assign wire4121 = ( ng1211  &  (~ ng1196)  &  ng1218  &  (~ ng1243) ) ;
 assign wire4133 = ( ng1312  &  wire4685 ) | ( ng1312  &  wire4686 ) | ( ng1312  &  wire4687 ) ;
 assign wire4135 = ( wire3221  &  (~ wire35515)  &  (~ wire35516)  &  (~ wire35517) ) ;
 assign wire4155 = ( ng823  &  wire35911 ) | ( ng823  &  wire35912 ) | ( ng823  &  wire35913 ) ;
 assign wire4214 = ( (~ ng13165)  &  ng22381 ) | ( (~ ng13165)  &  wire31236 ) | ( (~ ng13165)  &  (~ ng22381)  &  wire31235 ) ;
 assign wire4215 = ( ng823  &  (~ ng24676)  &  wire35876 ) | ( ng823  &  (~ ng24676)  &  wire35877 ) ;
 assign wire4217 = ( ng823  &  (~ ng2257)  &  (~ ng11935) ) | ( ng823  &  (~ ng17985)  &  (~ ng11935) ) | ( ng823  &  ng2257  &  (~ ng17985)  &  ng11935 ) ;
 assign wire4239 = ( ng1315  &  wire30883 ) | ( ng1315  &  ng21851  &  wire30881 ) ;
 assign wire4250 = ( (~ pg3234)  &  (~ ng3018) ) | ( (~ pg3234)  &  ng3036 ) ;
 assign wire4254 = ( ng12008  &  wire3230  &  (~ wire36171) ) | ( (~ wire3341)  &  wire3230  &  (~ wire36171) ) ;
 assign wire4255 = ( ng11965  &  wire3198  &  (~ wire36172) ) | ( (~ wire3341)  &  wire3198  &  (~ wire36172) ) ;
 assign wire4265 = ( (~ ng1890)  &  ng1913  &  (~ ng1937)  &  ng1905 ) ;
 assign wire4271 = ( ng1211  &  ng1217  &  (~ ng1196)  &  (~ ng1243) ) ;
 assign wire4282 = ( ng1315  &  wire4685 ) | ( ng1315  &  wire4686 ) | ( ng1315  &  wire4687 ) ;
 assign wire4284 = ( wire3220  &  (~ wire35515)  &  (~ wire35516)  &  (~ wire35517) ) ;
 assign wire4286 = ( ng2563  &  ng2562  &  ng2561 ) ;
 assign wire4287 = ( (~ ng1309)  &  ng2562  &  ng2561 ) ;
 assign wire4288 = ( (~ ng1315)  &  ng2563  &  ng2561 ) ;
 assign wire4291 = ( (~ ng1312)  &  (~ ng1309)  &  ng2562 ) ;
 assign wire4292 = ( (~ ng1315)  &  (~ ng1309)  &  ng2561 ) ;
 assign wire4302 = ( ng23521  &  wire6720  &  wire36140 ) | ( ng23521  &  wire34440  &  wire36140 ) ;
 assign wire4305 = ( (~ wire33770)  &  (~ wire33771)  &  (~ wire33772)  &  wire36145 ) ;
 assign wire4306 = ( (~ wire33786)  &  (~ wire33787)  &  (~ wire33788)  &  wire36146 ) ;
 assign wire4309 = ( ng853  &  (~ ng2257)  &  (~ ng12121) ) | ( ng853  &  (~ ng12121)  &  (~ ng18325) ) | ( ng853  &  ng2257  &  ng12121  &  (~ ng18325) ) ;
 assign wire4315 = ( ng823  &  (~ ng2257)  &  (~ ng12057) ) | ( ng823  &  (~ ng18218)  &  (~ ng12057) ) | ( ng823  &  ng2257  &  (~ ng18218)  &  ng12057 ) ;
 assign wire4319 = ( (~ ng28556)  &  (~ ng26918)  &  wire32701 ) | ( (~ ng28556)  &  (~ ng26918)  &  wire32702 ) ;
 assign wire4320 = ( (~ ng28556)  &  ng26918  &  (~ wire32701)  &  (~ wire32702) ) ;
 assign wire4321 = ( wire3180  &  (~ wire32816)  &  (~ wire32817) ) ;
 assign wire4323 = ( ng826  &  wire35911 ) | ( ng826  &  wire35912 ) | ( ng826  &  wire35913 ) ;
 assign wire4345 = ( ng1164  &  ng1165  &  ng1166 ) ;
 assign wire4346 = ( (~ ng1312)  &  ng1165  &  ng1166 ) ;
 assign wire4347 = ( (~ ng1315)  &  ng1164  &  ng1166 ) ;
 assign wire4348 = ( (~ ng1309)  &  ng1164  &  ng1165 ) ;
 assign wire4349 = ( (~ ng1312)  &  (~ ng1315)  &  ng1166 ) ;
 assign wire4350 = ( (~ ng1312)  &  (~ ng1309)  &  ng1165 ) ;
 assign wire4351 = ( (~ ng1315)  &  (~ ng1309)  &  ng1164 ) ;
 assign wire4359 = ( ng11600  &  (~ wire36120)  &  wire36121 ) | ( (~ ng27729)  &  (~ wire36120)  &  wire36121 ) ;
 assign wire4360 = ( wire36120  &  wire36122 ) | ( (~ ng11600)  &  ng27729  &  wire36122 ) ;
 assign wire4376 = ( ng12043  &  wire3117  &  wire36111 ) | ( ng12043  &  ng12090  &  wire36111 ) | ( wire3117  &  (~ ng12090)  &  wire36111 ) ;
 assign wire4379 = ( pg3229  &  (~ wire36109)  &  (~ wire36110) ) ;
 assign wire4380 = ( ng1085  &  ng1075  &  (~ ng853) ) ;
 assign wire4381 = ( ng1075  &  ng1078  &  (~ ng826) ) ;
 assign wire4382 = ( ng1085  &  ng1078  &  (~ ng823) ) ;
 assign wire4383 = ( ng1085  &  ng1075  &  ng1078 ) ;
 assign wire4384 = ( ng1078  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire4385 = ( ng1085  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire4386 = ( ng1075  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire4397 = ( ng797  &  wire32131 ) | ( ng797  &  ng27850  &  wire32130 ) ;
 assign wire4415 = ( wire6933  &  wire36083 ) | ( wire6934  &  wire36083 ) | ( wire34262  &  wire36083 ) ;
 assign wire4416 = ( ng18548  &  (~ wire34243)  &  (~ wire34244)  &  wire36084 ) ;
 assign wire4420 = ( (~ ng1309)  &  ng487  &  ng486 ) ;
 assign wire4425 = ( (~ ng1312)  &  (~ ng1309)  &  ng487 ) ;
 assign wire4426 = ( (~ ng1315)  &  (~ ng1309)  &  ng486 ) ;
 assign wire4432 = ( (~ ng15950)  &  ng22381 ) | ( (~ ng15950)  &  wire31236 ) | ( (~ ng15950)  &  (~ ng22381)  &  wire31235 ) ;
 assign wire4434 = ( ng853  &  (~ ng24676)  &  wire35876 ) | ( ng853  &  (~ ng24676)  &  wire35877 ) ;
 assign wire4436 = ( ng826  &  (~ ng2257)  &  (~ ng11935) ) | ( ng826  &  (~ ng17985)  &  (~ ng11935) ) | ( ng826  &  ng2257  &  (~ ng17985)  &  ng11935 ) ;
 assign wire4467 = ( ng1312  &  wire30883 ) | ( ng1312  &  ng21851  &  wire30881 ) ;
 assign wire4476 = ( (~ pg3234)  &  (~ wire35758)  &  wire36057 ) | ( (~ pg3234)  &  (~ wire35759)  &  wire36057 ) ;
 assign wire4477 = ( (~ pg3234)  &  (~ wire35758)  &  wire36058 ) | ( (~ pg3234)  &  (~ wire35759)  &  wire36058 ) ;
 assign wire4478 = ( (~ pg3234)  &  wire35758  &  wire35759 ) ;
 assign wire4479 = ( ng12271  &  wire3230  &  (~ wire36054) ) | ( (~ wire3338)  &  wire3230  &  (~ wire36054) ) ;
 assign wire4487 = ( (~ ng1890)  &  (~ ng1937)  &  ng1905  &  ng1910 ) ;
 assign wire4493 = ( ng1211  &  ng1216  &  (~ ng1196)  &  (~ ng1243) ) ;
 assign wire4506 = ( wire34390  &  wire36045 ) | ( ng21435  &  wire34389  &  wire36045 ) ;
 assign wire4560 = ( ng823  &  (~ ng2257)  &  (~ ng12121) ) | ( ng823  &  (~ ng12121)  &  (~ ng18325) ) | ( ng823  &  ng2257  &  ng12121  &  (~ ng18325) ) ;
 assign wire4568 = ( ng853  &  (~ ng24712)  &  wire35163 ) | ( ng853  &  (~ ng24712)  &  wire35164 ) ;
 assign wire4571 = ( ng826  &  wire4932 ) | ( ng826  &  wire35795 ) | ( ng826  &  wire35796 ) ;
 assign wire4588 = ( wire3142  &  (~ wire32534)  &  (~ wire32535)  &  (~ wire32536) ) ;
 assign wire4610 = ( (~ ng13165)  &  wire3353  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire4647 = ( ng12306  &  wire3230  &  (~ wire35957) ) | ( (~ wire3341)  &  wire3230  &  (~ wire35957) ) ;
 assign wire4648 = ( (~ ng2631)  &  (~ ng2584)  &  ng2599  &  ng2603 ) ;
 assign wire4654 = ( (~ ng1890)  &  ng1911  &  (~ ng1937)  &  ng1905 ) ;
 assign wire4662 = ( ng1211  &  ng1215  &  (~ ng1196)  &  (~ ng1243) ) ;
 assign wire4673 = ( wire3049  &  wire35840 ) | ( wire3049  &  wire35841 ) | ( wire3049  &  wire35845 ) ;
 assign wire4683 = ( ng1309  &  wire4685 ) | ( ng1309  &  wire4686 ) | ( ng1309  &  wire4687 ) ;
 assign wire4685 = ( (~ wire5231)  &  (~ wire5232)  &  (~ wire35551)  &  wire35932 ) ;
 assign wire4686 = ( (~ wire5231)  &  (~ wire5232)  &  (~ wire35551)  &  wire35934 ) ;
 assign wire4687 = ( (~ ng13055)  &  (~ wire33977)  &  (~ wire33978) ) ;
 assign wire4690 = ( ng2559  &  ng2539  &  ng2555 ) ;
 assign wire4691 = ( (~ ng1315)  &  ng2539  &  ng2555 ) ;
 assign wire4692 = ( (~ ng1309)  &  ng2559  &  ng2555 ) ;
 assign wire4695 = ( (~ ng1312)  &  (~ ng1309)  &  ng2559 ) ;
 assign wire4696 = ( (~ ng1315)  &  (~ ng1309)  &  ng2555 ) ;
 assign wire4703 = ( wire32253  &  wire35915 ) | ( ng21346  &  wire32252  &  wire35915 ) ;
 assign wire4708 = ( ng826  &  (~ ng2257)  &  (~ ng12121) ) | ( ng826  &  (~ ng12121)  &  (~ ng18325) ) | ( ng826  &  ng2257  &  ng12121  &  (~ ng18325) ) ;
 assign wire4721 = ( ng823  &  wire4932 ) | ( ng823  &  wire35795 ) | ( ng823  &  wire35796 ) ;
 assign wire4722 = ( ng853  &  wire35911 ) | ( ng853  &  wire35912 ) | ( ng853  &  wire35913 ) ;
 assign wire4748 = ( wire3221  &  (~ wire32534)  &  (~ wire32535)  &  (~ wire32536) ) ;
 assign wire4757 = ( ng767  &  (~ ng17031)  &  (~ ng23513) ) ;
 assign wire4770 = ( ng484  &  ng464  &  ng480 ) ;
 assign wire4771 = ( (~ ng1315)  &  ng464  &  ng480 ) ;
 assign wire4772 = ( (~ ng1309)  &  ng484  &  ng480 ) ;
 assign wire4775 = ( (~ ng1312)  &  (~ ng1309)  &  ng484 ) ;
 assign wire4776 = ( (~ ng1315)  &  (~ ng1309)  &  ng480 ) ;
 assign wire4780 = ( ng826  &  (~ ng24676)  &  wire35876 ) | ( ng826  &  (~ ng24676)  &  wire35877 ) ;
 assign wire4784 = ( (~ ng15950)  &  wire3353  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire4807 = ( (~ pg3234)  &  (~ wire35758)  &  wire35866 ) | ( (~ pg3234)  &  (~ wire35759)  &  wire35866 ) ;
 assign wire4808 = ( (~ pg3234)  &  (~ wire35758)  &  wire35867 ) | ( (~ pg3234)  &  (~ wire35759)  &  wire35867 ) ;
 assign wire4809 = ( ng12184  &  wire3230  &  (~ wire35864) ) | ( (~ wire3338)  &  wire3230  &  (~ wire35864) ) ;
 assign wire4810 = ( (~ ng2631)  &  (~ ng2584)  &  ng2599  &  ng2606 ) ;
 assign wire4869 = ( ng1425  &  (~ ng1315)  &  ng1424 ) ;
 assign wire4872 = ( ng1425  &  ng1423  &  (~ ng1309) ) ;
 assign wire4873 = ( (~ ng1312)  &  (~ ng1315)  &  ng1424 ) ;
 assign wire4874 = ( ng1423  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire4875 = ( ng1425  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire4888 = ( (~ ng21851)  &  wire3138  &  (~ wire34028)  &  wire35802 ) ;
 assign wire4889 = ( (~ ng21851)  &  wire3138  &  (~ wire34028)  &  wire35806 ) ;
 assign wire4918 = ( (~ ng13165)  &  (~ wire33906)  &  (~ wire33907)  &  wire35395 ) ;
 assign wire4928 = ( ng853  &  wire4932 ) | ( ng853  &  wire35795 ) | ( ng853  &  wire35796 ) ;
 assign wire4932 = ( wire3180  &  (~ wire32828)  &  (~ wire32829) ) ;
 assign wire4947 = ( (~ ng1339)  &  wire35792 ) | ( (~ ng1319)  &  wire35792 ) | ( (~ wire32567)  &  wire35792 ) ;
 assign wire4955 = ( wire3220  &  (~ wire32534)  &  (~ wire32535)  &  (~ wire32536) ) ;
 assign wire4961 = ( (~ ng28529)  &  (~ ng11647)  &  wire31817  &  wire35777 ) ;
 assign wire4964 = ( ng813  &  wire32131 ) | ( ng813  &  ng27850  &  wire32130 ) ;
 assign wire4975 = ( wire3220  &  (~ wire34164)  &  (~ wire34165)  &  (~ wire34166) ) ;
 assign wire4983 = ( ng323  &  (~ ng2257)  &  ng17051 ) | ( ng323  &  (~ ng17051)  &  ng23495 ) ;
 assign wire4985 = ( (~ ng15970)  &  wire3353  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire5013 = ( ng12233  &  wire3230  &  (~ wire35752) ) | ( (~ wire3341)  &  wire3230  &  (~ wire35752) ) ;
 assign wire5021 = ( ng2631  &  (~ ng2584)  &  ng30072 ) | ( ng2631  &  (~ ng2584)  &  wire35748 ) ;
 assign wire5029 = ( ng2812  &  ng2813  &  ng2811 ) ;
 assign wire5030 = ( (~ ng1309)  &  ng2813  &  ng2811 ) ;
 assign wire5031 = ( (~ ng1312)  &  ng2812  &  ng2811 ) ;
 assign wire5034 = ( (~ ng1312)  &  (~ ng1309)  &  ng2811 ) ;
 assign wire5035 = ( (~ ng1315)  &  (~ ng1309)  &  ng2813 ) ;
 assign wire5049 = ( (~ ng1890)  &  (~ ng1937)  &  ng1905  &  ng1909 ) ;
 assign wire5060 = ( wire3049  &  wire35694 ) | ( wire3049  &  wire35695 ) | ( wire3049  &  wire35699 ) ;
 assign wire5069 = ( ng2117  &  ng2119  &  ng2118 ) ;
 assign wire5070 = ( (~ ng1315)  &  ng2119  &  ng2118 ) ;
 assign wire5071 = ( (~ ng1312)  &  ng2117  &  ng2118 ) ;
 assign wire5072 = ( (~ ng1309)  &  ng2117  &  ng2119 ) ;
 assign wire5073 = ( (~ ng1312)  &  (~ ng1315)  &  ng2118 ) ;
 assign wire5074 = ( (~ ng1312)  &  (~ ng1309)  &  ng2117 ) ;
 assign wire5075 = ( (~ ng1315)  &  (~ ng1309)  &  ng2119 ) ;
 assign wire5088 = ( (~ ng1315)  &  ng2080  &  ng2079 ) ;
 assign wire5091 = ( ng2078  &  ng2080  &  (~ ng1309) ) ;
 assign wire5092 = ( (~ ng1312)  &  (~ ng1315)  &  ng2079 ) ;
 assign wire5093 = ( ng2078  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire5094 = ( (~ ng1315)  &  ng2080  &  (~ ng1309) ) ;
 assign wire5096 = ( (~ ng1309)  &  ng2093  &  ng2095 ) ;
 assign wire5101 = ( (~ ng1312)  &  (~ ng1309)  &  ng2093 ) ;
 assign wire5102 = ( (~ ng1315)  &  (~ ng1309)  &  ng2095 ) ;
 assign wire5104 = ( (~ ng1309)  &  ng2081  &  ng2083 ) ;
 assign wire5109 = ( (~ ng1312)  &  (~ ng1309)  &  ng2081 ) ;
 assign wire5110 = ( (~ ng1315)  &  (~ ng1309)  &  ng2083 ) ;
 assign wire5112 = ( ng2085  &  ng2086  &  ng2084 ) ;
 assign wire5113 = ( (~ ng1315)  &  ng2085  &  ng2086 ) ;
 assign wire5114 = ( (~ ng1309)  &  ng2086  &  ng2084 ) ;
 assign wire5117 = ( (~ ng1312)  &  (~ ng1309)  &  ng2084 ) ;
 assign wire5118 = ( (~ ng1315)  &  (~ ng1309)  &  ng2086 ) ;
 assign wire5120 = ( ng2104  &  (~ ng1309)  &  ng2102 ) ;
 assign wire5125 = ( (~ ng1312)  &  (~ ng1309)  &  ng2102 ) ;
 assign wire5126 = ( ng2104  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire5128 = ( ng2089  &  ng2087  &  ng2088 ) ;
 assign wire5129 = ( (~ ng1312)  &  ng2087  &  ng2088 ) ;
 assign wire5130 = ( (~ ng1315)  &  ng2089  &  ng2088 ) ;
 assign wire5131 = ( (~ ng1309)  &  ng2089  &  ng2087 ) ;
 assign wire5132 = ( (~ ng1312)  &  (~ ng1315)  &  ng2088 ) ;
 assign wire5133 = ( (~ ng1312)  &  (~ ng1309)  &  ng2087 ) ;
 assign wire5134 = ( (~ ng1315)  &  (~ ng1309)  &  ng2089 ) ;
 assign wire5136 = ( (~ ng1315)  &  ng2091  &  ng2092 ) ;
 assign wire5141 = ( ng2090  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire5142 = ( (~ ng1315)  &  (~ ng1309)  &  ng2092 ) ;
 assign wire5144 = ( ng2113  &  ng2111  &  ng2112 ) ;
 assign wire5145 = ( (~ ng1312)  &  ng2111  &  ng2112 ) ;
 assign wire5146 = ( (~ ng1315)  &  ng2113  &  ng2112 ) ;
 assign wire5147 = ( ng2113  &  (~ ng1309)  &  ng2111 ) ;
 assign wire5148 = ( (~ ng1312)  &  (~ ng1315)  &  ng2112 ) ;
 assign wire5149 = ( (~ ng1312)  &  (~ ng1309)  &  ng2111 ) ;
 assign wire5150 = ( (~ ng1315)  &  ng2113  &  (~ ng1309) ) ;
 assign wire5152 = ( ng2096  &  ng2098  &  ng2097 ) ;
 assign wire5153 = ( (~ ng1315)  &  ng2098  &  ng2097 ) ;
 assign wire5154 = ( (~ ng1312)  &  ng2096  &  ng2097 ) ;
 assign wire5155 = ( (~ ng1309)  &  ng2096  &  ng2098 ) ;
 assign wire5156 = ( (~ ng1312)  &  (~ ng1315)  &  ng2097 ) ;
 assign wire5157 = ( (~ ng1312)  &  (~ ng1309)  &  ng2096 ) ;
 assign wire5158 = ( (~ ng1315)  &  (~ ng1309)  &  ng2098 ) ;
 assign wire5160 = ( ng2107  &  ng2105  &  ng2106 ) ;
 assign wire5161 = ( (~ ng1309)  &  ng2107  &  ng2105 ) ;
 assign wire5162 = ( (~ ng1312)  &  ng2105  &  ng2106 ) ;
 assign wire5165 = ( (~ ng1312)  &  (~ ng1309)  &  ng2105 ) ;
 assign wire5166 = ( (~ ng1315)  &  (~ ng1309)  &  ng2107 ) ;
 assign wire5168 = ( ng2100  &  ng2099  &  ng2101 ) ;
 assign wire5169 = ( (~ ng1309)  &  ng2099  &  ng2101 ) ;
 assign wire5170 = ( (~ ng1315)  &  ng2100  &  ng2101 ) ;
 assign wire5173 = ( (~ ng1312)  &  (~ ng1309)  &  ng2099 ) ;
 assign wire5174 = ( (~ ng1315)  &  (~ ng1309)  &  ng2101 ) ;
 assign wire5176 = ( wire3224  &  ng11830  &  (~ wire35564) ) | ( wire3224  &  (~ wire3336)  &  (~ wire35564) ) ;
 assign wire5177 = ( ng12195  &  wire3140  &  (~ wire35565) ) | ( wire3140  &  (~ wire3336)  &  (~ wire35565) ) ;
 assign wire5199 = ( ng18639  &  (~ wire35462)  &  (~ wire35463)  &  wire35519 ) ;
 assign wire5200 = ( wire5231  &  wire35554 ) | ( wire5232  &  wire35554 ) | ( wire35551  &  wire35554 ) ;
 assign wire5202 = ( (~ ng2661)  &  (~ ng2664)  &  (~ ng185)  &  (~ ng2667) ) ;
 assign wire5203 = ( (~ ng1315)  &  (~ ng2661)  &  (~ ng2664)  &  (~ ng185) ) ;
 assign wire5204 = ( (~ ng1312)  &  (~ ng2661)  &  (~ ng185)  &  (~ ng2667) ) ;
 assign wire5205 = ( (~ ng1309)  &  (~ ng2664)  &  (~ ng185)  &  (~ ng2667) ) ;
 assign wire5206 = ( wire34948  &  wire35473 ) | ( wire34949  &  wire35473 ) ;
 assign wire5210 = ( (~ ng2598)  &  (~ ng2661)  &  (~ ng2664)  &  (~ ng2667) ) ;
 assign wire5211 = ( (~ ng1315)  &  (~ ng2598)  &  (~ ng2661)  &  (~ ng2664) ) ;
 assign wire5212 = ( (~ ng1312)  &  (~ ng2598)  &  (~ ng2661)  &  (~ ng2667) ) ;
 assign wire5213 = ( (~ ng1309)  &  (~ ng2598)  &  (~ ng2664)  &  (~ ng2667) ) ;
 assign wire5214 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2661)  &  (~ ng185) ) ;
 assign wire5216 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2598)  &  (~ ng2661) ) ;
 assign wire5217 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng185)  &  (~ ng2667) ) ;
 assign wire5219 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2598)  &  (~ ng2667) ) ;
 assign wire5220 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2664)  &  (~ ng185) ) ;
 assign wire5222 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2598)  &  (~ ng2664) ) ;
 assign wire5223 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire5224 = ( wire3049  &  wire34948 ) | ( wire3049  &  wire34949 ) ;
 assign wire5225 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng2598) ) ;
 assign wire5226 = ( (~ wire35408)  &  (~ wire35409)  &  wire35521  &  wire35522 ) ;
 assign wire5227 = ( wire35408  &  wire35524  &  wire35525 ) | ( wire35409  &  wire35524  &  wire35525 ) ;
 assign wire5228 = ( wire35408  &  wire35527  &  wire35528 ) | ( wire35409  &  wire35527  &  wire35528 ) ;
 assign wire5229 = ( wire3945  &  (~ wire35408)  &  (~ wire35409)  &  wire35530 ) ;
 assign wire5230 = ( wire3351  &  (~ wire35428)  &  (~ wire35429)  &  wire35532 ) ;
 assign wire5231 = ( (~ ng10822)  &  (~ wire35462)  &  (~ wire35463)  &  wire35534 ) ;
 assign wire5232 = ( ng10839  &  (~ wire35462)  &  (~ wire35463)  &  wire35536 ) ;
 assign wire5237 = ( (~ wire34008)  &  (~ wire34009)  &  wire35542 ) ;
 assign wire5238 = ( wire3351  &  wire3945  &  wire35430 ) ;
 assign wire5239 = ( wire3352  &  wire3926  &  wire35442 ) ;
 assign wire5244 = ( wire3352  &  wire3945  &  (~ wire34008)  &  (~ wire34009) ) ;
 assign wire5245 = ( wire3351  &  wire3926  &  wire35440 ) | ( wire3351  &  wire3926  &  wire35441 ) ;
 assign wire5248 = ( (~ ng1312)  &  (~ ng2428)  &  (~ ng2424) ) ;
 assign wire5251 = ( (~ ng2426)  &  (~ ng1309)  &  (~ ng2428) ) ;
 assign wire5252 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2424) ) ;
 assign wire5253 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2428) ) ;
 assign wire5254 = ( (~ ng2426)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire5256 = ( (~ ng2439)  &  (~ ng2443)  &  (~ ng2441) ) ;
 assign wire5257 = ( (~ ng1309)  &  (~ ng2443)  &  (~ ng2441) ) ;
 assign wire5258 = ( (~ ng1315)  &  (~ ng2439)  &  (~ ng2441) ) ;
 assign wire5261 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2443) ) ;
 assign wire5262 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2441) ) ;
 assign wire5264 = ( (~ ng1312)  &  (~ ng2458)  &  (~ ng2454) ) ;
 assign wire5267 = ( (~ ng2456)  &  (~ ng1309)  &  (~ ng2458) ) ;
 assign wire5268 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2454) ) ;
 assign wire5269 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2458) ) ;
 assign wire5270 = ( (~ ng2456)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire5272 = ( (~ ng2399)  &  (~ ng2469)  &  (~ ng2471) ) ;
 assign wire5273 = ( (~ ng1315)  &  (~ ng2469)  &  (~ ng2471) ) ;
 assign wire5274 = ( (~ ng1312)  &  (~ ng2399)  &  (~ ng2469) ) ;
 assign wire5275 = ( (~ ng1309)  &  (~ ng2399)  &  (~ ng2471) ) ;
 assign wire5276 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2469) ) ;
 assign wire5277 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2399) ) ;
 assign wire5278 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2471) ) ;
 assign wire5286 = ( (~ ng24723)  &  (~ ng23533)  &  wire35397 ) | ( (~ ng24723)  &  (~ ng23521)  &  wire35397 ) ;
 assign wire5287 = ( ng11687  &  ng11653  &  (~ ng11678)  &  (~ ng24723) ) ;
 assign wire5288 = ( (~ ng15950)  &  (~ wire33906)  &  (~ wire33907)  &  wire35395 ) ;
 assign wire5303 = ( ng1501  &  wire32947 ) | ( ng1501  &  ng27875  &  wire32946 ) ;
 assign wire5326 = ( ng801  &  wire32131 ) | ( ng801  &  ng27850  &  wire32130 ) ;
 assign wire5335 = ( wire3221  &  (~ wire34164)  &  (~ wire34165)  &  (~ wire34166) ) ;
 assign wire5341 = ( ng322  &  (~ ng2257)  &  ng17051 ) | ( ng322  &  (~ ng17051)  &  ng23495 ) ;
 assign wire5351 = ( ng113  &  wire31274 ) | ( ng113  &  ng27834  &  wire31273 ) ;
 assign wire5356 = ( ng97  &  wire31274 ) | ( ng97  &  ng27834  &  wire31273 ) ;
 assign wire5370 = ( wire3224  &  ng11863  &  (~ wire35367) ) | ( wire3224  &  (~ wire3339)  &  (~ wire35367) ) ;
 assign wire5371 = ( wire3140  &  ng11831  &  (~ wire35368) ) | ( wire3140  &  (~ wire3339)  &  (~ wire35368) ) ;
 assign wire5382 = ( wire3221  &  (~ wire35273)  &  (~ wire35274)  &  (~ wire35275) ) ;
 assign wire5419 = ( ng1858  &  (~ ng1315)  &  ng1860 ) ;
 assign wire5422 = ( ng1858  &  ng1859  &  (~ ng1309) ) ;
 assign wire5423 = ( (~ ng1312)  &  (~ ng1315)  &  ng1860 ) ;
 assign wire5424 = ( ng1859  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire5425 = ( ng1858  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire5435 = ( (~ ng15970)  &  (~ wire33053)  &  (~ wire33054)  &  wire35160 ) ;
 assign wire5442 = ( ng12107  &  ng12162  &  wire35347 ) | ( ng12107  &  (~ wire3122)  &  wire35347 ) | ( (~ ng12162)  &  (~ wire3122)  &  wire35347 ) ;
 assign wire5443 = ( (~ pg3229)  &  ng12162  &  (~ wire33008)  &  (~ wire33009) ) ;
 assign wire5445 = ( pg3229  &  (~ wire34927)  &  (~ wire34928) ) ;
 assign wire5464 = ( (~ ng15950)  &  ng22396 ) | ( (~ ng15950)  &  wire32093 ) | ( (~ ng15950)  &  (~ ng22396)  &  wire32092 ) ;
 assign wire5469 = ( ng853  &  wire5902 ) | ( ng853  &  wire5903 ) | ( ng853  &  wire35144 ) ;
 assign wire5475 = ( (~ ng633)  &  wire35346 ) | ( (~ ng640)  &  wire35346 ) | ( (~ wire31592)  &  wire35346 ) ;
 assign wire5492 = ( wire3142  &  (~ wire35273)  &  (~ wire35274)  &  (~ wire35275) ) ;
 assign wire5512 = ( ng2165  &  wire33795 ) | ( ng2165  &  ng27892  &  wire33794 ) ;
 assign wire5525 = ( ng2026  &  wire33413  &  wire33414  &  wire35337 ) ;
 assign wire5526 = ( (~ ng2026)  &  wire35338 ) | ( (~ wire33413)  &  wire35338 ) | ( (~ wire33414)  &  wire35338 ) ;
 assign wire5527 = ( wire3220  &  (~ wire33231)  &  (~ wire33232)  &  (~ wire33233) ) ;
 assign wire5557 = ( wire3142  &  (~ wire32387)  &  (~ wire32388)  &  (~ wire32389) ) ;
 assign wire5564 = ( (~ ng13165)  &  ng22396 ) | ( (~ ng13165)  &  wire32093 ) | ( (~ ng13165)  &  (~ ng22396)  &  wire32092 ) ;
 assign wire5571 = ( ng17086  &  ng27850  &  wire3235 ) | ( (~ ng23511)  &  ng27850  &  wire3235 ) ;
 assign wire5572 = ( (~ wire32122)  &  (~ wire32123)  &  (~ wire32124)  &  wire35325 ) ;
 assign wire5573 = ( (~ wire32106)  &  (~ wire32107)  &  (~ wire32108)  &  wire35326 ) ;
 assign wire5577 = ( (~ ng2257)  &  wire35320 ) | ( (~ ng23511)  &  wire35320 ) ;
 assign wire5605 = ( wire3224  &  ng11938  &  (~ wire35309) ) | ( wire3224  &  (~ wire3339)  &  (~ wire35309) ) ;
 assign wire5606 = ( (~ ng557)  &  (~ ng510)  &  ng525  &  ng533 ) ;
 assign wire5619 = ( ng2396  &  (~ ng2257)  &  ng17151 ) | ( ng2396  &  ng23537  &  (~ ng17151) ) ;
 assign wire5626 = ( ng2147  &  (~ ng17031)  &  (~ ng23539) ) ;
 assign wire5673 = ( (~ ng13165)  &  (~ wire33053)  &  (~ wire33054)  &  wire35160 ) ;
 assign wire5694 = ( wire3221  &  (~ wire32387)  &  (~ wire32388)  &  (~ wire32389) ) ;
 assign wire5702 = ( ng853  &  (~ ng2257)  &  (~ ng11988) ) | ( ng853  &  (~ ng18102)  &  (~ ng11988) ) | ( ng853  &  ng2257  &  (~ ng18102)  &  ng11988 ) ;
 assign wire5707 = ( ng826  &  wire5902 ) | ( ng826  &  wire5903 ) | ( ng826  &  wire35144 ) ;
 assign wire5726 = ( ng121  &  wire31274 ) | ( ng121  &  ng27834  &  wire31273 ) ;
 assign wire5739 = ( wire3224  &  ng11896  &  (~ wire35277) ) | ( wire3224  &  (~ wire3336)  &  (~ wire35277) ) ;
 assign wire5740 = ( (~ ng557)  &  (~ ng510)  &  ng525  &  ng534 ) ;
 assign wire5749 = ( wire3220  &  (~ wire35273)  &  (~ wire35274)  &  (~ wire35275) ) ;
 assign wire5751 = ( (~ ng1312)  &  (~ ng2670)  &  (~ ng2676)  &  (~ ng185) ) ;
 assign wire5752 = ( (~ ng2670)  &  (~ ng2676)  &  (~ ng2673)  &  (~ ng185) ) ;
 assign wire5753 = ( (~ ng1315)  &  (~ ng2670)  &  (~ ng2673)  &  (~ ng185) ) ;
 assign wire5754 = ( (~ ng1309)  &  (~ ng2676)  &  (~ ng2673)  &  (~ ng185) ) ;
 assign wire5755 = ( wire35228  &  wire35231 ) | ( wire35229  &  wire35231 ) ;
 assign wire5759 = ( (~ ng2616)  &  (~ ng1312)  &  (~ ng2670)  &  (~ ng2676) ) ;
 assign wire5760 = ( (~ ng2616)  &  (~ ng2670)  &  (~ ng2676)  &  (~ ng2673) ) ;
 assign wire5761 = ( (~ ng2616)  &  (~ ng1315)  &  (~ ng2670)  &  (~ ng2673) ) ;
 assign wire5762 = ( (~ ng2616)  &  (~ ng1309)  &  (~ ng2676)  &  (~ ng2673) ) ;
 assign wire5763 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2670)  &  (~ ng185) ) ;
 assign wire5765 = ( (~ ng2616)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng2670) ) ;
 assign wire5766 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2676)  &  (~ ng185) ) ;
 assign wire5768 = ( (~ ng2616)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng2676) ) ;
 assign wire5769 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2673)  &  (~ ng185) ) ;
 assign wire5771 = ( (~ ng2616)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng2673) ) ;
 assign wire5772 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire5774 = ( (~ ng2616)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire5775 = ( (~ ng1309)  &  (~ ng2564)  &  (~ ng2641) ) ;
 assign wire5780 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2564) ) ;
 assign wire5781 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2641) ) ;
 assign wire5787 = ( ng2398  &  (~ ng2257)  &  ng17151 ) | ( ng2398  &  ng23537  &  (~ ng17151) ) ;
 assign wire5793 = ( (~ ng12224)  &  wire35208 ) | ( ng12179  &  wire3120  &  wire35208 ) | ( ng12179  &  ng12224  &  wire35208 ) ;
 assign wire5794 = ( (~ pg3229)  &  ng12224  &  (~ wire33860)  &  (~ wire33861) ) ;
 assign wire5795 = ( pg3229  &  (~ wire34421)  &  (~ wire34422) ) ;
 assign wire5804 = ( (~ ng28584)  &  ng26941  &  (~ wire33478)  &  (~ wire33479) ) ;
 assign wire5805 = ( ng2200  &  wire33795 ) | ( ng2200  &  ng27892  &  wire33794 ) ;
 assign wire5810 = ( ng2195  &  wire33795 ) | ( ng2195  &  ng27892  &  wire33794 ) ;
 assign wire5831 = ( ng1865  &  ng1845  &  ng1861 ) ;
 assign wire5832 = ( (~ ng1315)  &  ng1845  &  ng1861 ) ;
 assign wire5833 = ( (~ ng1309)  &  ng1865  &  ng1861 ) ;
 assign wire5836 = ( (~ ng1312)  &  (~ ng1309)  &  ng1865 ) ;
 assign wire5837 = ( (~ ng1315)  &  (~ ng1309)  &  ng1861 ) ;
 assign wire5849 = ( ng17124  &  ng27875  &  wire3234 ) | ( ng27875  &  wire3234  &  (~ ng23526) ) ;
 assign wire5850 = ( (~ wire32922)  &  (~ wire32923)  &  (~ wire32924)  &  wire35169 ) ;
 assign wire5851 = ( (~ wire32938)  &  (~ wire32939)  &  (~ wire32940)  &  wire35170 ) ;
 assign wire5854 = ( ng826  &  (~ ng24712)  &  wire35163 ) | ( ng826  &  (~ ng24712)  &  wire35164 ) ;
 assign wire5858 = ( (~ ng15950)  &  (~ wire33053)  &  (~ wire33054)  &  wire35160 ) ;
 assign wire5879 = ( wire3220  &  (~ wire32387)  &  (~ wire32388)  &  (~ wire32389) ) ;
 assign wire5883 = ( ng12152  &  ng12207  &  wire35150 ) | ( ng12152  &  wire3123  &  wire35150 ) | ( (~ ng12207)  &  wire3123  &  wire35150 ) ;
 assign wire5886 = ( pg3229  &  (~ wire32303)  &  (~ wire32304) ) ;
 assign wire5893 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire35146 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire35146 ) ;
 assign wire5894 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire35147 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire35147 ) ;
 assign wire5895 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire35148 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire35148 ) ;
 assign wire5899 = ( ng823  &  wire5902 ) | ( ng823  &  wire5903 ) | ( ng823  &  wire35144 ) ;
 assign wire5902 = ( (~ ng28529)  &  ng16655  &  wire31826 ) | ( (~ ng28529)  &  ng16655  &  wire31827 ) ;
 assign wire5903 = ( ng785  &  wire32131 ) | ( ng785  &  ng27850  &  wire32130 ) ;
 assign wire5963 = ( (~ ng28501)  &  (~ ng27462)  &  (~ wire30937)  &  (~ wire30938) ) ;
 assign wire5964 = ( (~ ng28501)  &  ng27462  &  wire30937 ) | ( (~ ng28501)  &  ng27462  &  wire30938 ) ;
 assign wire5965 = ( wire3175  &  (~ wire31201)  &  (~ wire31202) ) ;
 assign wire5973 = ( (~ ng28501)  &  ng26902  &  wire35043 ) ;
 assign wire5976 = ( ng117  &  wire31274 ) | ( ng117  &  ng27834  &  wire31273 ) ;
 assign wire5993 = ( wire3224  &  ng12035  &  (~ wire35023) ) | ( wire3224  &  (~ wire3339)  &  (~ wire35023) ) ;
 assign wire5994 = ( (~ ng557)  &  (~ ng510)  &  ng531  &  ng525 ) ;
 assign wire6005 = ( ng2720  &  wire34449  &  wire34450  &  wire35021 ) ;
 assign wire6006 = ( (~ ng2720)  &  wire35022 ) | ( (~ wire34449)  &  wire35022 ) | ( (~ wire34450)  &  wire35022 ) ;
 assign wire6015 = ( ng2397  &  (~ ng2257)  &  ng17151 ) | ( ng2397  &  ng23537  &  (~ ng17151) ) ;
 assign wire6043 = ( wire3220  &  (~ wire33296)  &  (~ wire33297)  &  (~ wire33298) ) ;
 assign wire6055 = ( ng1704  &  (~ ng2257)  &  ng17124 ) | ( ng1704  &  (~ ng17124)  &  ng23526 ) ;
 assign wire6057 = ( ng853  &  (~ ng2257)  &  (~ ng12057) ) | ( ng853  &  (~ ng18218)  &  (~ ng12057) ) | ( ng853  &  ng2257  &  (~ ng18218)  &  ng12057 ) ;
 assign wire6089 = ( ng1171  &  (~ ng1309)  &  ng1167 ) ;
 assign wire6094 = ( ng1171  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6095 = ( (~ ng1315)  &  (~ ng1309)  &  ng1167 ) ;
 assign wire6103 = ( ng1009  &  (~ ng2257)  &  ng17086 ) | ( ng1009  &  (~ ng17086)  &  ng23511 ) ;
 assign wire6105 = ( ng826  &  wire8487 ) | ( ng826  &  wire3150  &  wire32248 ) ;
 assign wire6107 = ( ng826  &  (~ ng2257)  &  (~ ng11988) ) | ( ng826  &  (~ ng18102)  &  (~ ng11988) ) | ( ng826  &  ng2257  &  (~ ng18102)  &  ng11988 ) ;
 assign wire6114 = ( ng11902  &  wire3930  &  (~ ng11807)  &  (~ wire32226) ) ;
 assign wire6138 = ( ng1309  &  wire6925 ) | ( ng1309  &  wire6926 ) | ( ng1309  &  wire6927 ) ;
 assign wire6140 = ( wire3220  &  (~ wire31587)  &  (~ wire31588)  &  (~ wire31589) ) ;
 assign wire6155 = ( ng79  &  (~ ng17031)  &  (~ ng23497) ) ;
 assign wire6170 = ( (~ ng3135)  &  ng3092  &  ng8430  &  (~ wire30903) ) ;
 assign wire6171 = ( ng3093  &  (~ wire3193)  &  (~ wire3247)  &  ng8430 ) ;
 assign wire6175 = ( (~ ng3135)  &  ng3091  &  ng8430  &  (~ wire30904) ) ;
 assign wire6176 = ( (~ ng3135)  &  ng3085  &  ng8430  &  (~ wire30900) ) ;
 assign wire6177 = ( (~ ng3135)  &  ng3084  &  ng8430  &  (~ wire30898) ) ;
 assign wire6178 = ( ng3094  &  (~ wire3247)  &  ng8430  &  (~ wire30899) ) ;
 assign wire6179 = ( ng3096  &  ng8430  &  (~ wire30902) ) ;
 assign wire6180 = ( ng3095  &  ng8430  &  (~ wire30905) ) ;
 assign wire6188 = ( ng1309  &  wire30883 ) | ( (~ ng1186)  &  ng1309  &  ng21851 ) ;
 assign wire6190 = ( wire3224  &  (~ wire3336)  &  (~ wire34962) ) | ( wire3224  &  ng11979  &  (~ wire34962) ) ;
 assign wire6207 = ( ng2554  &  ng2553  &  ng2552 ) ;
 assign wire6208 = ( (~ ng1309)  &  ng2553  &  ng2552 ) ;
 assign wire6209 = ( (~ ng1315)  &  ng2554  &  ng2552 ) ;
 assign wire6212 = ( (~ ng1312)  &  (~ ng1309)  &  ng2553 ) ;
 assign wire6213 = ( (~ ng1315)  &  (~ ng1309)  &  ng2552 ) ;
 assign wire6217 = ( (~ ng2647)  &  (~ ng2645)  &  (~ ng2643) ) ;
 assign wire6218 = ( (~ ng1312)  &  (~ ng2647)  &  (~ ng2643) ) ;
 assign wire6219 = ( (~ ng1315)  &  (~ ng2645)  &  (~ ng2643) ) ;
 assign wire6220 = ( (~ ng1309)  &  (~ ng2647)  &  (~ ng2645) ) ;
 assign wire6221 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2643) ) ;
 assign wire6222 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2647) ) ;
 assign wire6223 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2645) ) ;
 assign wire6240 = ( ng2185  &  wire33795 ) | ( ng2185  &  ng27892  &  wire33794 ) ;
 assign wire6255 = ( wire3221  &  (~ wire33296)  &  (~ wire33297)  &  (~ wire33298) ) ;
 assign wire6263 = ( ng1703  &  (~ ng2257)  &  ng17124 ) | ( ng1703  &  (~ ng17124)  &  ng23526 ) ;
 assign wire6278 = ( ng1769  &  ng1772  &  (~ ng826) ) ;
 assign wire6281 = ( ng1769  &  ng1779  &  (~ ng853) ) ;
 assign wire6282 = ( ng1772  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire6283 = ( ng1779  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire6284 = ( ng1769  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire6292 = ( ng1471  &  wire32947 ) | ( ng1471  &  ng27875  &  wire32946 ) ;
 assign wire6301 = ( wire34893  &  wire34898 ) | ( wire34894  &  wire34898 ) | ( wire34895  &  wire34898 ) ;
 assign wire6302 = ( wire34893  &  wire34900 ) | ( wire34894  &  wire34900 ) | ( wire34895  &  wire34900 ) ;
 assign wire6303 = ( wire34893  &  wire34902 ) | ( wire34894  &  wire34902 ) | ( wire34895  &  wire34902 ) ;
 assign wire6304 = ( wire34893  &  wire34904 ) | ( wire34894  &  wire34904 ) | ( wire34895  &  wire34904 ) ;
 assign wire6305 = ( wire34893  &  wire34905 ) | ( wire34894  &  wire34905 ) | ( wire34895  &  wire34905 ) ;
 assign wire6306 = ( wire34893  &  wire34906 ) | ( wire34894  &  wire34906 ) | ( wire34895  &  wire34906 ) ;
 assign wire6307 = ( wire34893  &  wire34907 ) | ( wire34894  &  wire34907 ) | ( wire34895  &  wire34907 ) ;
 assign wire6308 = ( wire3049  &  wire34893 ) | ( wire3049  &  wire34894 ) | ( wire3049  &  wire34895 ) ;
 assign wire6329 = ( ng1396  &  ng1398  &  ng1397 ) ;
 assign wire6330 = ( (~ ng1315)  &  ng1398  &  ng1397 ) ;
 assign wire6331 = ( (~ ng1312)  &  ng1396  &  ng1397 ) ;
 assign wire6332 = ( (~ ng1309)  &  ng1396  &  ng1398 ) ;
 assign wire6333 = ( (~ ng1312)  &  (~ ng1315)  &  ng1397 ) ;
 assign wire6334 = ( (~ ng1312)  &  (~ ng1309)  &  ng1396 ) ;
 assign wire6335 = ( (~ ng1315)  &  (~ ng1309)  &  ng1398 ) ;
 assign wire6337 = ( ng1404  &  ng1402  &  (~ ng1309) ) ;
 assign wire6342 = ( (~ ng1312)  &  ng1402  &  (~ ng1309) ) ;
 assign wire6343 = ( ng1404  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6345 = ( ng1389  &  ng1387  &  ng1388 ) ;
 assign wire6346 = ( (~ ng1312)  &  ng1387  &  ng1388 ) ;
 assign wire6347 = ( (~ ng1315)  &  ng1389  &  ng1388 ) ;
 assign wire6348 = ( (~ ng1309)  &  ng1389  &  ng1387 ) ;
 assign wire6349 = ( (~ ng1312)  &  (~ ng1315)  &  ng1388 ) ;
 assign wire6350 = ( (~ ng1312)  &  (~ ng1309)  &  ng1387 ) ;
 assign wire6351 = ( (~ ng1315)  &  (~ ng1309)  &  ng1389 ) ;
 assign wire6353 = ( ng1392  &  (~ ng1309)  &  ng1390 ) ;
 assign wire6358 = ( (~ ng1312)  &  (~ ng1309)  &  ng1390 ) ;
 assign wire6359 = ( ng1392  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6361 = ( ng1409  &  ng1410  &  ng1408 ) ;
 assign wire6362 = ( (~ ng1309)  &  ng1410  &  ng1408 ) ;
 assign wire6363 = ( (~ ng1312)  &  ng1409  &  ng1408 ) ;
 assign wire6366 = ( (~ ng1312)  &  (~ ng1309)  &  ng1408 ) ;
 assign wire6367 = ( (~ ng1315)  &  (~ ng1309)  &  ng1410 ) ;
 assign wire6369 = ( ng1384  &  ng1385  &  ng1386 ) ;
 assign wire6370 = ( (~ ng1315)  &  ng1385  &  ng1386 ) ;
 assign wire6371 = ( (~ ng1309)  &  ng1384  &  ng1386 ) ;
 assign wire6374 = ( (~ ng1312)  &  (~ ng1309)  &  ng1384 ) ;
 assign wire6375 = ( (~ ng1315)  &  (~ ng1309)  &  ng1386 ) ;
 assign wire6377 = ( ng1413  &  (~ ng1315)  &  ng1412 ) ;
 assign wire6380 = ( ng1411  &  ng1413  &  (~ ng1309) ) ;
 assign wire6381 = ( (~ ng1312)  &  (~ ng1315)  &  ng1412 ) ;
 assign wire6382 = ( ng1411  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6383 = ( ng1413  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6385 = ( ng1393  &  ng1395  &  ng1394 ) ;
 assign wire6386 = ( (~ ng1315)  &  ng1395  &  ng1394 ) ;
 assign wire6387 = ( (~ ng1312)  &  ng1393  &  ng1394 ) ;
 assign wire6388 = ( (~ ng1309)  &  ng1393  &  ng1395 ) ;
 assign wire6389 = ( (~ ng1312)  &  (~ ng1315)  &  ng1394 ) ;
 assign wire6390 = ( (~ ng1312)  &  (~ ng1309)  &  ng1393 ) ;
 assign wire6391 = ( (~ ng1315)  &  (~ ng1309)  &  ng1395 ) ;
 assign wire6393 = ( ng1400  &  ng1401  &  ng1399 ) ;
 assign wire6394 = ( (~ ng1309)  &  ng1401  &  ng1399 ) ;
 assign wire6395 = ( (~ ng1312)  &  ng1400  &  ng1399 ) ;
 assign wire6398 = ( (~ ng1312)  &  (~ ng1309)  &  ng1399 ) ;
 assign wire6399 = ( (~ ng1315)  &  (~ ng1309)  &  ng1401 ) ;
 assign wire6401 = ( ng1406  &  ng1407  &  ng1405 ) ;
 assign wire6402 = ( (~ ng1309)  &  ng1407  &  ng1405 ) ;
 assign wire6403 = ( (~ ng1312)  &  ng1406  &  ng1405 ) ;
 assign wire6406 = ( (~ ng1312)  &  (~ ng1309)  &  ng1405 ) ;
 assign wire6407 = ( (~ ng1315)  &  (~ ng1309)  &  ng1407 ) ;
 assign wire6409 = ( ng1418  &  ng1417  &  ng1419 ) ;
 assign wire6410 = ( (~ ng1309)  &  ng1417  &  ng1419 ) ;
 assign wire6411 = ( (~ ng1315)  &  ng1418  &  ng1419 ) ;
 assign wire6414 = ( (~ ng1312)  &  (~ ng1309)  &  ng1417 ) ;
 assign wire6415 = ( (~ ng1315)  &  (~ ng1309)  &  ng1419 ) ;
 assign wire6424 = ( wire32469  &  wire34747 ) | ( wire32470  &  wire34747 ) | ( wire32471  &  wire34747 ) ;
 assign wire6425 = ( (~ ng13055)  &  (~ wire32292)  &  (~ wire32293) ) ;
 assign wire6434 = ( ng1010  &  (~ ng2257)  &  ng17086 ) | ( ng1010  &  (~ ng17086)  &  ng23511 ) ;
 assign wire6441 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34716 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34716 ) ;
 assign wire6442 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34719 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34719 ) ;
 assign wire6443 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34722 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34722 ) ;
 assign wire6444 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34725 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34725 ) ;
 assign wire6445 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34727 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34727 ) ;
 assign wire6446 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34729 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34729 ) ;
 assign wire6447 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34731 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34731 ) ;
 assign wire6448 = ( (~ ng12044)  &  ng18102  &  ng11988  &  wire34732 ) | ( ng12044  &  (~ ng18102)  &  (~ ng11988)  &  wire34732 ) ;
 assign wire6452 = ( ng823  &  (~ ng2257)  &  (~ ng11988) ) | ( ng823  &  (~ ng18102)  &  (~ ng11988) ) | ( ng823  &  ng2257  &  (~ ng18102)  &  ng11988 ) ;
 assign wire6459 = ( ng866  &  ng867  &  (~ ng853) ) ;
 assign wire6464 = ( ng866  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire6465 = ( (~ ng826)  &  ng867  &  (~ ng853) ) ;
 assign wire6468 = ( (~ ng1119)  &  (~ ng1116)  &  (~ ng853) ) ;
 assign wire6473 = ( (~ ng1116)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire6474 = ( (~ ng1119)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire6488 = ( ng809  &  wire32131 ) | ( ng809  &  ng27850  &  wire32130 ) ;
 assign wire6508 = ( ng1312  &  wire6925 ) | ( ng1312  &  wire6926 ) | ( ng1312  &  wire6927 ) ;
 assign wire6514 = ( ng479  &  ng478  &  ng477 ) ;
 assign wire6515 = ( (~ ng1309)  &  ng478  &  ng477 ) ;
 assign wire6516 = ( (~ ng1315)  &  ng479  &  ng477 ) ;
 assign wire6519 = ( (~ ng1312)  &  (~ ng1309)  &  ng478 ) ;
 assign wire6520 = ( (~ ng1315)  &  (~ ng1309)  &  ng477 ) ;
 assign wire6532 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34642 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34642 ) ;
 assign wire6533 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34645 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34645 ) ;
 assign wire6534 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34648 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34648 ) ;
 assign wire6535 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34651 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34651 ) ;
 assign wire6536 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34653 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34653 ) ;
 assign wire6537 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34655 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34655 ) ;
 assign wire6538 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34657 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34657 ) ;
 assign wire6539 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire34658 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire34658 ) ;
 assign wire6544 = ( (~ ng12026)  &  wire34638 ) | ( ng11974  &  ng12026  &  wire34638 ) | ( ng11974  &  (~ wire3121)  &  wire34638 ) ;
 assign wire6545 = ( (~ pg3229)  &  ng12026  &  (~ wire31334)  &  (~ wire31335) ) ;
 assign wire6546 = ( pg3229  &  (~ wire34636)  &  (~ wire34637) ) ;
 assign wire6547 = ( ng388  &  ng398  &  (~ ng853) ) ;
 assign wire6552 = ( ng398  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire6553 = ( ng388  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire6564 = ( ng3110  &  (~ wire3246)  &  (~ ng8381)  &  (~ wire30892) ) ;
 assign wire6572 = ( wire3224  &  ng12146  &  (~ wire34619) ) | ( wire3224  &  (~ wire3339)  &  (~ wire34619) ) ;
 assign wire6581 = ( wire34598  &  wire34603 ) | ( wire34599  &  wire34603 ) | ( wire34600  &  wire34603 ) ;
 assign wire6582 = ( wire34598  &  wire34605 ) | ( wire34599  &  wire34605 ) | ( wire34600  &  wire34605 ) ;
 assign wire6583 = ( wire34598  &  wire34607 ) | ( wire34599  &  wire34607 ) | ( wire34600  &  wire34607 ) ;
 assign wire6584 = ( wire34598  &  wire34609 ) | ( wire34599  &  wire34609 ) | ( wire34600  &  wire34609 ) ;
 assign wire6585 = ( wire34598  &  wire34610 ) | ( wire34599  &  wire34610 ) | ( wire34600  &  wire34610 ) ;
 assign wire6586 = ( wire34598  &  wire34611 ) | ( wire34599  &  wire34611 ) | ( wire34600  &  wire34611 ) ;
 assign wire6587 = ( wire34598  &  wire34612 ) | ( wire34599  &  wire34612 ) | ( wire34600  &  wire34612 ) ;
 assign wire6588 = ( wire3049  &  wire34598 ) | ( wire3049  &  wire34599 ) | ( wire3049  &  wire34600 ) ;
 assign wire6609 = ( (~ ng1315)  &  ng2773  &  ng2774 ) ;
 assign wire6614 = ( ng2772  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6615 = ( (~ ng1315)  &  (~ ng1309)  &  ng2774 ) ;
 assign wire6617 = ( ng2779  &  ng2778  &  ng2780 ) ;
 assign wire6618 = ( (~ ng1309)  &  ng2778  &  ng2780 ) ;
 assign wire6619 = ( (~ ng1315)  &  ng2779  &  ng2780 ) ;
 assign wire6622 = ( (~ ng1312)  &  (~ ng1309)  &  ng2778 ) ;
 assign wire6623 = ( (~ ng1315)  &  (~ ng1309)  &  ng2780 ) ;
 assign wire6625 = ( ng2799  &  ng2801  &  ng2800 ) ;
 assign wire6626 = ( (~ ng1315)  &  ng2801  &  ng2800 ) ;
 assign wire6627 = ( (~ ng1312)  &  ng2799  &  ng2800 ) ;
 assign wire6628 = ( (~ ng1309)  &  ng2799  &  ng2801 ) ;
 assign wire6629 = ( (~ ng1312)  &  (~ ng1315)  &  ng2800 ) ;
 assign wire6630 = ( (~ ng1312)  &  (~ ng1309)  &  ng2799 ) ;
 assign wire6631 = ( (~ ng1315)  &  (~ ng1309)  &  ng2801 ) ;
 assign wire6633 = ( (~ ng1315)  &  ng2806  &  ng2807 ) ;
 assign wire6638 = ( ng2805  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6639 = ( (~ ng1315)  &  (~ ng1309)  &  ng2807 ) ;
 assign wire6641 = ( ng2786  &  (~ ng1315)  &  ng2785 ) ;
 assign wire6644 = ( ng2786  &  ng2784  &  (~ ng1309) ) ;
 assign wire6645 = ( (~ ng1312)  &  (~ ng1315)  &  ng2785 ) ;
 assign wire6646 = ( ng2784  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6647 = ( ng2786  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6649 = ( (~ ng1309)  &  ng2796  &  ng2798 ) ;
 assign wire6654 = ( (~ ng1312)  &  (~ ng1309)  &  ng2796 ) ;
 assign wire6655 = ( (~ ng1315)  &  (~ ng1309)  &  ng2798 ) ;
 assign wire6657 = ( (~ ng1315)  &  ng2795  &  ng2794 ) ;
 assign wire6660 = ( ng2793  &  ng2795  &  (~ ng1309) ) ;
 assign wire6661 = ( (~ ng1312)  &  (~ ng1315)  &  ng2794 ) ;
 assign wire6662 = ( ng2793  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6663 = ( (~ ng1315)  &  ng2795  &  (~ ng1309) ) ;
 assign wire6665 = ( ng2777  &  ng2776  &  ng2775 ) ;
 assign wire6666 = ( (~ ng1312)  &  ng2776  &  ng2775 ) ;
 assign wire6667 = ( ng2777  &  (~ ng1309)  &  ng2775 ) ;
 assign wire6670 = ( (~ ng1312)  &  (~ ng1309)  &  ng2775 ) ;
 assign wire6671 = ( (~ ng1315)  &  ng2777  &  (~ ng1309) ) ;
 assign wire6673 = ( ng2783  &  ng2782  &  ng2781 ) ;
 assign wire6674 = ( (~ ng1312)  &  ng2782  &  ng2781 ) ;
 assign wire6675 = ( (~ ng1309)  &  ng2783  &  ng2781 ) ;
 assign wire6678 = ( (~ ng1312)  &  (~ ng1309)  &  ng2781 ) ;
 assign wire6679 = ( (~ ng1315)  &  (~ ng1309)  &  ng2783 ) ;
 assign wire6681 = ( ng2792  &  ng2790  &  ng2791 ) ;
 assign wire6682 = ( (~ ng1312)  &  ng2790  &  ng2791 ) ;
 assign wire6683 = ( (~ ng1315)  &  ng2792  &  ng2791 ) ;
 assign wire6684 = ( (~ ng1309)  &  ng2792  &  ng2790 ) ;
 assign wire6685 = ( (~ ng1312)  &  (~ ng1315)  &  ng2791 ) ;
 assign wire6686 = ( (~ ng1312)  &  (~ ng1309)  &  ng2790 ) ;
 assign wire6687 = ( (~ ng1315)  &  (~ ng1309)  &  ng2792 ) ;
 assign wire6689 = ( ng2787  &  ng2788  &  ng2789 ) ;
 assign wire6690 = ( (~ ng1315)  &  ng2788  &  ng2789 ) ;
 assign wire6691 = ( (~ ng1309)  &  ng2787  &  ng2789 ) ;
 assign wire6694 = ( (~ ng1312)  &  (~ ng1309)  &  ng2787 ) ;
 assign wire6695 = ( (~ ng1315)  &  (~ ng1309)  &  ng2789 ) ;
 assign wire6702 = ( (~ ng2727)  &  wire34453 ) | ( (~ ng2707)  &  wire34453 ) | ( (~ wire34450)  &  wire34453 ) ;
 assign wire6720 = ( (~ ng23533)  &  wire34435 ) | ( (~ ng23521)  &  wire34435 ) ;
 assign wire6732 = ( ng2463  &  ng2473  &  (~ ng853) ) ;
 assign wire6737 = ( ng2473  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire6738 = ( ng2463  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire6771 = ( wire3221  &  (~ wire33231)  &  (~ wire33232)  &  (~ wire33233) ) ;
 assign wire6791 = ( ng1491  &  wire32947 ) | ( ng1491  &  ng27875  &  wire32946 ) ;
 assign wire6818 = ( ng1173  &  ng1174  &  (~ ng1309) ) ;
 assign wire6819 = ( ng1173  &  ng1175  &  (~ ng1315) ) ;
 assign wire6820 = ( ng1174  &  ng1175  &  (~ ng1312) ) ;
 assign wire6821 = ( ng1173  &  ng1174  &  ng1175 ) ;
 assign wire6822 = ( ng1175  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire6823 = ( ng1174  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire6824 = ( ng1173  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6875 = ( ng1008  &  (~ ng2257)  &  ng17086 ) | ( ng1008  &  (~ ng17086)  &  ng23511 ) ;
 assign wire6881 = ( ng853  &  wire8487 ) | ( ng853  &  wire3150  &  wire32248 ) ;
 assign wire6883 = ( (~ ng15950)  &  (~ wire32243)  &  (~ wire32244)  &  wire32245 ) ;
 assign wire6921 = ( ng646  &  wire31591  &  wire31592  &  wire34269 ) ;
 assign wire6922 = ( (~ ng646)  &  wire34270 ) | ( (~ wire31591)  &  wire34270 ) | ( (~ wire31592)  &  wire34270 ) ;
 assign wire6923 = ( ng1315  &  wire6925 ) | ( ng1315  &  wire6926 ) | ( ng1315  &  wire6927 ) ;
 assign wire6925 = ( (~ wire6933)  &  (~ wire6934)  &  (~ wire34262)  &  wire34265 ) ;
 assign wire6926 = ( (~ wire6933)  &  (~ wire6934)  &  (~ wire34262)  &  wire34267 ) ;
 assign wire6927 = ( (~ ng13055)  &  (~ wire31469)  &  (~ wire31470) ) ;
 assign wire6928 = ( (~ wire34196)  &  (~ wire34197)  &  wire34198  &  wire34199 ) ;
 assign wire6929 = ( wire34196  &  wire34201  &  wire34202 ) | ( wire34197  &  wire34201  &  wire34202 ) ;
 assign wire6930 = ( wire34196  &  wire34204  &  wire34205 ) | ( wire34197  &  wire34204  &  wire34205 ) ;
 assign wire6931 = ( wire3949  &  (~ wire34196)  &  (~ wire34197)  &  wire34217 ) ;
 assign wire6932 = ( wire3344  &  (~ wire34186)  &  (~ wire34187)  &  wire34219 ) ;
 assign wire6933 = ( (~ ng10784)  &  (~ wire34243)  &  (~ wire34244)  &  wire34245 ) ;
 assign wire6934 = ( ng10789  &  (~ wire34243)  &  (~ wire34244)  &  wire34247 ) ;
 assign wire6939 = ( wire34215  &  wire34253 ) | ( wire34216  &  wire34253 ) ;
 assign wire6940 = ( wire3344  &  wire3949  &  wire34221 ) ;
 assign wire6941 = ( wire3345  &  wire3929  &  wire34223 ) ;
 assign wire6946 = ( wire3345  &  wire3949  &  (~ wire31502)  &  (~ wire31503) ) ;
 assign wire6947 = ( wire3344  &  wire3929  &  wire34186 ) | ( wire3344  &  wire3929  &  wire34187 ) ;
 assign wire6950 = ( (~ ng349)  &  (~ ng353)  &  (~ ng351) ) ;
 assign wire6951 = ( (~ ng1309)  &  (~ ng353)  &  (~ ng351) ) ;
 assign wire6952 = ( (~ ng1315)  &  (~ ng349)  &  (~ ng351) ) ;
 assign wire6955 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng353) ) ;
 assign wire6956 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng351) ) ;
 assign wire6958 = ( (~ ng324)  &  (~ ng394)  &  (~ ng396) ) ;
 assign wire6959 = ( (~ ng1315)  &  (~ ng394)  &  (~ ng396) ) ;
 assign wire6960 = ( (~ ng1309)  &  (~ ng324)  &  (~ ng396) ) ;
 assign wire6963 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng324) ) ;
 assign wire6964 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng396) ) ;
 assign wire6966 = ( (~ ng1312)  &  (~ ng383)  &  (~ ng379) ) ;
 assign wire6969 = ( (~ ng381)  &  (~ ng383)  &  (~ ng1309) ) ;
 assign wire6970 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng379) ) ;
 assign wire6971 = ( (~ ng1312)  &  (~ ng383)  &  (~ ng1309) ) ;
 assign wire6972 = ( (~ ng381)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire6974 = ( (~ ng366)  &  (~ ng368)  &  (~ ng364) ) ;
 assign wire6975 = ( (~ ng1312)  &  (~ ng368)  &  (~ ng364) ) ;
 assign wire6976 = ( (~ ng1315)  &  (~ ng366)  &  (~ ng364) ) ;
 assign wire6977 = ( (~ ng1309)  &  (~ ng366)  &  (~ ng368) ) ;
 assign wire6978 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng364) ) ;
 assign wire6979 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng368) ) ;
 assign wire6980 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng366) ) ;
 assign wire6982 = ( (~ ng599)  &  (~ ng596)  &  (~ ng185)  &  (~ ng602) ) ;
 assign wire6983 = ( (~ ng1312)  &  (~ ng596)  &  (~ ng185)  &  (~ ng602) ) ;
 assign wire6984 = ( (~ ng1309)  &  (~ ng599)  &  (~ ng185)  &  (~ ng602) ) ;
 assign wire6985 = ( wire34117  &  wire34120 ) | ( wire34118  &  wire34120 ) ;
 assign wire6988 = ( (~ ng542)  &  (~ ng599)  &  (~ ng596)  &  (~ ng602) ) ;
 assign wire6989 = ( (~ ng542)  &  (~ ng1312)  &  (~ ng596)  &  (~ ng602) ) ;
 assign wire6990 = ( (~ ng542)  &  (~ ng1309)  &  (~ ng599)  &  (~ ng602) ) ;
 assign wire6991 = ( (~ ng1315)  &  (~ ng599)  &  (~ ng596)  &  (~ ng185) ) ;
 assign wire6993 = ( (~ ng542)  &  (~ ng1315)  &  (~ ng599)  &  (~ ng596) ) ;
 assign wire6994 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng596)  &  (~ ng185) ) ;
 assign wire6996 = ( (~ ng542)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng596) ) ;
 assign wire6997 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng185)  &  (~ ng602) ) ;
 assign wire6999 = ( (~ ng542)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng602) ) ;
 assign wire7000 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng599)  &  (~ ng185) ) ;
 assign wire7002 = ( (~ ng542)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng599) ) ;
 assign wire7003 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7005 = ( (~ ng542)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire7006 = ( (~ ng1309)  &  (~ ng489)  &  (~ ng567) ) ;
 assign wire7011 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng489) ) ;
 assign wire7012 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng567) ) ;
 assign wire7014 = ( wire3142  &  (~ wire31587)  &  (~ wire31588)  &  (~ wire31589) ) ;
 assign wire7026 = ( ng23478  &  wire9118  &  wire34089 ) | ( ng23478  &  wire31438  &  wire34089 ) ;
 assign wire7029 = ( (~ wire31249)  &  (~ wire31250)  &  (~ wire31251)  &  wire34094 ) ;
 assign wire7030 = ( (~ wire31265)  &  (~ wire31266)  &  (~ wire31267)  &  wire34095 ) ;
 assign wire7045 = ( ng3135  &  (~ ng3120)  &  ng8430  &  wire34081 ) ;
 assign wire7046 = ( ng3135  &  (~ ng3120)  &  ng8430  &  wire34082 ) ;
 assign wire7048 = ( (~ ng185)  &  (~ ng8381)  &  (~ wire30893) ) ;
 assign wire7057 = ( wire3224  &  ng12082  &  (~ wire34076) ) | ( wire3224  &  (~ wire3336)  &  (~ wire34076) ) ;
 assign wire7058 = ( (~ ng557)  &  (~ ng510)  &  ng530  &  ng525 ) ;
 assign wire7069 = ( wire34044  &  wire34068 ) | ( wire34045  &  wire34068 ) | ( wire34049  &  wire34068 ) ;
 assign wire7070 = ( (~ ng499)  &  wire3140 ) | ( ng21851  &  wire3140 ) | ( wire3140  &  wire34028 ) ;
 assign wire7078 = ( ng739  &  (~ ng1309)  &  ng737 ) ;
 assign wire7083 = ( (~ ng1312)  &  (~ ng1309)  &  ng737 ) ;
 assign wire7084 = ( (~ ng1315)  &  ng739  &  (~ ng1309) ) ;
 assign wire7111 = ( ng12305  &  ng12269  &  wire34020 ) | ( (~ ng12305)  &  wire3124  &  wire34020 ) | ( ng12269  &  wire3124  &  wire34020 ) ;
 assign wire7114 = ( pg3229  &  (~ wire33988)  &  (~ wire33989) ) ;
 assign wire7119 = ( ng2654  &  ng2653  &  ng2652 ) ;
 assign wire7120 = ( (~ ng1312)  &  ng2653  &  ng2652 ) ;
 assign wire7121 = ( ng2654  &  (~ ng1309)  &  ng2652 ) ;
 assign wire7124 = ( (~ ng1312)  &  (~ ng1309)  &  ng2652 ) ;
 assign wire7125 = ( (~ ng1315)  &  ng2654  &  (~ ng1309) ) ;
 assign wire7127 = ( ng2656  &  ng2657  &  ng2655 ) ;
 assign wire7128 = ( (~ ng1309)  &  ng2657  &  ng2655 ) ;
 assign wire7129 = ( (~ ng1312)  &  ng2656  &  ng2655 ) ;
 assign wire7132 = ( (~ ng1312)  &  (~ ng1309)  &  ng2655 ) ;
 assign wire7133 = ( (~ ng1315)  &  (~ ng1309)  &  ng2657 ) ;
 assign wire7135 = ( ng2651  &  (~ ng1315)  &  ng2650 ) ;
 assign wire7138 = ( ng2649  &  ng2651  &  (~ ng1309) ) ;
 assign wire7139 = ( (~ ng1312)  &  (~ ng1315)  &  ng2650 ) ;
 assign wire7140 = ( ng2649  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire7141 = ( ng2651  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire7143 = ( ng2659  &  ng2660  &  ng2658 ) ;
 assign wire7144 = ( (~ ng1309)  &  ng2660  &  ng2658 ) ;
 assign wire7145 = ( (~ ng1312)  &  ng2659  &  ng2658 ) ;
 assign wire7148 = ( (~ ng1312)  &  (~ ng1309)  &  ng2658 ) ;
 assign wire7149 = ( (~ ng1315)  &  (~ ng1309)  &  ng2660 ) ;
 assign wire7152 = ( (~ wire31471)  &  wire33977 ) | ( (~ wire31472)  &  wire33977 ) | ( (~ wire31471)  &  wire33978 ) | ( (~ wire31472)  &  wire33978 ) ;
 assign wire7153 = ( (~ wire31471)  &  wire33967 ) | ( (~ wire31472)  &  wire33967 ) | ( (~ wire31471)  &  wire33968 ) | ( (~ wire31472)  &  wire33968 ) ;
 assign wire7154 = ( (~ ng1309)  &  (~ ng2685)  &  (~ ng2682) ) ;
 assign wire7159 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2685) ) ;
 assign wire7160 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2682) ) ;
 assign wire7162 = ( (~ ng2571)  &  (~ ng2568)  &  (~ ng2565) ) ;
 assign wire7163 = ( (~ ng1315)  &  (~ ng2568)  &  (~ ng2565) ) ;
 assign wire7164 = ( (~ ng1312)  &  (~ ng2571)  &  (~ ng2565) ) ;
 assign wire7165 = ( (~ ng1309)  &  (~ ng2571)  &  (~ ng2568) ) ;
 assign wire7166 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2565) ) ;
 assign wire7167 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2571) ) ;
 assign wire7168 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2568) ) ;
 assign wire7170 = ( (~ ng1315)  &  (~ ng2691)  &  (~ ng2688) ) ;
 assign wire7175 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2694) ) ;
 assign wire7176 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2691) ) ;
 assign wire7190 = ( (~ ng12180)  &  ng12121  &  ng18325  &  wire33940 ) | ( ng12180  &  (~ ng12121)  &  (~ ng18325)  &  wire33940 ) ;
 assign wire7191 = ( (~ ng12180)  &  ng12121  &  ng18325  &  wire33941 ) | ( ng12180  &  (~ ng12121)  &  (~ ng18325)  &  wire33941 ) ;
 assign wire7192 = ( (~ ng12180)  &  ng12121  &  ng18325  &  wire33942 ) | ( ng12180  &  (~ ng12121)  &  (~ ng18325)  &  wire33942 ) ;
 assign wire7196 = ( (~ ng2504)  &  (~ ng2507)  &  (~ ng853) ) ;
 assign wire7201 = ( (~ ng2504)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7202 = ( (~ ng826)  &  (~ ng2507)  &  (~ ng853) ) ;
 assign wire7204 = ( ng2255  &  ng2254  &  (~ ng853) ) ;
 assign wire7209 = ( ng2254  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7210 = ( ng2255  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7213 = ( (~ ng853)  &  (~ ng2513)  &  (~ ng2516) ) ;
 assign wire7218 = ( (~ ng823)  &  (~ ng853)  &  (~ ng2513) ) ;
 assign wire7219 = ( (~ ng826)  &  (~ ng853)  &  (~ ng2516) ) ;
 assign wire7225 = ( ng12005  &  (~ ng11917)  &  wire3925  &  (~ wire33878) ) ;
 assign wire7227 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33892 ) ;
 assign wire7228 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33894 ) ;
 assign wire7229 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33896 ) ;
 assign wire7230 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33898 ) ;
 assign wire7231 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33899 ) ;
 assign wire7232 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33900 ) ;
 assign wire7233 = ( ng2257  &  (~ ng25099)  &  (~ ng11962)  &  wire33901 ) ;
 assign wire7234 = ( ng2257  &  wire3046  &  (~ ng25099)  &  (~ ng11962) ) ;
 assign wire7235 = ( (~ ng2486)  &  (~ ng2483)  &  (~ ng853) ) ;
 assign wire7240 = ( (~ ng2483)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7241 = ( (~ ng2486)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7246 = ( (~ ng2495)  &  (~ ng826)  &  (~ ng2498) ) ;
 assign wire7249 = ( (~ ng2495)  &  (~ ng2492)  &  (~ ng853) ) ;
 assign wire7250 = ( (~ ng826)  &  (~ ng823)  &  (~ ng2498) ) ;
 assign wire7251 = ( (~ ng2492)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7252 = ( (~ ng2495)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7262 = ( ng2418  &  ng2429  &  (~ ng853) ) ;
 assign wire7267 = ( ng2429  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7268 = ( ng2418  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7270 = ( ng2448  &  ng2451  &  (~ ng826) ) ;
 assign wire7273 = ( ng2448  &  ng2459  &  (~ ng853) ) ;
 assign wire7274 = ( ng2451  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7275 = ( ng2459  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7276 = ( ng2448  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7278 = ( ng2444  &  ng2433  &  (~ ng853) ) ;
 assign wire7283 = ( ng2444  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7284 = ( ng2433  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7307 = ( (~ ng28584)  &  ng26941  &  wire33813 ) ;
 assign wire7308 = ( ng2190  &  wire33795 ) | ( ng2190  &  ng27892  &  wire33794 ) ;
 assign wire7327 = ( wire3925  &  (~ wire33538)  &  (~ wire33539) ) ;
 assign wire7331 = ( (~ ng2398)  &  ng823 ) ;
 assign wire7336 = ( (~ ng22400)  &  wire33548  &  wire33792 ) | ( (~ ng22400)  &  wire33549  &  wire33792 ) ;
 assign wire7337 = ( (~ ng18319)  &  (~ ng18053)  &  (~ ng18231) ) | ( (~ ng18606)  &  (~ ng18053)  &  (~ ng18231) ) ;
 assign wire7342 = ( (~ ng18319)  &  (~ ng18231)  &  wire3066 ) ;
 assign wire7343 = ( (~ ng18606)  &  (~ ng18053)  &  wire3066 ) ;
 assign wire7344 = ( (~ ng18319)  &  (~ ng18606)  &  wire3066 ) ;
 assign wire7359 = ( (~ ng18395)  &  (~ ng18578)  &  wire3055 ) | ( (~ ng18478)  &  (~ ng18578)  &  wire3055 ) ;
 assign wire7364 = ( (~ ng18395)  &  wire3055  &  wire3105 ) ;
 assign wire7365 = ( (~ ng18478)  &  (~ ng18578)  &  wire3105 ) ;
 assign wire7366 = ( (~ ng18395)  &  (~ ng18478)  &  wire3105 ) ;
 assign wire7383 = ( ng2221  &  ng2222  &  (~ ng853)  &  ng2180 ) ;
 assign wire7384 = ( ng2221  &  ng2220  &  (~ ng823)  &  ng2180 ) ;
 assign wire7385 = ( (~ ng823)  &  ng2224  &  ng2223  &  ng2185 ) ;
 assign wire7386 = ( (~ ng853)  &  ng2224  &  ng2225  &  ng2185 ) ;
 assign wire7387 = ( (~ ng826)  &  ng2220  &  (~ ng823)  &  ng2180 ) ;
 assign wire7388 = ( (~ ng826)  &  (~ ng823)  &  ng2223  &  ng2185 ) ;
 assign wire7389 = ( ng2221  &  (~ ng823)  &  (~ ng853)  &  ng2180 ) ;
 assign wire7390 = ( (~ ng823)  &  (~ ng853)  &  ng2224  &  ng2185 ) ;
 assign wire7391 = ( (~ ng826)  &  ng2222  &  (~ ng853)  &  ng2180 ) ;
 assign wire7392 = ( (~ ng826)  &  (~ ng853)  &  ng2225  &  ng2185 ) ;
 assign wire7393 = ( (~ ng2220)  &  ng853  &  (~ ng2180) ) ;
 assign wire7394 = ( (~ ng2222)  &  ng823  &  (~ ng2180) ) ;
 assign wire7395 = ( ng853  &  (~ ng2223)  &  (~ ng2185) ) ;
 assign wire7396 = ( ng823  &  (~ ng2225)  &  (~ ng2185) ) ;
 assign wire7397 = ( ng826  &  (~ ng2224)  &  (~ ng2185) ) ;
 assign wire7398 = ( (~ ng2221)  &  ng826  &  (~ ng2180) ) ;
 assign wire7399 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2180 ) ;
 assign wire7400 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2185 ) ;
 assign wire7409 = ( ng2245  &  ng2246  &  (~ ng853) ) ;
 assign wire7414 = ( ng2245  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7415 = ( ng2246  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7417 = ( (~ ng826)  &  ng2210  &  ng2208 ) ;
 assign wire7422 = ( ng2209  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7423 = ( (~ ng826)  &  (~ ng853)  &  ng2210 ) ;
 assign wire7425 = ( (~ ng853)  &  ng2218  &  ng2219 ) ;
 assign wire7430 = ( (~ ng823)  &  (~ ng853)  &  ng2218 ) ;
 assign wire7431 = ( (~ ng826)  &  (~ ng853)  &  ng2219 ) ;
 assign wire7435 = ( (~ ng853)  &  ng2227  &  ng2228  &  ng2190 ) ;
 assign wire7436 = ( (~ ng823)  &  ng2227  &  ng2226  &  ng2190 ) ;
 assign wire7437 = ( ng2233  &  (~ ng853)  &  ng2234  &  ng2200 ) ;
 assign wire7438 = ( ng2233  &  (~ ng823)  &  ng2232  &  ng2200 ) ;
 assign wire7439 = ( (~ ng826)  &  (~ ng823)  &  ng2226  &  ng2190 ) ;
 assign wire7440 = ( (~ ng826)  &  (~ ng823)  &  ng2232  &  ng2200 ) ;
 assign wire7441 = ( (~ ng823)  &  (~ ng853)  &  ng2227  &  ng2190 ) ;
 assign wire7442 = ( ng2233  &  (~ ng823)  &  (~ ng853)  &  ng2200 ) ;
 assign wire7443 = ( (~ ng826)  &  (~ ng853)  &  ng2228  &  ng2190 ) ;
 assign wire7444 = ( (~ ng826)  &  (~ ng853)  &  ng2234  &  ng2200 ) ;
 assign wire7445 = ( ng823  &  (~ ng2228)  &  (~ ng2190) ) ;
 assign wire7446 = ( ng853  &  (~ ng2226)  &  (~ ng2190) ) ;
 assign wire7447 = ( ng823  &  (~ ng2234)  &  (~ ng2200) ) ;
 assign wire7448 = ( ng853  &  (~ ng2232)  &  (~ ng2200) ) ;
 assign wire7449 = ( ng826  &  (~ ng2233)  &  (~ ng2200) ) ;
 assign wire7450 = ( ng826  &  (~ ng2227)  &  (~ ng2190) ) ;
 assign wire7451 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2190 ) ;
 assign wire7452 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2200 ) ;
 assign wire7455 = ( wire33630  &  (~ wire33640)  &  (~ wire33641) ) | ( wire33631  &  (~ wire33640)  &  (~ wire33641) ) ;
 assign wire7456 = ( (~ wire33630)  &  (~ wire33631)  &  wire33640 ) | ( (~ wire33630)  &  (~ wire33631)  &  wire33641 ) ;
 assign wire7459 = ( ng2239  &  ng2240  &  (~ ng853) ) ;
 assign wire7464 = ( ng2239  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7465 = ( ng2240  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7467 = ( ng2248  &  (~ ng853)  &  ng2249 ) ;
 assign wire7472 = ( ng2248  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7473 = ( (~ ng826)  &  (~ ng853)  &  ng2249 ) ;
 assign wire7475 = ( ng2231  &  ng2230  &  (~ ng853) ) ;
 assign wire7480 = ( ng2230  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7481 = ( ng2231  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7483 = ( ng2237  &  (~ ng853)  &  ng2236 ) ;
 assign wire7488 = ( (~ ng823)  &  (~ ng853)  &  ng2236 ) ;
 assign wire7489 = ( ng2237  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7491 = ( ng2207  &  ng2206  &  (~ ng853) ) ;
 assign wire7496 = ( ng2206  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7497 = ( ng2207  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7500 = ( (~ ng25969)  &  wire33574  &  wire33575  &  wire33579 ) ;
 assign wire7504 = ( ng2387  &  ng2388  &  (~ ng853) ) ;
 assign wire7509 = ( ng2387  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7510 = ( (~ ng826)  &  ng2388  &  (~ ng853) ) ;
 assign wire7512 = ( (~ ng853)  &  ng2391  &  ng2390 ) ;
 assign wire7517 = ( (~ ng823)  &  (~ ng853)  &  ng2390 ) ;
 assign wire7518 = ( (~ ng826)  &  (~ ng853)  &  ng2391 ) ;
 assign wire7520 = ( ng2394  &  (~ ng853)  &  ng2393 ) ;
 assign wire7521 = ( ng2394  &  ng2395  &  (~ ng826) ) ;
 assign wire7522 = ( ng2395  &  (~ ng823)  &  ng2393 ) ;
 assign wire7523 = ( ng2394  &  ng2395  &  ng2393 ) ;
 assign wire7524 = ( ng2395  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7525 = ( (~ ng823)  &  (~ ng853)  &  ng2393 ) ;
 assign wire7526 = ( ng2394  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7528 = ( (~ ng2264)  &  (~ ng826)  &  (~ ng2267) ) ;
 assign wire7531 = ( (~ ng2261)  &  (~ ng2264)  &  (~ ng853) ) ;
 assign wire7532 = ( (~ ng826)  &  (~ ng823)  &  (~ ng2267) ) ;
 assign wire7533 = ( (~ ng2261)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7534 = ( (~ ng2264)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7536 = ( (~ ng2282)  &  (~ ng853)  &  (~ ng2279) ) ;
 assign wire7541 = ( (~ ng823)  &  (~ ng853)  &  (~ ng2279) ) ;
 assign wire7542 = ( (~ ng2282)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7544 = ( (~ ng2306)  &  (~ ng2309)  &  (~ ng853) ) ;
 assign wire7549 = ( (~ ng2306)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7550 = ( (~ ng2309)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7552 = ( (~ ng2291)  &  (~ ng2288)  &  (~ ng853) ) ;
 assign wire7553 = ( (~ ng2294)  &  (~ ng2291)  &  (~ ng826) ) ;
 assign wire7554 = ( (~ ng2294)  &  (~ ng2288)  &  (~ ng823) ) ;
 assign wire7555 = ( (~ ng2294)  &  (~ ng2291)  &  (~ ng2288) ) ;
 assign wire7556 = ( (~ ng2294)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7557 = ( (~ ng2288)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7558 = ( (~ ng2291)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7560 = ( (~ ng2315)  &  (~ ng2318)  &  (~ ng853) ) ;
 assign wire7565 = ( (~ ng2315)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7566 = ( (~ ng2318)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7568 = ( (~ ng2333)  &  (~ ng853)  &  (~ ng2336) ) ;
 assign wire7573 = ( (~ ng2333)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7574 = ( (~ ng826)  &  (~ ng853)  &  (~ ng2336) ) ;
 assign wire7576 = ( (~ ng2327)  &  (~ ng2324)  &  (~ ng853) ) ;
 assign wire7577 = ( (~ ng2327)  &  (~ ng2330)  &  (~ ng826) ) ;
 assign wire7578 = ( (~ ng2324)  &  (~ ng2330)  &  (~ ng823) ) ;
 assign wire7579 = ( (~ ng2327)  &  (~ ng2324)  &  (~ ng2330) ) ;
 assign wire7580 = ( (~ ng2330)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7581 = ( (~ ng2324)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7582 = ( (~ ng2327)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7584 = ( (~ ng2297)  &  (~ ng2300)  &  (~ ng853) ) ;
 assign wire7585 = ( (~ ng2300)  &  (~ ng2303)  &  (~ ng826) ) ;
 assign wire7586 = ( (~ ng2297)  &  (~ ng2303)  &  (~ ng823) ) ;
 assign wire7587 = ( (~ ng2297)  &  (~ ng2300)  &  (~ ng2303) ) ;
 assign wire7588 = ( (~ ng2303)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7589 = ( (~ ng2297)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7590 = ( (~ ng2300)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7592 = ( (~ ng2270)  &  (~ ng2273)  &  (~ ng853) ) ;
 assign wire7597 = ( (~ ng2270)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7598 = ( (~ ng2273)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7600 = ( (~ ng2342)  &  (~ ng2345)  &  (~ ng853) ) ;
 assign wire7601 = ( (~ ng2345)  &  (~ ng2348)  &  (~ ng826) ) ;
 assign wire7602 = ( (~ ng2342)  &  (~ ng2348)  &  (~ ng823) ) ;
 assign wire7603 = ( (~ ng2342)  &  (~ ng2345)  &  (~ ng2348) ) ;
 assign wire7604 = ( (~ ng2348)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7605 = ( (~ ng2342)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7606 = ( (~ ng2345)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7612 = ( ng2251  &  ng2252  &  (~ ng853) ) ;
 assign wire7617 = ( ng2251  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7618 = ( ng2252  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7627 = ( (~ ng2033)  &  wire33417 ) | ( (~ ng2020)  &  wire33417 ) | ( (~ wire33414)  &  wire33417 ) ;
 assign wire7633 = ( ng1315  &  wire7635 ) | ( ng1315  &  wire7636 ) | ( ng1315  &  wire7637 ) ;
 assign wire7635 = ( (~ wire7640)  &  (~ wire33399)  &  (~ wire33401)  &  wire33403 ) ;
 assign wire7636 = ( (~ wire7640)  &  (~ wire33399)  &  (~ wire33401)  &  wire33405 ) ;
 assign wire7637 = ( (~ ng13055)  &  (~ wire33167)  &  (~ wire33168) ) ;
 assign wire7638 = ( wire33338  &  wire33340  &  wire33341 ) | ( wire33339  &  wire33340  &  wire33341 ) ;
 assign wire7639 = ( wire3440  &  wire33328  &  wire33343 ) | ( wire3440  &  wire33329  &  wire33343 ) ;
 assign wire7640 = ( wire3437  &  (~ wire33376)  &  (~ wire33377)  &  wire33378 ) ;
 assign wire7641 = ( (~ wire3233)  &  (~ wire33353)  &  (~ wire33354)  &  wire33380 ) ;
 assign wire7644 = ( wire3354  &  wire3437  &  (~ wire33117)  &  (~ wire33118) ) ;
 assign wire7649 = ( wire33353  &  wire33391 ) | ( wire33354  &  wire33391 ) ;
 assign wire7650 = ( wire3354  &  wire3440  &  wire33355 ) ;
 assign wire7651 = ( wire3364  &  wire3437  &  wire33357 ) ;
 assign wire7652 = ( wire3364  &  (~ wire33353)  &  (~ wire33354)  &  wire33359 ) ;
 assign wire7653 = ( wire3354  &  wire33127  &  wire33361 ) | ( wire3354  &  wire33128  &  wire33361 ) ;
 assign wire7660 = ( ng1966  &  ng1965  &  ng1964 ) ;
 assign wire7661 = ( (~ ng1312)  &  ng1965  &  ng1964 ) ;
 assign wire7662 = ( (~ ng1309)  &  ng1966  &  ng1964 ) ;
 assign wire7665 = ( (~ ng1312)  &  (~ ng1309)  &  ng1964 ) ;
 assign wire7666 = ( (~ ng1315)  &  (~ ng1309)  &  ng1966 ) ;
 assign wire7668 = ( (~ ng1705)  &  (~ ng1777)  &  (~ ng1775) ) ;
 assign wire7669 = ( (~ ng1315)  &  (~ ng1777)  &  (~ ng1775) ) ;
 assign wire7670 = ( (~ ng1312)  &  (~ ng1705)  &  (~ ng1775) ) ;
 assign wire7671 = ( (~ ng1309)  &  (~ ng1705)  &  (~ ng1777) ) ;
 assign wire7672 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1775) ) ;
 assign wire7673 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1705) ) ;
 assign wire7674 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1777) ) ;
 assign wire7676 = ( (~ ng1730)  &  (~ ng1732)  &  (~ ng1734) ) ;
 assign wire7677 = ( (~ ng1309)  &  (~ ng1732)  &  (~ ng1734) ) ;
 assign wire7678 = ( (~ ng1312)  &  (~ ng1730)  &  (~ ng1734) ) ;
 assign wire7681 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1734) ) ;
 assign wire7682 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1732) ) ;
 assign wire7684 = ( (~ ng1749)  &  (~ ng1747)  &  (~ ng1745) ) ;
 assign wire7685 = ( (~ ng1312)  &  (~ ng1749)  &  (~ ng1745) ) ;
 assign wire7686 = ( (~ ng1315)  &  (~ ng1747)  &  (~ ng1745) ) ;
 assign wire7687 = ( (~ ng1309)  &  (~ ng1749)  &  (~ ng1747) ) ;
 assign wire7688 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1745) ) ;
 assign wire7689 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1749) ) ;
 assign wire7690 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1747) ) ;
 assign wire7692 = ( (~ ng1760)  &  (~ ng1764)  &  (~ ng1762) ) ;
 assign wire7693 = ( (~ ng1309)  &  (~ ng1764)  &  (~ ng1762) ) ;
 assign wire7694 = ( (~ ng1315)  &  (~ ng1760)  &  (~ ng1762) ) ;
 assign wire7697 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1764) ) ;
 assign wire7698 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1762) ) ;
 assign wire7700 = ( (~ ng1979)  &  (~ ng1309)  &  (~ ng185)  &  (~ ng1982) ) ;
 assign wire7701 = ( (~ ng1979)  &  (~ ng1976)  &  (~ ng185)  &  (~ ng1982) ) ;
 assign wire7702 = ( (~ ng1312)  &  (~ ng1976)  &  (~ ng185)  &  (~ ng1982) ) ;
 assign wire7703 = ( (~ ng1315)  &  (~ ng1979)  &  (~ ng1976)  &  (~ ng185) ) ;
 assign wire7704 = ( wire33251  &  wire33254 ) | ( wire33252  &  wire33254 ) ;
 assign wire7708 = ( (~ ng1922)  &  (~ ng1979)  &  (~ ng1309)  &  (~ ng1982) ) ;
 assign wire7709 = ( (~ ng1922)  &  (~ ng1979)  &  (~ ng1976)  &  (~ ng1982) ) ;
 assign wire7710 = ( (~ ng1922)  &  (~ ng1312)  &  (~ ng1976)  &  (~ ng1982) ) ;
 assign wire7711 = ( (~ ng1922)  &  (~ ng1315)  &  (~ ng1979)  &  (~ ng1976) ) ;
 assign wire7712 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1976)  &  (~ ng185) ) ;
 assign wire7714 = ( (~ ng1922)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1976) ) ;
 assign wire7715 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng185)  &  (~ ng1982) ) ;
 assign wire7717 = ( (~ ng1922)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng1982) ) ;
 assign wire7718 = ( (~ ng1315)  &  (~ ng1979)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7720 = ( (~ ng1922)  &  (~ ng1315)  &  (~ ng1979)  &  (~ ng1309) ) ;
 assign wire7721 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7723 = ( (~ ng1922)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire7724 = ( (~ ng1947)  &  (~ ng1309)  &  (~ ng1870) ) ;
 assign wire7729 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1870) ) ;
 assign wire7730 = ( (~ ng1315)  &  (~ ng1947)  &  (~ ng1309) ) ;
 assign wire7732 = ( wire3142  &  (~ wire33231)  &  (~ wire33232)  &  (~ wire33233) ) ;
 assign wire7734 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1967)  &  (~ ng185) ) ;
 assign wire7735 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1967)  &  (~ ng185) ) ;
 assign wire7736 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1967)  &  (~ ng185) ) ;
 assign wire7737 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7738 = ( wire33186  &  wire33189 ) | ( wire33187  &  wire33189 ) ;
 assign wire7741 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1904)  &  (~ ng1967) ) ;
 assign wire7742 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1904)  &  (~ ng1967) ) ;
 assign wire7743 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1904)  &  (~ ng1967) ) ;
 assign wire7745 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1309)  &  (~ ng1904) ) ;
 assign wire7746 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1967)  &  (~ ng185) ) ;
 assign wire7748 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1904)  &  (~ ng1967) ) ;
 assign wire7749 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7751 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng1904) ) ;
 assign wire7752 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7754 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng1904) ) ;
 assign wire7755 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire7756 = ( wire3049  &  wire33186 ) | ( wire3049  &  wire33187 ) ;
 assign wire7757 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng1904) ) ;
 assign wire7758 = ( (~ ng1949)  &  (~ ng1951)  &  (~ ng1953) ) ;
 assign wire7759 = ( (~ ng1309)  &  (~ ng1951)  &  (~ ng1953) ) ;
 assign wire7760 = ( (~ ng1312)  &  (~ ng1949)  &  (~ ng1953) ) ;
 assign wire7763 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1953) ) ;
 assign wire7764 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1951) ) ;
 assign wire7769 = ( (~ wire31471)  &  wire33157 ) | ( (~ wire31472)  &  wire33157 ) | ( (~ wire31471)  &  wire33158 ) | ( (~ wire31472)  &  wire33158 ) ;
 assign wire7770 = ( (~ wire31471)  &  wire33167 ) | ( (~ wire31472)  &  wire33167 ) | ( (~ wire31471)  &  wire33168 ) | ( (~ wire31472)  &  wire33168 ) ;
 assign wire7771 = ( (~ ng1874)  &  (~ ng1309)  &  (~ ng1877) ) ;
 assign wire7776 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1877) ) ;
 assign wire7777 = ( (~ ng1315)  &  (~ ng1874)  &  (~ ng1309) ) ;
 assign wire7779 = ( (~ ng1312)  &  (~ ng1994)  &  (~ ng2000) ) ;
 assign wire7784 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2000) ) ;
 assign wire7785 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1997) ) ;
 assign wire7787 = ( (~ ng1315)  &  (~ ng1985)  &  (~ ng1988) ) ;
 assign wire7792 = ( (~ ng1991)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire7793 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1988) ) ;
 assign wire7797 = ( ng1960  &  ng1958  &  (~ ng1309) ) ;
 assign wire7802 = ( (~ ng1312)  &  ng1958  &  (~ ng1309) ) ;
 assign wire7803 = ( ng1960  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire7807 = ( ng1956  &  ng1957  &  ng1955 ) ;
 assign wire7808 = ( (~ ng1309)  &  ng1957  &  ng1955 ) ;
 assign wire7809 = ( (~ ng1312)  &  ng1956  &  ng1955 ) ;
 assign wire7812 = ( (~ ng1312)  &  (~ ng1309)  &  ng1955 ) ;
 assign wire7813 = ( (~ ng1315)  &  (~ ng1309)  &  ng1957 ) ;
 assign wire7815 = ( ng1962  &  ng1963  &  ng1961 ) ;
 assign wire7816 = ( (~ ng1309)  &  ng1963  &  ng1961 ) ;
 assign wire7817 = ( (~ ng1312)  &  ng1962  &  ng1961 ) ;
 assign wire7820 = ( (~ ng1312)  &  (~ ng1309)  &  ng1961 ) ;
 assign wire7821 = ( (~ ng1315)  &  (~ ng1309)  &  ng1963 ) ;
 assign wire7829 = ( ng11630  &  (~ wire33106)  &  wire33107 ) | ( (~ ng27730)  &  (~ wire33106)  &  wire33107 ) ;
 assign wire7830 = ( wire33106  &  wire33108 ) | ( (~ ng11630)  &  ng27730  &  wire33108 ) ;
 assign wire7837 = ( (~ ng2257)  &  wire33103 ) | ( (~ ng23526)  &  wire33103 ) ;
 assign wire7844 = ( (~ ng12108)  &  ng18218  &  ng12057  &  wire33087 ) | ( ng12108  &  (~ ng18218)  &  (~ ng12057)  &  wire33087 ) ;
 assign wire7845 = ( (~ ng12108)  &  ng18218  &  ng12057  &  wire33088 ) | ( ng12108  &  (~ ng18218)  &  (~ ng12057)  &  wire33088 ) ;
 assign wire7846 = ( (~ ng12108)  &  ng18218  &  ng12057  &  wire33089 ) | ( ng12108  &  (~ ng18218)  &  (~ ng12057)  &  wire33089 ) ;
 assign wire7850 = ( (~ ng853)  &  (~ ng1813)  &  (~ ng1810) ) ;
 assign wire7855 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1810) ) ;
 assign wire7856 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1813) ) ;
 assign wire7858 = ( ng1560  &  ng1561  &  (~ ng853) ) ;
 assign wire7863 = ( ng1560  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7864 = ( ng1561  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7867 = ( (~ ng1822)  &  (~ ng1819)  &  (~ ng853) ) ;
 assign wire7868 = ( (~ ng1825)  &  (~ ng1822)  &  (~ ng826) ) ;
 assign wire7869 = ( (~ ng1825)  &  (~ ng1819)  &  (~ ng823) ) ;
 assign wire7870 = ( (~ ng1825)  &  (~ ng1822)  &  (~ ng1819) ) ;
 assign wire7871 = ( (~ ng1825)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7872 = ( (~ ng1819)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7873 = ( (~ ng1822)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7879 = ( ng11952  &  (~ ng11875)  &  wire3935  &  (~ wire33025) ) ;
 assign wire7881 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33039 ) ;
 assign wire7882 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33041 ) ;
 assign wire7883 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33043 ) ;
 assign wire7884 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33045 ) ;
 assign wire7885 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33046 ) ;
 assign wire7886 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33047 ) ;
 assign wire7887 = ( ng2257  &  (~ ng11912)  &  (~ ng25091)  &  wire33048 ) ;
 assign wire7888 = ( ng2257  &  wire3046  &  (~ ng11912)  &  (~ ng25091) ) ;
 assign wire7892 = ( (~ ng1792)  &  (~ ng853)  &  (~ ng1789) ) ;
 assign wire7897 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1789) ) ;
 assign wire7898 = ( (~ ng1792)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7900 = ( (~ ng1798)  &  (~ ng1801)  &  (~ ng853) ) ;
 assign wire7901 = ( (~ ng1801)  &  (~ ng1804)  &  (~ ng826) ) ;
 assign wire7902 = ( (~ ng1798)  &  (~ ng1804)  &  (~ ng823) ) ;
 assign wire7903 = ( (~ ng1798)  &  (~ ng1801)  &  (~ ng1804) ) ;
 assign wire7904 = ( (~ ng1804)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7905 = ( (~ ng1798)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7906 = ( (~ ng1801)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7914 = ( (~ ng826)  &  ng1724  &  ng1727 ) ;
 assign wire7919 = ( ng1735  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7920 = ( (~ ng826)  &  ng1724  &  (~ ng853) ) ;
 assign wire7922 = ( ng1765  &  ng1754  &  (~ ng853) ) ;
 assign wire7927 = ( ng1765  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7928 = ( ng1754  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7930 = ( ng1739  &  ng1750  &  (~ ng853) ) ;
 assign wire7931 = ( ng1739  &  ng1742  &  (~ ng826) ) ;
 assign wire7932 = ( ng1750  &  ng1742  &  (~ ng823) ) ;
 assign wire7933 = ( ng1739  &  ng1750  &  ng1742 ) ;
 assign wire7934 = ( ng1742  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire7935 = ( ng1750  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire7936 = ( ng1739  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire7941 = ( ng1453  &  (~ ng17031)  &  (~ ng23528) ) ;
 assign wire7954 = ( (~ ng28556)  &  (~ ng26918)  &  wire32681 ) | ( (~ ng28556)  &  (~ ng26918)  &  wire32682 ) ;
 assign wire7955 = ( ng1506  &  wire32947 ) | ( ng1506  &  ng27875  &  wire32946 ) ;
 assign wire7972 = ( wire3935  &  (~ wire32640)  &  (~ wire32641) ) ;
 assign wire7976 = ( (~ ng1704)  &  ng823 ) ;
 assign wire7977 = ( (~ wire32902)  &  (~ wire32903)  &  (~ wire32904)  &  wire32906 ) ;
 assign wire7978 = ( (~ wire32902)  &  (~ wire32903)  &  (~ wire32904)  &  wire32907 ) ;
 assign wire7979 = ( (~ wire32902)  &  (~ wire32903)  &  (~ wire32904)  &  wire32908 ) ;
 assign wire7981 = ( ng17124  &  (~ wire32902)  &  (~ wire32903)  &  (~ wire32904) ) ;
 assign wire7982 = ( (~ ng17942)  &  (~ ng18212)  &  (~ ng18115) ) | ( (~ ng18556)  &  (~ ng18212)  &  (~ ng18115) ) ;
 assign wire7987 = ( (~ ng17942)  &  (~ ng18115)  &  wire3108 ) ;
 assign wire7988 = ( (~ ng18556)  &  (~ ng18212)  &  wire3108 ) ;
 assign wire7989 = ( (~ ng17942)  &  (~ ng18556)  &  wire3108 ) ;
 assign wire8004 = ( (~ ng18561)  &  (~ ng18514)  &  (~ ng18383) ) | ( (~ ng18458)  &  (~ ng18514)  &  (~ ng18383) ) ;
 assign wire8009 = ( (~ ng18561)  &  (~ ng18383)  &  wire3068 ) ;
 assign wire8010 = ( (~ ng18458)  &  (~ ng18514)  &  wire3068 ) ;
 assign wire8011 = ( (~ ng18561)  &  (~ ng18458)  &  wire3068 ) ;
 assign wire8026 = ( (~ wire32816)  &  (~ wire32817)  &  wire32819 ) ;
 assign wire8027 = ( (~ wire32828)  &  (~ wire32829)  &  wire32831 ) ;
 assign wire8028 = ( (~ wire32816)  &  (~ wire32817)  &  wire32833 ) ;
 assign wire8029 = ( (~ wire32828)  &  (~ wire32829)  &  wire32835 ) ;
 assign wire8030 = ( (~ wire32816)  &  (~ wire32817)  &  wire32837 ) ;
 assign wire8035 = ( (~ wire32828)  &  (~ wire32829)  &  wire32843 ) ;
 assign wire8036 = ( (~ wire32816)  &  (~ wire32817)  &  wire32844 ) ;
 assign wire8041 = ( (~ ng1545)  &  ng826  &  wire32828 ) | ( (~ ng1545)  &  ng826  &  wire32829 ) ;
 assign wire8042 = ( (~ ng1543)  &  ng823  &  wire32816 ) | ( (~ ng1543)  &  ng823  &  wire32817 ) ;
 assign wire8043 = ( (~ ng1546)  &  ng823  &  wire32828 ) | ( (~ ng1546)  &  ng823  &  wire32829 ) ;
 assign wire8044 = ( wire3046  &  (~ wire32816)  &  (~ wire32817) ) ;
 assign wire8046 = ( (~ ng1506)  &  (~ wire32858)  &  (~ wire32859) ) ;
 assign wire8047 = ( ng1506  &  wire32858 ) | ( ng1506  &  wire32859 ) ;
 assign wire8050 = ( (~ ng1501)  &  (~ wire32878)  &  (~ wire32879) ) ;
 assign wire8051 = ( ng1501  &  wire32878 ) | ( ng1501  &  wire32879 ) ;
 assign wire8054 = ( ng1552  &  ng1551  &  (~ ng853) ) ;
 assign wire8055 = ( ng1552  &  ng1550  &  (~ ng826) ) ;
 assign wire8056 = ( ng1551  &  ng1550  &  (~ ng823) ) ;
 assign wire8057 = ( ng1552  &  ng1551  &  ng1550 ) ;
 assign wire8058 = ( ng1550  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8059 = ( ng1551  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8060 = ( ng1552  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8062 = ( ng1539  &  ng1540  &  (~ ng853) ) ;
 assign wire8067 = ( ng1539  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8068 = ( ng1540  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8070 = ( ng1534  &  ng1533  &  (~ ng853) ) ;
 assign wire8075 = ( ng1533  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8076 = ( ng1534  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8086 = ( ng823  &  (~ ng1516)  &  (~ ng1476) ) ;
 assign wire8087 = ( ng853  &  (~ ng1514)  &  (~ ng1476) ) ;
 assign wire8088 = ( (~ ng1529)  &  ng853  &  (~ ng1491) ) ;
 assign wire8089 = ( (~ ng1530)  &  ng826  &  (~ ng1491) ) ;
 assign wire8090 = ( (~ ng1531)  &  ng823  &  (~ ng1491) ) ;
 assign wire8094 = ( (~ ng1486)  &  (~ wire32778)  &  (~ wire32779) ) ;
 assign wire8095 = ( ng1486  &  wire32778 ) | ( ng1486  &  wire32779 ) ;
 assign wire8098 = ( ng1512  &  ng1513  &  (~ ng853) ) ;
 assign wire8103 = ( ng1512  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8104 = ( ng1513  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8106 = ( ng1527  &  ng1528  &  (~ ng853) ) ;
 assign wire8111 = ( ng1527  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8112 = ( ng1528  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8114 = ( ng1525  &  ng1524  &  (~ ng853) ) ;
 assign wire8119 = ( ng1524  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8120 = ( ng1525  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8122 = ( ng1536  &  ng1537  &  (~ ng853) ) ;
 assign wire8127 = ( ng1536  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8128 = ( ng1537  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8130 = ( ng1557  &  ng1558  &  ng1556 ) ;
 assign wire8131 = ( (~ ng826)  &  ng1558  &  ng1556 ) ;
 assign wire8132 = ( (~ ng823)  &  ng1557  &  ng1556 ) ;
 assign wire8133 = ( (~ ng853)  &  ng1557  &  ng1558 ) ;
 assign wire8134 = ( (~ ng826)  &  (~ ng823)  &  ng1556 ) ;
 assign wire8135 = ( (~ ng823)  &  (~ ng853)  &  ng1557 ) ;
 assign wire8136 = ( (~ ng826)  &  (~ ng853)  &  ng1558 ) ;
 assign wire8138 = ( ng1555  &  (~ ng826)  &  ng1553 ) ;
 assign wire8141 = ( ng1554  &  ng1555  &  (~ ng853) ) ;
 assign wire8142 = ( (~ ng826)  &  (~ ng823)  &  ng1553 ) ;
 assign wire8143 = ( ng1554  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8144 = ( ng1555  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8146 = ( ng25964  &  wire32721  &  wire32722 ) ;
 assign wire8147 = ( (~ ng25964)  &  wire32726  &  wire32727  &  wire32731 ) ;
 assign wire8151 = ( ng1696  &  ng1697  &  (~ ng853) ) ;
 assign wire8156 = ( ng1696  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8157 = ( ng1697  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8159 = ( ng1693  &  (~ ng853)  &  ng1694 ) ;
 assign wire8164 = ( ng1693  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8165 = ( (~ ng826)  &  (~ ng853)  &  ng1694 ) ;
 assign wire8167 = ( ng1700  &  ng1699  &  (~ ng853) ) ;
 assign wire8168 = ( ng1700  &  ng1701  &  (~ ng826) ) ;
 assign wire8169 = ( ng1701  &  ng1699  &  (~ ng823) ) ;
 assign wire8170 = ( ng1700  &  ng1701  &  ng1699 ) ;
 assign wire8171 = ( ng1701  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8172 = ( ng1699  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8173 = ( ng1700  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8175 = ( (~ ng853)  &  (~ ng1606)  &  (~ ng1603) ) ;
 assign wire8180 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1603) ) ;
 assign wire8181 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1606) ) ;
 assign wire8183 = ( (~ ng853)  &  (~ ng1615)  &  (~ ng1612) ) ;
 assign wire8188 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1612) ) ;
 assign wire8189 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1615) ) ;
 assign wire8191 = ( (~ ng1597)  &  (~ ng1594)  &  (~ ng853) ) ;
 assign wire8196 = ( (~ ng1594)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8197 = ( (~ ng1597)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8199 = ( (~ ng826)  &  (~ ng1624)  &  (~ ng1627) ) ;
 assign wire8202 = ( (~ ng1624)  &  (~ ng1621)  &  (~ ng853) ) ;
 assign wire8203 = ( (~ ng826)  &  (~ ng823)  &  (~ ng1627) ) ;
 assign wire8204 = ( (~ ng1621)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8205 = ( (~ ng826)  &  (~ ng1624)  &  (~ ng853) ) ;
 assign wire8207 = ( (~ ng1579)  &  (~ ng853)  &  (~ ng1576) ) ;
 assign wire8212 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1576) ) ;
 assign wire8213 = ( (~ ng1579)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8215 = ( (~ ng853)  &  (~ ng1630)  &  (~ ng1633) ) ;
 assign wire8220 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1630) ) ;
 assign wire8221 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1633) ) ;
 assign wire8223 = ( (~ ng823)  &  (~ ng1645)  &  (~ ng1639) ) ;
 assign wire8228 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1639) ) ;
 assign wire8229 = ( (~ ng1642)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8231 = ( (~ ng1651)  &  (~ ng1648)  &  (~ ng853) ) ;
 assign wire8236 = ( (~ ng1648)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8237 = ( (~ ng826)  &  (~ ng1651)  &  (~ ng853) ) ;
 assign wire8239 = ( (~ ng1567)  &  (~ ng853)  &  (~ ng1570) ) ;
 assign wire8244 = ( (~ ng1567)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8245 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1570) ) ;
 assign wire8247 = ( (~ ng1585)  &  (~ ng853)  &  (~ ng1588) ) ;
 assign wire8252 = ( (~ ng1585)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8253 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1588) ) ;
 assign wire8274 = ( ng1332  &  wire32566  &  wire32567  &  wire32568 ) ;
 assign wire8275 = ( (~ ng1332)  &  wire32569 ) | ( (~ wire32566)  &  wire32569 ) | ( (~ wire32567)  &  wire32569 ) ;
 assign wire8280 = ( (~ ng13055)  &  (~ wire32272)  &  (~ wire32273) ) ;
 assign wire8281 = ( (~ ng1273)  &  (~ ng1276)  &  (~ ng1279)  &  (~ ng185) ) ;
 assign wire8282 = ( (~ ng1312)  &  (~ ng1273)  &  (~ ng1279)  &  (~ ng185) ) ;
 assign wire8283 = ( (~ ng1309)  &  (~ ng1276)  &  (~ ng1279)  &  (~ ng185) ) ;
 assign wire8284 = ( (~ ng1315)  &  (~ ng1273)  &  (~ ng1276)  &  (~ ng185) ) ;
 assign wire8285 = ( wire32489  &  wire32492 ) | ( wire32490  &  wire32492 ) ;
 assign wire8287 = ( (~ ng1210)  &  (~ ng1273)  &  (~ ng1276)  &  (~ ng1279) ) ;
 assign wire8288 = ( (~ ng1210)  &  (~ ng1312)  &  (~ ng1273)  &  (~ ng1279) ) ;
 assign wire8290 = ( (~ ng1210)  &  (~ ng1309)  &  (~ ng1276)  &  (~ ng1279) ) ;
 assign wire8292 = ( (~ ng1210)  &  (~ ng1315)  &  (~ ng1273)  &  (~ ng1276) ) ;
 assign wire8293 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1273)  &  (~ ng185) ) ;
 assign wire8295 = ( (~ ng1210)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1273) ) ;
 assign wire8296 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1279)  &  (~ ng185) ) ;
 assign wire8298 = ( (~ ng1210)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng1279) ) ;
 assign wire8299 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1276)  &  (~ ng185) ) ;
 assign wire8301 = ( (~ ng1210)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng1276) ) ;
 assign wire8302 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire8304 = ( (~ ng1210)  &  (~ ng1312)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8305 = ( (~ ng1309)  &  (~ ng1259)  &  (~ ng1257) ) ;
 assign wire8310 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1259) ) ;
 assign wire8311 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1257) ) ;
 assign wire8314 = ( (~ ng12207)  &  wire32445  &  wire32446 ) | ( wire8332  &  wire32445  &  wire32446 ) ;
 assign wire8315 = ( (~ wire8334)  &  (~ wire8335)  &  wire32448  &  wire32449 ) ;
 assign wire8316 = ( wire32313  &  wire32451  &  wire32452 ) | ( wire32314  &  wire32451  &  wire32452 ) ;
 assign wire8317 = ( ng10793  &  (~ ng12152)  &  ng10801  &  ng12207 ) ;
 assign wire8318 = ( ng10814  &  (~ wire8334)  &  (~ wire8335)  &  wire32456 ) ;
 assign wire8323 = ( (~ wire8334)  &  (~ wire8335)  &  wire32540  &  wire32541 ) ;
 assign wire8324 = ( wire3288  &  (~ wire32313)  &  (~ wire32314)  &  wire32543 ) ;
 assign wire8326 = ( ng10801  &  (~ ng12207)  &  wire32547 ) | ( ng10801  &  wire8332  &  wire32547 ) ;
 assign wire8327 = ( (~ ng10801)  &  wire8334  &  wire32549 ) | ( (~ ng10801)  &  wire8335  &  wire32549 ) ;
 assign wire8329 = ( wire8332  &  wire32553 ) | ( (~ wire32429)  &  (~ wire32430)  &  wire32553 ) ;
 assign wire8330 = ( wire8334  &  wire32554 ) | ( wire8335  &  wire32554 ) ;
 assign wire8332 = ( wire32303  &  (~ wire32399)  &  (~ wire32400) ) | ( wire32304  &  (~ wire32399)  &  (~ wire32400) ) ;
 assign wire8334 = ( wire32313  &  wire32399 ) | ( wire32314  &  wire32399 ) | ( wire32313  &  wire32400 ) | ( wire32314  &  wire32400 ) ;
 assign wire8335 = ( (~ wire32399)  &  (~ wire32400)  &  (~ wire32429)  &  (~ wire32430) ) ;
 assign wire8336 = ( ng1267  &  ng1269  &  (~ ng1309) ) ;
 assign wire8337 = ( ng1269  &  ng1268  &  (~ ng1315) ) ;
 assign wire8338 = ( ng1267  &  ng1268  &  (~ ng1312) ) ;
 assign wire8339 = ( ng1267  &  ng1269  &  ng1268 ) ;
 assign wire8340 = ( ng1268  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire8341 = ( ng1267  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire8342 = ( ng1269  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8344 = ( (~ ng1053)  &  (~ ng1315)  &  (~ ng1051) ) ;
 assign wire8347 = ( (~ ng1053)  &  (~ ng1055)  &  (~ ng1309) ) ;
 assign wire8348 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1051) ) ;
 assign wire8349 = ( (~ ng1055)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire8350 = ( (~ ng1053)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8352 = ( (~ ng1083)  &  (~ ng1309)  &  (~ ng1011) ) ;
 assign wire8357 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1011) ) ;
 assign wire8358 = ( (~ ng1083)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8360 = ( (~ ng1070)  &  (~ ng1066)  &  (~ ng1068) ) ;
 assign wire8361 = ( (~ ng1315)  &  (~ ng1066)  &  (~ ng1068) ) ;
 assign wire8362 = ( (~ ng1309)  &  (~ ng1070)  &  (~ ng1068) ) ;
 assign wire8365 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1070) ) ;
 assign wire8366 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1068) ) ;
 assign wire8368 = ( (~ ng1309)  &  (~ ng1038)  &  (~ ng1040) ) ;
 assign wire8373 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1040) ) ;
 assign wire8374 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1038) ) ;
 assign wire8376 = ( wire32334  &  wire32337 ) | ( wire32335  &  wire32337 ) ;
 assign wire8380 = ( (~ ng1315)  &  (~ ng1282)  &  (~ ng1285)  &  (~ ng1228) ) ;
 assign wire8381 = ( (~ ng1282)  &  (~ ng1285)  &  (~ ng1288)  &  (~ ng1228) ) ;
 assign wire8382 = ( (~ ng1309)  &  (~ ng1285)  &  (~ ng1288)  &  (~ ng1228) ) ;
 assign wire8383 = ( (~ ng1312)  &  (~ ng1282)  &  (~ ng1288)  &  (~ ng1228) ) ;
 assign wire8384 = ( (~ ng1315)  &  (~ ng1282)  &  (~ ng1285)  &  (~ ng185) ) ;
 assign wire8385 = ( (~ ng1282)  &  (~ ng1285)  &  (~ ng1288)  &  (~ ng185) ) ;
 assign wire8386 = ( (~ ng1309)  &  (~ ng1285)  &  (~ ng1288)  &  (~ ng185) ) ;
 assign wire8387 = ( (~ ng1312)  &  (~ ng1282)  &  (~ ng1288)  &  (~ ng185) ) ;
 assign wire8389 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1282)  &  (~ ng1228) ) ;
 assign wire8390 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1282)  &  (~ ng185) ) ;
 assign wire8392 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1288)  &  (~ ng1228) ) ;
 assign wire8393 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1288)  &  (~ ng185) ) ;
 assign wire8395 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1285)  &  (~ ng1228) ) ;
 assign wire8396 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1285)  &  (~ ng185) ) ;
 assign wire8397 = ( wire3049  &  wire32334 ) | ( wire3049  &  wire32335 ) ;
 assign wire8398 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng1228) ) ;
 assign wire8399 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire8400 = ( (~ ng1251)  &  (~ ng1253)  &  (~ ng1176) ) ;
 assign wire8401 = ( (~ ng1309)  &  (~ ng1253)  &  (~ ng1176) ) ;
 assign wire8402 = ( (~ ng1312)  &  (~ ng1251)  &  (~ ng1176) ) ;
 assign wire8405 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1176) ) ;
 assign wire8406 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1253) ) ;
 assign wire8414 = ( ng1263  &  ng1262  &  ng1261 ) ;
 assign wire8415 = ( (~ ng1312)  &  ng1262  &  ng1261 ) ;
 assign wire8416 = ( (~ ng1309)  &  ng1263  &  ng1261 ) ;
 assign wire8419 = ( (~ ng1312)  &  (~ ng1309)  &  ng1261 ) ;
 assign wire8420 = ( (~ ng1315)  &  (~ ng1309)  &  ng1263 ) ;
 assign wire8422 = ( ng1264  &  ng1266  &  ng1265 ) ;
 assign wire8423 = ( (~ ng1315)  &  ng1266  &  ng1265 ) ;
 assign wire8424 = ( (~ ng1312)  &  ng1264  &  ng1265 ) ;
 assign wire8425 = ( ng1264  &  (~ ng1309)  &  ng1266 ) ;
 assign wire8426 = ( (~ ng1312)  &  (~ ng1315)  &  ng1265 ) ;
 assign wire8427 = ( (~ ng1312)  &  ng1264  &  (~ ng1309) ) ;
 assign wire8428 = ( (~ ng1315)  &  (~ ng1309)  &  ng1266 ) ;
 assign wire8430 = ( ng1270  &  ng1272  &  ng1271 ) ;
 assign wire8431 = ( (~ ng1315)  &  ng1272  &  ng1271 ) ;
 assign wire8432 = ( (~ ng1312)  &  ng1270  &  ng1271 ) ;
 assign wire8433 = ( (~ ng1309)  &  ng1270  &  ng1272 ) ;
 assign wire8434 = ( (~ ng1312)  &  (~ ng1315)  &  ng1271 ) ;
 assign wire8435 = ( (~ ng1312)  &  (~ ng1309)  &  ng1270 ) ;
 assign wire8436 = ( (~ ng1315)  &  (~ ng1309)  &  ng1272 ) ;
 assign wire8439 = ( (~ wire31471)  &  wire32292 ) | ( (~ wire31472)  &  wire32292 ) | ( (~ wire31471)  &  wire32293 ) | ( (~ wire31472)  &  wire32293 ) ;
 assign wire8440 = ( (~ wire31471)  &  wire32282 ) | ( (~ wire31472)  &  wire32282 ) | ( (~ wire31471)  &  wire32283 ) | ( (~ wire31472)  &  wire32283 ) ;
 assign wire8441 = ( (~ ng1309)  &  (~ ng1294)  &  (~ ng1297) ) ;
 assign wire8446 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1297) ) ;
 assign wire8447 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1294) ) ;
 assign wire8449 = ( (~ ng1183)  &  (~ ng1180)  &  (~ ng1177) ) ;
 assign wire8450 = ( (~ ng1315)  &  (~ ng1180)  &  (~ ng1177) ) ;
 assign wire8451 = ( (~ ng1312)  &  (~ ng1183)  &  (~ ng1177) ) ;
 assign wire8452 = ( (~ ng1309)  &  (~ ng1183)  &  (~ ng1180) ) ;
 assign wire8453 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1177) ) ;
 assign wire8454 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1183) ) ;
 assign wire8455 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1180) ) ;
 assign wire8457 = ( (~ ng1303)  &  (~ ng1315)  &  (~ ng1300) ) ;
 assign wire8460 = ( (~ ng1303)  &  (~ ng1306)  &  (~ ng1309) ) ;
 assign wire8461 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1300) ) ;
 assign wire8462 = ( (~ ng1306)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire8463 = ( (~ ng1303)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8469 = ( (~ ng1125)  &  (~ ng853)  &  (~ ng1128) ) ;
 assign wire8474 = ( (~ ng1125)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8475 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1128) ) ;
 assign wire8482 = ( (~ ng15970)  &  ng22396 ) | ( (~ ng15970)  &  wire32093 ) | ( (~ ng15970)  &  (~ ng22396)  &  wire32092 ) ;
 assign wire8484 = ( ng823  &  wire8487 ) | ( ng823  &  wire3150  &  wire32248 ) ;
 assign wire8487 = ( (~ wire8594)  &  (~ wire32093)  &  wire32249 ) ;
 assign wire8488 = ( (~ ng13165)  &  (~ wire32243)  &  (~ wire32244)  &  wire32245 ) ;
 assign wire8491 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32229 ) ;
 assign wire8492 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32231 ) ;
 assign wire8493 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32233 ) ;
 assign wire8494 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32235 ) ;
 assign wire8495 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32236 ) ;
 assign wire8496 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32237 ) ;
 assign wire8497 = ( ng2257  &  (~ ng11870)  &  (~ ng25082)  &  wire32238 ) ;
 assign wire8498 = ( ng2257  &  wire3046  &  (~ ng11870)  &  (~ ng25082) ) ;
 assign wire8502 = ( (~ ng1107)  &  (~ ng1104)  &  (~ ng1110) ) ;
 assign wire8503 = ( (~ ng823)  &  (~ ng1104)  &  (~ ng1110) ) ;
 assign wire8504 = ( (~ ng826)  &  (~ ng1107)  &  (~ ng1110) ) ;
 assign wire8505 = ( (~ ng853)  &  (~ ng1107)  &  (~ ng1104) ) ;
 assign wire8506 = ( (~ ng826)  &  (~ ng823)  &  (~ ng1110) ) ;
 assign wire8507 = ( (~ ng823)  &  (~ ng853)  &  (~ ng1104) ) ;
 assign wire8508 = ( (~ ng826)  &  (~ ng853)  &  (~ ng1107) ) ;
 assign wire8510 = ( (~ ng1095)  &  (~ ng1098)  &  (~ ng853) ) ;
 assign wire8515 = ( (~ ng1095)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8516 = ( (~ ng1098)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8524 = ( (~ ng826)  &  ng1033  &  ng1030 ) ;
 assign wire8529 = ( ng1041  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8530 = ( (~ ng826)  &  (~ ng853)  &  ng1030 ) ;
 assign wire8532 = ( ng1063  &  ng1071  &  ng1060 ) ;
 assign wire8533 = ( ng1063  &  (~ ng826)  &  ng1060 ) ;
 assign wire8534 = ( ng1063  &  (~ ng823)  &  ng1071 ) ;
 assign wire8535 = ( (~ ng853)  &  ng1071  &  ng1060 ) ;
 assign wire8536 = ( ng1063  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8537 = ( (~ ng823)  &  (~ ng853)  &  ng1071 ) ;
 assign wire8538 = ( (~ ng826)  &  (~ ng853)  &  ng1060 ) ;
 assign wire8540 = ( ng1048  &  (~ ng826)  &  ng1045 ) ;
 assign wire8543 = ( ng1056  &  ng1045  &  (~ ng853) ) ;
 assign wire8544 = ( ng1048  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8545 = ( ng1056  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8546 = ( (~ ng826)  &  ng1045  &  (~ ng853) ) ;
 assign wire8556 = ( (~ ng26925)  &  (~ wire32142)  &  (~ wire32155)  &  wire32156 ) ;
 assign wire8557 = ( (~ ng26925)  &  (~ wire32142)  &  (~ wire32155)  &  wire32157 ) ;
 assign wire8566 = ( (~ ng28529)  &  (~ ng11647)  &  wire31817  &  wire32147 ) ;
 assign wire8569 = ( ng805  &  wire32131 ) | ( ng805  &  ng27850  &  wire32130 ) ;
 assign wire8591 = ( (~ ng1010)  &  ng823 ) ;
 assign wire8594 = ( (~ ng1091)  &  ng823  &  (~ wire32088)  &  (~ wire32089) ) ;
 assign wire8596 = ( ng11647  &  (~ wire32088)  &  (~ wire32089)  &  wire32128 ) ;
 assign wire8597 = ( (~ ng18096)  &  (~ ng18492)  &  wire3056 ) | ( (~ ng17998)  &  (~ ng18492)  &  wire3056 ) ;
 assign wire8602 = ( (~ ng17998)  &  wire3056  &  wire3107 ) ;
 assign wire8603 = ( (~ ng18096)  &  (~ ng18492)  &  wire3107 ) ;
 assign wire8604 = ( (~ ng18096)  &  (~ ng17998)  &  wire3107 ) ;
 assign wire8619 = ( (~ ng18363)  &  (~ ng18441)  &  (~ ng18290) ) | ( (~ ng18441)  &  (~ ng18195)  &  (~ ng18290) ) ;
 assign wire8624 = ( (~ ng18363)  &  (~ ng18290)  &  wire3067 ) ;
 assign wire8625 = ( (~ ng18441)  &  (~ ng18195)  &  wire3067 ) ;
 assign wire8626 = ( (~ ng18363)  &  (~ ng18195)  &  wire3067 ) ;
 assign wire8641 = ( (~ wire32020)  &  (~ wire32021)  &  wire32023 ) ;
 assign wire8649 = ( ng826  &  (~ ng842)  &  (~ ng809) ) ;
 assign wire8650 = ( ng823  &  (~ ng843)  &  (~ ng809) ) ;
 assign wire8663 = ( ng857  &  ng858  &  (~ ng853) ) ;
 assign wire8668 = ( ng857  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8669 = ( (~ ng826)  &  ng858  &  (~ ng853) ) ;
 assign wire8671 = ( ng839  &  ng840  &  (~ ng853) ) ;
 assign wire8676 = ( ng839  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8677 = ( ng840  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8679 = ( ng860  &  ng861  &  (~ ng853) ) ;
 assign wire8684 = ( ng860  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8685 = ( ng861  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8689 = ( ng830  &  ng831  &  (~ ng853)  &  ng793 ) ;
 assign wire8690 = ( ng831  &  (~ ng826)  &  ng829  &  ng793 ) ;
 assign wire8691 = ( (~ ng853)  &  ng834  &  ng833  &  ng797 ) ;
 assign wire8692 = ( (~ ng826)  &  ng834  &  ng832  &  ng797 ) ;
 assign wire8693 = ( (~ ng826)  &  (~ ng823)  &  ng829  &  ng793 ) ;
 assign wire8694 = ( (~ ng826)  &  (~ ng823)  &  ng832  &  ng797 ) ;
 assign wire8695 = ( ng830  &  (~ ng823)  &  (~ ng853)  &  ng793 ) ;
 assign wire8696 = ( (~ ng823)  &  (~ ng853)  &  ng833  &  ng797 ) ;
 assign wire8697 = ( ng831  &  (~ ng826)  &  (~ ng853)  &  ng793 ) ;
 assign wire8698 = ( (~ ng826)  &  (~ ng853)  &  ng834  &  ng797 ) ;
 assign wire8699 = ( ng853  &  (~ ng829)  &  (~ ng793) ) ;
 assign wire8700 = ( (~ ng830)  &  ng826  &  (~ ng793) ) ;
 assign wire8701 = ( ng826  &  (~ ng833)  &  (~ ng797) ) ;
 assign wire8702 = ( ng853  &  (~ ng832)  &  (~ ng797) ) ;
 assign wire8703 = ( ng823  &  (~ ng834)  &  (~ ng797) ) ;
 assign wire8704 = ( (~ ng831)  &  ng823  &  (~ ng793) ) ;
 assign wire8705 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng793 ) ;
 assign wire8706 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng797 ) ;
 assign wire8709 = ( (~ ng785)  &  (~ wire31976)  &  (~ wire31977) ) ;
 assign wire8710 = ( ng785  &  wire31976 ) | ( ng785  &  wire31977 ) ;
 assign wire8713 = ( ng821  &  ng822  &  (~ ng853) ) ;
 assign wire8718 = ( ng821  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8719 = ( ng822  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8721 = ( (~ ng853)  &  ng819  &  ng818 ) ;
 assign wire8726 = ( (~ ng823)  &  (~ ng853)  &  ng818 ) ;
 assign wire8727 = ( (~ ng826)  &  (~ ng853)  &  ng819 ) ;
 assign wire8729 = ( ng836  &  ng837  &  (~ ng853) ) ;
 assign wire8734 = ( ng836  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8735 = ( ng837  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8737 = ( ng849  &  ng848  &  (~ ng853) ) ;
 assign wire8738 = ( ng849  &  ng847  &  (~ ng826) ) ;
 assign wire8739 = ( ng848  &  ng847  &  (~ ng823) ) ;
 assign wire8740 = ( ng849  &  ng848  &  ng847 ) ;
 assign wire8741 = ( ng847  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8742 = ( ng848  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8743 = ( ng849  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8745 = ( ng846  &  (~ ng853)  &  ng845 ) ;
 assign wire8750 = ( (~ ng823)  &  (~ ng853)  &  ng845 ) ;
 assign wire8751 = ( ng846  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8754 = ( (~ ng25958)  &  wire31920  &  wire31921  &  wire31925 ) ;
 assign wire8757 = ( (~ ng882)  &  (~ ng885)  &  (~ ng853) ) ;
 assign wire8762 = ( (~ ng882)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8763 = ( (~ ng885)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8765 = ( (~ ng912)  &  (~ ng909)  &  (~ ng853) ) ;
 assign wire8770 = ( (~ ng909)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8771 = ( (~ ng912)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8773 = ( (~ ng853)  &  (~ ng927)  &  (~ ng930) ) ;
 assign wire8774 = ( (~ ng826)  &  (~ ng930)  &  (~ ng933) ) ;
 assign wire8775 = ( (~ ng823)  &  (~ ng927)  &  (~ ng933) ) ;
 assign wire8776 = ( (~ ng927)  &  (~ ng930)  &  (~ ng933) ) ;
 assign wire8777 = ( (~ ng826)  &  (~ ng823)  &  (~ ng933) ) ;
 assign wire8778 = ( (~ ng823)  &  (~ ng853)  &  (~ ng927) ) ;
 assign wire8779 = ( (~ ng826)  &  (~ ng853)  &  (~ ng930) ) ;
 assign wire8781 = ( (~ ng900)  &  (~ ng853)  &  (~ ng903) ) ;
 assign wire8786 = ( (~ ng900)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8787 = ( (~ ng826)  &  (~ ng853)  &  (~ ng903) ) ;
 assign wire8789 = ( (~ ng939)  &  (~ ng936)  &  (~ ng853) ) ;
 assign wire8790 = ( (~ ng939)  &  (~ ng942)  &  (~ ng826) ) ;
 assign wire8791 = ( (~ ng936)  &  (~ ng942)  &  (~ ng823) ) ;
 assign wire8792 = ( (~ ng939)  &  (~ ng936)  &  (~ ng942) ) ;
 assign wire8793 = ( (~ ng942)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8794 = ( (~ ng936)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8795 = ( (~ ng939)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8797 = ( (~ ng876)  &  (~ ng873)  &  (~ ng853) ) ;
 assign wire8802 = ( (~ ng873)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8803 = ( (~ ng876)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8805 = ( (~ ng921)  &  (~ ng918)  &  (~ ng853) ) ;
 assign wire8806 = ( (~ ng924)  &  (~ ng921)  &  (~ ng826) ) ;
 assign wire8807 = ( (~ ng924)  &  (~ ng918)  &  (~ ng823) ) ;
 assign wire8808 = ( (~ ng924)  &  (~ ng921)  &  (~ ng918) ) ;
 assign wire8809 = ( (~ ng924)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8810 = ( (~ ng918)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8811 = ( (~ ng921)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8813 = ( (~ ng853)  &  (~ ng948)  &  (~ ng945) ) ;
 assign wire8818 = ( (~ ng823)  &  (~ ng853)  &  (~ ng945) ) ;
 assign wire8819 = ( (~ ng826)  &  (~ ng853)  &  (~ ng948) ) ;
 assign wire8821 = ( (~ ng954)  &  (~ ng957)  &  (~ ng853) ) ;
 assign wire8822 = ( (~ ng957)  &  (~ ng826)  &  (~ ng960) ) ;
 assign wire8823 = ( (~ ng954)  &  (~ ng823)  &  (~ ng960) ) ;
 assign wire8824 = ( (~ ng954)  &  (~ ng957)  &  (~ ng960) ) ;
 assign wire8825 = ( (~ ng826)  &  (~ ng823)  &  (~ ng960) ) ;
 assign wire8826 = ( (~ ng954)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8827 = ( (~ ng957)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8829 = ( ng1007  &  ng1006  &  ng1005 ) ;
 assign wire8830 = ( (~ ng853)  &  ng1006  &  ng1005 ) ;
 assign wire8831 = ( (~ ng823)  &  ng1007  &  ng1005 ) ;
 assign wire8834 = ( (~ ng823)  &  (~ ng853)  &  ng1005 ) ;
 assign wire8835 = ( (~ ng826)  &  (~ ng853)  &  ng1006 ) ;
 assign wire8837 = ( ng1003  &  (~ ng826)  &  ng1004 ) ;
 assign wire8840 = ( ng1002  &  ng1003  &  (~ ng853) ) ;
 assign wire8841 = ( (~ ng826)  &  (~ ng823)  &  ng1004 ) ;
 assign wire8842 = ( ng1002  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8843 = ( ng1003  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8845 = ( ng1000  &  ng999  &  (~ ng853) ) ;
 assign wire8846 = ( ng1000  &  ng1001  &  (~ ng826) ) ;
 assign wire8847 = ( ng1001  &  ng999  &  (~ ng823) ) ;
 assign wire8848 = ( ng1000  &  ng1001  &  ng999 ) ;
 assign wire8849 = ( ng1001  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire8850 = ( ng999  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8851 = ( ng1000  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8853 = ( (~ ng894)  &  (~ ng853)  &  (~ ng891) ) ;
 assign wire8858 = ( (~ ng823)  &  (~ ng853)  &  (~ ng891) ) ;
 assign wire8859 = ( (~ ng894)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire8865 = ( ng863  &  (~ ng853)  &  ng864 ) ;
 assign wire8870 = ( ng863  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire8871 = ( (~ ng826)  &  (~ ng853)  &  ng864 ) ;
 assign wire8879 = ( wire31741  &  wire31746 ) | ( wire31742  &  wire31746 ) | ( wire31743  &  wire31746 ) ;
 assign wire8880 = ( wire31741  &  wire31748 ) | ( wire31742  &  wire31748 ) | ( wire31743  &  wire31748 ) ;
 assign wire8881 = ( wire31741  &  wire31750 ) | ( wire31742  &  wire31750 ) | ( wire31743  &  wire31750 ) ;
 assign wire8882 = ( wire31741  &  wire31752 ) | ( wire31742  &  wire31752 ) | ( wire31743  &  wire31752 ) ;
 assign wire8883 = ( wire31741  &  wire31753 ) | ( wire31742  &  wire31753 ) | ( wire31743  &  wire31753 ) ;
 assign wire8884 = ( wire31741  &  wire31754 ) | ( wire31742  &  wire31754 ) | ( wire31743  &  wire31754 ) ;
 assign wire8885 = ( wire31741  &  wire31755 ) | ( wire31742  &  wire31755 ) | ( wire31743  &  wire31755 ) ;
 assign wire8886 = ( wire3049  &  wire31741 ) | ( wire3049  &  wire31742 ) | ( wire3049  &  wire31743 ) ;
 assign wire8907 = ( ng732  &  ng733  &  ng731 ) ;
 assign wire8908 = ( (~ ng1309)  &  ng733  &  ng731 ) ;
 assign wire8909 = ( (~ ng1312)  &  ng732  &  ng731 ) ;
 assign wire8912 = ( (~ ng1312)  &  (~ ng1309)  &  ng731 ) ;
 assign wire8913 = ( (~ ng1315)  &  (~ ng1309)  &  ng733 ) ;
 assign wire8915 = ( (~ ng1312)  &  ng710  &  ng711 ) ;
 assign wire8918 = ( ng712  &  ng710  &  (~ ng1309) ) ;
 assign wire8919 = ( (~ ng1312)  &  (~ ng1315)  &  ng711 ) ;
 assign wire8920 = ( (~ ng1312)  &  ng710  &  (~ ng1309) ) ;
 assign wire8921 = ( ng712  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8923 = ( ng718  &  ng716  &  ng717 ) ;
 assign wire8924 = ( (~ ng1312)  &  ng716  &  ng717 ) ;
 assign wire8925 = ( (~ ng1315)  &  ng718  &  ng717 ) ;
 assign wire8926 = ( (~ ng1309)  &  ng718  &  ng716 ) ;
 assign wire8927 = ( (~ ng1312)  &  (~ ng1315)  &  ng717 ) ;
 assign wire8928 = ( (~ ng1312)  &  (~ ng1309)  &  ng716 ) ;
 assign wire8929 = ( (~ ng1315)  &  (~ ng1309)  &  ng718 ) ;
 assign wire8931 = ( ng698  &  ng700  &  ng699 ) ;
 assign wire8932 = ( (~ ng1315)  &  ng700  &  ng699 ) ;
 assign wire8933 = ( (~ ng1312)  &  ng698  &  ng699 ) ;
 assign wire8934 = ( (~ ng1309)  &  ng698  &  ng700 ) ;
 assign wire8935 = ( (~ ng1312)  &  (~ ng1315)  &  ng699 ) ;
 assign wire8936 = ( (~ ng1312)  &  (~ ng1309)  &  ng698 ) ;
 assign wire8937 = ( (~ ng1315)  &  (~ ng1309)  &  ng700 ) ;
 assign wire8939 = ( ng707  &  ng709  &  ng708 ) ;
 assign wire8940 = ( (~ ng1315)  &  ng709  &  ng708 ) ;
 assign wire8941 = ( (~ ng1312)  &  ng707  &  ng708 ) ;
 assign wire8942 = ( (~ ng1309)  &  ng707  &  ng709 ) ;
 assign wire8943 = ( (~ ng1312)  &  (~ ng1315)  &  ng708 ) ;
 assign wire8944 = ( (~ ng1312)  &  (~ ng1309)  &  ng707 ) ;
 assign wire8945 = ( (~ ng1315)  &  (~ ng1309)  &  ng709 ) ;
 assign wire8947 = ( ng703  &  ng701  &  (~ ng1309) ) ;
 assign wire8952 = ( (~ ng1312)  &  ng701  &  (~ ng1309) ) ;
 assign wire8953 = ( ng703  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8955 = ( ng725  &  ng727  &  ng726 ) ;
 assign wire8956 = ( (~ ng1315)  &  ng727  &  ng726 ) ;
 assign wire8957 = ( (~ ng1312)  &  ng725  &  ng726 ) ;
 assign wire8958 = ( (~ ng1309)  &  ng725  &  ng727 ) ;
 assign wire8959 = ( (~ ng1312)  &  (~ ng1315)  &  ng726 ) ;
 assign wire8960 = ( (~ ng1312)  &  (~ ng1309)  &  ng725 ) ;
 assign wire8961 = ( (~ ng1315)  &  (~ ng1309)  &  ng727 ) ;
 assign wire8963 = ( (~ ng1309)  &  ng704  &  ng706 ) ;
 assign wire8968 = ( (~ ng1312)  &  (~ ng1309)  &  ng704 ) ;
 assign wire8969 = ( (~ ng1315)  &  (~ ng1309)  &  ng706 ) ;
 assign wire8971 = ( ng719  &  ng721  &  ng720 ) ;
 assign wire8972 = ( (~ ng1315)  &  ng721  &  ng720 ) ;
 assign wire8973 = ( (~ ng1312)  &  ng719  &  ng720 ) ;
 assign wire8974 = ( ng719  &  (~ ng1309)  &  ng721 ) ;
 assign wire8975 = ( (~ ng1312)  &  (~ ng1315)  &  ng720 ) ;
 assign wire8976 = ( (~ ng1312)  &  ng719  &  (~ ng1309) ) ;
 assign wire8977 = ( (~ ng1315)  &  (~ ng1309)  &  ng721 ) ;
 assign wire8979 = ( ng715  &  (~ ng1309)  &  ng713 ) ;
 assign wire8984 = ( (~ ng1312)  &  (~ ng1309)  &  ng713 ) ;
 assign wire8985 = ( ng715  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire8987 = ( ng722  &  ng724  &  (~ ng1309) ) ;
 assign wire8988 = ( ng724  &  ng723  &  (~ ng1315) ) ;
 assign wire8989 = ( ng722  &  ng723  &  (~ ng1312) ) ;
 assign wire8990 = ( ng722  &  ng724  &  ng723 ) ;
 assign wire8991 = ( ng723  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire8992 = ( ng722  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire8993 = ( ng724  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire9005 = ( wire3221  &  (~ wire31587)  &  (~ wire31588)  &  (~ wire31589) ) ;
 assign wire9007 = ( (~ ng590)  &  (~ ng593)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire9008 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng587)  &  (~ ng185) ) ;
 assign wire9009 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng587)  &  (~ ng185) ) ;
 assign wire9010 = ( (~ ng590)  &  (~ ng593)  &  (~ ng587)  &  (~ ng185) ) ;
 assign wire9011 = ( (~ ng590)  &  (~ ng593)  &  (~ ng1309)  &  (~ ng524) ) ;
 assign wire9012 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng587)  &  (~ ng524) ) ;
 assign wire9013 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng587)  &  (~ ng524) ) ;
 assign wire9014 = ( (~ ng590)  &  (~ ng593)  &  (~ ng587)  &  (~ ng524) ) ;
 assign wire9015 = ( wire31550  &  wire31553 ) | ( wire31551  &  wire31553 ) ;
 assign wire9019 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng587)  &  (~ ng185) ) ;
 assign wire9020 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng587)  &  (~ ng524) ) ;
 assign wire9022 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire9023 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng1309)  &  (~ ng524) ) ;
 assign wire9025 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire9026 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng524) ) ;
 assign wire9028 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng185) ) ;
 assign wire9029 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1309)  &  (~ ng524) ) ;
 assign wire9030 = ( wire3049  &  wire31550 ) | ( wire3049  &  wire31551 ) ;
 assign wire9031 = ( (~ ng573)  &  (~ ng571)  &  (~ ng569) ) ;
 assign wire9032 = ( (~ ng1315)  &  (~ ng571)  &  (~ ng569) ) ;
 assign wire9033 = ( (~ ng1312)  &  (~ ng573)  &  (~ ng569) ) ;
 assign wire9034 = ( (~ ng573)  &  (~ ng1309)  &  (~ ng571) ) ;
 assign wire9035 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng569) ) ;
 assign wire9036 = ( (~ ng1312)  &  (~ ng573)  &  (~ ng1309) ) ;
 assign wire9037 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng571) ) ;
 assign wire9041 = ( ng12145  &  ng12080  &  wire31514 ) | ( (~ ng12145)  &  wire3118  &  wire31514 ) | ( ng12080  &  wire3118  &  wire31514 ) ;
 assign wire9044 = ( pg3229  &  (~ wire31482)  &  (~ wire31483) ) ;
 assign wire9049 = ( ng580  &  (~ ng1309)  &  ng578 ) ;
 assign wire9054 = ( (~ ng1312)  &  (~ ng1309)  &  ng578 ) ;
 assign wire9055 = ( ng580  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire9057 = ( ng577  &  (~ ng1315)  &  ng576 ) ;
 assign wire9060 = ( ng575  &  ng577  &  (~ ng1309) ) ;
 assign wire9061 = ( (~ ng1312)  &  (~ ng1315)  &  ng576 ) ;
 assign wire9062 = ( ng575  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire9063 = ( ng577  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire9065 = ( (~ ng1315)  &  ng585  &  ng586 ) ;
 assign wire9070 = ( ng584  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire9071 = ( (~ ng1315)  &  (~ ng1309)  &  ng586 ) ;
 assign wire9073 = ( ng582  &  ng583  &  ng581 ) ;
 assign wire9074 = ( (~ ng1309)  &  ng583  &  ng581 ) ;
 assign wire9075 = ( (~ ng1312)  &  ng582  &  ng581 ) ;
 assign wire9078 = ( (~ ng1312)  &  (~ ng1309)  &  ng581 ) ;
 assign wire9079 = ( (~ ng1315)  &  (~ ng1309)  &  ng583 ) ;
 assign wire9082 = ( wire31469  &  (~ wire31471) ) | ( wire31470  &  (~ wire31471) ) | ( wire31469  &  (~ wire31472) ) | ( wire31470  &  (~ wire31472) ) ;
 assign wire9083 = ( wire31459  &  (~ wire31471) ) | ( wire31460  &  (~ wire31471) ) | ( wire31459  &  (~ wire31472) ) | ( wire31460  &  (~ wire31472) ) ;
 assign wire9084 = ( (~ ng611)  &  (~ ng608)  &  (~ ng1309) ) ;
 assign wire9085 = ( (~ ng608)  &  (~ ng1315)  &  (~ ng605) ) ;
 assign wire9086 = ( (~ ng611)  &  (~ ng1312)  &  (~ ng605) ) ;
 assign wire9087 = ( (~ ng611)  &  (~ ng608)  &  (~ ng605) ) ;
 assign wire9088 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng605) ) ;
 assign wire9089 = ( (~ ng611)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire9090 = ( (~ ng608)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire9092 = ( (~ ng1309)  &  (~ ng493)  &  (~ ng496) ) ;
 assign wire9097 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng496) ) ;
 assign wire9098 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng493) ) ;
 assign wire9100 = ( (~ ng620)  &  (~ ng617)  &  (~ ng614) ) ;
 assign wire9101 = ( (~ ng1312)  &  (~ ng620)  &  (~ ng614) ) ;
 assign wire9102 = ( (~ ng1315)  &  (~ ng617)  &  (~ ng614) ) ;
 assign wire9103 = ( (~ ng1309)  &  (~ ng620)  &  (~ ng617) ) ;
 assign wire9104 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng614) ) ;
 assign wire9105 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng620) ) ;
 assign wire9106 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng617) ) ;
 assign wire9118 = ( (~ ng23486)  &  ng11624  &  (~ wire31067) ) | ( ng11624  &  (~ ng23478)  &  (~ wire31067) ) ;
 assign wire9128 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire31418 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire31418 ) ;
 assign wire9129 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire31419 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire31419 ) ;
 assign wire9130 = ( (~ ng11975)  &  ng17985  &  ng11935  &  wire31420 ) | ( ng11975  &  (~ ng17985)  &  (~ ng11935)  &  wire31420 ) ;
 assign wire9134 = ( (~ ng441)  &  (~ ng853)  &  (~ ng438) ) ;
 assign wire9139 = ( (~ ng823)  &  (~ ng853)  &  (~ ng438) ) ;
 assign wire9140 = ( (~ ng441)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9142 = ( (~ ng429)  &  (~ ng432)  &  (~ ng435) ) ;
 assign wire9143 = ( (~ ng826)  &  (~ ng432)  &  (~ ng435) ) ;
 assign wire9144 = ( (~ ng429)  &  (~ ng823)  &  (~ ng435) ) ;
 assign wire9145 = ( (~ ng429)  &  (~ ng853)  &  (~ ng432) ) ;
 assign wire9146 = ( (~ ng826)  &  (~ ng823)  &  (~ ng435) ) ;
 assign wire9147 = ( (~ ng429)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9148 = ( (~ ng826)  &  (~ ng853)  &  (~ ng432) ) ;
 assign wire9150 = ( (~ ng826)  &  ng179  &  ng177 ) ;
 assign wire9153 = ( ng178  &  ng179  &  (~ ng853) ) ;
 assign wire9154 = ( (~ ng826)  &  (~ ng823)  &  ng177 ) ;
 assign wire9155 = ( ng178  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9156 = ( (~ ng826)  &  ng179  &  (~ ng853) ) ;
 assign wire9165 = ( (~ ng11781)  &  ng25078  &  (~ wire31362)  &  wire31365 ) ;
 assign wire9167 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31368 ) ;
 assign wire9168 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31370 ) ;
 assign wire9169 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31372 ) ;
 assign wire9170 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31374 ) ;
 assign wire9171 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31375 ) ;
 assign wire9172 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31376 ) ;
 assign wire9173 = ( ng2257  &  (~ ng11828)  &  (~ ng25078)  &  wire31377 ) ;
 assign wire9174 = ( ng2257  &  wire3046  &  (~ ng11828)  &  (~ ng25078) ) ;
 assign wire9178 = ( (~ ng423)  &  (~ ng420)  &  (~ ng417) ) ;
 assign wire9179 = ( (~ ng853)  &  (~ ng420)  &  (~ ng417) ) ;
 assign wire9180 = ( (~ ng823)  &  (~ ng423)  &  (~ ng417) ) ;
 assign wire9183 = ( (~ ng823)  &  (~ ng853)  &  (~ ng417) ) ;
 assign wire9184 = ( (~ ng826)  &  (~ ng853)  &  (~ ng420) ) ;
 assign wire9186 = ( (~ ng411)  &  (~ ng408)  &  (~ ng853) ) ;
 assign wire9187 = ( (~ ng414)  &  (~ ng411)  &  (~ ng826) ) ;
 assign wire9188 = ( (~ ng414)  &  (~ ng408)  &  (~ ng823) ) ;
 assign wire9189 = ( (~ ng414)  &  (~ ng411)  &  (~ ng408) ) ;
 assign wire9190 = ( (~ ng414)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire9191 = ( (~ ng408)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9192 = ( (~ ng411)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9202 = ( ng343  &  ng354  &  (~ ng853) ) ;
 assign wire9207 = ( ng354  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9208 = ( ng343  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9210 = ( ng373  &  ng384  &  (~ ng853) ) ;
 assign wire9215 = ( ng384  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9216 = ( ng373  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9218 = ( ng358  &  ng361  &  (~ ng826) ) ;
 assign wire9221 = ( ng369  &  ng358  &  (~ ng853) ) ;
 assign wire9222 = ( ng361  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire9223 = ( ng369  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9224 = ( ng358  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9238 = ( (~ ng28501)  &  ng26902  &  (~ wire31008)  &  (~ wire31009) ) ;
 assign wire9239 = ( ng125  &  wire31274 ) | ( ng125  &  ng27834  &  wire31273 ) ;
 assign wire9260 = ( (~ ng323)  &  ng823 ) ;
 assign wire9263 = ( (~ ng404)  &  ng823  &  (~ wire31231)  &  (~ wire31232) ) ;
 assign wire9265 = ( ng11624  &  (~ wire31231)  &  (~ wire31232)  &  wire31271 ) ;
 assign wire9266 = ( (~ ng18419)  &  (~ ng17807)  &  (~ ng17729) ) | ( (~ ng17887)  &  (~ ng17807)  &  (~ ng17729) ) ;
 assign wire9271 = ( (~ ng17887)  &  (~ ng17729)  &  wire3106 ) ;
 assign wire9272 = ( (~ ng18419)  &  (~ ng17807)  &  wire3106 ) ;
 assign wire9273 = ( (~ ng18419)  &  (~ ng17887)  &  wire3106 ) ;
 assign wire9288 = ( (~ ng18079)  &  (~ ng18183)  &  wire3054 ) | ( (~ ng18183)  &  (~ ng18346)  &  wire3054 ) ;
 assign wire9293 = ( (~ ng18079)  &  wire3054  &  wire3065 ) ;
 assign wire9294 = ( (~ ng18183)  &  (~ ng18346)  &  wire3065 ) ;
 assign wire9295 = ( (~ ng18079)  &  (~ ng18346)  &  wire3065 ) ;
 assign wire9313 = ( (~ wire31159)  &  (~ wire31160)  &  wire31162 ) ;
 assign wire9318 = ( ng823  &  (~ ng152)  &  (~ ng117) ) ;
 assign wire9319 = ( ng853  &  (~ ng150)  &  (~ ng117) ) ;
 assign wire9332 = ( ng170  &  ng169  &  (~ ng853) ) ;
 assign wire9337 = ( ng169  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9338 = ( ng170  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9340 = ( ng158  &  ng157  &  (~ ng853) ) ;
 assign wire9345 = ( ng157  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9346 = ( ng158  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9356 = ( ng853  &  (~ ng132)  &  (~ ng101) ) ;
 assign wire9357 = ( (~ ng134)  &  ng823  &  (~ ng101) ) ;
 assign wire9358 = ( ng853  &  (~ ng147)  &  (~ ng113) ) ;
 assign wire9359 = ( ng826  &  (~ ng148)  &  (~ ng113) ) ;
 assign wire9360 = ( (~ ng149)  &  ng823  &  (~ ng113) ) ;
 assign wire9364 = ( (~ ng109)  &  (~ wire31115)  &  (~ wire31116) ) ;
 assign wire9365 = ( ng109  &  wire31115 ) | ( ng109  &  wire31116 ) ;
 assign wire9368 = ( (~ ng853)  &  ng142  &  ng143 ) ;
 assign wire9373 = ( (~ ng823)  &  (~ ng853)  &  ng142 ) ;
 assign wire9374 = ( (~ ng826)  &  (~ ng853)  &  ng143 ) ;
 assign wire9376 = ( ng145  &  ng146  &  (~ ng853) ) ;
 assign wire9381 = ( ng145  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9382 = ( ng146  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9384 = ( ng130  &  ng131  &  (~ ng853) ) ;
 assign wire9389 = ( ng130  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9390 = ( ng131  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9392 = ( ng155  &  ng154  &  (~ ng853) ) ;
 assign wire9393 = ( ng155  &  ng153  &  (~ ng826) ) ;
 assign wire9394 = ( ng154  &  ng153  &  (~ ng823) ) ;
 assign wire9395 = ( ng155  &  ng154  &  ng153 ) ;
 assign wire9396 = ( ng153  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire9397 = ( ng154  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9398 = ( ng155  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9400 = ( (~ ng826)  &  ng171  &  ng173 ) ;
 assign wire9405 = ( ng172  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9406 = ( (~ ng826)  &  (~ ng853)  &  ng173 ) ;
 assign wire9408 = ( ng164  &  (~ ng853)  &  ng163 ) ;
 assign wire9413 = ( (~ ng823)  &  (~ ng853)  &  ng163 ) ;
 assign wire9414 = ( ng164  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9416 = ( ng176  &  (~ ng853)  &  ng175 ) ;
 assign wire9421 = ( (~ ng823)  &  (~ ng853)  &  ng175 ) ;
 assign wire9422 = ( (~ ng826)  &  ng176  &  (~ ng853) ) ;
 assign wire9425 = ( (~ ng25954)  &  wire31061  &  wire31062  &  wire31066 ) ;
 assign wire9429 = ( ng312  &  (~ ng853)  &  ng313 ) ;
 assign wire9434 = ( ng312  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9435 = ( (~ ng826)  &  (~ ng853)  &  ng313 ) ;
 assign wire9437 = ( ng318  &  ng319  &  (~ ng853) ) ;
 assign wire9442 = ( ng318  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9443 = ( ng319  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9445 = ( (~ ng853)  &  ng316  &  ng315 ) ;
 assign wire9450 = ( (~ ng823)  &  (~ ng853)  &  ng315 ) ;
 assign wire9451 = ( (~ ng826)  &  (~ ng853)  &  ng316 ) ;
 assign wire9453 = ( (~ ng853)  &  (~ ng186)  &  (~ ng189) ) ;
 assign wire9458 = ( (~ ng823)  &  (~ ng853)  &  (~ ng186) ) ;
 assign wire9459 = ( (~ ng826)  &  (~ ng853)  &  (~ ng189) ) ;
 assign wire9461 = ( (~ ng826)  &  (~ ng225)  &  (~ ng228) ) ;
 assign wire9464 = ( (~ ng222)  &  (~ ng225)  &  (~ ng853) ) ;
 assign wire9465 = ( (~ ng826)  &  (~ ng823)  &  (~ ng228) ) ;
 assign wire9466 = ( (~ ng222)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9467 = ( (~ ng826)  &  (~ ng225)  &  (~ ng853) ) ;
 assign wire9469 = ( (~ ng198)  &  (~ ng826)  &  (~ ng201) ) ;
 assign wire9472 = ( (~ ng195)  &  (~ ng198)  &  (~ ng853) ) ;
 assign wire9473 = ( (~ ng826)  &  (~ ng823)  &  (~ ng201) ) ;
 assign wire9474 = ( (~ ng195)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9475 = ( (~ ng198)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9477 = ( (~ ng270)  &  (~ ng853)  &  (~ ng267) ) ;
 assign wire9482 = ( (~ ng823)  &  (~ ng853)  &  (~ ng267) ) ;
 assign wire9483 = ( (~ ng270)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9485 = ( (~ ng231)  &  (~ ng234)  &  (~ ng853) ) ;
 assign wire9490 = ( (~ ng231)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9491 = ( (~ ng234)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9493 = ( (~ ng252)  &  (~ ng249)  &  (~ ng853) ) ;
 assign wire9498 = ( (~ ng249)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9499 = ( (~ ng252)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9501 = ( (~ ng207)  &  (~ ng204)  &  (~ ng853) ) ;
 assign wire9506 = ( (~ ng204)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9507 = ( (~ ng207)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9509 = ( (~ ng240)  &  (~ ng853)  &  (~ ng243) ) ;
 assign wire9514 = ( (~ ng240)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9515 = ( (~ ng826)  &  (~ ng853)  &  (~ ng243) ) ;
 assign wire9517 = ( (~ ng258)  &  (~ ng261)  &  (~ ng853) ) ;
 assign wire9518 = ( (~ ng261)  &  (~ ng264)  &  (~ ng826) ) ;
 assign wire9519 = ( (~ ng258)  &  (~ ng264)  &  (~ ng823) ) ;
 assign wire9520 = ( (~ ng258)  &  (~ ng261)  &  (~ ng264) ) ;
 assign wire9521 = ( (~ ng264)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire9522 = ( (~ ng258)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9523 = ( (~ ng261)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9525 = ( (~ ng213)  &  (~ ng216)  &  (~ ng853) ) ;
 assign wire9530 = ( (~ ng213)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire9531 = ( (~ ng216)  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire9538 = ( ng3179  &  (~ wire3193)  &  (~ wire3247)  &  ng8430 ) ;
 assign wire9542 = ( (~ ng3135)  &  ng3161  &  ng8430  &  (~ wire30898) ) ;
 assign wire9543 = ( ng3182  &  (~ wire3247)  &  ng8430  &  (~ wire30899) ) ;
 assign wire9544 = ( (~ ng3135)  &  ng3164  &  ng8430  &  (~ wire30900) ) ;
 assign wire9547 = ( (~ ng3135)  &  ng3176  &  ng8430  &  (~ wire30903) ) ;
 assign wire9548 = ( (~ ng3135)  &  ng3173  &  ng8430  &  (~ wire30904) ) ;
 assign wire9549 = ( ng3185  &  ng8430  &  (~ wire30905) ) ;
 assign wire9550 = ( ng3135  &  (~ ng3120)  &  (~ wire3246)  &  (~ ng8381) ) ;
 assign wire9559 = ( wire30883  &  wire30884 ) | ( ng21851  &  wire30881  &  wire30884 ) ;
 assign wire30881 = ( ng1309  &  (~ ng1186) ) ;
 assign wire30883 = ( ng1186  &  ng1230 ) | ( (~ ng1186)  &  ng1234  &  (~ ng1309) ) ;
 assign wire30884 = ( (~ ng1880)  &  ng1309 ) ;
 assign wire30886 = ( ng1880  &  ng1924 ) | ( (~ ng1309)  &  (~ ng1880)  &  ng1928 ) ;
 assign wire30887 = ( (~ ng2574)  &  ng1309 ) ;
 assign wire30889 = ( ng2618  &  ng2574 ) | ( (~ ng1309)  &  (~ ng2574)  &  ng2622 ) ;
 assign wire30892 = ( ng3120 ) | ( ng3135 ) ;
 assign wire30893 = ( (~ ng3135) ) | ( ng3139 ) | ( (~ ng3120) ) | ( ng3147 ) ;
 assign wire30896 = ( ng3147 ) | ( (~ ng3139) ) ;
 assign wire30897 = ( (~ ng3147) ) | ( (~ ng3139) ) ;
 assign wire30898 = ( ng3139 ) | ( (~ ng3120) ) | ( ng3147 ) ;
 assign wire30899 = ( ng3147 ) | ( (~ ng3139) ) ;
 assign wire30900 = ( (~ ng3139) ) | ( (~ ng3120) ) | ( ng3147 ) ;
 assign wire30902 = ( (~ ng3135) ) | ( (~ ng3139) ) | ( (~ ng3120) ) | ( ng3147 ) ;
 assign wire30903 = ( (~ ng3139) ) | ( (~ ng3120) ) | ( (~ ng3147) ) ;
 assign wire30904 = ( ng3139 ) | ( (~ ng3120) ) | ( (~ ng3147) ) ;
 assign wire30905 = ( (~ ng3135) ) | ( ng3139 ) | ( (~ ng3120) ) | ( ng3147 ) ;
 assign wire30906 = ( ng17973 ) | ( ng3088  &  ng8430  &  (~ wire30902) ) ;
 assign wire30911 = ( wire30906 ) | ( ng3135  &  wire3217 ) ;
 assign wire30912 = ( ng3167  &  (~ ng15719) ) | ( ng3158  &  (~ ng15841) ) ;
 assign wire30913 = ( ng3155  &  (~ ng15830) ) | ( ng3170  &  (~ ng15757) ) ;
 assign wire30914 = ( wire9538 ) | ( wire9542 ) | ( wire9543 ) | ( wire9549 ) ;
 assign wire30915 = ( wire9544 ) | ( wire9547 ) | ( wire9548 ) | ( wire9550 ) ;
 assign wire30918 = ( wire30911 ) | ( wire30912 ) | ( wire30915 ) ;
 assign wire30924 = ( (~ ng240)  &  (~ ng823)  &  (~ ng246) ) | ( (~ ng240)  &  (~ ng246)  &  (~ ng243) ) ;
 assign wire30925 = ( (~ ng826)  &  (~ ng823)  &  (~ ng246) ) | ( (~ ng826)  &  (~ ng246)  &  (~ ng243) ) ;
 assign wire30927 = ( wire3046 ) | ( wire9509 ) | ( wire30924 ) ;
 assign wire30928 = ( wire9514 ) | ( wire9515 ) | ( wire30925 ) ;
 assign wire30934 = ( (~ ng270)  &  (~ ng273)  &  (~ ng267) ) | ( (~ ng273)  &  (~ ng823)  &  (~ ng267) ) ;
 assign wire30935 = ( (~ ng270)  &  (~ ng273)  &  (~ ng826) ) | ( (~ ng273)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire30937 = ( wire3046 ) | ( wire9477 ) | ( wire30934 ) ;
 assign wire30938 = ( wire9482 ) | ( wire9483 ) | ( wire30935 ) ;
 assign wire30944 = ( (~ ng213)  &  (~ ng216)  &  (~ ng219) ) | ( (~ ng216)  &  (~ ng219)  &  (~ ng826) ) ;
 assign wire30945 = ( (~ ng213)  &  (~ ng219)  &  (~ ng823) ) | ( (~ ng219)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire30947 = ( wire3046 ) | ( wire9525 ) | ( wire30944 ) ;
 assign wire30948 = ( wire9530 ) | ( wire9531 ) | ( wire30945 ) ;
 assign wire30954 = ( ng318  &  ng319  &  ng320 ) | ( ng319  &  (~ ng826)  &  ng320 ) ;
 assign wire30955 = ( ng318  &  ng320  &  (~ ng823) ) | ( (~ ng826)  &  ng320  &  (~ ng823) ) ;
 assign wire30957 = ( wire3046 ) | ( wire9437 ) | ( wire30954 ) ;
 assign wire30958 = ( wire9442 ) | ( wire9443 ) | ( wire30955 ) ;
 assign wire30964 = ( ng312  &  ng314  &  ng313 ) | ( (~ ng826)  &  ng314  &  ng313 ) ;
 assign wire30965 = ( ng312  &  ng314  &  (~ ng823) ) | ( (~ ng826)  &  ng314  &  (~ ng823) ) ;
 assign wire30967 = ( wire3046 ) | ( wire9429 ) | ( wire30964 ) ;
 assign wire30968 = ( wire9434 ) | ( wire9435 ) | ( wire30965 ) ;
 assign wire30974 = ( ng317  &  (~ ng823)  &  ng315 ) | ( ng317  &  ng316  &  ng315 ) ;
 assign wire30975 = ( ng317  &  (~ ng826)  &  (~ ng823) ) | ( ng317  &  (~ ng826)  &  ng316 ) ;
 assign wire30977 = ( wire3046 ) | ( wire9445 ) | ( wire30974 ) ;
 assign wire30978 = ( wire9450 ) | ( wire9451 ) | ( wire30975 ) ;
 assign wire30979 = ( wire30957  &  wire30967 ) | ( wire30958  &  wire30967 ) | ( wire30957  &  wire30968 ) | ( wire30958  &  wire30968 ) ;
 assign wire30985 = ( (~ ng207)  &  (~ ng204)  &  (~ ng210) ) | ( (~ ng207)  &  (~ ng826)  &  (~ ng210) ) ;
 assign wire30986 = ( (~ ng204)  &  (~ ng210)  &  (~ ng823) ) | ( (~ ng826)  &  (~ ng210)  &  (~ ng823) ) ;
 assign wire30988 = ( wire3046 ) | ( wire9501 ) | ( wire30985 ) ;
 assign wire30989 = ( wire9506 ) | ( wire9507 ) | ( wire30986 ) ;
 assign wire30995 = ( (~ ng255)  &  (~ ng252)  &  (~ ng249) ) | ( (~ ng255)  &  (~ ng252)  &  (~ ng826) ) ;
 assign wire30996 = ( (~ ng255)  &  (~ ng249)  &  (~ ng823) ) | ( (~ ng255)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire30998 = ( wire3046 ) | ( wire9493 ) | ( wire30995 ) ;
 assign wire30999 = ( wire9498 ) | ( wire9499 ) | ( wire30996 ) ;
 assign wire31008 = ( wire3046 ) | ( wire9517 ) | ( wire9518 ) | ( wire9519 ) ;
 assign wire31009 = ( wire9520 ) | ( wire9521 ) | ( wire9522 ) | ( wire9523 ) ;
 assign wire31015 = ( (~ ng231)  &  (~ ng234)  &  (~ ng237) ) | ( (~ ng234)  &  (~ ng826)  &  (~ ng237) ) ;
 assign wire31016 = ( (~ ng231)  &  (~ ng237)  &  (~ ng823) ) | ( (~ ng826)  &  (~ ng237)  &  (~ ng823) ) ;
 assign wire31018 = ( wire3046 ) | ( wire9485 ) | ( wire31015 ) ;
 assign wire31019 = ( wire9490 ) | ( wire9491 ) | ( wire31016 ) ;
 assign wire31025 = ( (~ ng195)  &  (~ ng198)  &  (~ ng201) ) | ( (~ ng195)  &  (~ ng823)  &  (~ ng201) ) ;
 assign wire31028 = ( wire3046 ) | ( wire9469 ) | ( wire31025 ) ;
 assign wire31029 = ( wire9472 ) | ( wire9473 ) | ( wire9474 ) | ( wire9475 ) ;
 assign wire31035 = ( (~ ng222)  &  (~ ng225)  &  (~ ng228) ) | ( (~ ng222)  &  (~ ng823)  &  (~ ng228) ) ;
 assign wire31038 = ( wire3046 ) | ( wire9461 ) | ( wire31035 ) ;
 assign wire31039 = ( wire9464 ) | ( wire9465 ) | ( wire9466 ) | ( wire9467 ) ;
 assign wire31045 = ( (~ ng192)  &  (~ ng826)  &  (~ ng189) ) | ( (~ ng192)  &  (~ ng186)  &  (~ ng189) ) ;
 assign wire31046 = ( (~ ng192)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng192)  &  (~ ng823)  &  (~ ng186) ) ;
 assign wire31048 = ( wire3046 ) | ( wire9453 ) | ( wire31045 ) ;
 assign wire31049 = ( wire9458 ) | ( wire9459 ) | ( wire31046 ) ;
 assign wire31050 = ( (~ wire30927)  &  (~ wire30928)  &  (~ wire30937)  &  (~ wire30938) ) ;
 assign wire31051 = ( wire30947  &  wire30988 ) | ( wire30948  &  wire30988 ) | ( wire30947  &  wire30989 ) | ( wire30948  &  wire30989 ) ;
 assign wire31052 = ( wire30998  &  wire31008 ) | ( wire30999  &  wire31008 ) | ( wire30998  &  wire31009 ) | ( wire30999  &  wire31009 ) ;
 assign wire31053 = ( (~ wire31018)  &  (~ wire31019)  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire31054 = ( (~ wire31038)  &  (~ wire31039)  &  wire31048 ) | ( (~ wire31038)  &  (~ wire31039)  &  wire31049 ) ;
 assign wire31057 = ( (~ wire30977)  &  (~ wire30978)  &  wire30979  &  wire31054 ) ;
 assign wire31058 = ( wire31050  &  wire31051  &  wire31052  &  wire31053 ) ;
 assign wire31059 = ( wire30927  &  wire30937 ) | ( wire30928  &  wire30937 ) | ( wire30927  &  wire30938 ) | ( wire30928  &  wire30938 ) ;
 assign wire31060 = ( wire30947  &  wire30988 ) | ( wire30948  &  wire30988 ) | ( wire30947  &  wire30989 ) | ( wire30948  &  wire30989 ) ;
 assign wire31061 = ( wire30998  &  wire31008 ) | ( wire30999  &  wire31008 ) | ( wire30998  &  wire31009 ) | ( wire30999  &  wire31009 ) ;
 assign wire31062 = ( wire31018  &  wire31028 ) | ( wire31019  &  wire31028 ) | ( wire31018  &  wire31029 ) | ( wire31019  &  wire31029 ) ;
 assign wire31063 = ( wire31038  &  wire31048 ) | ( wire31039  &  wire31048 ) | ( wire31038  &  wire31049 ) | ( wire31039  &  wire31049 ) ;
 assign wire31065 = ( wire31062  &  wire31061 ) ;
 assign wire31066 = ( wire31059  &  wire31060  &  wire31063 ) ;
 assign wire31067 = ( wire30957  &  wire30967 ) | ( wire30958  &  wire30967 ) | ( wire30957  &  wire30968 ) | ( wire30958  &  wire30968 ) ;
 assign wire31074 = ( ng168  &  ng170  &  ng169 ) | ( ng168  &  ng169  &  (~ ng823) ) ;
 assign wire31075 = ( ng168  &  ng170  &  (~ ng826) ) | ( ng168  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31077 = ( wire3046 ) | ( wire9332 ) | ( wire31074 ) ;
 assign wire31078 = ( wire9337 ) | ( wire9338 ) | ( wire31075 ) ;
 assign wire31079 = ( ng147  &  ng148 ) ;
 assign wire31081 = ( ng147  &  (~ ng826) ) ;
 assign wire31083 = ( (~ ng853)  &  ng148 ) ;
 assign wire31084 = ( ng149  &  ng113 ) | ( (~ ng823)  &  ng113 ) ;
 assign wire31085 = ( ng132  &  ng134 ) ;
 assign wire31086 = ( (~ ng826)  &  ng101 ) | ( ng133  &  ng101 ) ;
 assign wire31087 = ( ng132  &  (~ ng823) ) ;
 assign wire31089 = ( (~ ng853)  &  ng134 ) ;
 assign wire31091 = ( (~ ng826)  &  (~ ng853)  &  ng113 ) ;
 assign wire31092 = ( (~ ng823)  &  (~ ng853)  &  ng101 ) ;
 assign wire31102 = ( ng141  &  (~ ng826)  &  ng143 ) | ( ng141  &  ng142  &  ng143 ) ;
 assign wire31103 = ( ng141  &  (~ ng826)  &  (~ ng823) ) | ( ng141  &  (~ ng823)  &  ng142 ) ;
 assign wire31106 = ( wire9373 ) | ( wire9374 ) | ( wire31103 ) ;
 assign wire31112 = ( ng145  &  ng144  &  ng146 ) | ( ng144  &  ng146  &  (~ ng826) ) ;
 assign wire31113 = ( ng145  &  ng144  &  (~ ng823) ) | ( ng144  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31115 = ( wire3046 ) | ( wire9376 ) | ( wire31112 ) ;
 assign wire31116 = ( wire9381 ) | ( wire9382 ) | ( wire31113 ) ;
 assign wire31122 = ( ng130  &  ng131  &  ng129 ) | ( ng131  &  ng129  &  (~ ng826) ) ;
 assign wire31123 = ( ng130  &  ng129  &  (~ ng823) ) | ( ng129  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31126 = ( wire9389 ) | ( wire9390 ) | ( wire31123 ) ;
 assign wire31129 = ( wire9360 ) | ( ng826  &  (~ ng133)  &  (~ ng101) ) ;
 assign wire31130 = ( ng113  &  wire3308  &  wire31079 ) | ( ng113  &  wire3308  &  wire31081 ) ;
 assign wire31131 = ( wire31083  &  wire31084 ) | ( wire31085  &  wire31086 ) ;
 assign wire31132 = ( ng101  &  wire3307  &  wire31087 ) | ( ng101  &  wire3307  &  wire31089 ) ;
 assign wire31133 = ( wire3308  &  wire31091 ) | ( wire3307  &  wire31092 ) ;
 assign wire31134 = ( wire9356 ) | ( wire9357 ) | ( wire9358 ) | ( wire9359 ) ;
 assign wire31137 = ( wire31134 ) | ( wire31133 ) ;
 assign wire31138 = ( wire31129 ) | ( wire31130 ) | ( wire31131 ) | ( wire31132 ) ;
 assign wire31143 = ( wire9364 ) | ( wire31137 ) | ( ng105  &  ng11744 ) | ( (~ ng105)  &  (~ ng11744) ) ;
 assign wire31144 = ( wire9365 ) | ( wire31138 ) | ( ng97  &  ng11889 ) | ( (~ ng97)  &  (~ ng11889) ) ;
 assign wire31145 = ( ng152  &  ng150 ) ;
 assign wire31147 = ( ng152  &  (~ ng853) ) ;
 assign wire31149 = ( ng150  &  (~ ng823) ) ;
 assign wire31156 = ( ng174  &  ng176  &  ng175 ) | ( ng174  &  (~ ng823)  &  ng175 ) ;
 assign wire31157 = ( ng174  &  (~ ng826)  &  ng176 ) | ( ng174  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31159 = ( wire3046 ) | ( wire9416 ) | ( wire31156 ) ;
 assign wire31160 = ( wire9421 ) | ( wire9422 ) | ( wire31157 ) ;
 assign wire31162 = ( ng159  &  ng160  &  ng161 ) | ( (~ ng853)  &  ng160  &  ng161 ) ;
 assign wire31164 = ( (~ ng826)  &  ng159  &  ng161 ) | ( (~ ng826)  &  (~ ng853)  &  ng161 ) ;
 assign wire31166 = ( ng159  &  (~ ng823)  &  ng160 ) | ( (~ ng823)  &  (~ ng853)  &  ng160 ) ;
 assign wire31167 = ( (~ ng823)  &  (~ ng853)  &  ng117 ) ;
 assign wire31168 = ( (~ ng826)  &  ng159  &  (~ ng823) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire31171 = ( (~ ng161)  &  ng823 ) ;
 assign wire31172 = ( (~ ng160)  &  ng826 ) ;
 assign wire31178 = ( ng158  &  ng156  &  ng157 ) | ( ng156  &  ng157  &  (~ ng823) ) ;
 assign wire31179 = ( ng158  &  ng156  &  (~ ng826) ) | ( ng156  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31181 = ( wire3046 ) | ( wire9340 ) | ( wire31178 ) ;
 assign wire31182 = ( wire9345 ) | ( wire9346 ) | ( wire31179 ) ;
 assign wire31191 = ( wire3046 ) | ( wire9392 ) | ( wire9393 ) | ( wire9394 ) ;
 assign wire31192 = ( wire9395 ) | ( wire9396 ) | ( wire9397 ) | ( wire9398 ) ;
 assign wire31198 = ( ng172  &  (~ ng853)  &  ng173 ) | ( ng172  &  ng171  &  ng173 ) ;
 assign wire31199 = ( ng172  &  (~ ng823)  &  ng171 ) | ( (~ ng826)  &  (~ ng823)  &  ng171 ) ;
 assign wire31201 = ( wire3046 ) | ( wire9400 ) | ( wire31198 ) ;
 assign wire31202 = ( wire9405 ) | ( wire9406 ) | ( wire31199 ) ;
 assign wire31208 = ( ng164  &  ng162  &  ng163 ) | ( ng162  &  (~ ng823)  &  ng163 ) ;
 assign wire31209 = ( ng164  &  ng162  &  (~ ng826) ) | ( ng162  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31211 = ( wire3046 ) | ( wire9408 ) | ( wire31208 ) ;
 assign wire31212 = ( wire9413 ) | ( wire9414 ) | ( wire31209 ) ;
 assign wire31214 = ( ng826  &  (~ ng151)  &  (~ ng117) ) | ( (~ ng826)  &  ng117  &  wire31145 ) | ( ng151  &  ng117  &  wire31145 ) ;
 assign wire31215 = ( ng117  &  wire3287  &  wire31147 ) | ( ng117  &  wire3287  &  wire31149 ) ;
 assign wire31216 = ( wire9318 ) | ( wire9319 ) | ( wire3287  &  wire31167 ) ;
 assign wire31218 = ( wire31214 ) | ( wire31215 ) | ( wire31216 ) ;
 assign wire31220 = ( (~ wire31159)  &  (~ wire31160)  &  wire31164 ) | ( (~ wire31159)  &  (~ wire31160)  &  wire31166 ) ;
 assign wire31221 = ( wire31159  &  wire31171 ) | ( wire31160  &  wire31171 ) | ( (~ wire31159)  &  (~ wire31160)  &  wire31168 ) ;
 assign wire31222 = ( (~ wire3286)  &  wire31159 ) | ( (~ wire3286)  &  wire31160 ) | ( wire31159  &  wire31172 ) | ( wire31160  &  wire31172 ) ;
 assign wire31223 = ( ng125  &  wire31181 ) | ( ng125  &  wire31182 ) | ( (~ ng125)  &  (~ wire31181)  &  (~ wire31182) ) ;
 assign wire31224 = ( ng121  &  wire31191 ) | ( ng121  &  wire31192 ) | ( (~ ng121)  &  (~ wire31191)  &  (~ wire31192) ) ;
 assign wire31225 = ( (~ wire31201)  &  (~ wire31202)  &  wire31211 ) | ( (~ wire31201)  &  (~ wire31202)  &  wire31212 ) | ( wire31201  &  (~ wire31211)  &  (~ wire31212) ) | ( wire31202  &  (~ wire31211)  &  (~ wire31212) ) ;
 assign wire31226 = ( wire3368 ) | ( wire9313 ) | ( wire31218 ) ;
 assign wire31227 = ( wire31221 ) | ( wire31220 ) ;
 assign wire31231 = ( wire31222 ) | ( wire31223 ) | ( wire31224 ) | ( wire31225 ) ;
 assign wire31232 = ( wire31143 ) | ( wire31144 ) | ( wire31226 ) | ( wire31227 ) ;
 assign wire31233 = ( (~ ng403)  &  ng826 ) ;
 assign wire31234 = ( (~ ng402)  &  ng853 ) ;
 assign wire31235 = ( ng823  &  (~ ng404) ) ;
 assign wire31236 = ( (~ wire31231)  &  (~ wire31232)  &  wire31233 ) | ( (~ wire31231)  &  (~ wire31232)  &  wire31234 ) ;
 assign wire31245 = ( wire3368 ) | ( (~ ng18183)  &  wire3054  &  wire3065 ) ;
 assign wire31248 = ( (~ ng18079)  &  (~ ng18183)  &  (~ ng18346) ) | ( (~ ng18079)  &  (~ ng18183)  &  wire3054 ) | ( (~ ng18079)  &  (~ ng18346)  &  wire3054 ) | ( (~ ng18183)  &  (~ ng18346)  &  wire3054 ) ;
 assign wire31249 = ( wire3065  &  wire3326 ) | ( (~ ng18079)  &  (~ ng18346)  &  wire3326 ) ;
 assign wire31250 = ( wire9293 ) | ( wire9294 ) | ( wire31245 ) ;
 assign wire31251 = ( wire9288 ) | ( wire9295 ) | ( wire31248 ) ;
 assign wire31261 = ( wire3368 ) | ( (~ ng17807)  &  (~ ng17729)  &  wire3106 ) ;
 assign wire31264 = ( (~ ng18419)  &  (~ ng17887)  &  (~ ng17807) ) | ( (~ ng18419)  &  (~ ng17887)  &  (~ ng17729) ) | ( (~ ng18419)  &  (~ ng17807)  &  (~ ng17729) ) | ( (~ ng17887)  &  (~ ng17807)  &  (~ ng17729) ) ;
 assign wire31265 = ( wire3106  &  wire3284 ) | ( (~ ng18419)  &  (~ ng17887)  &  wire3284 ) ;
 assign wire31266 = ( wire9271 ) | ( wire9272 ) | ( wire31261 ) ;
 assign wire31267 = ( wire9266 ) | ( wire9273 ) | ( wire31264 ) ;
 assign wire31269 = ( wire30957  &  (~ wire30967)  &  (~ wire30968) ) | ( wire30958  &  (~ wire30967)  &  (~ wire30968) ) ;
 assign wire31270 = ( (~ wire31231)  &  (~ wire31232)  &  wire31269 ) ;
 assign wire31271 = ( (~ wire30957)  &  (~ wire30958)  &  (~ wire30967)  &  (~ wire30968) ) ;
 assign wire31272 = ( (~ ng322)  &  ng826 ) | ( ng853  &  (~ ng321) ) ;
 assign wire31273 = ( wire9260  &  wire30977 ) | ( wire9260  &  wire30978 ) | ( wire30977  &  wire31272 ) | ( wire30978  &  wire31272 ) ;
 assign wire31274 = ( wire9263 ) | ( wire31236 ) | ( (~ ng13378)  &  wire3936 ) ;
 assign wire31279 = ( (~ wire30927)  &  (~ wire30928)  &  wire31028 ) | ( (~ wire30927)  &  (~ wire30928)  &  wire31029 ) | ( wire30927  &  (~ wire31028)  &  (~ wire31029) ) | ( wire30928  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire31281 = ( (~ ng12967)  &  ng12849 ) | ( ng11624  &  (~ ng12849) ) | ( (~ ng12849)  &  (~ wire30979) ) | ( (~ ng11624)  &  ng12967  &  wire30979 ) ;
 assign wire31283 = ( (~ ng12698)  &  ng12880 ) | ( ng11624  &  (~ ng12880) ) | ( (~ ng12880)  &  (~ wire30979) ) | ( (~ ng11624)  &  ng12698  &  wire30979 ) ;
 assign wire31284 = ( (~ ng12698)  &  (~ wire30977)  &  (~ wire30978)  &  wire30979 ) ;
 assign wire31285 = ( ng27563  &  (~ wire31279)  &  (~ wire31281)  &  wire31284 ) ;
 assign wire31287 = ( (~ ng12880)  &  (~ wire30977)  &  (~ wire30978)  &  wire30979 ) ;
 assign wire31289 = ( (~ wire30947)  &  (~ wire30948)  &  (~ wire31008)  &  (~ wire31009) ) ;
 assign wire31292 = ( (~ ng28501)  &  ng26892  &  wire31285 ) | ( (~ ng28501)  &  ng26892  &  wire31287 ) ;
 assign wire31293 = ( (~ ng28501)  &  (~ ng16643)  &  (~ ng26892) ) | ( (~ ng28501)  &  ng26892  &  wire31289 ) ;
 assign wire31297 = ( (~ ng2903)  &  (~ ng2892) ) ;
 assign wire31298 = ( (~ ng2900)  &  (~ ng2896)  &  (~ ng2908) ) ;
 assign wire31311 = ( ng373  &  ng376  &  ng384 ) | ( ng373  &  ng376  &  (~ ng826) ) ;
 assign wire31312 = ( ng376  &  ng384  &  (~ ng823) ) | ( ng376  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31314 = ( wire3046 ) | ( wire9210 ) | ( wire31311 ) ;
 assign wire31315 = ( wire9215 ) | ( wire9216 ) | ( wire31312 ) ;
 assign wire31321 = ( ng343  &  ng346  &  ng354 ) | ( ng343  &  ng346  &  (~ ng826) ) ;
 assign wire31322 = ( ng346  &  ng354  &  (~ ng823) ) | ( ng346  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31324 = ( wire3046 ) | ( wire9202 ) | ( wire31321 ) ;
 assign wire31325 = ( wire9207 ) | ( wire9208 ) | ( wire31322 ) ;
 assign wire31331 = ( ng369  &  ng358  &  ng361 ) | ( ng369  &  ng361  &  (~ ng823) ) ;
 assign wire31334 = ( wire3046 ) | ( wire9218 ) | ( wire31331 ) ;
 assign wire31335 = ( wire9221 ) | ( wire9222 ) | ( wire9223 ) | ( wire9224 ) ;
 assign wire31336 = ( (~ wire30957)  &  (~ wire30958)  &  wire30967 ) | ( (~ wire30957)  &  (~ wire30958)  &  wire30968 ) ;
 assign wire31345 = ( wire3046 ) | ( wire9186 ) | ( wire9187 ) | ( wire9188 ) ;
 assign wire31346 = ( wire9189 ) | ( wire9190 ) | ( wire9191 ) | ( wire9192 ) ;
 assign wire31353 = ( (~ ng826)  &  (~ ng823)  &  (~ ng423) ) | ( (~ ng826)  &  (~ ng423)  &  (~ ng420) ) ;
 assign wire31355 = ( wire3046 ) | ( wire9178 ) | ( wire9179 ) | ( wire9180 ) ;
 assign wire31356 = ( wire9183 ) | ( wire9184 ) | ( wire31353 ) ;
 assign wire31360 = ( ng113  &  ng117  &  ng97  &  ng125 ) ;
 assign wire31361 = ( ng121  &  ng101  &  ng105  &  ng109 ) ;
 assign wire31362 = ( wire31159 ) | ( wire31160 ) | ( (~ wire31360) ) | ( (~ wire31361) ) ;
 assign wire31365 = ( ng2257  &  wire31355 ) | ( ng2257  &  wire31356 ) ;
 assign wire31368 = ( ng427  &  ng428  &  (~ ng853) ) ;
 assign wire31370 = ( ng428  &  (~ ng826)  &  ng426 ) ;
 assign wire31372 = ( ng427  &  ng428  &  ng426 ) ;
 assign wire31374 = ( ng427  &  ng426  &  (~ ng823) ) ;
 assign wire31375 = ( (~ ng826)  &  ng426  &  (~ ng823) ) ;
 assign wire31376 = ( ng427  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire31377 = ( ng428  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire31382 = ( wire9167 ) | ( wire9168 ) | ( wire9169 ) | ( wire9170 ) ;
 assign wire31383 = ( wire9171 ) | ( wire9172 ) | ( wire9173 ) | ( wire9174 ) ;
 assign wire31391 = ( (~ ng441)  &  (~ ng444)  &  (~ ng438) ) | ( (~ ng444)  &  (~ ng823)  &  (~ ng438) ) ;
 assign wire31392 = ( (~ ng441)  &  (~ ng444)  &  (~ ng826) ) | ( (~ ng444)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31394 = ( wire3046 ) | ( wire9134 ) | ( wire31391 ) ;
 assign wire31395 = ( wire9139 ) | ( wire9140 ) | ( wire31392 ) ;
 assign wire31404 = ( wire3046 ) | ( wire9142 ) | ( wire9143 ) | ( wire9144 ) ;
 assign wire31405 = ( wire9145 ) | ( wire9146 ) | ( wire9147 ) | ( wire9148 ) ;
 assign wire31411 = ( ng178  &  ng179  &  ng177 ) | ( ng178  &  (~ ng823)  &  ng177 ) ;
 assign wire31414 = ( wire3046 ) | ( wire9150 ) | ( (~ wire31360) ) | ( (~ wire31361) ) ;
 assign wire31415 = ( wire9153 ) | ( wire9154 ) | ( wire31411 ) ;
 assign wire31418 = ( (~ ng449)  &  ng823  &  ng2257 ) ;
 assign wire31419 = ( (~ ng447)  &  ng853  &  ng2257 ) ;
 assign wire31420 = ( (~ ng448)  &  ng826  &  ng2257 ) ;
 assign wire31426 = ( (~ ng101)  &  (~ ng17729)  &  wire31018 ) | ( (~ ng101)  &  (~ ng17729)  &  wire31019 ) | ( ng101  &  (~ ng17729)  &  (~ wire31018)  &  (~ wire31019) ) ;
 assign wire31427 = ( (~ ng18079)  &  (~ ng18183)  &  (~ ng18346)  &  wire3054 ) ;
 assign wire31428 = ( wire3065  &  (~ ng18419)  &  (~ ng17887)  &  (~ ng17807) ) ;
 assign wire31431 = ( (~ ng13378)  &  (~ ng11624)  &  wire30957 ) | ( (~ ng13378)  &  (~ ng11624)  &  wire30958 ) ;
 assign wire31432 = ( ng23495  &  (~ wire30957)  &  (~ wire30958) ) ;
 assign wire31436 = ( (~ ng11644)  &  ng13378 ) | ( (~ ng2257)  &  ng11644  &  (~ ng13378) ) | ( (~ ng11644)  &  (~ ng13378)  &  ng11624 ) ;
 assign wire31437 = ( wire31436 ) | ( (~ ng23495)  &  wire31431 ) ;
 assign wire31438 = ( wire31437 ) | ( ng23486  &  ng23478  &  wire31432 ) ;
 assign wire31449 = ( wire3049 ) | ( wire9100 ) | ( wire9101 ) | ( wire9102 ) ;
 assign wire31450 = ( wire9103 ) | ( wire9104 ) | ( wire9105 ) | ( wire9106 ) ;
 assign wire31456 = ( (~ ng490)  &  (~ ng1315)  &  (~ ng493) ) | ( (~ ng490)  &  (~ ng493)  &  (~ ng496) ) ;
 assign wire31457 = ( (~ ng490)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng490)  &  (~ ng1312)  &  (~ ng496) ) ;
 assign wire31459 = ( wire3049 ) | ( wire9092 ) | ( wire31456 ) ;
 assign wire31460 = ( wire9097 ) | ( wire9098 ) | ( wire31457 ) ;
 assign wire31469 = ( wire3049 ) | ( wire9084 ) | ( wire9085 ) | ( wire9086 ) ;
 assign wire31470 = ( wire9087 ) | ( wire9088 ) | ( wire9089 ) | ( wire9090 ) ;
 assign wire31471 = ( (~ ng3002)  &  (~ ng3013) ) ;
 assign wire31472 = ( (~ ng3006)  &  (~ ng3024)  &  (~ ng3010) ) ;
 assign wire31479 = ( ng584  &  (~ ng1309)  &  ng586 ) | ( ng584  &  ng585  &  ng586 ) ;
 assign wire31480 = ( ng584  &  (~ ng1312)  &  ng585 ) | ( (~ ng1312)  &  (~ ng1315)  &  ng585 ) ;
 assign wire31482 = ( wire3049 ) | ( wire9065 ) | ( wire31479 ) ;
 assign wire31483 = ( wire9070 ) | ( wire9071 ) | ( wire31480 ) ;
 assign wire31489 = ( ng575  &  ng577  &  ng576 ) | ( ng575  &  (~ ng1312)  &  ng576 ) ;
 assign wire31492 = ( wire3049 ) | ( wire9057 ) | ( wire31489 ) ;
 assign wire31493 = ( wire9060 ) | ( wire9061 ) | ( wire9062 ) | ( wire9063 ) ;
 assign wire31500 = ( (~ ng1312)  &  (~ ng1315)  &  ng582 ) | ( (~ ng1315)  &  ng582  &  ng583 ) ;
 assign wire31502 = ( wire3049 ) | ( wire9073 ) | ( wire9074 ) | ( wire9075 ) ;
 assign wire31503 = ( wire9078 ) | ( wire9079 ) | ( wire31500 ) ;
 assign wire31509 = ( ng580  &  ng579  &  ng578 ) | ( (~ ng1312)  &  ng579  &  ng578 ) ;
 assign wire31510 = ( ng580  &  (~ ng1315)  &  ng579 ) | ( (~ ng1312)  &  (~ ng1315)  &  ng579 ) ;
 assign wire31512 = ( wire3049 ) | ( wire9049 ) | ( wire31509 ) ;
 assign wire31513 = ( wire9054 ) | ( wire9055 ) | ( wire31510 ) ;
 assign wire31514 = ( wire31482  &  (~ wire31492)  &  (~ wire31493) ) | ( wire31483  &  (~ wire31492)  &  (~ wire31493) ) ;
 assign wire31518 = ( pg3229  &  (~ ng12145)  &  (~ ng12033) ) | ( (~ pg3229)  &  ng12145  &  (~ ng12080) ) ;
 assign wire31522 = ( ng3018  &  (~ ng2993)  &  (~ ng3036) ) ;
 assign wire31523 = ( ng3013  &  ng3002  &  (~ ng3006)  &  (~ ng3010) ) ;
 assign wire31524 = ( ng2998  &  ng3028  &  ng3024  &  (~ ng3032) ) ;
 assign wire31550 = ( wire3049 ) | ( wire9031 ) | ( wire9032 ) | ( wire9033 ) ;
 assign wire31551 = ( wire9034 ) | ( wire9035 ) | ( wire9036 ) | ( wire9037 ) ;
 assign wire31553 = ( (~ ng590)  &  (~ ng593)  &  (~ ng1309) ) ;
 assign wire31555 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng587) ) ;
 assign wire31557 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng587) ) ;
 assign wire31559 = ( (~ ng590)  &  (~ ng593)  &  (~ ng587) ) ;
 assign wire31562 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng587) ) ;
 assign wire31565 = ( (~ ng593)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire31568 = ( (~ ng590)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire31577 = ( wire9007 ) | ( wire9008 ) | ( wire9009 ) | ( wire9010 ) ;
 assign wire31578 = ( wire9011 ) | ( wire9012 ) | ( wire9013 ) | ( wire9014 ) ;
 assign wire31579 = ( wire9019 ) | ( wire9020 ) | ( wire9022 ) | ( wire9023 ) ;
 assign wire31580 = ( wire9025 ) | ( wire9026 ) | ( wire9028 ) | ( wire9029 ) ;
 assign wire31582 = ( wire31580 ) | ( wire31579 ) ;
 assign wire31584 = ( wire31550  &  wire31555 ) | ( wire31551  &  wire31555 ) | ( wire31550  &  wire31557 ) | ( wire31551  &  wire31557 ) ;
 assign wire31585 = ( wire31550  &  wire31559 ) | ( wire31551  &  wire31559 ) | ( wire31550  &  wire31562 ) | ( wire31551  &  wire31562 ) ;
 assign wire31586 = ( wire31550  &  wire31565 ) | ( wire31551  &  wire31565 ) | ( wire31550  &  wire31568 ) | ( wire31551  &  wire31568 ) ;
 assign wire31587 = ( wire9030 ) | ( wire31579 ) | ( wire31580 ) ;
 assign wire31588 = ( wire9015 ) | ( wire31577 ) | ( wire31578 ) | ( wire31584 ) ;
 assign wire31589 = ( wire31586 ) | ( wire31585 ) ;
 assign wire31591 = ( ng640  &  ng633 ) ;
 assign wire31592 = ( ng1315  &  (~ ng659)  &  ng653 ) ;
 assign wire31602 = ( ng712  &  (~ ng1315)  &  ng711 ) | ( ng712  &  ng710  &  ng711 ) ;
 assign wire31605 = ( wire3049 ) | ( wire8915 ) | ( wire31602 ) ;
 assign wire31606 = ( wire8918 ) | ( wire8919 ) | ( wire8920 ) | ( wire8921 ) ;
 assign wire31613 = ( (~ ng1312)  &  (~ ng1315)  &  ng732 ) | ( (~ ng1315)  &  ng732  &  ng733 ) ;
 assign wire31615 = ( wire3049 ) | ( wire8907 ) | ( wire8908 ) | ( wire8909 ) ;
 assign wire31616 = ( wire8912 ) | ( wire8913 ) | ( wire31613 ) ;
 assign wire31627 = ( wire3049 ) | ( wire8923 ) | ( wire8924 ) | ( wire8925 ) ;
 assign wire31628 = ( wire8926 ) | ( wire8927 ) | ( wire8928 ) | ( wire8929 ) ;
 assign wire31639 = ( wire3049 ) | ( wire8931 ) | ( wire8932 ) | ( wire8933 ) ;
 assign wire31640 = ( wire8934 ) | ( wire8935 ) | ( wire8936 ) | ( wire8937 ) ;
 assign wire31651 = ( wire3049 ) | ( wire8939 ) | ( wire8940 ) | ( wire8941 ) ;
 assign wire31652 = ( wire8942 ) | ( wire8943 ) | ( wire8944 ) | ( wire8945 ) ;
 assign wire31663 = ( wire3049 ) | ( wire8955 ) | ( wire8956 ) | ( wire8957 ) ;
 assign wire31664 = ( wire8958 ) | ( wire8959 ) | ( wire8960 ) | ( wire8961 ) ;
 assign wire31672 = ( ng703  &  ng702  &  ng701 ) | ( ng702  &  (~ ng1312)  &  ng701 ) ;
 assign wire31673 = ( ng703  &  ng702  &  (~ ng1315) ) | ( ng702  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire31675 = ( wire3049 ) | ( wire8947 ) | ( wire31672 ) ;
 assign wire31676 = ( wire8952 ) | ( wire8953 ) | ( wire31673 ) ;
 assign wire31684 = ( ng705  &  (~ ng1315)  &  ng706 ) | ( ng705  &  ng704  &  ng706 ) ;
 assign wire31685 = ( ng705  &  (~ ng1312)  &  (~ ng1315) ) | ( ng705  &  (~ ng1312)  &  ng704 ) ;
 assign wire31687 = ( wire3049 ) | ( wire8963 ) | ( wire31684 ) ;
 assign wire31688 = ( wire8968 ) | ( wire8969 ) | ( wire31685 ) ;
 assign wire31699 = ( wire3049 ) | ( wire8971 ) | ( wire8972 ) | ( wire8973 ) ;
 assign wire31700 = ( wire8974 ) | ( wire8975 ) | ( wire8976 ) | ( wire8977 ) ;
 assign wire31708 = ( ng714  &  ng715  &  ng713 ) | ( ng714  &  (~ ng1312)  &  ng713 ) ;
 assign wire31709 = ( ng714  &  ng715  &  (~ ng1315) ) | ( ng714  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire31711 = ( wire3049 ) | ( wire8979 ) | ( wire31708 ) ;
 assign wire31712 = ( wire8984 ) | ( wire8985 ) | ( wire31709 ) ;
 assign wire31723 = ( wire3049 ) | ( wire8987 ) | ( wire8988 ) | ( wire8989 ) ;
 assign wire31724 = ( wire8990 ) | ( wire8991 ) | ( wire8992 ) | ( wire8993 ) ;
 assign wire31727 = ( ng660  &  ng12036  &  wire31605 ) | ( ng660  &  ng12036  &  wire31606 ) | ( (~ ng660)  &  ng12036  &  (~ wire31605)  &  (~ wire31606) ) ;
 assign wire31728 = ( ng666  &  ng12036  &  wire31627 ) | ( ng666  &  ng12036  &  wire31628 ) | ( (~ ng666)  &  ng12036  &  (~ wire31627)  &  (~ wire31628) ) ;
 assign wire31729 = ( ng640  &  ng12036  &  wire31639 ) | ( ng640  &  ng12036  &  wire31640 ) | ( (~ ng640)  &  ng12036  &  (~ wire31639)  &  (~ wire31640) ) ;
 assign wire31730 = ( ng646  &  ng12036  &  wire31651 ) | ( ng646  &  ng12036  &  wire31652 ) | ( (~ ng646)  &  ng12036  &  (~ wire31651)  &  (~ wire31652) ) ;
 assign wire31731 = ( ng692  &  ng12036  &  wire31663 ) | ( ng692  &  ng12036  &  wire31664 ) | ( (~ ng692)  &  ng12036  &  (~ wire31663)  &  (~ wire31664) ) ;
 assign wire31732 = ( ng633  &  ng12036  &  wire31675 ) | ( ng633  &  ng12036  &  wire31676 ) | ( (~ ng633)  &  ng12036  &  (~ wire31675)  &  (~ wire31676) ) ;
 assign wire31733 = ( ng653  &  ng12036  &  wire31687 ) | ( ng653  &  ng12036  &  wire31688 ) | ( (~ ng653)  &  ng12036  &  (~ wire31687)  &  (~ wire31688) ) ;
 assign wire31734 = ( ng679  &  ng12036  &  wire31699 ) | ( ng679  &  ng12036  &  wire31700 ) | ( (~ ng679)  &  ng12036  &  (~ wire31699)  &  (~ wire31700) ) ;
 assign wire31735 = ( ng672  &  ng12036  &  wire31711 ) | ( ng672  &  ng12036  &  wire31712 ) | ( (~ ng672)  &  ng12036  &  (~ wire31711)  &  (~ wire31712) ) ;
 assign wire31741 = ( wire31735 ) | ( ng686  &  ng12195  &  ng12036 ) | ( (~ ng686)  &  (~ ng12195)  &  ng12036 ) ;
 assign wire31742 = ( wire31727 ) | ( wire31728 ) | ( wire31729 ) | ( wire31730 ) ;
 assign wire31743 = ( wire31731 ) | ( wire31732 ) | ( wire31733 ) | ( wire31734 ) ;
 assign wire31746 = ( ng730  &  ng728  &  ng729 ) ;
 assign wire31748 = ( (~ ng1312)  &  ng728  &  ng729 ) ;
 assign wire31750 = ( (~ ng1315)  &  ng730  &  ng729 ) ;
 assign wire31752 = ( (~ ng1309)  &  ng730  &  ng728 ) ;
 assign wire31753 = ( (~ ng1312)  &  (~ ng1315)  &  ng729 ) ;
 assign wire31754 = ( (~ ng1312)  &  (~ ng1309)  &  ng728 ) ;
 assign wire31755 = ( (~ ng1315)  &  (~ ng1309)  &  ng730 ) ;
 assign wire31760 = ( wire8879 ) | ( wire8880 ) | ( wire8881 ) | ( wire8882 ) ;
 assign wire31761 = ( wire8883 ) | ( wire8884 ) | ( wire8885 ) | ( wire8886 ) ;
 assign wire31767 = ( ng863  &  ng862  &  ng864 ) | ( ng862  &  (~ ng826)  &  ng864 ) ;
 assign wire31768 = ( ng863  &  ng862  &  (~ ng823) ) | ( ng862  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31770 = ( wire3046 ) | ( wire8865 ) | ( wire31767 ) ;
 assign wire31771 = ( wire8870 ) | ( wire8871 ) | ( wire31768 ) ;
 assign wire31774 = ( (~ ng2920)  &  ng2924 ) ;
 assign wire31775 = ( (~ ng2888)  &  ng2883  &  (~ ng2912)  &  (~ ng2917) ) ;
 assign wire31785 = ( wire3046 ) | ( wire8805 ) | ( wire8806 ) | ( wire8807 ) ;
 assign wire31786 = ( wire8808 ) | ( wire8809 ) | ( wire8810 ) | ( wire8811 ) ;
 assign wire31793 = ( (~ ng826)  &  (~ ng823)  &  ng1007 ) | ( (~ ng826)  &  ng1007  &  ng1006 ) ;
 assign wire31795 = ( wire3046 ) | ( wire8829 ) | ( wire8830 ) | ( wire8831 ) ;
 assign wire31796 = ( wire8834 ) | ( wire8835 ) | ( wire31793 ) ;
 assign wire31805 = ( wire3046 ) | ( wire8845 ) | ( wire8846 ) | ( wire8847 ) ;
 assign wire31806 = ( wire8848 ) | ( wire8849 ) | ( wire8850 ) | ( wire8851 ) ;
 assign wire31812 = ( ng1002  &  ng1003  &  ng1004 ) | ( ng1002  &  (~ ng823)  &  ng1004 ) ;
 assign wire31815 = ( wire3046 ) | ( wire8837 ) | ( wire31812 ) ;
 assign wire31816 = ( wire8840 ) | ( wire8841 ) | ( wire8842 ) | ( wire8843 ) ;
 assign wire31817 = ( wire31795  &  wire31805 ) | ( wire31796  &  wire31805 ) | ( wire31795  &  wire31806 ) | ( wire31796  &  wire31806 ) ;
 assign wire31823 = ( (~ ng876)  &  (~ ng873)  &  (~ ng879) ) | ( (~ ng876)  &  (~ ng879)  &  (~ ng826) ) ;
 assign wire31824 = ( (~ ng873)  &  (~ ng879)  &  (~ ng823) ) | ( (~ ng879)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31826 = ( wire3046 ) | ( wire8797 ) | ( wire31823 ) ;
 assign wire31827 = ( wire8802 ) | ( wire8803 ) | ( wire31824 ) ;
 assign wire31828 = ( wire31795  &  wire31805 ) | ( wire31796  &  wire31805 ) | ( wire31795  &  wire31806 ) | ( wire31796  &  wire31806 ) ;
 assign wire31834 = ( (~ ng882)  &  (~ ng885)  &  (~ ng888) ) | ( (~ ng885)  &  (~ ng888)  &  (~ ng826) ) ;
 assign wire31835 = ( (~ ng882)  &  (~ ng888)  &  (~ ng823) ) | ( (~ ng888)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31837 = ( wire3046 ) | ( wire8757 ) | ( wire31834 ) ;
 assign wire31838 = ( wire8762 ) | ( wire8763 ) | ( wire31835 ) ;
 assign wire31844 = ( (~ ng894)  &  (~ ng897)  &  (~ ng826) ) | ( (~ ng894)  &  (~ ng897)  &  (~ ng891) ) ;
 assign wire31845 = ( (~ ng897)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng897)  &  (~ ng823)  &  (~ ng891) ) ;
 assign wire31847 = ( wire3046 ) | ( wire8853 ) | ( wire31844 ) ;
 assign wire31848 = ( wire8858 ) | ( wire8859 ) | ( wire31845 ) ;
 assign wire31854 = ( (~ ng900)  &  (~ ng906)  &  (~ ng903) ) | ( (~ ng826)  &  (~ ng906)  &  (~ ng903) ) ;
 assign wire31855 = ( (~ ng900)  &  (~ ng823)  &  (~ ng906) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng906) ) ;
 assign wire31857 = ( wire3046 ) | ( wire8781 ) | ( wire31854 ) ;
 assign wire31858 = ( wire8786 ) | ( wire8787 ) | ( wire31855 ) ;
 assign wire31867 = ( wire3046 ) | ( wire8821 ) | ( wire8822 ) | ( wire8823 ) ;
 assign wire31868 = ( wire8824 ) | ( wire8825 ) | ( wire8826 ) | ( wire8827 ) ;
 assign wire31874 = ( (~ ng951)  &  (~ ng826)  &  (~ ng948) ) | ( (~ ng951)  &  (~ ng948)  &  (~ ng945) ) ;
 assign wire31875 = ( (~ ng951)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng951)  &  (~ ng823)  &  (~ ng945) ) ;
 assign wire31877 = ( wire3046 ) | ( wire8813 ) | ( wire31874 ) ;
 assign wire31878 = ( wire8818 ) | ( wire8819 ) | ( wire31875 ) ;
 assign wire31887 = ( wire3046 ) | ( wire8789 ) | ( wire8790 ) | ( wire8791 ) ;
 assign wire31888 = ( wire8792 ) | ( wire8793 ) | ( wire8794 ) | ( wire8795 ) ;
 assign wire31897 = ( wire3046 ) | ( wire8773 ) | ( wire8774 ) | ( wire8775 ) ;
 assign wire31898 = ( wire8776 ) | ( wire8777 ) | ( wire8778 ) | ( wire8779 ) ;
 assign wire31904 = ( (~ ng912)  &  (~ ng915)  &  (~ ng909) ) | ( (~ ng912)  &  (~ ng915)  &  (~ ng826) ) ;
 assign wire31905 = ( (~ ng915)  &  (~ ng909)  &  (~ ng823) ) | ( (~ ng915)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31907 = ( wire3046 ) | ( wire8765 ) | ( wire31904 ) ;
 assign wire31908 = ( wire8770 ) | ( wire8771 ) | ( wire31905 ) ;
 assign wire31909 = ( (~ wire31785)  &  (~ wire31786)  &  (~ wire31837)  &  (~ wire31838) ) ;
 assign wire31910 = ( wire31847  &  wire31857 ) | ( wire31848  &  wire31857 ) | ( wire31847  &  wire31858 ) | ( wire31848  &  wire31858 ) ;
 assign wire31911 = ( (~ wire31867)  &  (~ wire31868)  &  wire31877 ) | ( (~ wire31867)  &  (~ wire31868)  &  wire31878 ) ;
 assign wire31912 = ( wire31887  &  (~ wire31897)  &  (~ wire31898) ) | ( wire31888  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign wire31915 = ( (~ wire31815)  &  (~ wire31816)  &  wire31817  &  wire31912 ) ;
 assign wire31916 = ( (~ ng12789)  &  wire31909  &  wire31910  &  wire31911 ) ;
 assign wire31918 = ( wire31785  &  wire31837 ) | ( wire31786  &  wire31837 ) | ( wire31785  &  wire31838 ) | ( wire31786  &  wire31838 ) ;
 assign wire31919 = ( wire31826  &  wire31847 ) | ( wire31827  &  wire31847 ) | ( wire31826  &  wire31848 ) | ( wire31827  &  wire31848 ) ;
 assign wire31920 = ( wire31857  &  wire31867 ) | ( wire31858  &  wire31867 ) | ( wire31857  &  wire31868 ) | ( wire31858  &  wire31868 ) ;
 assign wire31921 = ( wire31877  &  wire31887 ) | ( wire31878  &  wire31887 ) | ( wire31877  &  wire31888 ) | ( wire31878  &  wire31888 ) ;
 assign wire31922 = ( wire31897  &  wire31907 ) | ( wire31898  &  wire31907 ) | ( wire31897  &  wire31908 ) | ( wire31898  &  wire31908 ) ;
 assign wire31924 = ( wire31921  &  wire31920 ) ;
 assign wire31925 = ( wire31918  &  wire31919  &  wire31922 ) ;
 assign wire31931 = ( ng856  &  (~ ng826)  &  ng858 ) | ( ng856  &  ng857  &  ng858 ) ;
 assign wire31932 = ( ng856  &  (~ ng826)  &  (~ ng823) ) | ( ng856  &  ng857  &  (~ ng823) ) ;
 assign wire31934 = ( wire3046 ) | ( wire8663 ) | ( wire31931 ) ;
 assign wire31935 = ( wire8668 ) | ( wire8669 ) | ( wire31932 ) ;
 assign wire31936 = ( ng833  &  ng832 ) ;
 assign wire31937 = ( (~ ng823)  &  ng797 ) | ( ng834  &  ng797 ) ;
 assign wire31938 = ( ng829  &  ng830 ) ;
 assign wire31939 = ( ng831  &  ng793 ) | ( (~ ng823)  &  ng793 ) ;
 assign wire31963 = ( ng835  &  ng836  &  ng837 ) | ( ng835  &  ng837  &  (~ ng826) ) ;
 assign wire31964 = ( ng835  &  ng836  &  (~ ng823) ) | ( ng835  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31967 = ( wire8734 ) | ( wire8735 ) | ( wire31964 ) ;
 assign wire31973 = ( ng817  &  (~ ng823)  &  ng818 ) | ( ng817  &  ng819  &  ng818 ) ;
 assign wire31974 = ( ng817  &  (~ ng826)  &  (~ ng823) ) | ( ng817  &  (~ ng826)  &  ng819 ) ;
 assign wire31976 = ( wire3046 ) | ( wire8721 ) | ( wire31973 ) ;
 assign wire31977 = ( wire8726 ) | ( wire8727 ) | ( wire31974 ) ;
 assign wire31983 = ( ng821  &  ng820  &  ng822 ) | ( ng820  &  ng822  &  (~ ng826) ) ;
 assign wire31984 = ( ng821  &  ng820  &  (~ ng823) ) | ( ng820  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire31987 = ( wire8718 ) | ( wire8719 ) | ( wire31984 ) ;
 assign wire31996 = ( wire31936  &  wire31937 ) | ( wire31938  &  wire31939 ) ;
 assign wire31997 = ( wire8706 ) | ( wire8705 ) ;
 assign wire31998 = ( wire8689 ) | ( wire8690 ) | ( wire8691 ) | ( wire8692 ) ;
 assign wire31999 = ( wire8693 ) | ( wire8694 ) | ( wire8695 ) | ( wire8696 ) ;
 assign wire32000 = ( wire8697 ) | ( wire8698 ) | ( wire8699 ) | ( wire8700 ) ;
 assign wire32001 = ( wire8701 ) | ( wire8702 ) | ( wire8703 ) | ( wire8704 ) ;
 assign wire32004 = ( wire32001 ) | ( wire32000 ) ;
 assign wire32005 = ( wire31996 ) | ( wire31997 ) | ( wire31998 ) | ( wire31999 ) ;
 assign wire32010 = ( wire8709 ) | ( wire32004 ) | ( ng801  &  ng11784 ) | ( (~ ng801)  &  (~ ng11784) ) ;
 assign wire32011 = ( wire8710 ) | ( wire32005 ) | ( ng789  &  ng11981 ) | ( (~ ng789)  &  (~ ng11981) ) ;
 assign wire32017 = ( ng860  &  ng861  &  ng859 ) | ( ng861  &  ng859  &  (~ ng826) ) ;
 assign wire32018 = ( ng860  &  ng859  &  (~ ng823) ) | ( ng859  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32020 = ( wire3046 ) | ( wire8679 ) | ( wire32017 ) ;
 assign wire32021 = ( wire8684 ) | ( wire8685 ) | ( wire32018 ) ;
 assign wire32023 = ( ng852  &  (~ ng853)  &  ng851 ) | ( (~ ng823)  &  (~ ng853)  &  ng851 ) ;
 assign wire32025 = ( ng852  &  ng850  &  ng851 ) | ( ng850  &  (~ ng823)  &  ng851 ) ;
 assign wire32027 = ( ng852  &  ng850  &  (~ ng826) ) | ( ng850  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32028 = ( ng842  &  ng843 ) ;
 assign wire32030 = ( ng842  &  (~ ng823) ) ;
 assign wire32032 = ( ng843  &  (~ ng826) ) ;
 assign wire32034 = ( ng852  &  (~ ng826)  &  (~ ng853) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire32035 = ( (~ ng826)  &  (~ ng823)  &  ng809 ) ;
 assign wire32038 = ( (~ ng851)  &  ng826 ) ;
 assign wire32039 = ( ng853  &  (~ ng850) ) ;
 assign wire32045 = ( ng839  &  ng840  &  ng838 ) | ( ng840  &  ng838  &  (~ ng826) ) ;
 assign wire32046 = ( ng839  &  ng838  &  (~ ng823) ) | ( ng838  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32048 = ( wire3046 ) | ( wire8671 ) | ( wire32045 ) ;
 assign wire32049 = ( wire8676 ) | ( wire8677 ) | ( wire32046 ) ;
 assign wire32058 = ( wire3046 ) | ( wire8737 ) | ( wire8738 ) | ( wire8739 ) ;
 assign wire32059 = ( wire8740 ) | ( wire8741 ) | ( wire8742 ) | ( wire8743 ) ;
 assign wire32065 = ( ng844  &  ng846  &  ng845 ) | ( ng844  &  (~ ng823)  &  ng845 ) ;
 assign wire32066 = ( ng844  &  ng846  &  (~ ng826) ) | ( ng844  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32068 = ( wire3046 ) | ( wire8745 ) | ( wire32065 ) ;
 assign wire32069 = ( wire8750 ) | ( wire8751 ) | ( wire32066 ) ;
 assign wire32071 = ( ng853  &  (~ ng841)  &  (~ ng809) ) | ( (~ ng853)  &  ng809  &  wire32028 ) | ( ng841  &  ng809  &  wire32028 ) ;
 assign wire32072 = ( ng809  &  wire3315  &  wire32030 ) | ( ng809  &  wire3315  &  wire32032 ) ;
 assign wire32073 = ( wire8649 ) | ( wire8650 ) | ( wire3315  &  wire32035 ) ;
 assign wire32075 = ( wire32071 ) | ( wire32072 ) | ( wire32073 ) ;
 assign wire32077 = ( (~ wire32020)  &  (~ wire32021)  &  wire32025 ) | ( (~ wire32020)  &  (~ wire32021)  &  wire32027 ) ;
 assign wire32078 = ( wire32020  &  wire32038 ) | ( wire32021  &  wire32038 ) | ( (~ wire32020)  &  (~ wire32021)  &  wire32034 ) ;
 assign wire32079 = ( (~ wire3316)  &  wire32020 ) | ( (~ wire3316)  &  wire32021 ) | ( wire32020  &  wire32039 ) | ( wire32021  &  wire32039 ) ;
 assign wire32080 = ( ng805  &  wire32048 ) | ( ng805  &  wire32049 ) | ( (~ ng805)  &  (~ wire32048)  &  (~ wire32049) ) ;
 assign wire32081 = ( (~ wire31770)  &  (~ wire31771)  &  wire32058 ) | ( (~ wire31770)  &  (~ wire31771)  &  wire32059 ) | ( wire31770  &  (~ wire32058)  &  (~ wire32059) ) | ( wire31771  &  (~ wire32058)  &  (~ wire32059) ) ;
 assign wire32082 = ( ng813  &  wire32068 ) | ( ng813  &  wire32069 ) | ( (~ ng813)  &  (~ wire32068)  &  (~ wire32069) ) ;
 assign wire32083 = ( wire3375 ) | ( wire8641 ) | ( wire32075 ) ;
 assign wire32084 = ( wire32078 ) | ( wire32077 ) ;
 assign wire32088 = ( wire32079 ) | ( wire32080 ) | ( wire32081 ) | ( wire32082 ) ;
 assign wire32089 = ( wire32010 ) | ( wire32011 ) | ( wire32083 ) | ( wire32084 ) ;
 assign wire32090 = ( ng853  &  (~ ng1089) ) ;
 assign wire32091 = ( ng826  &  (~ ng1090) ) ;
 assign wire32092 = ( ng823  &  (~ ng1091) ) ;
 assign wire32093 = ( (~ wire32088)  &  (~ wire32089)  &  wire32090 ) | ( (~ wire32088)  &  (~ wire32089)  &  wire32091 ) ;
 assign wire32102 = ( wire3375 ) | ( (~ ng18441)  &  (~ ng18290)  &  wire3067 ) ;
 assign wire32105 = ( (~ ng18363)  &  (~ ng18441)  &  (~ ng18195) ) | ( (~ ng18363)  &  (~ ng18441)  &  (~ ng18290) ) | ( (~ ng18363)  &  (~ ng18195)  &  (~ ng18290) ) | ( (~ ng18441)  &  (~ ng18195)  &  (~ ng18290) ) ;
 assign wire32106 = ( wire3067  &  wire3285 ) | ( (~ ng18363)  &  (~ ng18195)  &  wire3285 ) ;
 assign wire32107 = ( wire8624 ) | ( wire8625 ) | ( wire32102 ) ;
 assign wire32108 = ( wire8619 ) | ( wire8626 ) | ( wire32105 ) ;
 assign wire32118 = ( wire3375 ) | ( (~ ng18492)  &  wire3056  &  wire3107 ) ;
 assign wire32121 = ( (~ ng18096)  &  (~ ng17998)  &  (~ ng18492) ) | ( (~ ng18096)  &  (~ ng17998)  &  wire3056 ) | ( (~ ng18096)  &  (~ ng18492)  &  wire3056 ) | ( (~ ng17998)  &  (~ ng18492)  &  wire3056 ) ;
 assign wire32122 = ( wire3107  &  wire3328 ) | ( (~ ng18096)  &  (~ ng17998)  &  wire3328 ) ;
 assign wire32123 = ( wire8602 ) | ( wire8603 ) | ( wire32118 ) ;
 assign wire32124 = ( wire8597 ) | ( wire8604 ) | ( wire32121 ) ;
 assign wire32126 = ( wire31795  &  (~ wire31805)  &  (~ wire31806) ) | ( wire31796  &  (~ wire31805)  &  (~ wire31806) ) ;
 assign wire32127 = ( (~ wire32088)  &  (~ wire32089)  &  wire32126 ) ;
 assign wire32128 = ( (~ wire31795)  &  (~ wire31796)  &  (~ wire31805)  &  (~ wire31806) ) ;
 assign wire32129 = ( (~ ng1009)  &  ng826 ) | ( (~ ng1008)  &  ng853 ) ;
 assign wire32130 = ( wire8591  &  wire31815 ) | ( wire8591  &  wire31816 ) | ( wire31815  &  wire32129 ) | ( wire31816  &  wire32129 ) ;
 assign wire32131 = ( wire8594 ) | ( wire32093 ) | ( (~ ng11600)  &  wire3930 ) ;
 assign wire32135 = ( (~ ng28529)  &  (~ ng25958)  &  wire31785 ) | ( (~ ng28529)  &  (~ ng25958)  &  wire31786 ) | ( (~ ng28529)  &  ng25958  &  (~ wire31785)  &  (~ wire31786) ) ;
 assign wire32136 = ( ng789  &  ng27743 ) | ( (~ ng16655)  &  ng25818  &  (~ ng27743) ) ;
 assign wire32140 = ( (~ ng12968)  &  ng11647 ) | ( ng12968  &  (~ ng12852) ) | ( (~ ng12968)  &  (~ wire31817) ) | ( (~ ng11647)  &  ng12852  &  wire31817 ) ;
 assign wire32142 = ( (~ ng12991)  &  ng12890 ) | ( ng11647  &  (~ ng12890) ) | ( (~ ng12890)  &  (~ wire31817) ) | ( (~ ng11647)  &  ng12991  &  wire31817 ) ;
 assign wire32144 = ( (~ ng26925)  &  (~ wire31847)  &  (~ wire31848)  &  wire32142 ) ;
 assign wire32145 = ( (~ wire31847)  &  (~ wire31848)  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign wire32146 = ( ng26925  &  wire32145 ) | ( wire32142  &  wire32145 ) ;
 assign wire32147 = ( ng26925  &  (~ wire31887)  &  (~ wire31888) ) | ( (~ wire31887)  &  (~ wire31888)  &  wire32142 ) ;
 assign wire32148 = ( (~ ng26925)  &  wire31887  &  (~ wire32142) ) | ( (~ ng26925)  &  wire31888  &  (~ wire32142) ) ;
 assign wire32149 = ( ng26925  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign wire32150 = ( (~ ng28529)  &  wire32146 ) | ( (~ ng28529)  &  wire32148 ) ;
 assign wire32151 = ( (~ ng28529)  &  wire32149 ) | ( (~ ng28529)  &  ng16655  &  wire32144 ) ;
 assign wire32155 = ( ng11647  &  (~ ng12755) ) | ( ng12755  &  (~ ng12920) ) | ( (~ ng12755)  &  (~ wire31817) ) | ( (~ ng11647)  &  ng12920  &  wire31817 ) ;
 assign wire32156 = ( (~ ng12789)  &  (~ wire31815)  &  (~ wire31816)  &  wire31817 ) ;
 assign wire32157 = ( ng12789  &  wire31815 ) | ( ng12789  &  wire31816 ) | ( ng12789  &  (~ wire31817) ) ;
 assign wire32160 = ( (~ ng28529)  &  ng27482  &  wire31867 ) | ( (~ ng28529)  &  ng27482  &  wire31868 ) | ( (~ ng28529)  &  (~ ng27482)  &  (~ wire31867)  &  (~ wire31868) ) ;
 assign wire32161 = ( ng27743  &  (~ ng11807) ) | ( (~ ng16655)  &  ng25818  &  (~ ng27743) ) ;
 assign wire32164 = ( ng767  &  ng776  &  ng771  &  ng780 ) ;
 assign wire32166 = ( ng749  &  ng753  &  ng758 ) ;
 assign wire32174 = ( ng1048  &  ng1056  &  ng1045 ) | ( ng1048  &  ng1056  &  (~ ng823) ) ;
 assign wire32177 = ( wire3046 ) | ( wire8540 ) | ( wire32174 ) ;
 assign wire32178 = ( wire8543 ) | ( wire8544 ) | ( wire8545 ) | ( wire8546 ) ;
 assign wire32184 = ( ng1041  &  (~ ng853)  &  ng1030 ) | ( ng1041  &  ng1033  &  ng1030 ) ;
 assign wire32185 = ( ng1041  &  (~ ng823)  &  ng1033 ) | ( (~ ng826)  &  (~ ng823)  &  ng1033 ) ;
 assign wire32187 = ( wire3046 ) | ( wire8524 ) | ( wire32184 ) ;
 assign wire32188 = ( wire8529 ) | ( wire8530 ) | ( wire32185 ) ;
 assign wire32197 = ( wire3046 ) | ( wire8532 ) | ( wire8533 ) | ( wire8534 ) ;
 assign wire32198 = ( wire8535 ) | ( wire8536 ) | ( wire8537 ) | ( wire8538 ) ;
 assign wire32199 = ( wire32177  &  wire32197 ) | ( wire32178  &  wire32197 ) | ( wire32177  &  wire32198 ) | ( wire32178  &  wire32198 ) ;
 assign wire32200 = ( (~ wire31795)  &  (~ wire31796)  &  wire31805 ) | ( (~ wire31795)  &  (~ wire31796)  &  wire31806 ) ;
 assign wire32206 = ( (~ ng1095)  &  (~ ng1098)  &  (~ ng1101) ) | ( (~ ng1098)  &  (~ ng1101)  &  (~ ng826) ) ;
 assign wire32207 = ( (~ ng1095)  &  (~ ng1101)  &  (~ ng823) ) | ( (~ ng1101)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32209 = ( wire3046 ) | ( wire8510 ) | ( wire32206 ) ;
 assign wire32210 = ( wire8515 ) | ( wire8516 ) | ( wire32207 ) ;
 assign wire32219 = ( wire3046 ) | ( wire8502 ) | ( wire8503 ) | ( wire8504 ) ;
 assign wire32220 = ( wire8505 ) | ( wire8506 ) | ( wire8507 ) | ( wire8508 ) ;
 assign wire32224 = ( ng809  &  ng789  &  ng801  &  ng813 ) ;
 assign wire32225 = ( ng805  &  ng785  &  ng793  &  ng797 ) ;
 assign wire32226 = ( wire31770 ) | ( wire31771 ) | ( (~ wire32224) ) | ( (~ wire32225) ) ;
 assign wire32229 = ( ng1115  &  (~ ng853)  &  ng1114 ) ;
 assign wire32231 = ( ng1113  &  (~ ng823)  &  ng1114 ) ;
 assign wire32233 = ( ng1113  &  ng1115  &  ng1114 ) ;
 assign wire32235 = ( ng1113  &  ng1115  &  (~ ng826) ) ;
 assign wire32236 = ( ng1113  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32237 = ( (~ ng823)  &  (~ ng853)  &  ng1114 ) ;
 assign wire32238 = ( ng1115  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire32243 = ( wire8491 ) | ( wire8492 ) | ( wire8493 ) | ( wire8494 ) ;
 assign wire32244 = ( wire8495 ) | ( wire8496 ) | ( wire8497 ) | ( wire8498 ) ;
 assign wire32245 = ( (~ ng25082)  &  wire32209 ) | ( (~ ng25082)  &  wire32210 ) ;
 assign wire32246 = ( ng1113  &  (~ ng853) ) | ( ng1113  &  (~ wire32243)  &  (~ wire32244) ) ;
 assign wire32247 = ( (~ ng11600)  &  (~ ng11647) ) | ( (~ ng11600)  &  wire31795 ) | ( (~ ng11600)  &  wire31796 ) ;
 assign wire32248 = ( (~ wire8594)  &  (~ wire32093)  &  wire32247 ) ;
 assign wire32249 = ( ng11600  &  (~ ng11647)  &  wire31795 ) | ( ng11600  &  (~ ng11647)  &  wire31796 ) ;
 assign wire32252 = ( ng823  &  ng986 ) ;
 assign wire32253 = ( (~ ng986)  &  (~ ng985) ) | ( ng992  &  ng986  &  (~ ng823) ) ;
 assign wire32259 = ( (~ ng1125)  &  (~ ng1128)  &  (~ ng1131) ) | ( (~ ng826)  &  (~ ng1128)  &  (~ ng1131) ) ;
 assign wire32260 = ( (~ ng1125)  &  (~ ng823)  &  (~ ng1131) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng1131) ) ;
 assign wire32262 = ( wire3046 ) | ( wire8469 ) | ( wire32259 ) ;
 assign wire32263 = ( wire8474 ) | ( wire8475 ) | ( wire32260 ) ;
 assign wire32269 = ( (~ ng1303)  &  (~ ng1306)  &  (~ ng1300) ) | ( (~ ng1306)  &  (~ ng1312)  &  (~ ng1300) ) ;
 assign wire32272 = ( wire3049 ) | ( wire8457 ) | ( wire32269 ) ;
 assign wire32273 = ( wire8460 ) | ( wire8461 ) | ( wire8462 ) | ( wire8463 ) ;
 assign wire32282 = ( wire3049 ) | ( wire8449 ) | ( wire8450 ) | ( wire8451 ) ;
 assign wire32283 = ( wire8452 ) | ( wire8453 ) | ( wire8454 ) | ( wire8455 ) ;
 assign wire32289 = ( (~ ng1291)  &  (~ ng1312)  &  (~ ng1297) ) | ( (~ ng1291)  &  (~ ng1294)  &  (~ ng1297) ) ;
 assign wire32290 = ( (~ ng1291)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng1291)  &  (~ ng1315)  &  (~ ng1294) ) ;
 assign wire32292 = ( wire3049 ) | ( wire8441 ) | ( wire32289 ) ;
 assign wire32293 = ( wire8446 ) | ( wire8447 ) | ( wire32290 ) ;
 assign wire32303 = ( wire3049 ) | ( wire8430 ) | ( wire8431 ) | ( wire8432 ) ;
 assign wire32304 = ( wire8433 ) | ( wire8434 ) | ( wire8435 ) | ( wire8436 ) ;
 assign wire32313 = ( wire3049 ) | ( wire8422 ) | ( wire8423 ) | ( wire8424 ) ;
 assign wire32314 = ( wire8425 ) | ( wire8426 ) | ( wire8427 ) | ( wire8428 ) ;
 assign wire32321 = ( (~ ng1312)  &  (~ ng1315)  &  ng1262 ) | ( (~ ng1315)  &  ng1263  &  ng1262 ) ;
 assign wire32323 = ( wire3049 ) | ( wire8414 ) | ( wire8415 ) | ( wire8416 ) ;
 assign wire32324 = ( wire8419 ) | ( wire8420 ) | ( wire32321 ) ;
 assign wire32332 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1251) ) | ( (~ ng1315)  &  (~ ng1251)  &  (~ ng1253) ) ;
 assign wire32334 = ( wire3049 ) | ( wire8400 ) | ( wire8401 ) | ( wire8402 ) ;
 assign wire32335 = ( wire8405 ) | ( wire8406 ) | ( wire32332 ) ;
 assign wire32337 = ( (~ ng1315)  &  (~ ng1282)  &  (~ ng1285) ) ;
 assign wire32339 = ( (~ ng1282)  &  (~ ng1285)  &  (~ ng1288) ) ;
 assign wire32341 = ( (~ ng1309)  &  (~ ng1285)  &  (~ ng1288) ) ;
 assign wire32343 = ( (~ ng1312)  &  (~ ng1282)  &  (~ ng1288) ) ;
 assign wire32360 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1282) ) ;
 assign wire32363 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1288) ) ;
 assign wire32366 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1285) ) ;
 assign wire32377 = ( wire8380 ) | ( wire8381 ) | ( wire8382 ) | ( wire8383 ) ;
 assign wire32378 = ( wire8384 ) | ( wire8385 ) | ( wire8386 ) | ( wire8387 ) ;
 assign wire32379 = ( wire8389 ) | ( wire8390 ) | ( wire8392 ) | ( wire8393 ) ;
 assign wire32380 = ( wire8395 ) | ( wire8396 ) | ( wire8398 ) | ( wire8399 ) ;
 assign wire32384 = ( wire32334  &  wire32339 ) | ( wire32335  &  wire32339 ) | ( wire32334  &  wire32341 ) | ( wire32335  &  wire32341 ) ;
 assign wire32385 = ( wire32334  &  wire32343 ) | ( wire32335  &  wire32343 ) | ( wire32334  &  wire32360 ) | ( wire32335  &  wire32360 ) ;
 assign wire32386 = ( wire32334  &  wire32363 ) | ( wire32335  &  wire32363 ) | ( wire32334  &  wire32366 ) | ( wire32335  &  wire32366 ) ;
 assign wire32387 = ( wire8397 ) | ( wire32379 ) | ( wire32380 ) ;
 assign wire32388 = ( wire8376 ) | ( wire32377 ) | ( wire32378 ) | ( wire32384 ) ;
 assign wire32389 = ( wire32386 ) | ( wire32385 ) ;
 assign wire32396 = ( (~ ng1315)  &  (~ ng1036)  &  (~ ng1038) ) | ( (~ ng1036)  &  (~ ng1038)  &  (~ ng1040) ) ;
 assign wire32397 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1036) ) | ( (~ ng1312)  &  (~ ng1036)  &  (~ ng1040) ) ;
 assign wire32399 = ( wire3049 ) | ( wire8368 ) | ( wire32396 ) ;
 assign wire32400 = ( wire8373 ) | ( wire8374 ) | ( wire32397 ) ;
 assign wire32407 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1066) ) | ( (~ ng1312)  &  (~ ng1070)  &  (~ ng1066) ) ;
 assign wire32409 = ( wire3049 ) | ( wire8360 ) | ( wire8361 ) | ( wire8362 ) ;
 assign wire32410 = ( wire8365 ) | ( wire8366 ) | ( wire32407 ) ;
 assign wire32416 = ( (~ ng1053)  &  (~ ng1055)  &  (~ ng1051) ) | ( (~ ng1055)  &  (~ ng1312)  &  (~ ng1051) ) ;
 assign wire32419 = ( wire3049 ) | ( wire8344 ) | ( wire32416 ) ;
 assign wire32420 = ( wire8347 ) | ( wire8348 ) | ( wire8349 ) | ( wire8350 ) ;
 assign wire32429 = ( wire3049 ) | ( wire8336 ) | ( wire8337 ) | ( wire8338 ) ;
 assign wire32430 = ( wire8339 ) | ( wire8340 ) | ( wire8341 ) | ( wire8342 ) ;
 assign wire32431 = ( wire32303  &  wire32399 ) | ( wire32304  &  wire32399 ) | ( wire32303  &  wire32400 ) | ( wire32304  &  wire32400 ) ;
 assign wire32432 = ( (~ wire32323)  &  (~ wire32324)  &  (~ wire32409)  &  (~ wire32410) ) ;
 assign wire32434 = ( wire8334  &  wire32432 ) | ( wire8335  &  wire32432 ) ;
 assign wire32440 = ( (~ ng1083)  &  (~ ng1081)  &  (~ ng1011) ) | ( (~ ng1312)  &  (~ ng1081)  &  (~ ng1011) ) ;
 assign wire32441 = ( (~ ng1083)  &  (~ ng1315)  &  (~ ng1081) ) | ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1081) ) ;
 assign wire32443 = ( wire3049 ) | ( wire8352 ) | ( wire32440 ) ;
 assign wire32444 = ( wire8357 ) | ( wire8358 ) | ( wire32441 ) ;
 assign wire32445 = ( (~ wire32323)  &  (~ wire32324)  &  wire32399 ) | ( (~ wire32323)  &  (~ wire32324)  &  wire32400 ) ;
 assign wire32446 = ( (~ wire32419)  &  (~ wire32420)  &  (~ wire32443)  &  (~ wire32444) ) ;
 assign wire32448 = ( wire32323  &  (~ wire32443)  &  (~ wire32444) ) | ( wire32324  &  (~ wire32443)  &  (~ wire32444) ) ;
 assign wire32449 = ( wire32313  &  (~ wire32419)  &  (~ wire32420) ) | ( wire32314  &  (~ wire32419)  &  (~ wire32420) ) ;
 assign wire32451 = ( wire32303  &  (~ wire32399)  &  (~ wire32400) ) | ( wire32304  &  (~ wire32399)  &  (~ wire32400) ) ;
 assign wire32452 = ( wire32323  &  wire32409 ) | ( wire32324  &  wire32409 ) | ( wire32323  &  wire32410 ) | ( wire32324  &  wire32410 ) ;
 assign wire32456 = ( (~ wire32323)  &  (~ wire32324)  &  wire32399 ) | ( (~ wire32323)  &  (~ wire32324)  &  wire32400 ) ;
 assign wire32458 = ( (~ wire32303)  &  (~ wire32304)  &  (~ wire32399)  &  (~ wire32400) ) ;
 assign wire32459 = ( (~ wire32409)  &  (~ wire32410)  &  (~ wire32419)  &  (~ wire32420) ) ;
 assign wire32460 = ( wire32323  &  (~ wire32409)  &  (~ wire32410) ) | ( wire32324  &  (~ wire32409)  &  (~ wire32410) ) ;
 assign wire32461 = ( (~ wire32313)  &  (~ wire32314)  &  wire32419 ) | ( (~ wire32313)  &  (~ wire32314)  &  wire32420 ) ;
 assign wire32462 = ( (~ wire32323)  &  (~ wire32324)  &  wire32443 ) | ( (~ wire32323)  &  (~ wire32324)  &  wire32444 ) ;
 assign wire32463 = ( wire32313  &  wire32429 ) | ( wire32314  &  wire32429 ) | ( wire32313  &  wire32430 ) | ( wire32314  &  wire32430 ) ;
 assign wire32464 = ( wire32323  &  (~ wire32399)  &  (~ wire32400) ) | ( wire32324  &  (~ wire32399)  &  (~ wire32400) ) ;
 assign wire32465 = ( wire32458  &  wire32459 ) | ( wire32460  &  wire32461 ) ;
 assign wire32466 = ( wire32462  &  wire32463 ) | ( (~ wire3288)  &  wire32464 ) ;
 assign wire32469 = ( wire32465 ) | ( wire8318 ) ;
 assign wire32470 = ( wire32466 ) | ( (~ ng10801)  &  wire32431  &  wire32434 ) ;
 assign wire32471 = ( wire8314 ) | ( wire8315 ) | ( wire8316 ) | ( wire8317 ) ;
 assign wire32486 = ( (~ ng1255)  &  (~ ng1315)  &  (~ ng1257) ) | ( (~ ng1255)  &  (~ ng1259)  &  (~ ng1257) ) ;
 assign wire32487 = ( (~ ng1255)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng1255)  &  (~ ng1312)  &  (~ ng1259) ) ;
 assign wire32489 = ( wire3049 ) | ( wire8305 ) | ( wire32486 ) ;
 assign wire32490 = ( wire8310 ) | ( wire8311 ) | ( wire32487 ) ;
 assign wire32492 = ( (~ ng1273)  &  (~ ng1276)  &  (~ ng1279) ) ;
 assign wire32494 = ( (~ ng1312)  &  (~ ng1273)  &  (~ ng1279) ) ;
 assign wire32500 = ( (~ ng1309)  &  (~ ng1276)  &  (~ ng1279) ) ;
 assign wire32504 = ( (~ ng1315)  &  (~ ng1273)  &  (~ ng1276) ) ;
 assign wire32508 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1273) ) ;
 assign wire32511 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1279) ) ;
 assign wire32514 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng1276) ) ;
 assign wire32524 = ( wire8281 ) | ( wire8282 ) | ( wire8283 ) | ( wire8284 ) ;
 assign wire32525 = ( wire8287 ) | ( wire8288 ) | ( wire8290 ) | ( wire8292 ) ;
 assign wire32526 = ( wire8293 ) | ( wire8295 ) | ( wire8296 ) | ( wire8298 ) ;
 assign wire32527 = ( wire8299 ) | ( wire8301 ) | ( wire8302 ) | ( wire8304 ) ;
 assign wire32529 = ( wire32527 ) | ( wire32526 ) ;
 assign wire32531 = ( wire32489  &  wire32494 ) | ( wire32490  &  wire32494 ) | ( wire32489  &  wire32500 ) | ( wire32490  &  wire32500 ) ;
 assign wire32532 = ( wire32489  &  wire32504 ) | ( wire32490  &  wire32504 ) | ( wire32489  &  wire32508 ) | ( wire32490  &  wire32508 ) ;
 assign wire32533 = ( wire32489  &  wire32511 ) | ( wire32490  &  wire32511 ) | ( wire32489  &  wire32514 ) | ( wire32490  &  wire32514 ) ;
 assign wire32534 = ( wire3049 ) | ( wire32526 ) | ( wire32527 ) ;
 assign wire32535 = ( wire8285 ) | ( wire32524 ) | ( wire32525 ) | ( wire32531 ) ;
 assign wire32536 = ( wire32533 ) | ( wire32532 ) ;
 assign wire32538 = ( ng13055  &  (~ wire32387)  &  (~ wire32388)  &  (~ wire32389) ) ;
 assign wire32539 = ( wire32534  &  wire32538 ) | ( wire32535  &  wire32538 ) | ( wire32536  &  wire32538 ) ;
 assign wire32540 = ( (~ wire32399)  &  (~ wire32400)  &  (~ wire32443)  &  (~ wire32444) ) ;
 assign wire32541 = ( (~ wire32313)  &  (~ wire32314)  &  (~ wire32419)  &  (~ wire32420) ) ;
 assign wire32543 = ( (~ wire32399)  &  (~ wire32400)  &  wire32409 ) | ( (~ wire32399)  &  (~ wire32400)  &  wire32410 ) ;
 assign wire32545 = ( wire32409  &  (~ wire32419)  &  (~ wire32420) ) | ( wire32410  &  (~ wire32419)  &  (~ wire32420) ) ;
 assign wire32546 = ( wire8334  &  wire32545 ) | ( wire8335  &  wire32545 ) ;
 assign wire32547 = ( (~ wire32323)  &  (~ wire32324)  &  (~ wire32409)  &  (~ wire32410) ) ;
 assign wire32549 = ( wire32323  &  (~ wire32409)  &  (~ wire32410) ) | ( wire32324  &  (~ wire32409)  &  (~ wire32410) ) ;
 assign wire32552 = ( (~ wire32323)  &  (~ wire32324)  &  (~ wire32443)  &  (~ wire32444) ) ;
 assign wire32553 = ( wire32323  &  wire32443 ) | ( wire32324  &  wire32443 ) | ( wire32323  &  wire32444 ) | ( wire32324  &  wire32444 ) ;
 assign wire32554 = ( (~ wire32323)  &  (~ wire32324)  &  wire32419 ) | ( (~ wire32323)  &  (~ wire32324)  &  wire32420 ) ;
 assign wire32556 = ( ng10793  &  (~ ng12248)  &  ng10814 ) | ( ng10793  &  (~ ng12248)  &  wire32552 ) ;
 assign wire32559 = ( wire8329 ) | ( wire8334  &  wire32554 ) | ( wire8335  &  wire32554 ) ;
 assign wire32560 = ( wire32556 ) | ( ng12207  &  (~ wire8332)  &  wire32546 ) ;
 assign wire32561 = ( wire8323 ) | ( wire8324 ) | ( wire8326 ) | ( wire8327 ) ;
 assign wire32563 = ( ng13055  &  wire32387 ) | ( ng13055  &  wire32388 ) | ( ng13055  &  wire32389 ) ;
 assign wire32564 = ( wire32559  &  wire32563 ) | ( wire32560  &  wire32563 ) | ( wire32561  &  wire32563 ) ;
 assign wire32566 = ( ng1319  &  ng1339 ) ;
 assign wire32567 = ( ng1315  &  (~ ng1345)  &  ng1326 ) ;
 assign wire32568 = ( (~ ng1312)  &  (~ ng1346) ) | ( (~ ng1346)  &  (~ ng1316) ) ;
 assign wire32569 = ( (~ ng1312)  &  ng1346 ) | ( ng1346  &  (~ ng1316) ) ;
 assign wire32575 = ( ng1352  &  ng1358  &  ng1346 ) ;
 assign wire32576 = ( (~ ng1312)  &  ng1358 ) | ( ng1358  &  (~ ng1316) ) ;
 assign wire32578 = ( ng1352  &  (~ ng1312) ) | ( ng1352  &  (~ ng1316) ) ;
 assign wire32587 = ( (~ ng1654)  &  (~ ng1651)  &  (~ ng1648) ) | ( (~ ng1654)  &  (~ ng1648)  &  (~ ng823) ) ;
 assign wire32588 = ( (~ ng1654)  &  (~ ng826)  &  (~ ng1651) ) | ( (~ ng1654)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32590 = ( wire3046 ) | ( wire8231 ) | ( wire32587 ) ;
 assign wire32591 = ( wire8236 ) | ( wire8237 ) | ( wire32588 ) ;
 assign wire32597 = ( (~ ng1585)  &  (~ ng1588)  &  (~ ng1591) ) | ( (~ ng826)  &  (~ ng1588)  &  (~ ng1591) ) ;
 assign wire32598 = ( (~ ng1585)  &  (~ ng823)  &  (~ ng1591) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng1591) ) ;
 assign wire32600 = ( wire3046 ) | ( wire8247 ) | ( wire32597 ) ;
 assign wire32601 = ( wire8252 ) | ( wire8253 ) | ( wire32598 ) ;
 assign wire32607 = ( (~ ng1582)  &  (~ ng1579)  &  (~ ng1576) ) | ( (~ ng1582)  &  (~ ng823)  &  (~ ng1576) ) ;
 assign wire32608 = ( (~ ng1582)  &  (~ ng1579)  &  (~ ng826) ) | ( (~ ng1582)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32610 = ( wire3046 ) | ( wire8207 ) | ( wire32607 ) ;
 assign wire32611 = ( wire8212 ) | ( wire8213 ) | ( wire32608 ) ;
 assign wire32617 = ( (~ ng1642)  &  (~ ng853)  &  (~ ng1639) ) | ( (~ ng1642)  &  (~ ng1645)  &  (~ ng1639) ) ;
 assign wire32618 = ( (~ ng1642)  &  (~ ng826)  &  (~ ng1645) ) | ( (~ ng826)  &  (~ ng823)  &  (~ ng1645) ) ;
 assign wire32620 = ( wire3046 ) | ( wire8223 ) | ( wire32617 ) ;
 assign wire32621 = ( wire8228 ) | ( wire8229 ) | ( wire32618 ) ;
 assign wire32630 = ( wire3046 ) | ( wire8167 ) | ( wire8168 ) | ( wire8169 ) ;
 assign wire32631 = ( wire8170 ) | ( wire8171 ) | ( wire8172 ) | ( wire8173 ) ;
 assign wire32637 = ( ng1693  &  ng1695  &  ng1694 ) | ( (~ ng826)  &  ng1695  &  ng1694 ) ;
 assign wire32638 = ( ng1693  &  ng1695  &  (~ ng823) ) | ( (~ ng826)  &  ng1695  &  (~ ng823) ) ;
 assign wire32640 = ( wire3046 ) | ( wire8159 ) | ( wire32637 ) ;
 assign wire32641 = ( wire8164 ) | ( wire8165 ) | ( wire32638 ) ;
 assign wire32647 = ( ng1696  &  ng1697  &  ng1698 ) | ( ng1697  &  ng1698  &  (~ ng826) ) ;
 assign wire32648 = ( ng1696  &  ng1698  &  (~ ng823) ) | ( ng1698  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32650 = ( wire3046 ) | ( wire8151 ) | ( wire32647 ) ;
 assign wire32651 = ( wire8156 ) | ( wire8157 ) | ( wire32648 ) ;
 assign wire32652 = ( wire32630  &  wire32640 ) | ( wire32631  &  wire32640 ) | ( wire32630  &  wire32641 ) | ( wire32631  &  wire32641 ) ;
 assign wire32658 = ( (~ ng826)  &  (~ ng1636)  &  (~ ng1633) ) | ( (~ ng1636)  &  (~ ng1630)  &  (~ ng1633) ) ;
 assign wire32659 = ( (~ ng826)  &  (~ ng1636)  &  (~ ng823) ) | ( (~ ng1636)  &  (~ ng823)  &  (~ ng1630) ) ;
 assign wire32661 = ( wire3046 ) | ( wire8215 ) | ( wire32658 ) ;
 assign wire32662 = ( wire8220 ) | ( wire8221 ) | ( wire32659 ) ;
 assign wire32668 = ( (~ ng1624)  &  (~ ng1621)  &  (~ ng1627) ) | ( (~ ng1621)  &  (~ ng823)  &  (~ ng1627) ) ;
 assign wire32671 = ( wire3046 ) | ( wire8199 ) | ( wire32668 ) ;
 assign wire32672 = ( wire8202 ) | ( wire8203 ) | ( wire8204 ) | ( wire8205 ) ;
 assign wire32678 = ( (~ ng1597)  &  (~ ng1600)  &  (~ ng826) ) | ( (~ ng1597)  &  (~ ng1600)  &  (~ ng1594) ) ;
 assign wire32679 = ( (~ ng1600)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng1600)  &  (~ ng1594)  &  (~ ng823) ) ;
 assign wire32681 = ( wire3046 ) | ( wire8191 ) | ( wire32678 ) ;
 assign wire32682 = ( wire8196 ) | ( wire8197 ) | ( wire32679 ) ;
 assign wire32688 = ( (~ ng826)  &  (~ ng1615)  &  (~ ng1618) ) | ( (~ ng1615)  &  (~ ng1612)  &  (~ ng1618) ) ;
 assign wire32689 = ( (~ ng826)  &  (~ ng823)  &  (~ ng1618) ) | ( (~ ng823)  &  (~ ng1612)  &  (~ ng1618) ) ;
 assign wire32691 = ( wire3046 ) | ( wire8183 ) | ( wire32688 ) ;
 assign wire32692 = ( wire8188 ) | ( wire8189 ) | ( wire32689 ) ;
 assign wire32698 = ( (~ ng826)  &  (~ ng1609)  &  (~ ng1606) ) | ( (~ ng1609)  &  (~ ng1606)  &  (~ ng1603) ) ;
 assign wire32699 = ( (~ ng826)  &  (~ ng823)  &  (~ ng1609) ) | ( (~ ng823)  &  (~ ng1609)  &  (~ ng1603) ) ;
 assign wire32701 = ( wire3046 ) | ( wire8175 ) | ( wire32698 ) ;
 assign wire32702 = ( wire8180 ) | ( wire8181 ) | ( wire32699 ) ;
 assign wire32703 = ( wire32630  &  wire32640 ) | ( wire32631  &  wire32640 ) | ( wire32630  &  wire32641 ) | ( wire32631  &  wire32641 ) ;
 assign wire32709 = ( (~ ng1573)  &  (~ ng1567)  &  (~ ng823) ) | ( (~ ng1573)  &  (~ ng1567)  &  (~ ng1570) ) ;
 assign wire32710 = ( (~ ng1573)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng1573)  &  (~ ng826)  &  (~ ng1570) ) ;
 assign wire32712 = ( wire3046 ) | ( wire8239 ) | ( wire32709 ) ;
 assign wire32713 = ( wire8244 ) | ( wire8245 ) | ( wire32710 ) ;
 assign wire32715 = ( (~ wire32590)  &  (~ wire32591)  &  wire32600 ) | ( (~ wire32590)  &  (~ wire32591)  &  wire32601 ) ;
 assign wire32716 = ( (~ wire32610)  &  (~ wire32611)  &  wire32620 ) | ( (~ wire32610)  &  (~ wire32611)  &  wire32621 ) ;
 assign wire32717 = ( wire32661  &  (~ wire32671)  &  (~ wire32672) ) | ( wire32662  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire32718 = ( wire32681  &  (~ wire32691)  &  (~ wire32692) ) | ( wire32682  &  (~ wire32691)  &  (~ wire32692) ) ;
 assign wire32721 = ( (~ wire32650)  &  (~ wire32651)  &  wire32652  &  wire32718 ) ;
 assign wire32722 = ( (~ ng12828)  &  wire32715  &  wire32716  &  wire32717 ) ;
 assign wire32724 = ( wire32590  &  wire32712 ) | ( wire32591  &  wire32712 ) | ( wire32590  &  wire32713 ) | ( wire32591  &  wire32713 ) ;
 assign wire32725 = ( wire32600  &  wire32610 ) | ( wire32601  &  wire32610 ) | ( wire32600  &  wire32611 ) | ( wire32601  &  wire32611 ) ;
 assign wire32726 = ( wire32620  &  wire32661 ) | ( wire32621  &  wire32661 ) | ( wire32620  &  wire32662 ) | ( wire32621  &  wire32662 ) ;
 assign wire32727 = ( wire32671  &  wire32681 ) | ( wire32672  &  wire32681 ) | ( wire32671  &  wire32682 ) | ( wire32672  &  wire32682 ) ;
 assign wire32728 = ( wire32691  &  wire32701 ) | ( wire32692  &  wire32701 ) | ( wire32691  &  wire32702 ) | ( wire32692  &  wire32702 ) ;
 assign wire32730 = ( wire32727  &  wire32726 ) ;
 assign wire32731 = ( wire32724  &  wire32725  &  wire32728 ) ;
 assign wire32740 = ( wire3046 ) | ( wire8054 ) | ( wire8055 ) | ( wire8056 ) ;
 assign wire32741 = ( wire8057 ) | ( wire8058 ) | ( wire8059 ) | ( wire8060 ) ;
 assign wire32742 = ( (~ ng853)  &  ng1530 ) ;
 assign wire32744 = ( ng1529  &  (~ ng826) ) ;
 assign wire32746 = ( ng1529  &  ng1530 ) ;
 assign wire32747 = ( ng1531  &  ng1491 ) | ( (~ ng823)  &  ng1491 ) ;
 assign wire32748 = ( ng1516  &  ng1514 ) ;
 assign wire32749 = ( ng1515  &  ng1476 ) | ( (~ ng826)  &  ng1476 ) ;
 assign wire32750 = ( ng1516  &  (~ ng853) ) ;
 assign wire32752 = ( ng1514  &  (~ ng823) ) ;
 assign wire32754 = ( (~ ng826)  &  (~ ng853)  &  ng1491 ) ;
 assign wire32755 = ( (~ ng823)  &  (~ ng853)  &  ng1476 ) ;
 assign wire32765 = ( ng1511  &  ng1512  &  ng1513 ) | ( ng1511  &  ng1513  &  (~ ng826) ) ;
 assign wire32766 = ( ng1511  &  ng1512  &  (~ ng823) ) | ( ng1511  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32769 = ( wire8103 ) | ( wire8104 ) | ( wire32766 ) ;
 assign wire32775 = ( ng1527  &  ng1526  &  ng1528 ) | ( ng1526  &  ng1528  &  (~ ng826) ) ;
 assign wire32776 = ( ng1527  &  ng1526  &  (~ ng823) ) | ( ng1526  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32778 = ( wire3046 ) | ( wire8106 ) | ( wire32775 ) ;
 assign wire32779 = ( wire8111 ) | ( wire8112 ) | ( wire32776 ) ;
 assign wire32785 = ( ng1523  &  ng1525  &  ng1524 ) | ( ng1523  &  ng1525  &  (~ ng826) ) ;
 assign wire32786 = ( ng1523  &  ng1524  &  (~ ng823) ) | ( ng1523  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32789 = ( wire8119 ) | ( wire8120 ) | ( wire32786 ) ;
 assign wire32792 = ( wire8090 ) | ( (~ ng1515)  &  ng826  &  (~ ng1476) ) ;
 assign wire32793 = ( ng1491  &  wire3321  &  wire32742 ) | ( ng1491  &  wire3321  &  wire32744 ) ;
 assign wire32794 = ( wire32746  &  wire32747 ) | ( wire32748  &  wire32749 ) ;
 assign wire32795 = ( ng1476  &  wire3320  &  wire32750 ) | ( ng1476  &  wire3320  &  wire32752 ) ;
 assign wire32796 = ( wire3321  &  wire32754 ) | ( wire3320  &  wire32755 ) ;
 assign wire32797 = ( wire8086 ) | ( wire8087 ) | ( wire8088 ) | ( wire8089 ) ;
 assign wire32800 = ( wire32797 ) | ( wire32796 ) ;
 assign wire32801 = ( wire32792 ) | ( wire32793 ) | ( wire32794 ) | ( wire32795 ) ;
 assign wire32806 = ( wire8094 ) | ( wire32800 ) | ( ng1471  &  ng11992 ) | ( (~ ng1471)  &  (~ ng11992) ) ;
 assign wire32807 = ( wire8095 ) | ( wire32801 ) | ( ng1481  &  ng11773 ) | ( (~ ng1481)  &  (~ ng11773) ) ;
 assign wire32816 = ( wire3046 ) | ( wire8130 ) | ( wire8131 ) | ( wire8132 ) ;
 assign wire32817 = ( wire8133 ) | ( wire8134 ) | ( wire8135 ) | ( wire8136 ) ;
 assign wire32819 = ( ng1541  &  ng1543  &  ng1542 ) | ( ng1541  &  ng1542  &  (~ ng823) ) ;
 assign wire32825 = ( ng1554  &  ng1555  &  ng1553 ) | ( ng1554  &  (~ ng823)  &  ng1553 ) ;
 assign wire32828 = ( wire3046 ) | ( wire8138 ) | ( wire32825 ) ;
 assign wire32829 = ( wire8141 ) | ( wire8142 ) | ( wire8143 ) | ( wire8144 ) ;
 assign wire32831 = ( ng1545  &  ng1544  &  ng1546 ) | ( ng1545  &  ng1544  &  (~ ng823) ) ;
 assign wire32833 = ( ng1543  &  ng1542  &  (~ ng853) ) ;
 assign wire32835 = ( ng1545  &  ng1546  &  (~ ng853) ) ;
 assign wire32837 = ( ng1541  &  (~ ng826)  &  ng1543 ) ;
 assign wire32839 = ( ng1544  &  ng1546  &  (~ ng826) ) ;
 assign wire32840 = ( ng1544  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32841 = ( ng1541  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32842 = ( ng1542  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire32843 = ( ng1545  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire32844 = ( (~ ng826)  &  ng1543  &  (~ ng853) ) ;
 assign wire32845 = ( ng1546  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire32846 = ( ng853  &  (~ ng1544) ) ;
 assign wire32847 = ( ng853  &  (~ ng1541) ) ;
 assign wire32848 = ( (~ ng1542)  &  ng826 ) ;
 assign wire32855 = ( ng1539  &  ng1540  &  ng1538 ) | ( ng1540  &  ng1538  &  (~ ng826) ) ;
 assign wire32856 = ( ng1539  &  ng1538  &  (~ ng823) ) | ( ng1538  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32858 = ( wire3046 ) | ( wire8062 ) | ( wire32855 ) ;
 assign wire32859 = ( wire8067 ) | ( wire8068 ) | ( wire32856 ) ;
 assign wire32865 = ( ng1534  &  ng1532  &  ng1533 ) | ( ng1532  &  ng1533  &  (~ ng823) ) ;
 assign wire32866 = ( ng1534  &  ng1532  &  (~ ng826) ) | ( ng1532  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32869 = ( wire8075 ) | ( wire8076 ) | ( wire32866 ) ;
 assign wire32875 = ( ng1535  &  ng1536  &  ng1537 ) | ( ng1535  &  ng1537  &  (~ ng826) ) ;
 assign wire32876 = ( ng1535  &  ng1536  &  (~ ng823) ) | ( ng1535  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32878 = ( wire3046 ) | ( wire8122 ) | ( wire32875 ) ;
 assign wire32879 = ( wire8127 ) | ( wire8128 ) | ( wire32876 ) ;
 assign wire32883 = ( (~ wire32828)  &  (~ wire32829)  &  wire32839 ) | ( (~ wire32828)  &  (~ wire32829)  &  wire32840 ) ;
 assign wire32884 = ( (~ wire32816)  &  (~ wire32817)  &  wire32841 ) | ( (~ wire32816)  &  (~ wire32817)  &  wire32842 ) ;
 assign wire32886 = ( wire32828  &  wire32846 ) | ( wire32829  &  wire32846 ) | ( (~ wire32828)  &  (~ wire32829)  &  wire32845 ) ;
 assign wire32887 = ( wire32816  &  wire32847 ) | ( wire32817  &  wire32847 ) | ( wire32816  &  wire32848 ) | ( wire32817  &  wire32848 ) ;
 assign wire32893 = ( wire3386 ) | ( wire8026 ) | ( wire8051 ) ;
 assign wire32894 = ( wire8027 ) | ( wire8028 ) | ( wire8029 ) | ( wire8030 ) ;
 assign wire32895 = ( wire32884 ) | ( wire32883 ) ;
 assign wire32896 = ( wire8035 ) | ( wire8036 ) | ( wire32886 ) ;
 assign wire32897 = ( wire8041 ) | ( wire8042 ) | ( wire32887 ) ;
 assign wire32898 = ( wire8043 ) | ( wire8044 ) | ( wire8046 ) ;
 assign wire32899 = ( wire8047 ) | ( wire8050 ) | ( ng1496  &  ng11839 ) | ( (~ ng1496)  &  (~ ng11839) ) ;
 assign wire32902 = ( wire8041 ) | ( wire8042 ) | ( wire32887 ) | ( wire32898 ) ;
 assign wire32903 = ( wire32806 ) | ( wire32807 ) | ( wire32899 ) ;
 assign wire32904 = ( wire32893 ) | ( wire32894 ) | ( wire32895 ) | ( wire32896 ) ;
 assign wire32906 = ( ng853  &  (~ ng1783) ) ;
 assign wire32907 = ( (~ ng1784)  &  ng826 ) ;
 assign wire32908 = ( ng823  &  (~ ng1785) ) ;
 assign wire32918 = ( wire3386 ) | ( (~ ng18514)  &  (~ ng18383)  &  wire3068 ) ;
 assign wire32921 = ( (~ ng18561)  &  (~ ng18458)  &  (~ ng18514) ) | ( (~ ng18561)  &  (~ ng18458)  &  (~ ng18383) ) | ( (~ ng18561)  &  (~ ng18514)  &  (~ ng18383) ) | ( (~ ng18458)  &  (~ ng18514)  &  (~ ng18383) ) ;
 assign wire32922 = ( wire3068  &  wire3291 ) | ( (~ ng18561)  &  (~ ng18458)  &  wire3291 ) ;
 assign wire32923 = ( wire8009 ) | ( wire8010 ) | ( wire32918 ) ;
 assign wire32924 = ( wire8004 ) | ( wire8011 ) | ( wire32921 ) ;
 assign wire32934 = ( wire3386 ) | ( (~ ng18212)  &  (~ ng18115)  &  wire3108 ) ;
 assign wire32937 = ( (~ ng17942)  &  (~ ng18556)  &  (~ ng18212) ) | ( (~ ng17942)  &  (~ ng18556)  &  (~ ng18115) ) | ( (~ ng17942)  &  (~ ng18212)  &  (~ ng18115) ) | ( (~ ng18556)  &  (~ ng18212)  &  (~ ng18115) ) ;
 assign wire32938 = ( wire3108  &  wire3297 ) | ( (~ ng17942)  &  (~ ng18556)  &  wire3297 ) ;
 assign wire32939 = ( wire7987 ) | ( wire7988 ) | ( wire32934 ) ;
 assign wire32940 = ( wire7982 ) | ( wire7989 ) | ( wire32937 ) ;
 assign wire32942 = ( wire32630  &  (~ wire32640)  &  (~ wire32641) ) | ( wire32631  &  (~ wire32640)  &  (~ wire32641) ) ;
 assign wire32943 = ( (~ wire32902)  &  (~ wire32903)  &  (~ wire32904)  &  wire32942 ) ;
 assign wire32944 = ( (~ wire32630)  &  (~ wire32631)  &  (~ wire32640)  &  (~ wire32641) ) ;
 assign wire32945 = ( (~ ng1703)  &  ng826 ) | ( ng853  &  (~ ng1702) ) ;
 assign wire32946 = ( wire7976  &  wire32650 ) | ( wire7976  &  wire32651 ) | ( wire32650  &  wire32945 ) | ( wire32651  &  wire32945 ) ;
 assign wire32947 = ( wire7972 ) | ( wire7977 ) | ( wire7978 ) | ( wire7979 ) ;
 assign wire32952 = ( (~ wire32610)  &  (~ wire32611)  &  wire32671 ) | ( (~ wire32610)  &  (~ wire32611)  &  wire32672 ) | ( wire32610  &  (~ wire32671)  &  (~ wire32672) ) | ( wire32611  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire32954 = ( (~ ng13001)  &  ng12930 ) | ( ng11666  &  (~ ng12930) ) | ( (~ ng12930)  &  (~ wire32652) ) | ( ng13001  &  (~ ng11666)  &  wire32652 ) ;
 assign wire32956 = ( (~ ng12949)  &  ng12797 ) | ( ng11666  &  (~ ng12797) ) | ( (~ ng12797)  &  (~ wire32652) ) | ( (~ ng11666)  &  ng12949  &  wire32652 ) ;
 assign wire32957 = ( (~ ng12797)  &  (~ wire32650)  &  (~ wire32651)  &  wire32652 ) ;
 assign wire32958 = ( ng27582  &  (~ wire32952)  &  (~ wire32954)  &  wire32957 ) ;
 assign wire32959 = ( (~ wire32620)  &  (~ wire32621)  &  (~ wire32681)  &  (~ wire32682) ) ;
 assign wire32960 = ( (~ ng12949)  &  (~ wire32650)  &  (~ wire32651)  &  wire32652 ) ;
 assign wire32961 = ( (~ ng12949)  &  (~ ng27582) ) | ( (~ ng12949)  &  wire32952 ) | ( (~ ng12949)  &  wire32954 ) ;
 assign wire32962 = ( (~ ng28556)  &  wire32961 ) | ( (~ ng28556)  &  ng26918  &  wire32958 ) ;
 assign wire32963 = ( (~ ng28556)  &  ng26918  &  wire32959 ) | ( (~ ng28556)  &  ng26918  &  wire32960 ) ;
 assign wire32975 = ( ng1453  &  ng1466  &  ng1457  &  ng1462 ) ;
 assign wire32977 = ( ng1457  &  (~ ng17031)  &  (~ ng23528) ) ;
 assign wire32979 = ( (~ wire32630)  &  (~ wire32631)  &  wire32640 ) | ( (~ wire32630)  &  (~ wire32631)  &  wire32641 ) ;
 assign wire32985 = ( ng1765  &  ng1757  &  ng1754 ) | ( ng1757  &  ng1754  &  (~ ng826) ) ;
 assign wire32986 = ( ng1765  &  ng1757  &  (~ ng823) ) | ( ng1757  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire32988 = ( wire3046 ) | ( wire7922 ) | ( wire32985 ) ;
 assign wire32989 = ( wire7927 ) | ( wire7928 ) | ( wire32986 ) ;
 assign wire32995 = ( ng1735  &  ng1724  &  (~ ng853) ) | ( ng1735  &  ng1724  &  ng1727 ) ;
 assign wire32996 = ( ng1735  &  (~ ng823)  &  ng1727 ) | ( (~ ng826)  &  (~ ng823)  &  ng1727 ) ;
 assign wire32998 = ( wire3046 ) | ( wire7914 ) | ( wire32995 ) ;
 assign wire32999 = ( wire7919 ) | ( wire7920 ) | ( wire32996 ) ;
 assign wire33008 = ( wire3046 ) | ( wire7930 ) | ( wire7931 ) | ( wire7932 ) ;
 assign wire33009 = ( wire7933 ) | ( wire7934 ) | ( wire7935 ) | ( wire7936 ) ;
 assign wire33018 = ( wire3046 ) | ( wire7900 ) | ( wire7901 ) | ( wire7902 ) ;
 assign wire33019 = ( wire7903 ) | ( wire7904 ) | ( wire7905 ) | ( wire7906 ) ;
 assign wire33023 = ( ng1481  &  ng1486  &  ng1491  &  ng1506 ) ;
 assign wire33024 = ( ng1496  &  ng1471  &  ng1476  &  ng1501 ) ;
 assign wire33025 = ( wire32828 ) | ( wire32829 ) | ( (~ wire33023) ) | ( (~ wire33024) ) ;
 assign wire33033 = ( (~ ng1792)  &  (~ ng1795)  &  (~ ng1789) ) | ( (~ ng1795)  &  (~ ng823)  &  (~ ng1789) ) ;
 assign wire33034 = ( (~ ng1792)  &  (~ ng1795)  &  (~ ng826) ) | ( (~ ng1795)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33036 = ( wire3046 ) | ( wire7892 ) | ( wire33033 ) ;
 assign wire33037 = ( wire7897 ) | ( wire7898 ) | ( wire33034 ) ;
 assign wire33039 = ( ng1809  &  ng1808  &  (~ ng853) ) ;
 assign wire33041 = ( ng1809  &  ng1807  &  (~ ng826) ) ;
 assign wire33043 = ( ng1809  &  ng1807  &  ng1808 ) ;
 assign wire33045 = ( ng1807  &  ng1808  &  (~ ng823) ) ;
 assign wire33046 = ( ng1807  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33047 = ( ng1808  &  (~ ng823)  &  (~ ng853) ) ;
 assign wire33048 = ( ng1809  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire33053 = ( wire7881 ) | ( wire7882 ) | ( wire7883 ) | ( wire7884 ) ;
 assign wire33054 = ( wire7885 ) | ( wire7886 ) | ( wire7887 ) | ( wire7888 ) ;
 assign wire33063 = ( wire3046 ) | ( wire7867 ) | ( wire7868 ) | ( wire7869 ) ;
 assign wire33064 = ( wire7870 ) | ( wire7871 ) | ( wire7872 ) | ( wire7873 ) ;
 assign wire33070 = ( (~ ng1816)  &  (~ ng823)  &  (~ ng1810) ) | ( (~ ng1816)  &  (~ ng1813)  &  (~ ng1810) ) ;
 assign wire33071 = ( (~ ng1816)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng1816)  &  (~ ng826)  &  (~ ng1813) ) ;
 assign wire33074 = ( wire7855 ) | ( wire7856 ) | ( wire33071 ) ;
 assign wire33080 = ( ng1560  &  ng1561  &  ng1559 ) | ( ng1561  &  (~ ng826)  &  ng1559 ) ;
 assign wire33081 = ( ng1560  &  ng1559  &  (~ ng823) ) | ( (~ ng826)  &  ng1559  &  (~ ng823) ) ;
 assign wire33083 = ( wire3046 ) | ( wire7858 ) | ( (~ wire33023) ) | ( (~ wire33024) ) ;
 assign wire33084 = ( wire33081 ) | ( wire33080 ) ;
 assign wire33087 = ( (~ ng1830)  &  ng823  &  ng2257 ) ;
 assign wire33088 = ( (~ ng1829)  &  ng826  &  ng2257 ) ;
 assign wire33089 = ( (~ ng1828)  &  ng853  &  ng2257 ) ;
 assign wire33091 = ( wire32650  &  (~ wire32703) ) | ( wire32651  &  (~ wire32703) ) ;
 assign wire33097 = ( (~ ng1496)  &  (~ ng18115)  &  wire32661 ) | ( (~ ng1496)  &  (~ ng18115)  &  wire32662 ) | ( ng1496  &  (~ ng18115)  &  (~ wire32661)  &  (~ wire32662) ) ;
 assign wire33098 = ( (~ ng18561)  &  (~ ng17942)  &  (~ ng18458)  &  (~ ng18514) ) ;
 assign wire33099 = ( (~ ng18383)  &  wire3068  &  (~ ng18556)  &  (~ ng18212) ) ;
 assign wire33101 = ( (~ wire32630)  &  (~ wire32631)  &  (~ wire32650)  &  (~ wire32651) ) ;
 assign wire33102 = ( ng23526  &  wire33101 ) ;
 assign wire33103 = ( wire32630  &  (~ wire32650)  &  (~ wire32651) ) | ( wire32631  &  (~ wire32650)  &  (~ wire32651) ) ;
 assign wire33105 = ( (~ ng11675)  &  ng11630 ) | ( (~ ng2257)  &  (~ ng11675)  &  ng11666 ) | ( (~ ng2257)  &  (~ ng11630)  &  ng11666 ) | ( (~ ng11675)  &  (~ ng11630)  &  ng11666 ) ;
 assign wire33106 = ( wire33105 ) | ( (~ ng23518)  &  wire33091 ) | ( (~ ng23505)  &  wire33091 ) ;
 assign wire33107 = ( (~ ng11675)  &  (~ wire7977)  &  (~ wire7978)  &  (~ wire7979) ) ;
 assign wire33108 = ( ng11675  &  (~ wire7977)  &  (~ wire7978)  &  (~ wire7979) ) ;
 assign wire33115 = ( (~ ng1312)  &  (~ ng1315)  &  ng1962 ) | ( (~ ng1315)  &  ng1962  &  ng1963 ) ;
 assign wire33117 = ( wire3049 ) | ( wire7815 ) | ( wire7816 ) | ( wire7817 ) ;
 assign wire33118 = ( wire7820 ) | ( wire7821 ) | ( wire33115 ) ;
 assign wire33124 = ( ng1959  &  ng1960  &  ng1958 ) | ( ng1959  &  (~ ng1312)  &  ng1958 ) ;
 assign wire33125 = ( ng1959  &  ng1960  &  (~ ng1315) ) | ( ng1959  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire33127 = ( wire3049 ) | ( wire7797 ) | ( wire33124 ) ;
 assign wire33128 = ( wire7802 ) | ( wire7803 ) | ( wire33125 ) ;
 assign wire33135 = ( (~ ng1312)  &  (~ ng1315)  &  ng1956 ) | ( (~ ng1315)  &  ng1956  &  ng1957 ) ;
 assign wire33137 = ( wire3049 ) | ( wire7807 ) | ( wire7808 ) | ( wire7809 ) ;
 assign wire33138 = ( wire7812 ) | ( wire7813 ) | ( wire33135 ) ;
 assign wire33144 = ( (~ ng1309)  &  (~ ng1997)  &  (~ ng2000) ) | ( (~ ng1994)  &  (~ ng1997)  &  (~ ng2000) ) ;
 assign wire33145 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1994) ) | ( (~ ng1315)  &  (~ ng1994)  &  (~ ng1997) ) ;
 assign wire33147 = ( wire3049 ) | ( wire7779 ) | ( wire33144 ) ;
 assign wire33148 = ( wire7784 ) | ( wire7785 ) | ( wire33145 ) ;
 assign wire33154 = ( (~ ng1871)  &  (~ ng1312)  &  (~ ng1877) ) | ( (~ ng1871)  &  (~ ng1874)  &  (~ ng1877) ) ;
 assign wire33155 = ( (~ ng1871)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng1871)  &  (~ ng1315)  &  (~ ng1874) ) ;
 assign wire33157 = ( wire3049 ) | ( wire7771 ) | ( wire33154 ) ;
 assign wire33158 = ( wire7776 ) | ( wire7777 ) | ( wire33155 ) ;
 assign wire33164 = ( (~ ng1991)  &  (~ ng1309)  &  (~ ng1988) ) | ( (~ ng1991)  &  (~ ng1985)  &  (~ ng1988) ) ;
 assign wire33165 = ( (~ ng1991)  &  (~ ng1312)  &  (~ ng1985) ) | ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1985) ) ;
 assign wire33167 = ( wire3049 ) | ( wire7787 ) | ( wire33164 ) ;
 assign wire33168 = ( wire7792 ) | ( wire7793 ) | ( wire33165 ) ;
 assign wire33184 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1949) ) | ( (~ ng1315)  &  (~ ng1949)  &  (~ ng1951) ) ;
 assign wire33186 = ( wire3049 ) | ( wire7758 ) | ( wire7759 ) | ( wire7760 ) ;
 assign wire33187 = ( wire7763 ) | ( wire7764 ) | ( wire33184 ) ;
 assign wire33189 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1967) ) ;
 assign wire33191 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1967) ) ;
 assign wire33193 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1967) ) ;
 assign wire33201 = ( (~ ng1973)  &  (~ ng1970)  &  (~ ng1309) ) ;
 assign wire33205 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1967) ) ;
 assign wire33208 = ( (~ ng1973)  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire33211 = ( (~ ng1970)  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire33221 = ( wire7734 ) | ( wire7735 ) | ( wire7736 ) | ( wire7737 ) ;
 assign wire33222 = ( wire7741 ) | ( wire7742 ) | ( wire7743 ) | ( wire7745 ) ;
 assign wire33223 = ( wire7746 ) | ( wire7748 ) | ( wire7749 ) | ( wire7751 ) ;
 assign wire33224 = ( wire7752 ) | ( wire7754 ) | ( wire7755 ) | ( wire7757 ) ;
 assign wire33226 = ( wire33224 ) | ( wire33223 ) ;
 assign wire33228 = ( wire33186  &  wire33191 ) | ( wire33187  &  wire33191 ) | ( wire33186  &  wire33193 ) | ( wire33187  &  wire33193 ) ;
 assign wire33229 = ( wire33186  &  wire33201 ) | ( wire33187  &  wire33201 ) | ( wire33186  &  wire33205 ) | ( wire33187  &  wire33205 ) ;
 assign wire33230 = ( wire33186  &  wire33208 ) | ( wire33187  &  wire33208 ) | ( wire33186  &  wire33211 ) | ( wire33187  &  wire33211 ) ;
 assign wire33231 = ( wire7756 ) | ( wire33223 ) | ( wire33224 ) ;
 assign wire33232 = ( wire7738 ) | ( wire33221 ) | ( wire33222 ) | ( wire33228 ) ;
 assign wire33233 = ( wire33230 ) | ( wire33229 ) ;
 assign wire33248 = ( (~ ng1945)  &  (~ ng1312)  &  (~ ng1870) ) | ( (~ ng1945)  &  (~ ng1947)  &  (~ ng1870) ) ;
 assign wire33249 = ( (~ ng1945)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng1945)  &  (~ ng1315)  &  (~ ng1947) ) ;
 assign wire33251 = ( wire3049 ) | ( wire7724 ) | ( wire33248 ) ;
 assign wire33252 = ( wire7729 ) | ( wire7730 ) | ( wire33249 ) ;
 assign wire33254 = ( (~ ng1979)  &  (~ ng1309)  &  (~ ng1982) ) ;
 assign wire33256 = ( (~ ng1979)  &  (~ ng1976)  &  (~ ng1982) ) ;
 assign wire33258 = ( (~ ng1312)  &  (~ ng1976)  &  (~ ng1982) ) ;
 assign wire33260 = ( (~ ng1315)  &  (~ ng1979)  &  (~ ng1976) ) ;
 assign wire33270 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1976) ) ;
 assign wire33273 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng1982) ) ;
 assign wire33276 = ( (~ ng1315)  &  (~ ng1979)  &  (~ ng1309) ) ;
 assign wire33286 = ( wire7700 ) | ( wire7701 ) | ( wire7702 ) | ( wire7703 ) ;
 assign wire33287 = ( wire7708 ) | ( wire7709 ) | ( wire7710 ) | ( wire7711 ) ;
 assign wire33288 = ( wire7712 ) | ( wire7714 ) | ( wire7715 ) | ( wire7717 ) ;
 assign wire33289 = ( wire7718 ) | ( wire7720 ) | ( wire7721 ) | ( wire7723 ) ;
 assign wire33293 = ( wire33251  &  wire33256 ) | ( wire33252  &  wire33256 ) | ( wire33251  &  wire33258 ) | ( wire33252  &  wire33258 ) ;
 assign wire33294 = ( wire33251  &  wire33260 ) | ( wire33252  &  wire33260 ) | ( wire33251  &  wire33270 ) | ( wire33252  &  wire33270 ) ;
 assign wire33295 = ( wire33251  &  wire33273 ) | ( wire33252  &  wire33273 ) | ( wire33251  &  wire33276 ) | ( wire33252  &  wire33276 ) ;
 assign wire33296 = ( wire3049 ) | ( wire33288 ) | ( wire33289 ) ;
 assign wire33297 = ( wire7704 ) | ( wire33286 ) | ( wire33287 ) | ( wire33293 ) ;
 assign wire33298 = ( wire33295 ) | ( wire33294 ) ;
 assign wire33306 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1760) ) | ( (~ ng1312)  &  (~ ng1760)  &  (~ ng1764) ) ;
 assign wire33308 = ( wire3049 ) | ( wire7692 ) | ( wire7693 ) | ( wire7694 ) ;
 assign wire33309 = ( wire7697 ) | ( wire7698 ) | ( wire33306 ) ;
 assign wire33318 = ( wire3049 ) | ( wire7684 ) | ( wire7685 ) | ( wire7686 ) ;
 assign wire33319 = ( wire7687 ) | ( wire7688 ) | ( wire7689 ) | ( wire7690 ) ;
 assign wire33326 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng1730) ) | ( (~ ng1315)  &  (~ ng1730)  &  (~ ng1732) ) ;
 assign wire33328 = ( wire3049 ) | ( wire7676 ) | ( wire7677 ) | ( wire7678 ) ;
 assign wire33329 = ( wire7681 ) | ( wire7682 ) | ( wire33326 ) ;
 assign wire33336 = ( (~ ng1312)  &  (~ ng1315)  &  ng1965 ) | ( (~ ng1315)  &  ng1966  &  ng1965 ) ;
 assign wire33338 = ( wire3049 ) | ( wire7660 ) | ( wire7661 ) | ( wire7662 ) ;
 assign wire33339 = ( wire7665 ) | ( wire7666 ) | ( wire33336 ) ;
 assign wire33340 = ( (~ wire33308)  &  (~ wire33309)  &  wire33318 ) | ( (~ wire33308)  &  (~ wire33309)  &  wire33319 ) ;
 assign wire33341 = ( (~ wire33137)  &  (~ wire33138)  &  (~ wire33328)  &  (~ wire33329) ) ;
 assign wire33343 = ( wire33308  &  (~ wire33318)  &  (~ wire33319) ) | ( wire33309  &  (~ wire33318)  &  (~ wire33319) ) ;
 assign wire33353 = ( wire3049 ) | ( wire7668 ) | ( wire7669 ) | ( wire7670 ) ;
 assign wire33354 = ( wire7671 ) | ( wire7672 ) | ( wire7673 ) | ( wire7674 ) ;
 assign wire33355 = ( (~ wire33318)  &  (~ wire33319)  &  (~ wire33353)  &  (~ wire33354) ) ;
 assign wire33357 = ( wire33127  &  wire33338 ) | ( wire33128  &  wire33338 ) | ( wire33127  &  wire33339 ) | ( wire33128  &  wire33339 ) ;
 assign wire33359 = ( (~ wire33117)  &  (~ wire33118)  &  (~ wire33318)  &  (~ wire33319) ) ;
 assign wire33361 = ( wire33308  &  wire33338 ) | ( wire33309  &  wire33338 ) | ( wire33308  &  wire33339 ) | ( wire33309  &  wire33339 ) ;
 assign wire33363 = ( (~ wire33308)  &  (~ wire33309)  &  wire33318 ) | ( (~ wire33308)  &  (~ wire33309)  &  wire33319 ) ;
 assign wire33364 = ( (~ wire33127)  &  (~ wire33128)  &  wire33137 ) | ( (~ wire33127)  &  (~ wire33128)  &  wire33138 ) ;
 assign wire33365 = ( (~ wire33137)  &  (~ wire33138)  &  wire33353 ) | ( (~ wire33137)  &  (~ wire33138)  &  wire33354 ) ;
 assign wire33366 = ( (~ wire33328)  &  (~ wire33329)  &  (~ wire33338)  &  (~ wire33339) ) ;
 assign wire33367 = ( (~ wire33127)  &  (~ wire33128)  &  wire33308 ) | ( (~ wire33127)  &  (~ wire33128)  &  wire33309 ) ;
 assign wire33368 = ( (~ wire33117)  &  (~ wire33118)  &  wire33318 ) | ( (~ wire33117)  &  (~ wire33118)  &  wire33319 ) ;
 assign wire33369 = ( wire33318  &  wire33328 ) | ( wire33319  &  wire33328 ) | ( wire33318  &  wire33329 ) | ( wire33319  &  wire33329 ) ;
 assign wire33370 = ( wire33363  &  wire33364 ) | ( wire3440  &  wire33365 ) ;
 assign wire33371 = ( wire3437  &  wire33366 ) | ( wire3364  &  wire33367 ) ;
 assign wire33372 = ( wire3354  &  wire33368 ) | ( (~ wire3233)  &  wire33369 ) ;
 assign wire33376 = ( wire7650 ) | ( wire7651 ) | ( wire33372 ) ;
 assign wire33377 = ( wire7652 ) | ( wire7653 ) | ( wire33370 ) | ( wire33371 ) ;
 assign wire33378 = ( wire33127  &  wire33137 ) | ( wire33128  &  wire33137 ) | ( wire33127  &  wire33138 ) | ( wire33128  &  wire33138 ) ;
 assign wire33380 = ( (~ wire33318)  &  (~ wire33319)  &  (~ wire33328)  &  (~ wire33329) ) ;
 assign wire33382 = ( wire33308  &  (~ wire33328)  &  (~ wire33329) ) | ( wire33309  &  (~ wire33328)  &  (~ wire33329) ) ;
 assign wire33383 = ( (~ wire33127)  &  (~ wire33128)  &  wire33382 ) ;
 assign wire33384 = ( (~ wire33117)  &  (~ wire33118)  &  wire33318 ) | ( (~ wire33117)  &  (~ wire33118)  &  wire33319 ) ;
 assign wire33385 = ( (~ wire33137)  &  (~ wire33138)  &  wire33384 ) ;
 assign wire33387 = ( wire33127  &  wire33318 ) | ( wire33128  &  wire33318 ) | ( wire33127  &  wire33319 ) | ( wire33128  &  wire33319 ) ;
 assign wire33388 = ( (~ wire33338)  &  (~ wire33339)  &  (~ wire33353)  &  (~ wire33354) ) ;
 assign wire33390 = ( wire33308  &  wire33328 ) | ( wire33309  &  wire33328 ) | ( wire33308  &  wire33329 ) | ( wire33309  &  wire33329 ) ;
 assign wire33391 = ( (~ wire33117)  &  (~ wire33118)  &  wire33137 ) | ( (~ wire33117)  &  (~ wire33118)  &  wire33138 ) ;
 assign wire33392 = ( wire3364  &  wire33387 ) | ( wire3364  &  wire33388 ) ;
 assign wire33393 = ( (~ ng12291)  &  wire33390 ) | ( ng10851  &  ng12291  &  wire3354 ) ;
 assign wire33398 = ( wire7639 ) | ( wire7641 ) | ( wire7644 ) | ( wire33392 ) ;
 assign wire33399 = ( wire7638 ) | ( wire7649 ) | ( wire33393 ) | ( wire33398 ) ;
 assign wire33401 = ( (~ wire33376)  &  (~ wire33377)  &  wire33383 ) | ( (~ wire33376)  &  (~ wire33377)  &  wire33385 ) ;
 assign wire33402 = ( ng13055  &  wire33296 ) | ( ng13055  &  wire33297 ) | ( ng13055  &  wire33298 ) ;
 assign wire33403 = ( (~ wire33231)  &  (~ wire33232)  &  (~ wire33233)  &  wire33402 ) ;
 assign wire33404 = ( ng13055  &  wire33231 ) | ( ng13055  &  wire33232 ) | ( ng13055  &  wire33233 ) ;
 assign wire33405 = ( wire33376  &  wire33404 ) | ( wire33377  &  wire33404 ) ;
 assign wire33413 = ( ng2020  &  ng2033 ) ;
 assign wire33414 = ( ng1315  &  ng2013  &  (~ ng2039) ) ;
 assign wire33415 = ( (~ ng1312)  &  ng2013 ) | ( ng2013  &  (~ ng2010) ) ;
 assign wire33416 = ( (~ ng2033)  &  wire33415 ) | ( (~ ng2020)  &  wire33415 ) | ( (~ wire33414)  &  wire33415 ) ;
 assign wire33417 = ( ng2033  &  (~ ng1312) ) | ( ng2033  &  (~ ng2010) ) ;
 assign wire33425 = ( ng2251  &  ng2250  &  ng2252 ) | ( ng2250  &  ng2252  &  (~ ng826) ) ;
 assign wire33426 = ( ng2251  &  ng2250  &  (~ ng823) ) | ( ng2250  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33428 = ( wire3046 ) | ( wire7612 ) | ( wire33425 ) ;
 assign wire33429 = ( wire7617 ) | ( wire7618 ) | ( wire33426 ) ;
 assign wire33438 = ( wire3046 ) | ( wire7600 ) | ( wire7601 ) | ( wire7602 ) ;
 assign wire33439 = ( wire7603 ) | ( wire7604 ) | ( wire7605 ) | ( wire7606 ) ;
 assign wire33445 = ( (~ ng2270)  &  (~ ng2273)  &  (~ ng2276) ) | ( (~ ng2273)  &  (~ ng2276)  &  (~ ng826) ) ;
 assign wire33446 = ( (~ ng2270)  &  (~ ng2276)  &  (~ ng823) ) | ( (~ ng2276)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33448 = ( wire3046 ) | ( wire7592 ) | ( wire33445 ) ;
 assign wire33449 = ( wire7597 ) | ( wire7598 ) | ( wire33446 ) ;
 assign wire33458 = ( wire3046 ) | ( wire7584 ) | ( wire7585 ) | ( wire7586 ) ;
 assign wire33459 = ( wire7587 ) | ( wire7588 ) | ( wire7589 ) | ( wire7590 ) ;
 assign wire33468 = ( wire3046 ) | ( wire7576 ) | ( wire7577 ) | ( wire7578 ) ;
 assign wire33469 = ( wire7579 ) | ( wire7580 ) | ( wire7581 ) | ( wire7582 ) ;
 assign wire33475 = ( (~ ng2339)  &  (~ ng826)  &  (~ ng2336) ) | ( (~ ng2339)  &  (~ ng2333)  &  (~ ng2336) ) ;
 assign wire33476 = ( (~ ng2339)  &  (~ ng826)  &  (~ ng823) ) | ( (~ ng2339)  &  (~ ng2333)  &  (~ ng823) ) ;
 assign wire33478 = ( wire3046 ) | ( wire7568 ) | ( wire33475 ) ;
 assign wire33479 = ( wire7573 ) | ( wire7574 ) | ( wire33476 ) ;
 assign wire33485 = ( (~ ng2315)  &  (~ ng2318)  &  (~ ng2321) ) | ( (~ ng2318)  &  (~ ng826)  &  (~ ng2321) ) ;
 assign wire33486 = ( (~ ng2315)  &  (~ ng2321)  &  (~ ng823) ) | ( (~ ng826)  &  (~ ng2321)  &  (~ ng823) ) ;
 assign wire33488 = ( wire3046 ) | ( wire7560 ) | ( wire33485 ) ;
 assign wire33489 = ( wire7565 ) | ( wire7566 ) | ( wire33486 ) ;
 assign wire33498 = ( wire3046 ) | ( wire7552 ) | ( wire7553 ) | ( wire7554 ) ;
 assign wire33499 = ( wire7555 ) | ( wire7556 ) | ( wire7557 ) | ( wire7558 ) ;
 assign wire33505 = ( (~ ng2312)  &  (~ ng2306)  &  (~ ng2309) ) | ( (~ ng2312)  &  (~ ng2309)  &  (~ ng826) ) ;
 assign wire33506 = ( (~ ng2312)  &  (~ ng2306)  &  (~ ng823) ) | ( (~ ng2312)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33508 = ( wire3046 ) | ( wire7544 ) | ( wire33505 ) ;
 assign wire33509 = ( wire7549 ) | ( wire7550 ) | ( wire33506 ) ;
 assign wire33515 = ( (~ ng2285)  &  (~ ng2282)  &  (~ ng2279) ) | ( (~ ng2285)  &  (~ ng823)  &  (~ ng2279) ) ;
 assign wire33516 = ( (~ ng2285)  &  (~ ng2282)  &  (~ ng826) ) | ( (~ ng2285)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33518 = ( wire3046 ) | ( wire7536 ) | ( wire33515 ) ;
 assign wire33519 = ( wire7541 ) | ( wire7542 ) | ( wire33516 ) ;
 assign wire33528 = ( wire3046 ) | ( wire7520 ) | ( wire7521 ) | ( wire7522 ) ;
 assign wire33529 = ( wire7523 ) | ( wire7524 ) | ( wire7525 ) | ( wire7526 ) ;
 assign wire33535 = ( ng2387  &  ng2389  &  ng2388 ) | ( (~ ng826)  &  ng2389  &  ng2388 ) ;
 assign wire33536 = ( ng2387  &  ng2389  &  (~ ng823) ) | ( (~ ng826)  &  ng2389  &  (~ ng823) ) ;
 assign wire33538 = ( wire3046 ) | ( wire7504 ) | ( wire33535 ) ;
 assign wire33539 = ( wire7509 ) | ( wire7510 ) | ( wire33536 ) ;
 assign wire33545 = ( (~ ng823)  &  ng2390  &  ng2392 ) | ( ng2391  &  ng2390  &  ng2392 ) ;
 assign wire33546 = ( (~ ng826)  &  (~ ng823)  &  ng2392 ) | ( (~ ng826)  &  ng2391  &  ng2392 ) ;
 assign wire33548 = ( wire3046 ) | ( wire7512 ) | ( wire33545 ) ;
 assign wire33549 = ( wire7517 ) | ( wire7518 ) | ( wire33546 ) ;
 assign wire33550 = ( wire33528  &  wire33538 ) | ( wire33529  &  wire33538 ) | ( wire33528  &  wire33539 ) | ( wire33529  &  wire33539 ) ;
 assign wire33551 = ( wire33528  &  wire33538 ) | ( wire33529  &  wire33538 ) | ( wire33528  &  wire33539 ) | ( wire33529  &  wire33539 ) ;
 assign wire33557 = ( (~ ng2261)  &  (~ ng2264)  &  (~ ng2267) ) | ( (~ ng2261)  &  (~ ng823)  &  (~ ng2267) ) ;
 assign wire33560 = ( wire3046 ) | ( wire7528 ) | ( wire33557 ) ;
 assign wire33561 = ( wire7531 ) | ( wire7532 ) | ( wire7533 ) | ( wire7534 ) ;
 assign wire33563 = ( (~ wire33438)  &  (~ wire33439)  &  (~ wire33448)  &  (~ wire33449) ) ;
 assign wire33564 = ( (~ wire33458)  &  (~ wire33459)  &  wire33468 ) | ( (~ wire33458)  &  (~ wire33459)  &  wire33469 ) ;
 assign wire33565 = ( wire33478  &  (~ wire33488)  &  (~ wire33489) ) | ( wire33479  &  (~ wire33488)  &  (~ wire33489) ) ;
 assign wire33566 = ( wire33498  &  (~ wire33508)  &  (~ wire33509) ) | ( wire33499  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign wire33569 = ( (~ wire33548)  &  (~ wire33549)  &  wire33550  &  wire33566 ) ;
 assign wire33570 = ( ng13022  &  wire33563  &  wire33564  &  wire33565 ) ;
 assign wire33572 = ( wire33438  &  wire33448 ) | ( wire33439  &  wire33448 ) | ( wire33438  &  wire33449 ) | ( wire33439  &  wire33449 ) ;
 assign wire33573 = ( wire33458  &  wire33468 ) | ( wire33459  &  wire33468 ) | ( wire33458  &  wire33469 ) | ( wire33459  &  wire33469 ) ;
 assign wire33574 = ( wire33478  &  wire33488 ) | ( wire33479  &  wire33488 ) | ( wire33478  &  wire33489 ) | ( wire33479  &  wire33489 ) ;
 assign wire33575 = ( wire33498  &  wire33508 ) | ( wire33499  &  wire33508 ) | ( wire33498  &  wire33509 ) | ( wire33499  &  wire33509 ) ;
 assign wire33576 = ( wire33518  &  wire33560 ) | ( wire33519  &  wire33560 ) | ( wire33518  &  wire33561 ) | ( wire33519  &  wire33561 ) ;
 assign wire33578 = ( wire33575  &  wire33574 ) ;
 assign wire33579 = ( wire33572  &  wire33573  &  wire33576 ) ;
 assign wire33585 = ( ng2245  &  ng2246  &  ng2244 ) | ( ng2246  &  ng2244  &  (~ ng826) ) ;
 assign wire33586 = ( ng2245  &  ng2244  &  (~ ng823) ) | ( ng2244  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33588 = ( wire3046 ) | ( wire7409 ) | ( wire33585 ) ;
 assign wire33589 = ( wire7414 ) | ( wire7415 ) | ( wire33586 ) ;
 assign wire33590 = ( ng2234  &  ng2232 ) ;
 assign wire33591 = ( (~ ng826)  &  ng2200 ) | ( ng2233  &  ng2200 ) ;
 assign wire33592 = ( ng2228  &  ng2226 ) ;
 assign wire33593 = ( (~ ng826)  &  ng2190 ) | ( ng2227  &  ng2190 ) ;
 assign wire33617 = ( ng2231  &  ng2230  &  ng2229 ) | ( ng2231  &  (~ ng826)  &  ng2229 ) ;
 assign wire33618 = ( ng2230  &  ng2229  &  (~ ng823) ) | ( (~ ng826)  &  ng2229  &  (~ ng823) ) ;
 assign wire33621 = ( wire7480 ) | ( wire7481 ) | ( wire33618 ) ;
 assign wire33627 = ( ng2247  &  ng2248  &  ng2249 ) | ( ng2247  &  (~ ng826)  &  ng2249 ) ;
 assign wire33628 = ( ng2247  &  ng2248  &  (~ ng823) ) | ( ng2247  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33630 = ( wire3046 ) | ( wire7467 ) | ( wire33627 ) ;
 assign wire33631 = ( wire7472 ) | ( wire7473 ) | ( wire33628 ) ;
 assign wire33637 = ( ng2239  &  ng2240  &  ng2238 ) | ( ng2240  &  ng2238  &  (~ ng826) ) ;
 assign wire33638 = ( ng2239  &  ng2238  &  (~ ng823) ) | ( ng2238  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33640 = ( wire3046 ) | ( wire7459 ) | ( wire33637 ) ;
 assign wire33641 = ( wire7464 ) | ( wire7465 ) | ( wire33638 ) ;
 assign wire33647 = ( ng2237  &  ng2235  &  ng2236 ) | ( ng2235  &  (~ ng823)  &  ng2236 ) ;
 assign wire33648 = ( ng2237  &  ng2235  &  (~ ng826) ) | ( ng2235  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33651 = ( wire7488 ) | ( wire7489 ) | ( wire33648 ) ;
 assign wire33660 = ( wire33590  &  wire33591 ) | ( wire33592  &  wire33593 ) ;
 assign wire33661 = ( wire7452 ) | ( wire7451 ) ;
 assign wire33662 = ( wire7435 ) | ( wire7436 ) | ( wire7437 ) | ( wire7438 ) ;
 assign wire33663 = ( wire7439 ) | ( wire7440 ) | ( wire7441 ) | ( wire7442 ) ;
 assign wire33664 = ( wire7443 ) | ( wire7444 ) | ( wire7445 ) | ( wire7446 ) ;
 assign wire33665 = ( wire7447 ) | ( wire7448 ) | ( wire7449 ) | ( wire7450 ) ;
 assign wire33668 = ( wire33665 ) | ( wire33664 ) ;
 assign wire33669 = ( wire33660 ) | ( wire33661 ) | ( wire33662 ) | ( wire33663 ) ;
 assign wire33674 = ( wire7455 ) | ( wire33668 ) | ( ng2195  &  ng11916 ) | ( (~ ng2195)  &  (~ ng11916) ) ;
 assign wire33675 = ( wire7456 ) | ( wire33669 ) | ( (~ ng11917)  &  ng12000 ) | ( ng11917  &  (~ ng12000) ) ;
 assign wire33676 = ( ng2223  &  ng2225 ) ;
 assign wire33677 = ( (~ ng826)  &  ng2185 ) | ( ng2224  &  ng2185 ) ;
 assign wire33678 = ( ng2220  &  ng2222 ) ;
 assign wire33679 = ( ng2221  &  ng2180 ) | ( (~ ng826)  &  ng2180 ) ;
 assign wire33703 = ( ng2205  &  ng2207  &  ng2206 ) | ( ng2205  &  ng2207  &  (~ ng826) ) ;
 assign wire33704 = ( ng2205  &  ng2206  &  (~ ng823) ) | ( ng2205  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33706 = ( wire3046 ) | ( wire7491 ) | ( wire33703 ) ;
 assign wire33707 = ( wire7496 ) | ( wire7497 ) | ( wire33704 ) ;
 assign wire33713 = ( ng2217  &  (~ ng826)  &  ng2219 ) | ( ng2217  &  ng2218  &  ng2219 ) ;
 assign wire33714 = ( ng2217  &  (~ ng826)  &  (~ ng823) ) | ( ng2217  &  (~ ng823)  &  ng2218 ) ;
 assign wire33716 = ( wire3046 ) | ( wire7425 ) | ( wire33713 ) ;
 assign wire33717 = ( wire7430 ) | ( wire7431 ) | ( wire33714 ) ;
 assign wire33723 = ( ng2209  &  (~ ng853)  &  ng2210 ) | ( ng2209  &  ng2210  &  ng2208 ) ;
 assign wire33724 = ( ng2209  &  (~ ng823)  &  ng2208 ) | ( (~ ng826)  &  (~ ng823)  &  ng2208 ) ;
 assign wire33726 = ( wire3046 ) | ( wire7417 ) | ( wire33723 ) ;
 assign wire33727 = ( wire7422 ) | ( wire7423 ) | ( wire33724 ) ;
 assign wire33736 = ( wire33676  &  wire33677 ) | ( wire33678  &  wire33679 ) ;
 assign wire33737 = ( wire7400 ) | ( wire7399 ) ;
 assign wire33738 = ( wire7383 ) | ( wire7384 ) | ( wire7385 ) | ( wire7386 ) ;
 assign wire33739 = ( wire7387 ) | ( wire7388 ) | ( wire7389 ) | ( wire7390 ) ;
 assign wire33740 = ( wire7391 ) | ( wire7392 ) | ( wire7393 ) | ( wire7394 ) ;
 assign wire33741 = ( wire7395 ) | ( wire7396 ) | ( wire7397 ) | ( wire7398 ) ;
 assign wire33744 = ( wire33741 ) | ( wire33740 ) ;
 assign wire33745 = ( wire33736 ) | ( wire33737 ) | ( wire33738 ) | ( wire33739 ) ;
 assign wire33747 = ( ng2165  &  wire33706 ) | ( ng2165  &  wire33707 ) | ( (~ ng2165)  &  (~ wire33706)  &  (~ wire33707) ) ;
 assign wire33749 = ( ng2170  &  wire33726 ) | ( ng2170  &  wire33727 ) | ( (~ ng2170)  &  (~ wire33726)  &  (~ wire33727) ) ;
 assign wire33751 = ( wire33747 ) | ( ng2175  &  wire33716 ) | ( ng2175  &  wire33717 ) | ( (~ ng2175)  &  (~ wire33716)  &  (~ wire33717) ) ;
 assign wire33752 = ( wire3369 ) | ( wire33744 ) | ( wire33745 ) | ( wire33749 ) ;
 assign wire33754 = ( ng853  &  (~ ng2477) ) ;
 assign wire33755 = ( ng826  &  (~ ng2478) ) ;
 assign wire33756 = ( ng823  &  (~ ng2479) ) ;
 assign wire33766 = ( wire3369 ) | ( (~ ng18578)  &  wire3055  &  wire3105 ) ;
 assign wire33769 = ( (~ ng18395)  &  (~ ng18478)  &  (~ ng18578) ) | ( (~ ng18395)  &  (~ ng18478)  &  wire3055 ) | ( (~ ng18395)  &  (~ ng18578)  &  wire3055 ) | ( (~ ng18478)  &  (~ ng18578)  &  wire3055 ) ;
 assign wire33770 = ( wire3105  &  wire3327 ) | ( (~ ng18395)  &  (~ ng18478)  &  wire3327 ) ;
 assign wire33771 = ( wire7364 ) | ( wire7365 ) | ( wire33766 ) ;
 assign wire33772 = ( wire7359 ) | ( wire7366 ) | ( wire33769 ) ;
 assign wire33782 = ( wire3369 ) | ( (~ ng18053)  &  (~ ng18231)  &  wire3066 ) ;
 assign wire33785 = ( (~ ng18319)  &  (~ ng18606)  &  (~ ng18053) ) | ( (~ ng18319)  &  (~ ng18606)  &  (~ ng18231) ) | ( (~ ng18319)  &  (~ ng18053)  &  (~ ng18231) ) | ( (~ ng18606)  &  (~ ng18053)  &  (~ ng18231) ) ;
 assign wire33786 = ( wire3066  &  wire3289 ) | ( (~ ng18319)  &  (~ ng18606)  &  wire3289 ) ;
 assign wire33787 = ( wire7342 ) | ( wire7343 ) | ( wire33782 ) ;
 assign wire33788 = ( wire7337 ) | ( wire7344 ) | ( wire33785 ) ;
 assign wire33790 = ( wire33528  &  (~ wire33538)  &  (~ wire33539) ) | ( wire33529  &  (~ wire33538)  &  (~ wire33539) ) ;
 assign wire33791 = ( (~ ng22400)  &  wire33790 ) ;
 assign wire33792 = ( (~ wire33528)  &  (~ wire33529)  &  (~ wire33538)  &  (~ wire33539) ) ;
 assign wire33793 = ( (~ ng2397)  &  ng826 ) | ( (~ ng2396)  &  ng853 ) ;
 assign wire33794 = ( wire7331  &  wire33548 ) | ( wire7331  &  wire33549 ) | ( wire33548  &  wire33793 ) | ( wire33549  &  wire33793 ) ;
 assign wire33795 = ( ng24723 ) | ( wire3925  &  (~ wire33538)  &  (~ wire33539) ) ;
 assign wire33799 = ( (~ ng28584)  &  (~ ng25969)  &  wire33508 ) | ( (~ ng28584)  &  (~ ng25969)  &  wire33509 ) | ( (~ ng28584)  &  ng25969  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign wire33800 = ( ng2170  &  ng27756 ) | ( ng25874  &  (~ ng27756)  &  (~ ng16693) ) ;
 assign wire33805 = ( ng11678  &  (~ wire33488)  &  (~ wire33489) ) | ( (~ ng11678)  &  wire33488  &  wire33550 ) | ( (~ ng11678)  &  wire33489  &  wire33550 ) | ( (~ wire33488)  &  (~ wire33489)  &  (~ wire33550) ) ;
 assign wire33807 = ( (~ ng12959)  &  ng13022 ) | ( (~ ng13022)  &  ng11678 ) | ( (~ ng13022)  &  (~ wire33550) ) | ( ng12959  &  (~ ng11678)  &  wire33550 ) ;
 assign wire33808 = ( (~ ng11678)  &  (~ wire33518)  &  (~ wire33519)  &  wire33550 ) ;
 assign wire33809 = ( ng27585  &  (~ wire33805)  &  wire33808 ) ;
 assign wire33811 = ( (~ wire33468)  &  (~ wire33469)  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire33812 = ( (~ ng27585)  &  (~ wire33468)  &  (~ wire33469) ) | ( (~ wire33468)  &  (~ wire33469)  &  wire33805 ) ;
 assign wire33813 = ( (~ ng11678)  &  (~ wire33468)  &  (~ wire33469)  &  wire33550 ) ;
 assign wire33814 = ( ng13022  &  (~ ng28584)  &  (~ ng26941) ) | ( (~ ng28584)  &  ng26941  &  wire33809 ) ;
 assign wire33815 = ( (~ ng28584)  &  ng26941  &  wire33811 ) | ( (~ ng28584)  &  ng26941  &  wire33812 ) ;
 assign wire33819 = ( (~ ng12978)  &  ng12836 ) | ( (~ ng12836)  &  ng11678 ) | ( (~ ng12836)  &  (~ wire33550) ) | ( ng12978  &  (~ ng11678)  &  wire33550 ) ;
 assign wire33823 = ( (~ ng28584)  &  (~ wire3426)  &  wire33438 ) | ( (~ ng28584)  &  (~ wire3426)  &  wire33439 ) | ( (~ ng28584)  &  wire3426  &  (~ wire33438)  &  (~ wire33439) ) ;
 assign wire33824 = ( ng27756  &  (~ ng11882) ) | ( ng25874  &  (~ ng27756)  &  (~ ng16693) ) ;
 assign wire33827 = ( ng2160  &  ng2147  &  ng2156  &  ng2151 ) ;
 assign wire33829 = ( ng2129  &  ng2133  &  ng2138 ) ;
 assign wire33837 = ( ng2418  &  ng2421  &  ng2429 ) | ( ng2418  &  ng2421  &  (~ ng826) ) ;
 assign wire33838 = ( ng2421  &  ng2429  &  (~ ng823) ) | ( ng2421  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33840 = ( wire3046 ) | ( wire7262 ) | ( wire33837 ) ;
 assign wire33841 = ( wire7267 ) | ( wire7268 ) | ( wire33838 ) ;
 assign wire33847 = ( ng2448  &  ng2459  &  ng2451 ) | ( ng2459  &  ng2451  &  (~ ng823) ) ;
 assign wire33850 = ( wire3046 ) | ( wire7270 ) | ( wire33847 ) ;
 assign wire33851 = ( wire7273 ) | ( wire7274 ) | ( wire7275 ) | ( wire7276 ) ;
 assign wire33857 = ( ng2436  &  ng2444  &  ng2433 ) | ( ng2436  &  ng2433  &  (~ ng826) ) ;
 assign wire33858 = ( ng2436  &  ng2444  &  (~ ng823) ) | ( ng2436  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33860 = ( wire3046 ) | ( wire7278 ) | ( wire33857 ) ;
 assign wire33861 = ( wire7283 ) | ( wire7284 ) | ( wire33858 ) ;
 assign wire33862 = ( (~ wire33528)  &  (~ wire33529)  &  wire33538 ) | ( (~ wire33528)  &  (~ wire33529)  &  wire33539 ) ;
 assign wire33868 = ( (~ ng2495)  &  (~ ng2492)  &  (~ ng2498) ) | ( (~ ng2492)  &  (~ ng823)  &  (~ ng2498) ) ;
 assign wire33871 = ( wire3046 ) | ( wire7246 ) | ( wire33868 ) ;
 assign wire33872 = ( wire7249 ) | ( wire7250 ) | ( wire7251 ) | ( wire7252 ) ;
 assign wire33876 = ( ng2200  &  ng2170  &  ng2175  &  ng2185 ) ;
 assign wire33877 = ( ng2180  &  ng2165  &  ng2190  &  ng2195 ) ;
 assign wire33878 = ( wire33630 ) | ( wire33631 ) | ( (~ wire33876) ) | ( (~ wire33877) ) ;
 assign wire33886 = ( (~ ng2489)  &  (~ ng2486)  &  (~ ng2483) ) | ( (~ ng2489)  &  (~ ng2486)  &  (~ ng826) ) ;
 assign wire33887 = ( (~ ng2489)  &  (~ ng2483)  &  (~ ng823) ) | ( (~ ng2489)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33889 = ( wire3046 ) | ( wire7235 ) | ( wire33886 ) ;
 assign wire33890 = ( wire7240 ) | ( wire7241 ) | ( wire33887 ) ;
 assign wire33892 = ( ng2503  &  (~ ng853)  &  ng2502 ) ;
 assign wire33894 = ( ng2503  &  ng2501  &  ng2502 ) ;
 assign wire33896 = ( ng2501  &  (~ ng823)  &  ng2502 ) ;
 assign wire33898 = ( ng2503  &  ng2501  &  (~ ng826) ) ;
 assign wire33899 = ( ng2501  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33900 = ( (~ ng823)  &  (~ ng853)  &  ng2502 ) ;
 assign wire33901 = ( ng2503  &  (~ ng826)  &  (~ ng853) ) ;
 assign wire33906 = ( wire7227 ) | ( wire7228 ) | ( wire7229 ) | ( wire7230 ) ;
 assign wire33907 = ( wire7231 ) | ( wire7232 ) | ( wire7233 ) | ( wire7234 ) ;
 assign wire33913 = ( (~ ng826)  &  (~ ng2507)  &  (~ ng2510) ) | ( (~ ng2504)  &  (~ ng2507)  &  (~ ng2510) ) ;
 assign wire33914 = ( (~ ng826)  &  (~ ng823)  &  (~ ng2510) ) | ( (~ ng2504)  &  (~ ng823)  &  (~ ng2510) ) ;
 assign wire33917 = ( wire7201 ) | ( wire7202 ) | ( wire33914 ) ;
 assign wire33923 = ( ng2255  &  ng2254  &  ng2253 ) | ( ng2255  &  ng2253  &  (~ ng826) ) ;
 assign wire33924 = ( ng2254  &  ng2253  &  (~ ng823) ) | ( ng2253  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire33926 = ( wire3046 ) | ( wire7204 ) | ( (~ wire33876) ) | ( (~ wire33877) ) ;
 assign wire33927 = ( wire33924 ) | ( wire33923 ) ;
 assign wire33934 = ( (~ ng823)  &  (~ ng2513)  &  (~ ng2519) ) | ( (~ ng2513)  &  (~ ng2516)  &  (~ ng2519) ) ;
 assign wire33935 = ( (~ ng826)  &  (~ ng823)  &  (~ ng2519) ) | ( (~ ng826)  &  (~ ng2516)  &  (~ ng2519) ) ;
 assign wire33937 = ( wire3046 ) | ( wire7213 ) | ( wire33934 ) ;
 assign wire33938 = ( wire7218 ) | ( wire7219 ) | ( wire33935 ) ;
 assign wire33940 = ( ng823  &  (~ ng2524)  &  ng2257 ) ;
 assign wire33941 = ( (~ ng2522)  &  ng853  &  ng2257 ) ;
 assign wire33942 = ( (~ ng2523)  &  ng826  &  ng2257 ) ;
 assign wire33944 = ( ng2257  &  (~ ng12180)  &  ng12121  &  ng18325 ) | ( ng2257  &  ng12180  &  (~ ng12121)  &  (~ ng18325) ) ;
 assign wire33948 = ( ng2257  &  (~ ng12180)  &  (~ ng12121)  &  ng18325 ) | ( ng2257  &  ng12180  &  ng12121  &  (~ ng18325) ) ;
 assign wire33954 = ( (~ ng1309)  &  (~ ng2691)  &  (~ ng2694) ) | ( (~ ng2691)  &  (~ ng2688)  &  (~ ng2694) ) ;
 assign wire33955 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2688) ) | ( (~ ng1312)  &  (~ ng2688)  &  (~ ng2694) ) ;
 assign wire33957 = ( wire3049 ) | ( wire7170 ) | ( wire33954 ) ;
 assign wire33958 = ( wire7175 ) | ( wire7176 ) | ( wire33955 ) ;
 assign wire33967 = ( wire3049 ) | ( wire7162 ) | ( wire7163 ) | ( wire7164 ) ;
 assign wire33968 = ( wire7165 ) | ( wire7166 ) | ( wire7167 ) | ( wire7168 ) ;
 assign wire33974 = ( (~ ng1312)  &  (~ ng2679)  &  (~ ng2685) ) | ( (~ ng2679)  &  (~ ng2685)  &  (~ ng2682) ) ;
 assign wire33975 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2679) ) | ( (~ ng1315)  &  (~ ng2679)  &  (~ ng2682) ) ;
 assign wire33977 = ( wire3049 ) | ( wire7154 ) | ( wire33974 ) ;
 assign wire33978 = ( wire7159 ) | ( wire7160 ) | ( wire33975 ) ;
 assign wire33986 = ( (~ ng1312)  &  (~ ng1315)  &  ng2659 ) | ( (~ ng1315)  &  ng2659  &  ng2660 ) ;
 assign wire33988 = ( wire3049 ) | ( wire7143 ) | ( wire7144 ) | ( wire7145 ) ;
 assign wire33989 = ( wire7148 ) | ( wire7149 ) | ( wire33986 ) ;
 assign wire33995 = ( ng2649  &  ng2651  &  ng2650 ) | ( ng2649  &  (~ ng1312)  &  ng2650 ) ;
 assign wire33998 = ( wire3049 ) | ( wire7135 ) | ( wire33995 ) ;
 assign wire33999 = ( wire7138 ) | ( wire7139 ) | ( wire7140 ) | ( wire7141 ) ;
 assign wire34006 = ( (~ ng1312)  &  (~ ng1315)  &  ng2656 ) | ( (~ ng1315)  &  ng2656  &  ng2657 ) ;
 assign wire34008 = ( wire3049 ) | ( wire7127 ) | ( wire7128 ) | ( wire7129 ) ;
 assign wire34009 = ( wire7132 ) | ( wire7133 ) | ( wire34006 ) ;
 assign wire34016 = ( (~ ng1312)  &  (~ ng1315)  &  ng2653 ) | ( (~ ng1315)  &  ng2654  &  ng2653 ) ;
 assign wire34018 = ( wire3049 ) | ( wire7119 ) | ( wire7120 ) | ( wire7121 ) ;
 assign wire34019 = ( wire7124 ) | ( wire7125 ) | ( wire34016 ) ;
 assign wire34020 = ( wire33988  &  (~ wire33998)  &  (~ wire33999) ) | ( wire33989  &  (~ wire33998)  &  (~ wire33999) ) ;
 assign wire34024 = ( pg3229  &  (~ ng12231)  &  (~ ng12305) ) | ( (~ pg3229)  &  ng12305  &  (~ ng12269) ) ;
 assign wire34028 = ( pg563 ) | ( ng559 ) | ( ng1309  &  (~ ng499) ) ;
 assign wire34034 = ( ng738  &  (~ ng1312)  &  ng737 ) | ( ng738  &  ng739  &  ng737 ) ;
 assign wire34035 = ( ng738  &  (~ ng1312)  &  (~ ng1315) ) | ( ng738  &  (~ ng1315)  &  ng739 ) ;
 assign wire34037 = ( wire3049 ) | ( wire7078 ) | ( wire34034 ) ;
 assign wire34038 = ( wire7083 ) | ( wire7084 ) | ( wire34035 ) ;
 assign wire34040 = ( wire31723 ) | ( wire31724 ) | ( (~ wire31711)  &  (~ wire31712) ) ;
 assign wire34041 = ( wire31687 ) | ( wire31688 ) | ( (~ wire31699)  &  (~ wire31700) ) ;
 assign wire34042 = ( wire31663 ) | ( wire31664 ) | ( wire31675 ) | ( wire31676 ) ;
 assign wire34043 = ( wire31651 ) | ( wire31652 ) | ( (~ wire31639)  &  (~ wire31640) ) ;
 assign wire34044 = ( (~ wire31605)  &  (~ wire31606) ) | ( (~ wire31627)  &  (~ wire31628) ) ;
 assign wire34045 = ( wire31615 ) | ( wire31616 ) | ( wire34037 ) | ( wire34038 ) ;
 assign wire34048 = ( wire34045 ) | ( wire34044 ) ;
 assign wire34049 = ( wire34040 ) | ( wire34041 ) | ( wire34042 ) | ( wire34043 ) ;
 assign wire34051 = ( ng736  &  (~ ng1315)  &  ng735 ) ;
 assign wire34052 = ( ng557  &  (~ ng510)  &  wire34051 ) ;
 assign wire34054 = ( ng734  &  (~ ng1312)  &  ng735 ) ;
 assign wire34055 = ( ng557  &  (~ ng510)  &  wire34054 ) ;
 assign wire34057 = ( ng736  &  ng734  &  ng735 ) ;
 assign wire34058 = ( ng557  &  (~ ng510)  &  wire34057 ) ;
 assign wire34060 = ( ng736  &  ng734  &  (~ ng1309) ) ;
 assign wire34061 = ( ng557  &  (~ ng510)  &  wire34060 ) ;
 assign wire34062 = ( (~ ng1312)  &  (~ ng1315)  &  ng735 ) ;
 assign wire34063 = ( ng557  &  (~ ng510)  &  wire34062 ) ;
 assign wire34064 = ( ng734  &  (~ ng1312)  &  (~ ng1309) ) ;
 assign wire34065 = ( ng557  &  (~ ng510)  &  wire34064 ) ;
 assign wire34066 = ( ng736  &  (~ ng1315)  &  (~ ng1309) ) ;
 assign wire34067 = ( ng557  &  (~ ng510)  &  wire34066 ) ;
 assign wire34068 = ( ng557  &  (~ ng510)  &  wire3049 ) ;
 assign wire34069 = ( wire7070 ) | ( wire34048  &  wire34052 ) | ( wire34049  &  wire34052 ) ;
 assign wire34070 = ( wire34048  &  wire34055 ) | ( wire34049  &  wire34055 ) | ( wire34048  &  wire34058 ) | ( wire34049  &  wire34058 ) ;
 assign wire34071 = ( wire34048  &  wire34061 ) | ( wire34049  &  wire34061 ) | ( wire34048  &  wire34063 ) | ( wire34049  &  wire34063 ) ;
 assign wire34072 = ( wire34048  &  wire34065 ) | ( wire34049  &  wire34065 ) | ( wire34048  &  wire34067 ) | ( wire34049  &  wire34067 ) ;
 assign wire34074 = ( wire34071 ) | ( wire34070 ) ;
 assign wire34075 = ( wire7069 ) | ( wire34069 ) | ( wire34072 ) ;
 assign wire34076 = ( ng12082  &  wire3188 ) | ( wire3188  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire34079 = ( ng3135 ) | ( ng3139 ) | ( ng3120 ) | ( ng3147 ) ;
 assign wire34081 = ( ng3139  &  (~ ng185)  &  ng3147 ) ;
 assign wire34082 = ( (~ ng3139)  &  (~ ng2991)  &  (~ ng2992)  &  ng3147 ) ;
 assign wire34083 = ( ng3135  &  (~ ng3120)  &  (~ ng3147) ) ;
 assign wire34084 = ( (~ pg3233) ) | ( pg3230 ) | ( (~ ng8381)  &  (~ wire34079) ) ;
 assign wire34087 = ( wire7045 ) | ( wire34084 ) | ( (~ ng8381)  &  wire34083 ) ;
 assign wire34088 = ( (~ wire30967)  &  (~ wire30968)  &  (~ wire30977)  &  (~ wire30978) ) ;
 assign wire34089 = ( (~ ng23495)  &  wire34088 ) ;
 assign wire34091 = ( ng2257  &  wire30957 ) | ( ng2257  &  wire30958 ) ;
 assign wire34093 = ( (~ ng23495)  &  wire3237 ) | ( ng11624  &  wire3237  &  wire31271 ) ;
 assign wire34094 = ( (~ wire30967)  &  (~ wire30968)  &  (~ wire30977)  &  (~ wire30978) ) ;
 assign wire34095 = ( wire30957  &  wire30977 ) | ( wire30958  &  wire30977 ) | ( wire30957  &  wire30978 ) | ( wire30958  &  wire30978 ) ;
 assign wire34096 = ( ng11644  &  ng13378  &  ng11624 ) | ( (~ ng11644)  &  (~ ng13378)  &  ng11624  &  wire3936 ) ;
 assign wire34097 = ( wire34096 ) | ( ng11624  &  ng23495  &  wire34091 ) ;
 assign wire34099 = ( wire7029 ) | ( wire7030 ) | ( wire34097 ) ;
 assign wire34100 = ( wire34099 ) | ( ng27834  &  wire34093 ) ;
 assign wire34114 = ( (~ ng565)  &  (~ ng1315)  &  (~ ng567) ) | ( (~ ng565)  &  (~ ng489)  &  (~ ng567) ) ;
 assign wire34115 = ( (~ ng565)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng565)  &  (~ ng1312)  &  (~ ng489) ) ;
 assign wire34117 = ( wire3049 ) | ( wire7006 ) | ( wire34114 ) ;
 assign wire34118 = ( wire7011 ) | ( wire7012 ) | ( wire34115 ) ;
 assign wire34120 = ( (~ ng599)  &  (~ ng596)  &  (~ ng602) ) ;
 assign wire34122 = ( (~ ng1312)  &  (~ ng596)  &  (~ ng602) ) ;
 assign wire34124 = ( (~ ng1309)  &  (~ ng599)  &  (~ ng602) ) ;
 assign wire34134 = ( (~ ng1315)  &  (~ ng599)  &  (~ ng596) ) ;
 assign wire34138 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng596) ) ;
 assign wire34141 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng602) ) ;
 assign wire34144 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng599) ) ;
 assign wire34154 = ( wire6982 ) | ( wire6983 ) | ( wire6984 ) | ( wire6988 ) ;
 assign wire34155 = ( wire6989 ) | ( wire6990 ) | ( wire6991 ) | ( wire6993 ) ;
 assign wire34156 = ( wire6994 ) | ( wire6996 ) | ( wire6997 ) | ( wire6999 ) ;
 assign wire34157 = ( wire7000 ) | ( wire7002 ) | ( wire7003 ) | ( wire7005 ) ;
 assign wire34161 = ( wire34117  &  wire34122 ) | ( wire34118  &  wire34122 ) | ( wire34117  &  wire34124 ) | ( wire34118  &  wire34124 ) ;
 assign wire34162 = ( wire34117  &  wire34134 ) | ( wire34118  &  wire34134 ) | ( wire34117  &  wire34138 ) | ( wire34118  &  wire34138 ) ;
 assign wire34163 = ( wire34117  &  wire34141 ) | ( wire34118  &  wire34141 ) | ( wire34117  &  wire34144 ) | ( wire34118  &  wire34144 ) ;
 assign wire34164 = ( wire3049 ) | ( wire34156 ) | ( wire34157 ) ;
 assign wire34165 = ( wire6985 ) | ( wire34154 ) | ( wire34155 ) | ( wire34161 ) ;
 assign wire34166 = ( wire34163 ) | ( wire34162 ) ;
 assign wire34176 = ( wire3049 ) | ( wire6974 ) | ( wire6975 ) | ( wire6976 ) ;
 assign wire34177 = ( wire6977 ) | ( wire6978 ) | ( wire6979 ) | ( wire6980 ) ;
 assign wire34183 = ( (~ ng381)  &  (~ ng1315)  &  (~ ng379) ) | ( (~ ng381)  &  (~ ng383)  &  (~ ng379) ) ;
 assign wire34186 = ( wire3049 ) | ( wire6966 ) | ( wire34183 ) ;
 assign wire34187 = ( wire6969 ) | ( wire6970 ) | ( wire6971 ) | ( wire6972 ) ;
 assign wire34194 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng349) ) | ( (~ ng1312)  &  (~ ng349)  &  (~ ng353) ) ;
 assign wire34196 = ( wire3049 ) | ( wire6950 ) | ( wire6951 ) | ( wire6952 ) ;
 assign wire34197 = ( wire6955 ) | ( wire6956 ) | ( wire34194 ) ;
 assign wire34198 = ( wire31482  &  (~ wire31492)  &  (~ wire31493) ) | ( wire31483  &  (~ wire31492)  &  (~ wire31493) ) ;
 assign wire34199 = ( wire34176  &  (~ wire34186)  &  (~ wire34187) ) | ( wire34177  &  (~ wire34186)  &  (~ wire34187) ) ;
 assign wire34201 = ( wire31492  &  (~ wire34176)  &  (~ wire34177) ) | ( wire31493  &  (~ wire34176)  &  (~ wire34177) ) ;
 assign wire34202 = ( wire31512  &  (~ wire34186)  &  (~ wire34187) ) | ( wire31513  &  (~ wire34186)  &  (~ wire34187) ) ;
 assign wire34204 = ( wire31502  &  (~ wire34176)  &  (~ wire34177) ) | ( wire31503  &  (~ wire34176)  &  (~ wire34177) ) ;
 assign wire34205 = ( wire31512  &  wire34186 ) | ( wire31513  &  wire34186 ) | ( wire31512  &  wire34187 ) | ( wire31513  &  wire34187 ) ;
 assign wire34213 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng394) ) | ( (~ ng1312)  &  (~ ng324)  &  (~ ng394) ) ;
 assign wire34215 = ( wire3049 ) | ( wire6958 ) | ( wire6959 ) | ( wire6960 ) ;
 assign wire34216 = ( wire6963 ) | ( wire6964 ) | ( wire34213 ) ;
 assign wire34217 = ( wire31502  &  (~ wire31512)  &  (~ wire31513) ) | ( wire31503  &  (~ wire31512)  &  (~ wire31513) ) ;
 assign wire34219 = ( (~ wire31502)  &  (~ wire31503)  &  (~ wire34176)  &  (~ wire34177) ) ;
 assign wire34221 = ( wire31502  &  wire31512 ) | ( wire31503  &  wire31512 ) | ( wire31502  &  wire31513 ) | ( wire31503  &  wire31513 ) ;
 assign wire34223 = ( (~ wire34176)  &  (~ wire34177)  &  (~ wire34186)  &  (~ wire34187) ) ;
 assign wire34225 = ( (~ wire31482)  &  (~ wire31483)  &  (~ wire34176)  &  (~ wire34177) ) ;
 assign wire34226 = ( (~ wire34186)  &  (~ wire34187)  &  (~ wire34196)  &  (~ wire34197) ) ;
 assign wire34227 = ( wire31502  &  wire34176 ) | ( wire31503  &  wire34176 ) | ( wire31502  &  wire34177 ) | ( wire31503  &  wire34177 ) ;
 assign wire34228 = ( (~ wire31512)  &  (~ wire31513)  &  wire34196 ) | ( (~ wire31512)  &  (~ wire31513)  &  wire34197 ) ;
 assign wire34229 = ( (~ wire31492)  &  (~ wire31493)  &  wire31502 ) | ( (~ wire31492)  &  (~ wire31493)  &  wire31503 ) ;
 assign wire34230 = ( wire31512  &  wire34215 ) | ( wire31513  &  wire34215 ) | ( wire31512  &  wire34216 ) | ( wire31513  &  wire34216 ) ;
 assign wire34231 = ( wire31492  &  wire34176 ) | ( wire31493  &  wire34176 ) | ( wire31492  &  wire34177 ) | ( wire31493  &  wire34177 ) ;
 assign wire34232 = ( (~ wire31512)  &  (~ wire31513)  &  (~ wire34186)  &  (~ wire34187) ) ;
 assign wire34235 = ( (~ wire31512)  &  (~ wire31513)  &  wire34186 ) | ( (~ wire31512)  &  (~ wire31513)  &  wire34187 ) ;
 assign wire34236 = ( (~ wire31502)  &  (~ wire31503)  &  wire34176 ) | ( (~ wire31502)  &  (~ wire31503)  &  wire34177 ) ;
 assign wire34237 = ( wire34225  &  wire34226 ) | ( wire34227  &  wire34228 ) ;
 assign wire34238 = ( wire34229  &  wire34230 ) | ( wire34231  &  wire34232 ) ;
 assign wire34239 = ( (~ ng12033)  &  ng10784  &  wire34235 ) | ( ng12033  &  (~ ng10784)  &  wire34236 ) ;
 assign wire34243 = ( wire6940 ) | ( wire6941 ) | ( wire34239 ) ;
 assign wire34244 = ( wire6946 ) | ( wire6947 ) | ( wire34237 ) | ( wire34238 ) ;
 assign wire34245 = ( (~ wire31512)  &  (~ wire31513)  &  wire34186 ) | ( (~ wire31512)  &  (~ wire31513)  &  wire34187 ) ;
 assign wire34247 = ( (~ wire31492)  &  (~ wire31493)  &  (~ wire31502)  &  (~ wire31503) ) ;
 assign wire34249 = ( (~ wire31482)  &  (~ wire31483)  &  (~ wire34215)  &  (~ wire34216) ) ;
 assign wire34250 = ( wire31512  &  wire34176 ) | ( wire31513  &  wire34176 ) | ( wire31512  &  wire34177 ) | ( wire31513  &  wire34177 ) ;
 assign wire34251 = ( wire31482  &  wire34215 ) | ( wire31483  &  wire34215 ) | ( wire31482  &  wire34216 ) | ( wire31483  &  wire34216 ) ;
 assign wire34252 = ( (~ wire31482)  &  (~ wire31483)  &  wire34186 ) | ( (~ wire31482)  &  (~ wire31483)  &  wire34187 ) ;
 assign wire34253 = ( wire31492  &  (~ wire31502)  &  (~ wire31503) ) | ( wire31493  &  (~ wire31502)  &  (~ wire31503) ) ;
 assign wire34254 = ( wire3345  &  wire34249 ) | ( wire3345  &  wire34250 ) ;
 assign wire34255 = ( ng10784  &  wire34252 ) | ( ng12033  &  (~ ng10784)  &  wire34251 ) ;
 assign wire34260 = ( wire6928 ) | ( wire6929 ) | ( wire6930 ) | ( wire6939 ) ;
 assign wire34261 = ( wire6931 ) | ( wire6932 ) | ( wire34254 ) | ( wire34255 ) ;
 assign wire34262 = ( wire34261 ) | ( wire34260 ) ;
 assign wire34264 = ( ng13055  &  wire34164 ) | ( ng13055  &  wire34165 ) | ( ng13055  &  wire34166 ) ;
 assign wire34265 = ( (~ wire31587)  &  (~ wire31588)  &  (~ wire31589)  &  wire34264 ) ;
 assign wire34266 = ( ng13055  &  wire31587 ) | ( ng13055  &  wire31588 ) | ( ng13055  &  wire31589 ) ;
 assign wire34267 = ( wire34243  &  wire34266 ) | ( wire34244  &  wire34266 ) ;
 assign wire34269 = ( (~ ng660)  &  (~ ng1312) ) | ( (~ ng660)  &  (~ ng630) ) ;
 assign wire34270 = ( ng660  &  (~ ng1312) ) | ( ng660  &  (~ ng630) ) ;
 assign wire34273 = ( (~ ng28529)  &  ng26327  &  wire31837 ) | ( (~ ng28529)  &  ng26327  &  wire31838 ) | ( (~ ng28529)  &  (~ ng26327)  &  (~ wire31837)  &  (~ wire31838) ) ;
 assign wire34274 = ( ng793  &  ng27743 ) | ( (~ ng16655)  &  ng25818  &  (~ ng27743) ) ;
 assign wire34281 = ( (~ ng17031)  &  ng753 ) ;
 assign wire34283 = ( (~ ng17031)  &  ng749 ) ;
 assign wire34284 = ( ng1115  &  (~ ng823) ) | ( ng1115  &  (~ wire32243)  &  (~ wire32244) ) ;
 assign wire34289 = ( (~ ng805)  &  wire3056  &  wire31887 ) | ( (~ ng805)  &  wire3056  &  wire31888 ) | ( ng805  &  wire3056  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign wire34290 = ( (~ ng18363)  &  (~ ng18441)  &  (~ ng18195)  &  (~ ng18290) ) ;
 assign wire34291 = ( wire3067  &  (~ ng18096)  &  (~ ng17998)  &  (~ ng18492) ) ;
 assign wire34293 = ( (~ ng23511)  &  (~ wire32128) ) | ( (~ ng23511)  &  (~ wire31815)  &  (~ wire31816) ) ;
 assign wire34294 = ( wire6875 ) | ( ng1008  &  (~ ng853) ) ;
 assign wire34295 = ( wire34294 ) | ( (~ ng13165)  &  ng17086  &  (~ ng27850) ) ;
 assign wire34296 = ( (~ ng771)  &  (~ wire31837)  &  (~ wire31838) ) ;
 assign wire34297 = ( (~ ng771)  &  (~ wire31837)  &  (~ wire31838) ) ;
 assign wire34298 = ( ng771  &  wire31837 ) | ( ng771  &  wire31838 ) ;
 assign wire34299 = ( ng771  &  wire31837 ) | ( ng771  &  wire31838 ) ;
 assign wire34300 = ( (~ ng744)  &  (~ wire31907)  &  (~ wire31908) ) ;
 assign wire34301 = ( (~ ng744)  &  (~ wire31907)  &  (~ wire31908) ) ;
 assign wire34302 = ( ng744  &  wire31907 ) | ( ng744  &  wire31908 ) ;
 assign wire34303 = ( ng744  &  wire31907 ) | ( ng744  &  wire31908 ) ;
 assign wire34304 = ( (~ ng767)  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign wire34305 = ( (~ ng767)  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign wire34306 = ( ng767  &  wire31897 ) | ( ng767  &  wire31898 ) ;
 assign wire34307 = ( ng767  &  wire31897 ) | ( ng767  &  wire31898 ) ;
 assign wire34308 = ( (~ ng753)  &  (~ wire31857)  &  (~ wire31858) ) ;
 assign wire34309 = ( (~ ng753)  &  (~ wire31857)  &  (~ wire31858) ) ;
 assign wire34310 = ( ng753  &  wire31857 ) | ( ng753  &  wire31858 ) ;
 assign wire34311 = ( ng753  &  wire31857 ) | ( ng753  &  wire31858 ) ;
 assign wire34312 = ( (~ ng740)  &  (~ wire31867)  &  (~ wire31868) ) ;
 assign wire34313 = ( (~ ng740)  &  (~ wire31867)  &  (~ wire31868) ) ;
 assign wire34314 = ( ng740  &  wire31867 ) | ( ng740  &  wire31868 ) ;
 assign wire34315 = ( ng740  &  wire31867 ) | ( ng740  &  wire31868 ) ;
 assign wire34316 = ( (~ ng776)  &  (~ wire31785)  &  (~ wire31786) ) ;
 assign wire34317 = ( (~ ng776)  &  (~ wire31785)  &  (~ wire31786) ) ;
 assign wire34318 = ( ng776  &  wire31785 ) | ( ng776  &  wire31786 ) ;
 assign wire34319 = ( ng776  &  wire31785 ) | ( ng776  &  wire31786 ) ;
 assign wire34320 = ( (~ ng780)  &  (~ wire31826)  &  (~ wire31827) ) ;
 assign wire34321 = ( (~ ng780)  &  (~ wire31826)  &  (~ wire31827) ) ;
 assign wire34322 = ( ng780  &  wire31826 ) | ( ng780  &  wire31827 ) ;
 assign wire34323 = ( ng780  &  wire31826 ) | ( ng780  &  wire31827 ) ;
 assign wire34324 = ( (~ ng758)  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign wire34325 = ( (~ ng758)  &  (~ wire31887)  &  (~ wire31888) ) ;
 assign wire34326 = ( ng758  &  wire31887 ) | ( ng758  &  wire31888 ) ;
 assign wire34327 = ( ng758  &  wire31887 ) | ( ng758  &  wire31888 ) ;
 assign wire34328 = ( (~ ng762)  &  (~ wire31847)  &  (~ wire31848) ) ;
 assign wire34329 = ( ng762  &  wire31847 ) | ( ng762  &  wire31848 ) ;
 assign wire34330 = ( (~ ng749)  &  (~ wire31877)  &  (~ wire31878) ) ;
 assign wire34331 = ( ng749  &  wire31877 ) | ( ng749  &  wire31878 ) ;
 assign wire34332 = ( (~ ng762)  &  (~ wire31847)  &  (~ wire31848) ) ;
 assign wire34333 = ( ng762  &  wire31847 ) | ( ng762  &  wire31848 ) ;
 assign wire34334 = ( (~ ng749)  &  (~ wire31877)  &  (~ wire31878) ) ;
 assign wire34335 = ( ng749  &  wire31877 ) | ( ng749  &  wire31878 ) ;
 assign wire34336 = ( (~ ng11663)  &  wire34296 ) | ( (~ ng11600)  &  wire34296 ) | ( (~ ng11647)  &  wire34296 ) | ( (~ ng11663)  &  ng11600  &  (~ ng11647) ) ;
 assign wire34337 = ( (~ ng11647)  &  wire34298 ) | ( (~ wire31828)  &  wire34298 ) | ( (~ ng11647)  &  wire34300 ) | ( (~ wire31828)  &  wire34300 ) ;
 assign wire34338 = ( (~ ng11647)  &  wire34302 ) | ( (~ wire31828)  &  wire34302 ) | ( (~ ng11647)  &  wire34304 ) | ( (~ wire31828)  &  wire34304 ) ;
 assign wire34339 = ( (~ ng11647)  &  wire34306 ) | ( (~ wire31828)  &  wire34306 ) | ( (~ ng11647)  &  wire34308 ) | ( (~ wire31828)  &  wire34308 ) ;
 assign wire34340 = ( (~ ng11647)  &  wire34310 ) | ( (~ wire31828)  &  wire34310 ) | ( (~ ng11647)  &  wire34312 ) | ( (~ wire31828)  &  wire34312 ) ;
 assign wire34341 = ( (~ ng11647)  &  wire34314 ) | ( (~ wire31828)  &  wire34314 ) | ( (~ ng11647)  &  wire34316 ) | ( (~ wire31828)  &  wire34316 ) ;
 assign wire34342 = ( (~ ng11647)  &  wire34318 ) | ( (~ wire31828)  &  wire34318 ) | ( (~ ng11647)  &  wire34320 ) | ( (~ wire31828)  &  wire34320 ) ;
 assign wire34343 = ( (~ ng11647)  &  wire34322 ) | ( (~ wire31828)  &  wire34322 ) | ( (~ ng11647)  &  wire34324 ) | ( (~ wire31828)  &  wire34324 ) ;
 assign wire34344 = ( (~ ng11647)  &  wire34326 ) | ( (~ wire31828)  &  wire34326 ) | ( (~ ng11647)  &  wire34328 ) | ( (~ wire31828)  &  wire34328 ) ;
 assign wire34345 = ( (~ ng11647)  &  wire34329 ) | ( (~ wire31828)  &  wire34329 ) | ( (~ ng11647)  &  wire34330 ) | ( (~ wire31828)  &  wire34330 ) ;
 assign wire34346 = ( (~ ng11647)  &  ng10711 ) | ( ng10711  &  (~ wire31828) ) | ( (~ ng11647)  &  wire34331 ) | ( (~ wire31828)  &  wire34331 ) ;
 assign wire34351 = ( wire34345 ) | ( wire34344 ) ;
 assign wire34352 = ( wire34346 ) | ( (~ wire31924)  &  wire34297 ) | ( (~ wire31925)  &  wire34297 ) ;
 assign wire34353 = ( (~ wire31924)  &  wire34299 ) | ( (~ wire31925)  &  wire34299 ) | ( (~ wire31924)  &  wire34301 ) | ( (~ wire31925)  &  wire34301 ) ;
 assign wire34354 = ( (~ wire31924)  &  wire34303 ) | ( (~ wire31925)  &  wire34303 ) | ( (~ wire31924)  &  wire34305 ) | ( (~ wire31925)  &  wire34305 ) ;
 assign wire34355 = ( (~ wire31924)  &  wire34307 ) | ( (~ wire31925)  &  wire34307 ) | ( (~ wire31924)  &  wire34309 ) | ( (~ wire31925)  &  wire34309 ) ;
 assign wire34356 = ( (~ wire31924)  &  wire34311 ) | ( (~ wire31925)  &  wire34311 ) | ( (~ wire31924)  &  wire34313 ) | ( (~ wire31925)  &  wire34313 ) ;
 assign wire34357 = ( (~ wire31924)  &  wire34315 ) | ( (~ wire31925)  &  wire34315 ) | ( (~ wire31924)  &  wire34317 ) | ( (~ wire31925)  &  wire34317 ) ;
 assign wire34358 = ( (~ wire31924)  &  wire34319 ) | ( (~ wire31925)  &  wire34319 ) | ( (~ wire31924)  &  wire34321 ) | ( (~ wire31925)  &  wire34321 ) ;
 assign wire34359 = ( (~ wire31924)  &  wire34323 ) | ( (~ wire31925)  &  wire34323 ) | ( (~ wire31924)  &  wire34325 ) | ( (~ wire31925)  &  wire34325 ) ;
 assign wire34360 = ( (~ wire31924)  &  wire34327 ) | ( (~ wire31925)  &  wire34327 ) | ( (~ wire31924)  &  wire34332 ) | ( (~ wire31925)  &  wire34332 ) ;
 assign wire34361 = ( (~ wire31924)  &  wire34333 ) | ( (~ wire31925)  &  wire34333 ) | ( (~ wire31924)  &  wire34334 ) | ( (~ wire31925)  &  wire34334 ) ;
 assign wire34362 = ( ng10711  &  (~ wire31924) ) | ( ng10711  &  (~ wire31925) ) | ( (~ wire31924)  &  wire34335 ) | ( (~ wire31925)  &  wire34335 ) ;
 assign wire34363 = ( wire34336 ) | ( wire34337 ) | ( wire34338 ) | ( wire34339 ) ;
 assign wire34364 = ( wire34340 ) | ( wire34341 ) | ( wire34342 ) | ( wire34343 ) ;
 assign wire34371 = ( wire34364 ) | ( wire34363 ) ;
 assign wire34372 = ( wire34351 ) | ( wire34352 ) | ( wire34353 ) | ( wire34354 ) ;
 assign wire34373 = ( wire34355 ) | ( wire34356 ) | ( wire34357 ) | ( wire34358 ) ;
 assign wire34374 = ( wire34359 ) | ( wire34360 ) | ( wire34361 ) | ( wire34362 ) ;
 assign wire34385 = ( wire3049 ) | ( wire6818 ) | ( wire6819 ) | ( wire6820 ) ;
 assign wire34386 = ( wire6821 ) | ( wire6822 ) | ( wire6823 ) | ( wire6824 ) ;
 assign wire34389 = ( (~ ng1192)  &  ng1312 ) ;
 assign wire34390 = ( ng1193  &  ng1192 ) | ( pg16355  &  (~ ng1312)  &  (~ ng1192) ) ;
 assign wire34395 = ( (~ ng28556)  &  (~ ng26938)  &  wire32600 ) | ( (~ ng28556)  &  (~ ng26938)  &  wire32601 ) | ( (~ ng28556)  &  ng26938  &  (~ wire32600)  &  (~ wire32601) ) ;
 assign wire34402 = ( (~ ng28584)  &  ng26417  &  wire33448 ) | ( (~ ng28584)  &  ng26417  &  wire33449 ) | ( (~ ng28584)  &  (~ ng26417)  &  (~ wire33448)  &  (~ wire33449) ) ;
 assign wire34403 = ( ng2175  &  ng27756 ) | ( ng25874  &  (~ ng27756)  &  (~ ng16693) ) ;
 assign wire34410 = ( (~ ng17031)  &  ng2133 ) ;
 assign wire34412 = ( (~ ng17031)  &  ng2129 ) ;
 assign wire34418 = ( ng2466  &  ng2463  &  ng2473 ) | ( ng2466  &  ng2463  &  (~ ng826) ) ;
 assign wire34419 = ( ng2466  &  ng2473  &  (~ ng823) ) | ( ng2466  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire34421 = ( wire3046 ) | ( wire6732 ) | ( wire34418 ) ;
 assign wire34422 = ( wire6737 ) | ( wire6738 ) | ( wire34419 ) ;
 assign wire34428 = ( (~ ng2185)  &  wire3066  &  wire33518 ) | ( (~ ng2185)  &  wire3066  &  wire33519 ) | ( ng2185  &  wire3066  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire34429 = ( (~ ng18319)  &  (~ ng18395)  &  (~ ng18478)  &  (~ ng18578) ) ;
 assign wire34430 = ( (~ ng18606)  &  (~ ng18053)  &  (~ ng18231)  &  wire3055 ) ;
 assign wire34432 = ( wire33528  &  (~ wire33538)  &  (~ wire33539) ) | ( wire33529  &  (~ wire33538)  &  (~ wire33539) ) ;
 assign wire34434 = ( ng23537  &  (~ wire33528)  &  (~ wire33529) ) ;
 assign wire34435 = ( (~ wire33538)  &  (~ wire33539)  &  wire33548 ) | ( (~ wire33538)  &  (~ wire33539)  &  wire33549 ) ;
 assign wire34438 = ( (~ ng11687)  &  ng11653 ) | ( (~ ng2257)  &  ng11687  &  (~ ng11653) ) | ( (~ ng11687)  &  (~ ng11653)  &  ng11678 ) ;
 assign wire34439 = ( wire34438 ) | ( (~ ng23537)  &  (~ ng11678)  &  wire34432 ) ;
 assign wire34440 = ( wire34439 ) | ( ng23533  &  ng23521  &  wire34434 ) ;
 assign wire34449 = ( ng2707  &  ng2727 ) ;
 assign wire34450 = ( ng1315  &  ng2714  &  (~ ng2733) ) ;
 assign wire34451 = ( (~ ng1312)  &  ng2707 ) | ( (~ ng2704)  &  ng2707 ) ;
 assign wire34452 = ( (~ ng2727)  &  wire34451 ) | ( (~ ng2707)  &  wire34451 ) | ( (~ wire34450)  &  wire34451 ) ;
 assign wire34453 = ( ng2727  &  (~ ng1312) ) | ( ng2727  &  (~ ng2704) ) ;
 assign wire34459 = ( ng2805  &  (~ ng1309)  &  ng2807 ) | ( ng2805  &  ng2806  &  ng2807 ) ;
 assign wire34460 = ( ng2805  &  (~ ng1312)  &  ng2806 ) | ( (~ ng1312)  &  (~ ng1315)  &  ng2806 ) ;
 assign wire34462 = ( wire3049 ) | ( wire6633 ) | ( wire34459 ) ;
 assign wire34463 = ( wire6638 ) | ( wire6639 ) | ( wire34460 ) ;
 assign wire34469 = ( ng2772  &  (~ ng1309)  &  ng2774 ) | ( ng2772  &  ng2773  &  ng2774 ) ;
 assign wire34470 = ( ng2772  &  (~ ng1312)  &  ng2773 ) | ( (~ ng1312)  &  (~ ng1315)  &  ng2773 ) ;
 assign wire34472 = ( wire3049 ) | ( wire6609 ) | ( wire34469 ) ;
 assign wire34473 = ( wire6614 ) | ( wire6615 ) | ( wire34470 ) ;
 assign wire34482 = ( (~ ng1312)  &  (~ ng1315)  &  ng2779 ) | ( (~ ng1312)  &  ng2779  &  ng2778 ) ;
 assign wire34484 = ( wire3049 ) | ( wire6617 ) | ( wire6618 ) | ( wire6619 ) ;
 assign wire34485 = ( wire6622 ) | ( wire6623 ) | ( wire34482 ) ;
 assign wire34496 = ( wire3049 ) | ( wire6625 ) | ( wire6626 ) | ( wire6627 ) ;
 assign wire34497 = ( wire6628 ) | ( wire6629 ) | ( wire6630 ) | ( wire6631 ) ;
 assign wire34505 = ( ng2786  &  ng2784  &  ng2785 ) | ( ng2784  &  (~ ng1312)  &  ng2785 ) ;
 assign wire34508 = ( wire3049 ) | ( wire6641 ) | ( wire34505 ) ;
 assign wire34509 = ( wire6644 ) | ( wire6645 ) | ( wire6646 ) | ( wire6647 ) ;
 assign wire34517 = ( ng2797  &  (~ ng1315)  &  ng2798 ) | ( ng2797  &  ng2796  &  ng2798 ) ;
 assign wire34518 = ( ng2797  &  (~ ng1312)  &  (~ ng1315) ) | ( ng2797  &  (~ ng1312)  &  ng2796 ) ;
 assign wire34520 = ( wire3049 ) | ( wire6649 ) | ( wire34517 ) ;
 assign wire34521 = ( wire6654 ) | ( wire6655 ) | ( wire34518 ) ;
 assign wire34530 = ( (~ ng1312)  &  (~ ng1315)  &  ng2788 ) | ( (~ ng1312)  &  ng2787  &  ng2788 ) ;
 assign wire34532 = ( wire3049 ) | ( wire6689 ) | ( wire6690 ) | ( wire6691 ) ;
 assign wire34533 = ( wire6694 ) | ( wire6695 ) | ( wire34530 ) ;
 assign wire34544 = ( wire3049 ) | ( wire6681 ) | ( wire6682 ) | ( wire6683 ) ;
 assign wire34545 = ( wire6684 ) | ( wire6685 ) | ( wire6686 ) | ( wire6687 ) ;
 assign wire34553 = ( ng2793  &  (~ ng1312)  &  ng2794 ) | ( ng2793  &  ng2795  &  ng2794 ) ;
 assign wire34556 = ( wire3049 ) | ( wire6657 ) | ( wire34553 ) ;
 assign wire34557 = ( wire6660 ) | ( wire6661 ) | ( wire6662 ) | ( wire6663 ) ;
 assign wire34566 = ( (~ ng1312)  &  (~ ng1315)  &  ng2776 ) | ( (~ ng1315)  &  ng2777  &  ng2776 ) ;
 assign wire34568 = ( wire3049 ) | ( wire6665 ) | ( wire6666 ) | ( wire6667 ) ;
 assign wire34569 = ( wire6670 ) | ( wire6671 ) | ( wire34566 ) ;
 assign wire34578 = ( (~ ng1312)  &  (~ ng1315)  &  ng2782 ) | ( (~ ng1315)  &  ng2783  &  ng2782 ) ;
 assign wire34580 = ( wire3049 ) | ( wire6673 ) | ( wire6674 ) | ( wire6675 ) ;
 assign wire34581 = ( wire6678 ) | ( wire6679 ) | ( wire34578 ) ;
 assign wire34584 = ( ng2714  &  ng11964  &  wire34462 ) | ( (~ ng2714)  &  (~ ng11964)  &  wire34462 ) | ( ng2714  &  ng11964  &  wire34463 ) | ( (~ ng2714)  &  (~ ng11964)  &  wire34463 ) ;
 assign wire34585 = ( ng2727  &  ng12068  &  wire34462 ) | ( (~ ng2727)  &  (~ ng12068)  &  wire34462 ) | ( ng2727  &  ng12068  &  wire34463 ) | ( (~ ng2727)  &  (~ ng12068)  &  wire34463 ) ;
 assign wire34586 = ( ng2766  &  ng11965  &  wire34462 ) | ( (~ ng2766)  &  (~ ng11965)  &  wire34462 ) | ( ng2766  &  ng11965  &  wire34463 ) | ( (~ ng2766)  &  (~ ng11965)  &  wire34463 ) ;
 assign wire34587 = ( ng2734  &  ng12234  &  wire34508 ) | ( ng2734  &  ng12234  &  wire34509 ) | ( (~ ng2734)  &  ng12234  &  (~ wire34508)  &  (~ wire34509) ) ;
 assign wire34588 = ( ng2760  &  ng12234  &  wire34520 ) | ( ng2760  &  ng12234  &  wire34521 ) | ( (~ ng2760)  &  ng12234  &  (~ wire34520)  &  (~ wire34521) ) ;
 assign wire34589 = ( ng2746  &  ng12234  &  wire34532 ) | ( ng2746  &  ng12234  &  wire34533 ) | ( (~ ng2746)  &  ng12234  &  (~ wire34532)  &  (~ wire34533) ) ;
 assign wire34590 = ( ng2740  &  ng12234  &  wire34544 ) | ( ng2740  &  ng12234  &  wire34545 ) | ( (~ ng2740)  &  ng12234  &  (~ wire34544)  &  (~ wire34545) ) ;
 assign wire34591 = ( ng2753  &  ng12234  &  wire34556 ) | ( ng2753  &  ng12234  &  wire34557 ) | ( (~ ng2753)  &  ng12234  &  (~ wire34556)  &  (~ wire34557) ) ;
 assign wire34592 = ( ng2707  &  ng12234  &  wire34568 ) | ( ng2707  &  ng12234  &  wire34569 ) | ( (~ ng2707)  &  ng12234  &  (~ wire34568)  &  (~ wire34569) ) ;
 assign wire34598 = ( wire34592 ) | ( ng2720  &  ng12124  &  ng12234 ) | ( (~ ng2720)  &  (~ ng12124)  &  ng12234 ) ;
 assign wire34599 = ( wire34584 ) | ( wire34585 ) | ( wire34586 ) | ( wire34587 ) ;
 assign wire34600 = ( wire34588 ) | ( wire34589 ) | ( wire34590 ) | ( wire34591 ) ;
 assign wire34603 = ( ng2804  &  ng2803  &  ng2802 ) ;
 assign wire34605 = ( (~ ng1312)  &  ng2803  &  ng2802 ) ;
 assign wire34607 = ( (~ ng1309)  &  ng2804  &  ng2802 ) ;
 assign wire34609 = ( (~ ng1315)  &  ng2804  &  ng2803 ) ;
 assign wire34610 = ( (~ ng1312)  &  (~ ng1315)  &  ng2803 ) ;
 assign wire34611 = ( (~ ng1312)  &  (~ ng1309)  &  ng2802 ) ;
 assign wire34612 = ( (~ ng1315)  &  (~ ng1309)  &  ng2804 ) ;
 assign wire34617 = ( wire6581 ) | ( wire6582 ) | ( wire6583 ) | ( wire6584 ) ;
 assign wire34618 = ( wire6585 ) | ( wire6586 ) | ( wire6587 ) | ( wire6588 ) ;
 assign wire34619 = ( ng12146  &  wire3174 ) | ( wire3174  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire34620 = ( ng529  &  wire3138 ) | ( ng21851  &  wire3138 ) | ( wire3138  &  wire34028 ) ;
 assign wire34622 = ( ng17973 ) | ( (~ ng3125)  &  (~ ng8381)  &  (~ wire30893) ) ;
 assign wire34625 = ( ng83  &  ng88  &  ng79  &  ng92 ) ;
 assign wire34633 = ( ng391  &  ng388  &  ng398 ) | ( ng391  &  ng388  &  (~ ng826) ) ;
 assign wire34634 = ( ng391  &  ng398  &  (~ ng823) ) | ( ng391  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire34636 = ( wire3046 ) | ( wire6547 ) | ( wire34633 ) ;
 assign wire34637 = ( wire6552 ) | ( wire6553 ) | ( wire34634 ) ;
 assign wire34638 = ( (~ wire31324)  &  (~ wire31325)  &  wire34636 ) | ( (~ wire31324)  &  (~ wire31325)  &  wire34637 ) ;
 assign wire34642 = ( ng448  &  ng449  &  (~ ng853)  &  ng2257 ) ;
 assign wire34645 = ( ng449  &  (~ ng826)  &  ng447  &  ng2257 ) ;
 assign wire34648 = ( ng448  &  ng449  &  ng447  &  ng2257 ) ;
 assign wire34651 = ( ng448  &  ng447  &  (~ ng823)  &  ng2257 ) ;
 assign wire34653 = ( (~ ng826)  &  ng447  &  (~ ng823)  &  ng2257 ) ;
 assign wire34655 = ( ng448  &  (~ ng823)  &  (~ ng853)  &  ng2257 ) ;
 assign wire34657 = ( ng449  &  (~ ng826)  &  (~ ng853)  &  ng2257 ) ;
 assign wire34658 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2257 ) ;
 assign wire34663 = ( wire6532 ) | ( wire6533 ) | ( wire6534 ) | ( wire6535 ) ;
 assign wire34664 = ( wire6536 ) | ( wire6537 ) | ( wire6538 ) | ( wire6539 ) ;
 assign wire34668 = ( ng2257  &  ng11975  &  (~ ng17985)  &  ng11935 ) | ( ng2257  &  (~ ng11975)  &  ng17985  &  (~ ng11935) ) ;
 assign wire34675 = ( (~ ng1312)  &  (~ ng1315)  &  ng479 ) | ( (~ ng1312)  &  ng479  &  ng478 ) ;
 assign wire34677 = ( wire3049 ) | ( wire6514 ) | ( wire6515 ) | ( wire6516 ) ;
 assign wire34679 = ( wire31502  &  wire31512 ) | ( wire31503  &  wire31512 ) | ( wire31502  &  wire31513 ) | ( wire31503  &  wire31513 ) ;
 assign wire34686 = ( (~ ng28529)  &  (~ ng26915)  &  wire31857 ) | ( (~ ng28529)  &  (~ ng26915)  &  wire31858 ) | ( (~ ng28529)  &  ng26915  &  (~ wire31857)  &  (~ wire31858) ) ;
 assign wire34689 = ( (~ ng28529)  &  (~ ng26906)  &  wire31907 ) | ( (~ ng28529)  &  (~ ng26906)  &  wire31908 ) | ( (~ ng28529)  &  ng26906  &  (~ wire31907)  &  (~ wire31908) ) ;
 assign wire34690 = ( (~ ng11833)  &  ng27743 ) | ( (~ ng16655)  &  ng25818  &  (~ ng27743) ) ;
 assign wire34696 = ( (~ ng1119)  &  (~ ng1116)  &  (~ ng1122) ) | ( (~ ng1119)  &  (~ ng1122)  &  (~ ng826) ) ;
 assign wire34697 = ( (~ ng1116)  &  (~ ng1122)  &  (~ ng823) ) | ( (~ ng1122)  &  (~ ng826)  &  (~ ng823) ) ;
 assign wire34700 = ( wire6473 ) | ( wire6474 ) | ( wire34697 ) ;
 assign wire34706 = ( ng866  &  ng865  &  ng867 ) | ( (~ ng826)  &  ng865  &  ng867 ) ;
 assign wire34707 = ( ng866  &  ng865  &  (~ ng823) ) | ( (~ ng826)  &  ng865  &  (~ ng823) ) ;
 assign wire34709 = ( wire3046 ) | ( wire6459 ) | ( (~ wire32224) ) | ( (~ wire32225) ) ;
 assign wire34710 = ( wire34707 ) | ( wire34706 ) ;
 assign wire34716 = ( (~ ng853)  &  ng1135  &  ng1136  &  ng2257 ) ;
 assign wire34719 = ( ng1134  &  ng1135  &  ng1136  &  ng2257 ) ;
 assign wire34722 = ( ng1134  &  (~ ng826)  &  ng1136  &  ng2257 ) ;
 assign wire34725 = ( ng1134  &  (~ ng823)  &  ng1135  &  ng2257 ) ;
 assign wire34727 = ( ng1134  &  (~ ng826)  &  (~ ng823)  &  ng2257 ) ;
 assign wire34729 = ( (~ ng823)  &  (~ ng853)  &  ng1135  &  ng2257 ) ;
 assign wire34731 = ( (~ ng826)  &  (~ ng853)  &  ng1136  &  ng2257 ) ;
 assign wire34732 = ( (~ ng826)  &  (~ ng823)  &  (~ ng853)  &  ng2257 ) ;
 assign wire34737 = ( wire6441 ) | ( wire6442 ) | ( wire6443 ) | ( wire6444 ) ;
 assign wire34738 = ( wire6445 ) | ( wire6446 ) | ( wire6447 ) | ( wire6448 ) ;
 assign wire34741 = ( ng2257  &  ng12044  &  (~ ng18102)  &  ng11988 ) | ( ng2257  &  (~ ng12044)  &  ng18102  &  (~ ng11988) ) ;
 assign wire34742 = ( wire6434 ) | ( ng1010  &  (~ ng823) ) ;
 assign wire34743 = ( wire34742 ) | ( (~ ng15950)  &  ng17086  &  (~ ng27850) ) ;
 assign wire34744 = ( ng13055  &  wire32387 ) | ( ng13055  &  wire32388 ) | ( ng13055  &  wire32389 ) ;
 assign wire34746 = ( ng13055  &  wire32534 ) | ( ng13055  &  wire32535 ) | ( ng13055  &  wire32536 ) ;
 assign wire34747 = ( (~ wire32559)  &  (~ wire32560)  &  (~ wire32561)  &  wire34746 ) ;
 assign wire34748 = ( wire6425 ) | ( (~ ng23071)  &  (~ ng18598)  &  wire34744 ) ;
 assign wire34755 = ( (~ ng1312)  &  (~ ng1315)  &  ng1418 ) | ( (~ ng1312)  &  ng1418  &  ng1417 ) ;
 assign wire34757 = ( wire3049 ) | ( wire6409 ) | ( wire6410 ) | ( wire6411 ) ;
 assign wire34758 = ( wire6414 ) | ( wire6415 ) | ( wire34755 ) ;
 assign wire34767 = ( wire3049 ) | ( wire6329 ) | ( wire6330 ) | ( wire6331 ) ;
 assign wire34768 = ( wire6332 ) | ( wire6333 ) | ( wire6334 ) | ( wire6335 ) ;
 assign wire34776 = ( ng1403  &  ng1404  &  ng1402 ) | ( ng1403  &  (~ ng1312)  &  ng1402 ) ;
 assign wire34777 = ( ng1403  &  ng1404  &  (~ ng1315) ) | ( ng1403  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire34779 = ( wire3049 ) | ( wire6337 ) | ( wire34776 ) ;
 assign wire34780 = ( wire6342 ) | ( wire6343 ) | ( wire34777 ) ;
 assign wire34791 = ( wire3049 ) | ( wire6345 ) | ( wire6346 ) | ( wire6347 ) ;
 assign wire34792 = ( wire6348 ) | ( wire6349 ) | ( wire6350 ) | ( wire6351 ) ;
 assign wire34800 = ( ng1392  &  ng1391  &  ng1390 ) | ( ng1391  &  (~ ng1312)  &  ng1390 ) ;
 assign wire34801 = ( ng1392  &  ng1391  &  (~ ng1315) ) | ( ng1391  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire34803 = ( wire3049 ) | ( wire6353 ) | ( wire34800 ) ;
 assign wire34804 = ( wire6358 ) | ( wire6359 ) | ( wire34801 ) ;
 assign wire34813 = ( (~ ng1312)  &  (~ ng1315)  &  ng1409 ) | ( (~ ng1315)  &  ng1409  &  ng1410 ) ;
 assign wire34815 = ( wire3049 ) | ( wire6361 ) | ( wire6362 ) | ( wire6363 ) ;
 assign wire34816 = ( wire6366 ) | ( wire6367 ) | ( wire34813 ) ;
 assign wire34825 = ( (~ ng1312)  &  (~ ng1315)  &  ng1385 ) | ( (~ ng1312)  &  ng1384  &  ng1385 ) ;
 assign wire34827 = ( wire3049 ) | ( wire6369 ) | ( wire6370 ) | ( wire6371 ) ;
 assign wire34828 = ( wire6374 ) | ( wire6375 ) | ( wire34825 ) ;
 assign wire34836 = ( ng1411  &  ng1413  &  ng1412 ) | ( ng1411  &  (~ ng1312)  &  ng1412 ) ;
 assign wire34839 = ( wire3049 ) | ( wire6377 ) | ( wire34836 ) ;
 assign wire34840 = ( wire6380 ) | ( wire6381 ) | ( wire6382 ) | ( wire6383 ) ;
 assign wire34851 = ( wire3049 ) | ( wire6385 ) | ( wire6386 ) | ( wire6387 ) ;
 assign wire34852 = ( wire6388 ) | ( wire6389 ) | ( wire6390 ) | ( wire6391 ) ;
 assign wire34861 = ( (~ ng1312)  &  (~ ng1315)  &  ng1400 ) | ( (~ ng1315)  &  ng1400  &  ng1401 ) ;
 assign wire34863 = ( wire3049 ) | ( wire6393 ) | ( wire6394 ) | ( wire6395 ) ;
 assign wire34864 = ( wire6398 ) | ( wire6399 ) | ( wire34861 ) ;
 assign wire34873 = ( (~ ng1312)  &  (~ ng1315)  &  ng1406 ) | ( (~ ng1315)  &  ng1406  &  ng1407 ) ;
 assign wire34875 = ( wire3049 ) | ( wire6401 ) | ( wire6402 ) | ( wire6403 ) ;
 assign wire34876 = ( wire6406 ) | ( wire6407 ) | ( wire34873 ) ;
 assign wire34879 = ( ng1346  &  ng12048  &  wire34757 ) | ( (~ ng1346)  &  (~ ng12048)  &  wire34757 ) | ( ng1346  &  ng12048  &  wire34758 ) | ( (~ ng1346)  &  (~ ng12048)  &  wire34758 ) ;
 assign wire34880 = ( ng1352  &  ng12154  &  wire34757 ) | ( (~ ng1352)  &  (~ ng12154)  &  wire34757 ) | ( ng1352  &  ng12154  &  wire34758 ) | ( (~ ng1352)  &  (~ ng12154)  &  wire34758 ) ;
 assign wire34881 = ( ng1319  &  ng11905  &  wire34757 ) | ( (~ ng1319)  &  (~ ng11905)  &  wire34757 ) | ( ng1319  &  ng11905  &  wire34758 ) | ( (~ ng1319)  &  (~ ng11905)  &  wire34758 ) ;
 assign wire34882 = ( ng1339  &  ng11946  &  wire34757 ) | ( (~ ng1339)  &  (~ ng11946)  &  wire34757 ) | ( ng1339  &  ng11946  &  wire34758 ) | ( (~ ng1339)  &  (~ ng11946)  &  wire34758 ) ;
 assign wire34883 = ( ng1372  &  ng12100  &  wire34815 ) | ( ng1372  &  ng12100  &  wire34816 ) | ( (~ ng1372)  &  ng12100  &  (~ wire34815)  &  (~ wire34816) ) ;
 assign wire34884 = ( ng1326  &  ng11872  &  wire34757 ) | ( (~ ng1326)  &  (~ ng11872)  &  wire34757 ) | ( ng1326  &  ng11872  &  wire34758 ) | ( (~ ng1326)  &  (~ ng11872)  &  wire34758 ) ;
 assign wire34885 = ( ng1378  &  ng12100  &  wire34839 ) | ( ng1378  &  ng12100  &  wire34840 ) | ( (~ ng1378)  &  ng12100  &  (~ wire34839)  &  (~ wire34840) ) ;
 assign wire34886 = ( ng1332  &  ng11991  &  wire34757 ) | ( (~ ng1332)  &  (~ ng11991)  &  wire34757 ) | ( ng1332  &  ng11991  &  wire34758 ) | ( (~ ng1332)  &  (~ ng11991)  &  wire34758 ) ;
 assign wire34887 = ( ng1358  &  ng12099  &  wire34757 ) | ( (~ ng1358)  &  (~ ng12099)  &  wire34757 ) | ( ng1358  &  ng12099  &  wire34758 ) | ( (~ ng1358)  &  (~ ng12099)  &  wire34758 ) ;
 assign wire34893 = ( wire34887 ) | ( ng1365  &  ng12100  &  ng12208 ) | ( (~ ng1365)  &  ng12100  &  (~ ng12208) ) ;
 assign wire34894 = ( wire34879 ) | ( wire34880 ) | ( wire34881 ) | ( wire34882 ) ;
 assign wire34895 = ( wire34883 ) | ( wire34884 ) | ( wire34885 ) | ( wire34886 ) ;
 assign wire34898 = ( ng1416  &  ng1415  &  ng1414 ) ;
 assign wire34900 = ( (~ ng1312)  &  ng1415  &  ng1414 ) ;
 assign wire34902 = ( ng1416  &  (~ ng1309)  &  ng1414 ) ;
 assign wire34904 = ( (~ ng1315)  &  ng1416  &  ng1415 ) ;
 assign wire34905 = ( (~ ng1312)  &  (~ ng1315)  &  ng1415 ) ;
 assign wire34906 = ( (~ ng1312)  &  (~ ng1309)  &  ng1414 ) ;
 assign wire34907 = ( (~ ng1315)  &  ng1416  &  (~ ng1309) ) ;
 assign wire34912 = ( wire6301 ) | ( wire6302 ) | ( wire6303 ) | ( wire6304 ) ;
 assign wire34913 = ( wire6305 ) | ( wire6306 ) | ( wire6307 ) | ( wire6308 ) ;
 assign wire34916 = ( (~ ng28556)  &  wire3302  &  wire32712 ) | ( (~ ng28556)  &  wire3302  &  wire32713 ) | ( (~ ng28556)  &  (~ wire3302)  &  (~ wire32712)  &  (~ wire32713) ) ;
 assign wire34924 = ( ng1769  &  ng1779  &  ng1772 ) | ( ng1779  &  ng1772  &  (~ ng823) ) ;
 assign wire34927 = ( wire3046 ) | ( wire6278 ) | ( wire34924 ) ;
 assign wire34928 = ( wire6281 ) | ( wire6282 ) | ( wire6283 ) | ( wire6284 ) ;
 assign wire34932 = ( (~ ng23526)  &  (~ wire32944) ) | ( (~ ng23526)  &  (~ wire32650)  &  (~ wire32651) ) ;
 assign wire34933 = ( wire6263 ) | ( ng1703  &  (~ ng826) ) ;
 assign wire34934 = ( wire34933 ) | ( (~ ng15970)  &  ng17124  &  (~ ng27875) ) ;
 assign wire34937 = ( (~ ng28584)  &  (~ ng26947)  &  wire33518 ) | ( (~ ng28584)  &  (~ ng26947)  &  wire33519 ) | ( (~ ng28584)  &  ng26947  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire34948 = ( wire3049 ) | ( wire6217 ) | ( wire6218 ) | ( wire6219 ) ;
 assign wire34949 = ( wire6220 ) | ( wire6221 ) | ( wire6222 ) | ( wire6223 ) ;
 assign wire34956 = ( (~ ng1312)  &  (~ ng1315)  &  ng2554 ) | ( (~ ng1312)  &  ng2554  &  ng2553 ) ;
 assign wire34958 = ( wire3049 ) | ( wire6207 ) | ( wire6208 ) | ( wire6209 ) ;
 assign wire34962 = ( wire3188  &  ng11979 ) | ( wire3188  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire34963 = ( ng532  &  wire3138 ) | ( ng21851  &  wire3138 ) | ( wire3138  &  wire34028 ) ;
 assign wire34965 = ( ng17973 ) | ( wire3282  &  (~ ng8381)  &  (~ wire34079) ) ;
 assign wire34969 = ( wire6178 ) | ( wire6177 ) ;
 assign wire34970 = ( wire6179 ) | ( wire6180 ) | ( wire34965 ) ;
 assign wire34971 = ( ng3120  &  wire3217 ) | ( ng3120  &  wire3397 ) ;
 assign wire34972 = ( ng3087  &  (~ ng15757) ) | ( ng3211  &  (~ ng15841) ) ;
 assign wire34973 = ( ng3210  &  (~ ng15830) ) | ( ng3086  &  (~ ng15719) ) ;
 assign wire34974 = ( wire6170 ) | ( wire6171 ) | ( wire6175 ) | ( wire6176 ) ;
 assign wire34978 = ( wire34969 ) | ( wire34970 ) | ( wire34971 ) | ( wire34972 ) ;
 assign wire34982 = ( (~ ng28501)  &  (~ ng26892)  &  wire31038 ) | ( (~ ng28501)  &  (~ ng26892)  &  wire31039 ) | ( (~ ng28501)  &  ng26892  &  (~ wire31038)  &  (~ wire31039) ) ;
 assign wire34983 = ( (~ ng11800)  &  ng27738 ) | ( (~ ng16643)  &  ng25764  &  (~ ng27738) ) ;
 assign wire34985 = ( ng83  &  (~ ng17031)  &  (~ ng23497) ) ;
 assign wire34987 = ( wire31314  &  wire31334 ) | ( wire31315  &  wire31334 ) | ( wire31314  &  wire31335 ) | ( wire31315  &  wire31335 ) ;
 assign wire34989 = ( ng660  &  ng672  &  ng666 ) ;
 assign wire34990 = ( ng672  &  (~ ng1312) ) | ( ng672  &  (~ ng630) ) ;
 assign wire34992 = ( (~ ng1312)  &  ng666 ) | ( ng666  &  (~ ng630) ) ;
 assign wire34996 = ( wire6103 ) | ( ng1009  &  (~ ng826) ) ;
 assign wire34997 = ( wire34996 ) | ( (~ ng15970)  &  ng17086  &  (~ ng27850) ) ;
 assign wire35003 = ( ng1151  &  ng1171  &  ng1167 ) | ( ng1151  &  (~ ng1315)  &  ng1167 ) ;
 assign wire35004 = ( ng1151  &  ng1171  &  (~ ng1312) ) | ( ng1151  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire35007 = ( wire6094 ) | ( wire6095 ) | ( wire35004 ) ;
 assign wire35013 = ( wire6055 ) | ( ng1704  &  (~ ng823) ) ;
 assign wire35014 = ( wire35013 ) | ( (~ ng15950)  &  ng17124  &  (~ ng27875) ) ;
 assign wire35018 = ( (~ ng23537)  &  (~ wire33792) ) | ( (~ ng23537)  &  (~ wire33548)  &  (~ wire33549) ) ;
 assign wire35019 = ( wire6015 ) | ( ng2397  &  (~ ng826) ) ;
 assign wire35020 = ( wire35019 ) | ( (~ ng15970)  &  ng17151  &  (~ ng27892) ) ;
 assign wire35021 = ( (~ ng1312)  &  (~ ng2734) ) | ( (~ ng2734)  &  (~ ng2704) ) ;
 assign wire35022 = ( (~ ng1312)  &  ng2734 ) | ( ng2734  &  (~ ng2704) ) ;
 assign wire35023 = ( ng12035  &  wire3174 ) | ( wire3174  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35029 = ( (~ ng2900)  &  ng2888  &  (~ ng2896)  &  ng2892 ) ;
 assign wire35030 = ( ng2950  &  ng2903  &  (~ ng2883)  &  ng2908 ) ;
 assign wire35032 = ( ng2950  &  ng2892 ) ;
 assign wire35033 = ( ng2888  &  ng2896  &  ng2883 ) ;
 assign wire35038 = ( (~ ng28501)  &  ng26283  &  wire31028 ) | ( (~ ng28501)  &  ng26283  &  wire31029 ) | ( (~ ng28501)  &  (~ ng26283)  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire35039 = ( ng105  &  ng27738 ) | ( (~ ng16643)  &  ng25764  &  (~ ng27738) ) ;
 assign wire35040 = ( (~ ng12967)  &  (~ wire30977)  &  (~ wire30978)  &  wire30979 ) ;
 assign wire35041 = ( ng27563  &  (~ wire31279)  &  wire35040 ) ;
 assign wire35042 = ( (~ ng12849)  &  (~ wire30977)  &  (~ wire30978)  &  wire30979 ) ;
 assign wire35043 = ( (~ wire30988)  &  (~ wire30989)  &  (~ wire30998)  &  (~ wire30999) ) ;
 assign wire35044 = ( (~ ng27563)  &  (~ wire30998)  &  (~ wire30999) ) | ( (~ wire30998)  &  (~ wire30999)  &  wire31279 ) ;
 assign wire35045 = ( ng27563  &  (~ ng16643)  &  (~ wire31279)  &  (~ wire31281) ) ;
 assign wire35046 = ( (~ ng28501)  &  wire35044 ) | ( (~ ng28501)  &  wire35045 ) ;
 assign wire35047 = ( (~ ng28501)  &  ng26902  &  wire35041 ) | ( (~ ng28501)  &  ng26902  &  wire35042 ) ;
 assign wire35057 = ( ng65  &  ng70  &  ng61 ) ;
 assign wire35060 = ( (~ ng92)  &  (~ wire31048)  &  (~ wire31049) ) ;
 assign wire35061 = ( (~ ng92)  &  (~ wire31048)  &  (~ wire31049) ) ;
 assign wire35062 = ( ng92  &  wire31048 ) | ( ng92  &  wire31049 ) ;
 assign wire35063 = ( ng92  &  wire31048 ) | ( ng92  &  wire31049 ) ;
 assign wire35064 = ( (~ ng56)  &  (~ wire31038)  &  (~ wire31039) ) ;
 assign wire35065 = ( (~ ng56)  &  (~ wire31038)  &  (~ wire31039) ) ;
 assign wire35066 = ( ng56  &  wire31038 ) | ( ng56  &  wire31039 ) ;
 assign wire35067 = ( ng56  &  wire31038 ) | ( ng56  &  wire31039 ) ;
 assign wire35068 = ( (~ ng83)  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire35069 = ( (~ ng83)  &  (~ wire31028)  &  (~ wire31029) ) ;
 assign wire35070 = ( ng83  &  wire31028 ) | ( ng83  &  wire31029 ) ;
 assign wire35071 = ( ng83  &  wire31028 ) | ( ng83  &  wire31029 ) ;
 assign wire35072 = ( (~ ng52)  &  (~ wire30937)  &  (~ wire30938) ) ;
 assign wire35073 = ( ng52  &  wire30937 ) | ( ng52  &  wire30938 ) ;
 assign wire35074 = ( (~ ng61)  &  (~ wire31008)  &  (~ wire31009) ) ;
 assign wire35075 = ( ng61  &  wire31008 ) | ( ng61  &  wire31009 ) ;
 assign wire35076 = ( (~ ng70)  &  (~ wire30998)  &  (~ wire30999) ) ;
 assign wire35077 = ( ng70  &  wire30998 ) | ( ng70  &  wire30999 ) ;
 assign wire35078 = ( (~ ng65)  &  (~ wire30947)  &  (~ wire30948) ) ;
 assign wire35079 = ( ng65  &  wire30947 ) | ( ng65  &  wire30948 ) ;
 assign wire35080 = ( (~ ng88)  &  (~ wire31018)  &  (~ wire31019) ) ;
 assign wire35081 = ( ng88  &  wire31018 ) | ( ng88  &  wire31019 ) ;
 assign wire35082 = ( (~ ng74)  &  (~ wire30988)  &  (~ wire30989) ) ;
 assign wire35083 = ( ng74  &  wire30988 ) | ( ng74  &  wire30989 ) ;
 assign wire35084 = ( (~ ng79)  &  (~ wire30927)  &  (~ wire30928) ) ;
 assign wire35085 = ( ng79  &  wire30927 ) | ( ng79  &  wire30928 ) ;
 assign wire35086 = ( (~ ng52)  &  (~ wire30937)  &  (~ wire30938) ) ;
 assign wire35087 = ( ng52  &  wire30937 ) | ( ng52  &  wire30938 ) ;
 assign wire35088 = ( (~ ng61)  &  (~ wire31008)  &  (~ wire31009) ) ;
 assign wire35089 = ( ng61  &  wire31008 ) | ( ng61  &  wire31009 ) ;
 assign wire35090 = ( (~ ng70)  &  (~ wire30998)  &  (~ wire30999) ) ;
 assign wire35091 = ( ng70  &  wire30998 ) | ( ng70  &  wire30999 ) ;
 assign wire35092 = ( (~ ng65)  &  (~ wire30947)  &  (~ wire30948) ) ;
 assign wire35093 = ( ng65  &  wire30947 ) | ( ng65  &  wire30948 ) ;
 assign wire35094 = ( (~ ng88)  &  (~ wire31018)  &  (~ wire31019) ) ;
 assign wire35095 = ( ng88  &  wire31018 ) | ( ng88  &  wire31019 ) ;
 assign wire35096 = ( (~ ng74)  &  (~ wire30988)  &  (~ wire30989) ) ;
 assign wire35097 = ( ng74  &  wire30988 ) | ( ng74  &  wire30989 ) ;
 assign wire35098 = ( (~ ng79)  &  (~ wire30927)  &  (~ wire30928) ) ;
 assign wire35099 = ( ng79  &  wire30927 ) | ( ng79  &  wire30928 ) ;
 assign wire35100 = ( (~ ng11644)  &  wire35060 ) | ( (~ ng13378)  &  wire35060 ) | ( (~ ng11624)  &  wire35060 ) | ( (~ ng11644)  &  ng13378  &  (~ ng11624) ) ;
 assign wire35101 = ( (~ ng11624)  &  wire35062 ) | ( (~ wire31067)  &  wire35062 ) | ( (~ ng11624)  &  wire35064 ) | ( (~ wire31067)  &  wire35064 ) ;
 assign wire35102 = ( (~ ng11624)  &  wire35066 ) | ( (~ wire31067)  &  wire35066 ) | ( (~ ng11624)  &  wire35068 ) | ( (~ wire31067)  &  wire35068 ) ;
 assign wire35103 = ( (~ ng11624)  &  wire35070 ) | ( (~ wire31067)  &  wire35070 ) | ( (~ ng11624)  &  wire35072 ) | ( (~ wire31067)  &  wire35072 ) ;
 assign wire35104 = ( (~ ng11624)  &  wire35073 ) | ( (~ wire31067)  &  wire35073 ) | ( (~ ng11624)  &  wire35074 ) | ( (~ wire31067)  &  wire35074 ) ;
 assign wire35105 = ( (~ ng11624)  &  wire35075 ) | ( (~ wire31067)  &  wire35075 ) | ( (~ ng11624)  &  wire35076 ) | ( (~ wire31067)  &  wire35076 ) ;
 assign wire35106 = ( (~ ng11624)  &  wire35077 ) | ( (~ wire31067)  &  wire35077 ) | ( (~ ng11624)  &  wire35078 ) | ( (~ wire31067)  &  wire35078 ) ;
 assign wire35107 = ( (~ ng11624)  &  wire35079 ) | ( (~ wire31067)  &  wire35079 ) | ( (~ ng11624)  &  wire35080 ) | ( (~ wire31067)  &  wire35080 ) ;
 assign wire35108 = ( (~ ng11624)  &  wire35081 ) | ( (~ wire31067)  &  wire35081 ) | ( (~ ng11624)  &  wire35082 ) | ( (~ wire31067)  &  wire35082 ) ;
 assign wire35109 = ( (~ ng11624)  &  wire35083 ) | ( (~ wire31067)  &  wire35083 ) | ( (~ ng11624)  &  wire35084 ) | ( (~ wire31067)  &  wire35084 ) ;
 assign wire35110 = ( (~ ng11624)  &  ng10711 ) | ( ng10711  &  (~ wire31067) ) | ( (~ ng11624)  &  wire35085 ) | ( (~ wire31067)  &  wire35085 ) ;
 assign wire35115 = ( wire35109 ) | ( wire35108 ) ;
 assign wire35116 = ( wire35110 ) | ( (~ wire31065)  &  wire35061 ) | ( (~ wire31066)  &  wire35061 ) ;
 assign wire35117 = ( (~ wire31065)  &  wire35063 ) | ( (~ wire31066)  &  wire35063 ) | ( (~ wire31065)  &  wire35065 ) | ( (~ wire31066)  &  wire35065 ) ;
 assign wire35118 = ( (~ wire31065)  &  wire35067 ) | ( (~ wire31066)  &  wire35067 ) | ( (~ wire31065)  &  wire35069 ) | ( (~ wire31066)  &  wire35069 ) ;
 assign wire35119 = ( (~ wire31065)  &  wire35071 ) | ( (~ wire31066)  &  wire35071 ) | ( (~ wire31065)  &  wire35086 ) | ( (~ wire31066)  &  wire35086 ) ;
 assign wire35120 = ( (~ wire31065)  &  wire35087 ) | ( (~ wire31066)  &  wire35087 ) | ( (~ wire31065)  &  wire35088 ) | ( (~ wire31066)  &  wire35088 ) ;
 assign wire35121 = ( (~ wire31065)  &  wire35089 ) | ( (~ wire31066)  &  wire35089 ) | ( (~ wire31065)  &  wire35090 ) | ( (~ wire31066)  &  wire35090 ) ;
 assign wire35122 = ( (~ wire31065)  &  wire35091 ) | ( (~ wire31066)  &  wire35091 ) | ( (~ wire31065)  &  wire35092 ) | ( (~ wire31066)  &  wire35092 ) ;
 assign wire35123 = ( (~ wire31065)  &  wire35093 ) | ( (~ wire31066)  &  wire35093 ) | ( (~ wire31065)  &  wire35094 ) | ( (~ wire31066)  &  wire35094 ) ;
 assign wire35124 = ( (~ wire31065)  &  wire35095 ) | ( (~ wire31066)  &  wire35095 ) | ( (~ wire31065)  &  wire35096 ) | ( (~ wire31066)  &  wire35096 ) ;
 assign wire35125 = ( (~ wire31065)  &  wire35097 ) | ( (~ wire31066)  &  wire35097 ) | ( (~ wire31065)  &  wire35098 ) | ( (~ wire31066)  &  wire35098 ) ;
 assign wire35126 = ( ng10711  &  (~ wire31065) ) | ( ng10711  &  (~ wire31066) ) | ( (~ wire31065)  &  wire35099 ) | ( (~ wire31066)  &  wire35099 ) ;
 assign wire35127 = ( wire35100 ) | ( wire35101 ) | ( wire35102 ) | ( wire35103 ) ;
 assign wire35128 = ( wire35104 ) | ( wire35105 ) | ( wire35106 ) | ( wire35107 ) ;
 assign wire35135 = ( wire35128 ) | ( wire35127 ) ;
 assign wire35136 = ( wire35115 ) | ( wire35116 ) | ( wire35117 ) | ( wire35118 ) ;
 assign wire35137 = ( wire35119 ) | ( wire35120 ) | ( wire35121 ) | ( wire35122 ) ;
 assign wire35138 = ( wire35123 ) | ( wire35124 ) | ( wire35125 ) | ( wire35126 ) ;
 assign wire35143 = ( (~ ng11600)  &  (~ ng12941) ) | ( (~ ng12941)  &  (~ wire31795)  &  (~ wire31796) ) ;
 assign wire35144 = ( (~ ng28529)  &  (~ wire3748) ) | ( (~ ng28529)  &  wire35143 ) ;
 assign wire35146 = ( ng823  &  (~ ng1136)  &  ng2257 ) ;
 assign wire35147 = ( ng826  &  (~ ng1135)  &  ng2257 ) ;
 assign wire35148 = ( (~ ng1134)  &  ng853  &  ng2257 ) ;
 assign wire35150 = ( wire32303  &  (~ wire32323)  &  (~ wire32324) ) | ( wire32304  &  (~ wire32323)  &  (~ wire32324) ) ;
 assign wire35154 = ( (~ pg3229)  &  (~ ng12152)  &  ng12207 ) | ( pg3229  &  (~ ng12097)  &  (~ ng12207) ) ;
 assign wire35156 = ( ng1444  &  ng1439  &  ng1435 ) ;
 assign wire35157 = ( (~ ng17031)  &  ng1439 ) ;
 assign wire35159 = ( (~ ng17031)  &  ng1435 ) ;
 assign wire35160 = ( (~ ng25091)  &  wire33036 ) | ( (~ ng25091)  &  wire33037 ) ;
 assign wire35161 = ( ng1809  &  (~ ng823) ) | ( ng1809  &  (~ wire33053)  &  (~ wire33054) ) ;
 assign wire35162 = ( (~ ng11630)  &  (~ ng11666) ) | ( (~ ng11630)  &  wire32630 ) | ( (~ ng11630)  &  wire32631 ) ;
 assign wire35163 = ( (~ ng23518)  &  wire35162 ) | ( (~ ng23505)  &  wire35162 ) ;
 assign wire35164 = ( ng11630  &  (~ ng11666)  &  wire32630 ) | ( ng11630  &  (~ ng11666)  &  wire32631 ) ;
 assign wire35165 = ( (~ ng23526)  &  (~ wire32640)  &  (~ wire32641) ) ;
 assign wire35167 = ( wire32630  &  wire32650 ) | ( wire32631  &  wire32650 ) | ( wire32630  &  wire32651 ) | ( wire32631  &  wire32651 ) ;
 assign wire35169 = ( (~ wire32640)  &  (~ wire32641)  &  (~ wire32650)  &  (~ wire32651) ) ;
 assign wire35170 = ( wire32630  &  wire32650 ) | ( wire32631  &  wire32650 ) | ( wire32630  &  wire32651 ) | ( wire32631  &  wire32651 ) ;
 assign wire35171 = ( ng11675  &  ng11630  &  ng11666 ) | ( (~ ng11675)  &  (~ ng11630)  &  ng11666  &  wire3935 ) ;
 assign wire35172 = ( wire35171 ) | ( ng2257  &  ng23526  &  wire35167 ) ;
 assign wire35174 = ( wire5850 ) | ( wire5851 ) | ( wire35172 ) ;
 assign wire35175 = ( wire35174 ) | ( ng23505  &  ng27730  &  wire35165 ) ;
 assign wire35184 = ( (~ ng1312)  &  (~ ng1315)  &  ng1845 ) | ( (~ ng1312)  &  ng1865  &  ng1845 ) ;
 assign wire35186 = ( wire3049 ) | ( wire5831 ) | ( wire5832 ) | ( wire5833 ) ;
 assign wire35190 = ( (~ ng28584)  &  ng27585  &  wire33488 ) | ( (~ ng28584)  &  ng27585  &  wire33489 ) | ( (~ ng28584)  &  (~ ng27585)  &  (~ wire33488)  &  (~ wire33489) ) ;
 assign wire35191 = ( ng2180  &  ng27756 ) | ( ng25874  &  (~ ng27756)  &  (~ ng16693) ) ;
 assign wire35193 = ( (~ ng28584)  &  (~ ng26941)  &  wire33498 ) | ( (~ ng28584)  &  (~ ng26941)  &  wire33499 ) | ( (~ ng28584)  &  ng26941  &  (~ wire33498)  &  (~ wire33499) ) ;
 assign wire35194 = ( (~ ng11678)  &  (~ wire33498)  &  (~ wire33499)  &  wire33550 ) ;
 assign wire35195 = ( ng27585  &  (~ wire33805)  &  (~ wire33807)  &  wire35194 ) ;
 assign wire35197 = ( (~ wire33478)  &  (~ wire33479)  &  (~ wire33498)  &  (~ wire33499) ) ;
 assign wire35199 = ( (~ wire33478)  &  (~ wire33479)  &  wire33498 ) | ( (~ wire33478)  &  (~ wire33479)  &  wire33499 ) ;
 assign wire35200 = ( (~ wire33548)  &  (~ wire33549)  &  wire33550  &  wire35199 ) ;
 assign wire35202 = ( (~ ng28584)  &  ng26931  &  wire35195 ) | ( (~ ng28584)  &  ng26931  &  wire35197 ) ;
 assign wire35203 = ( (~ ng28584)  &  wire35200 ) | ( ng12836  &  (~ ng28584)  &  (~ ng26931) ) ;
 assign wire35208 = ( (~ wire33840)  &  (~ wire33841)  &  wire34421 ) | ( (~ wire33840)  &  (~ wire33841)  &  wire34422 ) ;
 assign wire35210 = ( wire5787 ) | ( ng2398  &  (~ ng823) ) ;
 assign wire35211 = ( wire35210 ) | ( (~ ng15950)  &  ng17151  &  (~ ng27892) ) ;
 assign wire35225 = ( (~ ng2639)  &  (~ ng1312)  &  (~ ng2564) ) | ( (~ ng2639)  &  (~ ng2564)  &  (~ ng2641) ) ;
 assign wire35226 = ( (~ ng2639)  &  (~ ng1312)  &  (~ ng1315) ) | ( (~ ng2639)  &  (~ ng1315)  &  (~ ng2641) ) ;
 assign wire35228 = ( wire3049 ) | ( wire5775 ) | ( wire35225 ) ;
 assign wire35229 = ( wire5780 ) | ( wire5781 ) | ( wire35226 ) ;
 assign wire35231 = ( (~ ng1312)  &  (~ ng2670)  &  (~ ng2676) ) ;
 assign wire35233 = ( (~ ng2670)  &  (~ ng2676)  &  (~ ng2673) ) ;
 assign wire35235 = ( (~ ng1315)  &  (~ ng2670)  &  (~ ng2673) ) ;
 assign wire35237 = ( (~ ng1309)  &  (~ ng2676)  &  (~ ng2673) ) ;
 assign wire35247 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2670) ) ;
 assign wire35250 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2676) ) ;
 assign wire35253 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2673) ) ;
 assign wire35263 = ( wire5751 ) | ( wire5752 ) | ( wire5753 ) | ( wire5754 ) ;
 assign wire35264 = ( wire5759 ) | ( wire5760 ) | ( wire5761 ) | ( wire5762 ) ;
 assign wire35265 = ( wire5763 ) | ( wire5765 ) | ( wire5766 ) | ( wire5768 ) ;
 assign wire35266 = ( wire5769 ) | ( wire5771 ) | ( wire5772 ) | ( wire5774 ) ;
 assign wire35270 = ( wire35228  &  wire35233 ) | ( wire35229  &  wire35233 ) | ( wire35228  &  wire35235 ) | ( wire35229  &  wire35235 ) ;
 assign wire35271 = ( wire35228  &  wire35237 ) | ( wire35229  &  wire35237 ) | ( wire35228  &  wire35247 ) | ( wire35229  &  wire35247 ) ;
 assign wire35272 = ( wire35228  &  wire35250 ) | ( wire35229  &  wire35250 ) | ( wire35228  &  wire35253 ) | ( wire35229  &  wire35253 ) ;
 assign wire35273 = ( wire3049 ) | ( wire35265 ) | ( wire35266 ) ;
 assign wire35274 = ( wire5755 ) | ( wire35263 ) | ( wire35264 ) | ( wire35270 ) ;
 assign wire35275 = ( wire35272 ) | ( wire35271 ) ;
 assign wire35277 = ( ng11896  &  wire3188 ) | ( wire3188  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35278 = ( wire5740 ) | ( ng21851  &  ng17139 ) | ( ng17139  &  wire34028 ) ;
 assign wire35280 = ( (~ ng28501)  &  (~ ng26902)  &  wire30947 ) | ( (~ ng28501)  &  (~ ng26902)  &  wire30948 ) | ( (~ ng28501)  &  ng26902  &  (~ wire30947)  &  (~ wire30948) ) ;
 assign wire35281 = ( wire32313  &  wire32429 ) | ( wire32314  &  wire32429 ) | ( wire32313  &  wire32430 ) | ( wire32314  &  wire32430 ) ;
 assign wire35284 = ( ng1807  &  (~ ng853) ) | ( ng1807  &  (~ wire33053)  &  (~ wire33054) ) ;
 assign wire35285 = ( ng2257  &  (~ ng12108)  &  ng18218  &  ng12057 ) | ( ng2257  &  ng12108  &  (~ ng18218)  &  (~ ng12057) ) ;
 assign wire35288 = ( ng2257  &  ng12108  &  (~ ng18218)  &  ng12057 ) | ( ng2257  &  (~ ng12108)  &  ng18218  &  (~ ng12057) ) ;
 assign wire35294 = ( (~ ng28584)  &  (~ ng26931)  &  wire33458 ) | ( (~ ng28584)  &  (~ ng26931)  &  wire33459 ) | ( (~ ng28584)  &  ng26931  &  (~ wire33458)  &  (~ wire33459) ) ;
 assign wire35295 = ( ng27756  &  (~ ng11917) ) | ( ng25874  &  (~ ng27756)  &  (~ ng16693) ) ;
 assign wire35304 = ( ng2151  &  (~ ng17031)  &  (~ ng23539) ) ;
 assign wire35306 = ( wire33850  &  wire33860 ) | ( wire33851  &  wire33860 ) | ( wire33850  &  wire33861 ) | ( wire33851  &  wire33861 ) ;
 assign wire35307 = ( wire5619 ) | ( ng2396  &  (~ ng853) ) ;
 assign wire35308 = ( wire35307 ) | ( (~ ng13165)  &  ng17151  &  (~ ng27892) ) ;
 assign wire35309 = ( ng11938  &  wire3174 ) | ( wire3174  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35310 = ( wire5606 ) | ( ng21851  &  ng17139 ) | ( ng17139  &  wire34028 ) ;
 assign wire35318 = ( (~ wire31795)  &  (~ wire31796)  &  (~ wire31815)  &  (~ wire31816) ) ;
 assign wire35319 = ( ng23511  &  wire35318 ) ;
 assign wire35320 = ( wire31795  &  (~ wire31815)  &  (~ wire31816) ) | ( wire31796  &  (~ wire31815)  &  (~ wire31816) ) ;
 assign wire35321 = ( (~ ng23511)  &  (~ wire31805)  &  (~ wire31806) ) ;
 assign wire35323 = ( wire31795  &  wire31815 ) | ( wire31796  &  wire31815 ) | ( wire31795  &  wire31816 ) | ( wire31796  &  wire31816 ) ;
 assign wire35325 = ( wire31795  &  wire31815 ) | ( wire31796  &  wire31815 ) | ( wire31795  &  wire31816 ) | ( wire31796  &  wire31816 ) ;
 assign wire35326 = ( (~ wire31805)  &  (~ wire31806)  &  (~ wire31815)  &  (~ wire31816) ) ;
 assign wire35327 = ( ng11663  &  ng11600  &  ng11647 ) | ( (~ ng11663)  &  (~ ng11600)  &  ng11647  &  wire3930 ) ;
 assign wire35328 = ( wire35327 ) | ( ng2257  &  ng23511  &  wire35323 ) ;
 assign wire35330 = ( wire5572 ) | ( wire5573 ) | ( wire35328 ) ;
 assign wire35331 = ( wire35330 ) | ( ng23489  &  ng27729  &  wire35321 ) ;
 assign wire35336 = ( wire32988  &  wire33008 ) | ( wire32989  &  wire33008 ) | ( wire32988  &  wire33009 ) | ( wire32989  &  wire33009 ) ;
 assign wire35337 = ( (~ ng1312)  &  (~ ng2040) ) | ( (~ ng2040)  &  (~ ng2010) ) ;
 assign wire35338 = ( (~ ng1312)  &  ng2040 ) | ( ng2040  &  (~ ng2010) ) ;
 assign wire35341 = ( (~ ng28584)  &  wire3314  &  wire33560 ) | ( (~ ng28584)  &  wire3314  &  wire33561 ) | ( (~ ng28584)  &  (~ wire3314)  &  (~ wire33560)  &  (~ wire33561) ) ;
 assign wire35345 = ( (~ ng1312)  &  ng633  &  (~ ng653) ) | ( (~ ng630)  &  ng633  &  (~ ng653) ) ;
 assign wire35346 = ( (~ ng1312)  &  ng653 ) | ( (~ ng630)  &  ng653 ) ;
 assign wire35347 = ( (~ wire32998)  &  (~ wire32999)  &  wire34927 ) | ( (~ wire32998)  &  (~ wire32999)  &  wire34928 ) ;
 assign wire35349 = ( pg3229  &  (~ wire32988)  &  (~ wire32989) ) ;
 assign wire35350 = ( wire5445 ) | ( (~ wire32998)  &  (~ wire32999)  &  wire35349 ) ;
 assign wire35352 = ( ng1808  &  (~ ng826) ) | ( ng1808  &  (~ wire33053)  &  (~ wire33054) ) ;
 assign wire35358 = ( ng1858  &  ng1859  &  ng1860 ) | ( ng1859  &  (~ ng1312)  &  ng1860 ) ;
 assign wire35362 = ( wire5422 ) | ( wire5423 ) | ( wire5424 ) | ( wire5425 ) ;
 assign wire35367 = ( ng11863  &  wire3174 ) | ( wire3174  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35368 = ( ng11831  &  wire3174 ) | ( wire3174  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35369 = ( ng536  &  wire3138 ) | ( ng21851  &  wire3138 ) | ( wire3138  &  wire34028 ) ;
 assign wire35371 = ( (~ ng2950)  &  ng2883 ) | ( ng2950  &  (~ ng2883) ) ;
 assign wire35375 = ( (~ ng28501)  &  wire3317  &  wire31048 ) | ( (~ ng28501)  &  wire3317  &  wire31049 ) | ( (~ ng28501)  &  (~ wire3317)  &  (~ wire31048)  &  (~ wire31049) ) ;
 assign wire35378 = ( (~ ng28501)  &  (~ ng26911)  &  wire30988 ) | ( (~ ng28501)  &  (~ ng26911)  &  wire30989 ) | ( (~ ng28501)  &  ng26911  &  (~ wire30988)  &  (~ wire30989) ) ;
 assign wire35379 = ( (~ ng23495)  &  (~ wire31271) ) | ( (~ ng23495)  &  (~ wire30977)  &  (~ wire30978) ) ;
 assign wire35380 = ( wire5341 ) | ( ng322  &  (~ ng826) ) ;
 assign wire35381 = ( wire35380 ) | ( ng826  &  (~ ng27834)  &  wire35379 ) ;
 assign wire35384 = ( (~ ng28529)  &  (~ ng26925)  &  wire31847 ) | ( (~ ng28529)  &  (~ ng26925)  &  wire31848 ) | ( (~ ng28529)  &  ng26925  &  (~ wire31847)  &  (~ wire31848) ) ;
 assign wire35390 = ( (~ ng28556)  &  ng26374  &  wire32610 ) | ( (~ ng28556)  &  ng26374  &  wire32611 ) | ( (~ ng28556)  &  (~ ng26374)  &  (~ wire32610)  &  (~ wire32611) ) ;
 assign wire35391 = ( ng1481  &  ng27751 ) | ( ng25853  &  (~ ng27751)  &  (~ ng16672) ) ;
 assign wire35394 = ( (~ ng28556)  &  (~ ng26928)  &  wire32681 ) | ( (~ ng28556)  &  (~ ng26928)  &  wire32682 ) | ( (~ ng28556)  &  ng26928  &  (~ wire32681)  &  (~ wire32682) ) ;
 assign wire35395 = ( (~ ng25099)  &  wire33889 ) | ( (~ ng25099)  &  wire33890 ) ;
 assign wire35396 = ( ng2503  &  (~ ng823) ) | ( ng2503  &  (~ wire33906)  &  (~ wire33907) ) ;
 assign wire35397 = ( (~ ng11653)  &  (~ ng11678) ) | ( (~ ng11653)  &  wire33528 ) | ( (~ ng11653)  &  wire33529 ) ;
 assign wire35405 = ( (~ ng2426)  &  (~ ng1315)  &  (~ ng2424) ) | ( (~ ng2426)  &  (~ ng2428)  &  (~ ng2424) ) ;
 assign wire35408 = ( wire3049 ) | ( wire5248 ) | ( wire35405 ) ;
 assign wire35409 = ( wire5251 ) | ( wire5252 ) | ( wire5253 ) | ( wire5254 ) ;
 assign wire35418 = ( wire3049 ) | ( wire5272 ) | ( wire5273 ) | ( wire5274 ) ;
 assign wire35419 = ( wire5275 ) | ( wire5276 ) | ( wire5277 ) | ( wire5278 ) ;
 assign wire35426 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2439) ) | ( (~ ng1312)  &  (~ ng2439)  &  (~ ng2443) ) ;
 assign wire35428 = ( wire3049 ) | ( wire5256 ) | ( wire5257 ) | ( wire5258 ) ;
 assign wire35429 = ( wire5261 ) | ( wire5262 ) | ( wire35426 ) ;
 assign wire35430 = ( wire34008  &  wire34018 ) | ( wire34009  &  wire34018 ) | ( wire34008  &  wire34019 ) | ( wire34009  &  wire34019 ) ;
 assign wire35437 = ( (~ ng2456)  &  (~ ng1315)  &  (~ ng2454) ) | ( (~ ng2456)  &  (~ ng2458)  &  (~ ng2454) ) ;
 assign wire35440 = ( wire3049 ) | ( wire5264 ) | ( wire35437 ) ;
 assign wire35441 = ( wire5267 ) | ( wire5268 ) | ( wire5269 ) | ( wire5270 ) ;
 assign wire35442 = ( (~ wire35428)  &  (~ wire35429)  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35444 = ( (~ wire33988)  &  (~ wire33989)  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35445 = ( (~ wire35408)  &  (~ wire35409)  &  (~ wire35428)  &  (~ wire35429) ) ;
 assign wire35446 = ( wire34008  &  wire35428 ) | ( wire34009  &  wire35428 ) | ( wire34008  &  wire35429 ) | ( wire34009  &  wire35429 ) ;
 assign wire35447 = ( (~ wire34018)  &  (~ wire34019)  &  wire35408 ) | ( (~ wire34018)  &  (~ wire34019)  &  wire35409 ) ;
 assign wire35448 = ( wire33998  &  (~ wire35440)  &  (~ wire35441) ) | ( wire33999  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35449 = ( (~ wire34018)  &  (~ wire34019)  &  wire35428 ) | ( (~ wire34018)  &  (~ wire34019)  &  wire35429 ) ;
 assign wire35450 = ( (~ wire33998)  &  (~ wire33999)  &  wire35418 ) | ( (~ wire33998)  &  (~ wire33999)  &  wire35419 ) ;
 assign wire35451 = ( wire34008  &  wire34018 ) | ( wire34009  &  wire34018 ) | ( wire34008  &  wire34019 ) | ( wire34009  &  wire34019 ) ;
 assign wire35454 = ( (~ wire34018)  &  (~ wire34019)  &  wire35440 ) | ( (~ wire34018)  &  (~ wire34019)  &  wire35441 ) ;
 assign wire35455 = ( (~ wire34008)  &  (~ wire34009)  &  wire35428 ) | ( (~ wire34008)  &  (~ wire34009)  &  wire35429 ) ;
 assign wire35456 = ( wire35444  &  wire35445 ) | ( wire35446  &  wire35447 ) ;
 assign wire35457 = ( wire35448  &  wire35449 ) | ( wire35450  &  wire35451 ) ;
 assign wire35458 = ( (~ ng12231)  &  ng10822  &  wire35454 ) | ( ng12231  &  (~ ng10822)  &  wire35455 ) ;
 assign wire35462 = ( wire5238 ) | ( wire5239 ) | ( wire35458 ) ;
 assign wire35463 = ( wire5244 ) | ( wire5245 ) | ( wire35456 ) | ( wire35457 ) ;
 assign wire35473 = ( (~ ng2661)  &  (~ ng2664)  &  (~ ng2667) ) ;
 assign wire35475 = ( (~ ng1315)  &  (~ ng2661)  &  (~ ng2664) ) ;
 assign wire35477 = ( (~ ng1312)  &  (~ ng2661)  &  (~ ng2667) ) ;
 assign wire35479 = ( (~ ng1309)  &  (~ ng2664)  &  (~ ng2667) ) ;
 assign wire35489 = ( (~ ng1312)  &  (~ ng1315)  &  (~ ng2661) ) ;
 assign wire35492 = ( (~ ng1312)  &  (~ ng1309)  &  (~ ng2667) ) ;
 assign wire35495 = ( (~ ng1315)  &  (~ ng1309)  &  (~ ng2664) ) ;
 assign wire35505 = ( wire5202 ) | ( wire5203 ) | ( wire5204 ) | ( wire5205 ) ;
 assign wire35506 = ( wire5210 ) | ( wire5211 ) | ( wire5212 ) | ( wire5213 ) ;
 assign wire35507 = ( wire5214 ) | ( wire5216 ) | ( wire5217 ) | ( wire5219 ) ;
 assign wire35508 = ( wire5220 ) | ( wire5222 ) | ( wire5223 ) | ( wire5225 ) ;
 assign wire35510 = ( wire35508 ) | ( wire35507 ) ;
 assign wire35512 = ( wire34948  &  wire35475 ) | ( wire34949  &  wire35475 ) | ( wire34948  &  wire35477 ) | ( wire34949  &  wire35477 ) ;
 assign wire35513 = ( wire34948  &  wire35479 ) | ( wire34949  &  wire35479 ) | ( wire34948  &  wire35489 ) | ( wire34949  &  wire35489 ) ;
 assign wire35514 = ( wire34948  &  wire35492 ) | ( wire34949  &  wire35492 ) | ( wire34948  &  wire35495 ) | ( wire34949  &  wire35495 ) ;
 assign wire35515 = ( wire5224 ) | ( wire35507 ) | ( wire35508 ) ;
 assign wire35516 = ( wire5206 ) | ( wire35505 ) | ( wire35506 ) | ( wire35512 ) ;
 assign wire35517 = ( wire35514 ) | ( wire35513 ) ;
 assign wire35519 = ( ng13055  &  (~ wire35273)  &  (~ wire35274)  &  (~ wire35275) ) ;
 assign wire35521 = ( wire33988  &  (~ wire33998)  &  (~ wire33999) ) | ( wire33989  &  (~ wire33998)  &  (~ wire33999) ) ;
 assign wire35522 = ( wire35428  &  (~ wire35440)  &  (~ wire35441) ) | ( wire35429  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35524 = ( wire33998  &  (~ wire35440)  &  (~ wire35441) ) | ( wire33999  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35525 = ( wire34018  &  (~ wire35428)  &  (~ wire35429) ) | ( wire34019  &  (~ wire35428)  &  (~ wire35429) ) ;
 assign wire35527 = ( wire34008  &  wire35440 ) | ( wire34009  &  wire35440 ) | ( wire34008  &  wire35441 ) | ( wire34009  &  wire35441 ) ;
 assign wire35528 = ( wire34018  &  (~ wire35428)  &  (~ wire35429) ) | ( wire34019  &  (~ wire35428)  &  (~ wire35429) ) ;
 assign wire35530 = ( wire34008  &  (~ wire34018)  &  (~ wire34019) ) | ( wire34009  &  (~ wire34018)  &  (~ wire34019) ) ;
 assign wire35532 = ( (~ wire34008)  &  (~ wire34009)  &  (~ wire35440)  &  (~ wire35441) ) ;
 assign wire35534 = ( (~ wire34018)  &  (~ wire34019)  &  wire35440 ) | ( (~ wire34018)  &  (~ wire34019)  &  wire35441 ) ;
 assign wire35536 = ( (~ wire33998)  &  (~ wire33999)  &  (~ wire34008)  &  (~ wire34009) ) ;
 assign wire35538 = ( wire34018  &  wire35428 ) | ( wire34019  &  wire35428 ) | ( wire34018  &  wire35429 ) | ( wire34019  &  wire35429 ) ;
 assign wire35539 = ( (~ wire33988)  &  (~ wire33989)  &  (~ wire35418)  &  (~ wire35419) ) ;
 assign wire35540 = ( wire33988  &  wire35418 ) | ( wire33989  &  wire35418 ) | ( wire33988  &  wire35419 ) | ( wire33989  &  wire35419 ) ;
 assign wire35541 = ( (~ wire33988)  &  (~ wire33989)  &  wire35440 ) | ( (~ wire33988)  &  (~ wire33989)  &  wire35441 ) ;
 assign wire35542 = ( wire33998  &  wire35418 ) | ( wire33999  &  wire35418 ) | ( wire33998  &  wire35419 ) | ( wire33999  &  wire35419 ) ;
 assign wire35543 = ( wire3352  &  wire35538 ) | ( wire3352  &  wire35539 ) ;
 assign wire35544 = ( ng10822  &  wire35541 ) | ( ng12231  &  (~ ng10822)  &  wire35540 ) ;
 assign wire35549 = ( wire5226 ) | ( wire5227 ) | ( wire5228 ) | ( wire5237 ) ;
 assign wire35550 = ( wire5229 ) | ( wire5230 ) | ( wire35543 ) | ( wire35544 ) ;
 assign wire35551 = ( wire35550 ) | ( wire35549 ) ;
 assign wire35553 = ( ng13055  &  wire35273 ) | ( ng13055  &  wire35274 ) | ( ng13055  &  wire35275 ) ;
 assign wire35554 = ( (~ wire35462)  &  (~ wire35463)  &  wire35553 ) ;
 assign wire35555 = ( wire5199 ) | ( (~ ng13055)  &  (~ wire33957)  &  (~ wire33958) ) ;
 assign wire35557 = ( ng2734  &  ng2746  &  ng2740 ) ;
 assign wire35564 = ( ng11830  &  wire3188 ) | ( wire3188  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35565 = ( ng12195  &  wire3188 ) | ( wire3188  &  (~ wire34048)  &  (~ wire34049) ) ;
 assign wire35566 = ( ng537  &  wire3138 ) | ( ng21851  &  wire3138 ) | ( wire3138  &  wire34028 ) ;
 assign wire35568 = ( ng1939 ) | ( pg1943 ) ;
 assign wire35574 = ( ng2082  &  (~ ng1315)  &  ng2083 ) | ( ng2082  &  ng2081  &  ng2083 ) ;
 assign wire35575 = ( ng2082  &  (~ ng1312)  &  (~ ng1315) ) | ( ng2082  &  (~ ng1312)  &  ng2081 ) ;
 assign wire35577 = ( wire3049 ) | ( wire5104 ) | ( wire35574 ) ;
 assign wire35578 = ( wire5109 ) | ( wire5110 ) | ( wire35575 ) ;
 assign wire35585 = ( (~ ng1312)  &  (~ ng1315)  &  ng2106 ) | ( (~ ng1315)  &  ng2107  &  ng2106 ) ;
 assign wire35587 = ( wire3049 ) | ( wire5160 ) | ( wire5161 ) | ( wire5162 ) ;
 assign wire35588 = ( wire5165 ) | ( wire5166 ) | ( wire35585 ) ;
 assign wire35597 = ( wire3049 ) | ( wire5152 ) | ( wire5153 ) | ( wire5154 ) ;
 assign wire35598 = ( wire5155 ) | ( wire5156 ) | ( wire5157 ) | ( wire5158 ) ;
 assign wire35607 = ( wire3049 ) | ( wire5144 ) | ( wire5145 ) | ( wire5146 ) ;
 assign wire35608 = ( wire5147 ) | ( wire5148 ) | ( wire5149 ) | ( wire5150 ) ;
 assign wire35614 = ( ng2090  &  (~ ng1309)  &  ng2092 ) | ( ng2090  &  ng2091  &  ng2092 ) ;
 assign wire35615 = ( ng2090  &  (~ ng1312)  &  ng2091 ) | ( (~ ng1312)  &  (~ ng1315)  &  ng2091 ) ;
 assign wire35617 = ( wire3049 ) | ( wire5136 ) | ( wire35614 ) ;
 assign wire35618 = ( wire5141 ) | ( wire5142 ) | ( wire35615 ) ;
 assign wire35627 = ( wire3049 ) | ( wire5128 ) | ( wire5129 ) | ( wire5130 ) ;
 assign wire35628 = ( wire5131 ) | ( wire5132 ) | ( wire5133 ) | ( wire5134 ) ;
 assign wire35634 = ( ng2104  &  ng2103  &  ng2102 ) | ( ng2103  &  (~ ng1312)  &  ng2102 ) ;
 assign wire35635 = ( ng2104  &  ng2103  &  (~ ng1315) ) | ( ng2103  &  (~ ng1312)  &  (~ ng1315) ) ;
 assign wire35637 = ( wire3049 ) | ( wire5120 ) | ( wire35634 ) ;
 assign wire35638 = ( wire5125 ) | ( wire5126 ) | ( wire35635 ) ;
 assign wire35645 = ( (~ ng1312)  &  (~ ng1315)  &  ng2085 ) | ( (~ ng1312)  &  ng2085  &  ng2084 ) ;
 assign wire35647 = ( wire3049 ) | ( wire5112 ) | ( wire5113 ) | ( wire5114 ) ;
 assign wire35648 = ( wire5117 ) | ( wire5118 ) | ( wire35645 ) ;
 assign wire35655 = ( (~ ng1312)  &  (~ ng1315)  &  ng2100 ) | ( (~ ng1312)  &  ng2100  &  ng2099 ) ;
 assign wire35657 = ( wire3049 ) | ( wire5168 ) | ( wire5169 ) | ( wire5170 ) ;
 assign wire35658 = ( wire5173 ) | ( wire5174 ) | ( wire35655 ) ;
 assign wire35664 = ( ng2094  &  (~ ng1315)  &  ng2095 ) | ( ng2094  &  ng2093  &  ng2095 ) ;
 assign wire35665 = ( ng2094  &  (~ ng1312)  &  (~ ng1315) ) | ( ng2094  &  (~ ng1312)  &  ng2093 ) ;
 assign wire35667 = ( wire3049 ) | ( wire5096 ) | ( wire35664 ) ;
 assign wire35668 = ( wire5101 ) | ( wire5102 ) | ( wire35665 ) ;
 assign wire35674 = ( ng2078  &  (~ ng1312)  &  ng2079 ) | ( ng2078  &  ng2080  &  ng2079 ) ;
 assign wire35677 = ( wire3049 ) | ( wire5088 ) | ( wire35674 ) ;
 assign wire35678 = ( wire5091 ) | ( wire5092 ) | ( wire5093 ) | ( wire5094 ) ;
 assign wire35687 = ( wire3049 ) | ( wire5069 ) | ( wire5070 ) | ( wire5071 ) ;
 assign wire35688 = ( wire5072 ) | ( wire5073 ) | ( wire5074 ) | ( wire5075 ) ;
 assign wire35690 = ( wire35577 ) | ( wire35578 ) | ( wire35587 ) | ( wire35588 ) ;
 assign wire35691 = ( wire35607 ) | ( wire35608 ) | ( (~ wire35597)  &  (~ wire35598) ) ;
 assign wire35692 = ( wire35627 ) | ( wire35628 ) | ( (~ wire35617)  &  (~ wire35618) ) ;
 assign wire35693 = ( wire35637 ) | ( wire35638 ) | ( wire35647 ) | ( wire35648 ) ;
 assign wire35694 = ( (~ wire35657)  &  (~ wire35658) ) | ( (~ wire35667)  &  (~ wire35668) ) ;
 assign wire35695 = ( wire35687 ) | ( wire35688 ) | ( (~ wire35677)  &  (~ wire35678) ) ;
 assign wire35698 = ( wire35695 ) | ( wire35694 ) ;
 assign wire35699 = ( wire35690 ) | ( wire35691 ) | ( wire35692 ) | ( wire35693 ) ;
 assign wire35701 = ( ng2114  &  ng2116  &  ng2115 ) ;
 assign wire35703 = ( (~ ng1315)  &  ng2116  &  ng2115 ) ;
 assign wire35705 = ( (~ ng1312)  &  ng2114  &  ng2115 ) ;
 assign wire35707 = ( (~ ng1309)  &  ng2114  &  ng2116 ) ;
 assign wire35708 = ( (~ ng1312)  &  (~ ng1315)  &  ng2115 ) ;
 assign wire35709 = ( (~ ng1312)  &  (~ ng1309)  &  ng2114 ) ;
 assign wire35710 = ( (~ ng1315)  &  (~ ng1309)  &  ng2116 ) ;
 assign wire35711 = ( (~ ng1880) ) | ( wire35698  &  wire35701 ) | ( wire35699  &  wire35701 ) ;
 assign wire35712 = ( wire35698  &  wire35703 ) | ( wire35699  &  wire35703 ) | ( wire35698  &  wire35705 ) | ( wire35699  &  wire35705 ) ;
 assign wire35713 = ( wire35698  &  wire35707 ) | ( wire35699  &  wire35707 ) | ( wire35698  &  wire35708 ) | ( wire35699  &  wire35708 ) ;
 assign wire35714 = ( wire35698  &  wire35709 ) | ( wire35699  &  wire35709 ) | ( wire35698  &  wire35710 ) | ( wire35699  &  wire35710 ) ;
 assign wire35716 = ( wire35713 ) | ( wire35712 ) ;
 assign wire35717 = ( wire5060 ) | ( wire35711 ) | ( wire35714 ) ;
 assign wire35721 = ( ng1315  &  (~ ng2808)  &  ng2574 ) ;
 assign wire35723 = ( (~ ng2809)  &  ng1309  &  ng2574 ) ;
 assign wire35725 = ( ng1312  &  (~ ng2810)  &  ng2574 ) ;
 assign wire35732 = ( (~ ng1312)  &  (~ ng1315)  &  ng2812 ) | ( (~ ng1315)  &  ng2812  &  ng2813 ) ;
 assign wire35734 = ( wire3049 ) | ( wire5029 ) | ( wire5030 ) | ( wire5031 ) ;
 assign wire35735 = ( wire5034 ) | ( wire5035 ) | ( wire35732 ) ;
 assign wire35737 = ( (~ wire34532)  &  (~ wire34533) ) | ( (~ wire34544)  &  (~ wire34545) ) ;
 assign wire35738 = ( wire34568 ) | ( wire34569 ) | ( wire34580 ) | ( wire34581 ) ;
 assign wire35739 = ( wire34520 ) | ( wire34521 ) | ( (~ wire34556)  &  (~ wire34557) ) ;
 assign wire35740 = ( wire34462 ) | ( wire34463 ) | ( (~ wire34508)  &  (~ wire34509) ) ;
 assign wire35741 = ( wire34484 ) | ( wire34485 ) | ( wire34496 ) | ( wire34497 ) ;
 assign wire35742 = ( wire35734 ) | ( wire35735 ) | ( (~ wire34472)  &  (~ wire34473) ) ;
 assign wire35745 = ( wire35742 ) | ( wire35741 ) ;
 assign wire35746 = ( wire35737 ) | ( wire35738 ) | ( wire35739 ) | ( wire35740 ) ;
 assign wire35747 = ( ng2631  &  (~ ng2584)  &  ng2574 ) ;
 assign wire35748 = ( ng2633 ) | ( pg2637 ) ;
 assign wire35750 = ( wire3198  &  wire35721 ) | ( wire3198  &  wire35723 ) | ( wire3198  &  wire35725 ) ;
 assign wire35751 = ( wire35750 ) | ( (~ wire35745)  &  (~ wire35746)  &  wire35747 ) ;
 assign wire35752 = ( ng12233  &  wire3183 ) | ( wire3183  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire35753 = ( ng30072  &  wire3137 ) | ( ng2605  &  wire3137 ) | ( wire3137  &  wire35748 ) ;
 assign wire35755 = ( ng3006  &  ng3002 ) ;
 assign wire35758 = ( (~ ng3006)  &  ng3080  &  ng2998  &  (~ ng3010) ) ;
 assign wire35759 = ( ng3013  &  ng3002  &  ng3024  &  (~ ng2993) ) ;
 assign wire35768 = ( (~ ng28501)  &  (~ ng25954)  &  wire31018 ) | ( (~ ng28501)  &  (~ ng25954)  &  wire31019 ) | ( (~ ng28501)  &  ng25954  &  (~ wire31018)  &  (~ wire31019) ) ;
 assign wire35769 = ( ng101  &  ng27738 ) | ( (~ ng16643)  &  ng25764  &  (~ ng27738) ) ;
 assign wire35770 = ( ng427  &  (~ ng826) ) | ( ng427  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire35771 = ( wire4983 ) | ( ng323  &  (~ ng823) ) ;
 assign wire35772 = ( wire35771 ) | ( ng823  &  (~ ng27834)  &  wire35379 ) ;
 assign wire35774 = ( (~ ng12755)  &  (~ ng26925)  &  (~ wire32142)  &  wire32155 ) ;
 assign wire35775 = ( (~ wire31857)  &  (~ wire31858)  &  (~ wire31877)  &  (~ wire31878) ) ;
 assign wire35776 = ( ng26925  &  wire35775 ) | ( wire32142  &  wire35775 ) | ( wire32155  &  wire35775 ) ;
 assign wire35777 = ( (~ ng12920)  &  ng26925 ) | ( (~ ng12920)  &  wire32142 ) | ( (~ ng12920)  &  wire32155 ) ;
 assign wire35778 = ( ng26925  &  (~ wire31877)  &  (~ wire31878) ) | ( (~ wire31877)  &  (~ wire31878)  &  wire32142 ) ;
 assign wire35779 = ( ng12755  &  (~ ng26925)  &  (~ wire32142)  &  (~ wire32155) ) ;
 assign wire35780 = ( (~ ng28529)  &  wire35776 ) | ( (~ ng28529)  &  wire35778 ) ;
 assign wire35781 = ( (~ ng28529)  &  wire35779 ) | ( (~ ng28529)  &  ng16655  &  wire35774 ) ;
 assign wire35790 = ( (~ ng1312)  &  ng1319 ) | ( (~ ng1316)  &  ng1319 ) ;
 assign wire35791 = ( (~ ng1339)  &  wire35790 ) | ( (~ ng1319)  &  wire35790 ) | ( (~ wire32567)  &  wire35790 ) ;
 assign wire35792 = ( (~ ng1312)  &  ng1339 ) | ( ng1339  &  (~ ng1316) ) ;
 assign wire35794 = ( (~ ng12971)  &  ng11666  &  (~ ng12828) ) | ( (~ ng12971)  &  (~ ng12828)  &  (~ wire32652) ) | ( (~ ng12971)  &  (~ ng11666)  &  ng12828  &  wire32652 ) ;
 assign wire35795 = ( ng25853  &  (~ ng27751)  &  (~ ng16672) ) | ( (~ ng25853)  &  (~ ng27751)  &  wire35794 ) ;
 assign wire35796 = ( (~ ng28556)  &  (~ ng12971)  &  ng26918 ) | ( (~ ng28556)  &  ng12971  &  (~ wire3190)  &  (~ ng26918) ) ;
 assign wire35798 = ( ng2501  &  (~ ng853) ) | ( ng2501  &  (~ wire33906)  &  (~ wire33907) ) ;
 assign wire35799 = ( wire34008  &  wire34018 ) | ( wire34009  &  wire34018 ) | ( wire34008  &  wire34019 ) | ( wire34009  &  wire34019 ) ;
 assign wire35802 = ( pg3229  &  (~ ng557)  &  (~ ng510)  &  ng538 ) ;
 assign wire35806 = ( (~ pg3229)  &  (~ ng557)  &  (~ ng510)  &  ng541 ) ;
 assign wire35812 = ( wire4889 ) | ( wire4888 ) ;
 assign wire35814 = ( wire35812 ) | ( ng557  &  (~ ng26096)  &  ng26107 ) | ( ng557  &  ng26096  &  (~ ng26107) ) ;
 assign wire35816 = ( ng1245 ) | ( pg1249 ) ;
 assign wire35819 = ( (~ pg3229)  &  (~ ng1196)  &  ng1227  &  (~ ng1243) ) ;
 assign wire35823 = ( pg3229  &  ng1224  &  (~ ng1196)  &  (~ ng1243) ) ;
 assign wire35830 = ( ng1425  &  ng1423  &  ng1424 ) | ( ng1423  &  (~ ng1312)  &  ng1424 ) ;
 assign wire35833 = ( wire3049 ) | ( wire4869 ) | ( wire35830 ) ;
 assign wire35834 = ( wire4872 ) | ( wire4873 ) | ( wire4874 ) | ( wire4875 ) ;
 assign wire35836 = ( wire34815 ) | ( wire34816 ) | ( wire34839 ) | ( wire34840 ) ;
 assign wire35837 = ( wire34757 ) | ( wire34758 ) | ( wire34803 ) | ( wire34804 ) ;
 assign wire35838 = ( (~ wire34863)  &  (~ wire34864) ) | ( (~ wire34875)  &  (~ wire34876) ) ;
 assign wire35839 = ( wire34851 ) | ( wire34852 ) | ( (~ wire34827)  &  (~ wire34828) ) ;
 assign wire35840 = ( wire34791 ) | ( wire34792 ) | ( (~ wire34779)  &  (~ wire34780) ) ;
 assign wire35841 = ( wire35833 ) | ( wire35834 ) | ( (~ wire34767)  &  (~ wire34768) ) ;
 assign wire35844 = ( wire35841 ) | ( wire35840 ) ;
 assign wire35845 = ( wire35836 ) | ( wire35837 ) | ( wire35838 ) | ( wire35839 ) ;
 assign wire35860 = ( (~ ng27113)  &  wire3143  &  wire35819 ) | ( (~ ng27113)  &  wire3143  &  wire35823 ) ;
 assign wire35862 = ( wire35860 ) | ( ng1243  &  (~ ng27824)  &  ng27811 ) | ( ng1243  &  ng27824  &  (~ ng27811) ) ;
 assign wire35864 = ( ng12184  &  wire3189 ) | ( wire3189  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire35866 = ( (~ ng3006)  &  ng3080  &  ng2998  &  ng2993 ) ;
 assign wire35867 = ( ng3006  &  (~ ng3080) ) | ( ng3006  &  (~ ng2998) ) | ( ng3006  &  (~ ng2993) ) ;
 assign wire35872 = ( ng2896  &  (~ ng2892)  &  (~ ng20825) ) ;
 assign wire35873 = ( ng2892  &  (~ ng2950) ) | ( ng2892  &  (~ wire35033) ) ;
 assign wire35874 = ( ng428  &  (~ ng823) ) | ( ng428  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire35875 = ( (~ ng13378)  &  (~ ng11624) ) | ( (~ ng13378)  &  wire30957 ) | ( (~ ng13378)  &  wire30958 ) ;
 assign wire35876 = ( (~ ng23486)  &  wire35875 ) | ( (~ ng23478)  &  wire35875 ) ;
 assign wire35877 = ( ng13378  &  (~ ng11624)  &  wire30957 ) | ( ng13378  &  (~ ng11624)  &  wire30958 ) ;
 assign wire35884 = ( (~ ng1312)  &  (~ ng1315)  &  ng464 ) | ( (~ ng1312)  &  ng484  &  ng464 ) ;
 assign wire35886 = ( wire3049 ) | ( wire4770 ) | ( wire4771 ) | ( wire4772 ) ;
 assign wire35895 = ( ng771  &  (~ ng767) ) ;
 assign wire35900 = ( (~ ng28556)  &  ng27582  &  wire32671 ) | ( (~ ng28556)  &  ng27582  &  wire32672 ) | ( (~ ng28556)  &  (~ ng27582)  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire35901 = ( ng1486  &  ng27751 ) | ( ng25853  &  (~ ng27751)  &  (~ ng16672) ) ;
 assign wire35902 = ( (~ wire32600)  &  (~ wire32601)  &  wire32661 ) | ( (~ wire32600)  &  (~ wire32601)  &  wire32662 ) ;
 assign wire35903 = ( (~ wire32650)  &  (~ wire32651)  &  wire32652  &  wire35902 ) ;
 assign wire35904 = ( ng27582  &  (~ wire32952)  &  wire35903 ) ;
 assign wire35905 = ( (~ wire32600)  &  (~ wire32601)  &  (~ wire32661)  &  (~ wire32662) ) ;
 assign wire35906 = ( wire32650  &  wire35905 ) | ( wire32651  &  wire35905 ) | ( (~ wire32652)  &  wire35905 ) ;
 assign wire35907 = ( (~ ng12930)  &  (~ wire32650)  &  (~ wire32651)  &  wire32652 ) ;
 assign wire35908 = ( (~ ng27582)  &  wire35907 ) | ( wire32952  &  wire35907 ) | ( wire32954  &  wire35907 ) ;
 assign wire35909 = ( (~ ng27582)  &  (~ wire32661)  &  (~ wire32662) ) | ( (~ wire32661)  &  (~ wire32662)  &  wire32952 ) ;
 assign wire35910 = ( ng12930  &  ng27582  &  (~ wire32952)  &  (~ wire32954) ) ;
 assign wire35911 = ( (~ ng28556)  &  wire35904 ) | ( (~ ng28556)  &  wire35906 ) ;
 assign wire35912 = ( (~ ng28556)  &  wire35908 ) | ( (~ ng28556)  &  wire35909 ) ;
 assign wire35913 = ( ng1496  &  ng27751 ) | ( (~ ng25853)  &  (~ ng27751)  &  wire35910 ) ;
 assign wire35915 = ( ng1680  &  ng823 ) ;
 assign wire35917 = ( (~ ng1680)  &  (~ ng1679) ) | ( (~ ng823)  &  ng1680  &  ng1686 ) ;
 assign wire35918 = ( ng823  &  ng2374 ) ;
 assign wire35920 = ( (~ ng2374)  &  (~ ng2373) ) | ( ng2374  &  ng2380  &  (~ ng823) ) ;
 assign wire35927 = ( (~ ng1312)  &  (~ ng1315)  &  ng2539 ) | ( (~ ng1312)  &  ng2559  &  ng2539 ) ;
 assign wire35929 = ( wire3049 ) | ( wire4690 ) | ( wire4691 ) | ( wire4692 ) ;
 assign wire35931 = ( ng13055  &  wire35273 ) | ( ng13055  &  wire35274 ) | ( ng13055  &  wire35275 ) ;
 assign wire35932 = ( (~ wire35515)  &  (~ wire35516)  &  (~ wire35517)  &  wire35931 ) ;
 assign wire35933 = ( ng13055  &  wire35515 ) | ( ng13055  &  wire35516 ) | ( ng13055  &  wire35517 ) ;
 assign wire35934 = ( wire35462  &  wire35933 ) | ( wire35463  &  wire35933 ) ;
 assign wire35937 = ( ng1420  &  ng1421  &  ng1422 ) ;
 assign wire35939 = ( (~ ng1315)  &  ng1421  &  ng1422 ) ;
 assign wire35941 = ( ng1420  &  (~ ng1309)  &  ng1422 ) ;
 assign wire35943 = ( (~ ng1312)  &  ng1420  &  ng1421 ) ;
 assign wire35944 = ( (~ ng1312)  &  (~ ng1315)  &  ng1421 ) ;
 assign wire35945 = ( (~ ng1312)  &  ng1420  &  (~ ng1309) ) ;
 assign wire35946 = ( (~ ng1315)  &  (~ ng1309)  &  ng1422 ) ;
 assign wire35947 = ( (~ ng1186) ) | ( wire35844  &  wire35937 ) | ( wire35845  &  wire35937 ) ;
 assign wire35948 = ( wire35844  &  wire35939 ) | ( wire35845  &  wire35939 ) | ( wire35844  &  wire35941 ) | ( wire35845  &  wire35941 ) ;
 assign wire35949 = ( wire35844  &  wire35943 ) | ( wire35845  &  wire35943 ) | ( wire35844  &  wire35944 ) | ( wire35845  &  wire35944 ) ;
 assign wire35950 = ( wire35844  &  wire35945 ) | ( wire35845  &  wire35945 ) | ( wire35844  &  wire35946 ) | ( wire35845  &  wire35946 ) ;
 assign wire35952 = ( wire35949 ) | ( wire35948 ) ;
 assign wire35953 = ( wire4673 ) | ( wire35947 ) | ( wire35950 ) ;
 assign wire35957 = ( ng12306  &  wire3183 ) | ( wire3183  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire35961 = ( ng426  &  (~ ng853) ) | ( ng426  &  (~ wire31382)  &  (~ wire31383) ) ;
 assign wire35964 = ( (~ ng2160)  &  (~ wire33560)  &  (~ wire33561) ) ;
 assign wire35965 = ( (~ ng2160)  &  (~ wire33560)  &  (~ wire33561) ) ;
 assign wire35966 = ( ng2160  &  wire33560 ) | ( ng2160  &  wire33561 ) ;
 assign wire35967 = ( ng2160  &  wire33560 ) | ( ng2160  &  wire33561 ) ;
 assign wire35968 = ( (~ ng2142)  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire35969 = ( (~ ng2142)  &  (~ wire33518)  &  (~ wire33519) ) ;
 assign wire35970 = ( ng2142  &  wire33518 ) | ( ng2142  &  wire33519 ) ;
 assign wire35971 = ( ng2142  &  wire33518 ) | ( ng2142  &  wire33519 ) ;
 assign wire35972 = ( (~ ng2156)  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign wire35973 = ( (~ ng2156)  &  (~ wire33508)  &  (~ wire33509) ) ;
 assign wire35974 = ( ng2156  &  wire33508 ) | ( ng2156  &  wire33509 ) ;
 assign wire35975 = ( ng2156  &  wire33508 ) | ( ng2156  &  wire33509 ) ;
 assign wire35976 = ( (~ ng2133)  &  (~ wire33498)  &  (~ wire33499) ) ;
 assign wire35977 = ( (~ ng2133)  &  (~ wire33498)  &  (~ wire33499) ) ;
 assign wire35978 = ( ng2133  &  wire33498 ) | ( ng2133  &  wire33499 ) ;
 assign wire35979 = ( ng2133  &  wire33498 ) | ( ng2133  &  wire33499 ) ;
 assign wire35980 = ( (~ ng2147)  &  (~ wire33488)  &  (~ wire33489) ) ;
 assign wire35981 = ( ng2147  &  wire33488 ) | ( ng2147  &  wire33489 ) ;
 assign wire35982 = ( (~ ng2151)  &  (~ wire33448)  &  (~ wire33449) ) ;
 assign wire35983 = ( ng2151  &  wire33448 ) | ( ng2151  &  wire33449 ) ;
 assign wire35984 = ( (~ ng2129)  &  (~ wire33478)  &  (~ wire33479) ) ;
 assign wire35985 = ( ng2129  &  wire33478 ) | ( ng2129  &  wire33479 ) ;
 assign wire35986 = ( (~ ng2138)  &  (~ wire33468)  &  (~ wire33469) ) ;
 assign wire35987 = ( ng2138  &  wire33468 ) | ( ng2138  &  wire33469 ) ;
 assign wire35988 = ( (~ ng2124)  &  (~ wire33458)  &  (~ wire33459) ) ;
 assign wire35989 = ( ng2124  &  wire33458 ) | ( ng2124  &  wire33459 ) ;
 assign wire35990 = ( (~ ng2120)  &  (~ wire33438)  &  (~ wire33439) ) ;
 assign wire35991 = ( ng2120  &  wire33438 ) | ( ng2120  &  wire33439 ) ;
 assign wire35992 = ( (~ ng2147)  &  (~ wire33488)  &  (~ wire33489) ) ;
 assign wire35993 = ( ng2147  &  wire33488 ) | ( ng2147  &  wire33489 ) ;
 assign wire35994 = ( (~ ng2151)  &  (~ wire33448)  &  (~ wire33449) ) ;
 assign wire35995 = ( ng2151  &  wire33448 ) | ( ng2151  &  wire33449 ) ;
 assign wire35996 = ( (~ ng2129)  &  (~ wire33478)  &  (~ wire33479) ) ;
 assign wire35997 = ( ng2129  &  wire33478 ) | ( ng2129  &  wire33479 ) ;
 assign wire35998 = ( (~ ng2138)  &  (~ wire33468)  &  (~ wire33469) ) ;
 assign wire35999 = ( ng2138  &  wire33468 ) | ( ng2138  &  wire33469 ) ;
 assign wire36000 = ( (~ ng2124)  &  (~ wire33458)  &  (~ wire33459) ) ;
 assign wire36001 = ( ng2124  &  wire33458 ) | ( ng2124  &  wire33459 ) ;
 assign wire36002 = ( (~ ng2120)  &  (~ wire33438)  &  (~ wire33439) ) ;
 assign wire36003 = ( ng2120  &  wire33438 ) | ( ng2120  &  wire33439 ) ;
 assign wire36004 = ( (~ ng11687)  &  wire35964 ) | ( (~ ng11653)  &  wire35964 ) | ( (~ ng11678)  &  wire35964 ) | ( (~ ng11687)  &  ng11653  &  (~ ng11678) ) ;
 assign wire36005 = ( (~ ng11678)  &  wire35966 ) | ( (~ wire33551)  &  wire35966 ) | ( (~ ng11678)  &  wire35968 ) | ( (~ wire33551)  &  wire35968 ) ;
 assign wire36006 = ( (~ ng11678)  &  wire35970 ) | ( (~ wire33551)  &  wire35970 ) | ( (~ ng11678)  &  wire35972 ) | ( (~ wire33551)  &  wire35972 ) ;
 assign wire36007 = ( (~ ng11678)  &  wire35974 ) | ( (~ wire33551)  &  wire35974 ) | ( (~ ng11678)  &  wire35976 ) | ( (~ wire33551)  &  wire35976 ) ;
 assign wire36008 = ( (~ ng11678)  &  wire35978 ) | ( (~ wire33551)  &  wire35978 ) | ( (~ ng11678)  &  wire35980 ) | ( (~ wire33551)  &  wire35980 ) ;
 assign wire36009 = ( (~ ng11678)  &  wire35981 ) | ( (~ wire33551)  &  wire35981 ) | ( (~ ng11678)  &  wire35982 ) | ( (~ wire33551)  &  wire35982 ) ;
 assign wire36010 = ( (~ ng11678)  &  wire35983 ) | ( (~ wire33551)  &  wire35983 ) | ( (~ ng11678)  &  wire35984 ) | ( (~ wire33551)  &  wire35984 ) ;
 assign wire36011 = ( (~ ng11678)  &  wire35985 ) | ( (~ wire33551)  &  wire35985 ) | ( (~ ng11678)  &  wire35986 ) | ( (~ wire33551)  &  wire35986 ) ;
 assign wire36012 = ( (~ ng11678)  &  wire35987 ) | ( (~ wire33551)  &  wire35987 ) | ( (~ ng11678)  &  wire35988 ) | ( (~ wire33551)  &  wire35988 ) ;
 assign wire36013 = ( (~ ng11678)  &  wire35989 ) | ( (~ wire33551)  &  wire35989 ) | ( (~ ng11678)  &  wire35990 ) | ( (~ wire33551)  &  wire35990 ) ;
 assign wire36014 = ( (~ ng11678)  &  ng10711 ) | ( ng10711  &  (~ wire33551) ) | ( (~ ng11678)  &  wire35991 ) | ( (~ wire33551)  &  wire35991 ) ;
 assign wire36019 = ( wire36013 ) | ( wire36012 ) ;
 assign wire36020 = ( wire36014 ) | ( (~ wire33578)  &  wire35965 ) | ( (~ wire33579)  &  wire35965 ) ;
 assign wire36021 = ( (~ wire33578)  &  wire35967 ) | ( (~ wire33579)  &  wire35967 ) | ( (~ wire33578)  &  wire35969 ) | ( (~ wire33579)  &  wire35969 ) ;
 assign wire36022 = ( (~ wire33578)  &  wire35971 ) | ( (~ wire33579)  &  wire35971 ) | ( (~ wire33578)  &  wire35973 ) | ( (~ wire33579)  &  wire35973 ) ;
 assign wire36023 = ( (~ wire33578)  &  wire35975 ) | ( (~ wire33579)  &  wire35975 ) | ( (~ wire33578)  &  wire35977 ) | ( (~ wire33579)  &  wire35977 ) ;
 assign wire36024 = ( (~ wire33578)  &  wire35979 ) | ( (~ wire33579)  &  wire35979 ) | ( (~ wire33578)  &  wire35992 ) | ( (~ wire33579)  &  wire35992 ) ;
 assign wire36025 = ( (~ wire33578)  &  wire35993 ) | ( (~ wire33579)  &  wire35993 ) | ( (~ wire33578)  &  wire35994 ) | ( (~ wire33579)  &  wire35994 ) ;
 assign wire36026 = ( (~ wire33578)  &  wire35995 ) | ( (~ wire33579)  &  wire35995 ) | ( (~ wire33578)  &  wire35996 ) | ( (~ wire33579)  &  wire35996 ) ;
 assign wire36027 = ( (~ wire33578)  &  wire35997 ) | ( (~ wire33579)  &  wire35997 ) | ( (~ wire33578)  &  wire35998 ) | ( (~ wire33579)  &  wire35998 ) ;
 assign wire36028 = ( (~ wire33578)  &  wire35999 ) | ( (~ wire33579)  &  wire35999 ) | ( (~ wire33578)  &  wire36000 ) | ( (~ wire33579)  &  wire36000 ) ;
 assign wire36029 = ( (~ wire33578)  &  wire36001 ) | ( (~ wire33579)  &  wire36001 ) | ( (~ wire33578)  &  wire36002 ) | ( (~ wire33579)  &  wire36002 ) ;
 assign wire36030 = ( ng10711  &  (~ wire33578) ) | ( ng10711  &  (~ wire33579) ) | ( (~ wire33578)  &  wire36003 ) | ( (~ wire33579)  &  wire36003 ) ;
 assign wire36031 = ( wire36004 ) | ( wire36005 ) | ( wire36006 ) | ( wire36007 ) ;
 assign wire36032 = ( wire36008 ) | ( wire36009 ) | ( wire36010 ) | ( wire36011 ) ;
 assign wire36039 = ( wire36032 ) | ( wire36031 ) ;
 assign wire36040 = ( wire36019 ) | ( wire36020 ) | ( wire36021 ) | ( wire36022 ) ;
 assign wire36041 = ( wire36023 ) | ( wire36024 ) | ( wire36025 ) | ( wire36026 ) ;
 assign wire36042 = ( wire36027 ) | ( wire36028 ) | ( wire36029 ) | ( wire36030 ) ;
 assign wire36045 = ( (~ ng1886)  &  ng1312 ) ;
 assign wire36047 = ( ng1886  &  ng1887 ) | ( pg16399  &  (~ ng1312)  &  (~ ng1886) ) ;
 assign wire36048 = ( (~ ng2580)  &  ng1312 ) ;
 assign wire36050 = ( ng2580  &  ng2581 ) | ( pg16437  &  (~ ng1312)  &  (~ ng2580) ) ;
 assign wire36054 = ( ng12271  &  wire3189 ) | ( wire3189  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36055 = ( ng30072  &  wire3137 ) | ( ng2604  &  wire3137 ) | ( wire3137  &  wire35748 ) ;
 assign wire36057 = ( (~ ng2993)  &  ng3080 ) ;
 assign wire36058 = ( ng2993  &  (~ ng3080) ) ;
 assign wire36064 = ( (~ ng28501)  &  ng27563  &  wire30927 ) | ( (~ ng28501)  &  ng27563  &  wire30928 ) | ( (~ ng28501)  &  (~ ng27563)  &  (~ wire30927)  &  (~ wire30928) ) ;
 assign wire36065 = ( ng109  &  ng27738 ) | ( (~ ng16643)  &  ng25764  &  (~ ng27738) ) ;
 assign wire36077 = ( (~ ng1315)  &  ng488  &  ng486 ) | ( ng488  &  ng487  &  ng486 ) ;
 assign wire36078 = ( (~ ng1312)  &  (~ ng1315)  &  ng488 ) | ( (~ ng1312)  &  ng488  &  ng487 ) ;
 assign wire36081 = ( wire4425 ) | ( wire4426 ) | ( wire36078 ) ;
 assign wire36082 = ( ng13055  &  wire34164 ) | ( ng13055  &  wire34165 ) | ( ng13055  &  wire34166 ) ;
 assign wire36083 = ( (~ wire34243)  &  (~ wire34244)  &  wire36082 ) ;
 assign wire36084 = ( ng13055  &  (~ wire34164)  &  (~ wire34165)  &  (~ wire34166) ) ;
 assign wire36086 = ( wire4416 ) | ( (~ ng13055)  &  (~ wire31449)  &  (~ wire31450) ) ;
 assign wire36089 = ( (~ wire31837)  &  (~ wire31838)  &  wire31897 ) | ( (~ wire31837)  &  (~ wire31838)  &  wire31898 ) ;
 assign wire36090 = ( (~ ng12820)  &  (~ ng25958)  &  ng16655  &  wire36089 ) | ( ng12820  &  (~ ng25958)  &  (~ ng16655)  &  wire36089 ) ;
 assign wire36091 = ( (~ wire31837)  &  (~ wire31838)  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign wire36093 = ( wire31837  &  (~ wire31897)  &  (~ wire31898) ) | ( wire31838  &  (~ wire31897)  &  (~ wire31898) ) ;
 assign wire36095 = ( ng25958  &  (~ ng12852) ) | ( ng12820  &  ng16655  &  (~ ng12852) ) | ( (~ ng12820)  &  (~ ng16655)  &  (~ ng12852) ) ;
 assign wire36096 = ( (~ ng28529)  &  ng12968  &  (~ ng26925) ) | ( (~ ng28529)  &  ng26925  &  wire36091 ) ;
 assign wire36097 = ( (~ ng16655)  &  ng25818  &  (~ ng27743) ) | ( (~ ng25818)  &  (~ ng27743)  &  wire36095 ) ;
 assign wire36098 = ( (~ ng28529)  &  ng16655  &  wire36090 ) | ( (~ ng28529)  &  ng16655  &  wire36093 ) ;
 assign wire36109 = ( wire3046 ) | ( wire4380 ) | ( wire4381 ) | ( wire4382 ) ;
 assign wire36110 = ( wire4383 ) | ( wire4384 ) | ( wire4385 ) | ( wire4386 ) ;
 assign wire36111 = ( (~ wire32187)  &  (~ wire32188)  &  wire36109 ) | ( (~ wire32187)  &  (~ wire32188)  &  wire36110 ) ;
 assign wire36115 = ( (~ pg3229)  &  (~ ng12043)  &  ng12090 ) | ( pg3229  &  (~ ng11987)  &  (~ ng12090) ) ;
 assign wire36116 = ( wire31815  &  (~ wire31828) ) | ( wire31816  &  (~ wire31828) ) ;
 assign wire36119 = ( (~ ng11663)  &  ng11647 ) | ( (~ ng2257)  &  (~ ng11600)  &  ng11647 ) | ( (~ ng11663)  &  ng11600  &  (~ ng11647) ) ;
 assign wire36120 = ( wire36119 ) | ( (~ ng23502)  &  wire36116 ) | ( (~ ng23489)  &  wire36116 ) ;
 assign wire36121 = ( (~ wire8594)  &  (~ wire31795)  &  (~ wire31796)  &  (~ wire32093) ) ;
 assign wire36122 = ( (~ wire8594)  &  wire31795  &  (~ wire32093) ) | ( (~ wire8594)  &  wire31796  &  (~ wire32093) ) ;
 assign wire36131 = ( wire3049 ) | ( wire4345 ) | ( wire4346 ) | ( wire4347 ) ;
 assign wire36132 = ( wire4348 ) | ( wire4349 ) | ( wire4350 ) | ( wire4351 ) ;
 assign wire36135 = ( (~ ng28556)  &  (~ ng25964)  &  wire32691 ) | ( (~ ng28556)  &  (~ ng25964)  &  wire32692 ) | ( (~ ng28556)  &  ng25964  &  (~ wire32691)  &  (~ wire32692) ) ;
 assign wire36136 = ( ng1476  &  ng27751 ) | ( ng25853  &  (~ ng27751)  &  (~ ng16672) ) ;
 assign wire36139 = ( (~ wire33538)  &  (~ wire33539)  &  (~ wire33548)  &  (~ wire33549) ) ;
 assign wire36140 = ( (~ ng23537)  &  wire36139 ) ;
 assign wire36142 = ( ng2257  &  wire33528 ) | ( ng2257  &  wire33529 ) ;
 assign wire36144 = ( (~ ng23537)  &  wire3236 ) | ( ng11678  &  wire3236  &  wire33792 ) ;
 assign wire36145 = ( (~ wire33538)  &  (~ wire33539)  &  (~ wire33548)  &  (~ wire33549) ) ;
 assign wire36146 = ( wire33528  &  wire33548 ) | ( wire33529  &  wire33548 ) | ( wire33528  &  wire33549 ) | ( wire33529  &  wire33549 ) ;
 assign wire36147 = ( ng11687  &  ng11653  &  ng11678 ) | ( (~ ng11687)  &  (~ ng11653)  &  ng11678  &  wire3925 ) ;
 assign wire36148 = ( wire36147 ) | ( ng23537  &  ng11678  &  wire36142 ) ;
 assign wire36150 = ( wire4305 ) | ( wire4306 ) | ( wire36148 ) ;
 assign wire36151 = ( wire36150 ) | ( ng27892  &  wire36144 ) ;
 assign wire36160 = ( (~ ng1312)  &  (~ ng1315)  &  ng2563 ) | ( (~ ng1312)  &  ng2563  &  ng2562 ) ;
 assign wire36162 = ( wire3049 ) | ( wire4286 ) | ( wire4287 ) | ( wire4288 ) ;
 assign wire36170 = ( wire3277 ) | ( wire4265 ) ;
 assign wire36171 = ( ng12008  &  wire3183 ) | ( wire3183  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36172 = ( ng11965  &  wire3183 ) | ( wire3183  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36173 = ( ng2610  &  wire3137 ) | ( ng30072  &  wire3137 ) | ( wire3137  &  wire35748 ) ;
 assign wire36175 = ( (~ pg3234)  &  ng3028 ) | ( (~ pg3234)  &  (~ ng3032) ) ;
 assign wire36176 = ( wire4250 ) | ( (~ pg3234)  &  ng3028 ) | ( (~ pg3234)  &  (~ ng3032) ) ;
 assign wire36177 = ( ng3018  &  (~ wire35758) ) | ( ng3018  &  (~ wire35759) ) | ( (~ ng3018)  &  wire35758  &  wire35759 ) ;
 assign wire36183 = ( (~ ng1312)  &  ng2746  &  (~ ng2740) ) | ( (~ ng2704)  &  ng2746  &  (~ ng2740) ) ;
 assign wire36184 = ( (~ ng1312)  &  ng2740 ) | ( (~ ng2704)  &  ng2740 ) ;
 assign wire36188 = ( ng11964  &  wire3189 ) | ( wire3189  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36189 = ( ng12329  &  wire3189 ) | ( wire3189  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36190 = ( ng30072  &  wire3137 ) | ( ng2611  &  wire3137 ) | ( wire3137  &  wire35748 ) ;
 assign wire36192 = ( wire4076 ) | ( (~ ng853)  &  ng321 ) ;
 assign wire36193 = ( wire36192 ) | ( ng853  &  (~ ng27834)  &  wire35379 ) ;
 assign wire36198 = ( (~ ng826)  &  ng1114 ) | ( ng1114  &  (~ wire32243)  &  (~ wire32244) ) ;
 assign wire36201 = ( (~ ng1430)  &  (~ wire32701)  &  (~ wire32702) ) ;
 assign wire36202 = ( (~ ng1430)  &  (~ wire32701)  &  (~ wire32702) ) ;
 assign wire36203 = ( ng1430  &  wire32701 ) | ( ng1430  &  wire32702 ) ;
 assign wire36204 = ( ng1430  &  wire32701 ) | ( ng1430  &  wire32702 ) ;
 assign wire36205 = ( (~ ng1462)  &  (~ wire32691)  &  (~ wire32692) ) ;
 assign wire36206 = ( (~ ng1462)  &  (~ wire32691)  &  (~ wire32692) ) ;
 assign wire36207 = ( ng1462  &  wire32691 ) | ( ng1462  &  wire32692 ) ;
 assign wire36208 = ( ng1462  &  wire32691 ) | ( ng1462  &  wire32692 ) ;
 assign wire36209 = ( (~ ng1439)  &  (~ wire32681)  &  (~ wire32682) ) ;
 assign wire36210 = ( (~ ng1439)  &  (~ wire32681)  &  (~ wire32682) ) ;
 assign wire36211 = ( ng1439  &  wire32681 ) | ( ng1439  &  wire32682 ) ;
 assign wire36212 = ( ng1439  &  wire32681 ) | ( ng1439  &  wire32682 ) ;
 assign wire36213 = ( (~ ng1453)  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire36214 = ( (~ ng1453)  &  (~ wire32671)  &  (~ wire32672) ) ;
 assign wire36215 = ( ng1453  &  wire32671 ) | ( ng1453  &  wire32672 ) ;
 assign wire36216 = ( ng1453  &  wire32671 ) | ( ng1453  &  wire32672 ) ;
 assign wire36217 = ( (~ ng1457)  &  (~ wire32610)  &  (~ wire32611) ) ;
 assign wire36218 = ( ng1457  &  wire32610 ) | ( ng1457  &  wire32611 ) ;
 assign wire36219 = ( (~ ng1444)  &  (~ wire32661)  &  (~ wire32662) ) ;
 assign wire36220 = ( ng1444  &  wire32661 ) | ( ng1444  &  wire32662 ) ;
 assign wire36221 = ( (~ ng1435)  &  (~ wire32620)  &  (~ wire32621) ) ;
 assign wire36222 = ( ng1435  &  wire32620 ) | ( ng1435  &  wire32621 ) ;
 assign wire36223 = ( (~ ng1426)  &  (~ wire32590)  &  (~ wire32591) ) ;
 assign wire36224 = ( ng1426  &  wire32590 ) | ( ng1426  &  wire32591 ) ;
 assign wire36225 = ( (~ ng1466)  &  (~ wire32712)  &  (~ wire32713) ) ;
 assign wire36226 = ( ng1466  &  wire32712 ) | ( ng1466  &  wire32713 ) ;
 assign wire36227 = ( (~ ng1448)  &  (~ wire32600)  &  (~ wire32601) ) ;
 assign wire36228 = ( ng1448  &  wire32600 ) | ( ng1448  &  wire32601 ) ;
 assign wire36229 = ( (~ ng1457)  &  (~ wire32610)  &  (~ wire32611) ) ;
 assign wire36230 = ( ng1457  &  wire32610 ) | ( ng1457  &  wire32611 ) ;
 assign wire36231 = ( (~ ng1444)  &  (~ wire32661)  &  (~ wire32662) ) ;
 assign wire36232 = ( ng1444  &  wire32661 ) | ( ng1444  &  wire32662 ) ;
 assign wire36233 = ( (~ ng1435)  &  (~ wire32620)  &  (~ wire32621) ) ;
 assign wire36234 = ( ng1435  &  wire32620 ) | ( ng1435  &  wire32621 ) ;
 assign wire36235 = ( (~ ng1426)  &  (~ wire32590)  &  (~ wire32591) ) ;
 assign wire36236 = ( ng1426  &  wire32590 ) | ( ng1426  &  wire32591 ) ;
 assign wire36237 = ( (~ ng1466)  &  (~ wire32712)  &  (~ wire32713) ) ;
 assign wire36238 = ( ng1466  &  wire32712 ) | ( ng1466  &  wire32713 ) ;
 assign wire36239 = ( (~ ng1448)  &  (~ wire32600)  &  (~ wire32601) ) ;
 assign wire36240 = ( ng1448  &  wire32600 ) | ( ng1448  &  wire32601 ) ;
 assign wire36241 = ( (~ ng11675)  &  wire36201 ) | ( (~ ng11630)  &  wire36201 ) | ( (~ ng11666)  &  wire36201 ) | ( (~ ng11675)  &  ng11630  &  (~ ng11666) ) ;
 assign wire36242 = ( (~ ng11666)  &  wire36203 ) | ( (~ wire32703)  &  wire36203 ) | ( (~ ng11666)  &  wire36205 ) | ( (~ wire32703)  &  wire36205 ) ;
 assign wire36243 = ( (~ ng11666)  &  wire36207 ) | ( (~ wire32703)  &  wire36207 ) | ( (~ ng11666)  &  wire36209 ) | ( (~ wire32703)  &  wire36209 ) ;
 assign wire36244 = ( (~ ng11666)  &  wire36211 ) | ( (~ wire32703)  &  wire36211 ) | ( (~ ng11666)  &  wire36213 ) | ( (~ wire32703)  &  wire36213 ) ;
 assign wire36245 = ( (~ ng11666)  &  wire36215 ) | ( (~ wire32703)  &  wire36215 ) | ( (~ ng11666)  &  wire36217 ) | ( (~ wire32703)  &  wire36217 ) ;
 assign wire36246 = ( (~ ng11666)  &  wire36218 ) | ( (~ wire32703)  &  wire36218 ) | ( (~ ng11666)  &  wire36219 ) | ( (~ wire32703)  &  wire36219 ) ;
 assign wire36247 = ( (~ ng11666)  &  wire36220 ) | ( (~ wire32703)  &  wire36220 ) | ( (~ ng11666)  &  wire36221 ) | ( (~ wire32703)  &  wire36221 ) ;
 assign wire36248 = ( (~ ng11666)  &  wire36222 ) | ( (~ wire32703)  &  wire36222 ) | ( (~ ng11666)  &  wire36223 ) | ( (~ wire32703)  &  wire36223 ) ;
 assign wire36249 = ( (~ ng11666)  &  wire36224 ) | ( (~ wire32703)  &  wire36224 ) | ( (~ ng11666)  &  wire36225 ) | ( (~ wire32703)  &  wire36225 ) ;
 assign wire36250 = ( (~ ng11666)  &  wire36226 ) | ( (~ wire32703)  &  wire36226 ) | ( (~ ng11666)  &  wire36227 ) | ( (~ wire32703)  &  wire36227 ) ;
 assign wire36251 = ( (~ ng11666)  &  ng10711 ) | ( ng10711  &  (~ wire32703) ) | ( (~ ng11666)  &  wire36228 ) | ( (~ wire32703)  &  wire36228 ) ;
 assign wire36256 = ( wire36250 ) | ( wire36249 ) ;
 assign wire36257 = ( wire36251 ) | ( (~ wire32730)  &  wire36202 ) | ( (~ wire32731)  &  wire36202 ) ;
 assign wire36258 = ( (~ wire32730)  &  wire36204 ) | ( (~ wire32731)  &  wire36204 ) | ( (~ wire32730)  &  wire36206 ) | ( (~ wire32731)  &  wire36206 ) ;
 assign wire36259 = ( (~ wire32730)  &  wire36208 ) | ( (~ wire32731)  &  wire36208 ) | ( (~ wire32730)  &  wire36210 ) | ( (~ wire32731)  &  wire36210 ) ;
 assign wire36260 = ( (~ wire32730)  &  wire36212 ) | ( (~ wire32731)  &  wire36212 ) | ( (~ wire32730)  &  wire36214 ) | ( (~ wire32731)  &  wire36214 ) ;
 assign wire36261 = ( (~ wire32730)  &  wire36216 ) | ( (~ wire32731)  &  wire36216 ) | ( (~ wire32730)  &  wire36229 ) | ( (~ wire32731)  &  wire36229 ) ;
 assign wire36262 = ( (~ wire32730)  &  wire36230 ) | ( (~ wire32731)  &  wire36230 ) | ( (~ wire32730)  &  wire36231 ) | ( (~ wire32731)  &  wire36231 ) ;
 assign wire36263 = ( (~ wire32730)  &  wire36232 ) | ( (~ wire32731)  &  wire36232 ) | ( (~ wire32730)  &  wire36233 ) | ( (~ wire32731)  &  wire36233 ) ;
 assign wire36264 = ( (~ wire32730)  &  wire36234 ) | ( (~ wire32731)  &  wire36234 ) | ( (~ wire32730)  &  wire36235 ) | ( (~ wire32731)  &  wire36235 ) ;
 assign wire36265 = ( (~ wire32730)  &  wire36236 ) | ( (~ wire32731)  &  wire36236 ) | ( (~ wire32730)  &  wire36237 ) | ( (~ wire32731)  &  wire36237 ) ;
 assign wire36266 = ( (~ wire32730)  &  wire36238 ) | ( (~ wire32731)  &  wire36238 ) | ( (~ wire32730)  &  wire36239 ) | ( (~ wire32731)  &  wire36239 ) ;
 assign wire36267 = ( ng10711  &  (~ wire32730) ) | ( ng10711  &  (~ wire32731) ) | ( (~ wire32730)  &  wire36240 ) | ( (~ wire32731)  &  wire36240 ) ;
 assign wire36268 = ( wire36241 ) | ( wire36242 ) | ( wire36243 ) | ( wire36244 ) ;
 assign wire36269 = ( wire36245 ) | ( wire36246 ) | ( wire36247 ) | ( wire36248 ) ;
 assign wire36276 = ( wire36269 ) | ( wire36268 ) ;
 assign wire36277 = ( wire36256 ) | ( wire36257 ) | ( wire36258 ) | ( wire36259 ) ;
 assign wire36278 = ( wire36260 ) | ( wire36261 ) | ( wire36262 ) | ( wire36263 ) ;
 assign wire36279 = ( wire36264 ) | ( wire36265 ) | ( wire36266 ) | ( wire36267 ) ;
 assign wire36284 = ( wire3902 ) | ( ng27113  &  ng17162 ) ;
 assign wire36287 = ( wire3893 ) | ( wire3894 ) ;
 assign wire36288 = ( wire36287 ) | ( (~ ng1890)  &  ng1937  &  (~ ng29710) ) ;
 assign wire36289 = ( ng12124  &  wire3183 ) | ( wire3183  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36290 = ( wire3886 ) | ( ng30072  &  ng17194 ) | ( ng17194  &  wire35748 ) ;
 assign wire36297 = ( ng17973 ) | ( wire3281  &  (~ ng8381)  &  (~ wire34079) ) ;
 assign wire36302 = ( wire3858 ) | ( wire3857 ) ;
 assign wire36303 = ( wire3846 ) | ( wire3852 ) | ( wire36297 ) ;
 assign wire36304 = ( ng3098  &  (~ ng15841) ) | ( ng3147  &  wire3397 ) ;
 assign wire36305 = ( ng3102  &  (~ ng15757) ) | ( ng3101  &  (~ ng15719) ) ;
 assign wire36306 = ( wire3845 ) | ( wire3856 ) | ( ng3097  &  (~ ng15830) ) ;
 assign wire36307 = ( wire3850 ) | ( wire3851 ) | ( wire3854 ) | ( wire3855 ) ;
 assign wire36311 = ( wire36302 ) | ( wire36303 ) | ( wire36304 ) | ( wire36305 ) ;
 assign wire36312 = ( (~ ng17031)  &  ng65 ) ;
 assign wire36314 = ( (~ ng17031)  &  ng61 ) ;
 assign wire36321 = ( wire3727 ) | ( ng27113  &  ng17162 ) ;
 assign wire36323 = ( wire3277 ) | ( wire3721 ) ;
 assign wire36324 = ( ng12068  &  wire3189 ) | ( wire3189  &  (~ wire35745)  &  (~ wire35746) ) ;
 assign wire36325 = ( wire3715 ) | ( ng30072  &  ng17194 ) | ( ng17194  &  wire35748 ) ;
 assign wire36326 = ( ng1222  &  wire3143 ) | ( ng27113  &  wire3143 ) ;
 assign wire36327 = ( wire36326 ) | ( (~ ng1196)  &  ng1243  &  (~ ng27811) ) ;
 assign wire36330 = ( (~ pg3229)  &  (~ ng1890)  &  (~ ng1937)  &  ng1921 ) ;
 assign wire36331 = ( (~ ng1890)  &  (~ ng1937)  &  ng1905  &  wire36330 ) ;
 assign wire36334 = ( pg3229  &  (~ ng1890)  &  (~ ng1937)  &  ng1918 ) ;
 assign wire36335 = ( (~ ng1890)  &  (~ ng1937)  &  ng1905  &  wire36334 ) ;
 assign wire36342 = ( wire3673 ) | ( wire3672 ) ;
 assign wire36344 = ( wire36342 ) | ( ng1937  &  (~ ng29710)  &  ng29718 ) | ( ng1937  &  ng29710  &  (~ ng29718) ) ;
 assign wire36346 = ( ng1223  &  wire3143 ) | ( ng27113  &  wire3143 ) ;
 assign wire36347 = ( wire36346 ) | ( (~ ng1196)  &  ng1243  &  (~ ng27824) ) ;
 assign wire36348 = ( wire3660 ) | ( wire3661 ) ;
 assign wire36349 = ( wire36348 ) | ( (~ ng1890)  &  ng1937  &  (~ ng29718) ) ;
 assign wire36352 = ( pg3229  &  (~ ng2631)  &  (~ ng2584)  &  ng2612 ) ;
 assign wire36353 = ( (~ ng2631)  &  (~ ng2584)  &  ng2599  &  wire36352 ) ;
 assign wire36356 = ( (~ pg3229)  &  (~ ng2631)  &  (~ ng2584)  &  ng2615 ) ;
 assign wire36357 = ( (~ ng2631)  &  (~ ng2584)  &  ng2599  &  wire36356 ) ;
 assign wire36362 = ( (~ ng30072)  &  (~ wire35748)  &  wire36353 ) | ( (~ ng30072)  &  (~ wire35748)  &  wire36357 ) ;
 assign wire36364 = ( wire36362 ) | ( ng2631  &  (~ ng30594)  &  ng30602 ) | ( ng2631  &  ng30594  &  (~ ng30602) ) ;
 assign wire36369 = ( ng3036  &  (~ ng3032) ) ;
 assign wire36370 = ( ng21796  &  (~ wire36177)  &  wire36369 ) | ( wire36176  &  (~ wire36177)  &  wire36369 ) ;
 assign wire36377 = ( (~ pg8021)  &  (~ ng2912) ) | ( (~ pg8021)  &  ng2917 ) ;
 assign wire36378 = ( wire3564 ) | ( (~ pg8021)  &  (~ ng2912) ) | ( (~ pg8021)  &  ng2917 ) ;
 assign wire36379 = ( ng2912  &  (~ wire35029) ) | ( ng2912  &  (~ wire35030) ) | ( (~ ng2912)  &  wire35029  &  wire35030 ) ;
 assign wire36380 = ( ng2917  &  (~ wire35029) ) | ( ng2917  &  (~ wire35030) ) ;
 assign wire36381 = ( ng2917  &  (~ ng2912) ) ;
 assign wire36382 = ( (~ ng2917)  &  wire35029  &  wire35030 ) ;
 assign wire36383 = ( (~ wire3139)  &  wire36380 ) | ( wire36378  &  wire36380 ) | ( (~ wire3139)  &  wire36381 ) | ( wire36378  &  wire36381 ) ;
 assign wire36385 = ( ng2917  &  (~ ng2924)  &  wire35029  &  wire35030 ) ;
 assign wire36386 = ( ng2924  &  (~ ng2917) ) ;
 assign wire36387 = ( wire3527 ) | ( (~ wire3139)  &  wire36386 ) | ( wire36378  &  wire36386 ) ;
 assign wire36388 = ( (~ ng826)  &  ng2502 ) | ( ng2502  &  (~ wire33906)  &  (~ wire33907) ) ;
 assign wire36389 = ( (~ ng2920)  &  ng2924 ) ;
 assign wire36390 = ( (~ wire3139)  &  (~ wire36379)  &  wire36389 ) | ( wire36378  &  (~ wire36379)  &  wire36389 ) ;
 assign wire36391 = ( wire3512 ) | ( (~ wire3529)  &  (~ wire36387)  &  wire36390 ) ;
 assign wire36412 = ( ng2020  &  ng11914  &  wire35607 ) | ( (~ ng2020)  &  (~ ng11914)  &  wire35607 ) | ( ng2020  &  ng11914  &  wire35608 ) | ( (~ ng2020)  &  (~ ng11914)  &  wire35608 ) ;
 assign wire36413 = ( ng2052  &  ng12171  &  wire35607 ) | ( (~ ng2052)  &  (~ ng12171)  &  wire35607 ) | ( ng2052  &  ng12171  &  wire35608 ) | ( (~ ng2052)  &  (~ ng12171)  &  wire35608 ) ;
 assign wire36414 = ( ng2059  &  ng12263  &  wire35607 ) | ( (~ ng2059)  &  (~ ng12263)  &  wire35607 ) | ( ng2059  &  ng12263  &  wire35608 ) | ( (~ ng2059)  &  (~ ng12263)  &  wire35608 ) ;
 assign wire36415 = ( ng2013  &  ng12172  &  wire35577 ) | ( ng2013  &  ng12172  &  wire35578 ) | ( (~ ng2013)  &  ng12172  &  (~ wire35577)  &  (~ wire35578) ) ;
 assign wire36416 = ( ng2033  &  ng11999  &  wire35607 ) | ( (~ ng2033)  &  (~ ng11999)  &  wire35607 ) | ( ng2033  &  ng11999  &  wire35608 ) | ( (~ ng2033)  &  (~ ng11999)  &  wire35608 ) ;
 assign wire36417 = ( ng2066  &  ng12293  &  wire35607 ) | ( (~ ng2066)  &  (~ ng12293)  &  wire35607 ) | ( ng2066  &  ng12293  &  wire35608 ) | ( (~ ng2066)  &  (~ ng12293)  &  wire35608 ) ;
 assign wire36418 = ( ng2072  &  ng12172  &  wire35587 ) | ( ng2072  &  ng12172  &  wire35588 ) | ( (~ ng2072)  &  ng12172  &  (~ wire35587)  &  (~ wire35588) ) ;
 assign wire36419 = ( ng2026  &  ng12060  &  wire35607 ) | ( (~ ng2026)  &  (~ ng12060)  &  wire35607 ) | ( ng2026  &  ng12060  &  wire35608 ) | ( (~ ng2026)  &  (~ ng12060)  &  wire35608 ) ;
 assign wire36420 = ( ng2040  &  ng12112  &  wire35607 ) | ( (~ ng2040)  &  (~ ng12112)  &  wire35607 ) | ( ng2040  &  ng12112  &  wire35608 ) | ( (~ ng2040)  &  (~ ng12112)  &  wire35608 ) ;
 assign wire36426 = ( wire36420 ) | ( ng2046  &  ng12216  &  ng12172 ) | ( (~ ng2046)  &  (~ ng12216)  &  ng12172 ) ;
 assign wire36427 = ( wire36412 ) | ( wire36413 ) | ( wire36414 ) | ( wire36415 ) ;
 assign wire36428 = ( wire36416 ) | ( wire36417 ) | ( wire36418 ) | ( wire36419 ) ;
 assign wire36431 = ( ng2108  &  ng2109  &  ng2110 ) ;
 assign wire36433 = ( (~ ng1315)  &  ng2109  &  ng2110 ) ;
 assign wire36435 = ( (~ ng1309)  &  ng2108  &  ng2110 ) ;
 assign wire36437 = ( (~ ng1312)  &  ng2108  &  ng2109 ) ;
 assign wire36438 = ( (~ ng1312)  &  (~ ng1315)  &  ng2109 ) ;
 assign wire36439 = ( (~ ng1312)  &  (~ ng1309)  &  ng2108 ) ;
 assign wire36440 = ( (~ ng1315)  &  (~ ng1309)  &  ng2110 ) ;
 assign wire36445 = ( wire3422 ) | ( wire3423 ) | ( wire3424 ) | ( wire3441 ) ;
 assign wire36446 = ( wire3448 ) | ( wire3449 ) | ( wire3450 ) | ( wire3451 ) ;
 assign wire36455 = ( wire3049 ) | ( wire3388 ) | ( wire3390 ) | ( wire3391 ) ;
 assign wire36456 = ( wire3392 ) | ( wire3393 ) | ( wire3394 ) | ( wire3396 ) ;
 assign wire36457 = ( wire3213 ) | ( (~ ng853)  &  ng1702 ) ;
 assign wire36458 = ( wire36457 ) | ( (~ ng13165)  &  ng17124  &  (~ ng27875) ) ;
 assign wire36459 = ( ng13055  &  (~ wire33296)  &  (~ wire33297)  &  (~ wire33298) ) ;
 assign wire36461 = ( ng13055  &  wire33296 ) | ( ng13055  &  wire33297 ) | ( ng13055  &  wire33298 ) ;
 assign wire36462 = ( (~ wire33376)  &  (~ wire33377)  &  wire36461 ) ;
 assign wire36463 = ( wire3167 ) | ( (~ ng13055)  &  (~ wire33147)  &  (~ wire33148) ) ;
 assign wire36465 = ( ng2040  &  ng2052  &  ng2046 ) ;
 assign wire36474 = ( (~ ng1312)  &  ng2052 ) | ( ng2052  &  (~ ng2010) ) ;
 assign wire36476 = ( (~ ng1312)  &  ng2046 ) | ( (~ ng2010)  &  ng2046 ) ;


endmodule

