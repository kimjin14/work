module seq (
	i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, 
	i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, 
	i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, 
	i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, 
	i_38_, i_29_, i_37_, o_1_, o_19_, o_2_, o_0_, o_29_, o_25_, o_12_, 
	o_26_, o_11_, o_27_, o_14_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, 
	o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, 
	o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

input i_40_;
input i_30_;
input i_20_;
input i_9_;
input i_10_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_27_;
input i_14_;
input i_3_;
input i_39_;
input i_28_;
input i_13_;
input i_4_;
input i_25_;
input i_12_;
input i_1_;
input i_26_;
input i_11_;
input i_2_;
input i_23_;
input i_18_;
input i_24_;
input i_17_;
input i_0_;
input i_21_;
input i_16_;
input i_22_;
input i_15_;
input i_32_;
input i_31_;
input i_34_;
input i_33_;
input i_19_;
input i_36_;
input i_35_;
input i_38_;
input i_29_;
input i_37_;
output o_1_;
output o_19_;
output o_2_;
output o_0_;
output o_29_;
output o_25_;
output o_12_;
output o_26_;
output o_11_;
output o_27_;
output o_14_;
output o_28_;
output o_13_;
output o_34_;
output o_21_;
output o_16_;
output o_33_;
output o_22_;
output o_15_;
output o_32_;
output o_23_;
output o_18_;
output o_31_;
output o_24_;
output o_17_;
output o_30_;
output o_20_;
output o_10_;
output o_9_;
output o_7_;
output o_8_;
output o_5_;
output o_6_;
output o_3_;
output o_4_;
wire n_n955;
wire n_n709;
wire wire66;
wire wire145;
wire wire363;
wire wire537;
wire wire543;
wire n_n1055;
wire n_n985;
wire n_n979;
wire n_n515;
wire n_n1008;
wire n_n842;
wire n_n1067;
wire n_n982;
wire n_n990;
wire wire88;
wire wire330;
wire n_n1373;
wire n_n1164;
wire n_n1165;
wire wire48;
wire wire241;
wire wire432;
wire wire491;
wire wire549;
wire n_n1083;
wire n_n978;
wire n_n883;
wire n_n998;
wire n_n1021;
wire n_n330;
wire n_n969;
wire n_n2487;
wire n_n973;
wire n_n158;
wire n_n2488;
wire n_n1084;
wire n_n1777;
wire wire35;
wire n_n469;
wire n_n1993;
wire wire553;
wire n_n2581;
wire n_n1971;
wire n_n1581;
wire n_n1603;
wire wire173;
wire wire223;
wire n_n685;
wire n_n2838;
wire n_n2836;
wire n_n1990;
wire n_n1951;
wire wire555;
wire n_n926;
wire n_n2213;
wire n_n1394;
wire wire92;
wire wire319;
wire wire422;
wire wire470;
wire wire556;
wire n_n761;
wire n_n760;
wire n_n1628;
wire n_n1630;
wire n_n1631;
wire wire175;
wire wire240;
wire wire323;
wire wire559;
wire wire225;
wire n_n1011;
wire n_n980;
wire n_n1006;
wire n_n989;
wire n_n983;
wire n_n1709;
wire n_n1711;
wire wire445;
wire wire560;
wire n_n865;
wire n_n1525;
wire wire47;
wire n_n971;
wire n_n1005;
wire n_n997;
wire n_n975;
wire n_n880;
wire wire390;
wire wire411;
wire wire436;
wire wire526;
wire wire566;
wire wire565;
wire n_n1014;
wire n_n1528;
wire n_n1530;
wire wire183;
wire wire251;
wire wire335;
wire wire354;
wire wire392;
wire n_n874;
wire n_n966;
wire n_n862;
wire n_n1549;
wire n_n1552;
wire wire490;
wire n_n1445;
wire wire346;
wire n_n1986;
wire n_n837;
wire wire245;
wire wire364;
wire wire371;
wire wire570;
wire n_n1571;
wire n_n1408;
wire n_n1409;
wire n_n1411;
wire n_n968;
wire n_n819;
wire n_n1651;
wire wire99;
wire wire365;
wire wire572;
wire wire571;
wire n_n1489;
wire wire182;
wire wire301;
wire wire574;
wire wire575;
wire n_n857;
wire n_n411;
wire n_n1372;
wire wire57;
wire wire84;
wire wire416;
wire wire512;
wire wire579;
wire n_n1072;
wire n_n937;
wire n_n1374;
wire wire120;
wire wire333;
wire wire386;
wire wire583;
wire wire581;
wire wire146;
wire n_n698;
wire wire131;
wire wire402;
wire wire493;
wire wire495;
wire n_n1330;
wire n_n1332;
wire n_n866;
wire n_n1323;
wire wire316;
wire wire587;
wire wire586;
wire n_n1187;
wire n_n1184;
wire wire45;
wire wire202;
wire wire406;
wire n_n1233;
wire n_n775;
wire n_n785;
wire n_n1242;
wire wire469;
wire n_n528;
wire n_n977;
wire n_n888;
wire n_n313;
wire wire227;
wire wire508;
wire wire594;
wire n_n1326;
wire wire68;
wire wire174;
wire wire300;
wire wire504;
wire n_n1283;
wire n_n833;
wire wire176;
wire wire395;
wire wire598;
wire wire596;
wire wire595;
wire n_n1280;
wire n_n1052;
wire n_n1064;
wire n_n525;
wire wire148;
wire wire329;
wire wire357;
wire wire408;
wire wire441;
wire wire542;
wire n_n764;
wire wire600;
wire n_n1272;
wire n_n799;
wire n_n1237;
wire n_n1239;
wire wire398;
wire wire602;
wire n_n1235;
wire n_n861;
wire n_n793;
wire wire420;
wire wire604;
wire wire407;
wire n_n1048;
wire wire349;
wire wire607;
wire n_n1094;
wire n_n2837;
wire n_n1958;
wire n_n1956;
wire n_n1957;
wire n_n964;
wire n_n1073;
wire n_n1009;
wire n_n1002;
wire n_n960;
wire n_n1001;
wire n_n993;
wire wire81;
wire wire46;
wire wire382;
wire n_n933;
wire n_n1066;
wire n_n967;
wire wire86;
wire n_n1074;
wire n_n642;
wire n_n1047;
wire n_n976;
wire n_n1015;
wire n_n795;
wire n_n848;
wire n_n945;
wire n_n853;
wire n_n559;
wire wire87;
wire wire320;
wire n_n535;
wire wire471;
wire n_n949;
wire n_n460;
wire n_n1061;
wire n_n1023;
wire wire359;
wire n_n952;
wire wire317;
wire wire78;
wire n_n947;
wire n_n935;
wire n_n329;
wire n_n527;
wire n_n710;
wire wire400;
wire n_n688;
wire n_n462;
wire n_n700;
wire n_n492;
wire wire100;
wire n_n1065;
wire n_n488;
wire n_n453;
wire wire77;
wire n_n1012;
wire wire334;
wire wire378;
wire n_n884;
wire wire326;
wire n_n970;
wire n_n928;
wire n_n951;
wire n_n860;
wire n_n560;
wire n_n484;
wire wire60;
wire wire76;
wire wire103;
wire wire531;
wire wire611;
wire n_n1416;
wire wire430;
wire wire612;
wire wire462;
wire n_n1203;
wire n_n1202;
wire n_n777;
wire n_n781;
wire wire37;
wire wire64;
wire wire94;
wire wire106;
wire wire321;
wire wire614;
wire n_n1057;
wire n_n1056;
wire wire61;
wire n_n629;
wire wire410;
wire wire50;
wire wire315;
wire n_n162;
wire n_n991;
wire n_n334;
wire n_n801;
wire n_n428;
wire n_n427;
wire n_n843;
wire n_n791;
wire n_n459;
wire n_n905;
wire n_n1414;
wire n_n1412;
wire wire467;
wire wire616;
wire wire615;
wire n_n475;
wire n_n164;
wire n_n1417;
wire wire113;
wire wire617;
wire wire506;
wire wire619;
wire wire433;
wire wire621;
wire n_n2439;
wire wire624;
wire wire623;
wire wire352;
wire wire421;
wire wire518;
wire wire524;
wire wire627;
wire n_n1197;
wire wire36;
wire n_n1193;
wire wire633;
wire n_n1195;
wire wire154;
wire wire635;
wire wire65;
wire wire637;
wire n_n1135;
wire n_n1053;
wire n_n582;
wire n_n850;
wire wire367;
wire n_n771;
wire wire368;
wire wire479;
wire wire369;
wire wire393;
wire wire468;
wire wire83;
wire wire356;
wire wire643;
wire n_n1285;
wire wire486;
wire wire648;
wire wire646;
wire n_n923;
wire n_n1196;
wire n_n1068;
wire wire303;
wire wire520;
wire wire655;
wire n_n864;
wire wire79;
wire wire238;
wire wire336;
wire n_n458;
wire n_n643;
wire n_n1611;
wire n_n836;
wire wire394;
wire wire660;
wire wire366;
wire wire662;
wire wire54;
wire wire80;
wire wire325;
wire wire463;
wire wire135;
wire wire666;
wire wire665;
wire wire664;
wire wire153;
wire wire184;
wire wire187;
wire wire667;
wire wire458;
wire wire669;
wire wire668;
wire wire73;
wire wire327;
wire wire670;
wire wire671;
wire wire672;
wire wire529;
wire wire370;
wire n_n918;
wire n_n556;
wire n_n798;
wire wire110;
wire n_n859;
wire wire351;
wire wire674;
wire wire403;
wire wire676;
wire wire675;
wire wire69;
wire wire332;
wire wire680;
wire wire679;
wire wire678;
wire wire413;
wire wire684;
wire wire484;
wire n_n1091;
wire n_n1113;
wire wire244;
wire wire688;
wire n_n1081;
wire n_n1088;
wire n_n1086;
wire n_n1108;
wire wire464;
wire wire689;
wire wire132;
wire wire690;
wire n_n927;
wire wire82;
wire n_n773;
wire n_n715;
wire wire337;
wire wire344;
wire wire692;
wire wire696;
wire wire695;
wire wire102;
wire wire697;
wire wire509;
wire wire396;
wire wire342;
wire wire380;
wire wire702;
wire wire701;
wire wire700;
wire n_n783;
wire wire376;
wire n_n668;
wire n_n550;
wire wire401;
wire wire704;
wire wire706;
wire wire710;
wire wire149;
wire wire155;
wire wire383;
wire wire429;
wire wire711;
wire n_n1577;
wire wire713;
wire n_n1488;
wire wire718;
wire wire717;
wire wire139;
wire n_n1453;
wire wire488;
wire wire723;
wire n_n1452;
wire wire724;
wire wire727;
wire wire473;
wire n_n1277;
wire n_n693;
wire wire361;
wire wire737;
wire wire739;
wire wire740;
wire n_n1134;
wire wire742;
wire wire741;
wire n_n673;
wire wire124;
wire wire744;
wire wire535;
wire wire748;
wire n_n790;
wire wire166;
wire wire752;
wire wire140;
wire wire156;
wire wire494;
wire wire758;
wire n_n765;
wire n_n907;
wire wire761;
wire wire763;
wire wire762;
wire wire766;
wire wire348;
wire n_n1607;
wire wire101;
wire wire127;
wire wire772;
wire wire373;
wire n_n1575;
wire wire775;
wire wire461;
wire wire777;
wire n_n1672;
wire n_n1572;
wire wire780;
wire wire779;
wire wire476;
wire wire782;
wire wire786;
wire wire787;
wire n_n1580;
wire wire59;
wire wire788;
wire wire795;
wire wire794;
wire n_n1716;
wire wire158;
wire n_n1670;
wire wire185;
wire wire803;
wire wire806;
wire wire805;
wire wire808;
wire wire807;
wire wire811;
wire wire810;
wire wire809;
wire wire814;
wire wire450;
wire wire817;
wire wire465;
wire wire475;
wire wire822;
wire wire825;
wire wire826;
wire wire38;
wire wire39;
wire wire42;
wire wire43;
wire wire44;
wire wire53;
wire wire55;
wire wire304;
wire wire63;
wire wire67;
wire wire318;
wire wire492;
wire wire70;
wire wire104;
wire wire115;
wire wire302;
wire wire121;
wire wire830;
wire wire829;
wire wire831;
wire wire233;
wire wire835;
wire wire837;
wire wire375;
wire wire482;
wire wire474;
wire wire478;
wire wire481;
wire wire840;
wire wire483;
wire wire496;
wire wire546;
wire wire548;
wire wire558;
wire wire589;
wire wire609;
wire wire613;
wire wire622;
wire wire636;
wire wire638;
wire wire642;
wire wire652;
wire wire650;
wire wire677;
wire wire681;
wire wire686;
wire wire687;
wire wire693;
wire wire715;
wire wire716;
wire wire721;
wire wire729;
wire wire732;
wire wire731;
wire wire738;
wire wire743;
wire wire749;
wire wire756;
wire wire765;
wire wire767;
wire wire781;
wire wire785;
wire wire793;
wire wire792;
wire wire797;
wire wire801;
wire wire813;
wire wire818;
wire wire820;
wire wire824;
wire wire828;
wire wire841;
wire wire56;
wire wire74;
wire wire129;
wire wire133;
wire wire136;
wire wire137;
wire wire138;
wire wire141;
wire wire142;
wire wire143;
wire wire144;
wire wire151;
wire wire160;
wire wire162;
wire wire163;
wire wire164;
wire wire165;
wire wire167;
wire wire169;
wire wire170;
wire wire171;
wire wire188;
wire wire189;
wire wire190;
wire wire191;
wire wire192;
wire wire193;
wire wire196;
wire wire197;
wire wire198;
wire wire199;
wire wire201;
wire wire203;
wire wire205;
wire wire206;
wire wire207;
wire wire208;
wire wire209;
wire wire210;
wire wire211;
wire wire213;
wire wire217;
wire wire218;
wire wire226;
wire wire229;
wire wire231;
wire wire232;
wire wire234;
wire wire235;
wire wire243;
wire wire248;
wire wire249;
wire wire250;
wire wire252;
wire wire254;
wire wire260;
wire wire261;
wire wire262;
wire wire263;
wire wire264;
wire wire271;
wire wire272;
wire wire274;
wire wire276;
wire wire277;
wire wire279;
wire wire283;
wire wire284;
wire wire285;
wire wire286;
wire wire287;
wire wire288;
wire wire289;
wire wire291;
wire wire294;
wire wire295;
wire wire297;
wire wire298;
wire wire299;
wire wire306;
wire wire307;
wire wire308;
wire wire309;
wire wire310;
wire wire311;
wire wire312;
wire wire414;
wire wire443;
wire wire444;
wire wire446;
wire wire447;
wire wire449;
wire wire451;
wire wire454;
wire wire455;
wire wire459;
wire wire519;
wire wire533;
wire wire536;
wire wire538;
wire wire843;
wire wire845;
wire wire846;
wire wire847;
wire wire849;
wire wire850;
wire wire855;
wire wire856;
wire wire857;
wire wire859;
wire wire860;
wire wire864;
wire wire865;
wire wire869;
wire wire872;
wire wire873;
wire wire875;
wire wire876;
wire wire882;
wire wire888;
wire wire890;
wire wire891;
wire wire892;
wire wire893;
wire wire894;
wire wire902;
wire wire904;
wire wire905;
wire wire906;
wire wire911;
wire wire912;
wire wire913;
wire wire920;
wire wire921;
wire wire922;
wire wire925;
wire wire926;
wire wire927;
wire wire928;
wire wire929;
wire wire930;
wire wire932;
wire wire934;
wire wire937;
wire wire939;
wire wire940;
wire wire942;
wire wire948;
wire wire950;
wire wire952;
wire wire957;
wire wire962;
wire wire964;
wire wire967;
wire wire973;
wire wire983;
wire wire985;
wire wire986;
wire wire987;
wire wire988;
wire wire999;
wire wire1000;
wire wire1008;
wire wire1010;
wire wire1019;
wire wire1020;
wire wire1021;
wire wire1022;
wire wire1029;
wire wire1031;
wire wire1038;
wire wire1039;
wire wire1040;
wire wire1043;
wire wire1044;
wire wire1046;
wire wire1048;
wire wire1049;
wire wire1050;
wire wire1051;
wire wire1058;
wire wire1059;
wire wire1060;
wire wire1061;
wire wire1062;
wire wire1063;
wire wire1065;
wire wire1067;
wire wire1073;
wire wire1075;
wire wire1078;
wire wire1083;
wire wire1084;
wire wire1085;
wire wire1088;
wire wire1089;
wire wire1090;
wire wire1091;
wire wire1092;
wire wire1093;
wire wire1099;
wire wire1104;
wire wire1106;
wire wire1107;
wire wire1109;
wire wire1112;
wire wire1113;
wire wire1114;
wire wire1119;
wire wire1120;
wire wire1122;
wire wire1132;
wire wire1139;
wire wire1155;
wire wire1156;
wire wire1158;
wire wire1160;
wire wire1163;
wire wire1164;
wire wire1165;
wire wire1168;
wire wire1169;
wire wire1173;
wire wire1174;
wire wire1179;
wire wire1181;
wire wire1182;
wire wire1183;
wire wire1186;
wire wire1189;
wire wire1192;
wire wire1196;
wire wire1197;
wire wire1198;
wire wire1199;
wire wire1200;
wire wire1204;
wire wire1205;
wire wire1206;
wire wire1208;
wire wire1210;
wire wire1213;
wire wire1219;
wire wire1222;
wire wire1230;
wire wire1238;
wire wire1246;
wire wire1247;
wire wire1251;
wire wire1252;
wire wire1253;
wire wire1254;
wire wire1255;
wire wire1256;
wire wire1257;
wire wire1262;
wire wire1264;
wire wire1265;
wire wire1269;
wire wire1271;
wire wire1277;
wire wire1284;
wire wire1285;
wire wire1286;
wire wire1289;
wire wire1291;
wire wire1294;
wire wire1295;
wire wire1299;
wire wire1300;
wire wire1305;
wire wire1306;
wire wire1307;
wire wire1309;
wire wire1311;
wire wire1312;
wire wire1316;
wire wire1317;
wire wire1326;
wire wire1328;
wire wire1329;
wire wire1330;
wire wire1340;
wire wire1341;
wire wire1342;
wire wire1343;
wire wire1344;
wire wire1346;
wire wire1347;
wire wire1348;
wire wire1349;
wire wire1353;
wire wire1354;
wire wire1356;
wire wire1357;
wire wire1358;
wire wire1362;
wire wire1364;
wire wire1365;
wire wire1366;
wire wire1367;
wire wire1371;
wire wire1372;
wire wire1374;
wire wire1375;
wire wire1381;
wire wire1383;
wire wire1386;
wire wire1388;
wire wire1389;
wire wire1390;
wire wire1400;
wire wire1402;
wire wire1412;
wire wire1415;
wire wire1416;
wire wire1417;
wire wire1423;
wire wire1428;
wire wire1429;
wire wire1430;
wire wire1435;
wire wire1438;
wire wire1441;
wire wire1442;
wire wire1443;
wire wire1444;
wire wire1447;
wire wire1448;
wire wire1449;
wire wire1450;
wire wire1451;
wire wire1452;
wire wire1453;
wire wire1454;
wire wire1455;
wire wire1459;
wire wire1466;
wire wire1467;
wire wire1468;
wire wire1472;
wire wire1475;
wire wire1483;
wire wire1484;
wire wire1487;
wire wire1489;
wire wire1496;
wire wire1499;
wire wire1501;
wire wire1505;
wire wire1506;
wire wire1509;
wire wire1510;
wire wire1518;
wire wire1520;
wire wire1521;
wire wire1522;
wire wire1524;
wire wire1525;
wire wire1539;
wire wire1540;
wire wire1541;
wire wire1542;
wire wire1544;
wire wire1545;
wire wire1546;
wire wire1547;
wire wire1548;
wire wire1550;
wire wire1551;
wire wire1552;
wire wire1555;
wire wire1557;
wire wire1562;
wire wire1563;
wire wire1565;
wire wire1566;
wire wire1568;
wire wire1570;
wire wire1571;
wire wire1575;
wire wire1577;
wire wire1578;
wire wire1579;
wire wire1583;
wire wire1584;
wire wire1588;
wire wire1592;
wire wire1610;
wire wire1617;
wire wire1619;
wire wire1620;
wire wire1624;
wire wire1626;
wire wire1630;
wire wire1632;
wire wire1635;
wire wire1650;
wire wire1651;
wire wire1653;
wire wire1655;
wire wire1657;
wire wire1661;
wire wire1662;
wire wire1666;
wire wire1681;
wire wire1682;
wire wire1693;
wire wire1700;
wire wire1701;
wire wire1704;
wire wire1705;
wire wire1706;
wire wire1707;
wire wire1708;
wire wire1709;
wire wire1715;
wire wire1730;
wire wire1731;
wire wire1741;
wire wire1742;
wire wire1747;
wire wire1749;
wire wire1751;
wire wire1758;
wire wire1766;
wire wire1780;
wire wire1786;
wire wire1789;
wire wire1791;
wire wire1792;
wire wire1793;
wire wire1795;
wire wire1797;
wire wire1798;
wire wire1803;
wire wire1804;
wire wire1805;
wire wire1806;
wire wire1807;
wire wire1810;
wire wire1812;
wire wire1821;
wire wire1822;
wire wire1823;
wire wire1832;
wire wire1834;
wire wire1835;
wire wire1836;
wire wire1838;
wire wire1839;
wire wire1842;
wire wire1844;
wire wire1845;
wire wire1846;
wire wire1847;
wire wire1850;
wire wire1852;
wire wire1853;
wire wire1854;
wire wire1855;
wire wire1860;
wire wire1861;
wire wire1862;
wire wire1863;
wire wire1867;
wire wire1868;
wire wire1870;
wire wire1871;
wire wire1872;
wire wire1875;
wire wire1878;
wire wire1880;
wire wire1881;
wire wire1882;
wire wire1883;
wire wire1884;
wire wire1890;
wire wire1891;
wire wire1896;
wire wire1901;
wire wire1902;
wire wire1905;
wire wire1909;
wire wire1910;
wire wire1911;
wire wire1912;
wire wire1913;
wire wire1914;
wire wire1915;
wire wire1916;
wire wire1919;
wire wire1920;
wire wire1923;
wire wire1926;
wire wire1933;
wire wire1934;
wire wire1935;
wire wire1936;
wire wire6716;
wire wire6719;
wire wire6722;
wire wire6723;
wire wire6724;
wire wire6726;
wire wire6727;
wire wire6728;
wire wire6729;
wire wire6731;
wire wire6734;
wire wire6736;
wire wire6739;
wire wire6740;
wire wire6741;
wire wire6746;
wire wire6747;
wire wire6749;
wire wire6750;
wire wire6751;
wire wire6753;
wire wire6754;
wire wire6757;
wire wire6758;
wire wire6759;
wire wire6764;
wire wire6765;
wire wire6766;
wire wire6767;
wire wire6770;
wire wire6772;
wire wire6773;
wire wire6774;
wire wire6778;
wire wire6779;
wire wire6780;
wire wire6786;
wire wire6788;
wire wire6789;
wire wire6790;
wire wire6791;
wire wire6793;
wire wire6794;
wire wire6798;
wire wire6800;
wire wire6801;
wire wire6804;
wire wire6806;
wire wire6807;
wire wire6808;
wire wire6813;
wire wire6818;
wire wire6821;
wire wire6824;
wire wire6828;
wire wire6831;
wire wire6832;
wire wire6837;
wire wire6839;
wire wire6841;
wire wire6842;
wire wire6844;
wire wire6845;
wire wire6849;
wire wire6850;
wire wire6851;
wire wire6853;
wire wire6854;
wire wire6856;
wire wire6857;
wire wire6858;
wire wire6859;
wire wire6860;
wire wire6861;
wire wire6863;
wire wire6865;
wire wire6866;
wire wire6868;
wire wire6869;
wire wire6870;
wire wire6873;
wire wire6874;
wire wire6877;
wire wire6878;
wire wire6879;
wire wire6884;
wire wire6886;
wire wire6887;
wire wire6888;
wire wire6889;
wire wire6890;
wire wire6894;
wire wire6897;
wire wire6901;
wire wire6902;
wire wire6904;
wire wire6907;
wire wire6908;
wire wire6909;
wire wire6910;
wire wire6911;
wire wire6913;
wire wire6914;
wire wire6915;
wire wire6920;
wire wire6924;
wire wire6925;
wire wire6927;
wire wire6929;
wire wire6930;
wire wire6932;
wire wire6933;
wire wire6934;
wire wire6935;
wire wire6938;
wire wire6940;
wire wire6941;
wire wire6942;
wire wire6945;
wire wire6948;
wire wire6949;
wire wire6950;
wire wire6951;
wire wire6952;
wire wire6955;
wire wire6956;
wire wire6957;
wire wire6958;
wire wire6960;
wire wire6961;
wire wire6964;
wire wire6965;
wire wire6968;
wire wire6969;
wire wire6970;
wire wire6971;
wire wire6974;
wire wire6975;
wire wire6976;
wire wire6978;
wire wire6979;
wire wire6980;
wire wire6981;
wire wire6982;
wire wire6984;
wire wire6985;
wire wire6987;
wire wire6991;
wire wire6993;
wire wire6994;
wire wire6998;
wire wire6999;
wire wire7000;
wire wire7001;
wire wire7002;
wire wire7005;
wire wire7007;
wire wire7008;
wire wire7011;
wire wire7012;
wire wire7014;
wire wire7016;
wire wire7018;
wire wire7020;
wire wire7021;
wire wire7025;
wire wire7026;
wire wire7029;
wire wire7030;
wire wire7033;
wire wire7034;
wire wire7035;
wire wire7038;
wire wire7040;
wire wire7043;
wire wire7044;
wire wire7048;
wire wire7050;
wire wire7051;
wire wire7052;
wire wire7053;
wire wire7055;
wire wire7057;
wire wire7058;
wire wire7062;
wire wire7063;
wire wire7064;
wire wire7066;
wire wire7067;
wire wire7069;
wire wire7071;
wire wire7073;
wire wire7074;
wire wire7077;
wire wire7079;
wire wire7086;
wire wire7087;
wire wire7089;
wire wire7090;
wire wire7092;
wire wire7094;
wire wire7095;
wire wire7097;
wire wire7100;
wire wire7102;
wire wire7103;
wire wire7104;
wire wire7105;
wire wire7108;
wire wire7109;
wire wire7110;
wire wire7115;
wire wire7118;
wire wire7119;
wire wire7121;
wire wire7122;
wire wire7123;
wire wire7124;
wire wire7125;
wire wire7127;
wire wire7128;
wire wire7129;
wire wire7130;
wire wire7131;
wire wire7132;
wire wire7133;
wire wire7135;
wire wire7137;
wire wire7139;
wire wire7140;
wire wire7142;
wire wire7143;
wire wire7145;
wire wire7146;
wire wire7148;
wire wire7150;
wire wire7151;
wire wire7152;
wire wire7153;
wire wire7154;
wire wire7157;
wire wire7160;
wire wire7161;
wire wire7164;
wire wire7165;
wire wire7170;
wire wire7171;
wire wire7175;
wire wire7176;
wire wire7178;
wire wire7180;
wire wire7181;
wire wire7182;
wire wire7184;
wire wire7185;
wire wire7187;
wire wire7189;
wire wire7190;
wire wire7191;
wire wire7193;
wire wire7194;
wire wire7195;
wire wire7197;
wire wire7200;
wire wire7201;
wire wire7204;
wire wire7205;
wire wire7208;
wire wire7210;
wire wire7211;
wire wire7214;
wire wire7218;
wire wire7219;
wire wire7220;
wire wire7223;
wire wire7227;
wire wire7230;
wire wire7231;
wire wire7233;
wire wire7234;
wire wire7237;
wire wire7239;
wire wire7245;
wire wire7246;
wire wire7252;
wire wire7253;
wire wire7256;
wire wire7257;
wire wire7258;
wire wire7260;
wire wire7261;
wire wire7263;
wire wire7265;
wire wire7266;
wire wire7269;
wire wire7270;
wire wire7271;
wire wire7275;
wire wire7276;
wire wire7278;
wire wire7279;
wire wire7281;
wire wire7284;
wire wire7285;
wire wire7286;
wire wire7291;
wire wire7293;
wire wire7295;
wire wire7299;
wire wire7301;
wire wire7302;
wire wire7304;
wire wire7305;
wire wire7306;
wire wire7308;
wire wire7309;
wire wire7311;
wire wire7314;
wire wire7317;
wire wire7319;
wire wire7320;
wire wire7321;
wire wire7323;
wire wire7324;
wire wire7325;
wire wire7329;
wire wire7330;
wire wire7332;
wire wire7333;
wire wire7334;
wire wire7336;
wire wire7337;
wire wire7339;
wire wire7341;
wire wire7342;
wire wire7343;
wire wire7344;
wire wire7345;
wire wire7347;
wire wire7348;
wire wire7349;
wire wire7350;
wire wire7353;
wire wire7354;
wire wire7355;
wire wire7356;
wire wire7359;
wire wire7360;
wire wire7362;
wire wire7363;
wire wire7367;
wire wire7371;
wire wire7372;
wire wire7373;
wire wire7375;
wire wire7377;
wire wire7378;
wire wire7383;
wire wire7384;
wire wire7388;
wire wire7389;
wire wire7390;
wire wire7392;
wire wire7394;
wire wire7396;
wire wire7397;
wire wire7398;
wire wire7399;
wire wire7403;
wire wire7405;
wire wire7406;
wire wire7411;
wire wire7412;
wire wire7414;
wire wire7415;
wire wire7416;
wire wire7417;
wire wire7420;
wire wire7421;
wire wire7423;
wire wire7427;
wire wire7428;
wire wire7430;
wire wire7432;
wire wire7435;
wire wire7440;
wire wire7441;
wire wire7442;
wire wire7443;
wire wire7444;
wire wire7445;
wire wire7446;
wire wire7447;
wire wire7450;
wire wire7451;
wire wire7452;
wire wire7453;
wire wire7454;
wire wire7456;
wire wire7458;
wire wire7459;
wire wire7460;
wire wire7463;
wire wire7466;
wire wire7467;
wire wire7473;
wire wire7474;
wire wire7476;
wire wire7478;
wire wire7479;
wire wire7482;
wire wire7487;
wire wire7488;
wire wire7492;
wire wire7493;
wire wire7494;
wire wire7495;
wire wire7498;
wire wire7500;
wire wire7504;
wire wire7506;
wire wire7508;
wire wire7509;
wire wire7510;
wire wire7511;
wire wire7512;
wire wire7514;
wire wire7517;
wire wire7518;
wire wire7519;
wire wire7521;
wire wire7522;
wire wire7523;
wire wire7524;
wire wire7529;
wire wire7530;
wire wire7531;
wire wire7535;
wire wire7536;
wire wire7538;
wire wire7540;
wire wire7541;
wire wire7542;
wire wire7544;
wire wire7545;
wire wire7547;
wire wire7548;
wire wire7550;
wire wire7554;
wire wire7555;
wire wire7557;
wire wire7558;
wire wire7559;
wire wire7560;
wire wire7562;
wire wire7563;
wire wire7564;
wire wire7565;
wire wire7566;
wire wire7568;
wire wire7570;
wire wire7571;
wire wire7572;
wire wire7574;
wire wire7576;
wire wire7577;
wire wire7578;
wire wire7582;
wire wire7583;
wire wire7586;
wire wire7588;
wire wire7590;
wire wire7591;
wire wire7593;
wire wire7596;
wire wire7597;
wire wire7601;
wire wire7602;
wire wire7605;
wire wire7610;
wire wire7612;
wire wire7614;
wire wire7615;
wire wire7616;
wire wire7620;
wire wire7624;
wire wire7625;
wire wire7626;
wire wire7627;
wire wire7630;
wire wire7631;
wire wire7632;
wire wire7634;
wire wire7636;
wire wire7637;
wire wire7639;
wire wire7640;
wire wire7641;
wire wire7643;
wire wire7645;
wire wire7646;
wire wire7647;
wire wire7648;
wire wire7649;
wire wire7650;
wire wire7654;
wire wire7655;
wire wire7658;
wire wire7659;
wire wire7661;
wire wire7663;
wire wire7664;
wire wire7666;
wire wire7667;
wire wire7669;
wire wire7670;
wire wire7673;
wire wire7674;
wire wire7676;
wire wire7677;
wire wire7679;
wire wire7680;
wire wire7681;
wire wire7683;
wire wire7686;
wire wire7689;
wire wire7692;
wire wire7694;
wire wire7698;
wire wire7704;
wire wire7705;
wire wire7707;
wire wire7715;
wire wire7717;
wire wire7722;
wire wire7726;
wire wire7728;
wire wire7730;
wire wire7734;
wire wire7737;
wire wire7738;
wire wire7741;
wire wire7742;
wire wire7743;
wire wire7745;
wire wire7747;
wire wire7750;
wire wire7754;
wire wire7755;
wire wire7756;
wire wire7757;
wire wire7760;
wire wire7761;
wire wire7762;
wire wire7763;
wire wire7764;
wire wire7767;
wire wire7770;
wire wire7771;
wire wire7772;
wire wire7774;
wire wire7775;
wire wire7777;
wire wire7784;
wire wire7785;
wire wire7786;
wire wire7791;
wire wire7793;
wire wire7795;
wire wire7796;
wire wire7799;
wire wire7800;
wire wire7803;
wire wire7805;
wire wire7806;
wire wire7807;
wire wire7808;
wire wire7809;
wire wire7811;
wire wire7812;
wire wire7814;
wire wire7815;
wire wire7816;
wire wire7817;
wire wire7818;
wire wire7819;
wire wire7820;
wire wire7821;
wire wire7822;
assign o_1_ = ( wire6758 ) | ( wire6759 ) ;
 assign o_19_ = ( wire1867 ) | ( wire1870 ) | ( wire6767 ) | ( wire6770 ) ;
 assign o_2_ = ( n_n1165 ) | ( wire6806 ) | ( wire6807 ) | ( wire6808 ) ;
 assign o_0_ = ( n_n1081 ) | ( wire6914 ) | ( wire6915 ) | ( wire6929 ) ;
 assign o_29_ = ( wire1693 ) | ( wire6933 ) | ( wire6934 ) | ( wire6935 ) ;
 assign o_25_ = ( n_n1581 ) | ( n_n1603 ) | ( wire223 ) | ( wire6987 ) ;
 assign o_12_ = ( n_n685  &  wire1650  &  wire6991 ) | ( n_n685  &  wire1651  &  wire6991 ) ;
 assign o_26_ = ( wire238 ) | ( wire6994 ) | ( wire6998 ) | ( wire7005 ) ;
 assign o_11_ = ( n_n1394 ) | ( wire1617 ) | ( wire1619 ) | ( wire7021 ) ;
 assign o_27_ = ( n_n1628 ) | ( n_n1630 ) | ( n_n1631 ) | ( wire7040 ) ;
 assign o_14_ = ( wire225 ) | ( wire1588 ) ;
 assign o_28_ = ( n_n1971 ) | ( wire7043 ) | ( wire335  &  wire396 ) ;
 assign o_13_ = ( wire225 ) | ( n_n1011  &  n_n1074  &  n_n864 ) ;
 assign o_34_ = ( n_n1711 ) | ( wire7094 ) | ( wire7095 ) ;
 assign o_21_ = ( n_n1525 ) | ( wire1505 ) | ( wire1506 ) | ( wire7110 ) ;
 assign o_16_ = ( wire7118 ) | ( wire7119 ) | ( n_n1005  &  wire566 ) ;
 assign o_33_ = ( n_n1672 ) | ( n_n1670 ) | ( wire7187 ) | ( wire7190 ) ;
 assign o_22_ = ( n_n1530 ) | ( wire7210 ) | ( wire7211 ) | ( wire7223 ) ;
 assign o_15_ = ( i_7_  &  i_33_ ) ;
 assign o_32_ = ( n_n979  &  wire88  &  n_n1005 ) ;
 assign o_23_ = ( n_n1549 ) | ( n_n1552 ) | ( wire7270 ) | ( wire7271 ) ;
 assign o_18_ = ( n_n1445 ) | ( wire7301 ) | ( wire7302 ) | ( wire7345 ) ;
 assign o_31_ = ( wire7359 ) | ( i_22_  &  wire570 ) ;
 assign o_24_ = ( n_n2581 ) | ( n_n2838 ) | ( n_n1571 ) ;
 assign o_17_ = ( n_n1408 ) | ( n_n1409 ) | ( n_n1411 ) | ( wire7447 ) ;
 assign o_30_ = ( n_n1651 ) | ( wire7463 ) | ( i_24_  &  wire571 ) ;
 assign o_20_ = ( n_n1488 ) | ( wire7478 ) | ( wire7508 ) ;
 assign o_10_ = ( wire1031 ) | ( wire1043 ) | ( wire1044 ) | ( wire7519 ) ;
 assign o_9_ = ( wire7529 ) | ( wire7530 ) ;
 assign o_7_ = ( wire7540 ) | ( wire7541 ) | ( wire7547 ) | ( wire7548 ) ;
 assign o_8_ = ( wire7550 ) | ( n_n883  &  n_n966  &  n_n1012 ) ;
 assign o_5_ = ( n_n1272 ) | ( wire7615 ) | ( wire7616 ) | ( wire7639 ) ;
 assign o_6_ = ( n_n1330 ) | ( n_n1332 ) | ( n_n1323 ) | ( wire7683 ) ;
 assign o_3_ = ( n_n1187 ) | ( n_n1184 ) | ( wire7763 ) | ( wire7764 ) ;
 assign o_4_ = ( n_n1233 ) | ( wire56 ) | ( wire7821 ) | ( wire7822 ) ;
 assign n_n955 = ( i_9_  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n709 = ( (~ i_38_)  &  (~ i_37_) ) ;
 assign wire66 = ( i_40_  &  i_39_ ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire145 = ( o_15_ ) | ( n_n883  &  n_n1074  &  wire334 ) ;
 assign wire363 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  n_n1012 ) ;
 assign wire537 = ( n_n1014  &  wire45  &  n_n1009  &  wire37 ) ;
 assign wire543 = ( (~ i_40_)  &  i_39_ ) | ( i_39_  &  (~ i_38_) ) ;
 assign n_n1055 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n985 = ( (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n979 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign n_n515 = ( (~ i_7_)  &  wire471  &  wire80 ) ;
 assign n_n1008 = ( (~ i_40_)  &  (~ i_39_) ) ;
 assign n_n842 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n1067 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n982 = ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n990 = ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire88 = ( (~ i_40_)  &  (~ i_7_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire330 = ( i_40_  &  i_39_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n1373 = ( wire1890  &  wire6772 ) | ( wire1891  &  wire6772 ) ;
 assign n_n1164 = ( wire1852 ) | ( wire1853 ) | ( wire1854 ) | ( wire1855 ) ;
 assign n_n1165 = ( wire1844 ) | ( wire1846 ) | ( wire6793 ) | ( wire6794 ) ;
 assign wire48 = ( (~ i_21_)  &  i_15_ ) ;
 assign wire241 = ( i_40_  &  (~ i_39_)  &  n_n1074  &  n_n1061 ) ;
 assign wire432 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire491 = ( i_23_  &  i_24_  &  i_22_  &  i_19_ ) ;
 assign wire549 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign n_n1083 = ( n_n2838 ) | ( n_n2836 ) | ( wire6813 ) | ( wire6818 ) ;
 assign n_n978 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n883 = ( i_40_  &  (~ i_39_)  &  i_38_ ) ;
 assign n_n998 = ( i_34_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n1021 = ( (~ i_40_)  &  i_39_ ) ;
 assign n_n330 = ( (~ i_7_)  &  (~ i_5_)  &  i_13_ ) ;
 assign n_n969 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n2487 = ( n_n997  &  n_n793  &  n_n1048  &  n_n1047 ) ;
 assign n_n973 = ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign n_n158 = ( i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n2488 = ( n_n977  &  n_n793  &  n_n1048  &  n_n1047 ) ;
 assign n_n1084 = ( wire1805 ) | ( wire6831 ) | ( wire6832 ) ;
 assign n_n1777 = ( (~ i_7_)  &  wire50  &  wire6920 ) ;
 assign wire35 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n469 = ( (~ i_40_)  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1993 = ( wire88  &  n_n1002  &  n_n795 ) ;
 assign wire553 = ( (~ i_21_)  &  i_15_  &  n_n853 ) | ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign n_n2581 = ( wire88  &  n_n975  &  wire6938 ) ;
 assign n_n1971 = ( n_n971  &  n_n967  &  wire79  &  (~ wire115) ) ;
 assign n_n1581 = ( wire127 ) | ( wire6940 ) | ( wire6941 ) | ( wire6942 ) ;
 assign n_n1603 = ( wire185 ) | ( wire6964 ) | ( wire6965 ) ;
 assign wire173 = ( n_n1993 ) | ( n_n1986 ) | ( wire1666 ) ;
 assign wire223 = ( n_n1607 ) | ( wire1653 ) | ( wire1655 ) | ( wire6981 ) ;
 assign n_n685 = ( (~ i_7_)  &  i_5_  &  (~ i_0_) ) ;
 assign n_n2838 = ( (~ i_7_)  &  i_4_  &  n_n926  &  wire80 ) ;
 assign n_n2836 = ( (~ i_7_)  &  i_1_  &  n_n926  &  wire80 ) ;
 assign n_n1990 = ( n_n883  &  n_n970  &  wire79  &  wire318 ) ;
 assign n_n1951 = ( n_n971  &  n_n1072  &  wire79  &  wire318 ) ;
 assign wire555 = ( n_n1074  &  wire6828 ) | ( n_n1074  &  wire6897 ) ;
 assign n_n926 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n2213 = ( n_n998  &  n_n861  &  wire325 ) ;
 assign n_n1394 = ( wire1626 ) | ( wire92  &  wire1630 ) | ( wire92  &  wire7012 ) ;
 assign wire92 = ( i_40_  &  i_39_  &  n_n1009 ) ;
 assign wire319 = ( i_16_  &  n_n933  &  n_n1066 ) ;
 assign wire422 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_  &  (~ i_35_) ) ;
 assign wire470 = ( (~ i_12_)  &  wire82 ) ;
 assign wire556 = ( i_40_  &  (~ i_39_)  &  i_38_ ) | ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n761 = ( (~ i_21_)  &  i_15_  &  wire50  &  n_n850 ) ;
 assign n_n760 = ( (~ i_22_)  &  wire87  &  wire50 ) ;
 assign n_n1628 = ( n_n2487 ) | ( n_n2488 ) | ( wire173 ) | ( n_n1611 ) ;
 assign n_n1630 = ( wire174 ) | ( wire1610 ) | ( wire7025 ) | ( wire7026 ) ;
 assign n_n1631 = ( wire300 ) | ( wire127 ) | ( wire7029 ) | ( wire7030 ) ;
 assign wire175 = ( (~ i_22_)  &  n_n833  &  wire50  &  wire82 ) ;
 assign wire240 = ( (~ i_24_)  &  wire50  &  wire54  &  wire82 ) ;
 assign wire323 = ( (~ i_40_)  &  i_39_  &  n_n1009 ) ;
 assign wire559 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire225 = ( o_15_ ) | ( n_n968  &  n_n1074  &  wire59 ) ;
 assign n_n1011 = ( (~ i_39_)  &  (~ i_38_) ) ;
 assign n_n980 = ( i_5_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1006 = ( i_5_  &  (~ i_0_)  &  (~ i_32_) ) ;
 assign n_n989 = ( (~ i_15_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n983 = ( (~ i_34_)  &  i_33_  &  (~ i_36_) ) ;
 assign n_n1709 = ( wire1583 ) | ( wire1584 ) | ( wire7048 ) ;
 assign n_n1711 = ( n_n1716 ) | ( wire1575 ) | ( wire7053 ) | ( wire7071 ) ;
 assign wire445 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire560 = ( n_n979  &  n_n978 ) | ( n_n973  &  n_n1012 ) ;
 assign n_n865 = ( i_36_  &  i_35_  &  i_37_ ) ;
 assign n_n1525 = ( wire1518 ) | ( (~ i_0_)  &  wire1520 ) | ( (~ i_0_)  &  wire1521 ) ;
 assign wire47 = ( (~ i_7_)  &  (~ i_5_) ) ;
 assign n_n971 = ( i_36_  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign n_n1005 = ( (~ i_39_)  &  i_38_  &  i_37_ ) ;
 assign n_n997 = ( i_39_  &  i_38_  &  i_37_ ) ;
 assign n_n975 = ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n880 = ( i_40_  &  (~ i_38_) ) ;
 assign wire390 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  n_n629 ) ;
 assign wire411 = ( n_n842  &  n_n1074  &  wire7115 ) ;
 assign wire436 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  n_n865 ) ;
 assign wire526 = ( (~ i_3_)  &  (~ i_4_)  &  n_n1067  &  wire79 ) ;
 assign wire566 = ( i_40_  &  n_n979  &  n_n861 ) | ( (~ i_40_)  &  n_n861  &  n_n991 ) ;
 assign wire565 = ( i_37_  &  wire346  &  wire326 ) | ( (~ i_37_)  &  n_n1072  &  wire326 ) ;
 assign n_n1014 = ( i_40_  &  i_39_ ) ;
 assign n_n1528 = ( wire1402 ) | ( wire7193  &  wire7195 ) | ( wire7194  &  wire7195 ) ;
 assign n_n1530 = ( wire7204 ) | ( (~ i_38_)  &  (~ i_37_)  &  wire780 ) ;
 assign wire183 = ( wire330  &  n_n976  &  n_n668 ) ;
 assign wire251 = ( n_n983  &  n_n975  &  n_n668 ) ;
 assign wire335 = ( i_38_  &  n_n865  &  n_n1074 ) ;
 assign wire354 = ( (~ i_7_)  &  (~ i_31_)  &  i_33_  &  n_n1047 ) ;
 assign wire392 = ( n_n685  &  n_n874  &  n_n1052 ) ;
 assign n_n874 = ( (~ i_32_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n966 = ( (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign n_n862 = ( (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n1549 = ( wire1356 ) | ( wire1357 ) | ( wire1358 ) | ( wire7237 ) ;
 assign n_n1552 = ( wire7260 ) | ( wire7261 ) | ( wire46  &  wire810 ) ;
 assign wire490 = ( (~ i_34_)  &  (~ i_35_) ) ;
 assign n_n1445 = ( n_n1453 ) | ( n_n1452 ) | ( wire7329 ) ;
 assign wire346 = ( (~ i_39_)  &  i_38_ ) ;
 assign n_n1986 = ( (~ i_24_)  &  wire371  &  wire87  &  wire50 ) ;
 assign n_n837 = ( (~ i_24_)  &  wire50  &  wire82 ) ;
 assign wire245 = ( (~ i_24_)  &  wire87  &  wire50  &  wire54 ) ;
 assign wire364 = ( i_21_  &  i_22_  &  i_15_  &  wire35 ) ;
 assign wire371 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire570 = ( wire348  &  wire7350 ) | ( wire348  &  wire44  &  wire492 ) ;
 assign n_n1571 = ( wire223 ) | ( n_n1572 ) | ( wire7383 ) | ( wire7384 ) ;
 assign n_n1408 = ( n_n1414 ) | ( n_n1412 ) | ( wire7412 ) ;
 assign n_n1409 = ( n_n1416 ) | ( n_n1417 ) | ( wire7432 ) ;
 assign n_n1411 = ( wire7444 ) | ( wire7445 ) ;
 assign n_n968 = ( (~ i_36_)  &  i_35_  &  (~ i_37_) ) ;
 assign n_n819 = ( i_24_  &  (~ i_22_)  &  n_n1074  &  wire82 ) ;
 assign n_n1651 = ( wire1132 ) | ( wire7453 ) | ( wire7454 ) ;
 assign wire99 = ( i_24_  &  n_n968  &  n_n1074 ) ;
 assign wire365 = ( (~ i_21_)  &  i_15_  &  n_n853 ) ;
 assign wire572 = ( (~ i_40_)  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign wire571 = ( wire348  &  wire7350 ) | ( wire348  &  wire44  &  wire492 ) ;
 assign n_n1489 = ( wire1061 ) | ( wire1062 ) | ( wire7498 ) ;
 assign wire182 = ( (~ i_7_)  &  wire45  &  n_n693  &  wire6821 ) ;
 assign wire301 = ( wire371  &  n_n1023  &  n_n668 ) | ( n_n833  &  n_n1023  &  n_n668 ) ;
 assign wire574 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire575 = ( wire364  &  wire7512 ) | ( wire474  &  wire7517 ) ;
 assign n_n857 = ( n_n978  &  n_n1074  &  wire6731 ) ;
 assign n_n411 = ( i_23_  &  i_24_  &  i_22_ ) ;
 assign n_n1372 = ( wire478  &  wire6798 ) | ( wire407  &  wire39  &  wire6798 ) ;
 assign wire57 = ( wire1834 ) | ( i_18_  &  wire42 ) ;
 assign wire84 = ( n_n1055  &  n_n1048  &  n_n1047 ) ;
 assign wire416 = ( i_16_  &  n_n1055  &  n_n1048  &  n_n1047 ) ;
 assign wire512 = ( wire48  &  n_n978  &  n_n1074  &  wire6731 ) ;
 assign wire579 = ( (~ i_12_)  &  i_11_  &  i_15_  &  wire317 ) | ( i_12_  &  (~ i_11_)  &  i_15_  &  wire317 ) ;
 assign n_n1072 = ( i_40_  &  i_39_  &  i_38_ ) ;
 assign n_n937 = ( n_n1074  &  n_n949  &  wire7128 ) ;
 assign n_n1374 = ( i_19_  &  wire473  &  wire739 ) ;
 assign wire120 = ( i_40_  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign wire333 = ( n_n1001  &  n_n945  &  wire6789  &  wire7133 ) ;
 assign wire386 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  wire6907 ) ;
 assign wire583 = ( n_n1074  &  n_n949  &  wire7128 ) | ( n_n1074  &  n_n947  &  wire7128 ) ;
 assign wire581 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire146 = ( wire45  &  n_n693  &  wire7531 ) ;
 assign n_n698 = ( i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire131 = ( n_n1056  &  wire325  &  wire7626 ) ;
 assign wire402 = ( i_40_  &  i_36_  &  (~ i_35_)  &  i_38_ ) ;
 assign wire493 = ( (~ i_36_)  &  i_37_ ) ;
 assign wire495 = ( i_40_  &  i_39_  &  (~ i_37_) ) ;
 assign n_n1330 = ( wire882 ) | ( wire7643 ) | ( n_n334  &  wire619 ) ;
 assign n_n1332 = ( wire7650 ) | ( wire621  &  wire7649 ) ;
 assign n_n866 = ( i_40_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n1323 = ( wire536 ) | ( wire849 ) | ( wire7669 ) | ( wire7674 ) ;
 assign wire316 = ( i_38_  &  (~ i_37_) ) ;
 assign wire587 = ( n_n848  &  n_n945  &  n_n853 ) | ( n_n848  &  n_n945  &  n_n850 ) ;
 assign wire586 = ( wire94  &  wire106 ) | ( wire44  &  wire7679 ) ;
 assign n_n1187 = ( n_n1197 ) | ( n_n1196 ) | ( wire277 ) | ( wire7730 ) ;
 assign n_n1184 = ( n_n1203 ) | ( n_n1202 ) | ( wire7737 ) | ( wire7738 ) ;
 assign wire45 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign wire202 = ( i_28_ ) | ( i_29_ ) ;
 assign wire406 = ( (~ i_5_)  &  n_n462 ) ;
 assign n_n1233 = ( n_n1237 ) | ( n_n1239 ) | ( wire7793 ) ;
 assign n_n775 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_  &  n_n1047 ) ;
 assign n_n785 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_)  &  wire400 ) ;
 assign n_n1242 = ( wire129 ) | ( wire136  &  wire7816 ) | ( wire137  &  wire7816 ) ;
 assign wire469 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n528 = ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) ;
 assign n_n977 = ( (~ i_40_)  &  i_39_  &  i_38_ ) ;
 assign n_n888 = ( (~ i_34_)  &  i_35_  &  (~ i_37_) ) ;
 assign n_n313 = ( i_13_  &  wire50  &  wire315 ) ;
 assign wire227 = ( n_n330  &  n_n989  &  n_n1066  &  wire6887 ) ;
 assign wire508 = ( (~ i_7_)  &  wire45  &  n_n1061  &  wire115 ) ;
 assign wire594 = ( i_40_  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1326 = ( wire227 ) | ( wire869 ) | ( wire7654 ) | ( wire7655 ) ;
 assign wire68 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_37_) ) ;
 assign wire174 = ( wire504  &  n_n960 ) | ( wire367  &  wire479 ) ;
 assign wire300 = ( i_39_  &  i_38_  &  wire430 ) | ( i_40_  &  (~ i_38_)  &  wire430 ) ;
 assign wire504 = ( n_n793  &  n_n1047  &  wire78  &  wire6858 ) ;
 assign n_n1283 = ( wire174 ) | ( wire957 ) | ( wire7577 ) | ( wire7578 ) ;
 assign n_n833 = ( i_39_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire176 = ( (~ i_22_)  &  n_n833  &  wire87  &  wire50 ) ;
 assign wire395 = ( wire80  &  wire7145 ) ;
 assign wire598 = ( wire87  &  wire50 ) | ( wire50  &  wire82 ) ;
 assign wire596 = ( (~ i_24_)  &  wire87  &  wire50 ) | ( (~ i_24_)  &  wire50  &  wire82 ) ;
 assign wire595 = ( n_n926 ) | ( wire983 ) ;
 assign n_n1280 = ( wire7559 ) | ( wire7560 ) | ( n_n833  &  wire596 ) ;
 assign n_n1052 = ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n1064 = ( i_40_  &  (~ i_39_) ) ;
 assign n_n525 = ( (~ i_13_)  &  wire50  &  wire315 ) ;
 assign wire148 = ( (~ i_7_)  &  n_n1052  &  wire80  &  wire464 ) ;
 assign wire329 = ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign wire357 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1009 ) ;
 assign wire408 = ( i_13_  &  wire315 ) ;
 assign wire441 = ( i_40_  &  (~ i_39_)  &  i_38_  &  i_37_ ) ;
 assign wire542 = ( n_n842  &  n_n966  &  n_n1073  &  n_n843 ) ;
 assign n_n764 = ( (~ i_22_)  &  wire50  &  wire82 ) ;
 assign wire600 = ( (~ i_21_)  &  i_15_  &  n_n853 ) | ( (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign n_n1272 = ( n_n1280 ) | ( wire7570 ) | ( wire7571 ) | ( wire7574 ) ;
 assign n_n799 = ( (~ i_40_)  &  i_39_  &  (~ i_38_) ) ;
 assign n_n1237 = ( wire7774 ) | ( wire7775 ) | ( wire366  &  wire662 ) ;
 assign n_n1239 = ( wire203 ) | ( wire7784 ) | ( wire7785 ) | ( wire7786 ) ;
 assign wire398 = ( n_n861  &  n_n710  &  n_n715 ) ;
 assign wire602 = ( i_40_  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n1235 = ( wire7799 ) | ( wire7800 ) | ( n_n795  &  wire612 ) ;
 assign n_n861 = ( (~ i_7_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n793 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign wire420 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire604 = ( wire160 ) | ( wire7807  &  wire7809 ) | ( wire7808  &  wire7809 ) ;
 assign wire407 = ( (~ i_5_)  &  i_17_  &  i_16_  &  i_15_ ) ;
 assign n_n1048 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire349 = ( i_24_  &  i_22_ ) ;
 assign wire607 = ( i_12_  &  (~ i_18_) ) | ( i_11_  &  (~ i_18_) ) | ( i_11_  &  (~ i_19_) ) ;
 assign n_n1094 = ( wire1789 ) | ( (~ i_23_)  &  wire1791 ) | ( (~ i_23_)  &  wire1792 ) ;
 assign n_n2837 = ( (~ i_7_)  &  i_3_  &  n_n926  &  wire80 ) ;
 assign n_n1958 = ( (~ i_7_)  &  i_4_  &  n_n833  &  wire80 ) ;
 assign n_n1956 = ( (~ i_7_)  &  i_3_  &  n_n833  &  wire80 ) ;
 assign n_n1957 = ( (~ i_7_)  &  i_1_  &  n_n833  &  wire80 ) ;
 assign n_n964 = ( (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n1073 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign n_n1009 = ( (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1002 = ( (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign n_n960 = ( i_39_  &  i_38_ ) ;
 assign n_n1001 = ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n993 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire81 = ( (~ i_38_)  &  i_37_ ) ;
 assign wire46 = ( (~ i_32_)  &  i_33_ ) ;
 assign wire382 = ( (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n933 = ( i_17_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1066 = ( (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n967 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire86 = ( i_11_  &  i_15_ ) ;
 assign n_n1074 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign n_n642 = ( i_17_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1047 = ( (~ i_34_)  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n976 = ( i_33_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign n_n1015 = ( i_39_  &  (~ i_38_) ) ;
 assign n_n795 = ( i_39_  &  (~ i_38_)  &  i_37_ ) ;
 assign n_n848 = ( i_21_  &  i_22_  &  i_15_ ) ;
 assign n_n945 = ( i_24_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n853 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n559 = ( n_n848  &  n_n945  &  n_n853 ) ;
 assign wire87 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign wire320 = ( (~ i_31_)  &  (~ i_34_)  &  i_33_  &  (~ i_35_) ) ;
 assign n_n535 = ( i_16_  &  wire87  &  wire320 ) ;
 assign wire471 = ( (~ i_3_)  &  (~ i_4_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n949 = ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign n_n460 = ( n_n979  &  n_n949  &  wire7405 ) ;
 assign n_n1061 = ( i_36_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1023 = ( (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire359 = ( i_40_  &  (~ i_39_)  &  n_n985 ) ;
 assign n_n952 = ( i_40_  &  (~ i_39_)  &  n_n985  &  n_n1023 ) ;
 assign wire317 = ( i_9_  &  (~ i_5_) ) ;
 assign wire78 = ( i_12_  &  i_15_ ) ;
 assign n_n947 = ( (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign n_n935 = ( n_n1074  &  n_n947  &  wire7128 ) ;
 assign n_n329 = ( n_n330  &  n_n989  &  n_n1066 ) ;
 assign n_n527 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign n_n710 = ( (~ i_4_)  &  (~ i_1_)  &  i_0_ ) ;
 assign wire400 = ( i_40_  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign n_n688 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign n_n462 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign n_n700 = ( (~ i_15_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n492 = ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire100 = ( i_38_  &  i_37_ ) ;
 assign n_n1065 = ( i_36_  &  i_38_  &  i_37_ ) ;
 assign n_n488 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n453 = ( i_3_  &  i_0_  &  (~ i_32_) ) ;
 assign wire77 = ( (~ i_32_)  &  i_33_  &  n_n998 ) ;
 assign n_n1012 = ( (~ i_36_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire334 = ( i_35_  &  (~ i_37_) ) ;
 assign wire378 = ( (~ i_5_)  &  (~ i_15_) ) ;
 assign n_n884 = ( (~ i_5_)  &  (~ i_13_)  &  (~ i_15_) ) ;
 assign wire326 = ( i_36_  &  (~ i_35_) ) ;
 assign n_n970 = ( i_36_  &  (~ i_35_)  &  i_37_ ) ;
 assign n_n928 = ( i_9_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign n_n951 = ( i_9_  &  (~ i_5_)  &  i_12_ ) ;
 assign n_n860 = ( i_9_  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign n_n560 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1012 ) ;
 assign n_n484 = ( (~ i_16_)  &  i_15_  &  n_n492  &  wire76 ) ;
 assign wire60 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire76 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire103 = ( wire401 ) | ( wire465 ) ;
 assign wire531 = ( n_n979  &  n_n949  &  n_n791 ) ;
 assign wire611 = ( n_n492  &  wire76  &  wire352 ) | ( n_n492  &  wire76  &  wire7414 ) ;
 assign n_n1416 = ( wire1179 ) | ( wire1181 ) | ( wire1183 ) | ( wire7417 ) ;
 assign wire430 = ( n_n793  &  wire86  &  n_n1047  &  wire6850 ) ;
 assign wire612 = ( n_n861  &  wire613 ) | ( (~ i_40_)  &  n_n998  &  n_n861 ) ;
 assign wire462 = ( (~ i_5_)  &  i_31_  &  (~ i_36_)  &  wire45 ) ;
 assign n_n1203 = ( wire274 ) | ( i_38_  &  wire462 ) | ( (~ i_37_)  &  wire462 ) ;
 assign n_n1202 = ( wire271 ) | ( wire272 ) | ( i_39_  &  wire462 ) ;
 assign n_n777 = ( i_11_  &  i_15_  &  n_n793  &  wire6850 ) ;
 assign n_n781 = ( (~ i_17_)  &  (~ i_16_)  &  n_n1048  &  wire87 ) ;
 assign wire37 = ( i_17_ ) | ( i_16_ ) ;
 assign wire64 = ( n_n1055  &  n_n1047 ) | ( n_n1047  &  wire6851 ) ;
 assign wire94 = ( i_40_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign wire106 = ( n_n848  &  n_n945  &  n_n853 ) | ( n_n848  &  n_n945  &  n_n850 ) ;
 assign wire321 = ( (~ i_31_)  &  wire45 ) ;
 assign wire614 = ( wire1786 ) | ( (~ i_18_)  &  wire35 ) ;
 assign n_n1057 = ( (~ i_3_)  &  i_4_  &  (~ i_32_) ) ;
 assign n_n1056 = ( (~ i_34_)  &  i_33_  &  i_36_ ) ;
 assign wire61 = ( i_12_ ) | ( i_11_ ) ;
 assign n_n629 = ( (~ i_7_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire410 = ( (~ i_1_)  &  i_0_ ) ;
 assign wire50 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire315 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign n_n162 = ( n_n979  &  n_n947  &  wire7390 ) ;
 assign n_n991 = ( (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign n_n334 = ( i_13_  &  wire76  &  wire315 ) ;
 assign n_n801 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_28_) ) ;
 assign n_n428 = ( i_24_  &  i_22_  &  (~ i_32_) ) ;
 assign n_n427 = ( i_40_  &  i_39_  &  n_n1009  &  n_n1023 ) ;
 assign n_n843 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign n_n791 = ( (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n459 = ( n_n979  &  n_n947  &  wire7399 ) ;
 assign n_n905 = ( n_n979  &  n_n907  &  wire6716 ) ;
 assign n_n1414 = ( wire1204 ) | ( wire1205 ) | ( wire1206 ) | ( wire7392 ) ;
 assign n_n1412 = ( wire1196 ) | ( wire1197 ) | ( wire1198 ) | ( wire7403 ) ;
 assign wire467 = ( i_28_  &  (~ i_29_)  &  n_n1066  &  wire7122 ) ;
 assign wire616 = ( wire531 ) | ( n_n162 ) | ( n_n164 ) | ( wire1192 ) ;
 assign wire615 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n475 = ( (~ i_16_)  &  i_15_  &  n_n488  &  wire76 ) ;
 assign n_n164 = ( n_n979  &  n_n949  &  wire7406 ) ;
 assign n_n1417 = ( wire7427 ) | ( n_n1011  &  n_n1012  &  wire696 ) ;
 assign wire113 = ( n_n488  &  wire76  &  wire352 ) | ( n_n488  &  wire76  &  wire7414 ) ;
 assign wire617 = ( wire401 ) | ( wire465 ) ;
 assign wire506 = ( i_40_  &  i_39_  &  n_n1052  &  wire315 ) ;
 assign wire619 = ( i_40_  &  i_39_  &  n_n1073 ) | ( i_39_  &  (~ i_38_)  &  n_n1073 ) | ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  n_n1073 ) ;
 assign wire433 = ( n_n945  &  n_n860  &  wire6789 ) ;
 assign wire621 = ( wire622  &  wire7647 ) | ( wire44  &  wire7648 ) ;
 assign n_n2439 = ( n_n861  &  n_n1002  &  wire7330 ) ;
 assign wire624 = ( (~ i_34_)  &  i_36_  &  i_37_ ) | ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire623 = ( i_25_ ) | ( (~ i_26_) ) ;
 assign wire352 = ( (~ i_16_)  &  i_15_ ) ;
 assign wire421 = ( (~ i_32_)  &  i_33_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire518 = ( n_n1023  &  n_n1065  &  n_n1057 ) ;
 assign wire524 = ( n_n1057  &  n_n843  &  n_n1053 ) ;
 assign wire627 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n1197 = ( wire294 ) | ( wire295 ) | ( wire297 ) | ( wire7715 ) ;
 assign wire36 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign n_n1193 = ( wire451 ) | ( wire454 ) | ( wire459 ) | ( wire7692 ) ;
 assign wire633 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign n_n1195 = ( wire443 ) | ( wire444 ) | ( wire446 ) ;
 assign wire154 = ( wire45  &  n_n1061  &  wire7394 ) ;
 assign wire635 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire65 = ( i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire637 = ( n_n1055  &  n_n1047 ) | ( n_n1047  &  wire638 ) ;
 assign n_n1135 = ( wire1912 ) | ( wire1913 ) | ( wire6734 ) ;
 assign n_n1053 = ( i_34_  &  i_33_  &  (~ i_35_) ) ;
 assign n_n582 = ( (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign n_n850 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire367 = ( i_12_  &  i_15_  &  n_n793 ) ;
 assign n_n771 = ( i_12_  &  i_15_  &  n_n793  &  wire6858 ) ;
 assign wire368 = ( i_11_  &  i_15_  &  n_n793 ) ;
 assign wire479 = ( n_n1048  &  n_n1047  &  wire6859 ) ;
 assign wire369 = ( wire50  &  wire82 ) ;
 assign wire393 = ( n_n1052  &  n_n1057  &  n_n1053 ) ;
 assign wire468 = ( (~ i_31_)  &  wire45  &  wire7389 ) ;
 assign wire83 = ( n_n979  &  n_n791  &  wire6976 ) ;
 assign wire356 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_)  &  n_n967 ) ;
 assign wire643 = ( i_12_  &  i_15_  &  n_n793 ) | ( i_11_  &  i_15_  &  n_n793 ) ;
 assign n_n1285 = ( wire950 ) | ( wire952 ) | ( wire7582 ) | ( wire7583 ) ;
 assign wire486 = ( i_15_  &  wire35 ) ;
 assign wire648 = ( n_n1048  &  wire87  &  (~ wire37) ) | ( n_n1048  &  (~ wire37)  &  wire82 ) ;
 assign wire646 = ( n_n1072  &  n_n1073 ) | ( n_n1055  &  n_n1047 ) ;
 assign n_n923 = ( i_39_  &  (~ i_36_)  &  i_38_ ) ;
 assign n_n1196 = ( wire286 ) | ( wire287 ) | ( wire288 ) | ( wire289 ) ;
 assign n_n1068 = ( i_17_  &  i_16_  &  i_15_ ) ;
 assign wire303 = ( i_39_  &  i_38_  &  n_n968  &  n_n1074 ) ;
 assign wire520 = ( n_n1014  &  n_n874  &  n_n1009  &  (~ wire73) ) ;
 assign wire655 = ( (~ i_9_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_9_)  &  (~ i_5_)  &  i_11_ ) ;
 assign n_n864 = ( i_36_  &  i_35_  &  (~ i_37_) ) ;
 assign wire79 = ( (~ i_7_)  &  (~ i_32_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire238 = ( i_2_  &  wire835 ) ;
 assign wire336 = ( i_40_  &  i_39_  &  n_n966  &  n_n993 ) ;
 assign n_n458 = ( i_2_  &  i_0_  &  (~ i_32_) ) ;
 assign n_n643 = ( i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign n_n1611 = ( wire176 ) | ( wire1681 ) | ( wire1682 ) ;
 assign n_n836 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire394 = ( i_40_  &  (~ i_39_)  &  n_n1065 ) ;
 assign wire660 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire366 = ( (~ i_40_)  &  i_39_  &  (~ i_38_)  &  n_n1012 ) ;
 assign wire662 = ( wire46  &  wire43 ) | ( wire53  &  wire7772 ) ;
 assign wire54 = ( i_39_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire80 = ( (~ i_32_)  &  i_34_  &  i_33_  &  (~ i_35_) ) ;
 assign wire325 = ( i_40_  &  i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire463 = ( (~ i_14_)  &  wire87  &  wire351 ) ;
 assign wire135 = ( i_3_ ) | ( i_4_ ) ;
 assign wire666 = ( (~ i_40_)  &  i_38_ ) | ( i_39_  &  i_38_ ) ;
 assign wire665 = ( (~ i_40_)  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire664 = ( (~ i_5_)  &  (~ i_38_)  &  i_37_ ) | ( i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire153 = ( n_n977  &  n_n1074  &  n_n864 ) ;
 assign wire184 = ( (~ i_32_)  &  i_33_  &  n_n991  &  wire6773 ) ;
 assign wire187 = ( (~ i_32_)  &  i_33_  &  n_n991  &  wire6774 ) ;
 assign wire667 = ( i_25_ ) | ( i_26_ ) ;
 assign wire458 = ( i_40_  &  (~ i_5_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire669 = ( (~ i_30_)  &  i_29_ ) | ( i_28_  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) ;
 assign wire668 = ( (~ i_30_)  &  i_29_ ) | ( i_28_  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) | ( (~ i_28_)  &  (~ i_29_) ) ;
 assign wire73 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) ;
 assign wire327 = ( i_40_  &  i_39_  &  i_38_  &  n_n1073 ) ;
 assign wire670 = ( i_9_  &  i_17_  &  i_15_ ) | ( i_9_  &  i_16_  &  i_15_ ) | ( i_17_  &  i_16_  &  i_15_ ) ;
 assign wire671 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_37_) ) ;
 assign wire672 = ( wire371 ) | ( wire54 ) ;
 assign wire529 = ( i_30_  &  i_29_  &  wire76  &  n_n801 ) ;
 assign wire370 = ( wire87  &  wire50 ) ;
 assign n_n918 = ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign n_n556 = ( n_n848  &  n_n945  &  n_n850 ) ;
 assign n_n798 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_ ) ;
 assign wire110 = ( (~ i_17_) ) | ( (~ i_16_) ) ;
 assign n_n859 = ( i_11_  &  i_18_  &  i_15_ ) ;
 assign wire351 = ( i_17_  &  i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire674 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire403 = ( (~ i_40_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire676 = ( wire1160 ) | ( n_n1001  &  wire677 ) ;
 assign wire675 = ( i_3_ ) | ( i_1_ ) ;
 assign wire69 = ( (~ i_32_)  &  n_n1066  &  wire318 ) | ( (~ i_32_)  &  n_n1066  &  wire7397 ) ;
 assign wire332 = ( i_4_  &  i_0_  &  wire45 ) ;
 assign wire680 = ( n_n1023  &  wire681 ) | ( (~ i_32_)  &  n_n1023  &  wire410 ) ;
 assign wire679 = ( n_n1021  &  n_n862 ) | ( n_n960  &  n_n1012 ) ;
 assign wire678 = ( i_40_  &  i_39_  &  n_n1061 ) | ( i_40_  &  (~ i_39_)  &  n_n1065 ) ;
 assign wire413 = ( (~ i_34_)  &  (~ i_36_)  &  i_35_  &  wire7227 ) ;
 assign wire684 = ( (~ i_32_)  &  n_n1023  &  wire7397 ) | ( (~ i_32_)  &  n_n1023  &  wire7750 ) ;
 assign wire484 = ( i_9_  &  (~ i_5_)  &  i_12_  &  i_15_ ) ;
 assign n_n1091 = ( wire1766 ) | ( wire6868 ) | ( wire6869 ) | ( wire6870 ) ;
 assign n_n1113 = ( n_n837  &  wire371 ) | ( n_n837  &  wire54 ) ;
 assign wire244 = ( n_n330  &  n_n926  &  n_n989  &  n_n1066 ) ;
 assign wire688 = ( wire87  &  wire50 ) | ( wire50  &  wire82 ) ;
 assign n_n1081 = ( n_n1091 ) | ( wire6878 ) | ( wire6879 ) ;
 assign n_n1088 = ( n_n1986 ) | ( wire1751 ) | ( wire6886 ) ;
 assign n_n1086 = ( wire149 ) | ( wire155 ) | ( wire6894 ) ;
 assign n_n1108 = ( n_n1971 ) | ( n_n1074  &  wire711  &  wire6897 ) ;
 assign wire464 = ( (~ i_3_)  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire689 = ( i_30_  &  (~ i_28_)  &  i_29_  &  wire47 ) | ( (~ i_30_)  &  i_28_  &  (~ i_29_)  &  wire47 ) ;
 assign wire132 = ( n_n1074  &  wire87  &  wire6908 ) | ( n_n1074  &  wire82  &  wire6908 ) ;
 assign wire690 = ( n_n1048  &  wire87  &  (~ wire37) ) | ( n_n1048  &  (~ wire37)  &  wire82 ) ;
 assign n_n927 = ( i_16_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire82 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign n_n773 = ( (~ i_17_)  &  (~ i_16_)  &  n_n1048  &  wire82 ) ;
 assign n_n715 = ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire337 = ( i_40_  &  i_39_  &  n_n985  &  wire80 ) ;
 assign wire344 = ( i_9_  &  (~ i_7_) ) ;
 assign wire692 = ( (~ i_12_)  &  n_n642 ) | ( (~ i_12_)  &  n_n643 ) | ( n_n642  &  wire693 ) | ( n_n643  &  wire693 ) ;
 assign wire696 = ( n_n484 ) | ( wire113 ) | ( wire1173 ) | ( wire1174 ) ;
 assign wire695 = ( n_n492  &  wire76  &  wire352 ) | ( n_n488  &  wire76  &  wire352 ) ;
 assign wire102 = ( wire43 ) | ( wire1291 ) ;
 assign wire697 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_40_  &  i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire509 = ( i_40_  &  (~ i_39_)  &  n_n862 ) ;
 assign wire396 = ( (~ i_7_)  &  (~ i_3_)  &  i_4_  &  n_n843 ) ;
 assign wire342 = ( i_40_  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire380 = ( i_18_  &  wire36 ) ;
 assign wire702 = ( (~ i_40_)  &  i_39_  &  i_38_  &  (~ i_37_) ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire701 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire700 = ( n_n1048  &  n_n1047  &  n_n527 ) | ( n_n1048  &  n_n1047  &  wire6884 ) ;
 assign n_n783 = ( i_12_  &  i_15_  &  n_n793  &  wire6968 ) ;
 assign wire376 = ( (~ i_7_)  &  (~ i_32_) ) ;
 assign n_n668 = ( (~ i_7_)  &  i_5_  &  (~ i_32_) ) ;
 assign n_n550 = ( n_n1068  &  (~ wire73)  &  wire7309 ) ;
 assign wire401 = ( i_40_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire704 = ( wire855 ) | ( wire315  &  wire856 ) | ( wire315  &  wire857 ) ;
 assign wire706 = ( wire133 ) | ( i_18_  &  wire35 ) ;
 assign wire710 = ( wire371 ) | ( wire54 ) ;
 assign wire149 = ( wire1749 ) | ( i_0_  &  wire79  &  wire6888 ) ;
 assign wire155 = ( wire1747 ) | ( i_0_  &  wire79  &  wire6889 ) ;
 assign wire383 = ( (~ i_36_)  &  (~ i_37_) ) ;
 assign wire429 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  wire6897 ) ;
 assign wire711 = ( i_37_  &  n_n883  &  wire326 ) | ( (~ i_37_)  &  n_n1072  &  wire326 ) ;
 assign n_n1577 = ( n_n1108 ) | ( wire155 ) | ( wire7362 ) | ( wire7363 ) ;
 assign wire713 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) | ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) | ( (~ i_36_)  &  i_38_  &  i_37_ ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign n_n1488 = ( wire1104 ) | ( (~ i_15_)  &  wire1106 ) | ( (~ i_15_)  &  wire1107 ) ;
 assign wire718 = ( wire1099 ) | ( wire7473 ) | ( wire7474 ) ;
 assign wire717 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire139 = ( i_40_  &  i_38_  &  n_n979 ) | ( (~ i_38_)  &  i_37_  &  n_n979 ) ;
 assign n_n1453 = ( wire1277 ) | ( wire7311 ) | ( n_n559  &  wire139 ) ;
 assign wire488 = ( (~ i_31_)  &  i_33_ ) ;
 assign wire723 = ( i_16_  &  wire87  &  wire320 ) | ( i_16_  &  wire320  &  wire82 ) ;
 assign n_n1452 = ( wire7319 ) | ( wire7320 ) | ( wire7321 ) ;
 assign wire724 = ( wire402 ) | ( wire1269 ) ;
 assign wire727 = ( i_18_  &  wire35 ) | ( n_n860  &  wire61 ) ;
 assign wire473 = ( n_n985  &  n_n1064  &  n_n1023  &  wire7124 ) ;
 assign n_n1277 = ( wire925 ) | ( wire926 ) | ( wire927 ) | ( wire7605 ) ;
 assign n_n693 = ( i_36_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire361 = ( (~ i_34_)  &  i_33_  &  (~ i_35_)  &  wire7122 ) ;
 assign wire737 = ( wire450  &  wire38 ) | ( wire351  &  wire738 ) ;
 assign wire739 = ( wire484 ) | ( i_18_  &  wire36 ) ;
 assign wire740 = ( i_39_  &  i_38_  &  i_37_ ) | ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign n_n1134 = ( wire6740 ) | ( wire6741 ) | ( (~ n_n1055)  &  wire462 ) ;
 assign wire742 = ( wire363 ) | ( wire303 ) | ( wire1901 ) | ( wire1902 ) ;
 assign wire741 = ( i_37_  &  n_n973  &  n_n964 ) | ( (~ i_37_)  &  n_n964  &  n_n967 ) ;
 assign n_n673 = ( (~ i_31_)  &  n_n1047  &  wire7191  &  wire7201 ) ;
 assign wire124 = ( i_40_  &  (~ i_38_)  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire744 = ( (~ i_24_)  &  wire87  &  wire50 ) | ( (~ i_24_)  &  wire50  &  wire82 ) ;
 assign wire535 = ( (~ i_30_)  &  (~ i_29_)  &  wire76  &  n_n798 ) ;
 assign wire748 = ( n_n985  &  (~ n_n1014) ) | ( i_35_  &  wire749 ) ;
 assign n_n790 = ( i_11_  &  i_15_  &  n_n793  &  wire6974 ) ;
 assign wire166 = ( (~ i_12_) ) | ( (~ i_11_) ) | ( (~ i_15_) ) ;
 assign wire752 = ( n_n979  &  n_n861 ) | ( (~ i_40_)  &  n_n861  &  n_n991 ) ;
 assign wire140 = ( wire382  &  n_n976  &  wire458  &  wire7154 ) ;
 assign wire156 = ( wire36  &  wire80  &  wire7145  &  wire7146 ) ;
 assign wire494 = ( (~ i_7_)  &  (~ i_5_)  &  i_29_ ) ;
 assign wire758 = ( i_34_  &  n_n1073  &  wire46 ) | ( (~ i_34_)  &  wire46  &  wire6731 ) ;
 assign n_n765 = ( (~ i_21_)  &  i_15_  &  n_n853  &  wire50 ) ;
 assign n_n907 = ( (~ i_5_)  &  (~ i_12_)  &  (~ i_11_) ) ;
 assign wire761 = ( (~ i_36_)  &  i_38_  &  i_37_  &  n_n1008 ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_)  &  n_n1008 ) ;
 assign wire763 = ( i_40_  &  (~ i_39_)  &  (~ i_36_)  &  i_37_ ) | ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire762 = ( wire86  &  wire320  &  n_n860 ) | ( wire320  &  wire78  &  n_n860 ) ;
 assign wire766 = ( n_n861  &  wire767 ) | ( (~ i_40_)  &  n_n861  &  wire100 ) ;
 assign wire348 = ( (~ i_23_)  &  n_n978  &  n_n1074  &  wire6731 ) ;
 assign n_n1607 = ( wire1661 ) | ( wire1662 ) | ( wire6970 ) | ( wire6971 ) ;
 assign wire101 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire127 = ( n_n775  &  n_n781 ) | ( wire329  &  wire348 ) ;
 assign wire772 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) ;
 assign wire373 = ( (~ i_40_)  &  (~ i_38_) ) ;
 assign n_n1575 = ( wire7367 ) | ( wire7371 ) | ( i_2_  &  wire835 ) ;
 assign wire775 = ( n_n969  &  wire334 ) | ( (~ i_36_)  &  n_n1014  &  wire334 ) ;
 assign wire461 = ( i_16_  &  n_n933  &  n_n1066  &  wire7132 ) ;
 assign wire777 = ( n_n926 ) | ( wire1487 ) ;
 assign n_n1672 = ( wire1489 ) | ( wire7129 ) | ( wire7139 ) | ( wire7140 ) ;
 assign n_n1572 = ( n_n1577 ) | ( n_n1575 ) | ( wire7375 ) ;
 assign wire780 = ( wire354  &  wire781 ) | ( wire354  &  wire7200 ) | ( wire354  &  wire7201 ) ;
 assign wire779 = ( (~ i_40_)  &  i_39_  &  i_35_  &  i_38_ ) | ( i_40_  &  (~ i_39_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire476 = ( i_24_  &  (~ i_22_)  &  n_n1074 ) ;
 assign wire782 = ( n_n998  &  n_n973 ) | ( n_n969  &  n_n888 ) ;
 assign wire786 = ( n_n926  &  wire67 ) | ( n_n923  &  wire7150 ) ;
 assign wire787 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign n_n1580 = ( wire6950 ) | ( wire6951 ) | ( wire6952 ) ;
 assign wire59 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) | ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign wire788 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_ ) | ( i_40_  &  i_39_  &  (~ i_38_) ) ;
 assign wire795 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) | ( (~ i_15_) ) ;
 assign wire794 = ( i_39_ ) | ( i_38_ ) | ( (~ i_37_) ) ;
 assign n_n1716 = ( wire7062 ) | ( wire76  &  wire826 ) ;
 assign wire158 = ( i_11_  &  wire46  &  n_n991  &  wire325 ) ;
 assign n_n1670 = ( wire1443 ) | ( wire7171 ) | ( wire7175 ) | ( wire7176 ) ;
 assign wire185 = ( wire6956 ) | ( wire6957 ) | ( wire6958 ) ;
 assign wire803 = ( wire490  &  n_n700 ) | ( n_n1074  &  wire326 ) ;
 assign wire806 = ( (~ i_12_)  &  (~ i_11_) ) | ( (~ i_9_)  &  (~ i_16_) ) ;
 assign wire805 = ( n_n880  &  wire45 ) | ( wire316  &  wire421 ) ;
 assign wire808 = ( i_3_ ) | ( i_4_ ) | ( i_1_ ) ;
 assign wire807 = ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire811 = ( i_34_  &  n_n1073  &  wire46 ) | ( (~ i_34_)  &  wire46  &  wire7258 ) ;
 assign wire810 = ( wire464  &  wire7256 ) | ( n_n1047  &  wire7257 ) ;
 assign wire809 = ( (~ i_38_)  &  wire464 ) | ( i_2_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire814 = ( wire63 ) | ( i_9_  &  (~ i_5_)  &  (~ i_15_) ) ;
 assign wire450 = ( i_9_  &  (~ i_14_) ) ;
 assign wire817 = ( n_n971  &  n_n977 ) | ( wire818  &  wire7074 ) ;
 assign wire465 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire475 = ( i_24_  &  n_n968  &  n_n1074  &  wire7452 ) ;
 assign wire822 = ( (~ i_40_)  &  i_39_  &  i_38_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_) ) ;
 assign wire825 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) | ( (~ i_40_)  &  i_39_  &  n_n1009 ) ;
 assign wire826 = ( wire1570 ) | ( (~ wire61)  &  wire1571 ) | ( (~ wire61)  &  wire7058 ) ;
 assign wire38 = ( i_17_  &  (~ i_32_)  &  i_33_ ) | ( i_16_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire39 = ( (~ i_12_)  &  i_11_ ) | ( i_12_  &  (~ i_11_) ) ;
 assign wire42 = ( i_9_  &  (~ i_5_)  &  i_12_ ) | ( i_9_  &  (~ i_5_)  &  i_11_ ) ;
 assign wire43 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_  &  i_29_ ) | ( (~ i_7_)  &  (~ i_5_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire44 = ( wire469 ) | ( i_18_  &  wire35 ) ;
 assign wire53 = ( (~ i_30_)  &  i_29_ ) | ( i_30_  &  (~ i_29_) ) ;
 assign wire55 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire304 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire63 = ( i_9_  &  (~ i_5_)  &  (~ i_12_) ) | ( i_9_  &  (~ i_5_)  &  (~ i_11_) ) ;
 assign wire67 = ( (~ i_14_) ) | ( (~ i_12_) ) ;
 assign wire318 = ( i_1_  &  i_0_ ) ;
 assign wire492 = ( (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign wire70 = ( wire1795 ) | ( (~ i_21_)  &  wire1797 ) | ( (~ i_21_)  &  wire1798 ) ;
 assign wire104 = ( n_n642  &  wire7818 ) | ( n_n643  &  wire7818 ) | ( n_n643  &  wire7819 ) ;
 assign wire115 = ( (~ i_10_) ) | ( (~ i_27_) ) ;
 assign wire302 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  wire6828 ) ;
 assign wire121 = ( (~ i_40_)  &  (~ i_38_)  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire830 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) | ( (~ i_40_)  &  i_39_  &  n_n1009 ) ;
 assign wire829 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire831 = ( n_n1048  &  wire87  &  (~ wire37) ) | ( n_n1048  &  (~ wire37)  &  wire82 ) ;
 assign wire233 = ( i_40_  &  i_39_  &  n_n985  &  n_n874 ) ;
 assign wire835 = ( (~ i_7_)  &  n_n926  &  wire80 ) | ( (~ i_7_)  &  n_n833  &  wire80 ) ;
 assign wire837 = ( i_39_  &  i_38_ ) | ( i_40_  &  (~ i_38_) ) ;
 assign wire375 = ( (~ i_30_)  &  (~ i_29_) ) ;
 assign wire482 = ( i_24_  &  i_22_  &  n_n968  &  n_n1074 ) ;
 assign wire474 = ( i_24_  &  n_n968  &  n_n1074  &  wire7510 ) ;
 assign wire478 = ( (~ i_12_)  &  i_17_  &  i_15_  &  n_n955 ) ;
 assign wire481 = ( i_16_  &  wire320  &  wire82 ) ;
 assign wire840 = ( (~ i_14_)  &  wire469 ) | ( i_16_  &  wire841 ) ;
 assign wire483 = ( wire840  &  wire7817 ) ;
 assign wire496 = ( n_n977  &  n_n1073  &  wire79 ) ;
 assign wire546 = ( n_n1061  &  wire50 ) | ( n_n582  &  wire80 ) ;
 assign wire548 = ( (~ i_40_)  &  (~ i_38_) ) | ( (~ i_39_)  &  (~ i_38_) ) ;
 assign wire558 = ( n_n933  &  n_n1066 ) | ( n_n1066  &  n_n927 ) ;
 assign wire589 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( (~ i_40_)  &  i_39_  &  n_n1009 ) ;
 assign wire609 = ( i_12_  &  i_18_  &  i_15_ ) | ( i_11_  &  i_18_  &  i_15_ ) ;
 assign wire613 = ( i_40_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) | ( i_40_  &  (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire622 = ( n_n859 ) | ( wire1797 ) | ( wire1798 ) ;
 assign wire636 = ( (~ i_34_)  &  n_n865  &  wire46 ) | ( i_34_  &  n_n1073  &  wire46 ) ;
 assign wire638 = ( i_40_  &  i_39_  &  (~ i_37_) ) | ( i_40_  &  (~ i_38_)  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire642 = ( wire330  &  n_n998 ) | ( n_n979  &  wire60 ) ;
 assign wire652 = ( n_n998  &  n_n866 ) | ( n_n977  &  n_n888 ) ;
 assign wire650 = ( (~ i_5_)  &  i_12_  &  i_15_ ) | ( (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire677 = ( i_3_ ) | ( i_4_ ) | ( i_1_ ) | ( i_2_ ) ;
 assign wire681 = ( i_3_  &  i_0_  &  (~ i_32_) ) | ( i_2_  &  i_0_  &  (~ i_32_) ) ;
 assign wire686 = ( i_12_  &  wire407 ) | ( wire484  &  wire687 ) ;
 assign wire687 = ( i_17_ ) | ( i_16_ ) ;
 assign wire693 = ( (~ i_14_) ) | ( (~ i_11_) ) ;
 assign wire715 = ( n_n976  &  n_n795 ) | ( n_n983  &  wire716 ) ;
 assign wire716 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire721 = ( i_37_  &  n_n1011  &  n_n964 ) | ( (~ i_37_)  &  n_n1072  &  n_n964 ) ;
 assign wire729 = ( n_n927  &  wire7007 ) | ( wire39  &  wire7008 ) ;
 assign wire732 = ( wire1048 ) | ( (~ i_32_)  &  n_n952 ) | ( (~ i_32_)  &  n_n427 ) ;
 assign wire731 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire738 = ( (~ i_14_) ) | ( (~ i_12_) ) | ( (~ i_11_) ) ;
 assign wire743 = ( i_40_  &  i_39_ ) | ( i_40_  &  (~ i_38_) ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire749 = ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) | ( (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire756 = ( wire845 ) | ( wire47  &  wire846 ) | ( wire47  &  wire847 ) ;
 assign wire765 = ( wire43 ) | ( wire1300 ) ;
 assign wire767 = ( i_40_  &  (~ i_39_)  &  (~ i_38_) ) | ( i_40_  &  (~ i_39_)  &  (~ i_37_) ) ;
 assign wire781 = ( wire1400 ) | ( i_11_  &  i_16_  &  i_15_ ) ;
 assign wire785 = ( i_40_  &  i_39_  &  (~ i_37_) ) | ( i_39_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire793 = ( i_13_  &  wire371 ) | ( i_9_  &  n_n833 ) ;
 assign wire792 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire797 = ( wire1563 ) | ( i_40_  &  (~ i_39_)  &  n_n1065 ) ;
 assign wire801 = ( (~ i_37_)  &  wire66  &  n_n964 ) | ( i_37_  &  n_n1011  &  n_n964 ) ;
 assign wire813 = ( n_n933  &  wire63 ) | ( n_n927  &  wire7182 ) ;
 assign wire818 = ( (~ i_9_)  &  (~ i_17_) ) | ( (~ i_9_)  &  (~ i_16_) ) | ( (~ i_17_)  &  (~ i_16_) ) ;
 assign wire820 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_ ) | ( i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire824 = ( n_n969  &  n_n968 ) | ( n_n978  &  wire6907 ) ;
 assign wire828 = ( i_40_  &  i_39_ ) | ( i_39_  &  (~ i_38_) ) ;
 assign wire841 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_)  &  i_11_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  (~ i_11_) ) ;
 assign wire56 = ( n_n785  &  wire463 ) | ( n_n785  &  wire483 ) | ( n_n785  &  wire7820 ) ;
 assign wire74 = ( wire48  &  wire469  &  n_n428  &  n_n427 ) ;
 assign wire129 = ( wire48  &  n_n428  &  n_n427  &  wire706 ) ;
 assign wire133 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_11_ ) ;
 assign wire136 = ( n_n945  &  wire138  &  wire6789 ) | ( n_n945  &  wire141  &  wire6789 ) ;
 assign wire137 = ( n_n945  &  n_n860  &  wire70  &  wire6789 ) ;
 assign wire138 = ( i_11_  &  i_18_  &  i_15_  &  wire7815 ) ;
 assign wire141 = ( i_18_  &  wire35  &  wire492 ) ;
 assign wire142 = ( n_n883  &  n_n861  &  wire7803 ) ;
 assign wire143 = ( n_n979  &  n_n861  &  wire7805 ) ;
 assign wire144 = ( i_31_  &  (~ i_36_)  &  wire45  &  wire7806 ) ;
 assign wire151 = ( wire420  &  n_n1047  &  wire6728 ) ;
 assign wire160 = ( i_31_  &  (~ i_36_)  &  wire45  &  (~ wire37) ) ;
 assign wire162 = ( (~ i_36_)  &  (~ i_35_)  &  i_38_  &  i_37_ ) ;
 assign wire163 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  (~ i_38_) ) ;
 assign wire164 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire165 = ( (~ i_7_)  &  wire50  &  n_n693  &  wire7795 ) ;
 assign wire167 = ( n_n1047  &  wire6728  &  wire7796 ) ;
 assign wire169 = ( n_n982  &  wire88  &  n_n998 ) ;
 assign wire170 = ( wire88  &  n_n997  &  n_n991 ) ;
 assign wire171 = ( n_n469  &  n_n861  &  n_n1002 ) ;
 assign wire188 = ( n_n979  &  n_n330  &  wire602  &  n_n700 ) ;
 assign wire189 = ( n_n978  &  wire196 ) | ( n_n978  &  wire197 ) ;
 assign wire190 = ( wire45  &  n_n462  &  n_n801  &  wire375 ) ;
 assign wire191 = ( n_n977  &  n_n861  &  n_n710  &  n_n715 ) ;
 assign wire192 = ( n_n998  &  n_n799  &  n_n861  &  n_n710 ) ;
 assign wire193 = ( n_n883  &  n_n861  &  n_n1002  &  n_n710 ) ;
 assign wire196 = ( n_n968  &  wire420  &  n_n1074 ) ;
 assign wire197 = ( i_24_  &  wire47  &  n_n968  &  n_n1074 ) ;
 assign wire198 = ( i_13_  &  wire315  &  wire80  &  wire7777 ) ;
 assign wire199 = ( n_n975  &  wire46  &  wire94  &  wire315 ) ;
 assign wire201 = ( n_n1047  &  n_n700  &  wire325  &  wire7276 ) ;
 assign wire203 = ( i_40_  &  wire206 ) | ( i_40_  &  wire207 ) ;
 assign wire205 = ( i_13_  &  wire50  &  wire315  &  wire54 ) ;
 assign wire206 = ( i_13_  &  n_n985  &  wire50  &  wire315 ) ;
 assign wire207 = ( n_n998  &  n_n975  &  n_n861  &  n_n710 ) ;
 assign wire208 = ( n_n973  &  wire79  &  wire7767 ) ;
 assign wire209 = ( n_n998  &  n_n330  &  n_n795  &  n_n700 ) ;
 assign wire210 = ( (~ i_7_)  &  wire50  &  n_n693  &  wire7770 ) ;
 assign wire211 = ( i_31_  &  (~ i_36_)  &  wire45  &  wire7771 ) ;
 assign wire213 = ( (~ i_40_)  &  (~ i_7_)  &  wire50  &  wire6920 ) ;
 assign wire217 = ( (~ i_5_)  &  wire45  &  wire202  &  n_n462 ) ;
 assign wire218 = ( n_n874  &  wire226 ) | ( n_n874  &  n_n884  &  wire589 ) ;
 assign wire226 = ( i_40_  &  (~ i_39_)  &  n_n985  &  wire7760 ) ;
 assign wire229 = ( (~ i_9_)  &  (~ i_5_)  &  n_n997  &  wire45 ) ;
 assign wire231 = ( (~ i_25_)  &  n_n975  &  n_n1002  &  wire46 ) ;
 assign wire232 = ( n_n883  &  n_n1074  &  n_n864 ) ;
 assign wire234 = ( i_1_  &  n_n1055  &  n_n998  &  wire46 ) ;
 assign wire235 = ( n_n978  &  n_n966  &  n_n1012 ) ;
 assign wire243 = ( wire7741  &  wire7743 ) | ( wire7742  &  wire7743 ) ;
 assign wire248 = ( n_n1023  &  n_n458  &  wire403 ) ;
 assign wire249 = ( wire45  &  wire254 ) | ( n_n973  &  wire45  &  wire7745 ) ;
 assign wire250 = ( (~ i_40_)  &  i_39_  &  n_n979  &  wire7227 ) ;
 assign wire252 = ( i_2_  &  n_n1055  &  n_n998  &  wire46 ) ;
 assign wire254 = ( i_30_  &  (~ i_5_)  &  n_n462 ) ;
 assign wire260 = ( n_n1074  &  wire665  &  wire6731 ) ;
 assign wire261 = ( n_n966  &  n_n1073  &  wire666 ) ;
 assign wire262 = ( i_39_  &  n_n1074  &  n_n970 ) ;
 assign wire263 = ( n_n1055  &  n_n998  &  wire46  &  wire135 ) ;
 assign wire264 = ( (~ i_12_)  &  n_n1074  &  wire6739 ) ;
 assign wire271 = ( i_40_  &  (~ i_38_)  &  n_n1074  &  n_n970 ) ;
 assign wire272 = ( (~ i_14_)  &  n_n1074  &  wire6739 ) ;
 assign wire274 = ( (~ i_15_)  &  n_n1074  &  wire6739 ) ;
 assign wire276 = ( n_n926  &  wire45  &  n_n947  &  (~ wire37) ) ;
 assign wire277 = ( i_15_  &  wire283 ) | ( i_15_  &  wire520  &  wire7726 ) ;
 assign wire279 = ( wire445  &  n_n492  &  wire352  &  wire421 ) ;
 assign wire283 = ( n_n488  &  wire284 ) | ( n_n488  &  wire285 ) ;
 assign wire284 = ( (~ i_17_)  &  n_n926  &  wire45 ) ;
 assign wire285 = ( (~ i_16_)  &  wire445  &  wire421 ) ;
 assign wire286 = ( wire45  &  n_n488  &  n_n923  &  wire7717 ) ;
 assign wire287 = ( n_n791  &  wire291 ) | ( n_n791  &  wire652  &  wire650 ) ;
 assign wire288 = ( n_n979  &  n_n969  &  n_n949  &  n_n791 ) ;
 assign wire289 = ( n_n979  &  n_n1001  &  n_n949  &  wire7406 ) ;
 assign wire291 = ( n_n979  &  n_n969  &  n_n947 ) ;
 assign wire294 = ( (~ i_36_)  &  wire45  &  wire627  &  wire7707 ) ;
 assign wire295 = ( n_n947  &  wire400  &  (~ wire37)  &  wire421 ) ;
 assign wire297 = ( wire45  &  wire306 ) | ( wire45  &  wire307 ) | ( wire45  &  wire308 ) ;
 assign wire298 = ( n_n1023  &  n_n1065  &  n_n1057  &  n_n843 ) ;
 assign wire299 = ( (~ i_40_)  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire306 = ( (~ i_9_)  &  (~ i_11_)  &  n_n947  &  n_n923 ) ;
 assign wire307 = ( (~ i_16_)  &  i_15_  &  n_n985  &  n_n488 ) ;
 assign wire308 = ( (~ i_16_)  &  i_15_  &  n_n492  &  n_n918 ) ;
 assign wire309 = ( (~ i_36_)  &  wire45  &  n_n488  &  wire7698 ) ;
 assign wire310 = ( n_n1021  &  n_n862  &  n_n1074  &  wire635 ) ;
 assign wire311 = ( n_n710  &  wire414 ) | ( n_n1008  &  n_n710  &  wire636 ) ;
 assign wire312 = ( n_n1055  &  n_n1047  &  wire39  &  wire7689 ) ;
 assign wire414 = ( i_40_  &  i_39_  &  n_n1074  &  n_n1065 ) ;
 assign wire443 = ( wire633  &  wire447 ) | ( wire633  &  wire449 ) ;
 assign wire444 = ( n_n969  &  n_n162 ) | ( n_n969  &  n_n164 ) ;
 assign wire446 = ( n_n1001  &  n_n460 ) | ( n_n1001  &  n_n162 ) | ( n_n1001  &  n_n459 ) ;
 assign wire447 = ( n_n977  &  n_n888  &  wire7694 ) ;
 assign wire449 = ( (~ i_22_)  &  n_n998  &  n_n866  &  wire46 ) ;
 assign wire451 = ( n_n1021  &  n_n874  &  n_n1009  &  wire7686 ) ;
 assign wire454 = ( n_n979  &  wire81  &  n_n791  &  wire36 ) ;
 assign wire455 = ( n_n1073  &  n_n960  &  wire39  &  wire7689 ) ;
 assign wire459 = ( (~ i_39_)  &  (~ i_38_)  &  n_n460 ) | ( (~ i_39_)  &  (~ i_38_)  &  n_n459 ) ;
 assign wire519 = ( wire87  &  wire50  &  wire7670 ) | ( wire50  &  wire82  &  wire7670 ) ;
 assign wire533 = ( n_n1066  &  n_n462  &  wire494  &  wire7122 ) ;
 assign wire536 = ( (~ i_40_)  &  wire843 ) | ( (~ i_40_)  &  n_n795  &  wire756 ) ;
 assign wire538 = ( n_n883  &  n_n861  &  n_n1002  &  n_n710 ) ;
 assign wire843 = ( n_n861  &  n_n1002  &  n_n710  &  wire100 ) ;
 assign wire845 = ( (~ i_31_)  &  wire45  &  wire43 ) ;
 assign wire846 = ( i_30_  &  (~ i_31_)  &  (~ i_29_)  &  wire45 ) ;
 assign wire847 = ( i_29_  &  n_n1066  &  wire7122 ) ;
 assign wire849 = ( (~ i_36_)  &  (~ i_38_)  &  i_37_  &  wire704 ) ;
 assign wire850 = ( i_13_  &  wire76  &  wire315  &  wire401 ) ;
 assign wire855 = ( i_40_  &  (~ i_13_)  &  wire50  &  wire315 ) ;
 assign wire856 = ( i_40_  &  i_39_  &  (~ i_13_)  &  wire80 ) ;
 assign wire857 = ( i_40_  &  (~ i_39_)  &  (~ i_31_)  &  wire45 ) ;
 assign wire859 = ( wire420  &  n_n1048  &  n_n1047  &  wire697 ) ;
 assign wire860 = ( wire330  &  n_n998  &  n_n700  &  wire7276 ) ;
 assign wire864 = ( n_n998  &  wire441  &  n_n861 ) ;
 assign wire865 = ( (~ i_38_)  &  (~ i_37_)  &  n_n861  &  n_n1002 ) ;
 assign wire869 = ( n_n979  &  wire594  &  n_n700  &  wire7276 ) ;
 assign wire872 = ( i_13_  &  n_n528  &  wire50  &  wire315 ) ;
 assign wire873 = ( n_n977  &  n_n861  &  n_n1002  &  n_n710 ) ;
 assign wire875 = ( i_40_  &  (~ i_39_)  &  n_n330  &  n_n700 ) ;
 assign wire876 = ( n_n969  &  n_n700  &  wire7276 ) ;
 assign wire882 = ( wire888  &  wire7640 ) | ( n_n989  &  n_n1066  &  wire7640 ) ;
 assign wire888 = ( (~ i_12_)  &  (~ i_31_)  &  wire45 ) | ( (~ i_11_)  &  (~ i_31_)  &  wire45 ) ;
 assign wire890 = ( (~ i_7_)  &  wire493  &  wire50  &  wire7627 ) ;
 assign wire891 = ( wire302  &  wire7630 ) | ( wire902  &  wire7630 ) | ( wire1810  &  wire7630 ) ;
 assign wire892 = ( wire402  &  wire7632 ) | ( wire402  &  wire79  &  wire7631 ) ;
 assign wire893 = ( n_n998  &  wire495  &  n_n861 ) ;
 assign wire894 = ( (~ i_7_)  &  i_2_  &  n_n926  &  wire80 ) ;
 assign wire902 = ( (~ i_1_)  &  i_0_  &  wire79 ) ;
 assign wire904 = ( i_40_  &  n_n861  &  n_n991  &  wire740 ) ;
 assign wire905 = ( n_n1056  &  wire325  &  wire7620 ) ;
 assign wire906 = ( n_n982  &  wire88  &  n_n998 ) ;
 assign wire911 = ( n_n975  &  n_n700  &  wire94  &  wire7276 ) ;
 assign wire912 = ( n_n976  &  wire920 ) | ( n_n976  &  wire921 ) ;
 assign wire913 = ( n_n469  &  wire922 ) | ( n_n469  &  wire7610 ) ;
 assign wire920 = ( n_n330  &  n_n989  &  wire445 ) ;
 assign wire921 = ( (~ i_32_)  &  (~ i_31_)  &  wire315  &  wire325 ) ;
 assign wire922 = ( n_n1048  &  n_n1047  &  n_n527 ) ;
 assign wire925 = ( n_n973  &  wire420  &  n_n1048  &  n_n1073 ) ;
 assign wire926 = ( wire402  &  n_n1074  &  wire6897 ) | ( n_n1074  &  wire930  &  wire6897 ) ;
 assign wire927 = ( (~ i_40_)  &  i_39_  &  wire398 ) | ( (~ i_40_)  &  i_39_  &  wire932 ) ;
 assign wire928 = ( n_n971  &  wire346  &  wire79  &  (~ wire115) ) ;
 assign wire929 = ( (~ i_7_)  &  i_2_  &  n_n833  &  wire80 ) ;
 assign wire930 = ( (~ i_40_)  &  i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire932 = ( n_n1048  &  wire934  &  wire7602 ) | ( n_n1048  &  wire7601  &  wire7602 ) ;
 assign wire934 = ( i_30_  &  (~ i_7_)  &  (~ i_5_) ) ;
 assign wire937 = ( n_n1066  &  n_n462  &  wire7122  &  wire7593 ) ;
 assign wire939 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  wire744 ) ;
 assign wire940 = ( n_n998  &  n_n861  &  n_n710  &  wire124 ) ;
 assign wire942 = ( wire84  &  n_n853  &  wire7586 ) | ( n_n853  &  wire948  &  wire7586 ) ;
 assign wire948 = ( n_n1072  &  n_n1048  &  n_n1073 ) ;
 assign wire950 = ( n_n1055  &  n_n979  &  n_n783 ) | ( n_n1055  &  n_n979  &  n_n790 ) ;
 assign wire952 = ( n_n1055  &  n_n1047  &  n_n777 ) | ( n_n1055  &  n_n1047  &  n_n771 ) ;
 assign wire957 = ( wire68  &  wire504 ) ;
 assign wire962 = ( n_n833  &  n_n764 ) | ( n_n764  &  wire967 ) | ( n_n833  &  wire7572 ) | ( wire967  &  wire7572 ) ;
 assign wire964 = ( (~ i_22_)  &  n_n926  &  wire50  &  wire82 ) ;
 assign wire967 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire973 = ( wire441  &  n_n861  &  n_n1002  &  n_n710 ) ;
 assign wire983 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire985 = ( n_n799  &  n_n861  &  wire624 ) ;
 assign wire986 = ( (~ i_7_)  &  wire50  &  wire623  &  n_n693 ) ;
 assign wire987 = ( (~ i_38_)  &  i_37_  &  n_n979  &  wire88 ) ;
 assign wire988 = ( n_n990  &  n_n861  &  n_n1002 ) ;
 assign wire999 = ( n_n1072  &  wire380  &  wire482 ) | ( n_n1072  &  wire482  &  wire7127 ) ;
 assign wire1000 = ( n_n978  &  n_n937  &  wire6907 ) ;
 assign wire1008 = ( n_n883  &  n_n1074  &  n_n864 ) ;
 assign wire1010 = ( n_n973  &  n_n966  &  n_n1073 ) ;
 assign wire1019 = ( wire512  &  wire7521 ) ;
 assign wire1020 = ( wire1842  &  wire7522 ) | ( wire48  &  n_n951  &  wire7522 ) ;
 assign wire1021 = ( wire416  &  wire579 ) ;
 assign wire1022 = ( wire84  &  wire478 ) | ( wire84  &  wire1029 ) ;
 assign wire1029 = ( i_12_  &  i_17_  &  i_15_  &  n_n928 ) ;
 assign wire1031 = ( i_20_  &  i_21_  &  wire1038 ) | ( i_20_  &  i_21_  &  wire1039 ) ;
 assign wire1038 = ( n_n952  &  wire7514 ) | ( n_n427  &  wire7514 ) | ( wire1040  &  wire7514 ) ;
 assign wire1039 = ( i_15_  &  wire35  &  n_n411  &  wire303 ) ;
 assign wire1040 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052  &  n_n1023 ) ;
 assign wire1043 = ( wire1046  &  wire7511 ) | ( wire732  &  wire7509  &  wire7511 ) ;
 assign wire1044 = ( i_20_  &  wire35  &  n_n848  &  wire7512 ) ;
 assign wire1046 = ( (~ i_7_)  &  (~ i_5_)  &  i_12_  &  wire474 ) ;
 assign wire1048 = ( (~ i_40_)  &  (~ i_39_)  &  n_n1052  &  wire50 ) ;
 assign wire1049 = ( n_n980  &  wire574  &  n_n1047  &  wire7500 ) ;
 assign wire1050 = ( (~ i_15_)  &  wire1058 ) | ( (~ i_15_)  &  wire1059 ) ;
 assign wire1051 = ( i_38_  &  n_n685  &  n_n865  &  n_n1074 ) ;
 assign wire1058 = ( (~ i_7_)  &  n_n1008  &  wire45  &  n_n1009 ) ;
 assign wire1059 = ( (~ i_7_)  &  n_n1008  &  n_n1052  &  wire50 ) ;
 assign wire1060 = ( n_n469  &  n_n983  &  n_n668 ) ;
 assign wire1061 = ( (~ i_40_)  &  wire392 ) | ( (~ i_40_)  &  wire1065 ) ;
 assign wire1062 = ( (~ i_15_)  &  wire1067 ) | ( (~ i_15_)  &  wire79  &  wire793 ) ;
 assign wire1063 = ( (~ i_39_)  &  n_n685  &  n_n874  &  n_n1052 ) ;
 assign wire1065 = ( n_n685  &  n_n1074  &  n_n923 ) ;
 assign wire1067 = ( (~ i_7_)  &  wire45  &  wire792 ) ;
 assign wire1073 = ( i_9_  &  (~ i_11_)  &  wire496 ) | ( i_9_  &  (~ i_11_)  &  wire1078 ) ;
 assign wire1075 = ( n_n685  &  n_n971  &  n_n1072  &  n_n1074 ) ;
 assign wire1078 = ( (~ i_7_)  &  n_n1001  &  n_n1047  &  wire38 ) ;
 assign wire1083 = ( (~ i_12_)  &  wire1084 ) | ( (~ i_12_)  &  wire1085 ) ;
 assign wire1084 = ( n_n1001  &  n_n1047  &  wire344  &  wire38 ) ;
 assign wire1085 = ( i_9_  &  n_n977  &  n_n1073  &  wire79 ) ;
 assign wire1088 = ( n_n980  &  n_n1001  &  wire674  &  wire7479 ) ;
 assign wire1089 = ( n_n1055  &  n_n1047  &  wire351  &  wire7482 ) ;
 assign wire1090 = ( n_n969  &  n_n968  &  n_n1074  &  n_n629 ) ;
 assign wire1091 = ( n_n685  &  n_n1064  &  n_n1074  &  n_n1065 ) ;
 assign wire1092 = ( n_n1073  &  n_n967  &  n_n1074  &  n_n629 ) ;
 assign wire1093 = ( (~ i_7_)  &  n_n1047  &  wire717  &  wire6728 ) ;
 assign wire1099 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire1104 = ( n_n1066  &  n_n668  &  wire713 ) ;
 assign wire1106 = ( i_40_  &  wire1109 ) | ( i_40_  &  wire376  &  wire715 ) ;
 assign wire1107 = ( (~ i_7_)  &  n_n833  &  wire50 ) ;
 assign wire1109 = ( (~ i_7_)  &  wire45  &  n_n836 ) ;
 assign wire1112 = ( wire363  &  n_n629 ) | ( n_n629  &  wire303 ) | ( n_n629  &  wire233 ) ;
 assign wire1113 = ( wire390  &  wire1114 ) | ( wire390  &  wire7466 ) | ( wire390  &  wire7467 ) ;
 assign wire1114 = ( (~ i_36_)  &  wire1119 ) | ( (~ i_36_)  &  wire1120 ) ;
 assign wire1119 = ( i_40_  &  (~ i_39_)  &  i_13_  &  (~ i_38_) ) ;
 assign wire1120 = ( i_9_  &  i_39_  &  i_38_  &  (~ i_37_) ) ;
 assign wire1122 = ( n_n969  &  n_n968  &  n_n819 ) ;
 assign wire1132 = ( wire87  &  wire475 ) | ( wire87  &  wire476  &  wire824 ) ;
 assign wire1139 = ( i_4_  &  n_n1055  &  n_n998  &  wire46 ) ;
 assign wire1155 = ( wire50  &  wire403  &  wire7435 ) ;
 assign wire1156 = ( n_n1055  &  n_n998  &  wire46  &  wire675 ) ;
 assign wire1158 = ( n_n865  &  n_n799  &  n_n1074 ) ;
 assign wire1160 = ( (~ i_39_)  &  i_2_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire1163 = ( n_n949  &  wire1168 ) | ( n_n949  &  wire1169 ) ;
 assign wire1164 = ( n_n979  &  n_n469  &  n_n949  &  wire7347 ) ;
 assign wire1165 = ( n_n979  &  n_n949  &  wire60  &  wire7406 ) ;
 assign wire1168 = ( wire330  &  n_n998  &  n_n791 ) ;
 assign wire1169 = ( (~ i_22_)  &  wire330  &  n_n998  &  wire46 ) ;
 assign wire1173 = ( (~ i_17_)  &  (~ i_16_)  &  n_n949  &  wire76 ) ;
 assign wire1174 = ( (~ i_17_)  &  i_15_  &  n_n492  &  wire76 ) ;
 assign wire1179 = ( wire611  &  wire7415 ) ;
 assign wire1181 = ( n_n985  &  wire467  &  wire7121 ) | ( n_n985  &  wire468  &  wire7121 ) ;
 assign wire1182 = ( n_n979  &  n_n949  &  wire60  &  n_n791 ) ;
 assign wire1183 = ( n_n484  &  wire401 ) | ( n_n484  &  wire465 ) ;
 assign wire1186 = ( n_n979  &  n_n949  &  wire615  &  wire7405 ) ;
 assign wire1189 = ( n_n979  &  n_n975  &  n_n947  &  wire7399 ) ;
 assign wire1192 = ( n_n979  &  n_n947  &  n_n791 ) ;
 assign wire1196 = ( wire69  &  wire7398 ) | ( n_n1066  &  n_n458  &  wire7398 ) ;
 assign wire1197 = ( n_n979  &  n_n947  &  wire660  &  wire7399 ) ;
 assign wire1198 = ( n_n1057  &  n_n843  &  n_n1053  &  n_n836 ) ;
 assign wire1199 = ( n_n1023  &  n_n1065  &  n_n1057  &  n_n843 ) ;
 assign wire1200 = ( n_n1064  &  n_n1066  &  n_n1065  &  n_n458 ) ;
 assign wire1204 = ( n_n1052  &  n_n1057  &  n_n1053  &  wire7388 ) ;
 assign wire1205 = ( n_n947  &  wire1210 ) | ( n_n947  &  n_n791  &  wire642 ) ;
 assign wire1206 = ( n_n979  &  n_n469  &  n_n947  &  wire7347 ) ;
 assign wire1208 = ( n_n979  &  n_n947  &  wire60  &  wire7390 ) ;
 assign wire1210 = ( (~ i_22_)  &  wire330  &  n_n998  &  wire46 ) ;
 assign wire1213 = ( n_n865  &  wire373  &  wire1219 ) | ( n_n865  &  wire373  &  wire7372 ) ;
 assign wire1219 = ( (~ i_4_)  &  i_0_  &  wire79 ) | ( (~ i_1_)  &  i_0_  &  wire79 ) ;
 assign wire1222 = ( n_n842  &  n_n993  &  n_n843  &  wire7360 ) ;
 assign wire1230 = ( (~ i_24_)  &  wire371  &  wire50  &  wire82 ) ;
 assign wire1238 = ( (~ i_39_)  &  i_38_  &  n_n998  &  n_n861 ) ;
 assign wire1246 = ( n_n979  &  n_n861  &  n_n795 ) ;
 assign wire1247 = ( n_n977  &  n_n861  &  n_n991 ) ;
 assign wire1251 = ( (~ i_40_)  &  (~ i_10_)  &  i_38_ ) | ( (~ i_40_)  &  (~ i_27_)  &  i_38_ ) ;
 assign wire1252 = ( i_40_  &  (~ i_11_)  &  (~ i_38_) ) ;
 assign wire1253 = ( n_n998  &  n_n861  &  wire7332 ) ;
 assign wire1254 = ( n_n861  &  wire7334 ) | ( n_n969  &  n_n971  &  n_n861 ) ;
 assign wire1255 = ( i_38_  &  i_37_  &  n_n861  &  wire94 ) ;
 assign wire1256 = ( (~ i_38_)  &  i_37_  &  n_n979  &  wire88 ) ;
 assign wire1257 = ( n_n979  &  n_n1005  &  n_n861 ) ;
 assign wire1262 = ( n_n883  &  n_n888  &  n_n861 ) ;
 assign wire1264 = ( n_n535  &  wire7324 ) | ( wire481  &  wire7324 ) | ( wire7323  &  wire7324 ) ;
 assign wire1265 = ( wire481  &  wire7325 ) | ( wire7323  &  wire7325 ) ;
 assign wire1269 = ( i_40_  &  (~ i_39_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire1271 = ( n_n862  &  n_n860  &  (~ wire166)  &  wire7314 ) ;
 assign wire1277 = ( i_17_  &  wire721  &  wire7308 ) | ( i_16_  &  wire721  &  wire7308 ) ;
 assign wire1284 = ( n_n528  &  n_n525 ) | ( n_n528  &  wire1289 ) ;
 assign wire1285 = ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_)  &  wire723 ) ;
 assign wire1286 = ( n_n998  &  n_n799  &  n_n861  &  n_n710 ) ;
 assign wire1289 = ( i_24_  &  i_15_  &  wire35  &  wire50 ) ;
 assign wire1291 = ( i_30_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire1294 = ( (~ i_7_)  &  wire471  &  wire80  &  wire763 ) ;
 assign wire1295 = ( (~ i_40_)  &  wire1299 ) | ( (~ i_40_)  &  wire765  &  wire7291 ) ;
 assign wire1299 = ( i_16_  &  wire87  &  wire320  &  n_n688 ) ;
 assign wire1300 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_5_)  &  i_29_ ) | ( i_30_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire1305 = ( (~ i_7_)  &  wire471  &  wire80  &  wire7275 ) ;
 assign wire1306 = ( n_n888  &  n_n1064  &  n_n700  &  wire7276 ) ;
 assign wire1307 = ( n_n998  &  n_n861  &  n_n710  &  wire7278 ) ;
 assign wire1309 = ( i_38_  &  n_n861  &  n_n710  &  n_n715 ) ;
 assign wire1311 = ( n_n1047  &  wire494  &  wire7279 ) ;
 assign wire1312 = ( i_39_  &  i_38_  &  n_n1012  &  wire7281 ) ;
 assign wire1316 = ( (~ i_40_)  &  n_n966  &  n_n862 ) | ( (~ i_39_)  &  n_n966  &  n_n862 ) ;
 assign wire1317 = ( n_n874  &  n_n462 ) | ( n_n874  &  wire1326 ) ;
 assign wire1326 = ( i_40_  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire1328 = ( (~ i_36_)  &  wire45  &  wire7253 ) ;
 assign wire1329 = ( (~ i_12_)  &  (~ i_11_)  &  wire45  &  n_n918 ) ;
 assign wire1330 = ( (~ i_38_)  &  (~ i_37_)  &  n_n1006  &  n_n976 ) ;
 assign wire1340 = ( (~ i_40_)  &  (~ i_38_)  &  n_n715  &  wire7246 ) ;
 assign wire1341 = ( n_n998  &  wire81  &  wire46  &  wire808 ) ;
 assign wire1342 = ( n_n966  &  n_n1012  &  wire807 ) ;
 assign wire1343 = ( i_35_  &  (~ i_37_)  &  n_n977  &  n_n1074 ) ;
 assign wire1344 = ( (~ i_40_)  &  i_39_  &  n_n698  &  n_n1074 ) ;
 assign wire1346 = ( (~ i_12_)  &  n_n1073  &  wire7239 ) | ( (~ i_11_)  &  n_n1073  &  wire7239 ) ;
 assign wire1347 = ( (~ i_39_)  &  i_38_  &  n_n971  &  n_n1074 ) ;
 assign wire1348 = ( i_39_  &  (~ i_38_)  &  n_n1047  &  n_n700 ) ;
 assign wire1349 = ( wire806  &  wire805 ) ;
 assign wire1353 = ( i_5_  &  (~ i_0_)  &  (~ i_32_)  &  wire7231 ) ;
 assign wire1354 = ( (~ i_40_)  &  (~ i_39_)  &  n_n874  &  n_n693 ) ;
 assign wire1356 = ( i_38_  &  wire1362 ) | ( i_38_  &  wire7234 ) ;
 assign wire1357 = ( i_39_  &  n_n1074  &  n_n970 ) ;
 assign wire1358 = ( (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire1362 = ( i_0_  &  (~ i_32_)  &  i_33_  &  n_n991 ) ;
 assign wire1364 = ( (~ i_32_)  &  (~ i_34_)  &  i_33_  &  wire748 ) ;
 assign wire1365 = ( (~ i_38_)  &  n_n1074  &  n_n864 ) ;
 assign wire1366 = ( i_40_  &  n_n1074  &  wire6731 ) | ( (~ i_39_)  &  n_n1074  &  wire6731 ) ;
 assign wire1367 = ( i_38_  &  n_n966  &  n_n1073 ) ;
 assign wire1371 = ( (~ i_31_)  &  n_n1047  &  wire7191  &  wire7214 ) ;
 assign wire1372 = ( i_32_  &  n_n1047  &  wire7191 ) | ( n_n1047  &  wire1381  &  wire7191 ) ;
 assign wire1374 = ( n_n685  &  (~ n_n1014)  &  n_n874  &  n_n1052 ) ;
 assign wire1375 = ( i_38_  &  n_n685  &  n_n865  &  n_n1074 ) ;
 assign wire1381 = ( (~ i_9_)  &  i_5_  &  (~ i_17_) ) | ( (~ i_9_)  &  i_5_  &  (~ i_16_) ) ;
 assign wire1383 = ( wire320  &  wire383  &  (~ wire166)  &  wire7205 ) ;
 assign wire1386 = ( n_n685  &  n_n971  &  n_n1072  &  n_n1074 ) ;
 assign wire1388 = ( i_11_  &  i_16_  &  i_15_ ) ;
 assign wire1389 = ( i_9_  &  i_12_  &  i_15_ ) ;
 assign wire1390 = ( i_37_  &  n_n685  &  n_n1074  &  wire779 ) ;
 assign wire1400 = ( i_9_  &  i_12_  &  i_15_ ) ;
 assign wire1402 = ( n_n1066  &  wire166  &  wire7197 ) ;
 assign wire1412 = ( (~ i_39_)  &  i_38_  &  n_n966  &  n_n1073 ) ;
 assign wire1415 = ( n_n998  &  wire46  &  wire471  &  wire7181 ) ;
 assign wire1416 = ( n_n923  &  wire1423 ) | ( n_n1066  &  n_n923  &  wire813 ) ;
 assign wire1417 = ( n_n979  &  wire342  &  n_n907  &  wire6716 ) ;
 assign wire1423 = ( n_n1066  &  n_n928  &  n_n927 ) ;
 assign wire1428 = ( n_n880  &  n_n1048  &  n_n1047  &  n_n907 ) ;
 assign wire1429 = ( wire76  &  wire1435 ) | ( wire378  &  wire76  &  wire801 ) ;
 assign wire1430 = ( n_n857  &  n_n884 ) | ( n_n884  &  wire303 ) | ( n_n884  &  wire1438 ) ;
 assign wire1435 = ( i_39_  &  i_38_  &  wire317  &  n_n1012 ) ;
 assign wire1438 = ( i_35_  &  (~ i_37_)  &  n_n969  &  n_n1074 ) ;
 assign wire1441 = ( n_n1008  &  wire422  &  n_n1009  &  wire378 ) ;
 assign wire1442 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire7164 ) ;
 assign wire1443 = ( i_40_  &  wire1447 ) | ( i_40_  &  wire1448 ) | ( i_40_  &  wire1449 ) ;
 assign wire1444 = ( n_n1014  &  n_n966  &  n_n993  &  n_n884 ) ;
 assign wire1447 = ( (~ i_32_)  &  i_33_  &  n_n991  &  wire7165 ) ;
 assign wire1448 = ( (~ i_5_)  &  (~ i_15_)  &  n_n993  &  wire76 ) ;
 assign wire1449 = ( i_6_  &  wire1450 ) | ( i_6_  &  wire1451 ) ;
 assign wire1450 = ( i_38_  &  (~ i_37_)  &  n_n1002  &  wire46 ) ;
 assign wire1451 = ( (~ i_32_)  &  i_33_  &  n_n998  &  wire100 ) ;
 assign wire1452 = ( n_n973  &  wire7157 ) | ( n_n973  &  n_n865  &  n_n1074 ) ;
 assign wire1453 = ( (~ i_40_)  &  i_39_  &  n_n1074  &  n_n1061 ) ;
 assign wire1454 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1074  &  n_n864 ) ;
 assign wire1455 = ( n_n969  &  n_n1074  &  n_n970 ) ;
 assign wire1459 = ( n_n1023  &  n_n1057  &  wire7063  &  wire7148 ) ;
 assign wire1466 = ( n_n1067  &  wire518 ) | ( n_n1067  &  wire393 ) ;
 assign wire1467 = ( n_n907  &  wire1472 ) | ( n_n907  &  wire7142 ) ;
 assign wire1468 = ( n_n979  &  n_n1001  &  n_n907  &  wire6716 ) ;
 assign wire1472 = ( n_n1048  &  n_n1073  &  n_n967 ) ;
 assign wire1475 = ( n_n926  &  wire1483 ) | ( n_n926  &  wire1484 ) ;
 assign wire1483 = ( n_n933  &  n_n1066  &  n_n928 ) ;
 assign wire1484 = ( n_n1066  &  n_n927  &  wire63 ) ;
 assign wire1487 = ( i_40_  &  i_39_  &  (~ i_36_)  &  i_38_ ) ;
 assign wire1489 = ( n_n1014  &  wire380  &  wire482 ) | ( n_n1014  &  wire482  &  wire7127 ) ;
 assign wire1496 = ( n_n971  &  n_n880  &  n_n1074  &  n_n629 ) ;
 assign wire1499 = ( wire88  &  n_n998  &  n_n997 ) ;
 assign wire1501 = ( n_n975  &  n_n861  &  n_n991 ) ;
 assign wire1505 = ( wire7103  &  wire7105 ) | ( wire7104  &  wire7105 ) ;
 assign wire1506 = ( (~ i_7_)  &  wire1509 ) | ( (~ i_7_)  &  wire1510 ) ;
 assign wire1509 = ( (~ i_6_)  &  i_34_  &  n_n1072  &  n_n1012 ) ;
 assign wire1510 = ( i_32_  &  wire7109 ) | ( i_32_  &  n_n693  &  wire7108 ) ;
 assign wire1518 = ( n_n1072  &  n_n864  &  wire7097 ) ;
 assign wire1520 = ( (~ i_7_)  &  (~ i_5_)  &  wire400  &  n_n991 ) ;
 assign wire1521 = ( (~ i_7_)  &  (~ i_34_)  &  n_n969  &  n_n865 ) ;
 assign wire1522 = ( n_n989  &  n_n983  &  wire445 ) ;
 assign wire1524 = ( n_n1006  &  wire7089 ) | ( n_n1006  &  wire7090 ) ;
 assign wire1525 = ( n_n926  &  n_n989  &  n_n1066 ) ;
 assign wire1539 = ( i_9_  &  (~ i_15_)  &  wire76  &  wire465 ) ;
 assign wire1540 = ( n_n1006  &  wire441  &  n_n1056 ) ;
 assign wire1541 = ( (~ i_12_)  &  (~ i_11_)  &  wire76  &  wire401 ) ;
 assign wire1542 = ( n_n989  &  n_n1066  &  wire1546 ) | ( n_n989  &  n_n1066  &  wire1547 ) ;
 assign wire1544 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire820 ) ;
 assign wire1545 = ( (~ i_32_)  &  i_33_  &  n_n998  &  n_n997 ) ;
 assign wire1546 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire1547 = ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire1548 = ( n_n989  &  n_n1066  &  wire7073 ) ;
 assign wire1550 = ( n_n969  &  n_n1074  &  n_n970 ) ;
 assign wire1551 = ( n_n966  &  n_n967  &  n_n1012 ) ;
 assign wire1552 = ( n_n968  &  n_n1074  &  wire59 ) ;
 assign wire1555 = ( n_n1057  &  n_n1056  &  wire7063  &  wire7064 ) ;
 assign wire1557 = ( n_n1067  &  wire1562 ) | ( n_n1067  &  wire797  &  wire7067 ) ;
 assign wire1562 = ( (~ n_n1014)  &  n_n1052  &  n_n1057  &  n_n1053 ) ;
 assign wire1563 = ( i_39_  &  i_36_  &  i_38_  &  (~ i_37_) ) ;
 assign wire1565 = ( i_9_  &  n_n977  &  wire76  &  wire7055 ) ;
 assign wire1566 = ( n_n1055  &  n_n1048  &  n_n1047  &  wire7057 ) ;
 assign wire1568 = ( n_n1067  &  n_n1023  &  n_n1065  &  n_n1057 ) ;
 assign wire1570 = ( i_17_  &  i_16_  &  n_n1072  &  n_n1073 ) ;
 assign wire1571 = ( (~ i_36_)  &  (~ i_35_)  &  (~ i_37_)  &  wire828 ) ;
 assign wire1575 = ( i_17_  &  wire1577 ) | ( i_16_  &  wire1577 ) | ( i_17_  &  wire1578 ) | ( i_16_  &  wire1578 ) ;
 assign wire1577 = ( n_n1055  &  n_n1048  &  n_n1047  &  wire7052 ) ;
 assign wire1578 = ( i_9_  &  n_n1072  &  n_n1073  &  wire76 ) ;
 assign wire1579 = ( (~ i_12_)  &  i_16_ ) | ( (~ i_11_)  &  i_16_ ) ;
 assign wire1583 = ( i_5_  &  (~ i_36_)  &  wire45  &  wire795 ) ;
 assign wire1584 = ( n_n980  &  n_n1047  &  wire794 ) ;
 assign wire1588 = ( i_13_  &  n_n975  &  n_n1002  &  wire46 ) ;
 assign wire1592 = ( (~ i_22_)  &  wire559  &  wire87  &  wire50 ) ;
 assign wire1610 = ( wire68  &  wire504 ) ;
 assign wire1617 = ( (~ i_12_)  &  wire92  &  wire319  &  wire82 ) ;
 assign wire1619 = ( n_n926  &  wire7018 ) | ( n_n926  &  wire319  &  wire470 ) ;
 assign wire1620 = ( wire422  &  n_n462  &  n_n801  &  wire375 ) ;
 assign wire1624 = ( n_n933  &  n_n1066  &  n_n527  &  wire7016 ) ;
 assign wire1626 = ( wire48  &  n_n428  &  n_n427  &  wire727 ) ;
 assign wire1630 = ( n_n1066  &  n_n860  &  wire729 ) ;
 assign wire1632 = ( n_n1066  &  n_n860  &  n_n927  &  wire7011 ) ;
 assign wire1635 = ( wire555  &  wire6999 ) | ( wire555  &  n_n971  &  n_n1072 ) ;
 assign wire1650 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire100 ) ;
 assign wire1651 = ( (~ i_38_)  &  (~ i_37_)  &  n_n998  &  wire46 ) ;
 assign wire1653 = ( wire1657  &  wire6979 ) | ( wire6978  &  wire6979 ) ;
 assign wire1655 = ( n_n1047  &  wire400  &  wire831 ) ;
 assign wire1657 = ( (~ i_18_)  &  wire87 ) | ( (~ i_18_)  &  wire82 ) ;
 assign wire1661 = ( n_n777  &  wire64 ) | ( wire64  &  n_n771 ) ;
 assign wire1662 = ( (~ i_21_)  &  i_15_  &  n_n853  &  wire348 ) ;
 assign wire1666 = ( (~ i_24_)  &  n_n833  &  wire87  &  wire50 ) ;
 assign wire1681 = ( (~ i_24_)  &  wire87  &  wire50  &  wire6945 ) ;
 assign wire1682 = ( (~ i_24_)  &  wire371  &  wire50  &  wire82 ) ;
 assign wire1693 = ( wire48  &  wire35  &  wire1700 ) | ( wire48  &  wire35  &  wire1701 ) ;
 assign wire1700 = ( n_n966  &  n_n1012  &  wire6930 ) ;
 assign wire1701 = ( n_n945  &  wire304  &  wire6789 ) ;
 assign wire1704 = ( n_n998  &  n_n973  &  n_n158  &  wire35 ) ;
 assign wire1705 = ( n_n330  &  n_n969  &  n_n968  &  n_n1074 ) ;
 assign wire1706 = ( n_n865  &  wire429  &  wire373 ) | ( n_n865  &  wire373  &  wire1715 ) ;
 assign wire1707 = ( n_n979  &  n_n978  &  n_n330  &  n_n700 ) ;
 assign wire1708 = ( n_n883  &  n_n998  &  n_n861 ) ;
 assign wire1709 = ( (~ i_7_)  &  n_n1021  &  wire50  &  wire6920 ) ;
 assign wire1715 = ( (~ i_1_)  &  i_0_  &  wire79 ) ;
 assign wire1730 = ( (~ i_7_)  &  n_n1065  &  wire50  &  wire464 ) ;
 assign wire1731 = ( n_n469  &  wire420  &  n_n1048  &  n_n1047 ) ;
 assign wire1741 = ( n_n330  &  n_n989  &  n_n1066  &  wire6890 ) ;
 assign wire1742 = ( n_n979  &  n_n330  &  n_n700  &  wire65 ) ;
 assign wire1747 = ( n_n971  &  n_n1072  &  n_n1074  &  wire6828 ) ;
 assign wire1749 = ( n_n883  &  n_n1074  &  n_n970  &  wire6828 ) ;
 assign wire1751 = ( n_n979  &  n_n158  &  wire702  &  wire701 ) ;
 assign wire1758 = ( n_n330  &  n_n989  &  n_n1066  &  wire6874 ) ;
 assign wire1766 = ( (~ i_40_)  &  i_38_  &  n_n1073  &  n_n334 ) ;
 assign wire1780 = ( wire512  &  wire614  &  wire6842 ) ;
 assign wire1786 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  i_12_ ) ;
 assign wire1789 = ( wire512  &  n_n793  &  wire349  &  wire607 ) ;
 assign wire1791 = ( n_n793  &  n_n952  &  wire6837  &  wire6839 ) ;
 assign wire1792 = ( wire70  &  wire6841 ) | ( wire1793  &  wire6841 ) ;
 assign wire1793 = ( i_11_  &  i_18_  &  (~ i_21_)  &  i_15_ ) ;
 assign wire1795 = ( i_12_  &  (~ i_21_)  &  i_15_  &  i_19_ ) ;
 assign wire1797 = ( i_11_  &  i_15_  &  i_19_ ) ;
 assign wire1798 = ( i_12_  &  i_18_  &  i_15_ ) ;
 assign wire1803 = ( n_n864  &  wire79  &  wire6824 ) ;
 assign wire1804 = ( n_n330  &  n_n1014  &  n_n966  &  n_n993 ) ;
 assign wire1805 = ( n_n865  &  wire373  &  wire302 ) | ( n_n865  &  wire373  &  wire1810 ) ;
 assign wire1806 = ( n_n861  &  n_n1002  &  n_n710  &  wire100 ) ;
 assign wire1807 = ( n_n709  &  n_n998  &  n_n861  &  n_n710 ) ;
 assign wire1810 = ( (~ i_4_)  &  i_0_  &  wire79 ) ;
 assign wire1812 = ( wire88  &  n_n997  &  n_n991 ) ;
 assign wire1821 = ( wire1842  &  wire6800 ) | ( wire48  &  n_n951  &  wire6800 ) ;
 assign wire1822 = ( wire549  &  n_n1074  &  n_n970 ) ;
 assign wire1823 = ( wire48  &  wire1832 ) | ( wire48  &  wire57  &  wire6801 ) ;
 assign wire1832 = ( n_n1072  &  n_n945  &  wire42  &  wire6789 ) ;
 assign wire1834 = ( i_9_  &  (~ i_5_)  &  i_11_  &  i_19_ ) ;
 assign wire1835 = ( wire84  &  wire1838 ) | ( wire84  &  wire1839 ) ;
 assign wire1836 = ( i_12_  &  i_15_  &  wire416  &  n_n928 ) ;
 assign wire1838 = ( i_12_  &  i_17_  &  i_15_  &  n_n928 ) ;
 assign wire1839 = ( i_17_  &  n_n955  &  wire6751 ) | ( i_16_  &  n_n955  &  wire6751 ) ;
 assign wire1842 = ( i_18_  &  (~ i_21_)  &  wire36 ) ;
 assign wire1844 = ( i_18_  &  wire36  &  wire6791 ) ;
 assign wire1845 = ( (~ wire202)  &  n_n1048  &  n_n1047  &  wire458 ) ;
 assign wire1846 = ( n_n528  &  n_n905 ) | ( n_n528  &  wire1850 ) ;
 assign wire1847 = ( n_n998  &  wire46  &  wire471  &  wire342 ) ;
 assign wire1850 = ( n_n979  &  n_n945  &  n_n949 ) | ( n_n979  &  n_n945  &  n_n947 ) ;
 assign wire1852 = ( n_n799  &  n_n1012  &  wire668  &  wire6780 ) ;
 assign wire1853 = ( n_n1048  &  n_n1047  &  wire458  &  wire669 ) ;
 assign wire1854 = ( n_n968  &  n_n1064  &  n_n1074  &  n_n884 ) ;
 assign wire1855 = ( n_n998  &  n_n1001  &  wire46  &  wire471 ) ;
 assign wire1860 = ( n_n975  &  n_n1002  &  wire46  &  wire667 ) ;
 assign wire1861 = ( n_n966  &  n_n799  &  n_n1012 ) ;
 assign wire1862 = ( wire120  &  n_n1074  &  wire6731 ) ;
 assign wire1863 = ( n_n966  &  n_n1073  &  n_n967 ) ;
 assign wire1867 = ( n_n842  &  n_n1067  &  wire335 ) | ( n_n842  &  n_n1067  &  wire1878 ) ;
 assign wire1868 = ( n_n979  &  n_n982  &  wire88 ) ;
 assign wire1870 = ( i_6_  &  wire1875 ) | ( i_6_  &  wire546  &  wire6765 ) ;
 assign wire1871 = ( n_n990  &  n_n861  &  wire94 ) ;
 assign wire1872 = ( n_n1055  &  wire88  &  n_n991 ) ;
 assign wire1875 = ( (~ i_7_)  &  wire50  &  wire6766 ) ;
 assign wire1878 = ( n_n966  &  n_n1073  &  wire548 ) ;
 assign wire1880 = ( wire537  &  wire6749 ) ;
 assign wire1881 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire6750 ) ;
 assign wire1882 = ( wire543  &  n_n1074  &  n_n864 ) ;
 assign wire1883 = ( wire363  &  wire478 ) | ( wire363  &  wire1890 ) | ( wire363  &  wire1891 ) ;
 assign wire1884 = ( wire66  &  n_n1074  &  wire6731 ) ;
 assign wire1890 = ( i_12_  &  i_15_  &  n_n928  &  wire37 ) ;
 assign wire1891 = ( (~ i_12_)  &  i_16_  &  i_15_  &  n_n955 ) ;
 assign wire1896 = ( n_n979  &  n_n866  &  n_n907  &  wire6716 ) ;
 assign wire1901 = ( n_n1073  &  n_n1074  &  wire743 ) ;
 assign wire1902 = ( (~ i_39_)  &  (~ i_38_)  &  n_n968  &  n_n1074 ) ;
 assign wire1905 = ( (~ i_32_)  &  i_33_  &  n_n1002  &  wire6736 ) ;
 assign wire1909 = ( (~ i_12_)  &  n_n1074  &  wire6739 ) | ( (~ i_15_)  &  n_n1074  &  wire6739 ) ;
 assign wire1910 = ( n_n1056  &  wire325  &  wire6727 ) ;
 assign wire1911 = ( n_n1047  &  wire6728  &  wire6729 ) ;
 assign wire1912 = ( (~ i_5_)  &  wire1915 ) | ( (~ i_5_)  &  wire1916 ) ;
 assign wire1913 = ( n_n884  &  wire233 ) | ( n_n884  &  wire1919 ) | ( n_n884  &  wire1920 ) ;
 assign wire1914 = ( n_n1072  &  n_n1074  &  n_n970 ) ;
 assign wire1915 = ( n_n1047  &  wire55  &  wire6728 ) ;
 assign wire1916 = ( i_31_  &  wire445  &  wire421 ) ;
 assign wire1919 = ( (~ i_40_)  &  (~ i_39_)  &  n_n874  &  n_n1009 ) ;
 assign wire1920 = ( i_40_  &  (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire1923 = ( wire363  &  wire1926 ) | ( (~ i_14_)  &  wire363  &  wire686 ) ;
 assign wire1926 = ( (~ i_12_)  &  i_11_  &  wire407 ) | ( i_12_  &  (~ i_11_)  &  wire407 ) ;
 assign wire1933 = ( n_n979  &  n_n528  &  n_n945  &  wire36 ) ;
 assign wire1934 = ( wire637  &  n_n907  &  wire6716 ) ;
 assign wire1935 = ( n_n998  &  wire46  &  wire471  &  wire400 ) ;
 assign wire1936 = ( n_n979  &  wire65  &  n_n907  &  wire6716 ) ;
 assign wire6716 = ( (~ i_13_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire6719 = ( wire1933 ) | ( wire1935 ) | ( wire1936 ) ;
 assign wire6722 = ( n_n1072  &  n_n1073  &  wire670 ) ;
 assign wire6723 = ( i_40_  &  i_39_  &  n_n1009  &  (~ wire110) ) ;
 assign wire6724 = ( wire36  &  wire45 ) ;
 assign wire6726 = ( wire537  &  wire484 ) | ( wire6723  &  wire6724 ) ;
 assign wire6727 = ( i_12_  &  (~ i_11_)  &  (~ i_32_) ) ;
 assign wire6728 = ( (~ i_32_)  &  i_31_  &  i_33_ ) ;
 assign wire6729 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_16_) ) ;
 assign wire6731 = ( (~ i_36_)  &  i_35_  &  i_37_ ) ;
 assign wire6734 = ( wire1910 ) | ( wire1911 ) | ( wire1914 ) ;
 assign wire6736 = ( i_25_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire6739 = ( (~ i_5_)  &  i_31_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire6740 = ( wire1905 ) | ( n_n969  &  n_n971  &  n_n966 ) ;
 assign wire6741 = ( wire1909 ) | ( n_n967  &  wire758 ) ;
 assign wire6746 = ( wire1896 ) | ( wire741  &  n_n907  &  wire6716 ) ;
 assign wire6747 = ( wire6746 ) | ( n_n884  &  wire742 ) ;
 assign wire6749 = ( i_9_  &  (~ i_5_)  &  i_11_  &  i_15_ ) ;
 assign wire6750 = ( i_26_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire6751 = ( i_15_  &  (~ i_12_) ) ;
 assign wire6753 = ( wire1884 ) | ( n_n1074  &  (~ wire73)  &  wire6722 ) ;
 assign wire6754 = ( wire145 ) | ( wire1881 ) | ( wire1882 ) ;
 assign wire6757 = ( wire1880 ) | ( wire1934 ) | ( wire6719 ) | ( wire6753 ) ;
 assign wire6758 = ( wire1883 ) | ( wire1923 ) | ( wire6726 ) | ( wire6754 ) ;
 assign wire6759 = ( n_n1135 ) | ( n_n1134 ) | ( wire6747 ) | ( wire6757 ) ;
 assign wire6764 = ( (~ i_40_)  &  (~ i_39_)  &  n_n985 ) ;
 assign wire6765 = ( i_40_  &  (~ i_7_)  &  i_39_ ) ;
 assign wire6766 = ( i_40_  &  i_36_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire6767 = ( wire1868 ) | ( wire330  &  n_n861  &  n_n1002 ) ;
 assign wire6770 = ( wire1871 ) | ( wire1872 ) | ( n_n515  &  wire6764 ) ;
 assign wire6772 = ( n_n1048  &  n_n1047  &  wire400 ) ;
 assign wire6773 = ( (~ i_10_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire6774 = ( (~ i_27_)  &  (~ i_39_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire6778 = ( wire153 ) | ( wire184 ) | ( wire1860 ) ;
 assign wire6779 = ( wire187 ) | ( wire1861 ) | ( wire1862 ) | ( wire1863 ) ;
 assign wire6780 = ( (~ i_5_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire6786 = ( i_12_  &  (~ i_11_)  &  wire407 ) ;
 assign wire6788 = ( (~ i_12_)  &  i_11_  &  wire407 ) ;
 assign wire6789 = ( i_22_  &  (~ i_34_)  &  (~ i_36_)  &  i_35_ ) ;
 assign wire6790 = ( i_40_  &  i_39_  &  (~ i_21_)  &  i_38_ ) ;
 assign wire6791 = ( n_n945  &  wire6789  &  wire6790 ) ;
 assign wire6793 = ( (~ i_12_)  &  i_11_  &  wire84  &  wire407 ) | ( i_12_  &  (~ i_11_)  &  wire84  &  wire407 ) ;
 assign wire6794 = ( wire1847 ) | ( wire1845 ) ;
 assign wire6798 = ( n_n1048  &  n_n1047  &  wire400 ) ;
 assign wire6800 = ( wire491  &  n_n1011  &  n_n1074  &  wire6731 ) ;
 assign wire6801 = ( n_n1011  &  n_n411  &  n_n1074  &  wire6731 ) ;
 assign wire6804 = ( wire145 ) | ( wire241 ) | ( wire1822 ) ;
 assign wire6806 = ( n_n1164 ) | ( wire6778 ) | ( wire6779 ) ;
 assign wire6807 = ( n_n1373 ) | ( wire1821 ) | ( wire6804 ) ;
 assign wire6808 = ( n_n1372 ) | ( wire1823 ) | ( wire1835 ) | ( wire1836 ) ;
 assign wire6813 = ( n_n1993 ) | ( n_n2213 ) | ( wire1812 ) ;
 assign wire6818 = ( n_n2837 ) | ( n_n1958 ) | ( n_n1956 ) | ( n_n1957 ) ;
 assign wire6821 = ( i_40_  &  i_39_  &  i_11_ ) ;
 assign wire6824 = ( (~ i_39_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_38_) ) ;
 assign wire6828 = ( (~ i_7_)  &  i_3_  &  i_0_ ) ;
 assign wire6831 = ( wire182 ) | ( wire1803 ) | ( wire1807 ) ;
 assign wire6832 = ( wire1804 ) | ( wire1806 ) | ( i_2_  &  wire835 ) ;
 assign wire6837 = ( i_19_  &  (~ i_21_) ) ;
 assign wire6839 = ( i_24_  &  i_22_  &  (~ i_32_)  &  wire609 ) ;
 assign wire6841 = ( n_n945  &  n_n860  &  wire342  &  wire6789 ) ;
 assign wire6842 = ( i_24_  &  i_22_  &  (~ i_19_) ) ;
 assign wire6844 = ( (~ i_17_)  &  (~ i_16_)  &  n_n833 ) ;
 assign wire6845 = ( (~ i_12_)  &  (~ i_31_)  &  wire45  &  wire82 ) ;
 assign wire6849 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_  &  wire94 ) ;
 assign wire6850 = ( (~ i_16_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire6851 = ( (~ i_40_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire6853 = ( n_n785  &  n_n781 ) | ( n_n777  &  wire64 ) ;
 assign wire6854 = ( wire6844  &  wire6845 ) | ( wire106  &  wire6849 ) ;
 assign wire6856 = ( i_11_  &  (~ i_17_)  &  i_15_  &  n_n793 ) ;
 assign wire6857 = ( i_12_  &  (~ i_17_)  &  i_15_  &  n_n793 ) ;
 assign wire6858 = ( (~ i_16_)  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire6859 = ( i_39_  &  (~ i_17_)  &  i_38_ ) ;
 assign wire6860 = ( wire367  &  wire479 ) | ( wire504  &  wire671 ) ;
 assign wire6861 = ( wire103  &  n_n334 ) | ( n_n313  &  wire672 ) ;
 assign wire6863 = ( (~ i_37_)  &  i_39_ ) ;
 assign wire6865 = ( i_12_  &  (~ i_18_)  &  i_15_ ) | ( i_11_  &  (~ i_18_)  &  i_15_ ) ;
 assign wire6866 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  wire6865 ) ;
 assign wire6868 = ( wire368  &  wire479 ) | ( wire366  &  wire535 ) ;
 assign wire6869 = ( wire430  &  wire6863 ) | ( wire303  &  wire6866 ) ;
 assign wire6870 = ( n_n560  &  n_n334 ) | ( wire430  &  wire837 ) ;
 assign wire6873 = ( n_n833  &  i_21_ ) ;
 assign wire6874 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_  &  (~ i_37_) ) ;
 assign wire6877 = ( n_n837  &  wire710 ) | ( wire688  &  wire6873 ) ;
 assign wire6878 = ( wire175 ) | ( wire176 ) | ( wire244 ) | ( wire1758 ) ;
 assign wire6879 = ( wire6860 ) | ( wire6861 ) | ( wire6877 ) ;
 assign wire6884 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire6886 = ( wire245 ) | ( n_n469  &  wire700 ) ;
 assign wire6887 = ( i_40_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire6888 = ( i_4_  &  n_n883  &  n_n970 ) ;
 assign wire6889 = ( i_4_  &  n_n971  &  n_n1072 ) ;
 assign wire6890 = ( i_39_  &  (~ i_36_)  &  (~ i_37_) ) ;
 assign wire6894 = ( n_n1990 ) | ( wire227 ) | ( wire1741 ) | ( wire1742 ) ;
 assign wire6897 = ( (~ i_7_)  &  i_2_  &  i_0_ ) ;
 assign wire6901 = ( wire1730 ) | ( wire422  &  n_n462  &  wire689 ) ;
 assign wire6902 = ( n_n1971 ) | ( wire1731 ) | ( wire429  &  wire711 ) ;
 assign wire6904 = ( n_n1951 ) | ( wire148 ) | ( wire6901 ) | ( wire6902 ) ;
 assign wire6907 = ( (~ i_36_)  &  i_35_  &  i_37_ ) ;
 assign wire6908 = ( (~ i_22_)  &  i_24_ ) ;
 assign wire6909 = ( wire366  &  wire529 ) | ( wire84  &  wire6856 ) ;
 assign wire6910 = ( wire64  &  n_n771 ) | ( wire84  &  wire6857 ) ;
 assign wire6911 = ( wire386  &  wire132 ) | ( n_n775  &  wire690 ) ;
 assign wire6913 = ( wire6909 ) | ( wire6910 ) | ( wire6911 ) ;
 assign wire6914 = ( wire1780 ) | ( wire6853 ) | ( wire6854 ) | ( wire6913 ) ;
 assign wire6915 = ( n_n1094 ) | ( n_n1088 ) | ( n_n1086 ) | ( wire6904 ) ;
 assign wire6920 = ( i_0_  &  (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign wire6924 = ( n_n2487 ) | ( n_n2488 ) | ( wire1705 ) | ( wire1708 ) ;
 assign wire6925 = ( wire1704 ) | ( wire1707 ) | ( wire1709 ) ;
 assign wire6927 = ( wire1706 ) | ( wire6924 ) | ( wire6925 ) ;
 assign wire6929 = ( n_n1083 ) | ( n_n1084 ) | ( wire6927 ) ;
 assign wire6930 = ( i_40_  &  i_39_  &  i_22_  &  (~ i_38_) ) ;
 assign wire6932 = ( n_n469  &  n_n945  &  wire6789 ) ;
 assign wire6933 = ( n_n1993 ) | ( n_n799  &  n_n1012  &  wire529 ) ;
 assign wire6934 = ( wire529  &  wire509 ) | ( wire366  &  wire535 ) ;
 assign wire6935 = ( wire509  &  wire535 ) | ( wire553  &  wire6932 ) ;
 assign wire6938 = ( i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign wire6940 = ( n_n799  &  n_n1012  &  wire529 ) | ( n_n799  &  n_n1012  &  wire535 ) ;
 assign wire6941 = ( wire368  &  wire479 ) | ( n_n765  &  wire101 ) ;
 assign wire6942 = ( wire430  &  wire772 ) | ( i_39_  &  (~ i_37_)  &  wire430 ) ;
 assign wire6945 = ( (~ i_39_)  &  (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire6948 = ( wire82  &  (~ i_22_) ) ;
 assign wire6949 = ( (~ i_40_)  &  i_39_  &  (~ i_23_)  &  n_n1009 ) ;
 assign wire6950 = ( wire365  &  wire337 ) | ( (~ i_22_)  &  wire82  &  wire337 ) ;
 assign wire6951 = ( wire323  &  n_n765 ) | ( (~ i_23_)  &  wire323  &  wire369 ) ;
 assign wire6952 = ( wire504  &  wire671 ) | ( n_n764  &  wire787 ) ;
 assign wire6955 = ( (~ i_40_)  &  i_39_  &  (~ i_23_)  &  n_n1009 ) ;
 assign wire6956 = ( wire329  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire6957 = ( wire367  &  wire479 ) | ( wire370  &  wire6955 ) ;
 assign wire6958 = ( n_n761  &  wire830 ) | ( n_n760  &  wire829 ) ;
 assign wire6960 = ( n_n862  &  n_n1064  &  wire529 ) | ( n_n862  &  n_n1064  &  wire535 ) ;
 assign wire6961 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire6964 = ( wire175 ) | ( wire240 ) | ( wire6960 ) | ( wire6961 ) ;
 assign wire6965 = ( n_n1611 ) | ( wire6950 ) | ( wire6951 ) | ( wire6952 ) ;
 assign wire6968 = ( (~ i_18_)  &  (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire6969 = ( i_39_  &  i_38_  &  (~ i_37_)  &  n_n979 ) ;
 assign wire6970 = ( wire84  &  wire6856 ) | ( wire84  &  wire6857 ) ;
 assign wire6971 = ( n_n775  &  n_n773 ) | ( n_n783  &  wire6969 ) ;
 assign wire6974 = ( (~ i_18_)  &  (~ i_21_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire6975 = ( (~ i_39_)  &  (~ i_38_)  &  i_37_  &  wire94 ) ;
 assign wire6976 = ( (~ i_39_)  &  (~ i_19_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire6978 = ( i_12_  &  i_15_  &  n_n793 ) | ( i_11_  &  i_15_  &  n_n793 ) ;
 assign wire6979 = ( i_40_  &  n_n979  &  n_n791  &  wire6976 ) ;
 assign wire6980 = ( i_39_  &  i_38_  &  (~ i_37_)  &  n_n979 ) ;
 assign wire6981 = ( n_n783  &  wire6975 ) | ( n_n790  &  wire6975 ) | ( n_n790  &  wire6980 ) ;
 assign wire6982 = ( wire1653 ) | ( n_n1047  &  wire400  &  wire831 ) ;
 assign wire6984 = ( n_n2581 ) | ( n_n842  &  wire335  &  n_n843 ) ;
 assign wire6985 = ( n_n2487 ) | ( n_n2488 ) | ( n_n1971 ) ;
 assign wire6987 = ( wire173 ) | ( wire6984 ) | ( wire6985 ) ;
 assign wire6991 = ( i_8_  &  (~ i_40_) ) ;
 assign wire6993 = ( (~ i_4_)  &  n_n969  &  n_n865 ) | ( (~ i_1_)  &  n_n969  &  n_n865 ) ;
 assign wire6994 = ( i_0_  &  wire79  &  wire6888 ) | ( i_0_  &  wire79  &  wire6993 ) ;
 assign wire6998 = ( n_n2837 ) | ( n_n1958 ) | ( n_n1956 ) | ( n_n1957 ) ;
 assign wire6999 = ( n_n969  &  n_n865 ) | ( n_n883  &  n_n970 ) ;
 assign wire7000 = ( n_n1990 ) | ( wire88  &  n_n975  &  wire6938 ) ;
 assign wire7001 = ( n_n1951 ) | ( i_0_  &  wire79  &  wire6889 ) ;
 assign wire7002 = ( n_n2836 ) | ( n_n2838 ) ;
 assign wire7005 = ( wire1635 ) | ( wire7000 ) | ( wire7001 ) | ( wire7002 ) ;
 assign wire7007 = ( (~ i_12_)  &  i_11_  &  i_15_ ) ;
 assign wire7008 = ( i_17_  &  i_15_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire7011 = ( i_12_  &  (~ i_11_)  &  i_15_ ) ;
 assign wire7012 = ( wire1632 ) | ( wire319  &  wire78  &  n_n527 ) ;
 assign wire7014 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  i_15_ ) ;
 assign wire7016 = ( i_12_  &  i_16_  &  i_15_ ) ;
 assign wire7018 = ( wire1624 ) | ( wire39  &  wire558  &  wire7014 ) ;
 assign wire7020 = ( n_n998  &  wire556  &  n_n861 ) | ( n_n998  &  n_n861  &  wire325 ) ;
 assign wire7021 = ( wire7020 ) | ( wire1620 ) ;
 assign wire7025 = ( wire337  &  wire6948 ) | ( wire369  &  wire6949 ) ;
 assign wire7026 = ( n_n764  &  wire359 ) | ( n_n761  &  wire101 ) | ( n_n764  &  wire101 ) ;
 assign wire7029 = ( wire368  &  wire479 ) | ( wire365  &  wire337 ) ;
 assign wire7030 = ( n_n765  &  wire825 ) | ( wire430  &  wire6863 ) ;
 assign wire7033 = ( wire329  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire7034 = ( n_n761  &  wire323 ) | ( (~ i_23_)  &  wire323  &  wire370 ) ;
 assign wire7035 = ( wire240 ) | ( wire175 ) ;
 assign wire7038 = ( wire1592 ) | ( wire7033 ) | ( wire7034 ) | ( wire7035 ) ;
 assign wire7040 = ( n_n1607 ) | ( wire6981 ) | ( wire6982 ) | ( wire7038 ) ;
 assign wire7043 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire7044 = ( (~ i_36_)  &  (~ i_34_) ) ;
 assign wire7048 = ( o_15_ ) | ( n_n980  &  wire65  &  wire7044 ) ;
 assign wire7050 = ( i_9_  &  (~ i_14_) ) | ( i_9_  &  (~ i_11_) ) ;
 assign wire7051 = ( i_17_  &  wire1579 ) | ( i_17_  &  wire7050 ) ;
 assign wire7052 = ( (~ i_12_)  &  i_9_ ) ;
 assign wire7053 = ( wire84  &  wire7051 ) | ( i_16_  &  wire84  &  wire450 ) ;
 assign wire7055 = ( (~ i_12_)  &  (~ i_35_)  &  (~ i_37_) ) | ( (~ i_11_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire7057 = ( (~ i_14_)  &  i_17_  &  i_16_ ) ;
 assign wire7058 = ( n_n1008  &  n_n1009 ) | ( n_n1011  &  n_n1012 ) ;
 assign wire7062 = ( wire1565 ) | ( wire1566 ) | ( wire1568 ) ;
 assign wire7063 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire7064 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7066 = ( (~ i_11_)  &  i_9_ ) ;
 assign wire7067 = ( (~ i_3_)  &  (~ i_4_)  &  wire45 ) ;
 assign wire7069 = ( wire1555 ) | ( n_n1074  &  (~ wire73)  &  wire6722 ) ;
 assign wire7071 = ( wire1557 ) | ( wire7069 ) | ( wire416  &  wire7066 ) ;
 assign wire7073 = ( i_40_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire7074 = ( i_5_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire7077 = ( wire1548 ) | ( wire1550 ) | ( wire1551 ) | ( wire1552 ) ;
 assign wire7079 = ( i_6_  &  i_40_ ) ;
 assign wire7086 = ( wire1542 ) | ( wire1544  &  wire7079 ) | ( wire1545  &  wire7079 ) ;
 assign wire7087 = ( wire158 ) | ( wire1539 ) | ( wire1540 ) | ( wire1541 ) ;
 assign wire7089 = ( n_n983  &  n_n977 ) | ( n_n1023  &  n_n1065 ) ;
 assign wire7090 = ( n_n1001  &  n_n1066 ) | ( n_n976  &  wire121 ) ;
 assign wire7092 = ( wire1522 ) | ( wire1525 ) | ( n_n980  &  wire560 ) ;
 assign wire7094 = ( wire1524 ) | ( wire7077 ) | ( n_n1074  &  wire817 ) ;
 assign wire7095 = ( n_n1709 ) | ( wire7086 ) | ( wire7087 ) | ( wire7092 ) ;
 assign wire7097 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_34_) ) ;
 assign wire7100 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_34_) ) ;
 assign wire7102 = ( (~ i_34_)  &  i_36_  &  i_37_ ) ;
 assign wire7103 = ( n_n1002  &  wire100 ) | ( n_n883  &  wire7102 ) ;
 assign wire7104 = ( n_n977  &  n_n715 ) | ( n_n998  &  wire121 ) ;
 assign wire7105 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_0_) ) ;
 assign wire7108 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_35_) ) ;
 assign wire7109 = ( (~ i_34_)  &  i_36_ ) | ( (~ i_34_)  &  i_35_ ) | ( i_34_  &  (~ i_36_)  &  (~ i_35_) ) ;
 assign wire7110 = ( (~ i_33_) ) | ( n_n978  &  n_n865  &  wire7100 ) ;
 assign wire7115 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign wire7118 = ( wire1499 ) | ( wire526  &  wire565 ) ;
 assign wire7119 = ( wire1496 ) | ( wire1501 ) | ( wire411  &  wire436 ) ;
 assign wire7121 = ( (~ i_40_)  &  (~ i_5_)  &  i_39_ ) ;
 assign wire7122 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire7123 = ( (~ i_28_)  &  (~ i_29_)  &  n_n985  &  wire7121 ) ;
 assign wire7124 = ( i_23_  &  i_24_  &  i_22_  &  (~ i_32_) ) ;
 assign wire7125 = ( i_15_  &  wire1834 ) | ( i_18_  &  i_15_  &  wire42 ) ;
 assign wire7127 = ( wire42  &  i_15_ ) ;
 assign wire7128 = ( i_24_  &  i_21_  &  i_22_ ) ;
 assign wire7129 = ( wire386  &  n_n935 ) | ( n_n937  &  wire775 ) | ( n_n935  &  wire775 ) ;
 assign wire7130 = ( i_9_  &  (~ i_5_)  &  (~ i_14_) ) ;
 assign wire7131 = ( n_n1066  &  n_n927  &  wire7130 ) ;
 assign wire7132 = ( (~ i_5_)  &  (~ i_14_) ) | ( (~ i_5_)  &  (~ i_12_) ) | ( (~ i_5_)  &  (~ i_11_) ) ;
 assign wire7133 = ( i_21_  &  i_23_ ) ;
 assign wire7135 = ( wire361  &  wire7123 ) | ( wire777  &  wire7131 ) ;
 assign wire7137 = ( wire333  &  wire36 ) | ( wire92  &  wire461 ) ;
 assign wire7139 = ( n_n1374 ) | ( wire1475 ) | ( n_n937  &  wire386 ) ;
 assign wire7140 = ( wire7135 ) | ( wire7137 ) | ( wire473  &  wire7125 ) ;
 assign wire7142 = ( n_n1055  &  n_n1048  &  n_n1047 ) | ( n_n1048  &  n_n1047  &  wire785 ) ;
 assign wire7143 = ( wire1468 ) | ( n_n907  &  wire782  &  wire6716 ) ;
 assign wire7145 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire7146 = ( i_22_  &  i_21_ ) ;
 assign wire7148 = ( (~ i_40_)  &  (~ i_39_)  &  i_36_  &  (~ i_38_) ) ;
 assign wire7150 = ( (~ i_14_)  &  i_40_ ) ;
 assign wire7151 = ( i_9_  &  (~ i_5_)  &  n_n933  &  n_n1066 ) ;
 assign wire7152 = ( wire1459 ) | ( wire156 ) ;
 assign wire7153 = ( n_n926  &  wire461 ) | ( wire786  &  wire7151 ) ;
 assign wire7154 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire7157 = ( (~ i_34_)  &  n_n968  &  wire46 ) | ( i_34_  &  n_n1073  &  wire46 ) ;
 assign wire7160 = ( wire1455 ) | ( n_n968  &  n_n967  &  n_n1074 ) ;
 assign wire7161 = ( wire241 ) | ( wire187 ) | ( wire1453 ) | ( wire1454 ) ;
 assign wire7164 = ( i_40_  &  i_6_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7165 = ( i_39_  &  i_12_  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7170 = ( wire184 ) | ( wire1442 ) | ( wire1444 ) ;
 assign wire7171 = ( wire158 ) | ( wire1441 ) | ( wire7170 ) ;
 assign wire7175 = ( wire140 ) | ( wire1428 ) | ( wire1429 ) ;
 assign wire7176 = ( wire1430 ) | ( wire1452 ) | ( wire7160 ) | ( wire7161 ) ;
 assign wire7178 = ( (~ i_34_)  &  (~ i_35_)  &  (~ i_37_) ) ;
 assign wire7180 = ( n_n977  &  n_n1048  &  wire7178 ) ;
 assign wire7181 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7182 = ( i_9_  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire7184 = ( wire1415 ) | ( wire1417 ) | ( wire814  &  wire7180 ) ;
 assign wire7185 = ( wire1466 ) | ( wire1467 ) | ( wire7143 ) | ( wire7184 ) ;
 assign wire7187 = ( wire1416 ) | ( wire7152 ) | ( wire7153 ) | ( wire7185 ) ;
 assign wire7189 = ( o_15_ ) | ( n_n966  &  n_n862  &  n_n1064 ) ;
 assign wire7190 = ( wire1412 ) | ( wire7189 ) | ( i_32_  &  (~ i_33_) ) ;
 assign wire7191 = ( i_33_  &  (~ i_7_) ) ;
 assign wire7193 = ( (~ i_17_)  &  (~ i_16_) ) | ( i_38_  &  i_37_ ) ;
 assign wire7194 = ( (~ i_40_)  &  i_38_ ) | ( (~ i_39_)  &  i_38_ ) | ( i_39_  &  (~ i_38_) ) | ( (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7195 = ( (~ i_7_)  &  i_5_  &  i_33_  &  n_n1047 ) ;
 assign wire7197 = ( (~ i_7_)  &  i_5_  &  (~ i_36_) ) ;
 assign wire7200 = ( i_9_  &  i_11_  &  i_15_ ) ;
 assign wire7201 = ( i_12_  &  i_16_  &  i_15_ ) ;
 assign wire7204 = ( wire301 ) | ( wire1390 ) | ( n_n967  &  n_n673 ) ;
 assign wire7205 = ( (~ i_40_)  &  i_9_  &  (~ i_7_) ) ;
 assign wire7208 = ( wire59  &  wire1388 ) | ( wire59  &  wire1389 ) ;
 assign wire7210 = ( wire354  &  wire7208 ) | ( wire354  &  wire788  &  wire7200 ) ;
 assign wire7211 = ( wire1383 ) | ( wire1386 ) | ( n_n973  &  n_n673 ) ;
 assign wire7214 = ( (~ i_40_)  &  (~ i_39_)  &  i_38_  &  i_37_ ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7218 = ( wire1372 ) | ( (~ i_14_)  &  n_n1066  &  wire7197 ) ;
 assign wire7219 = ( wire1374 ) | ( wire1371 ) ;
 assign wire7220 = ( wire183 ) | ( wire251 ) | ( wire1375 ) ;
 assign wire7223 = ( n_n1528 ) | ( wire7218 ) | ( wire7219 ) | ( wire7220 ) ;
 assign wire7227 = ( i_0_  &  (~ i_32_)  &  i_33_  &  i_37_ ) ;
 assign wire7230 = ( wire413 ) | ( wire1365 ) | ( wire1366 ) | ( wire1367 ) ;
 assign wire7231 = ( (~ i_34_)  &  i_33_  &  i_38_  &  i_37_ ) ;
 assign wire7233 = ( (~ i_40_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7234 = ( n_n1073  &  n_n700 ) | ( n_n1074  &  wire7233 ) ;
 assign wire7237 = ( wire1353 ) | ( wire1354 ) | ( n_n880  &  wire803 ) ;
 assign wire7239 = ( i_39_  &  (~ i_32_)  &  i_33_  &  i_38_ ) ;
 assign wire7245 = ( wire303 ) | ( wire1346 ) | ( wire1347 ) | ( wire1348 ) ;
 assign wire7246 = ( i_0_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7252 = ( wire336 ) | ( wire1340 ) | ( wire1341 ) | ( wire1342 ) ;
 assign wire7253 = ( (~ i_9_)  &  i_39_  &  (~ i_16_) ) ;
 assign wire7256 = ( (~ i_34_)  &  i_35_  &  i_38_  &  i_37_ ) ;
 assign wire7257 = ( (~ i_9_)  &  i_39_  &  i_38_ ) ;
 assign wire7258 = ( i_35_  &  i_38_  &  i_37_ ) ;
 assign wire7260 = ( wire1328 ) | ( n_n710  &  wire811 ) ;
 assign wire7261 = ( wire1329 ) | ( wire1330 ) | ( wire77  &  wire809 ) ;
 assign wire7263 = ( (~ i_34_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7265 = ( i_7_  &  i_33_ ) | ( n_n1047  &  wire6728 ) ;
 assign wire7266 = ( n_n980  &  n_n1047 ) | ( n_n980  &  wire7263 ) ;
 assign wire7269 = ( wire1316 ) | ( wire1317 ) | ( wire7265 ) | ( wire7266 ) ;
 assign wire7270 = ( wire1349 ) | ( wire1364 ) | ( wire7230 ) | ( wire7245 ) ;
 assign wire7271 = ( wire1343 ) | ( wire1344 ) | ( wire7252 ) | ( wire7269 ) ;
 assign wire7275 = ( (~ i_40_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire7276 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_13_) ) ;
 assign wire7278 = ( (~ i_37_)  &  (~ i_39_) ) ;
 assign wire7279 = ( i_40_  &  (~ i_30_)  &  (~ i_39_)  &  i_38_ ) ;
 assign wire7281 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_34_) ) ;
 assign wire7284 = ( wire1307 ) | ( wire47  &  wire320  &  wire761 ) ;
 assign wire7285 = ( n_n2213 ) | ( wire1306 ) | ( wire1309 ) ;
 assign wire7286 = ( wire1305 ) | ( wire488  &  wire1311 ) | ( wire488  &  wire1312 ) ;
 assign wire7291 = ( (~ i_31_)  &  i_33_  &  n_n1047  &  n_n795 ) ;
 assign wire7293 = ( wire1294 ) | ( n_n1052  &  wire762 ) ;
 assign wire7295 = ( (~ i_31_)  &  i_33_  &  n_n883  &  n_n1047 ) ;
 assign wire7299 = ( wire1286 ) | ( wire43  &  wire7295 ) | ( wire1291  &  wire7295 ) ;
 assign wire7301 = ( wire7284 ) | ( wire7285 ) | ( wire7286 ) | ( wire7299 ) ;
 assign wire7302 = ( wire1284 ) | ( wire1285 ) | ( wire1295 ) | ( wire7293 ) ;
 assign wire7304 = ( i_23_  &  i_24_  &  n_n833 ) ;
 assign wire7305 = ( wire35  &  n_n848  &  wire50 ) ;
 assign wire7306 = ( i_15_  &  (~ i_34_)  &  i_33_ ) ;
 assign wire7308 = ( i_9_  &  (~ i_7_)  &  (~ wire73)  &  wire7306 ) ;
 assign wire7309 = ( (~ i_7_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire7311 = ( wire327  &  n_n550 ) | ( wire7304  &  wire7305 ) ;
 assign wire7314 = ( (~ i_40_)  &  (~ i_31_)  &  (~ i_34_)  &  i_33_ ) ;
 assign wire7317 = ( (~ i_39_)  &  (~ i_38_)  &  n_n888 ) ;
 assign wire7319 = ( wire1271 ) | ( n_n1008  &  wire411  &  n_n698 ) ;
 assign wire7320 = ( wire364  &  wire336 ) | ( n_n560  &  n_n550 ) ;
 assign wire7321 = ( n_n556  &  wire139 ) | ( n_n559  &  wire7317 ) | ( n_n556  &  wire7317 ) ;
 assign wire7323 = ( wire86  &  wire320  &  n_n860 ) | ( wire320  &  wire78  &  n_n860 ) ;
 assign wire7324 = ( i_40_  &  i_39_  &  (~ i_36_)  &  (~ i_38_) ) ;
 assign wire7325 = ( (~ i_40_)  &  (~ i_39_)  &  (~ i_36_)  &  i_38_ ) ;
 assign wire7329 = ( wire1264 ) | ( wire1265 ) | ( wire526  &  wire724 ) ;
 assign wire7330 = ( (~ i_40_)  &  i_39_  &  (~ i_37_) ) ;
 assign wire7332 = ( (~ i_40_)  &  i_39_  &  i_37_ ) ;
 assign wire7333 = ( i_37_  &  i_39_ ) ;
 assign wire7334 = ( n_n709  &  n_n1002 ) | ( n_n991  &  wire7333 ) ;
 assign wire7336 = ( n_n2439 ) | ( wire1257 ) | ( wire1262 ) ;
 assign wire7337 = ( wire1253 ) | ( wire1255 ) | ( wire1256 ) ;
 assign wire7339 = ( i_36_  &  wire1251 ) | ( i_36_  &  wire1252 ) ;
 assign wire7341 = ( n_n1777 ) | ( (~ i_7_)  &  wire45  &  wire7339 ) ;
 assign wire7342 = ( wire1246 ) | ( wire1247 ) | ( n_n991  &  wire766 ) ;
 assign wire7343 = ( wire1238 ) | ( i_32_  &  n_n1047  &  wire7191 ) ;
 assign wire7344 = ( wire1254 ) | ( wire7336 ) | ( wire7337 ) | ( wire7343 ) ;
 assign wire7345 = ( wire7341 ) | ( wire7342 ) | ( wire7344 ) ;
 assign wire7347 = ( (~ i_23_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7348 = ( n_n979  &  wire35  &  n_n848 ) ;
 assign wire7349 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_21_) ) ;
 assign wire7350 = ( n_n859  &  wire7349 ) | ( wire1797  &  wire7349 ) | ( wire1798  &  wire7349 ) ;
 assign wire7353 = ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) | ( (~ i_39_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire7354 = ( n_n1986 ) | ( wire240 ) ;
 assign wire7355 = ( wire245 ) | ( n_n469  &  wire7347  &  wire7348 ) ;
 assign wire7356 = ( n_n1971 ) | ( wire1230 ) | ( wire335  &  wire396 ) ;
 assign wire7359 = ( wire7353 ) | ( wire7354 ) | ( wire7355 ) | ( wire7356 ) ;
 assign wire7360 = ( (~ i_39_)  &  (~ i_32_)  &  i_34_  &  i_33_ ) ;
 assign wire7362 = ( n_n1951 ) | ( n_n842  &  wire335  &  n_n843 ) ;
 assign wire7363 = ( n_n1986 ) | ( wire1222 ) ;
 assign wire7367 = ( o_32_ ) | ( n_n1993 ) | ( n_n2836 ) ;
 assign wire7371 = ( n_n2837 ) | ( n_n1958 ) | ( n_n1956 ) | ( n_n1957 ) ;
 assign wire7372 = ( n_n1074  &  wire6828 ) | ( n_n1074  &  wire6897 ) ;
 assign wire7373 = ( n_n2487 ) | ( n_n2488 ) | ( n_n1990 ) ;
 assign wire7375 = ( wire149 ) | ( wire1213 ) | ( wire7373 ) ;
 assign wire7377 = ( n_n862  &  n_n1064  &  wire529 ) | ( n_n862  &  n_n1064  &  wire535 ) ;
 assign wire7378 = ( wire175 ) | ( (~ i_40_)  &  (~ i_38_)  &  wire542 ) ;
 assign wire7383 = ( wire245 ) | ( wire176 ) | ( wire185 ) | ( wire7378 ) ;
 assign wire7384 = ( n_n1581 ) | ( n_n1113 ) | ( n_n1580 ) | ( wire7377 ) ;
 assign wire7388 = ( (~ i_40_)  &  (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire7389 = ( i_30_  &  (~ i_28_)  &  i_29_ ) ;
 assign wire7390 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7392 = ( wire1208 ) | ( (~ i_5_)  &  n_n462  &  wire468 ) ;
 assign wire7394 = ( (~ i_40_)  &  i_10_  &  i_27_  &  (~ i_39_) ) ;
 assign wire7396 = ( i_0_  &  i_2_ ) ;
 assign wire7397 = ( i_0_  &  i_3_ ) ;
 assign wire7398 = ( i_40_  &  i_39_  &  n_n1061 ) ;
 assign wire7399 = ( (~ i_24_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7403 = ( wire154 ) | ( wire1199 ) | ( wire1200 ) ;
 assign wire7405 = ( (~ i_24_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7406 = ( (~ i_22_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7411 = ( wire1186 ) | ( wire1189 ) | ( wire406  &  wire467 ) ;
 assign wire7412 = ( wire7411 ) | ( n_n1001  &  wire616 ) ;
 assign wire7414 = ( i_15_  &  (~ i_17_) ) ;
 assign wire7415 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7416 = ( (~ i_39_)  &  (~ i_38_)  &  n_n1012  &  wire76 ) ;
 assign wire7417 = ( wire1182 ) | ( n_n947  &  (~ wire37)  &  wire7416 ) ;
 assign wire7420 = ( (~ i_17_)  &  (~ i_16_)  &  wire76 ) ;
 assign wire7421 = ( n_n1072  &  n_n1073  &  wire36 ) ;
 assign wire7423 = ( (~ i_40_)  &  i_38_  &  n_n1073 ) ;
 assign wire7427 = ( wire7420  &  wire7421 ) | ( wire695  &  wire7423 ) ;
 assign wire7428 = ( i_39_  &  (~ i_36_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7430 = ( wire1164 ) | ( wire1165 ) | ( n_n475  &  wire617 ) ;
 assign wire7432 = ( wire1163 ) | ( wire7430 ) | ( wire113  &  wire7428 ) ;
 assign wire7435 = ( (~ i_4_)  &  i_0_  &  i_36_ ) ;
 assign wire7440 = ( wire1156 ) | ( n_n998  &  wire46  &  wire676 ) ;
 assign wire7441 = ( (~ i_9_)  &  (~ i_5_)  &  wire76 ) ;
 assign wire7442 = ( (~ i_40_)  &  i_36_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7443 = ( i_0_  &  i_4_ ) ;
 assign wire7444 = ( wire332  &  wire678 ) | ( wire679  &  wire7441 ) ;
 assign wire7445 = ( wire394  &  wire69 ) | ( wire680  &  wire7442 ) ;
 assign wire7446 = ( wire1139 ) | ( i_7_  &  i_33_ ) ;
 assign wire7447 = ( wire1155 ) | ( wire1158 ) | ( wire7440 ) | ( wire7446 ) ;
 assign wire7450 = ( (~ i_21_)  &  i_15_  &  n_n850  &  wire822 ) ;
 assign wire7451 = ( i_39_  &  i_38_  &  n_n968 ) ;
 assign wire7452 = ( (~ i_40_)  &  i_39_  &  (~ i_23_)  &  i_38_ ) ;
 assign wire7453 = ( n_n819  &  wire386 ) | ( wire99  &  wire7450 ) ;
 assign wire7454 = ( wire82  &  wire475 ) | ( wire132  &  wire7451 ) ;
 assign wire7456 = ( (~ i_21_)  &  i_15_  &  wire572  &  n_n853 ) ;
 assign wire7458 = ( n_n1971 ) | ( wire48  &  n_n850  &  wire337 ) ;
 assign wire7459 = ( wire365  &  wire337 ) | ( (~ i_22_)  &  wire87  &  wire337 ) ;
 assign wire7460 = ( wire337  &  wire6948 ) | ( wire99  &  wire7456 ) ;
 assign wire7463 = ( wire1122 ) | ( wire7458 ) | ( wire7459 ) | ( wire7460 ) ;
 assign wire7466 = ( i_40_  &  (~ i_39_)  &  n_n985 ) | ( i_40_  &  i_39_  &  n_n1009 ) ;
 assign wire7467 = ( n_n1064  &  n_n993 ) | ( n_n1073  &  n_n1015 ) ;
 assign wire7473 = ( (~ i_39_)  &  (~ i_36_)  &  i_38_ ) | ( (~ i_36_)  &  (~ i_38_)  &  (~ i_37_) ) ;
 assign wire7474 = ( i_39_  &  (~ i_36_)  &  (~ i_38_) ) | ( (~ i_36_)  &  i_38_  &  i_37_ ) ;
 assign wire7476 = ( (~ i_7_)  &  i_31_  &  wire45 ) ;
 assign wire7478 = ( wire251 ) | ( wire1093 ) | ( wire718  &  wire7476 ) ;
 assign wire7479 = ( (~ i_7_)  &  (~ i_34_)  &  (~ i_36_) ) ;
 assign wire7482 = ( (~ i_7_)  &  (~ i_14_) ) | ( (~ i_7_)  &  (~ i_12_) ) | ( (~ i_7_)  &  (~ i_11_) ) ;
 assign wire7487 = ( wire1089 ) | ( wire1090 ) | ( wire1091 ) ;
 assign wire7488 = ( i_9_  &  (~ i_7_)  &  n_n1055  &  n_n1047 ) ;
 assign wire7492 = ( (~ i_7_)  &  n_n1047  &  wire400 ) ;
 assign wire7493 = ( wire1075 ) | ( wire737  &  wire7492 ) ;
 assign wire7494 = ( wire1073 ) | ( wire1088 ) | ( wire1092 ) | ( wire7487 ) ;
 assign wire7495 = ( wire1083 ) | ( wire7493 ) | ( wire692  &  wire7488 ) ;
 assign wire7498 = ( wire183 ) | ( wire1060 ) | ( wire1063 ) ;
 assign wire7500 = ( (~ i_38_)  &  (~ i_7_) ) ;
 assign wire7504 = ( wire182 ) | ( wire301 ) | ( wire1049 ) | ( wire1051 ) ;
 assign wire7506 = ( wire1050 ) | ( wire1112 ) | ( wire1113 ) | ( wire7504 ) ;
 assign wire7508 = ( n_n1489 ) | ( wire7494 ) | ( wire7495 ) | ( wire7506 ) ;
 assign wire7509 = ( wire731  &  i_24_ ) ;
 assign wire7510 = ( i_39_  &  i_23_  &  i_38_ ) ;
 assign wire7511 = ( i_25_  &  i_21_  &  i_22_  &  i_15_ ) ;
 assign wire7512 = ( (~ i_32_)  &  i_33_  &  n_n998  &  n_n973 ) ;
 assign wire7514 = ( wire87  &  n_n428 ) | ( n_n428  &  wire82 ) ;
 assign wire7517 = ( (~ i_7_)  &  (~ i_5_)  &  i_11_  &  n_n848 ) ;
 assign wire7518 = ( n_n982  &  n_n998  &  n_n861 ) | ( n_n998  &  n_n861  &  wire325 ) ;
 assign wire7519 = ( wire7518 ) | ( i_25_  &  wire575 ) ;
 assign wire7521 = ( n_n411  &  wire1834 ) | ( i_18_  &  n_n411  &  wire42 ) ;
 assign wire7522 = ( wire491  &  n_n978  &  n_n1074  &  wire6731 ) ;
 assign wire7523 = ( i_7_  &  i_33_ ) | ( wire84  &  wire6786 ) ;
 assign wire7524 = ( wire84  &  wire6788 ) | ( wire361  &  wire7123 ) ;
 assign wire7529 = ( n_n1373 ) | ( n_n1372 ) | ( wire1021 ) | ( wire1022 ) ;
 assign wire7530 = ( wire1019 ) | ( wire1020 ) | ( wire7523 ) | ( wire7524 ) ;
 assign wire7531 = ( i_40_  &  i_39_  &  i_12_  &  (~ i_11_) ) ;
 assign wire7535 = ( (~ i_12_)  &  i_11_  &  wire84  &  wire407 ) | ( i_12_  &  (~ i_11_)  &  wire84  &  wire407 ) ;
 assign wire7536 = ( wire140 ) | ( n_n1066  &  wire7122  &  wire7123 ) ;
 assign wire7538 = ( wire146 ) | ( wire153 ) | ( wire1008 ) | ( wire1010 ) ;
 assign wire7540 = ( wire156 ) | ( wire7536 ) | ( wire386  &  n_n935 ) ;
 assign wire7541 = ( wire1412 ) | ( wire7189 ) | ( wire7535 ) | ( wire7538 ) ;
 assign wire7542 = ( i_40_  &  i_39_  &  i_38_  &  n_n968 ) | ( (~ i_40_)  &  (~ i_39_)  &  (~ i_38_)  &  n_n968 ) ;
 assign wire7544 = ( wire333  &  wire581 ) | ( wire583  &  wire7542 ) ;
 assign wire7545 = ( wire473  &  wire7125 ) | ( i_19_  &  wire473  &  wire739 ) ;
 assign wire7547 = ( n_n1372 ) | ( wire999 ) | ( wire1835 ) | ( wire1836 ) ;
 assign wire7548 = ( n_n1373 ) | ( wire1000 ) | ( wire7544 ) | ( wire7545 ) ;
 assign wire7550 = ( o_15_ ) | ( wire45  &  n_n693  &  wire7531 ) ;
 assign wire7554 = ( n_n2439 ) | ( wire985 ) | ( wire987 ) | ( wire988 ) ;
 assign wire7555 = ( n_n2837 ) | ( n_n2838 ) ;
 assign wire7557 = ( (~ i_22_)  &  wire80  &  wire7145 ) ;
 assign wire7558 = ( n_n469  &  (~ i_23_) ) ;
 assign wire7559 = ( wire176 ) | ( wire87  &  wire7557 ) | ( wire82  &  wire7557 ) ;
 assign wire7560 = ( n_n760  &  wire595 ) | ( wire598  &  wire7558 ) ;
 assign wire7562 = ( (~ i_23_)  &  (~ i_21_)  &  i_15_  &  n_n850 ) ;
 assign wire7563 = ( (~ i_40_)  &  (~ i_39_)  &  wire422  &  n_n1009 ) ;
 assign wire7564 = ( i_40_  &  (~ i_39_)  &  n_n1052 ) ;
 assign wire7565 = ( wire529  &  wire509 ) | ( wire335  &  wire396 ) ;
 assign wire7566 = ( wire432  &  wire7562 ) | ( wire408  &  wire7563 ) ;
 assign wire7568 = ( n_n560  &  n_n334 ) | ( n_n525  &  wire7564 ) ;
 assign wire7570 = ( wire973 ) | ( wire7566 ) | ( (~ i_38_)  &  wire542 ) ;
 assign wire7571 = ( wire7565 ) | ( wire7568 ) | ( i_40_  &  wire148 ) ;
 assign wire7572 = ( wire48  &  n_n853  &  wire50 ) | ( wire48  &  wire50  &  n_n850 ) ;
 assign wire7574 = ( wire962 ) | ( wire964 ) | ( wire395  &  wire600 ) ;
 assign wire7576 = ( (~ i_23_)  &  (~ i_21_)  &  i_15_  &  n_n853 ) ;
 assign wire7577 = ( wire368  &  wire479 ) | ( wire432  &  wire7576 ) ;
 assign wire7578 = ( wire430  &  wire837 ) | ( i_39_  &  (~ i_37_)  &  wire430 ) ;
 assign wire7582 = ( wire84  &  wire6856 ) | ( wire84  &  wire6857 ) ;
 assign wire7583 = ( n_n777  &  wire356 ) | ( wire83  &  wire643 ) ;
 assign wire7586 = ( (~ i_14_)  &  i_12_  &  i_15_ ) ;
 assign wire7588 = ( (~ i_18_)  &  n_n979  &  n_n791  &  wire6976 ) ;
 assign wire7590 = ( wire648  &  wire646 ) | ( wire486  &  wire7588 ) ;
 assign wire7591 = ( wire942 ) | ( wire7590 ) | ( n_n771  &  wire356 ) ;
 assign wire7593 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_29_) ) ;
 assign wire7596 = ( n_n2487 ) | ( n_n2488 ) | ( wire937 ) ;
 assign wire7597 = ( wire940 ) | ( (~ i_36_)  &  wire68  &  n_n329 ) ;
 assign wire7601 = ( (~ i_7_)  &  (~ i_5_)  &  i_28_ ) | ( (~ i_7_)  &  (~ i_5_)  &  i_29_ ) ;
 assign wire7602 = ( (~ i_34_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7605 = ( wire929 ) | ( wire928 ) ;
 assign wire7610 = ( wire420  &  n_n1048  &  n_n1047 ) | ( n_n1048  &  n_n1047  &  wire6884 ) ;
 assign wire7612 = ( wire244 ) | ( wire911 ) | ( wire103  &  n_n334 ) ;
 assign wire7614 = ( wire939 ) | ( wire7596 ) | ( wire7597 ) | ( wire7612 ) ;
 assign wire7615 = ( n_n1277 ) | ( wire912 ) | ( wire913 ) ;
 assign wire7616 = ( n_n1283 ) | ( n_n1285 ) | ( wire7591 ) | ( wire7614 ) ;
 assign wire7620 = ( (~ i_7_)  &  i_12_  &  (~ i_32_) ) ;
 assign wire7624 = ( n_n1957 ) | ( wire904 ) | ( wire905 ) ;
 assign wire7625 = ( n_n2836 ) | ( n_n1958 ) | ( n_n1956 ) | ( wire906 ) ;
 assign wire7626 = ( (~ i_7_)  &  i_11_  &  (~ i_32_) ) ;
 assign wire7627 = ( (~ i_40_)  &  i_39_  &  i_0_ ) ;
 assign wire7630 = ( (~ i_40_)  &  i_35_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7631 = ( i_0_  &  i_4_ ) ;
 assign wire7632 = ( n_n1074  &  wire6828 ) | ( (~ i_7_)  &  n_n1074  &  wire318 ) ;
 assign wire7634 = ( wire894 ) | ( wire890 ) ;
 assign wire7636 = ( wire986 ) | ( wire7554 ) | ( wire7555 ) | ( wire7634 ) ;
 assign wire7637 = ( wire131 ) | ( wire891 ) | ( wire892 ) | ( wire893 ) ;
 assign wire7639 = ( wire7624 ) | ( wire7625 ) | ( wire7636 ) | ( wire7637 ) ;
 assign wire7640 = ( (~ i_40_)  &  i_39_  &  n_n1009  &  n_n860 ) ;
 assign wire7641 = ( (~ i_39_)  &  (~ i_38_)  &  n_n888 ) ;
 assign wire7643 = ( wire321  &  wire506 ) | ( wire106  &  wire7641 ) ;
 assign wire7645 = ( i_40_  &  i_38_  &  (~ i_37_) ) ;
 assign wire7646 = ( i_11_  &  i_15_  &  wire7645 ) ;
 assign wire7647 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  n_n411 ) ;
 assign wire7648 = ( wire491  &  i_15_ ) ;
 assign wire7649 = ( i_40_  &  (~ i_38_)  &  n_n1074  &  wire6731 ) ;
 assign wire7650 = ( wire7304  &  wire7305 ) | ( wire433  &  wire7646 ) ;
 assign wire7654 = ( wire873 ) | ( n_n888  &  wire875 ) | ( n_n888  &  wire876 ) ;
 assign wire7655 = ( wire872 ) | ( (~ i_40_)  &  (~ i_39_)  &  wire508 ) ;
 assign wire7658 = ( wire131 ) | ( n_n2439 ) | ( wire1262 ) ;
 assign wire7659 = ( wire864 ) | ( wire865 ) | ( n_n795  &  wire752 ) ;
 assign wire7661 = ( (~ i_31_)  &  wire45  &  n_n462 ) ;
 assign wire7663 = ( wire860 ) | ( n_n329  &  wire1546 ) | ( n_n329  &  wire1547 ) ;
 assign wire7664 = ( wire244 ) | ( wire859 ) | ( wire102  &  wire7661 ) ;
 assign wire7666 = ( wire357  &  n_n329 ) | ( n_n560  &  n_n334 ) ;
 assign wire7667 = ( wire850 ) | ( n_n833  &  n_n525 ) | ( n_n525  &  wire304 ) ;
 assign wire7669 = ( wire7666 ) | ( wire7667 ) | ( n_n515  &  wire92 ) ;
 assign wire7670 = ( i_40_  &  (~ i_39_)  &  i_24_  &  (~ i_37_) ) ;
 assign wire7673 = ( wire519 ) | ( wire533 ) | ( wire538 ) ;
 assign wire7674 = ( wire7663 ) | ( wire7664 ) | ( wire7673 ) ;
 assign wire7676 = ( i_40_  &  (~ i_38_)  &  i_37_  &  n_n979 ) ;
 assign wire7677 = ( n_n973  &  n_n966  &  n_n1012 ) ;
 assign wire7679 = ( i_40_  &  i_15_  &  n_n945  &  wire6789 ) ;
 assign wire7680 = ( wire587  &  wire7676 ) | ( wire364  &  wire7677 ) ;
 assign wire7681 = ( wire7680 ) | ( i_38_  &  (~ i_37_)  &  wire586 ) ;
 assign wire7683 = ( n_n1326 ) | ( wire7658 ) | ( wire7659 ) | ( wire7681 ) ;
 assign wire7686 = ( (~ i_5_)  &  (~ i_12_)  &  i_15_ ) ;
 assign wire7689 = ( (~ i_5_)  &  i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7692 = ( wire455 ) | ( wire81  &  n_n162 ) | ( wire81  &  n_n164 ) ;
 assign wire7694 = ( (~ i_23_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7698 = ( i_39_  &  (~ i_16_)  &  i_15_ ) ;
 assign wire7704 = ( wire154 ) | ( wire309 ) | ( wire310 ) | ( wire312 ) ;
 assign wire7705 = ( wire7704 ) | ( wire311 ) ;
 assign wire7707 = ( i_40_  &  (~ i_16_)  &  i_15_  &  (~ i_38_) ) ;
 assign wire7715 = ( wire298 ) | ( wire524  &  n_n836 ) | ( wire524  &  wire299 ) ;
 assign wire7717 = ( i_14_  &  i_15_ ) | ( (~ i_17_)  &  i_15_ ) ;
 assign wire7722 = ( (~ i_18_)  &  (~ i_21_)  &  i_15_ ) ;
 assign wire7726 = ( i_9_  &  i_17_ ) | ( i_9_  &  i_16_ ) ;
 assign wire7728 = ( wire276 ) | ( wire303  &  wire655  &  wire7722 ) ;
 assign wire7730 = ( wire279 ) | ( wire7728 ) | ( n_n1068  &  wire520 ) ;
 assign wire7734 = ( o_15_ ) | ( n_n1021  &  n_n1074  &  wire664 ) ;
 assign wire7737 = ( wire7734 ) | ( wire263 ) ;
 assign wire7738 = ( wire260 ) | ( wire261 ) | ( wire262 ) | ( wire264 ) ;
 assign wire7741 = ( n_n1066  &  n_n453 ) | ( n_n1066  &  n_n458 ) ;
 assign wire7742 = ( i_4_  &  i_0_  &  wire45 ) | ( i_1_  &  i_0_  &  wire45 ) ;
 assign wire7743 = ( i_40_  &  i_36_  &  i_37_ ) ;
 assign wire7745 = ( i_12_  &  (~ i_11_)  &  i_36_ ) ;
 assign wire7747 = ( wire248 ) | ( wire250 ) | ( wire252 ) ;
 assign wire7750 = ( (~ i_4_)  &  i_0_ ) | ( (~ i_1_)  &  i_0_ ) ;
 assign wire7754 = ( wire153 ) | ( wire229 ) | ( wire232 ) | ( wire235 ) ;
 assign wire7755 = ( wire231 ) | ( wire234 ) | ( wire403  &  wire684 ) ;
 assign wire7756 = ( (~ i_32_)  &  n_n1066  &  wire7396 ) | ( (~ i_32_)  &  n_n1066  &  wire7443 ) ;
 assign wire7757 = ( i_40_  &  i_39_  &  i_36_  &  i_38_ ) ;
 assign wire7760 = ( (~ i_5_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire7761 = ( wire217 ) | ( wire69  &  wire7757 ) | ( wire7756  &  wire7757 ) ;
 assign wire7762 = ( wire218 ) | ( wire7754 ) | ( wire7755 ) ;
 assign wire7763 = ( wire243 ) | ( wire249 ) | ( wire7747 ) | ( wire7761 ) ;
 assign wire7764 = ( n_n1193 ) | ( n_n1195 ) | ( wire7705 ) | ( wire7762 ) ;
 assign wire7767 = ( i_12_  &  (~ i_11_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7770 = ( i_25_  &  (~ i_39_) ) ;
 assign wire7771 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_16_) ) ;
 assign wire7772 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7774 = ( wire208 ) | ( wire209 ) | ( wire210 ) ;
 assign wire7775 = ( wire213 ) | ( wire211 ) ;
 assign wire7777 = ( i_39_  &  (~ i_36_)  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7784 = ( wire199 ) | ( wire198 ) ;
 assign wire7785 = ( wire201 ) | ( (~ i_13_)  &  wire45  &  wire506 ) ;
 assign wire7786 = ( wire205 ) | ( n_n1055  &  n_n1047  &  wire463 ) ;
 assign wire7791 = ( wire188 ) | ( wire190 ) | ( wire193 ) ;
 assign wire7793 = ( wire189 ) | ( wire191 ) | ( wire192 ) | ( wire7791 ) ;
 assign wire7795 = ( (~ i_26_)  &  (~ i_39_) ) ;
 assign wire7796 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_12_) ) ;
 assign wire7799 = ( n_n2581 ) | ( wire167 ) | ( wire170 ) ;
 assign wire7800 = ( wire165 ) | ( wire169 ) | ( wire171 ) ;
 assign wire7803 = ( (~ i_34_)  &  i_36_  &  (~ i_37_) ) ;
 assign wire7805 = ( (~ i_40_)  &  (~ i_39_)  &  i_37_ ) ;
 assign wire7806 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_17_) ) ;
 assign wire7807 = ( wire162 ) | ( (~ i_40_)  &  n_n862 ) | ( (~ i_39_)  &  n_n862 ) ;
 assign wire7808 = ( wire164 ) | ( wire163 ) ;
 assign wire7809 = ( (~ i_32_)  &  i_31_  &  (~ i_34_)  &  i_33_ ) ;
 assign wire7811 = ( wire142 ) | ( wire143 ) | ( wire151 ) ;
 assign wire7812 = ( wire144 ) | ( (~ i_39_)  &  wire508 ) ;
 assign wire7814 = ( wire7811 ) | ( wire7812 ) | ( wire47  &  wire604 ) ;
 assign wire7815 = ( i_9_  &  (~ i_7_)  &  (~ i_5_)  &  (~ i_21_) ) ;
 assign wire7816 = ( i_40_  &  i_23_  &  (~ i_38_)  &  i_37_ ) ;
 assign wire7817 = ( i_17_  &  i_15_  &  (~ i_32_)  &  i_33_ ) ;
 assign wire7818 = ( (~ i_12_)  &  i_11_  &  i_15_ ) ;
 assign wire7819 = ( (~ i_14_)  &  i_12_  &  i_15_ ) ;
 assign wire7820 = ( n_n860  &  wire104 ) | ( n_n860  &  wire38  &  wire7011 ) ;
 assign wire7821 = ( wire74 ) | ( n_n775  &  wire483 ) | ( n_n775  &  wire7820 ) ;
 assign wire7822 = ( n_n1242 ) | ( n_n1235 ) | ( wire7814 ) ;


endmodule

