module bigkey (
	pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_, pkey_243_, pcount_2_, 
	pkey_4_, pkey_132_, pkey_143_, pkey_158_, pkey_169_, pkey_231_, pkey_242_, pcount_1_, pkey_7_, pkey_146_, 
	pkey_159_, pkey_168_, pkey_245_, pcount_0_, pkey_6_, pkey_130_, pkey_145_, pkey_167_, pkey_244_, pkey_9_, 
	pkey_16_, pkey_27_, pkey_38_, pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_, pkey_221_, pkey_247_, 
	pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_39_, pkey_48_, pkey_110_, pkey_121_, pkey_147_, pkey_154_, 
	pkey_165_, pkey_220_, pkey_246_, pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_47_, pkey_111_, pkey_120_, 
	pkey_155_, pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_, pkey_37_, pkey_46_, pkey_112_, 
	pkey_149_, pkey_156_, pkey_163_, pkey_211_, pkey_248_, pkey_255_, pkey_56_, pkey_67_, pkey_78_, pkey_89_, 
	pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_, pkey_238_, pkey_57_, pkey_66_, pkey_79_, 
	pkey_88_, pkey_114_, pkey_125_, pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_239_, pkey_58_, pkey_69_, 
	pkey_76_, pkey_87_, pkey_115_, pkey_124_, pkey_137_, pkey_151_, pkey_160_, pkey_214_, pkey_223_, pkey_236_, 
	pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_, pkey_123_, pkey_138_, pkey_152_, pkey_215_, 
	pkey_222_, pkey_237_, pkey_251_, pkey_1_, pkey_96_, pkey_117_, pkey_135_, pkey_140_, pkey_216_, pkey_229_, 
	pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_, pkey_217_, pkey_228_, pkey_235_, pkey_3_, 
	pkey_98_, pkey_119_, pkey_128_, pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_, pkey_2_, 
	pkey_99_, pkey_127_, pkey_134_, pkey_141_, pkey_219_, pkey_226_, pkey_233_, pkey_240_, pkey_70_, pkey_81_, 
	pkey_92_, pkey_108_, pkey_180_, pkey_193_, pkey_207_, pkey_71_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, 
	pkey_206_, pclk, pkey_50_, pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_, pstart_0_, pkey_51_, 
	pkey_60_, pkey_95_, pkey_109_, pkey_181_, pkey_196_, pkey_208_, pkey_52_, pkey_63_, pkey_74_, pkey_85_, 
	pkey_104_, pkey_171_, pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_, pkey_75_, pkey_84_, pkey_103_, 
	pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_, pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_199_, 
	pkey_205_, pkey_55_, pkey_64_, pkey_73_, pkey_82_, pkey_91_, pkey_105_, pkey_170_, pkey_204_, pkey_12_, 
	pkey_23_, pkey_34_, pkey_45_, pkey_100_, pkey_175_, pkey_188_, pkey_13_, pkey_22_, pkey_35_, pkey_44_, 
	pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_, pkey_102_, pkey_173_, pkey_201_, pkey_15_, 
	pkey_24_, pkey_33_, pkey_42_, pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_, pkey_179_, 
	pkey_184_, pkey_31_, pkey_40_, pkey_183_, pkey_190_, pkey_10_, pkey_21_, pkey_177_, pkey_186_, pkey_191_, 
	pkey_11_, pkey_20_, pkey_178_, pkey_185_, pkey_192_, pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, 
	pksi_102_, pksi_115_, pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_, pksi_82_, pksi_95_, pksi_101_, 
	pksi_116_, pksi_127_, pksi_52_, pksi_63_, pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_, 
	pksi_62_, pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_, pksi_65_, pksi_76_, pksi_87_, 
	pksi_90_, pksi_119_, pksi_124_, pksi_191_, pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_, 
	pksi_56_, pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_, pksi_57_, pksi_66_, pksi_75_, 
	pksi_84_, pksi_93_, pksi_118_, pksi_125_, pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, 
	pksi_15_, pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_, pksi_27_, pksi_34_, pksi_45_, 
	pksi_108_, pksi_122_, pksi_17_, pksi_26_, pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, 
	pksi_32_, pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_, pksi_33_, pksi_42_, pksi_105_, 
	pksi_112_, pksi_12_, pksi_23_, pksi_30_, pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_, 
	pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_, pksi_164_, pksi_177_, pksi_2_, pksi_152_, 
	pksi_163_, pksi_178_, pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_, pksi_150_, pksi_165_, 
	pksi_187_, pksi_18_, pksi_29_, pksi_142_, pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_, 
	pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_, pksi_131_, pksi_140_, pksi_175_, pksi_184_, 
	pksi_39_, pksi_48_, pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_, pksi_133_, pksi_146_, 
	pksi_159_, pksi_182_, pksi_59_, pksi_68_, pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_, 
	pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_, pksi_8_, pksi_79_, pksi_88_, pksi_136_, 
	pksi_143_, pksi_158_, pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_, pksi_99_, 
	pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_, pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, 
	pksi_154_, pksi_161_);

input pcount_3_;
input pkey_5_;
input pkey_131_;
input pkey_144_;
input pkey_157_;
input pkey_230_;
input pkey_243_;
input pcount_2_;
input pkey_4_;
input pkey_132_;
input pkey_143_;
input pkey_158_;
input pkey_169_;
input pkey_231_;
input pkey_242_;
input pcount_1_;
input pkey_7_;
input pkey_146_;
input pkey_159_;
input pkey_168_;
input pkey_245_;
input pcount_0_;
input pkey_6_;
input pkey_130_;
input pkey_145_;
input pkey_167_;
input pkey_244_;
input pkey_9_;
input pkey_16_;
input pkey_27_;
input pkey_38_;
input pkey_49_;
input pkey_122_;
input pkey_148_;
input pkey_153_;
input pkey_166_;
input pkey_221_;
input pkey_247_;
input pkey_252_;
input pkey_8_;
input pkey_17_;
input pkey_26_;
input pkey_39_;
input pkey_48_;
input pkey_110_;
input pkey_121_;
input pkey_147_;
input pkey_154_;
input pkey_165_;
input pkey_220_;
input pkey_246_;
input pkey_253_;
input pkey_18_;
input pkey_29_;
input pkey_36_;
input pkey_47_;
input pkey_111_;
input pkey_120_;
input pkey_155_;
input pkey_164_;
input pkey_210_;
input pkey_249_;
input pkey_254_;
input pkey_19_;
input pkey_28_;
input pkey_37_;
input pkey_46_;
input pkey_112_;
input pkey_149_;
input pkey_156_;
input pkey_163_;
input pkey_211_;
input pkey_248_;
input pkey_255_;
input pkey_56_;
input pkey_67_;
input pkey_78_;
input pkey_89_;
input pkey_113_;
input pkey_126_;
input pkey_139_;
input pkey_162_;
input pkey_212_;
input pkey_225_;
input pkey_238_;
input pkey_57_;
input pkey_66_;
input pkey_79_;
input pkey_88_;
input pkey_114_;
input pkey_125_;
input pkey_150_;
input pkey_161_;
input pkey_213_;
input pkey_224_;
input pkey_239_;
input pkey_58_;
input pkey_69_;
input pkey_76_;
input pkey_87_;
input pkey_115_;
input pkey_124_;
input pkey_137_;
input pkey_151_;
input pkey_160_;
input pkey_214_;
input pkey_223_;
input pkey_236_;
input pkey_250_;
input pkey_59_;
input pkey_68_;
input pkey_77_;
input pkey_86_;
input pkey_116_;
input pkey_123_;
input pkey_138_;
input pkey_152_;
input pkey_215_;
input pkey_222_;
input pkey_237_;
input pkey_251_;
input pkey_1_;
input pkey_96_;
input pkey_117_;
input pkey_135_;
input pkey_140_;
input pkey_216_;
input pkey_229_;
input pkey_234_;
input pkey_0_;
input pkey_97_;
input pkey_118_;
input pkey_129_;
input pkey_136_;
input pkey_217_;
input pkey_228_;
input pkey_235_;
input pkey_3_;
input pkey_98_;
input pkey_119_;
input pkey_128_;
input pkey_133_;
input pkey_142_;
input pkey_218_;
input pkey_227_;
input pkey_232_;
input pkey_241_;
input pkey_2_;
input pkey_99_;
input pkey_127_;
input pkey_134_;
input pkey_141_;
input pkey_219_;
input pkey_226_;
input pkey_233_;
input pkey_240_;
input pkey_70_;
input pkey_81_;
input pkey_92_;
input pkey_108_;
input pkey_180_;
input pkey_193_;
input pkey_207_;
input pkey_71_;
input pkey_80_;
input pkey_93_;
input pkey_107_;
input pkey_194_;
input pkey_206_;
input pclk;
input pkey_50_;
input pkey_61_;
input pkey_94_;
input pkey_182_;
input pkey_195_;
input pkey_209_;
input pstart_0_;
input pkey_51_;
input pkey_60_;
input pkey_95_;
input pkey_109_;
input pkey_181_;
input pkey_196_;
input pkey_208_;
input pkey_52_;
input pkey_63_;
input pkey_74_;
input pkey_85_;
input pkey_104_;
input pkey_171_;
input pkey_197_;
input pkey_203_;
input pencrypt_0_;
input pkey_53_;
input pkey_62_;
input pkey_75_;
input pkey_84_;
input pkey_103_;
input pkey_172_;
input pkey_198_;
input pkey_202_;
input pkey_54_;
input pkey_65_;
input pkey_72_;
input pkey_83_;
input pkey_90_;
input pkey_106_;
input pkey_199_;
input pkey_205_;
input pkey_55_;
input pkey_64_;
input pkey_73_;
input pkey_82_;
input pkey_91_;
input pkey_105_;
input pkey_170_;
input pkey_204_;
input pkey_12_;
input pkey_23_;
input pkey_34_;
input pkey_45_;
input pkey_100_;
input pkey_175_;
input pkey_188_;
input pkey_13_;
input pkey_22_;
input pkey_35_;
input pkey_44_;
input pkey_176_;
input pkey_187_;
input pkey_14_;
input pkey_25_;
input pkey_32_;
input pkey_43_;
input pkey_102_;
input pkey_173_;
input pkey_201_;
input pkey_15_;
input pkey_24_;
input pkey_33_;
input pkey_42_;
input pkey_101_;
input pkey_174_;
input pkey_189_;
input pkey_200_;
input pkey_30_;
input pkey_41_;
input pkey_179_;
input pkey_184_;
input pkey_31_;
input pkey_40_;
input pkey_183_;
input pkey_190_;
input pkey_10_;
input pkey_21_;
input pkey_177_;
input pkey_186_;
input pkey_191_;
input pkey_11_;
input pkey_20_;
input pkey_178_;
input pkey_185_;
input pkey_192_;
output pksi_50_;
output pksi_61_;
output pksi_72_;
output pksi_83_;
output pksi_94_;
output pksi_102_;
output pksi_115_;
output pksi_128_;
output pdata_ready_0_;
output pksi_51_;
output pksi_60_;
output pksi_73_;
output pksi_82_;
output pksi_95_;
output pksi_101_;
output pksi_116_;
output pksi_127_;
output pksi_52_;
output pksi_63_;
output pksi_70_;
output pksi_81_;
output pksi_96_;
output pksi_100_;
output pksi_113_;
output pksi_53_;
output pksi_62_;
output pksi_71_;
output pksi_80_;
output pksi_97_;
output pksi_114_;
output pksi_129_;
output pksi_54_;
output pksi_65_;
output pksi_76_;
output pksi_87_;
output pksi_90_;
output pksi_119_;
output pksi_124_;
output pksi_191_;
output pksi_55_;
output pksi_64_;
output pksi_77_;
output pksi_86_;
output pksi_91_;
output pksi_123_;
output pksi_56_;
output pksi_67_;
output pksi_74_;
output pksi_85_;
output pksi_92_;
output pksi_117_;
output pksi_126_;
output pksi_57_;
output pksi_66_;
output pksi_75_;
output pksi_84_;
output pksi_93_;
output pksi_118_;
output pksi_125_;
output pksi_190_;
output pksi_14_;
output pksi_25_;
output pksi_36_;
output pksi_47_;
output pksi_120_;
output pksi_15_;
output pksi_24_;
output pksi_37_;
output pksi_46_;
output pksi_109_;
output pnew_count_3_;
output pksi_16_;
output pksi_27_;
output pksi_34_;
output pksi_45_;
output pksi_108_;
output pksi_122_;
output pksi_17_;
output pksi_26_;
output pksi_35_;
output pksi_44_;
output pksi_107_;
output pksi_121_;
output pksi_10_;
output pksi_21_;
output pksi_32_;
output pksi_43_;
output pksi_106_;
output pksi_111_;
output pnew_count_0_;
output pksi_11_;
output pksi_20_;
output pksi_33_;
output pksi_42_;
output pksi_105_;
output pksi_112_;
output pksi_12_;
output pksi_23_;
output pksi_30_;
output pksi_41_;
output pksi_104_;
output pnew_count_2_;
output pksi_13_;
output pksi_22_;
output pksi_31_;
output pksi_40_;
output pksi_103_;
output pksi_110_;
output pnew_count_1_;
output pksi_3_;
output pksi_151_;
output pksi_164_;
output pksi_177_;
output pksi_2_;
output pksi_152_;
output pksi_163_;
output pksi_178_;
output pksi_189_;
output pksi_1_;
output pksi_166_;
output pksi_179_;
output pksi_188_;
output pksi_0_;
output pksi_150_;
output pksi_165_;
output pksi_187_;
output pksi_18_;
output pksi_29_;
output pksi_142_;
output pksi_168_;
output pksi_173_;
output pksi_186_;
output pksi_19_;
output pksi_28_;
output pksi_130_;
output pksi_141_;
output pksi_167_;
output pksi_174_;
output pksi_185_;
output pksi_38_;
output pksi_49_;
output pksi_131_;
output pksi_140_;
output pksi_175_;
output pksi_184_;
output pksi_39_;
output pksi_48_;
output pksi_132_;
output pksi_169_;
output pksi_176_;
output pksi_183_;
output pksi_58_;
output pksi_69_;
output pksi_133_;
output pksi_146_;
output pksi_159_;
output pksi_182_;
output pksi_59_;
output pksi_68_;
output pksi_134_;
output pksi_145_;
output pksi_170_;
output pksi_181_;
output pksi_9_;
output pksi_78_;
output pksi_89_;
output pksi_135_;
output pksi_144_;
output pksi_157_;
output pksi_171_;
output pksi_180_;
output pksi_8_;
output pksi_79_;
output pksi_88_;
output pksi_136_;
output pksi_143_;
output pksi_158_;
output pksi_172_;
output pksi_7_;
output pksi_98_;
output pksi_137_;
output pksi_155_;
output pksi_160_;
output pksi_6_;
output pksi_99_;
output pksi_138_;
output pksi_149_;
output pksi_156_;
output pksi_5_;
output pksi_139_;
output pksi_148_;
output pksi_153_;
output pksi_162_;
output pksi_4_;
output pksi_147_;
output pksi_154_;
output pksi_161_;
wire n_n2854;
wire n_n2866;
wire n_n2878;
wire n_n2893;
wire n_n2905;
wire n_n2918;
wire n_n2969;
wire n_n2981;
wire n_n2855;
wire n_n2864;
wire n_n2880;
wire n_n2892;
wire n_n2906;
wire n_n2916;
wire n_n2970;
wire n_n2980;
wire n_n2856;
wire n_n2868;
wire n_n2875;
wire n_n2891;
wire n_n2928;
wire n_n2940;
wire n_n2971;
wire n_n2984;
wire n_n2992;
wire n_n2857;
wire n_n2867;
wire n_n2876;
wire n_n2890;
wire n_n2929;
wire n_n2939;
wire n_n2972;
wire n_n2983;
wire n_n2744;
wire n_n2849;
wire n_n2861;
wire n_n2873;
wire n_n2888;
wire n_n2952;
wire n_n2965;
wire n_n2977;
wire n_n2990;
wire n_n2850;
wire n_n2860;
wire n_n2874;
wire n_n2887;
wire n_n2953;
wire n_n2963;
wire n_n2966;
wire n_n2991;
wire n_n2851;
wire n_n2863;
wire n_n2871;
wire n_n2886;
wire n_n2967;
wire n_n2979;
wire n_n2852;
wire n_n2862;
wire n_n2872;
wire n_n2884;
wire n_n2968;
wire n_n2978;
wire n_n2989;
wire n_n2739;
wire n_n2896;
wire n_n2908;
wire n_n2922;
wire n_n2934;
wire n_n2947;
wire n_n2960;
wire n_n2740;
wire n_n2897;
wire n_n2907;
wire n_n2923;
wire n_n2933;
wire n_n2948;
wire n_n2959;
wire n_n2742;
wire n_n2898;
wire n_n2911;
wire n_n2919;
wire n_n2932;
wire n_n2949;
wire n_n2962;
wire n_n2743;
wire n_n2900;
wire n_n2910;
wire n_n2920;
wire n_n2930;
wire n_n2951;
wire n_n2961;
wire n_n2734;
wire n_n2858;
wire n_n2870;
wire n_n2901;
wire n_n2913;
wire n_n2926;
wire n_n2938;
wire n_n2941;
wire n_n2956;
wire n_n2973;
wire n_n2987;
wire n_n2735;
wire n_n2859;
wire n_n2869;
wire n_n2902;
wire n_n2912;
wire n_n2927;
wire n_n2937;
wire n_n2942;
wire n_n2955;
wire n_n2974;
wire n_n2985;
wire n_n2736;
wire n_n2882;
wire n_n2895;
wire n_n2903;
wire n_n2915;
wire n_n2924;
wire n_n2936;
wire n_n2944;
wire n_n2958;
wire n_n2975;
wire n_n2738;
wire n_n2883;
wire n_n2894;
wire n_n2904;
wire n_n2914;
wire n_n2925;
wire n_n2935;
wire n_n2946;
wire n_n2957;
wire n_n2988;
wire n_n2792;
wire n_n2804;
wire n_n2817;
wire n_n2829;
wire n_n2842;
wire n_n2793;
wire n_n2803;
wire n_n2818;
wire n_n2828;
wire n_n2844;
wire n_n2794;
wire n_n2807;
wire n_n2815;
wire n_n2827;
wire n_n2845;
wire n_n2733;
wire n_n2795;
wire n_n2805;
wire n_n2816;
wire n_n2826;
wire n_n2846;
wire n_n2745;
wire n_n2759;
wire n_n2771;
wire n_n2784;
wire n_n2847;
wire n_n2747;
wire n_n2758;
wire n_n2772;
wire n_n2783;
wire n_n2848;
wire n_n2748;
wire n_n2761;
wire n_n2768;
wire n_n2782;
wire n_n2750;
wire n_n2760;
wire n_n2769;
wire n_n2781;
wire n_n2751;
wire n_n2763;
wire n_n2776;
wire n_n2788;
wire n_n2800;
wire n_n2814;
wire n_n2752;
wire n_n2762;
wire n_n2777;
wire n_n2787;
wire n_n2801;
wire n_n2813;
wire n_n2753;
wire n_n2765;
wire n_n2773;
wire n_n2786;
wire n_n2824;
wire n_n2836;
wire n_n2754;
wire n_n2764;
wire n_n2775;
wire n_n2785;
wire n_n2825;
wire n_n2835;
wire n_n2755;
wire n_n2767;
wire n_n2796;
wire n_n2809;
wire n_n2822;
wire n_n2833;
wire n_n2837;
wire n_n2756;
wire n_n2766;
wire n_n2797;
wire n_n2808;
wire n_n2823;
wire n_n2832;
wire n_n2839;
wire n_n2778;
wire n_n2791;
wire n_n2798;
wire n_n2812;
wire n_n2819;
wire n_n2831;
wire n_n2840;
wire n_n2780;
wire n_n2790;
wire n_n2799;
wire n_n2810;
wire n_n2820;
wire n_n2830;
wire n_n2841;
wire wire891;
wire wire894;
wire wire775;
wire wire776;
wire wire777;
wire wire778;
wire wire779;
wire wire780;
wire wire781;
wire wire782;
wire wire783;
wire wire887;
wire wire890;
wire n_n2997;
wire wire774;
wire n_n2993;
wire wire784;
wire wire785;
wire wire786;
wire wire787;
wire wire788;
wire wire789;
wire wire790;
wire wire791;
wire wire792;
wire wire793;
wire wire794;
wire wire795;
wire wire796;
wire wire797;
wire wire798;
wire wire799;
wire wire800;
wire wire801;
wire wire802;
wire wire803;
wire wire804;
wire wire805;
wire wire806;
wire wire807;
wire wire808;
wire wire809;
wire wire810;
wire wire811;
wire wire812;
wire wire813;
wire wire814;
wire wire815;
wire wire816;
wire wire817;
wire wire818;
wire wire819;
wire wire820;
wire wire821;
wire wire822;
wire wire823;
wire wire824;
wire wire825;
wire wire826;
wire wire827;
wire wire828;
wire wire829;
wire wire830;
wire wire831;
wire wire832;
wire wire833;
wire wire834;
wire wire835;
wire wire836;
wire wire837;
wire wire838;
wire wire839;
wire wire840;
wire wire841;
wire wire842;
wire wire843;
wire wire844;
wire wire845;
wire wire846;
wire wire847;
wire wire848;
wire wire849;
wire wire850;
wire wire851;
wire wire852;
wire wire853;
wire wire854;
wire wire855;
wire wire856;
wire wire857;
wire wire858;
wire wire859;
wire wire860;
wire wire861;
wire wire862;
wire wire863;
wire wire864;
wire wire865;
wire wire866;
wire wire867;
wire wire868;
wire wire869;
wire wire870;
wire wire871;
wire wire872;
wire wire873;
wire wire874;
wire wire875;
wire wire876;
wire wire877;
wire wire878;
wire wire879;
wire wire880;
wire wire881;
wire wire882;
wire wire883;
wire wire884;
wire wire885;
wire wire886;
wire wire893;
wire wire907;
wire wire917;
wire wire919;
wire wire920;
wire wire923;
wire wire925;
wire wire926;
wire wire929;
wire wire931;
wire wire932;
wire wire935;
wire wire937;
wire wire938;
wire wire941;
wire wire943;
wire wire944;
wire wire947;
wire wire949;
wire wire950;
wire wire953;
wire wire955;
wire wire956;
wire wire959;
wire wire961;
wire wire962;
wire wire965;
wire wire967;
wire wire968;
wire wire971;
wire wire973;
wire wire974;
wire wire977;
wire wire979;
wire wire980;
wire wire983;
wire wire985;
wire wire986;
wire wire989;
wire wire991;
wire wire992;
wire wire995;
wire wire997;
wire wire998;
wire wire1001;
wire wire1003;
wire wire1004;
wire wire1007;
wire wire1009;
wire wire1010;
wire wire1013;
wire wire1015;
wire wire1016;
wire wire1019;
wire wire1021;
wire wire1022;
wire wire1025;
wire wire1027;
wire wire1028;
wire wire1031;
wire wire1033;
wire wire1034;
wire wire1037;
wire wire1039;
wire wire1040;
wire wire1043;
wire wire1045;
wire wire1046;
wire wire1049;
wire wire1051;
wire wire1052;
wire wire1055;
wire wire1057;
wire wire1058;
wire wire1061;
wire wire1063;
wire wire1064;
wire wire1067;
wire wire1069;
wire wire1070;
wire wire1073;
wire wire1075;
wire wire1076;
wire wire1079;
wire wire1081;
wire wire1082;
wire wire1085;
wire wire1087;
wire wire1088;
wire wire1091;
wire wire1093;
wire wire1094;
wire wire1097;
wire wire1099;
wire wire1100;
wire wire1103;
wire wire1105;
wire wire1106;
wire wire1109;
wire wire1111;
wire wire1112;
wire wire1115;
wire wire1117;
wire wire1118;
wire wire1121;
wire wire1123;
wire wire1124;
wire wire1127;
wire wire1129;
wire wire1130;
wire wire1133;
wire wire1135;
wire wire1136;
wire wire1139;
wire wire1141;
wire wire1142;
wire wire1145;
wire wire1147;
wire wire1148;
wire wire1151;
wire wire1153;
wire wire1154;
wire wire1157;
wire wire1159;
wire wire1160;
wire wire1163;
wire wire1165;
wire wire1166;
wire wire1169;
wire wire1171;
wire wire1172;
wire wire1175;
wire wire1177;
wire wire1178;
wire wire1181;
wire wire1183;
wire wire1184;
wire wire1187;
wire wire1189;
wire wire1190;
wire wire1193;
wire wire1195;
wire wire1196;
wire wire1199;
wire wire1201;
wire wire1202;
wire wire1205;
wire wire1207;
wire wire1208;
wire wire1211;
wire wire1213;
wire wire1214;
wire wire1217;
wire wire1219;
wire wire1220;
wire wire1223;
wire wire1225;
wire wire1226;
wire wire1229;
wire wire1231;
wire wire1232;
wire wire1235;
wire wire1237;
wire wire1238;
wire wire1241;
wire wire1243;
wire wire1244;
wire wire1247;
wire wire1249;
wire wire1250;
wire wire1253;
wire wire1255;
wire wire1256;
wire wire1259;
wire wire1261;
wire wire1262;
wire wire1265;
wire wire1267;
wire wire1268;
wire wire1271;
wire wire1273;
wire wire1274;
wire wire1277;
wire wire1279;
wire wire1280;
wire wire1283;
wire wire1285;
wire wire1286;
wire wire1289;
wire wire1291;
wire wire1292;
wire wire1295;
wire wire1297;
wire wire1298;
wire wire1301;
wire wire1303;
wire wire1304;
wire wire1307;
wire wire1309;
wire wire1310;
wire wire1313;
wire wire1315;
wire wire1316;
wire wire1319;
wire wire1321;
wire wire1322;
wire wire1325;
wire wire1327;
wire wire1328;
wire wire1331;
wire wire1333;
wire wire1334;
wire wire1337;
wire wire1339;
wire wire1340;
wire wire1343;
wire wire1345;
wire wire1346;
wire wire1349;
wire wire1351;
wire wire1352;
wire wire1355;
wire wire1357;
wire wire1358;
wire wire1361;
wire wire1363;
wire wire1364;
wire wire1367;
wire wire1369;
wire wire1370;
wire wire1373;
wire wire1375;
wire wire1376;
wire wire1379;
wire wire1381;
wire wire1382;
wire wire1385;
wire wire1387;
wire wire1388;
wire wire1391;
wire wire1393;
wire wire1394;
wire wire1397;
wire wire1399;
wire wire1400;
wire wire1403;
wire wire1405;
wire wire1406;
wire wire1409;
wire wire1411;
wire wire1412;
wire wire1415;
wire wire1417;
wire wire1418;
wire wire1421;
wire wire1423;
wire wire1424;
wire wire1427;
wire wire1429;
wire wire1430;
wire wire1433;
wire wire1435;
wire wire1436;
wire wire1439;
wire wire1441;
wire wire1442;
wire wire1445;
wire wire1447;
wire wire1448;
wire wire1451;
wire wire1453;
wire wire1454;
wire wire1457;
wire wire1459;
wire wire1460;
wire wire1463;
wire wire1465;
wire wire1466;
wire wire1469;
wire wire1471;
wire wire1472;
wire wire1477;
wire wire1479;
wire wire1480;
wire wire1485;
wire wire1487;
wire wire1488;
wire wire1493;
wire wire1495;
wire wire1496;
wire wire1501;
wire wire1503;
wire wire1504;
wire wire1509;
wire wire1511;
wire wire1512;
wire wire1517;
wire wire1519;
wire wire1520;
wire wire1525;
wire wire1527;
wire wire1528;
wire wire1533;
wire wire1535;
wire wire1536;
wire wire1539;
wire wire1541;
wire wire1542;
wire wire1547;
wire wire1549;
wire wire1550;
wire wire1555;
wire wire1557;
wire wire1558;
wire wire1563;
wire wire1565;
wire wire1566;
wire wire1571;
wire wire1573;
wire wire1574;
wire wire1579;
wire wire1581;
wire wire1582;
wire wire1587;
wire wire1589;
wire wire1590;
wire wire1595;
wire wire1597;
wire wire1598;
wire wire1603;
wire wire1605;
wire wire1606;
wire wire1611;
wire wire1613;
wire wire1614;
wire wire1617;
wire wire1619;
wire wire1620;
wire wire1623;
wire wire1625;
wire wire1626;
wire wire1631;
wire wire1633;
wire wire1634;
wire wire1639;
wire wire1641;
wire wire1642;
wire wire1647;
wire wire1649;
wire wire1650;
wire wire1655;
wire wire1657;
wire wire1658;
wire wire1663;
wire wire1665;
wire wire1666;
wire wire1671;
wire wire1673;
wire wire1674;
wire wire1679;
wire wire1681;
wire wire1682;
wire wire1685;
wire wire1687;
wire wire1688;
wire wire1691;
wire wire1693;
wire wire1694;
wire wire1697;
wire wire1699;
wire wire1700;
wire wire1703;
wire wire1705;
wire wire1706;
wire wire1711;
wire wire1713;
wire wire1714;
wire wire1719;
wire wire1721;
wire wire1722;
wire wire1727;
wire wire1729;
wire wire1730;
wire wire1735;
wire wire1737;
wire wire1738;
wire wire1743;
wire wire1745;
wire wire1746;
wire wire1751;
wire wire1753;
wire wire1754;
wire wire1759;
wire wire1761;
wire wire1762;
wire wire1765;
wire wire1767;
wire wire1768;
wire wire1771;
wire wire1773;
wire wire1774;
wire wire1777;
wire wire1779;
wire wire1780;
wire wire1785;
wire wire1787;
wire wire1788;
wire wire1793;
wire wire1795;
wire wire1796;
wire wire1801;
wire wire1803;
wire wire1804;
wire wire1809;
wire wire1811;
wire wire1812;
wire wire1817;
wire wire1819;
wire wire1820;
wire wire1825;
wire wire1827;
wire wire1828;
wire wire1831;
wire wire1833;
wire wire1834;
wire wire1839;
wire wire1841;
wire wire1842;
wire wire1847;
wire wire1849;
wire wire1850;
wire wire1855;
wire wire1857;
wire wire1858;
wire wire1863;
wire wire1865;
wire wire1866;
wire wire1871;
wire wire1873;
wire wire1874;
wire wire1879;
wire wire1881;
wire wire1882;
wire wire1887;
wire wire1889;
wire wire1890;
wire wire1895;
wire wire1897;
wire wire1898;
wire wire1903;
wire wire1905;
wire wire1906;
wire wire1911;
wire wire1913;
wire wire1914;
wire wire1919;
wire wire1921;
wire wire1922;
wire wire1927;
wire wire1929;
wire wire1930;
wire wire1935;
wire wire1937;
wire wire1938;
wire wire1943;
wire wire1945;
wire wire1946;
wire wire1951;
wire wire1953;
wire wire1954;
wire wire1959;
wire wire1961;
wire wire1962;
wire wire1967;
wire wire1969;
wire wire1970;
wire wire1975;
wire wire1977;
wire wire1978;
wire wire1983;
wire wire1985;
wire wire1986;
wire wire1991;
wire wire1993;
wire wire1994;
wire wire1997;
wire wire1999;
wire wire2000;
wire wire2005;
wire wire2007;
wire wire2008;
wire wire2013;
wire wire2015;
wire wire2016;
wire wire2021;
wire wire2023;
wire wire2024;
wire wire2029;
wire wire2031;
wire wire2032;
wire wire2035;
wire wire2037;
wire wire2038;
wire wire2043;
wire wire2045;
wire wire2046;
wire wire2049;
wire wire2051;
wire wire2052;
wire wire2055;
wire wire2057;
wire wire2058;
wire wire2063;
wire wire2065;
wire wire2066;
wire wire2071;
wire wire2073;
wire wire2074;
wire wire2079;
wire wire2081;
wire wire2082;
wire wire2087;
wire wire2089;
wire wire2090;
wire wire2093;
wire wire2095;
wire wire2096;
wire wire2099;
wire wire2101;
wire wire2102;
wire wire2107;
wire wire2109;
wire wire2110;
wire wire2115;
wire wire2117;
wire wire2118;
wire wire2123;
wire wire2125;
wire wire2126;
wire wire2131;
wire wire2133;
wire wire2134;
wire wire2139;
wire wire2141;
wire wire2142;
wire wire2147;
wire wire2149;
wire wire2150;
wire wire2153;
wire wire2155;
wire wire2156;
wire wire2161;
wire wire2163;
wire wire2164;
wire wire2169;
wire wire2171;
wire wire2172;
wire wire2177;
wire wire2179;
wire wire2180;
wire wire2185;
wire wire2187;
wire wire2188;
wire wire2193;
wire wire2195;
wire wire2196;
wire wire2201;
wire wire2203;
wire wire2204;
wire wire2207;
wire wire2209;
wire wire2210;
wire wire2215;
wire wire2217;
wire wire2218;
wire wire2223;
wire wire2225;
wire wire2226;
wire wire2231;
wire wire2233;
wire wire2234;
wire wire2239;
wire wire2241;
wire wire2242;
wire wire2247;
wire wire2249;
wire wire2250;
wire wire2255;
wire wire2257;
wire wire2258;
wire wire2263;
wire wire2265;
wire wire2266;
wire wire2271;
wire wire2273;
wire wire2274;
wire wire2279;
wire wire2281;
wire wire2282;
wire wire2287;
wire wire2289;
wire wire2290;
wire wire2295;
wire wire2297;
wire wire2298;
wire wire2301;
wire wire2303;
wire wire2304;
wire wire2309;
wire wire2311;
wire wire2312;
wire wire2317;
wire wire2319;
wire wire2320;
wire wire2325;
wire wire2327;
wire wire2328;
wire wire2333;
wire wire2335;
wire wire2336;
wire wire2341;
wire wire2343;
wire wire2344;
wire wire2349;
wire wire2351;
wire wire2352;
wire wire2357;
wire wire2359;
wire wire2360;
wire wire2365;
wire wire2367;
wire wire2368;
wire wire2373;
wire wire2375;
wire wire2376;
wire wire2381;
wire wire2383;
wire wire2384;
wire wire2389;
wire wire2391;
wire wire2392;
wire wire2397;
wire wire2399;
wire wire2400;
wire wire2405;
wire wire2407;
wire wire2408;
wire wire2413;
wire wire2415;
wire wire2416;
wire wire2421;
wire wire2423;
wire wire2424;
wire wire2429;
wire wire2431;
wire wire2432;
wire wire2437;
wire wire2439;
wire wire2440;
wire wire2445;
wire wire2447;
wire wire2448;
wire wire2453;
wire wire2455;
wire wire2456;
wire wire2461;
wire wire2463;
wire wire2464;
wire wire2469;
wire wire2471;
wire wire2472;
wire wire2477;
wire wire2479;
wire wire2480;
wire wire7760;
wire wire7763;
wire wire7764;
wire wire7765;
wire wire7766;
wire wire7767;
wire wire7770;
wire wire7771;
wire wire7772;
wire wire7773;
wire wire7776;
wire wire7777;
wire wire7778;
wire wire7781;
wire wire7782;
wire wire7783;
wire wire7786;
wire wire7787;
wire wire7788;
wire wire7791;
wire wire7792;
wire wire7793;
wire wire7796;
wire wire7797;
wire wire7798;
wire wire7801;
wire wire7802;
wire wire7803;
wire wire7806;
wire wire7807;
wire wire7808;
wire wire7811;
wire wire7812;
wire wire7813;
wire wire7816;
wire wire7817;
wire wire7818;
wire wire7821;
wire wire7822;
wire wire7823;
wire wire7826;
wire wire7827;
wire wire7828;
wire wire7831;
wire wire7832;
wire wire7833;
wire wire7836;
wire wire7837;
wire wire7838;
wire wire7841;
wire wire7842;
wire wire7843;
wire wire7846;
wire wire7847;
wire wire7848;
wire wire7851;
wire wire7852;
wire wire7853;
wire wire7856;
wire wire7857;
wire wire7858;
wire wire7861;
wire wire7862;
wire wire7863;
wire wire7866;
wire wire7867;
wire wire7868;
wire wire7871;
wire wire7872;
wire wire7873;
wire wire7876;
wire wire7877;
wire wire7878;
wire wire7881;
wire wire7882;
wire wire7883;
wire wire7886;
wire wire7887;
wire wire7888;
wire wire7891;
wire wire7892;
wire wire7893;
wire wire7896;
wire wire7897;
wire wire7898;
wire wire7901;
wire wire7902;
wire wire7903;
wire wire7906;
wire wire7907;
wire wire7908;
wire wire7911;
wire wire7912;
wire wire7913;
wire wire7916;
wire wire7917;
wire wire7918;
wire wire7921;
wire wire7922;
wire wire7923;
wire wire7926;
wire wire7927;
wire wire7928;
wire wire7931;
wire wire7932;
wire wire7933;
wire wire7936;
wire wire7937;
wire wire7938;
wire wire7941;
wire wire7942;
wire wire7943;
wire wire7946;
wire wire7947;
wire wire7948;
wire wire7951;
wire wire7952;
wire wire7953;
wire wire7956;
wire wire7957;
wire wire7958;
wire wire7961;
wire wire7962;
wire wire7963;
wire wire7966;
wire wire7967;
wire wire7968;
wire wire7971;
wire wire7972;
wire wire7973;
wire wire7976;
wire wire7977;
wire wire7978;
wire wire7981;
wire wire7982;
wire wire7983;
wire wire7986;
wire wire7987;
wire wire7988;
wire wire7991;
wire wire7992;
wire wire7993;
wire wire7996;
wire wire7997;
wire wire7998;
wire wire8001;
wire wire8002;
wire wire8003;
wire wire8006;
wire wire8007;
wire wire8008;
wire wire8011;
wire wire8012;
wire wire8013;
wire wire8016;
wire wire8017;
wire wire8018;
wire wire8021;
wire wire8022;
wire wire8023;
wire wire8026;
wire wire8027;
wire wire8028;
wire wire8031;
wire wire8032;
wire wire8033;
wire wire8036;
wire wire8037;
wire wire8038;
wire wire8041;
wire wire8042;
wire wire8043;
wire wire8046;
wire wire8047;
wire wire8048;
wire wire8051;
wire wire8052;
wire wire8053;
wire wire8056;
wire wire8057;
wire wire8058;
wire wire8061;
wire wire8062;
wire wire8063;
wire wire8066;
wire wire8067;
wire wire8068;
wire wire8071;
wire wire8072;
wire wire8073;
wire wire8076;
wire wire8077;
wire wire8078;
wire wire8081;
wire wire8082;
wire wire8083;
wire wire8086;
wire wire8087;
wire wire8088;
wire wire8091;
wire wire8092;
wire wire8093;
wire wire8096;
wire wire8097;
wire wire8098;
wire wire8101;
wire wire8102;
wire wire8103;
wire wire8106;
wire wire8107;
wire wire8108;
wire wire8111;
wire wire8112;
wire wire8113;
wire wire8116;
wire wire8117;
wire wire8118;
wire wire8121;
wire wire8122;
wire wire8123;
wire wire8126;
wire wire8127;
wire wire8128;
wire wire8131;
wire wire8132;
wire wire8133;
wire wire8136;
wire wire8137;
wire wire8138;
wire wire8141;
wire wire8142;
wire wire8143;
wire wire8146;
wire wire8147;
wire wire8148;
wire wire8151;
wire wire8152;
wire wire8153;
wire wire8156;
wire wire8157;
wire wire8158;
wire wire8161;
wire wire8162;
wire wire8163;
wire wire8166;
wire wire8167;
wire wire8168;
wire wire8171;
wire wire8172;
wire wire8173;
wire wire8176;
wire wire8177;
wire wire8178;
wire wire8181;
wire wire8182;
wire wire8183;
wire wire8186;
wire wire8187;
wire wire8188;
wire wire8191;
wire wire8192;
wire wire8193;
wire wire8196;
wire wire8197;
wire wire8198;
wire wire8201;
wire wire8202;
wire wire8203;
wire wire8206;
wire wire8207;
wire wire8208;
wire wire8211;
wire wire8212;
wire wire8213;
wire wire8216;
wire wire8217;
wire wire8218;
wire wire8221;
wire wire8222;
wire wire8223;
wire wire8226;
wire wire8227;
wire wire8228;
wire wire8231;
wire wire8232;
wire wire8233;
wire wire8236;
wire wire8237;
wire wire8238;
wire wire8241;
wire wire8242;
wire wire8243;
wire wire8246;
wire wire8247;
wire wire8248;
wire wire8251;
wire wire8252;
wire wire8253;
wire wire8256;
wire wire8257;
wire wire8258;
wire wire8261;
wire wire8262;
wire wire8263;
wire wire8266;
wire wire8267;
wire wire8268;
wire wire8271;
wire wire8272;
wire wire8273;
wire wire8276;
wire wire8277;
wire wire8278;
wire wire8281;
wire wire8282;
wire wire8283;
wire wire8286;
wire wire8287;
wire wire8288;
wire wire8291;
wire wire8292;
wire wire8293;
wire wire8296;
wire wire8297;
wire wire8298;
wire wire8301;
wire wire8302;
wire wire8303;
wire wire8306;
wire wire8307;
wire wire8308;
wire wire8311;
wire wire8312;
wire wire8313;
wire wire8316;
wire wire8317;
wire wire8318;
wire wire8321;
wire wire8322;
wire wire8323;
wire wire8326;
wire wire8327;
wire wire8328;
wire wire8331;
wire wire8332;
wire wire8333;
wire wire8336;
wire wire8337;
wire wire8338;
wire wire8341;
wire wire8342;
wire wire8343;
wire wire8346;
wire wire8347;
wire wire8348;
wire wire8351;
wire wire8352;
wire wire8353;
wire wire8356;
wire wire8357;
wire wire8358;
wire wire8361;
wire wire8362;
wire wire8363;
wire wire8366;
wire wire8367;
wire wire8368;
wire wire8371;
wire wire8372;
wire wire8373;
wire wire8376;
wire wire8377;
wire wire8378;
wire wire8381;
wire wire8382;
wire wire8383;
wire wire8386;
wire wire8387;
wire wire8388;
wire wire8391;
wire wire8392;
wire wire8393;
wire wire8396;
wire wire8397;
wire wire8398;
wire wire8401;
wire wire8402;
wire wire8403;
wire wire8406;
wire wire8407;
wire wire8408;
wire wire8411;
wire wire8412;
wire wire8413;
wire wire8416;
wire wire8417;
wire wire8418;
wire wire8421;
wire wire8422;
wire wire8423;
wire wire8426;
wire wire8427;
wire wire8428;
wire wire8431;
wire wire8432;
wire wire8433;
wire wire8436;
wire wire8437;
wire wire8438;
wire wire8441;
wire wire8442;
wire wire8443;
wire wire8446;
wire wire8447;
wire wire8448;
wire wire8451;
wire wire8452;
wire wire8453;
wire wire8456;
wire wire8457;
wire wire8458;
wire wire8461;
wire wire8462;
wire wire8463;
wire wire8466;
wire wire8467;
wire wire8468;
wire wire8471;
wire wire8472;
wire wire8473;
wire wire8476;
wire wire8477;
wire wire8478;
wire wire8481;
wire wire8482;
wire wire8483;
wire wire8486;
wire wire8487;
wire wire8488;
wire wire8491;
wire wire8492;
wire wire8493;
wire wire8496;
wire wire8497;
wire wire8498;
wire wire8501;
wire wire8502;
wire wire8503;
wire wire8506;
wire wire8507;
wire wire8508;
wire wire8511;
wire wire8512;
wire wire8513;
wire wire8516;
wire wire8517;
wire wire8518;
wire wire8521;
wire wire8522;
wire wire8523;
wire wire8526;
wire wire8527;
wire wire8528;
wire wire8531;
wire wire8532;
wire wire8533;
wire wire8536;
wire wire8537;
wire wire8538;
wire wire8541;
wire wire8542;
wire wire8543;
wire wire8546;
wire wire8547;
wire wire8548;
wire wire8551;
wire wire8552;
wire wire8553;
wire wire8556;
wire wire8557;
wire wire8558;
wire wire8561;
wire wire8562;
wire wire8563;
wire wire8566;
wire wire8567;
wire wire8568;
wire wire8571;
wire wire8572;
wire wire8573;
wire wire8576;
wire wire8577;
wire wire8578;
wire wire8581;
wire wire8582;
wire wire8583;
wire wire8586;
wire wire8587;
wire wire8588;
wire wire8591;
wire wire8592;
wire wire8593;
wire wire8596;
wire wire8597;
wire wire8598;
wire wire8601;
wire wire8602;
wire wire8603;
wire wire8606;
wire wire8607;
wire wire8608;
wire wire8611;
wire wire8612;
wire wire8613;
wire wire8616;
wire wire8617;
wire wire8618;
wire wire8621;
wire wire8622;
wire wire8623;
wire wire8626;
wire wire8627;
wire wire8628;
wire wire8631;
wire wire8632;
wire wire8633;
wire wire8636;
wire wire8637;
wire wire8638;
wire wire8641;
wire wire8642;
wire wire8643;
wire wire8646;
wire wire8647;
wire wire8648;
wire wire8651;
wire wire8652;
wire wire8653;
wire wire8656;
wire wire8657;
wire wire8658;
wire wire8661;
wire wire8662;
wire wire8663;
wire wire8666;
wire wire8667;
wire wire8668;
wire wire8671;
wire wire8672;
wire wire8673;
wire wire8676;
wire wire8677;
wire wire8678;
wire wire8681;
wire wire8682;
wire wire8683;
wire wire8686;
wire wire8687;
wire wire8688;
wire wire8691;
wire wire8692;
wire wire8693;
wire wire8696;
wire wire8697;
wire wire8698;
wire wire8701;
wire wire8702;
wire wire8703;
wire wire8706;
wire wire8707;
wire wire8708;
wire wire8711;
wire wire8712;
wire wire8713;
wire wire8716;
wire wire8717;
wire wire8718;
wire wire8721;
wire wire8722;
wire wire8723;
wire wire8726;
wire wire8727;
wire wire8728;
wire wire8731;
wire wire8732;
wire wire8733;
wire wire8736;
wire wire8737;
wire wire8738;
wire wire8741;
wire wire8742;
wire wire8743;
wire wire8746;
wire wire8747;
wire wire8748;
wire wire8751;
wire wire8752;
wire wire8753;
wire wire8756;
wire wire8757;
wire wire8758;
wire wire8761;
wire wire8762;
wire wire8763;
wire wire8766;
wire wire8767;
wire wire8768;
wire wire8771;
wire wire8772;
wire wire8773;
wire wire8776;
wire wire8777;
wire wire8778;
wire wire8781;
wire wire8782;
wire wire8783;
wire wire8786;
wire wire8787;
wire wire8788;
wire wire8791;
wire wire8792;
wire wire8793;
wire wire8796;
wire wire8797;
wire wire8798;
wire wire8801;
wire wire8802;
wire wire8803;
wire wire8806;
wire wire8807;
wire wire8808;
wire wire8811;
wire wire8812;
wire wire8813;
wire wire8816;
wire wire8817;
wire wire8818;
wire wire8821;
wire wire8822;
wire wire8823;
wire wire8826;
wire wire8827;
wire wire8828;
wire wire8831;
wire wire8832;
wire wire8833;
wire wire8836;
wire wire8837;
wire wire8838;
wire wire8841;
wire wire8842;
wire wire8843;
wire wire8846;
wire wire8847;
wire wire8848;
wire wire8851;
wire wire8852;
wire wire8853;
wire wire8856;
wire wire8857;
wire wire8858;
wire wire8861;
wire wire8862;
wire wire8863;
wire wire8866;
wire wire8867;
wire wire8868;
wire wire8871;
wire wire8872;
wire wire8873;
wire wire8876;
wire wire8877;
wire wire8878;
wire wire8881;
wire wire8882;
wire wire8883;
wire wire8889;
reg pksi_17_;

reg pksi_185_;

reg n_n2879;

reg pksi_170_;

reg pksi_155_;

reg pksi_147_;

reg pksi_109_;

reg n_n2982;

reg pksi_19_;

reg n_n2865;

reg n_n2881;

reg n_n2391;

reg pksi_148_;

reg n_n2917;

reg pksi_107_;

reg pksi_110_;

reg pksi_9_;

reg pksi_176_;

reg pksi_180_;

reg pksi_178_;

reg pksi_135_;

reg pksi_129_;

reg pksi_100_;

reg pksi_117_;

reg pksi_118_;

reg pksi_5_;

reg pksi_169_;

reg n_n2877;

reg pksi_184_;

reg pksi_125_;

reg pksi_138_;

reg pksi_114_;

reg pksi_99_;

reg pksi_85_;

reg pksi_14_;

reg pksi_4_;

reg pksi_186_;

reg n_n2889;

reg pksi_141_;

reg pksi_113_;

reg pksi_115_;

reg pksi_98_;

reg pksi_2_;

reg pksi_23_;

reg pksi_177_;

reg pksi_189_;

reg n_n2954;

reg n_n2964;

reg pksi_97_;

reg pksi_102_;

reg pksi_11_;

reg pksi_173_;

reg pksi_179_;

reg pksi_171_;

reg pksi_104_;

reg pksi_103_;

reg n_n2853;

reg pksi_183_;

reg pksi_172_;

reg n_n2885;

reg pksi_116_;

reg pksi_96_;

reg pksi_119_;

reg pksi_84_;

reg pksi_159_;

reg n_n2909;

reg pksi_160_;

reg pksi_128_;

reg pksi_127_;

reg pksi_142_;

reg n_n2741;

reg pksi_149_;

reg pksi_162_;

reg pksi_154_;

reg pksi_121_;

reg pksi_134_;

reg pksi_126_;

reg pksi_82_;

reg n_n2899;

reg pksi_153_;

reg pksi_165_;

reg pksi_137_;

reg n_n2950;

reg pksi_101_;

reg pksi_93_;

reg pksi_161_;

reg pksi_156_;

reg n_n2921;

reg n_n2931;

reg pksi_123_;

reg pksi_111_;

reg pksi_92_;

reg pksi_15_;

reg n_n2379;

reg pksi_145_;

reg pksi_144_;

reg pksi_150_;

reg pksi_124_;

reg pksi_132_;

reg pksi_130_;

reg pksi_105_;

reg pksi_112_;

reg n_n2280;

reg pksi_6_;

reg pksi_188_;

reg pksi_152_;

reg pksi_163_;

reg pksi_166_;

reg pksi_131_;

reg n_n2943;

reg pksi_136_;

reg pksi_108_;

reg n_n2986;

reg n_n2737;

reg pksi_175_;

reg pksi_190_;

reg pksi_164_;

reg pksi_158_;

reg pksi_167_;

reg pksi_133_;

reg n_n2945;

reg pksi_122_;

reg n_n2976;

reg pksi_75_;

reg pksi_182_;

reg pksi_174_;

reg pksi_157_;

reg pksi_151_;

reg pksi_146_;

reg pksi_140_;

reg pksi_120_;

reg n_n2438;

reg pksi_106_;

reg pksi_57_;

reg pksi_36_;

reg pksi_38_;

reg pksi_28_;

reg n_n2843;

reg pksi_53_;

reg pksi_27_;

reg pksi_26_;

reg pksi_47_;

reg pksi_1_;

reg pksi_63_;

reg pksi_34_;

reg pksi_24_;

reg pksi_30_;

reg pksi_18_;

reg pksi_79_;

reg pksi_54_;

reg n_n2806;

reg pksi_46_;

reg pksi_39_;

reg pksi_8_;

reg n_n2746;

reg pksi_91_;

reg pksi_51_;

reg pksi_70_;

reg pksi_0_;

reg pksi_73_;

reg pksi_89_;

reg pksi_60_;

reg pksi_48_;

reg pksi_22_;

reg n_n2749;

reg pksi_77_;

reg pksi_64_;

reg pksi_56_;

reg pksi_80_;

reg pksi_81_;

reg n_n2770;

reg pksi_66_;

reg pksi_72_;

reg pksi_78_;

reg pksi_69_;

reg n_n2789;

reg pksi_40_;

reg pksi_32_;

reg pksi_94_;

reg pksi_87_;

reg pksi_61_;

reg pksi_59_;

reg n_n2802;

reg pksi_42_;

reg pksi_86_;

reg pksi_76_;

reg n_n2774;

reg pksi_50_;

reg pksi_33_;

reg pksi_12_;

reg pksi_74_;

reg pksi_95_;

reg pksi_58_;

reg pksi_62_;

reg pksi_29_;

reg pksi_3_;

reg pksi_83_;

reg pksi_68_;

reg pksi_71_;

reg pksi_37_;

reg pksi_41_;

reg n_n2834;

reg n_n2838;

reg n_n2757;

reg pksi_55_;

reg pksi_52_;

reg pksi_45_;

reg pksi_43_;

reg pksi_16_;

reg pksi_10_;

reg n_n2779;

reg pksi_67_;

reg pksi_31_;

reg pksi_25_;

reg pksi_35_;

reg pksi_20_;

reg pksi_21_;

reg pksi_49_;

reg pksi_65_;

reg pksi_44_;

reg n_n2811;

reg n_n2821;

reg pksi_7_;

reg pksi_13_;

always  @(posedge pclk)
	pksi_17_<=n_n2854;

 always  @(posedge pclk)
	pksi_185_<=n_n2866;

 always  @(posedge pclk)
	n_n2879<=n_n2878;

 always  @(posedge pclk)
	pksi_170_<=n_n2893;

 always  @(posedge pclk)
	pksi_155_<=n_n2905;

 always  @(posedge pclk)
	pksi_147_<=n_n2918;

 always  @(posedge pclk)
	pksi_109_<=n_n2969;

 always  @(posedge pclk)
	n_n2982<=n_n2981;

 always  @(posedge pclk)
	pksi_19_<=n_n2855;

 always  @(posedge pclk)
	n_n2865<=n_n2864;

 always  @(posedge pclk)
	n_n2881<=n_n2880;

 always  @(posedge pclk)
	n_n2391<=n_n2892;

 always  @(posedge pclk)
	pksi_148_<=n_n2906;

 always  @(posedge pclk)
	n_n2917<=n_n2916;

 always  @(posedge pclk)
	pksi_107_<=n_n2970;

 always  @(posedge pclk)
	pksi_110_<=n_n2980;

 always  @(posedge pclk)
	pksi_9_<=n_n2856;

 always  @(posedge pclk)
	pksi_176_<=n_n2868;

 always  @(posedge pclk)
	pksi_180_<=n_n2875;

 always  @(posedge pclk)
	pksi_178_<=n_n2891;

 always  @(posedge pclk)
	pksi_135_<=n_n2928;

 always  @(posedge pclk)
	pksi_129_<=n_n2940;

 always  @(posedge pclk)
	pksi_100_<=n_n2971;

 always  @(posedge pclk)
	pksi_117_<=n_n2984;

 always  @(posedge pclk)
	pksi_118_<=n_n2992;

 always  @(posedge pclk)
	pksi_5_<=n_n2857;

 always  @(posedge pclk)
	pksi_169_<=n_n2867;

 always  @(posedge pclk)
	n_n2877<=n_n2876;

 always  @(posedge pclk)
	pksi_184_<=n_n2890;

 always  @(posedge pclk)
	pksi_125_<=n_n2929;

 always  @(posedge pclk)
	pksi_138_<=n_n2939;

 always  @(posedge pclk)
	pksi_114_<=n_n2972;

 always  @(posedge pclk)
	pksi_99_<=n_n2983;

 always  @(posedge pclk)
	pksi_85_<=n_n2744;

 always  @(posedge pclk)
	pksi_14_<=n_n2849;

 always  @(posedge pclk)
	pksi_4_<=n_n2861;

 always  @(posedge pclk)
	pksi_186_<=n_n2873;

 always  @(posedge pclk)
	n_n2889<=n_n2888;

 always  @(posedge pclk)
	pksi_141_<=n_n2952;

 always  @(posedge pclk)
	pksi_113_<=n_n2965;

 always  @(posedge pclk)
	pksi_115_<=n_n2977;

 always  @(posedge pclk)
	pksi_98_<=n_n2990;

 always  @(posedge pclk)
	pksi_2_<=n_n2850;

 always  @(posedge pclk)
	pksi_23_<=n_n2860;

 always  @(posedge pclk)
	pksi_177_<=n_n2874;

 always  @(posedge pclk)
	pksi_189_<=n_n2887;

 always  @(posedge pclk)
	n_n2954<=n_n2953;

 always  @(posedge pclk)
	n_n2964<=n_n2963;

 always  @(posedge pclk)
	pksi_97_<=n_n2966;

 always  @(posedge pclk)
	pksi_102_<=n_n2991;

 always  @(posedge pclk)
	pksi_11_<=n_n2851;

 always  @(posedge pclk)
	pksi_173_<=n_n2863;

 always  @(posedge pclk)
	pksi_179_<=n_n2871;

 always  @(posedge pclk)
	pksi_171_<=n_n2886;

 always  @(posedge pclk)
	pksi_104_<=n_n2967;

 always  @(posedge pclk)
	pksi_103_<=n_n2979;

 always  @(posedge pclk)
	n_n2853<=n_n2852;

 always  @(posedge pclk)
	pksi_183_<=n_n2862;

 always  @(posedge pclk)
	pksi_172_<=n_n2872;

 always  @(posedge pclk)
	n_n2885<=n_n2884;

 always  @(posedge pclk)
	pksi_116_<=n_n2968;

 always  @(posedge pclk)
	pksi_96_<=n_n2978;

 always  @(posedge pclk)
	pksi_119_<=n_n2989;

 always  @(posedge pclk)
	pksi_84_<=n_n2739;

 always  @(posedge pclk)
	pksi_159_<=n_n2896;

 always  @(posedge pclk)
	n_n2909<=n_n2908;

 always  @(posedge pclk)
	pksi_160_<=n_n2922;

 always  @(posedge pclk)
	pksi_128_<=n_n2934;

 always  @(posedge pclk)
	pksi_127_<=n_n2947;

 always  @(posedge pclk)
	pksi_142_<=n_n2960;

 always  @(posedge pclk)
	n_n2741<=n_n2740;

 always  @(posedge pclk)
	pksi_149_<=n_n2897;

 always  @(posedge pclk)
	pksi_162_<=n_n2907;

 always  @(posedge pclk)
	pksi_154_<=n_n2923;

 always  @(posedge pclk)
	pksi_121_<=n_n2933;

 always  @(posedge pclk)
	pksi_134_<=n_n2948;

 always  @(posedge pclk)
	pksi_126_<=n_n2959;

 always  @(posedge pclk)
	pksi_82_<=n_n2742;

 always  @(posedge pclk)
	n_n2899<=n_n2898;

 always  @(posedge pclk)
	pksi_153_<=n_n2911;

 always  @(posedge pclk)
	pksi_165_<=n_n2919;

 always  @(posedge pclk)
	pksi_137_<=n_n2932;

 always  @(posedge pclk)
	n_n2950<=n_n2949;

 always  @(posedge pclk)
	pksi_101_<=n_n2962;

 always  @(posedge pclk)
	pksi_93_<=n_n2743;

 always  @(posedge pclk)
	pksi_161_<=n_n2900;

 always  @(posedge pclk)
	pksi_156_<=n_n2910;

 always  @(posedge pclk)
	n_n2921<=n_n2920;

 always  @(posedge pclk)
	n_n2931<=n_n2930;

 always  @(posedge pclk)
	pksi_123_<=n_n2951;

 always  @(posedge pclk)
	pksi_111_<=n_n2961;

 always  @(posedge pclk)
	pksi_92_<=n_n2734;

 always  @(posedge pclk)
	pksi_15_<=n_n2858;

 always  @(posedge pclk)
	n_n2379<=n_n2870;

 always  @(posedge pclk)
	pksi_145_<=n_n2901;

 always  @(posedge pclk)
	pksi_144_<=n_n2913;

 always  @(posedge pclk)
	pksi_150_<=n_n2926;

 always  @(posedge pclk)
	pksi_124_<=n_n2938;

 always  @(posedge pclk)
	pksi_132_<=n_n2941;

 always  @(posedge pclk)
	pksi_130_<=n_n2956;

 always  @(posedge pclk)
	pksi_105_<=n_n2973;

 always  @(posedge pclk)
	pksi_112_<=n_n2987;

 always  @(posedge pclk)
	n_n2280<=n_n2735;

 always  @(posedge pclk)
	pksi_6_<=n_n2859;

 always  @(posedge pclk)
	pksi_188_<=n_n2869;

 always  @(posedge pclk)
	pksi_152_<=n_n2902;

 always  @(posedge pclk)
	pksi_163_<=n_n2912;

 always  @(posedge pclk)
	pksi_166_<=n_n2927;

 always  @(posedge pclk)
	pksi_131_<=n_n2937;

 always  @(posedge pclk)
	n_n2943<=n_n2942;

 always  @(posedge pclk)
	pksi_136_<=n_n2955;

 always  @(posedge pclk)
	pksi_108_<=n_n2974;

 always  @(posedge pclk)
	n_n2986<=n_n2985;

 always  @(posedge pclk)
	n_n2737<=n_n2736;

 always  @(posedge pclk)
	pksi_175_<=n_n2882;

 always  @(posedge pclk)
	pksi_190_<=n_n2895;

 always  @(posedge pclk)
	pksi_164_<=n_n2903;

 always  @(posedge pclk)
	pksi_158_<=n_n2915;

 always  @(posedge pclk)
	pksi_167_<=n_n2924;

 always  @(posedge pclk)
	pksi_133_<=n_n2936;

 always  @(posedge pclk)
	n_n2945<=n_n2944;

 always  @(posedge pclk)
	pksi_122_<=n_n2958;

 always  @(posedge pclk)
	n_n2976<=n_n2975;

 always  @(posedge pclk)
	pksi_75_<=n_n2738;

 always  @(posedge pclk)
	pksi_182_<=n_n2883;

 always  @(posedge pclk)
	pksi_174_<=n_n2894;

 always  @(posedge pclk)
	pksi_157_<=n_n2904;

 always  @(posedge pclk)
	pksi_151_<=n_n2914;

 always  @(posedge pclk)
	pksi_146_<=n_n2925;

 always  @(posedge pclk)
	pksi_140_<=n_n2935;

 always  @(posedge pclk)
	pksi_120_<=n_n2946;

 always  @(posedge pclk)
	n_n2438<=n_n2957;

 always  @(posedge pclk)
	pksi_106_<=n_n2988;

 always  @(posedge pclk)
	pksi_57_<=n_n2792;

 always  @(posedge pclk)
	pksi_36_<=n_n2804;

 always  @(posedge pclk)
	pksi_38_<=n_n2817;

 always  @(posedge pclk)
	pksi_28_<=n_n2829;

 always  @(posedge pclk)
	n_n2843<=n_n2842;

 always  @(posedge pclk)
	pksi_53_<=n_n2793;

 always  @(posedge pclk)
	pksi_27_<=n_n2803;

 always  @(posedge pclk)
	pksi_26_<=n_n2818;

 always  @(posedge pclk)
	pksi_47_<=n_n2828;

 always  @(posedge pclk)
	pksi_1_<=n_n2844;

 always  @(posedge pclk)
	pksi_63_<=n_n2794;

 always  @(posedge pclk)
	pksi_34_<=n_n2807;

 always  @(posedge pclk)
	pksi_24_<=n_n2815;

 always  @(posedge pclk)
	pksi_30_<=n_n2827;

 always  @(posedge pclk)
	pksi_18_<=n_n2845;

 always  @(posedge pclk)
	pksi_79_<=n_n2733;

 always  @(posedge pclk)
	pksi_54_<=n_n2795;

 always  @(posedge pclk)
	n_n2806<=n_n2805;

 always  @(posedge pclk)
	pksi_46_<=n_n2816;

 always  @(posedge pclk)
	pksi_39_<=n_n2826;

 always  @(posedge pclk)
	pksi_8_<=n_n2846;

 always  @(posedge pclk)
	n_n2746<=n_n2745;

 always  @(posedge pclk)
	pksi_91_<=n_n2759;

 always  @(posedge pclk)
	pksi_51_<=n_n2771;

 always  @(posedge pclk)
	pksi_70_<=n_n2784;

 always  @(posedge pclk)
	pksi_0_<=n_n2847;

 always  @(posedge pclk)
	pksi_73_<=n_n2747;

 always  @(posedge pclk)
	pksi_89_<=n_n2758;

 always  @(posedge pclk)
	pksi_60_<=n_n2772;

 always  @(posedge pclk)
	pksi_48_<=n_n2783;

 always  @(posedge pclk)
	pksi_22_<=n_n2848;

 always  @(posedge pclk)
	n_n2749<=n_n2748;

 always  @(posedge pclk)
	pksi_77_<=n_n2761;

 always  @(posedge pclk)
	pksi_64_<=n_n2768;

 always  @(posedge pclk)
	pksi_56_<=n_n2782;

 always  @(posedge pclk)
	pksi_80_<=n_n2750;

 always  @(posedge pclk)
	pksi_81_<=n_n2760;

 always  @(posedge pclk)
	n_n2770<=n_n2769;

 always  @(posedge pclk)
	pksi_66_<=n_n2781;

 always  @(posedge pclk)
	pksi_72_<=n_n2751;

 always  @(posedge pclk)
	pksi_78_<=n_n2763;

 always  @(posedge pclk)
	pksi_69_<=n_n2776;

 always  @(posedge pclk)
	n_n2789<=n_n2788;

 always  @(posedge pclk)
	pksi_40_<=n_n2800;

 always  @(posedge pclk)
	pksi_32_<=n_n2814;

 always  @(posedge pclk)
	pksi_94_<=n_n2752;

 always  @(posedge pclk)
	pksi_87_<=n_n2762;

 always  @(posedge pclk)
	pksi_61_<=n_n2777;

 always  @(posedge pclk)
	pksi_59_<=n_n2787;

 always  @(posedge pclk)
	n_n2802<=n_n2801;

 always  @(posedge pclk)
	pksi_42_<=n_n2813;

 always  @(posedge pclk)
	pksi_86_<=n_n2753;

 always  @(posedge pclk)
	pksi_76_<=n_n2765;

 always  @(posedge pclk)
	n_n2774<=n_n2773;

 always  @(posedge pclk)
	pksi_50_<=n_n2786;

 always  @(posedge pclk)
	pksi_33_<=n_n2824;

 always  @(posedge pclk)
	pksi_12_<=n_n2836;

 always  @(posedge pclk)
	pksi_74_<=n_n2754;

 always  @(posedge pclk)
	pksi_95_<=n_n2764;

 always  @(posedge pclk)
	pksi_58_<=n_n2775;

 always  @(posedge pclk)
	pksi_62_<=n_n2785;

 always  @(posedge pclk)
	pksi_29_<=n_n2825;

 always  @(posedge pclk)
	pksi_3_<=n_n2835;

 always  @(posedge pclk)
	pksi_83_<=n_n2755;

 always  @(posedge pclk)
	pksi_68_<=n_n2767;

 always  @(posedge pclk)
	pksi_71_<=n_n2796;

 always  @(posedge pclk)
	pksi_37_<=n_n2809;

 always  @(posedge pclk)
	pksi_41_<=n_n2822;

 always  @(posedge pclk)
	n_n2834<=n_n2833;

 always  @(posedge pclk)
	n_n2838<=n_n2837;

 always  @(posedge pclk)
	n_n2757<=n_n2756;

 always  @(posedge pclk)
	pksi_55_<=n_n2766;

 always  @(posedge pclk)
	pksi_52_<=n_n2797;

 always  @(posedge pclk)
	pksi_45_<=n_n2808;

 always  @(posedge pclk)
	pksi_43_<=n_n2823;

 always  @(posedge pclk)
	pksi_16_<=n_n2832;

 always  @(posedge pclk)
	pksi_10_<=n_n2839;

 always  @(posedge pclk)
	n_n2779<=n_n2778;

 always  @(posedge pclk)
	pksi_67_<=n_n2791;

 always  @(posedge pclk)
	pksi_31_<=n_n2798;

 always  @(posedge pclk)
	pksi_25_<=n_n2812;

 always  @(posedge pclk)
	pksi_35_<=n_n2819;

 always  @(posedge pclk)
	pksi_20_<=n_n2831;

 always  @(posedge pclk)
	pksi_21_<=n_n2840;

 always  @(posedge pclk)
	pksi_49_<=n_n2780;

 always  @(posedge pclk)
	pksi_65_<=n_n2790;

 always  @(posedge pclk)
	pksi_44_<=n_n2799;

 always  @(posedge pclk)
	n_n2811<=n_n2810;

 always  @(posedge pclk)
	n_n2821<=n_n2820;

 always  @(posedge pclk)
	pksi_7_<=n_n2830;

 always  @(posedge pclk)
	pksi_13_<=n_n2841;

 assign pdata_ready_0_ = ( (~ pstart_0_)  &  wire891 ) ;
 assign pnew_count_3_ = ( pstart_0_  &  (~ pencrypt_0_) ) | ( (~ pstart_0_)  &  wire907 ) | ( (~ pstart_0_)  &  wire8889 ) ;
 assign pnew_count_0_ = ( (~ pcount_0_)  &  (~ pstart_0_) ) | ( pstart_0_  &  (~ pencrypt_0_) ) ;
 assign pnew_count_2_ = ( pstart_0_  &  (~ pencrypt_0_) ) | ( (~ pstart_0_)  &  wire894 ) ;
 assign pnew_count_1_ = ( pstart_0_  &  (~ pencrypt_0_) ) | ( pcount_1_  &  pcount_0_  &  (~ pencrypt_0_) ) | ( (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) | ( (~ pcount_1_)  &  pcount_0_  &  (~ pstart_0_)  &  pencrypt_0_ ) | ( pcount_1_  &  (~ pcount_0_)  &  (~ pstart_0_)  &  pencrypt_0_ ) ;
 assign n_n2854 = ( wire2477 ) | ( wire2479 ) | ( wire2480 ) | ( wire7767 ) ;
 assign n_n2866 = ( wire2469 ) | ( wire2471 ) | ( wire2472 ) | ( wire7773 ) ;
 assign n_n2878 = ( wire2461 ) | ( wire2463 ) | ( wire2464 ) | ( wire7778 ) ;
 assign n_n2893 = ( wire2453 ) | ( wire2455 ) | ( wire2456 ) | ( wire7783 ) ;
 assign n_n2905 = ( wire2445 ) | ( wire2447 ) | ( wire2448 ) | ( wire7788 ) ;
 assign n_n2918 = ( wire2437 ) | ( wire2439 ) | ( wire2440 ) | ( wire7793 ) ;
 assign n_n2969 = ( wire2429 ) | ( wire2431 ) | ( wire2432 ) | ( wire7798 ) ;
 assign n_n2981 = ( wire2421 ) | ( wire2423 ) | ( wire2424 ) | ( wire7803 ) ;
 assign n_n2855 = ( wire2413 ) | ( wire2415 ) | ( wire2416 ) | ( wire7808 ) ;
 assign n_n2864 = ( wire2405 ) | ( wire2407 ) | ( wire2408 ) | ( wire7813 ) ;
 assign n_n2880 = ( wire2397 ) | ( wire2399 ) | ( wire2400 ) | ( wire7818 ) ;
 assign n_n2892 = ( wire2389 ) | ( wire2391 ) | ( wire2392 ) | ( wire7823 ) ;
 assign n_n2906 = ( wire2381 ) | ( wire2383 ) | ( wire2384 ) | ( wire7828 ) ;
 assign n_n2916 = ( wire2373 ) | ( wire2375 ) | ( wire2376 ) | ( wire7833 ) ;
 assign n_n2970 = ( wire2365 ) | ( wire2367 ) | ( wire2368 ) | ( wire7838 ) ;
 assign n_n2980 = ( wire2357 ) | ( wire2359 ) | ( wire2360 ) | ( wire7843 ) ;
 assign n_n2856 = ( wire2349 ) | ( wire2351 ) | ( wire2352 ) | ( wire7848 ) ;
 assign n_n2868 = ( wire2341 ) | ( wire2343 ) | ( wire2344 ) | ( wire7853 ) ;
 assign n_n2875 = ( wire2333 ) | ( wire2335 ) | ( wire2336 ) | ( wire7858 ) ;
 assign n_n2891 = ( wire2325 ) | ( wire2327 ) | ( wire2328 ) | ( wire7863 ) ;
 assign n_n2928 = ( wire2317 ) | ( wire2319 ) | ( wire2320 ) | ( wire7868 ) ;
 assign n_n2940 = ( wire2309 ) | ( wire2311 ) | ( wire2312 ) | ( wire7873 ) ;
 assign n_n2971 = ( wire2301 ) | ( wire2303 ) | ( wire2304 ) | ( wire7878 ) ;
 assign n_n2984 = ( wire2295 ) | ( wire2297 ) | ( wire2298 ) | ( wire7883 ) ;
 assign n_n2992 = ( wire2287 ) | ( wire2289 ) | ( wire2290 ) | ( wire7888 ) ;
 assign n_n2857 = ( wire2279 ) | ( wire2281 ) | ( wire2282 ) | ( wire7893 ) ;
 assign n_n2867 = ( wire2271 ) | ( wire2273 ) | ( wire2274 ) | ( wire7898 ) ;
 assign n_n2876 = ( wire2263 ) | ( wire2265 ) | ( wire2266 ) | ( wire7903 ) ;
 assign n_n2890 = ( wire2255 ) | ( wire2257 ) | ( wire2258 ) | ( wire7908 ) ;
 assign n_n2929 = ( wire2247 ) | ( wire2249 ) | ( wire2250 ) | ( wire7913 ) ;
 assign n_n2939 = ( wire2239 ) | ( wire2241 ) | ( wire2242 ) | ( wire7918 ) ;
 assign n_n2972 = ( wire2231 ) | ( wire2233 ) | ( wire2234 ) | ( wire7923 ) ;
 assign n_n2983 = ( wire2223 ) | ( wire2225 ) | ( wire2226 ) | ( wire7928 ) ;
 assign n_n2744 = ( wire2215 ) | ( wire2217 ) | ( wire2218 ) | ( wire7933 ) ;
 assign n_n2849 = ( wire2207 ) | ( wire2209 ) | ( wire2210 ) | ( wire7938 ) ;
 assign n_n2861 = ( wire2201 ) | ( wire2203 ) | ( wire2204 ) | ( wire7943 ) ;
 assign n_n2873 = ( wire2193 ) | ( wire2195 ) | ( wire2196 ) | ( wire7948 ) ;
 assign n_n2888 = ( wire2185 ) | ( wire2187 ) | ( wire2188 ) | ( wire7953 ) ;
 assign n_n2952 = ( wire2177 ) | ( wire2179 ) | ( wire2180 ) | ( wire7958 ) ;
 assign n_n2965 = ( wire2169 ) | ( wire2171 ) | ( wire2172 ) | ( wire7963 ) ;
 assign n_n2977 = ( wire2161 ) | ( wire2163 ) | ( wire2164 ) | ( wire7968 ) ;
 assign n_n2990 = ( wire2153 ) | ( wire2155 ) | ( wire2156 ) | ( wire7973 ) ;
 assign n_n2850 = ( wire2147 ) | ( wire2149 ) | ( wire2150 ) | ( wire7978 ) ;
 assign n_n2860 = ( wire2139 ) | ( wire2141 ) | ( wire2142 ) | ( wire7983 ) ;
 assign n_n2874 = ( wire2131 ) | ( wire2133 ) | ( wire2134 ) | ( wire7988 ) ;
 assign n_n2887 = ( wire2123 ) | ( wire2125 ) | ( wire2126 ) | ( wire7993 ) ;
 assign n_n2953 = ( wire2115 ) | ( wire2117 ) | ( wire2118 ) | ( wire7998 ) ;
 assign n_n2963 = ( wire2107 ) | ( wire2109 ) | ( wire2110 ) | ( wire8003 ) ;
 assign n_n2966 = ( wire2099 ) | ( wire2101 ) | ( wire2102 ) | ( wire8008 ) ;
 assign n_n2991 = ( wire2093 ) | ( wire2095 ) | ( wire2096 ) | ( wire8013 ) ;
 assign n_n2851 = ( wire2087 ) | ( wire2089 ) | ( wire2090 ) | ( wire8018 ) ;
 assign n_n2863 = ( wire2079 ) | ( wire2081 ) | ( wire2082 ) | ( wire8023 ) ;
 assign n_n2871 = ( wire2071 ) | ( wire2073 ) | ( wire2074 ) | ( wire8028 ) ;
 assign n_n2886 = ( wire2063 ) | ( wire2065 ) | ( wire2066 ) | ( wire8033 ) ;
 assign n_n2967 = ( wire2055 ) | ( wire2057 ) | ( wire2058 ) | ( wire8038 ) ;
 assign n_n2979 = ( wire2049 ) | ( wire2051 ) | ( wire2052 ) | ( wire8043 ) ;
 assign n_n2852 = ( wire2043 ) | ( wire2045 ) | ( wire2046 ) | ( wire8048 ) ;
 assign n_n2862 = ( wire2035 ) | ( wire2037 ) | ( wire2038 ) | ( wire8053 ) ;
 assign n_n2872 = ( wire2029 ) | ( wire2031 ) | ( wire2032 ) | ( wire8058 ) ;
 assign n_n2884 = ( wire2021 ) | ( wire2023 ) | ( wire2024 ) | ( wire8063 ) ;
 assign n_n2968 = ( wire2013 ) | ( wire2015 ) | ( wire2016 ) | ( wire8068 ) ;
 assign n_n2978 = ( wire2005 ) | ( wire2007 ) | ( wire2008 ) | ( wire8073 ) ;
 assign n_n2989 = ( wire1997 ) | ( wire1999 ) | ( wire2000 ) | ( wire8078 ) ;
 assign n_n2739 = ( wire1991 ) | ( wire1993 ) | ( wire1994 ) | ( wire8083 ) ;
 assign n_n2896 = ( wire1983 ) | ( wire1985 ) | ( wire1986 ) | ( wire8088 ) ;
 assign n_n2908 = ( wire1975 ) | ( wire1977 ) | ( wire1978 ) | ( wire8093 ) ;
 assign n_n2922 = ( wire1967 ) | ( wire1969 ) | ( wire1970 ) | ( wire8098 ) ;
 assign n_n2934 = ( wire1959 ) | ( wire1961 ) | ( wire1962 ) | ( wire8103 ) ;
 assign n_n2947 = ( wire1951 ) | ( wire1953 ) | ( wire1954 ) | ( wire8108 ) ;
 assign n_n2960 = ( wire1943 ) | ( wire1945 ) | ( wire1946 ) | ( wire8113 ) ;
 assign n_n2740 = ( wire1935 ) | ( wire1937 ) | ( wire1938 ) | ( wire8118 ) ;
 assign n_n2897 = ( wire1927 ) | ( wire1929 ) | ( wire1930 ) | ( wire8123 ) ;
 assign n_n2907 = ( wire1919 ) | ( wire1921 ) | ( wire1922 ) | ( wire8128 ) ;
 assign n_n2923 = ( wire1911 ) | ( wire1913 ) | ( wire1914 ) | ( wire8133 ) ;
 assign n_n2933 = ( wire1903 ) | ( wire1905 ) | ( wire1906 ) | ( wire8138 ) ;
 assign n_n2948 = ( wire1895 ) | ( wire1897 ) | ( wire1898 ) | ( wire8143 ) ;
 assign n_n2959 = ( wire1887 ) | ( wire1889 ) | ( wire1890 ) | ( wire8148 ) ;
 assign n_n2742 = ( wire1879 ) | ( wire1881 ) | ( wire1882 ) | ( wire8153 ) ;
 assign n_n2898 = ( wire1871 ) | ( wire1873 ) | ( wire1874 ) | ( wire8158 ) ;
 assign n_n2911 = ( wire1863 ) | ( wire1865 ) | ( wire1866 ) | ( wire8163 ) ;
 assign n_n2919 = ( wire1855 ) | ( wire1857 ) | ( wire1858 ) | ( wire8168 ) ;
 assign n_n2932 = ( wire1847 ) | ( wire1849 ) | ( wire1850 ) | ( wire8173 ) ;
 assign n_n2949 = ( wire1839 ) | ( wire1841 ) | ( wire1842 ) | ( wire8178 ) ;
 assign n_n2962 = ( wire1831 ) | ( wire1833 ) | ( wire1834 ) | ( wire8183 ) ;
 assign n_n2743 = ( wire1825 ) | ( wire1827 ) | ( wire1828 ) | ( wire8188 ) ;
 assign n_n2900 = ( wire1817 ) | ( wire1819 ) | ( wire1820 ) | ( wire8193 ) ;
 assign n_n2910 = ( wire1809 ) | ( wire1811 ) | ( wire1812 ) | ( wire8198 ) ;
 assign n_n2920 = ( wire1801 ) | ( wire1803 ) | ( wire1804 ) | ( wire8203 ) ;
 assign n_n2930 = ( wire1793 ) | ( wire1795 ) | ( wire1796 ) | ( wire8208 ) ;
 assign n_n2951 = ( wire1785 ) | ( wire1787 ) | ( wire1788 ) | ( wire8213 ) ;
 assign n_n2961 = ( wire1777 ) | ( wire1779 ) | ( wire1780 ) | ( wire8218 ) ;
 assign n_n2734 = ( wire1771 ) | ( wire1773 ) | ( wire1774 ) | ( wire8223 ) ;
 assign n_n2858 = ( wire1765 ) | ( wire1767 ) | ( wire1768 ) | ( wire8228 ) ;
 assign n_n2870 = ( wire1759 ) | ( wire1761 ) | ( wire1762 ) | ( wire8233 ) ;
 assign n_n2901 = ( wire1751 ) | ( wire1753 ) | ( wire1754 ) | ( wire8238 ) ;
 assign n_n2913 = ( wire1743 ) | ( wire1745 ) | ( wire1746 ) | ( wire8243 ) ;
 assign n_n2926 = ( wire1735 ) | ( wire1737 ) | ( wire1738 ) | ( wire8248 ) ;
 assign n_n2938 = ( wire1727 ) | ( wire1729 ) | ( wire1730 ) | ( wire8253 ) ;
 assign n_n2941 = ( wire1719 ) | ( wire1721 ) | ( wire1722 ) | ( wire8258 ) ;
 assign n_n2956 = ( wire1711 ) | ( wire1713 ) | ( wire1714 ) | ( wire8263 ) ;
 assign n_n2973 = ( wire1703 ) | ( wire1705 ) | ( wire1706 ) | ( wire8268 ) ;
 assign n_n2987 = ( wire1697 ) | ( wire1699 ) | ( wire1700 ) | ( wire8273 ) ;
 assign n_n2735 = ( wire1691 ) | ( wire1693 ) | ( wire1694 ) | ( wire8278 ) ;
 assign n_n2859 = ( wire1685 ) | ( wire1687 ) | ( wire1688 ) | ( wire8283 ) ;
 assign n_n2869 = ( wire1679 ) | ( wire1681 ) | ( wire1682 ) | ( wire8288 ) ;
 assign n_n2902 = ( wire1671 ) | ( wire1673 ) | ( wire1674 ) | ( wire8293 ) ;
 assign n_n2912 = ( wire1663 ) | ( wire1665 ) | ( wire1666 ) | ( wire8298 ) ;
 assign n_n2927 = ( wire1655 ) | ( wire1657 ) | ( wire1658 ) | ( wire8303 ) ;
 assign n_n2937 = ( wire1647 ) | ( wire1649 ) | ( wire1650 ) | ( wire8308 ) ;
 assign n_n2942 = ( wire1639 ) | ( wire1641 ) | ( wire1642 ) | ( wire8313 ) ;
 assign n_n2955 = ( wire1631 ) | ( wire1633 ) | ( wire1634 ) | ( wire8318 ) ;
 assign n_n2974 = ( wire1623 ) | ( wire1625 ) | ( wire1626 ) | ( wire8323 ) ;
 assign n_n2985 = ( wire1617 ) | ( wire1619 ) | ( wire1620 ) | ( wire8328 ) ;
 assign n_n2736 = ( wire1611 ) | ( wire1613 ) | ( wire1614 ) | ( wire8333 ) ;
 assign n_n2882 = ( wire1603 ) | ( wire1605 ) | ( wire1606 ) | ( wire8338 ) ;
 assign n_n2895 = ( wire1595 ) | ( wire1597 ) | ( wire1598 ) | ( wire8343 ) ;
 assign n_n2903 = ( wire1587 ) | ( wire1589 ) | ( wire1590 ) | ( wire8348 ) ;
 assign n_n2915 = ( wire1579 ) | ( wire1581 ) | ( wire1582 ) | ( wire8353 ) ;
 assign n_n2924 = ( wire1571 ) | ( wire1573 ) | ( wire1574 ) | ( wire8358 ) ;
 assign n_n2936 = ( wire1563 ) | ( wire1565 ) | ( wire1566 ) | ( wire8363 ) ;
 assign n_n2944 = ( wire1555 ) | ( wire1557 ) | ( wire1558 ) | ( wire8368 ) ;
 assign n_n2958 = ( wire1547 ) | ( wire1549 ) | ( wire1550 ) | ( wire8373 ) ;
 assign n_n2975 = ( wire1539 ) | ( wire1541 ) | ( wire1542 ) | ( wire8378 ) ;
 assign n_n2738 = ( wire1533 ) | ( wire1535 ) | ( wire1536 ) | ( wire8383 ) ;
 assign n_n2883 = ( wire1525 ) | ( wire1527 ) | ( wire1528 ) | ( wire8388 ) ;
 assign n_n2894 = ( wire1517 ) | ( wire1519 ) | ( wire1520 ) | ( wire8393 ) ;
 assign n_n2904 = ( wire1509 ) | ( wire1511 ) | ( wire1512 ) | ( wire8398 ) ;
 assign n_n2914 = ( wire1501 ) | ( wire1503 ) | ( wire1504 ) | ( wire8403 ) ;
 assign n_n2925 = ( wire1493 ) | ( wire1495 ) | ( wire1496 ) | ( wire8408 ) ;
 assign n_n2935 = ( wire1485 ) | ( wire1487 ) | ( wire1488 ) | ( wire8413 ) ;
 assign n_n2946 = ( wire1477 ) | ( wire1479 ) | ( wire1480 ) | ( wire8418 ) ;
 assign n_n2957 = ( wire1469 ) | ( wire1471 ) | ( wire1472 ) | ( wire8423 ) ;
 assign n_n2988 = ( wire1463 ) | ( wire1465 ) | ( wire1466 ) | ( wire8428 ) ;
 assign n_n2792 = ( wire1457 ) | ( wire1459 ) | ( wire1460 ) | ( wire8433 ) ;
 assign n_n2804 = ( wire1451 ) | ( wire1453 ) | ( wire1454 ) | ( wire8438 ) ;
 assign n_n2817 = ( wire1445 ) | ( wire1447 ) | ( wire1448 ) | ( wire8443 ) ;
 assign n_n2829 = ( wire1439 ) | ( wire1441 ) | ( wire1442 ) | ( wire8448 ) ;
 assign n_n2842 = ( wire1433 ) | ( wire1435 ) | ( wire1436 ) | ( wire8453 ) ;
 assign n_n2793 = ( wire1427 ) | ( wire1429 ) | ( wire1430 ) | ( wire8458 ) ;
 assign n_n2803 = ( wire1421 ) | ( wire1423 ) | ( wire1424 ) | ( wire8463 ) ;
 assign n_n2818 = ( wire1415 ) | ( wire1417 ) | ( wire1418 ) | ( wire8468 ) ;
 assign n_n2828 = ( wire1409 ) | ( wire1411 ) | ( wire1412 ) | ( wire8473 ) ;
 assign n_n2844 = ( wire1403 ) | ( wire1405 ) | ( wire1406 ) | ( wire8478 ) ;
 assign n_n2794 = ( wire1397 ) | ( wire1399 ) | ( wire1400 ) | ( wire8483 ) ;
 assign n_n2807 = ( wire1391 ) | ( wire1393 ) | ( wire1394 ) | ( wire8488 ) ;
 assign n_n2815 = ( wire1385 ) | ( wire1387 ) | ( wire1388 ) | ( wire8493 ) ;
 assign n_n2827 = ( wire1379 ) | ( wire1381 ) | ( wire1382 ) | ( wire8498 ) ;
 assign n_n2845 = ( wire1373 ) | ( wire1375 ) | ( wire1376 ) | ( wire8503 ) ;
 assign n_n2733 = ( wire1367 ) | ( wire1369 ) | ( wire1370 ) | ( wire8508 ) ;
 assign n_n2795 = ( wire1361 ) | ( wire1363 ) | ( wire1364 ) | ( wire8513 ) ;
 assign n_n2805 = ( wire1355 ) | ( wire1357 ) | ( wire1358 ) | ( wire8518 ) ;
 assign n_n2816 = ( wire1349 ) | ( wire1351 ) | ( wire1352 ) | ( wire8523 ) ;
 assign n_n2826 = ( wire1343 ) | ( wire1345 ) | ( wire1346 ) | ( wire8528 ) ;
 assign n_n2846 = ( wire1337 ) | ( wire1339 ) | ( wire1340 ) | ( wire8533 ) ;
 assign n_n2745 = ( wire1331 ) | ( wire1333 ) | ( wire1334 ) | ( wire8538 ) ;
 assign n_n2759 = ( wire1325 ) | ( wire1327 ) | ( wire1328 ) | ( wire8543 ) ;
 assign n_n2771 = ( wire1319 ) | ( wire1321 ) | ( wire1322 ) | ( wire8548 ) ;
 assign n_n2784 = ( wire1313 ) | ( wire1315 ) | ( wire1316 ) | ( wire8553 ) ;
 assign n_n2847 = ( wire1307 ) | ( wire1309 ) | ( wire1310 ) | ( wire8558 ) ;
 assign n_n2747 = ( wire1301 ) | ( wire1303 ) | ( wire1304 ) | ( wire8563 ) ;
 assign n_n2758 = ( wire1295 ) | ( wire1297 ) | ( wire1298 ) | ( wire8568 ) ;
 assign n_n2772 = ( wire1289 ) | ( wire1291 ) | ( wire1292 ) | ( wire8573 ) ;
 assign n_n2783 = ( wire1283 ) | ( wire1285 ) | ( wire1286 ) | ( wire8578 ) ;
 assign n_n2848 = ( wire1277 ) | ( wire1279 ) | ( wire1280 ) | ( wire8583 ) ;
 assign n_n2748 = ( wire1271 ) | ( wire1273 ) | ( wire1274 ) | ( wire8588 ) ;
 assign n_n2761 = ( wire1265 ) | ( wire1267 ) | ( wire1268 ) | ( wire8593 ) ;
 assign n_n2768 = ( wire1259 ) | ( wire1261 ) | ( wire1262 ) | ( wire8598 ) ;
 assign n_n2782 = ( wire1253 ) | ( wire1255 ) | ( wire1256 ) | ( wire8603 ) ;
 assign n_n2750 = ( wire1247 ) | ( wire1249 ) | ( wire1250 ) | ( wire8608 ) ;
 assign n_n2760 = ( wire1241 ) | ( wire1243 ) | ( wire1244 ) | ( wire8613 ) ;
 assign n_n2769 = ( wire1235 ) | ( wire1237 ) | ( wire1238 ) | ( wire8618 ) ;
 assign n_n2781 = ( wire1229 ) | ( wire1231 ) | ( wire1232 ) | ( wire8623 ) ;
 assign n_n2751 = ( wire1223 ) | ( wire1225 ) | ( wire1226 ) | ( wire8628 ) ;
 assign n_n2763 = ( wire1217 ) | ( wire1219 ) | ( wire1220 ) | ( wire8633 ) ;
 assign n_n2776 = ( wire1211 ) | ( wire1213 ) | ( wire1214 ) | ( wire8638 ) ;
 assign n_n2788 = ( wire1205 ) | ( wire1207 ) | ( wire1208 ) | ( wire8643 ) ;
 assign n_n2800 = ( wire1199 ) | ( wire1201 ) | ( wire1202 ) | ( wire8648 ) ;
 assign n_n2814 = ( wire1193 ) | ( wire1195 ) | ( wire1196 ) | ( wire8653 ) ;
 assign n_n2752 = ( wire1187 ) | ( wire1189 ) | ( wire1190 ) | ( wire8658 ) ;
 assign n_n2762 = ( wire1181 ) | ( wire1183 ) | ( wire1184 ) | ( wire8663 ) ;
 assign n_n2777 = ( wire1175 ) | ( wire1177 ) | ( wire1178 ) | ( wire8668 ) ;
 assign n_n2787 = ( wire1169 ) | ( wire1171 ) | ( wire1172 ) | ( wire8673 ) ;
 assign n_n2801 = ( wire1163 ) | ( wire1165 ) | ( wire1166 ) | ( wire8678 ) ;
 assign n_n2813 = ( wire1157 ) | ( wire1159 ) | ( wire1160 ) | ( wire8683 ) ;
 assign n_n2753 = ( wire1151 ) | ( wire1153 ) | ( wire1154 ) | ( wire8688 ) ;
 assign n_n2765 = ( wire1145 ) | ( wire1147 ) | ( wire1148 ) | ( wire8693 ) ;
 assign n_n2773 = ( wire1139 ) | ( wire1141 ) | ( wire1142 ) | ( wire8698 ) ;
 assign n_n2786 = ( wire1133 ) | ( wire1135 ) | ( wire1136 ) | ( wire8703 ) ;
 assign n_n2824 = ( wire1127 ) | ( wire1129 ) | ( wire1130 ) | ( wire8708 ) ;
 assign n_n2836 = ( wire1121 ) | ( wire1123 ) | ( wire1124 ) | ( wire8713 ) ;
 assign n_n2754 = ( wire1115 ) | ( wire1117 ) | ( wire1118 ) | ( wire8718 ) ;
 assign n_n2764 = ( wire1109 ) | ( wire1111 ) | ( wire1112 ) | ( wire8723 ) ;
 assign n_n2775 = ( wire1103 ) | ( wire1105 ) | ( wire1106 ) | ( wire8728 ) ;
 assign n_n2785 = ( wire1097 ) | ( wire1099 ) | ( wire1100 ) | ( wire8733 ) ;
 assign n_n2825 = ( wire1091 ) | ( wire1093 ) | ( wire1094 ) | ( wire8738 ) ;
 assign n_n2835 = ( wire1085 ) | ( wire1087 ) | ( wire1088 ) | ( wire8743 ) ;
 assign n_n2755 = ( wire1079 ) | ( wire1081 ) | ( wire1082 ) | ( wire8748 ) ;
 assign n_n2767 = ( wire1073 ) | ( wire1075 ) | ( wire1076 ) | ( wire8753 ) ;
 assign n_n2796 = ( wire1067 ) | ( wire1069 ) | ( wire1070 ) | ( wire8758 ) ;
 assign n_n2809 = ( wire1061 ) | ( wire1063 ) | ( wire1064 ) | ( wire8763 ) ;
 assign n_n2822 = ( wire1055 ) | ( wire1057 ) | ( wire1058 ) | ( wire8768 ) ;
 assign n_n2833 = ( wire1049 ) | ( wire1051 ) | ( wire1052 ) | ( wire8773 ) ;
 assign n_n2837 = ( wire1043 ) | ( wire1045 ) | ( wire1046 ) | ( wire8778 ) ;
 assign n_n2756 = ( wire1037 ) | ( wire1039 ) | ( wire1040 ) | ( wire8783 ) ;
 assign n_n2766 = ( wire1031 ) | ( wire1033 ) | ( wire1034 ) | ( wire8788 ) ;
 assign n_n2797 = ( wire1025 ) | ( wire1027 ) | ( wire1028 ) | ( wire8793 ) ;
 assign n_n2808 = ( wire1019 ) | ( wire1021 ) | ( wire1022 ) | ( wire8798 ) ;
 assign n_n2823 = ( wire1013 ) | ( wire1015 ) | ( wire1016 ) | ( wire8803 ) ;
 assign n_n2832 = ( wire1007 ) | ( wire1009 ) | ( wire1010 ) | ( wire8808 ) ;
 assign n_n2839 = ( wire1001 ) | ( wire1003 ) | ( wire1004 ) | ( wire8813 ) ;
 assign n_n2778 = ( wire995 ) | ( wire997 ) | ( wire998 ) | ( wire8818 ) ;
 assign n_n2791 = ( wire989 ) | ( wire991 ) | ( wire992 ) | ( wire8823 ) ;
 assign n_n2798 = ( wire983 ) | ( wire985 ) | ( wire986 ) | ( wire8828 ) ;
 assign n_n2812 = ( wire977 ) | ( wire979 ) | ( wire980 ) | ( wire8833 ) ;
 assign n_n2819 = ( wire971 ) | ( wire973 ) | ( wire974 ) | ( wire8838 ) ;
 assign n_n2831 = ( wire965 ) | ( wire967 ) | ( wire968 ) | ( wire8843 ) ;
 assign n_n2840 = ( wire959 ) | ( wire961 ) | ( wire962 ) | ( wire8848 ) ;
 assign n_n2780 = ( wire953 ) | ( wire955 ) | ( wire956 ) | ( wire8853 ) ;
 assign n_n2790 = ( wire947 ) | ( wire949 ) | ( wire950 ) | ( wire8858 ) ;
 assign n_n2799 = ( wire941 ) | ( wire943 ) | ( wire944 ) | ( wire8863 ) ;
 assign n_n2810 = ( wire935 ) | ( wire937 ) | ( wire938 ) | ( wire8868 ) ;
 assign n_n2820 = ( wire929 ) | ( wire931 ) | ( wire932 ) | ( wire8873 ) ;
 assign n_n2830 = ( wire923 ) | ( wire925 ) | ( wire926 ) | ( wire8878 ) ;
 assign n_n2841 = ( wire917 ) | ( wire919 ) | ( wire920 ) | ( wire8883 ) ;
 assign wire891 = ( (~ pcount_0_)  &  (~ pencrypt_0_)  &  wire887 ) | ( pcount_0_  &  pencrypt_0_  &  wire890 ) ;
 assign wire894 = ( pcount_2_  &  (~ pcount_1_)  &  pencrypt_0_ ) | ( pcount_2_  &  (~ pcount_0_)  &  pencrypt_0_ ) | ( pcount_2_  &  pcount_1_  &  (~ pencrypt_0_) ) | ( pcount_2_  &  pcount_0_  &  (~ pencrypt_0_) ) | ( (~ pcount_2_)  &  pcount_1_  &  pcount_0_  &  pencrypt_0_ ) | ( (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) ;
 assign wire775 = ( pksi_117_ ) | ( pksi_17_ ) ;
 assign wire776 = ( pksi_185_ ) | ( n_n2737 ) ;
 assign wire777 = ( pksi_72_ ) | ( n_n2879 ) ;
 assign wire778 = ( pksi_170_ ) | ( pksi_78_ ) ;
 assign wire779 = ( pksi_69_ ) | ( pksi_155_ ) ;
 assign wire780 = ( pksi_147_ ) | ( n_n2789 ) ;
 assign wire781 = ( pksi_109_ ) | ( pksi_10_ ) ;
 assign wire782 = ( pksi_11_ ) | ( n_n2982 ) ;
 assign wire783 = ( pksi_188_ ) | ( n_n2741 ) ;
 assign wire887 = ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_) ) ;
 assign wire890 = ( pcount_3_  &  pcount_2_  &  pcount_1_ ) ;
 assign n_n2997 = ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_) ) | ( (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_) ) | ( pcount_3_  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) ;
 assign wire774 = ( (~ pcount_3_)  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) ;
 assign n_n2993 = ( (~ pcount_3_)  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) | ( pcount_3_  &  pcount_2_  &  pcount_1_  &  (~ pcount_0_) ) | ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_) ) ;
 assign wire784 = ( pksi_94_ ) | ( n_n2881 ) ;
 assign wire785 = ( pksi_95_ ) | ( pksi_174_ ) ;
 assign wire786 = ( pksi_61_ ) | ( pksi_148_ ) ;
 assign wire787 = ( pksi_65_ ) | ( pksi_165_ ) ;
 assign wire788 = ( pksi_137_ ) | ( n_n2802 ) ;
 assign wire789 = ( pksi_122_ ) | ( pksi_30_ ) ;
 assign wire790 = ( pksi_114_ ) | ( n_n2843 ) ;
 assign wire791 = ( pksi_71_ ) | ( pksi_150_ ) ;
 assign wire792 = ( pksi_42_ ) | ( pksi_132_ ) ;
 assign wire793 = ( pksi_19_ ) | ( n_n2986 ) ;
 assign wire794 = ( n_n2865 ) | ( n_n2280 ) ;
 assign wire795 = ( pksi_87_ ) | ( n_n2391 ) ;
 assign wire796 = ( pksi_59_ ) | ( n_n2917 ) ;
 assign wire797 = ( pksi_107_ ) | ( pksi_21_ ) ;
 assign wire798 = ( pksi_110_ ) | ( pksi_2_ ) ;
 assign wire799 = ( pksi_84_ ) | ( pksi_176_ ) ;
 assign wire800 = ( pksi_86_ ) | ( pksi_175_ ) ;
 assign wire801 = ( pksi_162_ ) | ( n_n2779 ) ;
 assign wire802 = ( pksi_27_ ) | ( pksi_121_ ) ;
 assign wire803 = ( pksi_39_ ) | ( n_n2438 ) ;
 assign wire804 = ( pksi_105_ ) | ( pksi_1_ ) ;
 assign wire805 = ( pksi_52_ ) | ( pksi_166_ ) ;
 assign wire806 = ( pksi_129_ ) | ( pksi_25_ ) ;
 assign wire807 = ( pksi_126_ ) | ( pksi_47_ ) ;
 assign wire808 = ( pksi_100_ ) | ( pksi_13_ ) ;
 assign wire809 = ( pksi_112_ ) | ( pksi_9_ ) ;
 assign wire810 = ( pksi_180_ ) | ( n_n2749 ) ;
 assign wire811 = ( pksi_77_ ) | ( pksi_178_ ) ;
 assign wire812 = ( pksi_31_ ) | ( pksi_135_ ) ;
 assign wire813 = ( pksi_118_ ) | ( pksi_4_ ) ;
 assign wire814 = ( pksi_93_ ) | ( pksi_179_ ) ;
 assign wire815 = ( pksi_74_ ) | ( pksi_182_ ) ;
 assign wire816 = ( pksi_55_ ) | ( pksi_159_ ) ;
 assign wire817 = ( pksi_58_ ) | ( pksi_157_ ) ;
 assign wire818 = ( pksi_128_ ) | ( pksi_36_ ) ;
 assign wire819 = ( pksi_142_ ) | ( pksi_28_ ) ;
 assign wire820 = ( pksi_24_ ) | ( n_n2945 ) ;
 assign wire821 = ( pksi_106_ ) | ( pksi_5_ ) ;
 assign wire822 = ( pksi_75_ ) | ( pksi_169_ ) ;
 assign wire823 = ( pksi_80_ ) | ( n_n2877 ) ;
 assign wire824 = ( pksi_81_ ) | ( pksi_184_ ) ;
 assign wire825 = ( pksi_125_ ) | ( pksi_44_ ) ;
 assign wire826 = ( pksi_138_ ) | ( n_n2811 ) ;
 assign wire827 = ( pksi_99_ ) | ( n_n2853 ) ;
 assign wire828 = ( pksi_82_ ) | ( n_n2379 ) ;
 assign wire829 = ( pksi_83_ ) | ( n_n2885 ) ;
 assign wire830 = ( pksi_76_ ) | ( pksi_190_ ) ;
 assign wire831 = ( pksi_50_ ) | ( pksi_158_ ) ;
 assign wire832 = ( pksi_140_ ) | ( n_n2806 ) ;
 assign wire833 = ( pksi_32_ ) | ( n_n2943 ) ;
 assign wire834 = ( pksi_85_ ) | ( pksi_172_ ) ;
 assign wire835 = ( pksi_14_ ) | ( pksi_103_ ) ;
 assign wire836 = ( pksi_186_ ) | ( n_n2746 ) ;
 assign wire837 = ( pksi_91_ ) | ( n_n2889 ) ;
 assign wire838 = ( pksi_41_ ) | ( pksi_141_ ) ;
 assign wire839 = ( pksi_113_ ) | ( n_n2834 ) ;
 assign wire840 = ( pksi_115_ ) | ( pksi_0_ ) ;
 assign wire841 = ( pksi_98_ ) | ( pksi_6_ ) ;
 assign wire842 = ( pksi_34_ ) | ( pksi_133_ ) ;
 assign wire843 = ( pksi_43_ ) | ( n_n2954 ) ;
 assign wire844 = ( pksi_40_ ) | ( n_n2931 ) ;
 assign wire845 = ( pksi_45_ ) | ( pksi_131_ ) ;
 assign wire846 = ( pksi_102_ ) | ( pksi_23_ ) ;
 assign wire847 = ( pksi_73_ ) | ( pksi_177_ ) ;
 assign wire848 = ( pksi_189_ ) | ( pksi_89_ ) ;
 assign wire849 = ( pksi_16_ ) | ( n_n2964 ) ;
 assign wire850 = ( pksi_97_ ) | ( pksi_3_ ) ;
 assign wire851 = ( pksi_92_ ) | ( pksi_173_ ) ;
 assign wire852 = ( pksi_171_ ) | ( n_n2757 ) ;
 assign wire853 = ( pksi_12_ ) | ( pksi_104_ ) ;
 assign wire854 = ( pksi_29_ ) | ( pksi_130_ ) ;
 assign wire855 = ( pksi_183_ ) | ( pksi_79_ ) ;
 assign wire856 = ( pksi_116_ ) | ( n_n2838 ) ;
 assign wire857 = ( pksi_96_ ) | ( pksi_22_ ) ;
 assign wire858 = ( pksi_119_ ) | ( pksi_15_ ) ;
 assign wire859 = ( pksi_33_ ) | ( pksi_136_ ) ;
 assign wire860 = ( pksi_124_ ) | ( pksi_37_ ) ;
 assign wire861 = ( pksi_49_ ) | ( n_n2909 ) ;
 assign wire862 = ( pksi_57_ ) | ( pksi_160_ ) ;
 assign wire863 = ( pksi_127_ ) | ( pksi_38_ ) ;
 assign wire864 = ( pksi_164_ ) | ( n_n2774 ) ;
 assign wire865 = ( pksi_68_ ) | ( pksi_149_ ) ;
 assign wire866 = ( pksi_53_ ) | ( pksi_154_ ) ;
 assign wire867 = ( pksi_26_ ) | ( pksi_134_ ) ;
 assign wire868 = ( pksi_60_ ) | ( pksi_152_ ) ;
 assign wire869 = ( pksi_35_ ) | ( n_n2950 ) ;
 assign wire870 = ( pksi_101_ ) | ( pksi_20_ ) ;
 assign wire871 = ( pksi_64_ ) | ( n_n2899 ) ;
 assign wire872 = ( pksi_56_ ) | ( pksi_153_ ) ;
 assign wire873 = ( pksi_70_ ) | ( pksi_144_ ) ;
 assign wire874 = ( pksi_8_ ) | ( n_n2976 ) ;
 assign wire875 = ( pksi_123_ ) | ( n_n2821 ) ;
 assign wire876 = ( pksi_111_ ) | ( pksi_7_ ) ;
 assign wire877 = ( pksi_161_ ) | ( n_n2770 ) ;
 assign wire878 = ( pksi_66_ ) | ( pksi_156_ ) ;
 assign wire879 = ( pksi_67_ ) | ( n_n2921 ) ;
 assign wire880 = ( pksi_62_ ) | ( pksi_151_ ) ;
 assign wire881 = ( pksi_54_ ) | ( pksi_146_ ) ;
 assign wire882 = ( pksi_108_ ) | ( pksi_18_ ) ;
 assign wire883 = ( pksi_51_ ) | ( pksi_145_ ) ;
 assign wire884 = ( pksi_63_ ) | ( pksi_167_ ) ;
 assign wire885 = ( pksi_163_ ) | ( pksi_48_ ) ;
 assign wire886 = ( pksi_120_ ) | ( pksi_46_ ) ;
 assign wire893 = ( (~ pcount_2_)  &  pencrypt_0_ ) | ( (~ pcount_1_)  &  pencrypt_0_ ) | ( (~ pcount_0_)  &  pencrypt_0_ ) | ( pcount_2_  &  (~ pencrypt_0_) ) | ( pcount_1_  &  (~ pencrypt_0_) ) | ( pcount_0_  &  (~ pencrypt_0_) ) ;
 assign pksi_90_ = ( n_n2280 ) ;
 assign pksi_191_ = ( n_n2391 ) ;
 assign pksi_187_ = ( n_n2391 ) ;
 assign pksi_168_ = ( n_n2379 ) ;
 assign pksi_181_ = ( n_n2379 ) ;
 assign pksi_88_ = ( n_n2280 ) ;
 assign pksi_143_ = ( n_n2438 ) ;
 assign pksi_139_ = ( n_n2438 ) ;
 assign wire907 = ( pcount_3_  &  wire893 ) ;
 assign wire917 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8881 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8881 ) ;
 assign wire919 = ( pksi_100_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_13_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire920 = ( (~ pksi_100_)  &  pksi_13_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_100_  &  (~ pksi_13_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire923 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8876 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8876 ) ;
 assign wire925 = ( pksi_111_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_7_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire926 = ( (~ pksi_111_)  &  pksi_7_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_111_  &  (~ pksi_7_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire929 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8871 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8871 ) ;
 assign wire931 = ( pksi_123_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2821  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire932 = ( (~ pksi_123_)  &  n_n2821  &  (~ n_n2993)  &  wire7765 ) | ( pksi_123_  &  (~ n_n2821)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire935 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8866 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8866 ) ;
 assign wire937 = ( pksi_138_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2811  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire938 = ( (~ pksi_138_)  &  n_n2811  &  (~ n_n2993)  &  wire7765 ) | ( pksi_138_  &  (~ n_n2811)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire941 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8861 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8861 ) ;
 assign wire943 = ( pksi_125_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_44_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire944 = ( (~ pksi_125_)  &  pksi_44_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_125_  &  (~ pksi_44_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire947 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8856 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8856 ) ;
 assign wire949 = ( pksi_65_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_165_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire950 = ( (~ pksi_65_)  &  pksi_165_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_65_  &  (~ pksi_165_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire953 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8851 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8851 ) ;
 assign wire955 = ( pksi_49_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2909  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire956 = ( (~ pksi_49_)  &  n_n2909  &  (~ n_n2993)  &  wire7765 ) | ( pksi_49_  &  (~ n_n2909)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire959 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8846 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8846 ) ;
 assign wire961 = ( pksi_107_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_21_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire962 = ( (~ pksi_107_)  &  pksi_21_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_107_  &  (~ pksi_21_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire965 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8841 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8841 ) ;
 assign wire967 = ( pksi_101_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_20_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire968 = ( (~ pksi_101_)  &  pksi_20_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_101_  &  (~ pksi_20_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire971 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8836 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8836 ) ;
 assign wire973 = ( pksi_35_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2950  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire974 = ( (~ pksi_35_)  &  n_n2950  &  (~ n_n2993)  &  wire7765 ) | ( pksi_35_  &  (~ n_n2950)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire977 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8831 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8831 ) ;
 assign wire979 = ( pksi_129_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_25_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire980 = ( (~ pksi_129_)  &  pksi_25_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_129_  &  (~ pksi_25_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire983 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8826 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8826 ) ;
 assign wire985 = ( pksi_31_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_135_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire986 = ( (~ pksi_31_)  &  pksi_135_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_31_  &  (~ pksi_135_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire989 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8821 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8821 ) ;
 assign wire991 = ( pksi_67_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2921  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire992 = ( (~ pksi_67_)  &  n_n2921  &  (~ n_n2993)  &  wire7765 ) | ( pksi_67_  &  (~ n_n2921)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire995 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8816 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8816 ) ;
 assign wire997 = ( pksi_162_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2779  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire998 = ( (~ pksi_162_)  &  n_n2779  &  (~ n_n2993)  &  wire7765 ) | ( pksi_162_  &  (~ n_n2779)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1001 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8811 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8811 ) ;
 assign wire1003 = ( pksi_109_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_10_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1004 = ( (~ pksi_109_)  &  pksi_10_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_109_  &  (~ pksi_10_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1007 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8806 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8806 ) ;
 assign wire1009 = ( pksi_16_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2964  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1010 = ( (~ pksi_16_)  &  n_n2964  &  (~ n_n2993)  &  wire7765 ) | ( pksi_16_  &  (~ n_n2964)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1013 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8801 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8801 ) ;
 assign wire1015 = ( pksi_43_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2954  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1016 = ( (~ pksi_43_)  &  n_n2954  &  (~ n_n2993)  &  wire7765 ) | ( pksi_43_  &  (~ n_n2954)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1019 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8796 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8796 ) ;
 assign wire1021 = ( pksi_45_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_131_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1022 = ( (~ pksi_45_)  &  pksi_131_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_45_  &  (~ pksi_131_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1025 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8791 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8791 ) ;
 assign wire1027 = ( pksi_52_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_166_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1028 = ( (~ pksi_52_)  &  pksi_166_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_52_  &  (~ pksi_166_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1031 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8786 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8786 ) ;
 assign wire1033 = ( pksi_55_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_159_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1034 = ( (~ pksi_55_)  &  pksi_159_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_55_  &  (~ pksi_159_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1037 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8781 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8781 ) ;
 assign wire1039 = ( pksi_171_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2757  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1040 = ( (~ pksi_171_)  &  n_n2757  &  (~ n_n2993)  &  wire7765 ) | ( pksi_171_  &  (~ n_n2757)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1043 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8776 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8776 ) ;
 assign wire1045 = ( pksi_116_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2838  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1046 = ( (~ pksi_116_)  &  n_n2838  &  (~ n_n2993)  &  wire7765 ) | ( pksi_116_  &  (~ n_n2838)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1049 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8771 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8771 ) ;
 assign wire1051 = ( pksi_113_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2834  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1052 = ( (~ pksi_113_)  &  n_n2834  &  (~ n_n2993)  &  wire7765 ) | ( pksi_113_  &  (~ n_n2834)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1055 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8766 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8766 ) ;
 assign wire1057 = ( pksi_41_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_141_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1058 = ( (~ pksi_41_)  &  pksi_141_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_41_  &  (~ pksi_141_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1061 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8761 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8761 ) ;
 assign wire1063 = ( pksi_124_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_37_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1064 = ( (~ pksi_124_)  &  pksi_37_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_124_  &  (~ pksi_37_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1067 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8756 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8756 ) ;
 assign wire1069 = ( pksi_71_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_150_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1070 = ( (~ pksi_71_)  &  pksi_150_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_71_  &  (~ pksi_150_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1073 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8751 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8751 ) ;
 assign wire1075 = ( pksi_68_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_149_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1076 = ( (~ pksi_68_)  &  pksi_149_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_68_  &  (~ pksi_149_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1079 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8746 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8746 ) ;
 assign wire1081 = ( pksi_83_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2885  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1082 = ( (~ pksi_83_)  &  n_n2885  &  (~ n_n2993)  &  wire7765 ) | ( pksi_83_  &  (~ n_n2885)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1085 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8741 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8741 ) ;
 assign wire1087 = ( pksi_97_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_3_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1088 = ( (~ pksi_97_)  &  pksi_3_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_97_  &  (~ pksi_3_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1091 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8736 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8736 ) ;
 assign wire1093 = ( pksi_29_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_130_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1094 = ( (~ pksi_29_)  &  pksi_130_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_29_  &  (~ pksi_130_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1097 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8731 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8731 ) ;
 assign wire1099 = ( pksi_62_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_151_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1100 = ( (~ pksi_62_)  &  pksi_151_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_62_  &  (~ pksi_151_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1103 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8726 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8726 ) ;
 assign wire1105 = ( pksi_58_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_157_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1106 = ( (~ pksi_58_)  &  pksi_157_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_58_  &  (~ pksi_157_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1109 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8721 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8721 ) ;
 assign wire1111 = ( pksi_95_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_174_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1112 = ( (~ pksi_95_)  &  pksi_174_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_95_  &  (~ pksi_174_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1115 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8716 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8716 ) ;
 assign wire1117 = ( pksi_74_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_182_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1118 = ( (~ pksi_74_)  &  pksi_182_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_74_  &  (~ pksi_182_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1121 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8711 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8711 ) ;
 assign wire1123 = ( pksi_12_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_104_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1124 = ( (~ pksi_12_)  &  pksi_104_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_12_  &  (~ pksi_104_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1127 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8706 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8706 ) ;
 assign wire1129 = ( pksi_33_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_136_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1130 = ( (~ pksi_33_)  &  pksi_136_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_33_  &  (~ pksi_136_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1133 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8701 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8701 ) ;
 assign wire1135 = ( pksi_50_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_158_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1136 = ( (~ pksi_50_)  &  pksi_158_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_50_  &  (~ pksi_158_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1139 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8696 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8696 ) ;
 assign wire1141 = ( pksi_164_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2774  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1142 = ( (~ pksi_164_)  &  n_n2774  &  (~ n_n2993)  &  wire7765 ) | ( pksi_164_  &  (~ n_n2774)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1145 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8691 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8691 ) ;
 assign wire1147 = ( pksi_76_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_190_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1148 = ( (~ pksi_76_)  &  pksi_190_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_76_  &  (~ pksi_190_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1151 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8686 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8686 ) ;
 assign wire1153 = ( pksi_86_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_175_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1154 = ( (~ pksi_86_)  &  pksi_175_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_86_  &  (~ pksi_175_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1157 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8681 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8681 ) ;
 assign wire1159 = ( pksi_42_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_132_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1160 = ( (~ pksi_42_)  &  pksi_132_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_42_  &  (~ pksi_132_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1163 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8676 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8676 ) ;
 assign wire1165 = ( pksi_137_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2802  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1166 = ( (~ pksi_137_)  &  n_n2802  &  (~ n_n2993)  &  wire7765 ) | ( pksi_137_  &  (~ n_n2802)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1169 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8671 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8671 ) ;
 assign wire1171 = ( pksi_59_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2917  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1172 = ( (~ pksi_59_)  &  n_n2917  &  (~ n_n2993)  &  wire7765 ) | ( pksi_59_  &  (~ n_n2917)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1175 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8666 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8666 ) ;
 assign wire1177 = ( pksi_61_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_148_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1178 = ( (~ pksi_61_)  &  pksi_148_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_61_  &  (~ pksi_148_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1181 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8661 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8661 ) ;
 assign wire1183 = ( pksi_87_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2391  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1184 = ( (~ pksi_87_)  &  n_n2391  &  (~ n_n2993)  &  wire7765 ) | ( pksi_87_  &  (~ n_n2391)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1187 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8656 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8656 ) ;
 assign wire1189 = ( pksi_94_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2881  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1190 = ( (~ pksi_94_)  &  n_n2881  &  (~ n_n2993)  &  wire7765 ) | ( pksi_94_  &  (~ n_n2881)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1193 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8651 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8651 ) ;
 assign wire1195 = ( pksi_32_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2943  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1196 = ( (~ pksi_32_)  &  n_n2943  &  (~ n_n2993)  &  wire7765 ) | ( pksi_32_  &  (~ n_n2943)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1199 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8646 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8646 ) ;
 assign wire1201 = ( pksi_40_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2931  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1202 = ( (~ pksi_40_)  &  n_n2931  &  (~ n_n2993)  &  wire7765 ) | ( pksi_40_  &  (~ n_n2931)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1205 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8641 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8641 ) ;
 assign wire1207 = ( pksi_147_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2789  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1208 = ( (~ pksi_147_)  &  n_n2789  &  (~ n_n2993)  &  wire7765 ) | ( pksi_147_  &  (~ n_n2789)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1211 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8636 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8636 ) ;
 assign wire1213 = ( pksi_69_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_155_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1214 = ( (~ pksi_69_)  &  pksi_155_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_69_  &  (~ pksi_155_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1217 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8631 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8631 ) ;
 assign wire1219 = ( pksi_170_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_78_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1220 = ( (~ pksi_170_)  &  pksi_78_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_170_  &  (~ pksi_78_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1223 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8626 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8626 ) ;
 assign wire1225 = ( pksi_72_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2879  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1226 = ( (~ pksi_72_)  &  n_n2879  &  (~ n_n2993)  &  wire7765 ) | ( pksi_72_  &  (~ n_n2879)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1229 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8621 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8621 ) ;
 assign wire1231 = ( pksi_66_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_156_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1232 = ( (~ pksi_66_)  &  pksi_156_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_66_  &  (~ pksi_156_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1235 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8616 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8616 ) ;
 assign wire1237 = ( pksi_161_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2770  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1238 = ( (~ pksi_161_)  &  n_n2770  &  (~ n_n2993)  &  wire7765 ) | ( pksi_161_  &  (~ n_n2770)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1241 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8611 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8611 ) ;
 assign wire1243 = ( pksi_81_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_184_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1244 = ( (~ pksi_81_)  &  pksi_184_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_81_  &  (~ pksi_184_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1247 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8606 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8606 ) ;
 assign wire1249 = ( pksi_80_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2877  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1250 = ( (~ pksi_80_)  &  n_n2877  &  (~ n_n2993)  &  wire7765 ) | ( pksi_80_  &  (~ n_n2877)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1253 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8601 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8601 ) ;
 assign wire1255 = ( pksi_56_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_153_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1256 = ( (~ pksi_56_)  &  pksi_153_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_56_  &  (~ pksi_153_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1259 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8596 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8596 ) ;
 assign wire1261 = ( pksi_64_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2899  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1262 = ( (~ pksi_64_)  &  n_n2899  &  (~ n_n2993)  &  wire7765 ) | ( pksi_64_  &  (~ n_n2899)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1265 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8591 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8591 ) ;
 assign wire1267 = ( pksi_77_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_178_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1268 = ( (~ pksi_77_)  &  pksi_178_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_77_  &  (~ pksi_178_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1271 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8586 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8586 ) ;
 assign wire1273 = ( pksi_180_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2749  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1274 = ( (~ pksi_180_)  &  n_n2749  &  (~ n_n2993)  &  wire7765 ) | ( pksi_180_  &  (~ n_n2749)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1277 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8581 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8581 ) ;
 assign wire1279 = ( pksi_96_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_22_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1280 = ( (~ pksi_96_)  &  pksi_22_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_96_  &  (~ pksi_22_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1283 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8576 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8576 ) ;
 assign wire1285 = ( pksi_163_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_48_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1286 = ( (~ pksi_163_)  &  pksi_48_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_163_  &  (~ pksi_48_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1289 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8571 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8571 ) ;
 assign wire1291 = ( pksi_60_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_152_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1292 = ( (~ pksi_60_)  &  pksi_152_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_60_  &  (~ pksi_152_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1295 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8566 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8566 ) ;
 assign wire1297 = ( pksi_189_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_89_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1298 = ( (~ pksi_189_)  &  pksi_89_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_189_  &  (~ pksi_89_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1301 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8561 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8561 ) ;
 assign wire1303 = ( pksi_73_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_177_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1304 = ( (~ pksi_73_)  &  pksi_177_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_73_  &  (~ pksi_177_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1307 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8556 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8556 ) ;
 assign wire1309 = ( pksi_115_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_0_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1310 = ( (~ pksi_115_)  &  pksi_0_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_115_  &  (~ pksi_0_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1313 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8551 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8551 ) ;
 assign wire1315 = ( pksi_70_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_144_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1316 = ( (~ pksi_70_)  &  pksi_144_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_70_  &  (~ pksi_144_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1319 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8546 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8546 ) ;
 assign wire1321 = ( pksi_51_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_145_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1322 = ( (~ pksi_51_)  &  pksi_145_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_51_  &  (~ pksi_145_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1325 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8541 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8541 ) ;
 assign wire1327 = ( pksi_91_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2889  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1328 = ( (~ pksi_91_)  &  n_n2889  &  (~ n_n2993)  &  wire7765 ) | ( pksi_91_  &  (~ n_n2889)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1331 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8536 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8536 ) ;
 assign wire1333 = ( pksi_186_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2746  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1334 = ( (~ pksi_186_)  &  n_n2746  &  (~ n_n2993)  &  wire7765 ) | ( pksi_186_  &  (~ n_n2746)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1337 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8531 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8531 ) ;
 assign wire1339 = ( pksi_8_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2976  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1340 = ( (~ pksi_8_)  &  n_n2976  &  (~ n_n2993)  &  wire7765 ) | ( pksi_8_  &  (~ n_n2976)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1343 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8526 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8526 ) ;
 assign wire1345 = ( pksi_39_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2438  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1346 = ( (~ pksi_39_)  &  n_n2438  &  (~ n_n2993)  &  wire7765 ) | ( pksi_39_  &  (~ n_n2438)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1349 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8521 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8521 ) ;
 assign wire1351 = ( pksi_120_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_46_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1352 = ( (~ pksi_120_)  &  pksi_46_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_120_  &  (~ pksi_46_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1355 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8516 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8516 ) ;
 assign wire1357 = ( pksi_140_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2806  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1358 = ( (~ pksi_140_)  &  n_n2806  &  (~ n_n2993)  &  wire7765 ) | ( pksi_140_  &  (~ n_n2806)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1361 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8511 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8511 ) ;
 assign wire1363 = ( pksi_54_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_146_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1364 = ( (~ pksi_54_)  &  pksi_146_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_54_  &  (~ pksi_146_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1367 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8506 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8506 ) ;
 assign wire1369 = ( pksi_183_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_79_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1370 = ( (~ pksi_183_)  &  pksi_79_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_183_  &  (~ pksi_79_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1373 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8501 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8501 ) ;
 assign wire1375 = ( pksi_108_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_18_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1376 = ( (~ pksi_108_)  &  pksi_18_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_108_  &  (~ pksi_18_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1379 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8496 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8496 ) ;
 assign wire1381 = ( pksi_122_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_30_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1382 = ( (~ pksi_122_)  &  pksi_30_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_122_  &  (~ pksi_30_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1385 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8491 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8491 ) ;
 assign wire1387 = ( pksi_24_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2945  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1388 = ( (~ pksi_24_)  &  n_n2945  &  (~ n_n2993)  &  wire7765 ) | ( pksi_24_  &  (~ n_n2945)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1391 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8486 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8486 ) ;
 assign wire1393 = ( pksi_34_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_133_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1394 = ( (~ pksi_34_)  &  pksi_133_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_34_  &  (~ pksi_133_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1397 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8481 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8481 ) ;
 assign wire1399 = ( pksi_63_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_167_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1400 = ( (~ pksi_63_)  &  pksi_167_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_63_  &  (~ pksi_167_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1403 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8476 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8476 ) ;
 assign wire1405 = ( pksi_105_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_1_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1406 = ( (~ pksi_105_)  &  pksi_1_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_105_  &  (~ pksi_1_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1409 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8471 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8471 ) ;
 assign wire1411 = ( pksi_126_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_47_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1412 = ( (~ pksi_126_)  &  pksi_47_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_126_  &  (~ pksi_47_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1415 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8466 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8466 ) ;
 assign wire1417 = ( pksi_26_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_134_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1418 = ( (~ pksi_26_)  &  pksi_134_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_26_  &  (~ pksi_134_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1421 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8461 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8461 ) ;
 assign wire1423 = ( pksi_27_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_121_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1424 = ( (~ pksi_27_)  &  pksi_121_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_27_  &  (~ pksi_121_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1427 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8456 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8456 ) ;
 assign wire1429 = ( pksi_53_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_154_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1430 = ( (~ pksi_53_)  &  pksi_154_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_53_  &  (~ pksi_154_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1433 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8451 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8451 ) ;
 assign wire1435 = ( pksi_114_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2843  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1436 = ( (~ pksi_114_)  &  n_n2843  &  (~ n_n2993)  &  wire7765 ) | ( pksi_114_  &  (~ n_n2843)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1439 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8446 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8446 ) ;
 assign wire1441 = ( pksi_142_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_28_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1442 = ( (~ pksi_142_)  &  pksi_28_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_142_  &  (~ pksi_28_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1445 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8441 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8441 ) ;
 assign wire1447 = ( pksi_127_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_38_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1448 = ( (~ pksi_127_)  &  pksi_38_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_127_  &  (~ pksi_38_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1451 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8436 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8436 ) ;
 assign wire1453 = ( pksi_128_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_36_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1454 = ( (~ pksi_128_)  &  pksi_36_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_128_  &  (~ pksi_36_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1457 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8431 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8431 ) ;
 assign wire1459 = ( pksi_57_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_160_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1460 = ( (~ pksi_57_)  &  pksi_160_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_57_  &  (~ pksi_160_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1463 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8426 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8426 ) ;
 assign wire1465 = ( pksi_106_  &  n_n2997  &  wire7763 ) | ( pksi_5_  &  n_n2997  &  wire7763 ) ;
 assign wire1466 = ( (~ pksi_106_)  &  pksi_5_  &  n_n2993  &  wire7771 ) | ( pksi_106_  &  (~ pksi_5_)  &  n_n2993  &  wire7771 ) ;
 assign wire1469 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8421 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8421 ) ;
 assign wire1471 = ( pksi_39_  &  n_n2997  &  wire7763 ) | ( n_n2438  &  n_n2997  &  wire7763 ) ;
 assign wire1472 = ( (~ pksi_39_)  &  n_n2438  &  n_n2993  &  wire7771 ) | ( pksi_39_  &  (~ n_n2438)  &  n_n2993  &  wire7771 ) ;
 assign wire1477 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8416 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8416 ) ;
 assign wire1479 = ( pksi_120_  &  n_n2997  &  wire7763 ) | ( pksi_46_  &  n_n2997  &  wire7763 ) ;
 assign wire1480 = ( (~ pksi_120_)  &  pksi_46_  &  n_n2993  &  wire7771 ) | ( pksi_120_  &  (~ pksi_46_)  &  n_n2993  &  wire7771 ) ;
 assign wire1485 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8411 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8411 ) ;
 assign wire1487 = ( pksi_140_  &  n_n2997  &  wire7763 ) | ( n_n2806  &  n_n2997  &  wire7763 ) ;
 assign wire1488 = ( (~ pksi_140_)  &  n_n2806  &  n_n2993  &  wire7771 ) | ( pksi_140_  &  (~ n_n2806)  &  n_n2993  &  wire7771 ) ;
 assign wire1493 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8406 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8406 ) ;
 assign wire1495 = ( pksi_54_  &  n_n2997  &  wire7763 ) | ( pksi_146_  &  n_n2997  &  wire7763 ) ;
 assign wire1496 = ( (~ pksi_54_)  &  pksi_146_  &  n_n2993  &  wire7771 ) | ( pksi_54_  &  (~ pksi_146_)  &  n_n2993  &  wire7771 ) ;
 assign wire1501 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8401 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8401 ) ;
 assign wire1503 = ( pksi_62_  &  n_n2997  &  wire7763 ) | ( pksi_151_  &  n_n2997  &  wire7763 ) ;
 assign wire1504 = ( (~ pksi_62_)  &  pksi_151_  &  n_n2993  &  wire7771 ) | ( pksi_62_  &  (~ pksi_151_)  &  n_n2993  &  wire7771 ) ;
 assign wire1509 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8396 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8396 ) ;
 assign wire1511 = ( pksi_58_  &  n_n2997  &  wire7763 ) | ( pksi_157_  &  n_n2997  &  wire7763 ) ;
 assign wire1512 = ( (~ pksi_58_)  &  pksi_157_  &  n_n2993  &  wire7771 ) | ( pksi_58_  &  (~ pksi_157_)  &  n_n2993  &  wire7771 ) ;
 assign wire1517 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8391 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8391 ) ;
 assign wire1519 = ( pksi_95_  &  n_n2997  &  wire7763 ) | ( pksi_174_  &  n_n2997  &  wire7763 ) ;
 assign wire1520 = ( (~ pksi_95_)  &  pksi_174_  &  n_n2993  &  wire7771 ) | ( pksi_95_  &  (~ pksi_174_)  &  n_n2993  &  wire7771 ) ;
 assign wire1525 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8386 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8386 ) ;
 assign wire1527 = ( pksi_74_  &  n_n2997  &  wire7763 ) | ( pksi_182_  &  n_n2997  &  wire7763 ) ;
 assign wire1528 = ( (~ pksi_74_)  &  pksi_182_  &  n_n2993  &  wire7771 ) | ( pksi_74_  &  (~ pksi_182_)  &  n_n2993  &  wire7771 ) ;
 assign wire1533 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8381 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8381 ) ;
 assign wire1535 = ( pksi_75_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_169_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1536 = ( (~ pksi_75_)  &  pksi_169_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_75_  &  (~ pksi_169_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1539 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8376 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8376 ) ;
 assign wire1541 = ( pksi_8_  &  n_n2997  &  wire7763 ) | ( n_n2976  &  n_n2997  &  wire7763 ) ;
 assign wire1542 = ( (~ pksi_8_)  &  n_n2976  &  n_n2993  &  wire7771 ) | ( pksi_8_  &  (~ n_n2976)  &  n_n2993  &  wire7771 ) ;
 assign wire1547 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8371 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8371 ) ;
 assign wire1549 = ( pksi_122_  &  n_n2997  &  wire7763 ) | ( pksi_30_  &  n_n2997  &  wire7763 ) ;
 assign wire1550 = ( (~ pksi_122_)  &  pksi_30_  &  n_n2993  &  wire7771 ) | ( pksi_122_  &  (~ pksi_30_)  &  n_n2993  &  wire7771 ) ;
 assign wire1555 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8366 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8366 ) ;
 assign wire1557 = ( pksi_24_  &  n_n2997  &  wire7763 ) | ( n_n2945  &  n_n2997  &  wire7763 ) ;
 assign wire1558 = ( (~ pksi_24_)  &  n_n2945  &  n_n2993  &  wire7771 ) | ( pksi_24_  &  (~ n_n2945)  &  n_n2993  &  wire7771 ) ;
 assign wire1563 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8361 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8361 ) ;
 assign wire1565 = ( pksi_34_  &  n_n2997  &  wire7763 ) | ( pksi_133_  &  n_n2997  &  wire7763 ) ;
 assign wire1566 = ( (~ pksi_34_)  &  pksi_133_  &  n_n2993  &  wire7771 ) | ( pksi_34_  &  (~ pksi_133_)  &  n_n2993  &  wire7771 ) ;
 assign wire1571 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8356 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8356 ) ;
 assign wire1573 = ( pksi_63_  &  n_n2997  &  wire7763 ) | ( pksi_167_  &  n_n2997  &  wire7763 ) ;
 assign wire1574 = ( (~ pksi_63_)  &  pksi_167_  &  n_n2993  &  wire7771 ) | ( pksi_63_  &  (~ pksi_167_)  &  n_n2993  &  wire7771 ) ;
 assign wire1579 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8351 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8351 ) ;
 assign wire1581 = ( pksi_50_  &  n_n2997  &  wire7763 ) | ( pksi_158_  &  n_n2997  &  wire7763 ) ;
 assign wire1582 = ( (~ pksi_50_)  &  pksi_158_  &  n_n2993  &  wire7771 ) | ( pksi_50_  &  (~ pksi_158_)  &  n_n2993  &  wire7771 ) ;
 assign wire1587 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8346 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8346 ) ;
 assign wire1589 = ( pksi_164_  &  n_n2997  &  wire7763 ) | ( n_n2774  &  n_n2997  &  wire7763 ) ;
 assign wire1590 = ( (~ pksi_164_)  &  n_n2774  &  n_n2993  &  wire7771 ) | ( pksi_164_  &  (~ n_n2774)  &  n_n2993  &  wire7771 ) ;
 assign wire1595 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8341 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8341 ) ;
 assign wire1597 = ( pksi_76_  &  n_n2997  &  wire7763 ) | ( pksi_190_  &  n_n2997  &  wire7763 ) ;
 assign wire1598 = ( (~ pksi_76_)  &  pksi_190_  &  n_n2993  &  wire7771 ) | ( pksi_76_  &  (~ pksi_190_)  &  n_n2993  &  wire7771 ) ;
 assign wire1603 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8336 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8336 ) ;
 assign wire1605 = ( pksi_86_  &  n_n2997  &  wire7763 ) | ( pksi_175_  &  n_n2997  &  wire7763 ) ;
 assign wire1606 = ( (~ pksi_86_)  &  pksi_175_  &  n_n2993  &  wire7771 ) | ( pksi_86_  &  (~ pksi_175_)  &  n_n2993  &  wire7771 ) ;
 assign wire1611 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8331 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8331 ) ;
 assign wire1613 = ( pksi_185_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2737  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1614 = ( (~ pksi_185_)  &  n_n2737  &  (~ n_n2993)  &  wire7765 ) | ( pksi_185_  &  (~ n_n2737)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1617 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8326 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8326 ) ;
 assign wire1619 = ( pksi_19_  &  n_n2997  &  wire7763 ) | ( n_n2986  &  n_n2997  &  wire7763 ) ;
 assign wire1620 = ( (~ pksi_19_)  &  n_n2986  &  n_n2993  &  wire7771 ) | ( pksi_19_  &  (~ n_n2986)  &  n_n2993  &  wire7771 ) ;
 assign wire1623 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8321 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8321 ) ;
 assign wire1625 = ( pksi_108_  &  n_n2997  &  wire7763 ) | ( pksi_18_  &  n_n2997  &  wire7763 ) ;
 assign wire1626 = ( (~ pksi_108_)  &  pksi_18_  &  n_n2993  &  wire7771 ) | ( pksi_108_  &  (~ pksi_18_)  &  n_n2993  &  wire7771 ) ;
 assign wire1631 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8316 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8316 ) ;
 assign wire1633 = ( pksi_33_  &  n_n2997  &  wire7763 ) | ( pksi_136_  &  n_n2997  &  wire7763 ) ;
 assign wire1634 = ( (~ pksi_33_)  &  pksi_136_  &  n_n2993  &  wire7771 ) | ( pksi_33_  &  (~ pksi_136_)  &  n_n2993  &  wire7771 ) ;
 assign wire1639 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8311 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8311 ) ;
 assign wire1641 = ( pksi_32_  &  n_n2997  &  wire7763 ) | ( n_n2943  &  n_n2997  &  wire7763 ) ;
 assign wire1642 = ( (~ pksi_32_)  &  n_n2943  &  n_n2993  &  wire7771 ) | ( pksi_32_  &  (~ n_n2943)  &  n_n2993  &  wire7771 ) ;
 assign wire1647 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8306 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8306 ) ;
 assign wire1649 = ( pksi_45_  &  n_n2997  &  wire7763 ) | ( pksi_131_  &  n_n2997  &  wire7763 ) ;
 assign wire1650 = ( (~ pksi_45_)  &  pksi_131_  &  n_n2993  &  wire7771 ) | ( pksi_45_  &  (~ pksi_131_)  &  n_n2993  &  wire7771 ) ;
 assign wire1655 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8301 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8301 ) ;
 assign wire1657 = ( pksi_52_  &  n_n2997  &  wire7763 ) | ( pksi_166_  &  n_n2997  &  wire7763 ) ;
 assign wire1658 = ( (~ pksi_52_)  &  pksi_166_  &  n_n2993  &  wire7771 ) | ( pksi_52_  &  (~ pksi_166_)  &  n_n2993  &  wire7771 ) ;
 assign wire1663 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8296 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8296 ) ;
 assign wire1665 = ( pksi_163_  &  n_n2997  &  wire7763 ) | ( pksi_48_  &  n_n2997  &  wire7763 ) ;
 assign wire1666 = ( (~ pksi_163_)  &  pksi_48_  &  n_n2993  &  wire7771 ) | ( pksi_163_  &  (~ pksi_48_)  &  n_n2993  &  wire7771 ) ;
 assign wire1671 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8291 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8291 ) ;
 assign wire1673 = ( pksi_60_  &  n_n2997  &  wire7763 ) | ( pksi_152_  &  n_n2997  &  wire7763 ) ;
 assign wire1674 = ( (~ pksi_60_)  &  pksi_152_  &  n_n2993  &  wire7771 ) | ( pksi_60_  &  (~ pksi_152_)  &  n_n2993  &  wire7771 ) ;
 assign wire1679 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8286 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8286 ) ;
 assign wire1681 = ( pksi_188_  &  n_n2997  &  wire7763 ) | ( n_n2741  &  n_n2997  &  wire7763 ) ;
 assign wire1682 = ( (~ pksi_188_)  &  n_n2741  &  n_n2993  &  wire7771 ) | ( pksi_188_  &  (~ n_n2741)  &  n_n2993  &  wire7771 ) ;
 assign wire1685 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8281 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8281 ) ;
 assign wire1687 = ( pksi_98_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_6_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1688 = ( (~ pksi_98_)  &  pksi_6_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_98_  &  (~ pksi_6_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1691 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8276 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8276 ) ;
 assign wire1693 = ( n_n2865  &  (~ n_n2997)  &  wire7764 ) | ( n_n2280  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1694 = ( (~ n_n2865)  &  n_n2280  &  (~ n_n2993)  &  wire7765 ) | ( n_n2865  &  (~ n_n2280)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1697 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8271 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8271 ) ;
 assign wire1699 = ( pksi_112_  &  n_n2997  &  wire7763 ) | ( pksi_9_  &  n_n2997  &  wire7763 ) ;
 assign wire1700 = ( (~ pksi_112_)  &  pksi_9_  &  n_n2993  &  wire7771 ) | ( pksi_112_  &  (~ pksi_9_)  &  n_n2993  &  wire7771 ) ;
 assign wire1703 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8266 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8266 ) ;
 assign wire1705 = ( pksi_105_  &  n_n2997  &  wire7763 ) | ( pksi_1_  &  n_n2997  &  wire7763 ) ;
 assign wire1706 = ( (~ pksi_105_)  &  pksi_1_  &  n_n2993  &  wire7771 ) | ( pksi_105_  &  (~ pksi_1_)  &  n_n2993  &  wire7771 ) ;
 assign wire1711 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8261 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8261 ) ;
 assign wire1713 = ( pksi_29_  &  n_n2997  &  wire7763 ) | ( pksi_130_  &  n_n2997  &  wire7763 ) ;
 assign wire1714 = ( (~ pksi_29_)  &  pksi_130_  &  n_n2993  &  wire7771 ) | ( pksi_29_  &  (~ pksi_130_)  &  n_n2993  &  wire7771 ) ;
 assign wire1719 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8256 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8256 ) ;
 assign wire1721 = ( pksi_42_  &  n_n2997  &  wire7763 ) | ( pksi_132_  &  n_n2997  &  wire7763 ) ;
 assign wire1722 = ( (~ pksi_42_)  &  pksi_132_  &  n_n2993  &  wire7771 ) | ( pksi_42_  &  (~ pksi_132_)  &  n_n2993  &  wire7771 ) ;
 assign wire1727 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8251 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8251 ) ;
 assign wire1729 = ( pksi_124_  &  n_n2997  &  wire7763 ) | ( pksi_37_  &  n_n2997  &  wire7763 ) ;
 assign wire1730 = ( (~ pksi_124_)  &  pksi_37_  &  n_n2993  &  wire7771 ) | ( pksi_124_  &  (~ pksi_37_)  &  n_n2993  &  wire7771 ) ;
 assign wire1735 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8246 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8246 ) ;
 assign wire1737 = ( pksi_71_  &  n_n2997  &  wire7763 ) | ( pksi_150_  &  n_n2997  &  wire7763 ) ;
 assign wire1738 = ( (~ pksi_71_)  &  pksi_150_  &  n_n2993  &  wire7771 ) | ( pksi_71_  &  (~ pksi_150_)  &  n_n2993  &  wire7771 ) ;
 assign wire1743 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8241 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8241 ) ;
 assign wire1745 = ( pksi_70_  &  n_n2997  &  wire7763 ) | ( pksi_144_  &  n_n2997  &  wire7763 ) ;
 assign wire1746 = ( (~ pksi_70_)  &  pksi_144_  &  n_n2993  &  wire7771 ) | ( pksi_70_  &  (~ pksi_144_)  &  n_n2993  &  wire7771 ) ;
 assign wire1751 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8236 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8236 ) ;
 assign wire1753 = ( pksi_51_  &  n_n2997  &  wire7763 ) | ( pksi_145_  &  n_n2997  &  wire7763 ) ;
 assign wire1754 = ( (~ pksi_51_)  &  pksi_145_  &  n_n2993  &  wire7771 ) | ( pksi_51_  &  (~ pksi_145_)  &  n_n2993  &  wire7771 ) ;
 assign wire1759 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8231 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8231 ) ;
 assign wire1761 = ( pksi_82_  &  n_n2997  &  wire7763 ) | ( n_n2379  &  n_n2997  &  wire7763 ) ;
 assign wire1762 = ( (~ pksi_82_)  &  n_n2379  &  n_n2993  &  wire7771 ) | ( pksi_82_  &  (~ n_n2379)  &  n_n2993  &  wire7771 ) ;
 assign wire1765 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8226 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8226 ) ;
 assign wire1767 = ( pksi_119_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_15_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1768 = ( (~ pksi_119_)  &  pksi_15_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_119_  &  (~ pksi_15_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1771 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8221 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8221 ) ;
 assign wire1773 = ( pksi_92_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_173_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1774 = ( (~ pksi_92_)  &  pksi_173_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_92_  &  (~ pksi_173_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1777 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8216 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8216 ) ;
 assign wire1779 = ( pksi_111_  &  n_n2997  &  wire7763 ) | ( pksi_7_  &  n_n2997  &  wire7763 ) ;
 assign wire1780 = ( (~ pksi_111_)  &  pksi_7_  &  n_n2993  &  wire7771 ) | ( pksi_111_  &  (~ pksi_7_)  &  n_n2993  &  wire7771 ) ;
 assign wire1785 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8211 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8211 ) ;
 assign wire1787 = ( pksi_123_  &  n_n2997  &  wire7763 ) | ( n_n2821  &  n_n2997  &  wire7763 ) ;
 assign wire1788 = ( (~ pksi_123_)  &  n_n2821  &  n_n2993  &  wire7771 ) | ( pksi_123_  &  (~ n_n2821)  &  n_n2993  &  wire7771 ) ;
 assign wire1793 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8206 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8206 ) ;
 assign wire1795 = ( pksi_40_  &  n_n2997  &  wire7763 ) | ( n_n2931  &  n_n2997  &  wire7763 ) ;
 assign wire1796 = ( (~ pksi_40_)  &  n_n2931  &  n_n2993  &  wire7771 ) | ( pksi_40_  &  (~ n_n2931)  &  n_n2993  &  wire7771 ) ;
 assign wire1801 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8201 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8201 ) ;
 assign wire1803 = ( pksi_67_  &  n_n2997  &  wire7763 ) | ( n_n2921  &  n_n2997  &  wire7763 ) ;
 assign wire1804 = ( (~ pksi_67_)  &  n_n2921  &  n_n2993  &  wire7771 ) | ( pksi_67_  &  (~ n_n2921)  &  n_n2993  &  wire7771 ) ;
 assign wire1809 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8196 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8196 ) ;
 assign wire1811 = ( pksi_66_  &  n_n2997  &  wire7763 ) | ( pksi_156_  &  n_n2997  &  wire7763 ) ;
 assign wire1812 = ( (~ pksi_66_)  &  pksi_156_  &  n_n2993  &  wire7771 ) | ( pksi_66_  &  (~ pksi_156_)  &  n_n2993  &  wire7771 ) ;
 assign wire1817 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8191 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8191 ) ;
 assign wire1819 = ( pksi_161_  &  n_n2997  &  wire7763 ) | ( n_n2770  &  n_n2997  &  wire7763 ) ;
 assign wire1820 = ( (~ pksi_161_)  &  n_n2770  &  n_n2993  &  wire7771 ) | ( pksi_161_  &  (~ n_n2770)  &  n_n2993  &  wire7771 ) ;
 assign wire1825 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8186 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8186 ) ;
 assign wire1827 = ( pksi_93_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_179_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1828 = ( (~ pksi_93_)  &  pksi_179_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_93_  &  (~ pksi_179_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1831 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8181 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8181 ) ;
 assign wire1833 = ( pksi_101_  &  n_n2997  &  wire7763 ) | ( pksi_20_  &  n_n2997  &  wire7763 ) ;
 assign wire1834 = ( (~ pksi_101_)  &  pksi_20_  &  n_n2993  &  wire7771 ) | ( pksi_101_  &  (~ pksi_20_)  &  n_n2993  &  wire7771 ) ;
 assign wire1839 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8176 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8176 ) ;
 assign wire1841 = ( pksi_35_  &  n_n2997  &  wire7763 ) | ( n_n2950  &  n_n2997  &  wire7763 ) ;
 assign wire1842 = ( (~ pksi_35_)  &  n_n2950  &  n_n2993  &  wire7771 ) | ( pksi_35_  &  (~ n_n2950)  &  n_n2993  &  wire7771 ) ;
 assign wire1847 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8171 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8171 ) ;
 assign wire1849 = ( pksi_137_  &  n_n2997  &  wire7763 ) | ( n_n2802  &  n_n2997  &  wire7763 ) ;
 assign wire1850 = ( (~ pksi_137_)  &  n_n2802  &  n_n2993  &  wire7771 ) | ( pksi_137_  &  (~ n_n2802)  &  n_n2993  &  wire7771 ) ;
 assign wire1855 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8166 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8166 ) ;
 assign wire1857 = ( pksi_65_  &  n_n2997  &  wire7763 ) | ( pksi_165_  &  n_n2997  &  wire7763 ) ;
 assign wire1858 = ( (~ pksi_65_)  &  pksi_165_  &  n_n2993  &  wire7771 ) | ( pksi_65_  &  (~ pksi_165_)  &  n_n2993  &  wire7771 ) ;
 assign wire1863 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8161 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8161 ) ;
 assign wire1865 = ( pksi_56_  &  n_n2997  &  wire7763 ) | ( pksi_153_  &  n_n2997  &  wire7763 ) ;
 assign wire1866 = ( (~ pksi_56_)  &  pksi_153_  &  n_n2993  &  wire7771 ) | ( pksi_56_  &  (~ pksi_153_)  &  n_n2993  &  wire7771 ) ;
 assign wire1871 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8156 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8156 ) ;
 assign wire1873 = ( pksi_64_  &  n_n2997  &  wire7763 ) | ( n_n2899  &  n_n2997  &  wire7763 ) ;
 assign wire1874 = ( (~ pksi_64_)  &  n_n2899  &  n_n2993  &  wire7771 ) | ( pksi_64_  &  (~ n_n2899)  &  n_n2993  &  wire7771 ) ;
 assign wire1879 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8151 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8151 ) ;
 assign wire1881 = ( pksi_82_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2379  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1882 = ( (~ pksi_82_)  &  n_n2379  &  (~ n_n2993)  &  wire7765 ) | ( pksi_82_  &  (~ n_n2379)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1887 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8146 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8146 ) ;
 assign wire1889 = ( pksi_126_  &  n_n2997  &  wire7763 ) | ( pksi_47_  &  n_n2997  &  wire7763 ) ;
 assign wire1890 = ( (~ pksi_126_)  &  pksi_47_  &  n_n2993  &  wire7771 ) | ( pksi_126_  &  (~ pksi_47_)  &  n_n2993  &  wire7771 ) ;
 assign wire1895 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8141 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8141 ) ;
 assign wire1897 = ( pksi_26_  &  n_n2997  &  wire7763 ) | ( pksi_134_  &  n_n2997  &  wire7763 ) ;
 assign wire1898 = ( (~ pksi_26_)  &  pksi_134_  &  n_n2993  &  wire7771 ) | ( pksi_26_  &  (~ pksi_134_)  &  n_n2993  &  wire7771 ) ;
 assign wire1903 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8136 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8136 ) ;
 assign wire1905 = ( pksi_27_  &  n_n2997  &  wire7763 ) | ( pksi_121_  &  n_n2997  &  wire7763 ) ;
 assign wire1906 = ( (~ pksi_27_)  &  pksi_121_  &  n_n2993  &  wire7771 ) | ( pksi_27_  &  (~ pksi_121_)  &  n_n2993  &  wire7771 ) ;
 assign wire1911 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8131 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8131 ) ;
 assign wire1913 = ( pksi_53_  &  n_n2997  &  wire7763 ) | ( pksi_154_  &  n_n2997  &  wire7763 ) ;
 assign wire1914 = ( (~ pksi_53_)  &  pksi_154_  &  n_n2993  &  wire7771 ) | ( pksi_53_  &  (~ pksi_154_)  &  n_n2993  &  wire7771 ) ;
 assign wire1919 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8126 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8126 ) ;
 assign wire1921 = ( pksi_162_  &  n_n2997  &  wire7763 ) | ( n_n2779  &  n_n2997  &  wire7763 ) ;
 assign wire1922 = ( (~ pksi_162_)  &  n_n2779  &  n_n2993  &  wire7771 ) | ( pksi_162_  &  (~ n_n2779)  &  n_n2993  &  wire7771 ) ;
 assign wire1927 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8121 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8121 ) ;
 assign wire1929 = ( pksi_68_  &  n_n2997  &  wire7763 ) | ( pksi_149_  &  n_n2997  &  wire7763 ) ;
 assign wire1930 = ( (~ pksi_68_)  &  pksi_149_  &  n_n2993  &  wire7771 ) | ( pksi_68_  &  (~ pksi_149_)  &  n_n2993  &  wire7771 ) ;
 assign wire1935 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8116 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8116 ) ;
 assign wire1937 = ( pksi_188_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2741  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1938 = ( (~ pksi_188_)  &  n_n2741  &  (~ n_n2993)  &  wire7765 ) | ( pksi_188_  &  (~ n_n2741)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1943 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8111 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8111 ) ;
 assign wire1945 = ( pksi_142_  &  n_n2997  &  wire7763 ) | ( pksi_28_  &  n_n2997  &  wire7763 ) ;
 assign wire1946 = ( (~ pksi_142_)  &  pksi_28_  &  n_n2993  &  wire7771 ) | ( pksi_142_  &  (~ pksi_28_)  &  n_n2993  &  wire7771 ) ;
 assign wire1951 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8106 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8106 ) ;
 assign wire1953 = ( pksi_127_  &  n_n2997  &  wire7763 ) | ( pksi_38_  &  n_n2997  &  wire7763 ) ;
 assign wire1954 = ( (~ pksi_127_)  &  pksi_38_  &  n_n2993  &  wire7771 ) | ( pksi_127_  &  (~ pksi_38_)  &  n_n2993  &  wire7771 ) ;
 assign wire1959 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8101 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8101 ) ;
 assign wire1961 = ( pksi_128_  &  n_n2997  &  wire7763 ) | ( pksi_36_  &  n_n2997  &  wire7763 ) ;
 assign wire1962 = ( (~ pksi_128_)  &  pksi_36_  &  n_n2993  &  wire7771 ) | ( pksi_128_  &  (~ pksi_36_)  &  n_n2993  &  wire7771 ) ;
 assign wire1967 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8096 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8096 ) ;
 assign wire1969 = ( pksi_57_  &  n_n2997  &  wire7763 ) | ( pksi_160_  &  n_n2997  &  wire7763 ) ;
 assign wire1970 = ( (~ pksi_57_)  &  pksi_160_  &  n_n2993  &  wire7771 ) | ( pksi_57_  &  (~ pksi_160_)  &  n_n2993  &  wire7771 ) ;
 assign wire1975 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8091 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8091 ) ;
 assign wire1977 = ( pksi_49_  &  n_n2997  &  wire7763 ) | ( n_n2909  &  n_n2997  &  wire7763 ) ;
 assign wire1978 = ( (~ pksi_49_)  &  n_n2909  &  n_n2993  &  wire7771 ) | ( pksi_49_  &  (~ n_n2909)  &  n_n2993  &  wire7771 ) ;
 assign wire1983 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8086 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8086 ) ;
 assign wire1985 = ( pksi_55_  &  n_n2997  &  wire7763 ) | ( pksi_159_  &  n_n2997  &  wire7763 ) ;
 assign wire1986 = ( (~ pksi_55_)  &  pksi_159_  &  n_n2993  &  wire7771 ) | ( pksi_55_  &  (~ pksi_159_)  &  n_n2993  &  wire7771 ) ;
 assign wire1991 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8081 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8081 ) ;
 assign wire1993 = ( pksi_84_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_176_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire1994 = ( (~ pksi_84_)  &  pksi_176_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_84_  &  (~ pksi_176_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire1997 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8076 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8076 ) ;
 assign wire1999 = ( pksi_119_  &  n_n2997  &  wire7763 ) | ( pksi_15_  &  n_n2997  &  wire7763 ) ;
 assign wire2000 = ( (~ pksi_119_)  &  pksi_15_  &  n_n2993  &  wire7771 ) | ( pksi_119_  &  (~ pksi_15_)  &  n_n2993  &  wire7771 ) ;
 assign wire2005 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8071 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8071 ) ;
 assign wire2007 = ( pksi_96_  &  n_n2997  &  wire7763 ) | ( pksi_22_  &  n_n2997  &  wire7763 ) ;
 assign wire2008 = ( (~ pksi_96_)  &  pksi_22_  &  n_n2993  &  wire7771 ) | ( pksi_96_  &  (~ pksi_22_)  &  n_n2993  &  wire7771 ) ;
 assign wire2013 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8066 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8066 ) ;
 assign wire2015 = ( pksi_116_  &  n_n2997  &  wire7763 ) | ( n_n2838  &  n_n2997  &  wire7763 ) ;
 assign wire2016 = ( (~ pksi_116_)  &  n_n2838  &  n_n2993  &  wire7771 ) | ( pksi_116_  &  (~ n_n2838)  &  n_n2993  &  wire7771 ) ;
 assign wire2021 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8061 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8061 ) ;
 assign wire2023 = ( pksi_83_  &  n_n2997  &  wire7763 ) | ( n_n2885  &  n_n2997  &  wire7763 ) ;
 assign wire2024 = ( (~ pksi_83_)  &  n_n2885  &  n_n2993  &  wire7771 ) | ( pksi_83_  &  (~ n_n2885)  &  n_n2993  &  wire7771 ) ;
 assign wire2029 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8056 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8056 ) ;
 assign wire2031 = ( pksi_85_  &  n_n2997  &  wire7763 ) | ( pksi_172_  &  n_n2997  &  wire7763 ) ;
 assign wire2032 = ( (~ pksi_85_)  &  pksi_172_  &  n_n2993  &  wire7771 ) | ( pksi_85_  &  (~ pksi_172_)  &  n_n2993  &  wire7771 ) ;
 assign wire2035 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8051 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8051 ) ;
 assign wire2037 = ( pksi_183_  &  n_n2997  &  wire7763 ) | ( pksi_79_  &  n_n2997  &  wire7763 ) ;
 assign wire2038 = ( (~ pksi_183_)  &  pksi_79_  &  n_n2993  &  wire7771 ) | ( pksi_183_  &  (~ pksi_79_)  &  n_n2993  &  wire7771 ) ;
 assign wire2043 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8046 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8046 ) ;
 assign wire2045 = ( pksi_99_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2853  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2046 = ( (~ pksi_99_)  &  n_n2853  &  (~ n_n2993)  &  wire7765 ) | ( pksi_99_  &  (~ n_n2853)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2049 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8041 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8041 ) ;
 assign wire2051 = ( pksi_14_  &  n_n2997  &  wire7763 ) | ( pksi_103_  &  n_n2997  &  wire7763 ) ;
 assign wire2052 = ( (~ pksi_14_)  &  pksi_103_  &  n_n2993  &  wire7771 ) | ( pksi_14_  &  (~ pksi_103_)  &  n_n2993  &  wire7771 ) ;
 assign wire2055 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8036 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8036 ) ;
 assign wire2057 = ( pksi_12_  &  n_n2997  &  wire7763 ) | ( pksi_104_  &  n_n2997  &  wire7763 ) ;
 assign wire2058 = ( (~ pksi_12_)  &  pksi_104_  &  n_n2993  &  wire7771 ) | ( pksi_12_  &  (~ pksi_104_)  &  n_n2993  &  wire7771 ) ;
 assign wire2063 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8031 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8031 ) ;
 assign wire2065 = ( pksi_171_  &  n_n2997  &  wire7763 ) | ( n_n2757  &  n_n2997  &  wire7763 ) ;
 assign wire2066 = ( (~ pksi_171_)  &  n_n2757  &  n_n2993  &  wire7771 ) | ( pksi_171_  &  (~ n_n2757)  &  n_n2993  &  wire7771 ) ;
 assign wire2071 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8026 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8026 ) ;
 assign wire2073 = ( pksi_93_  &  n_n2997  &  wire7763 ) | ( pksi_179_  &  n_n2997  &  wire7763 ) ;
 assign wire2074 = ( (~ pksi_93_)  &  pksi_179_  &  n_n2993  &  wire7771 ) | ( pksi_93_  &  (~ pksi_179_)  &  n_n2993  &  wire7771 ) ;
 assign wire2079 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8021 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8021 ) ;
 assign wire2081 = ( pksi_92_  &  n_n2997  &  wire7763 ) | ( pksi_173_  &  n_n2997  &  wire7763 ) ;
 assign wire2082 = ( (~ pksi_92_)  &  pksi_173_  &  n_n2993  &  wire7771 ) | ( pksi_92_  &  (~ pksi_173_)  &  n_n2993  &  wire7771 ) ;
 assign wire2087 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8016 ) | ( (~ pstart_0_)  &  n_n2993  &  wire8016 ) ;
 assign wire2089 = ( pksi_11_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2982  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2090 = ( (~ pksi_11_)  &  n_n2982  &  (~ n_n2993)  &  wire7765 ) | ( pksi_11_  &  (~ n_n2982)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2093 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8011 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8011 ) ;
 assign wire2095 = ( pksi_102_  &  n_n2997  &  wire7763 ) | ( pksi_23_  &  n_n2997  &  wire7763 ) ;
 assign wire2096 = ( (~ pksi_102_)  &  pksi_23_  &  n_n2993  &  wire7771 ) | ( pksi_102_  &  (~ pksi_23_)  &  n_n2993  &  wire7771 ) ;
 assign wire2099 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8006 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8006 ) ;
 assign wire2101 = ( pksi_97_  &  n_n2997  &  wire7763 ) | ( pksi_3_  &  n_n2997  &  wire7763 ) ;
 assign wire2102 = ( (~ pksi_97_)  &  pksi_3_  &  n_n2993  &  wire7771 ) | ( pksi_97_  &  (~ pksi_3_)  &  n_n2993  &  wire7771 ) ;
 assign wire2107 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire8001 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire8001 ) ;
 assign wire2109 = ( pksi_16_  &  n_n2997  &  wire7763 ) | ( n_n2964  &  n_n2997  &  wire7763 ) ;
 assign wire2110 = ( (~ pksi_16_)  &  n_n2964  &  n_n2993  &  wire7771 ) | ( pksi_16_  &  (~ n_n2964)  &  n_n2993  &  wire7771 ) ;
 assign wire2115 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7996 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7996 ) ;
 assign wire2117 = ( pksi_43_  &  n_n2997  &  wire7763 ) | ( n_n2954  &  n_n2997  &  wire7763 ) ;
 assign wire2118 = ( (~ pksi_43_)  &  n_n2954  &  n_n2993  &  wire7771 ) | ( pksi_43_  &  (~ n_n2954)  &  n_n2993  &  wire7771 ) ;
 assign wire2123 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7991 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7991 ) ;
 assign wire2125 = ( pksi_189_  &  n_n2997  &  wire7763 ) | ( pksi_89_  &  n_n2997  &  wire7763 ) ;
 assign wire2126 = ( (~ pksi_189_)  &  pksi_89_  &  n_n2993  &  wire7771 ) | ( pksi_189_  &  (~ pksi_89_)  &  n_n2993  &  wire7771 ) ;
 assign wire2131 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7986 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7986 ) ;
 assign wire2133 = ( pksi_73_  &  n_n2997  &  wire7763 ) | ( pksi_177_  &  n_n2997  &  wire7763 ) ;
 assign wire2134 = ( (~ pksi_73_)  &  pksi_177_  &  n_n2993  &  wire7771 ) | ( pksi_73_  &  (~ pksi_177_)  &  n_n2993  &  wire7771 ) ;
 assign wire2139 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7981 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7981 ) ;
 assign wire2141 = ( pksi_102_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_23_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2142 = ( (~ pksi_102_)  &  pksi_23_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_102_  &  (~ pksi_23_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2147 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7976 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7976 ) ;
 assign wire2149 = ( pksi_110_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_2_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2150 = ( (~ pksi_110_)  &  pksi_2_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_110_  &  (~ pksi_2_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2153 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7971 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7971 ) ;
 assign wire2155 = ( pksi_98_  &  n_n2997  &  wire7763 ) | ( pksi_6_  &  n_n2997  &  wire7763 ) ;
 assign wire2156 = ( (~ pksi_98_)  &  pksi_6_  &  n_n2993  &  wire7771 ) | ( pksi_98_  &  (~ pksi_6_)  &  n_n2993  &  wire7771 ) ;
 assign wire2161 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7966 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7966 ) ;
 assign wire2163 = ( pksi_115_  &  n_n2997  &  wire7763 ) | ( pksi_0_  &  n_n2997  &  wire7763 ) ;
 assign wire2164 = ( (~ pksi_115_)  &  pksi_0_  &  n_n2993  &  wire7771 ) | ( pksi_115_  &  (~ pksi_0_)  &  n_n2993  &  wire7771 ) ;
 assign wire2169 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7961 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7961 ) ;
 assign wire2171 = ( pksi_113_  &  n_n2997  &  wire7763 ) | ( n_n2834  &  n_n2997  &  wire7763 ) ;
 assign wire2172 = ( (~ pksi_113_)  &  n_n2834  &  n_n2993  &  wire7771 ) | ( pksi_113_  &  (~ n_n2834)  &  n_n2993  &  wire7771 ) ;
 assign wire2177 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7956 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7956 ) ;
 assign wire2179 = ( pksi_41_  &  n_n2997  &  wire7763 ) | ( pksi_141_  &  n_n2997  &  wire7763 ) ;
 assign wire2180 = ( (~ pksi_41_)  &  pksi_141_  &  n_n2993  &  wire7771 ) | ( pksi_41_  &  (~ pksi_141_)  &  n_n2993  &  wire7771 ) ;
 assign wire2185 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7951 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7951 ) ;
 assign wire2187 = ( pksi_91_  &  n_n2997  &  wire7763 ) | ( n_n2889  &  n_n2997  &  wire7763 ) ;
 assign wire2188 = ( (~ pksi_91_)  &  n_n2889  &  n_n2993  &  wire7771 ) | ( pksi_91_  &  (~ n_n2889)  &  n_n2993  &  wire7771 ) ;
 assign wire2193 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7946 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7946 ) ;
 assign wire2195 = ( pksi_186_  &  n_n2997  &  wire7763 ) | ( n_n2746  &  n_n2997  &  wire7763 ) ;
 assign wire2196 = ( (~ pksi_186_)  &  n_n2746  &  n_n2993  &  wire7771 ) | ( pksi_186_  &  (~ n_n2746)  &  n_n2993  &  wire7771 ) ;
 assign wire2201 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7941 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7941 ) ;
 assign wire2203 = ( pksi_118_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_4_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2204 = ( (~ pksi_118_)  &  pksi_4_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_118_  &  (~ pksi_4_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2207 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7936 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7936 ) ;
 assign wire2209 = ( pksi_14_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_103_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2210 = ( (~ pksi_14_)  &  pksi_103_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_14_  &  (~ pksi_103_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2215 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7931 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7931 ) ;
 assign wire2217 = ( pksi_85_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_172_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2218 = ( (~ pksi_85_)  &  pksi_172_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_85_  &  (~ pksi_172_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2223 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7926 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7926 ) ;
 assign wire2225 = ( pksi_99_  &  n_n2997  &  wire7763 ) | ( n_n2853  &  n_n2997  &  wire7763 ) ;
 assign wire2226 = ( (~ pksi_99_)  &  n_n2853  &  n_n2993  &  wire7771 ) | ( pksi_99_  &  (~ n_n2853)  &  n_n2993  &  wire7771 ) ;
 assign wire2231 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7921 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7921 ) ;
 assign wire2233 = ( pksi_114_  &  n_n2997  &  wire7763 ) | ( n_n2843  &  n_n2997  &  wire7763 ) ;
 assign wire2234 = ( (~ pksi_114_)  &  n_n2843  &  n_n2993  &  wire7771 ) | ( pksi_114_  &  (~ n_n2843)  &  n_n2993  &  wire7771 ) ;
 assign wire2239 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7916 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7916 ) ;
 assign wire2241 = ( pksi_138_  &  n_n2997  &  wire7763 ) | ( n_n2811  &  n_n2997  &  wire7763 ) ;
 assign wire2242 = ( (~ pksi_138_)  &  n_n2811  &  n_n2993  &  wire7771 ) | ( pksi_138_  &  (~ n_n2811)  &  n_n2993  &  wire7771 ) ;
 assign wire2247 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7911 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7911 ) ;
 assign wire2249 = ( pksi_125_  &  n_n2997  &  wire7763 ) | ( pksi_44_  &  n_n2997  &  wire7763 ) ;
 assign wire2250 = ( (~ pksi_125_)  &  pksi_44_  &  n_n2993  &  wire7771 ) | ( pksi_125_  &  (~ pksi_44_)  &  n_n2993  &  wire7771 ) ;
 assign wire2255 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7906 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7906 ) ;
 assign wire2257 = ( pksi_81_  &  n_n2997  &  wire7763 ) | ( pksi_184_  &  n_n2997  &  wire7763 ) ;
 assign wire2258 = ( (~ pksi_81_)  &  pksi_184_  &  n_n2993  &  wire7771 ) | ( pksi_81_  &  (~ pksi_184_)  &  n_n2993  &  wire7771 ) ;
 assign wire2263 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7901 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7901 ) ;
 assign wire2265 = ( pksi_80_  &  n_n2997  &  wire7763 ) | ( n_n2877  &  n_n2997  &  wire7763 ) ;
 assign wire2266 = ( (~ pksi_80_)  &  n_n2877  &  n_n2993  &  wire7771 ) | ( pksi_80_  &  (~ n_n2877)  &  n_n2993  &  wire7771 ) ;
 assign wire2271 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7896 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7896 ) ;
 assign wire2273 = ( pksi_75_  &  n_n2997  &  wire7763 ) | ( pksi_169_  &  n_n2997  &  wire7763 ) ;
 assign wire2274 = ( (~ pksi_75_)  &  pksi_169_  &  n_n2993  &  wire7771 ) | ( pksi_75_  &  (~ pksi_169_)  &  n_n2993  &  wire7771 ) ;
 assign wire2279 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7891 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7891 ) ;
 assign wire2281 = ( pksi_106_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_5_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2282 = ( (~ pksi_106_)  &  pksi_5_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_106_  &  (~ pksi_5_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2287 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7886 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7886 ) ;
 assign wire2289 = ( pksi_118_  &  n_n2997  &  wire7763 ) | ( pksi_4_  &  n_n2997  &  wire7763 ) ;
 assign wire2290 = ( (~ pksi_118_)  &  pksi_4_  &  n_n2993  &  wire7771 ) | ( pksi_118_  &  (~ pksi_4_)  &  n_n2993  &  wire7771 ) ;
 assign wire2295 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7881 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7881 ) ;
 assign wire2297 = ( pksi_117_  &  n_n2997  &  wire7763 ) | ( pksi_17_  &  n_n2997  &  wire7763 ) ;
 assign wire2298 = ( (~ pksi_117_)  &  pksi_17_  &  n_n2993  &  wire7771 ) | ( pksi_117_  &  (~ pksi_17_)  &  n_n2993  &  wire7771 ) ;
 assign wire2301 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7876 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7876 ) ;
 assign wire2303 = ( pksi_100_  &  n_n2997  &  wire7763 ) | ( pksi_13_  &  n_n2997  &  wire7763 ) ;
 assign wire2304 = ( (~ pksi_100_)  &  pksi_13_  &  n_n2993  &  wire7771 ) | ( pksi_100_  &  (~ pksi_13_)  &  n_n2993  &  wire7771 ) ;
 assign wire2309 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7871 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7871 ) ;
 assign wire2311 = ( pksi_129_  &  n_n2997  &  wire7763 ) | ( pksi_25_  &  n_n2997  &  wire7763 ) ;
 assign wire2312 = ( (~ pksi_129_)  &  pksi_25_  &  n_n2993  &  wire7771 ) | ( pksi_129_  &  (~ pksi_25_)  &  n_n2993  &  wire7771 ) ;
 assign wire2317 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7866 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7866 ) ;
 assign wire2319 = ( pksi_31_  &  n_n2997  &  wire7763 ) | ( pksi_135_  &  n_n2997  &  wire7763 ) ;
 assign wire2320 = ( (~ pksi_31_)  &  pksi_135_  &  n_n2993  &  wire7771 ) | ( pksi_31_  &  (~ pksi_135_)  &  n_n2993  &  wire7771 ) ;
 assign wire2325 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7861 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7861 ) ;
 assign wire2327 = ( pksi_77_  &  n_n2997  &  wire7763 ) | ( pksi_178_  &  n_n2997  &  wire7763 ) ;
 assign wire2328 = ( (~ pksi_77_)  &  pksi_178_  &  n_n2993  &  wire7771 ) | ( pksi_77_  &  (~ pksi_178_)  &  n_n2993  &  wire7771 ) ;
 assign wire2333 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7856 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7856 ) ;
 assign wire2335 = ( pksi_180_  &  n_n2997  &  wire7763 ) | ( n_n2749  &  n_n2997  &  wire7763 ) ;
 assign wire2336 = ( (~ pksi_180_)  &  n_n2749  &  n_n2993  &  wire7771 ) | ( pksi_180_  &  (~ n_n2749)  &  n_n2993  &  wire7771 ) ;
 assign wire2341 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7851 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7851 ) ;
 assign wire2343 = ( pksi_84_  &  n_n2997  &  wire7763 ) | ( pksi_176_  &  n_n2997  &  wire7763 ) ;
 assign wire2344 = ( (~ pksi_84_)  &  pksi_176_  &  n_n2993  &  wire7771 ) | ( pksi_84_  &  (~ pksi_176_)  &  n_n2993  &  wire7771 ) ;
 assign wire2349 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7846 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7846 ) ;
 assign wire2351 = ( pksi_112_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_9_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2352 = ( (~ pksi_112_)  &  pksi_9_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_112_  &  (~ pksi_9_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2357 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7841 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7841 ) ;
 assign wire2359 = ( pksi_110_  &  n_n2997  &  wire7763 ) | ( pksi_2_  &  n_n2997  &  wire7763 ) ;
 assign wire2360 = ( (~ pksi_110_)  &  pksi_2_  &  n_n2993  &  wire7771 ) | ( pksi_110_  &  (~ pksi_2_)  &  n_n2993  &  wire7771 ) ;
 assign wire2365 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7836 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7836 ) ;
 assign wire2367 = ( pksi_107_  &  n_n2997  &  wire7763 ) | ( pksi_21_  &  n_n2997  &  wire7763 ) ;
 assign wire2368 = ( (~ pksi_107_)  &  pksi_21_  &  n_n2993  &  wire7771 ) | ( pksi_107_  &  (~ pksi_21_)  &  n_n2993  &  wire7771 ) ;
 assign wire2373 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7831 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7831 ) ;
 assign wire2375 = ( pksi_59_  &  n_n2997  &  wire7763 ) | ( n_n2917  &  n_n2997  &  wire7763 ) ;
 assign wire2376 = ( (~ pksi_59_)  &  n_n2917  &  n_n2993  &  wire7771 ) | ( pksi_59_  &  (~ n_n2917)  &  n_n2993  &  wire7771 ) ;
 assign wire2381 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7826 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7826 ) ;
 assign wire2383 = ( pksi_61_  &  n_n2997  &  wire7763 ) | ( pksi_148_  &  n_n2997  &  wire7763 ) ;
 assign wire2384 = ( (~ pksi_61_)  &  pksi_148_  &  n_n2993  &  wire7771 ) | ( pksi_61_  &  (~ pksi_148_)  &  n_n2993  &  wire7771 ) ;
 assign wire2389 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7821 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7821 ) ;
 assign wire2391 = ( pksi_87_  &  n_n2997  &  wire7763 ) | ( n_n2391  &  n_n2997  &  wire7763 ) ;
 assign wire2392 = ( (~ pksi_87_)  &  n_n2391  &  n_n2993  &  wire7771 ) | ( pksi_87_  &  (~ n_n2391)  &  n_n2993  &  wire7771 ) ;
 assign wire2397 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7816 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7816 ) ;
 assign wire2399 = ( pksi_94_  &  n_n2997  &  wire7763 ) | ( n_n2881  &  n_n2997  &  wire7763 ) ;
 assign wire2400 = ( (~ pksi_94_)  &  n_n2881  &  n_n2993  &  wire7771 ) | ( pksi_94_  &  (~ n_n2881)  &  n_n2993  &  wire7771 ) ;
 assign wire2405 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7811 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7811 ) ;
 assign wire2407 = ( n_n2865  &  n_n2997  &  wire7763 ) | ( n_n2280  &  n_n2997  &  wire7763 ) ;
 assign wire2408 = ( (~ n_n2865)  &  n_n2280  &  n_n2993  &  wire7771 ) | ( n_n2865  &  (~ n_n2280)  &  n_n2993  &  wire7771 ) ;
 assign wire2413 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7806 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7806 ) ;
 assign wire2415 = ( pksi_19_  &  (~ n_n2997)  &  wire7764 ) | ( n_n2986  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2416 = ( (~ pksi_19_)  &  n_n2986  &  (~ n_n2993)  &  wire7765 ) | ( pksi_19_  &  (~ n_n2986)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire2421 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7801 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7801 ) ;
 assign wire2423 = ( pksi_11_  &  n_n2997  &  wire7763 ) | ( n_n2982  &  n_n2997  &  wire7763 ) ;
 assign wire2424 = ( (~ pksi_11_)  &  n_n2982  &  n_n2993  &  wire7771 ) | ( pksi_11_  &  (~ n_n2982)  &  n_n2993  &  wire7771 ) ;
 assign wire2429 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7796 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7796 ) ;
 assign wire2431 = ( pksi_109_  &  n_n2997  &  wire7763 ) | ( pksi_10_  &  n_n2997  &  wire7763 ) ;
 assign wire2432 = ( (~ pksi_109_)  &  pksi_10_  &  n_n2993  &  wire7771 ) | ( pksi_109_  &  (~ pksi_10_)  &  n_n2993  &  wire7771 ) ;
 assign wire2437 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7791 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7791 ) ;
 assign wire2439 = ( pksi_147_  &  n_n2997  &  wire7763 ) | ( n_n2789  &  n_n2997  &  wire7763 ) ;
 assign wire2440 = ( (~ pksi_147_)  &  n_n2789  &  n_n2993  &  wire7771 ) | ( pksi_147_  &  (~ n_n2789)  &  n_n2993  &  wire7771 ) ;
 assign wire2445 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7786 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7786 ) ;
 assign wire2447 = ( pksi_69_  &  n_n2997  &  wire7763 ) | ( pksi_155_  &  n_n2997  &  wire7763 ) ;
 assign wire2448 = ( (~ pksi_69_)  &  pksi_155_  &  n_n2993  &  wire7771 ) | ( pksi_69_  &  (~ pksi_155_)  &  n_n2993  &  wire7771 ) ;
 assign wire2453 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7781 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7781 ) ;
 assign wire2455 = ( pksi_170_  &  n_n2997  &  wire7763 ) | ( pksi_78_  &  n_n2997  &  wire7763 ) ;
 assign wire2456 = ( (~ pksi_170_)  &  pksi_78_  &  n_n2993  &  wire7771 ) | ( pksi_170_  &  (~ pksi_78_)  &  n_n2993  &  wire7771 ) ;
 assign wire2461 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7776 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7776 ) ;
 assign wire2463 = ( pksi_72_  &  n_n2997  &  wire7763 ) | ( n_n2879  &  n_n2997  &  wire7763 ) ;
 assign wire2464 = ( (~ pksi_72_)  &  n_n2879  &  n_n2993  &  wire7771 ) | ( pksi_72_  &  (~ n_n2879)  &  n_n2993  &  wire7771 ) ;
 assign wire2469 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7770 ) | ( (~ pstart_0_)  &  (~ n_n2993)  &  wire7770 ) ;
 assign wire2471 = ( pksi_185_  &  n_n2997  &  wire7763 ) | ( n_n2737  &  n_n2997  &  wire7763 ) ;
 assign wire2472 = ( (~ pksi_185_)  &  n_n2737  &  n_n2993  &  wire7771 ) | ( pksi_185_  &  (~ n_n2737)  &  n_n2993  &  wire7771 ) ;
 assign wire2477 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  wire7760 ) | ( (~ pstart_0_)  &  n_n2993  &  wire7760 ) ;
 assign wire2479 = ( pksi_117_  &  (~ n_n2997)  &  wire7764 ) | ( pksi_17_  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire2480 = ( (~ pksi_117_)  &  pksi_17_  &  (~ n_n2993)  &  wire7765 ) | ( pksi_117_  &  (~ pksi_17_)  &  (~ n_n2993)  &  wire7765 ) ;
 assign wire7760 = ( pksi_17_  &  pksi_117_ ) ;
 assign wire7763 = ( (~ pencrypt_0_)  &  (~ pstart_0_) ) ;
 assign wire7764 = ( (~ pencrypt_0_)  &  (~ pstart_0_) ) ;
 assign wire7765 = ( pencrypt_0_  &  (~ pstart_0_) ) ;
 assign wire7766 = ( pkey_57_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_0_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7767 = ( wire7766 ) | ( (~ wire775)  &  n_n2997  &  wire7763 ) ;
 assign wire7770 = ( n_n2737  &  pksi_185_ ) ;
 assign wire7771 = ( pencrypt_0_  &  (~ pstart_0_) ) ;
 assign wire7772 = ( pkey_211_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_219_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7773 = ( wire7772 ) | ( (~ wire776)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7776 = ( n_n2879  &  pksi_72_ ) ;
 assign wire7777 = ( pkey_213_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_205_ ) ;
 assign wire7778 = ( wire7777 ) | ( (~ wire777)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7781 = ( pksi_78_  &  pksi_170_ ) ;
 assign wire7782 = ( pkey_230_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_238_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7783 = ( wire7782 ) | ( (~ wire778)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7786 = ( pksi_155_  &  pksi_69_ ) ;
 assign wire7787 = ( pkey_156_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_164_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7788 = ( wire7787 ) | ( (~ wire779)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7791 = ( n_n2789  &  pksi_147_ ) ;
 assign wire7792 = ( pstart_0_  &  pkey_181_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_189_ ) ;
 assign wire7793 = ( wire7792 ) | ( (~ wire780)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7796 = ( pksi_10_  &  pksi_109_ ) ;
 assign wire7797 = ( pkey_28_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_20_ ) ;
 assign wire7798 = ( wire7797 ) | ( (~ wire781)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7801 = ( n_n2982  &  pksi_11_ ) ;
 assign wire7802 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_53_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_45_ ) ;
 assign wire7803 = ( wire7802 ) | ( (~ wire782)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7806 = ( n_n2986  &  pksi_19_ ) ;
 assign wire7807 = ( pkey_0_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_8_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7808 = ( wire7807 ) | ( n_n2997  &  (~ wire793)  &  wire7763 ) ;
 assign wire7811 = ( n_n2280  &  n_n2865 ) ;
 assign wire7812 = ( pstart_0_  &  pkey_203_  &  pencrypt_0_ ) | ( pkey_211_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7813 = ( wire7812 ) | ( (~ n_n2997)  &  (~ wire794)  &  wire7764 ) ;
 assign wire7816 = ( n_n2881  &  pksi_94_ ) ;
 assign wire7817 = ( pkey_213_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_221_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7818 = ( wire7817 ) | ( (~ n_n2997)  &  (~ wire784)  &  wire7764 ) ;
 assign wire7821 = ( n_n2391  &  pksi_87_ ) ;
 assign wire7822 = ( pkey_222_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_230_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7823 = ( wire7822 ) | ( (~ n_n2997)  &  (~ wire795)  &  wire7764 ) ;
 assign wire7826 = ( pksi_148_  &  pksi_61_ ) ;
 assign wire7827 = ( pkey_164_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_172_ ) ;
 assign wire7828 = ( wire7827 ) | ( (~ n_n2997)  &  (~ wire786)  &  wire7764 ) ;
 assign wire7831 = ( n_n2917  &  pksi_59_ ) ;
 assign wire7832 = ( pstart_0_  &  pkey_181_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_173_ ) ;
 assign wire7833 = ( wire7832 ) | ( (~ n_n2997)  &  (~ wire796)  &  wire7764 ) ;
 assign wire7836 = ( pksi_21_  &  pksi_107_ ) ;
 assign wire7837 = ( pkey_28_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_36_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7838 = ( wire7837 ) | ( (~ n_n2997)  &  (~ wire797)  &  wire7764 ) ;
 assign wire7841 = ( pksi_2_  &  pksi_110_ ) ;
 assign wire7842 = ( pkey_37_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_45_ ) ;
 assign wire7843 = ( wire7842 ) | ( (~ n_n2997)  &  (~ wire798)  &  wire7764 ) ;
 assign wire7846 = ( pksi_9_  &  pksi_112_ ) ;
 assign wire7847 = ( pkey_8_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_16_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7848 = ( wire7847 ) | ( n_n2997  &  (~ wire809)  &  wire7763 ) ;
 assign wire7851 = ( pksi_176_  &  pksi_84_ ) ;
 assign wire7852 = ( pstart_0_  &  pkey_196_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_204_ ) ;
 assign wire7853 = ( wire7852 ) | ( (~ n_n2997)  &  (~ wire799)  &  wire7764 ) ;
 assign wire7856 = ( n_n2749  &  pksi_180_ ) ;
 assign wire7857 = ( pkey_252_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_197_  &  (~ pencrypt_0_) ) ;
 assign wire7858 = ( wire7857 ) | ( (~ n_n2997)  &  (~ wire810)  &  wire7764 ) ;
 assign wire7861 = ( pksi_178_  &  pksi_77_ ) ;
 assign wire7862 = ( pkey_214_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_222_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7863 = ( wire7862 ) | ( (~ n_n2997)  &  (~ wire811)  &  wire7764 ) ;
 assign wire7866 = ( pksi_135_  &  pksi_31_ ) ;
 assign wire7867 = ( pkey_67_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_190_ ) ;
 assign wire7868 = ( wire7867 ) | ( (~ n_n2997)  &  (~ wire812)  &  wire7764 ) ;
 assign wire7871 = ( pksi_25_  &  pksi_129_ ) ;
 assign wire7872 = ( pkey_116_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_124_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7873 = ( wire7872 ) | ( (~ n_n2997)  &  (~ wire806)  &  wire7764 ) ;
 assign wire7876 = ( pksi_13_  &  pksi_100_ ) ;
 assign wire7877 = ( pkey_36_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_44_ ) ;
 assign wire7878 = ( wire7877 ) | ( (~ n_n2997)  &  (~ wire808)  &  wire7764 ) ;
 assign wire7881 = ( pksi_17_  &  pksi_117_ ) ;
 assign wire7882 = ( pkey_61_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_6_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7883 = ( wire7882 ) | ( (~ wire775)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire7886 = ( pksi_4_  &  pksi_118_ ) ;
 assign wire7887 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_62_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_54_ ) ;
 assign wire7888 = ( wire7887 ) | ( (~ n_n2997)  &  (~ wire813)  &  wire7764 ) ;
 assign wire7891 = ( pksi_5_  &  pksi_106_ ) ;
 assign wire7892 = ( pkey_16_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_24_ ) ;
 assign wire7893 = ( wire7892 ) | ( n_n2997  &  (~ wire821)  &  wire7763 ) ;
 assign wire7896 = ( pksi_169_  &  pksi_75_ ) ;
 assign wire7897 = ( pkey_219_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_196_  &  (~ pencrypt_0_) ) ;
 assign wire7898 = ( wire7897 ) | ( (~ n_n2997)  &  (~ wire822)  &  wire7764 ) ;
 assign wire7901 = ( n_n2877  &  pksi_80_ ) ;
 assign wire7902 = ( pstart_0_  &  pkey_197_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_205_ ) ;
 assign wire7903 = ( wire7902 ) | ( (~ n_n2997)  &  (~ wire823)  &  wire7764 ) ;
 assign wire7906 = ( pksi_184_  &  pksi_81_ ) ;
 assign wire7907 = ( pkey_206_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_214_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7908 = ( wire7907 ) | ( (~ n_n2997)  &  (~ wire824)  &  wire7764 ) ;
 assign wire7911 = ( pksi_44_  &  pksi_125_ ) ;
 assign wire7912 = ( pkey_67_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_75_ ) ;
 assign wire7913 = ( wire7912 ) | ( (~ n_n2997)  &  (~ wire825)  &  wire7764 ) ;
 assign wire7916 = ( n_n2811  &  pksi_138_ ) ;
 assign wire7917 = ( pkey_116_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_44_ ) ;
 assign wire7918 = ( wire7917 ) | ( (~ n_n2997)  &  (~ wire826)  &  wire7764 ) ;
 assign wire7921 = ( n_n2843  &  pksi_114_ ) ;
 assign wire7922 = ( pstart_0_  &  pkey_52_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_44_ ) ;
 assign wire7923 = ( wire7922 ) | ( (~ n_n2997)  &  (~ wire790)  &  wire7764 ) ;
 assign wire7926 = ( n_n2853  &  pksi_99_ ) ;
 assign wire7927 = ( pkey_61_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_53_ ) ;
 assign wire7928 = ( wire7927 ) | ( (~ n_n2997)  &  (~ wire827)  &  wire7764 ) ;
 assign wire7931 = ( pksi_172_  &  pksi_85_ ) ;
 assign wire7932 = ( pkey_226_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_234_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7933 = ( wire7932 ) | ( n_n2997  &  (~ wire834)  &  wire7763 ) ;
 assign wire7936 = ( pksi_103_  &  pksi_14_ ) ;
 assign wire7937 = ( pstart_0_  &  pencrypt_0_  &  pkey_25_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_33_ ) ;
 assign wire7938 = ( wire7937 ) | ( n_n2997  &  (~ wire835)  &  wire7763 ) ;
 assign wire7941 = ( pksi_4_  &  pksi_118_ ) ;
 assign wire7942 = ( pkey_48_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_56_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7943 = ( wire7942 ) | ( n_n2997  &  (~ wire813)  &  wire7763 ) ;
 assign wire7946 = ( n_n2746  &  pksi_186_ ) ;
 assign wire7947 = ( pkey_244_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_172_ ) ;
 assign wire7948 = ( wire7947 ) | ( (~ n_n2997)  &  (~ wire836)  &  wire7764 ) ;
 assign wire7951 = ( n_n2889  &  pksi_91_ ) ;
 assign wire7952 = ( pkey_206_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_198_ ) ;
 assign wire7953 = ( wire7952 ) | ( (~ n_n2997)  &  (~ wire837)  &  wire7764 ) ;
 assign wire7956 = ( pksi_141_  &  pksi_41_ ) ;
 assign wire7957 = ( pkey_125_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_70_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7958 = ( wire7957 ) | ( (~ n_n2997)  &  (~ wire838)  &  wire7764 ) ;
 assign wire7961 = ( n_n2834  &  pksi_113_ ) ;
 assign wire7962 = ( pkey_19_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_27_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7963 = ( wire7962 ) | ( (~ n_n2997)  &  (~ wire839)  &  wire7764 ) ;
 assign wire7966 = ( pksi_0_  &  pksi_115_ ) ;
 assign wire7967 = ( pstart_0_  &  pencrypt_0_  &  pkey_13_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_21_ ) ;
 assign wire7968 = ( wire7967 ) | ( (~ n_n2997)  &  (~ wire840)  &  wire7764 ) ;
 assign wire7971 = ( pksi_6_  &  pksi_98_ ) ;
 assign wire7972 = ( pkey_38_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_46_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7973 = ( wire7972 ) | ( (~ n_n2997)  &  (~ wire841)  &  wire7764 ) ;
 assign wire7976 = ( pksi_2_  &  pksi_110_ ) ;
 assign wire7977 = ( pstart_0_  &  pencrypt_0_  &  pkey_33_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_41_ ) ;
 assign wire7978 = ( wire7977 ) | ( n_n2997  &  (~ wire798)  &  wire7763 ) ;
 assign wire7981 = ( pksi_23_  &  pksi_102_ ) ;
 assign wire7982 = ( pkey_48_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_40_ ) ;
 assign wire7983 = ( wire7982 ) | ( n_n2997  &  (~ wire846)  &  wire7763 ) ;
 assign wire7986 = ( pksi_177_  &  pksi_73_ ) ;
 assign wire7987 = ( pkey_244_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_252_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7988 = ( wire7987 ) | ( (~ n_n2997)  &  (~ wire847)  &  wire7764 ) ;
 assign wire7991 = ( pksi_89_  &  pksi_189_ ) ;
 assign wire7992 = ( pkey_253_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_198_ ) ;
 assign wire7993 = ( wire7992 ) | ( (~ n_n2997)  &  (~ wire848)  &  wire7764 ) ;
 assign wire7996 = ( n_n2954  &  pksi_43_ ) ;
 assign wire7997 = ( pkey_70_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_78_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7998 = ( wire7997 ) | ( (~ n_n2997)  &  (~ wire843)  &  wire7764 ) ;
 assign wire8001 = ( n_n2964  &  pksi_16_ ) ;
 assign wire8002 = ( pkey_19_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_11_ ) ;
 assign wire8003 = ( wire8002 ) | ( (~ n_n2997)  &  (~ wire849)  &  wire7764 ) ;
 assign wire8006 = ( pksi_3_  &  pksi_97_ ) ;
 assign wire8007 = ( pkey_27_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_4_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8008 = ( wire8007 ) | ( (~ n_n2997)  &  (~ wire850)  &  wire7764 ) ;
 assign wire8011 = ( pksi_23_  &  pksi_102_ ) ;
 assign wire8012 = ( pkey_46_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_54_ ) ;
 assign wire8013 = ( wire8012 ) | ( (~ n_n2997)  &  (~ wire846)  &  wire7764 ) ;
 assign wire8016 = ( n_n2982  &  pksi_11_ ) ;
 assign wire8017 = ( pkey_49_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_41_ ) ;
 assign wire8018 = ( wire8017 ) | ( (~ wire782)  &  n_n2997  &  wire7763 ) ;
 assign wire8021 = ( pksi_173_  &  pksi_92_ ) ;
 assign wire8022 = ( pkey_195_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_203_  &  (~ pencrypt_0_) ) ;
 assign wire8023 = ( wire8022 ) | ( (~ n_n2997)  &  (~ wire851)  &  wire7764 ) ;
 assign wire8026 = ( pksi_179_  &  pksi_93_ ) ;
 assign wire8027 = ( pkey_220_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_228_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8028 = ( wire8027 ) | ( (~ n_n2997)  &  (~ wire814)  &  wire7764 ) ;
 assign wire8031 = ( n_n2757  &  pksi_171_ ) ;
 assign wire8032 = ( pkey_245_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_253_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8033 = ( wire8032 ) | ( (~ n_n2997)  &  (~ wire852)  &  wire7764 ) ;
 assign wire8036 = ( pksi_104_  &  pksi_12_ ) ;
 assign wire8037 = ( pkey_4_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_12_ ) ;
 assign wire8038 = ( wire8037 ) | ( (~ n_n2997)  &  (~ wire853)  &  wire7764 ) ;
 assign wire8041 = ( pksi_103_  &  pksi_14_ ) ;
 assign wire8042 = ( pkey_29_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_37_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8043 = ( wire8042 ) | ( (~ n_n2997)  &  (~ wire835)  &  wire7764 ) ;
 assign wire8046 = ( n_n2853  &  pksi_99_ ) ;
 assign wire8047 = ( pkey_49_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_57_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8048 = ( wire8047 ) | ( n_n2997  &  (~ wire827)  &  wire7763 ) ;
 assign wire8051 = ( pksi_79_  &  pksi_183_ ) ;
 assign wire8052 = ( pkey_195_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_62_ ) ;
 assign wire8053 = ( wire8052 ) | ( (~ n_n2997)  &  (~ wire855)  &  wire7764 ) ;
 assign wire8056 = ( pksi_172_  &  pksi_85_ ) ;
 assign wire8057 = ( pkey_228_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_172_ ) ;
 assign wire8058 = ( wire8057 ) | ( (~ n_n2997)  &  (~ wire834)  &  wire7764 ) ;
 assign wire8061 = ( n_n2885  &  pksi_83_ ) ;
 assign wire8062 = ( pkey_237_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_245_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8063 = ( wire8062 ) | ( (~ n_n2997)  &  (~ wire829)  &  wire7764 ) ;
 assign wire8066 = ( n_n2838  &  pksi_116_ ) ;
 assign wire8067 = ( pstart_0_  &  pencrypt_0_  &  pkey_12_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_20_ ) ;
 assign wire8068 = ( wire8067 ) | ( (~ n_n2997)  &  (~ wire856)  &  wire7764 ) ;
 assign wire8071 = ( pksi_22_  &  pksi_96_ ) ;
 assign wire8072 = ( pkey_29_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_21_ ) ;
 assign wire8073 = ( wire8072 ) | ( (~ n_n2997)  &  (~ wire857)  &  wire7764 ) ;
 assign wire8076 = ( pksi_15_  &  pksi_119_ ) ;
 assign wire8077 = ( pkey_38_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_30_ ) ;
 assign wire8078 = ( wire8077 ) | ( (~ n_n2997)  &  (~ wire858)  &  wire7764 ) ;
 assign wire8081 = ( pksi_176_  &  pksi_84_ ) ;
 assign wire8082 = ( pkey_194_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_202_ ) ;
 assign wire8083 = ( wire8082 ) | ( n_n2997  &  (~ wire799)  &  wire7763 ) ;
 assign wire8086 = ( pksi_159_  &  pksi_55_ ) ;
 assign wire8087 = ( pkey_254_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_131_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8088 = ( wire8087 ) | ( (~ n_n2997)  &  (~ wire816)  &  wire7764 ) ;
 assign wire8091 = ( n_n2909  &  pksi_49_ ) ;
 assign wire8092 = ( pkey_180_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_188_ ) ;
 assign wire8093 = ( wire8092 ) | ( (~ n_n2997)  &  (~ wire861)  &  wire7764 ) ;
 assign wire8096 = ( pksi_160_  &  pksi_57_ ) ;
 assign wire8097 = ( pkey_142_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_150_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8098 = ( wire8097 ) | ( (~ n_n2997)  &  (~ wire862)  &  wire7764 ) ;
 assign wire8101 = ( pksi_36_  &  pksi_128_ ) ;
 assign wire8102 = ( pkey_68_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_76_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8103 = ( wire8102 ) | ( (~ n_n2997)  &  (~ wire818)  &  wire7764 ) ;
 assign wire8106 = ( pksi_38_  &  pksi_127_ ) ;
 assign wire8107 = ( pkey_93_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_101_ ) ;
 assign wire8108 = ( wire8107 ) | ( (~ n_n2997)  &  (~ wire863)  &  wire7764 ) ;
 assign wire8111 = ( pksi_28_  &  pksi_142_ ) ;
 assign wire8112 = ( pkey_118_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_126_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8113 = ( wire8112 ) | ( (~ n_n2997)  &  (~ wire819)  &  wire7764 ) ;
 assign wire8116 = ( n_n2741  &  pksi_188_ ) ;
 assign wire8117 = ( pkey_210_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_202_ ) ;
 assign wire8118 = ( wire8117 ) | ( (~ wire783)  &  n_n2997  &  wire7763 ) ;
 assign wire8121 = ( pksi_149_  &  pksi_68_ ) ;
 assign wire8122 = ( pkey_131_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_139_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8123 = ( wire8122 ) | ( (~ n_n2997)  &  (~ wire865)  &  wire7764 ) ;
 assign wire8126 = ( n_n2779  &  pksi_162_ ) ;
 assign wire8127 = ( pkey_180_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_172_ ) ;
 assign wire8128 = ( wire8127 ) | ( (~ n_n2997)  &  (~ wire801)  &  wire7764 ) ;
 assign wire8131 = ( pksi_154_  &  pksi_53_ ) ;
 assign wire8132 = ( pkey_150_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_158_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8133 = ( wire8132 ) | ( (~ n_n2997)  &  (~ wire866)  &  wire7764 ) ;
 assign wire8136 = ( pksi_121_  &  pksi_27_ ) ;
 assign wire8137 = ( pkey_68_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_91_ ) ;
 assign wire8138 = ( wire8137 ) | ( (~ n_n2997)  &  (~ wire802)  &  wire7764 ) ;
 assign wire8141 = ( pksi_134_  &  pksi_26_ ) ;
 assign wire8142 = ( pstart_0_  &  pkey_109_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_101_ ) ;
 assign wire8143 = ( wire8142 ) | ( (~ n_n2997)  &  (~ wire867)  &  wire7764 ) ;
 assign wire8146 = ( pksi_47_  &  pksi_126_ ) ;
 assign wire8147 = ( pkey_110_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_118_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8148 = ( wire8147 ) | ( (~ n_n2997)  &  (~ wire807)  &  wire7764 ) ;
 assign wire8151 = ( n_n2379  &  pksi_82_ ) ;
 assign wire8152 = ( pkey_210_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_218_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8153 = ( wire8152 ) | ( n_n2997  &  (~ wire828)  &  wire7763 ) ;
 assign wire8156 = ( n_n2899  &  pksi_64_ ) ;
 assign wire8157 = ( pkey_139_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_147_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8158 = ( wire8157 ) | ( (~ n_n2997)  &  (~ wire871)  &  wire7764 ) ;
 assign wire8161 = ( pksi_153_  &  pksi_56_ ) ;
 assign wire8162 = ( pkey_133_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_141_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8163 = ( wire8162 ) | ( (~ n_n2997)  &  (~ wire872)  &  wire7764 ) ;
 assign wire8166 = ( pksi_165_  &  pksi_65_ ) ;
 assign wire8167 = ( pkey_134_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_189_ ) ;
 assign wire8168 = ( wire8167 ) | ( (~ n_n2997)  &  (~ wire787)  &  wire7764 ) ;
 assign wire8171 = ( n_n2802  &  pksi_137_ ) ;
 assign wire8172 = ( pstart_0_  &  pencrypt_0_  &  pkey_83_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_91_ ) ;
 assign wire8173 = ( wire8172 ) | ( (~ n_n2997)  &  (~ wire788)  &  wire7764 ) ;
 assign wire8176 = ( n_n2950  &  pksi_35_ ) ;
 assign wire8177 = ( pstart_0_  &  pkey_109_  &  pencrypt_0_ ) | ( pkey_117_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8178 = ( wire8177 ) | ( (~ n_n2997)  &  (~ wire869)  &  wire7764 ) ;
 assign wire8181 = ( pksi_20_  &  pksi_101_ ) ;
 assign wire8182 = ( pkey_3_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_11_ ) ;
 assign wire8183 = ( wire8182 ) | ( (~ n_n2997)  &  (~ wire870)  &  wire7764 ) ;
 assign wire8186 = ( pksi_179_  &  pksi_93_ ) ;
 assign wire8187 = ( pkey_218_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_226_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8188 = ( wire8187 ) | ( n_n2997  &  (~ wire814)  &  wire7763 ) ;
 assign wire8191 = ( n_n2770  &  pksi_161_ ) ;
 assign wire8192 = ( pkey_147_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_155_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8193 = ( wire8192 ) | ( (~ n_n2997)  &  (~ wire877)  &  wire7764 ) ;
 assign wire8196 = ( pksi_156_  &  pksi_66_ ) ;
 assign wire8197 = ( pkey_133_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_188_ ) ;
 assign wire8198 = ( wire8197 ) | ( (~ n_n2997)  &  (~ wire878)  &  wire7764 ) ;
 assign wire8201 = ( n_n2921  &  pksi_67_ ) ;
 assign wire8202 = ( pkey_134_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_142_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8203 = ( wire8202 ) | ( (~ n_n2997)  &  (~ wire879)  &  wire7764 ) ;
 assign wire8206 = ( n_n2931  &  pksi_40_ ) ;
 assign wire8207 = ( pstart_0_  &  pencrypt_0_  &  pkey_75_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_83_ ) ;
 assign wire8208 = ( wire8207 ) | ( (~ n_n2997)  &  (~ wire844)  &  wire7764 ) ;
 assign wire8211 = ( n_n2821  &  pksi_123_ ) ;
 assign wire8212 = ( pkey_117_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_125_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8213 = ( wire8212 ) | ( (~ n_n2997)  &  (~ wire875)  &  wire7764 ) ;
 assign wire8216 = ( pksi_7_  &  pksi_111_ ) ;
 assign wire8217 = ( pkey_126_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_3_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8218 = ( wire8217 ) | ( (~ n_n2997)  &  (~ wire876)  &  wire7764 ) ;
 assign wire8221 = ( pksi_173_  &  pksi_92_ ) ;
 assign wire8222 = ( pkey_227_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_235_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8223 = ( wire8222 ) | ( n_n2997  &  (~ wire851)  &  wire7763 ) ;
 assign wire8226 = ( pksi_15_  &  pksi_119_ ) ;
 assign wire8227 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_32_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_24_ ) ;
 assign wire8228 = ( wire8227 ) | ( n_n2997  &  (~ wire858)  &  wire7763 ) ;
 assign wire8231 = ( n_n2379  &  pksi_82_ ) ;
 assign wire8232 = ( pkey_212_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_220_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8233 = ( wire8232 ) | ( (~ n_n2997)  &  (~ wire828)  &  wire7764 ) ;
 assign wire8236 = ( pksi_145_  &  pksi_51_ ) ;
 assign wire8237 = ( pkey_155_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_132_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8238 = ( wire8237 ) | ( (~ n_n2997)  &  (~ wire883)  &  wire7764 ) ;
 assign wire8241 = ( pksi_144_  &  pksi_70_ ) ;
 assign wire8242 = ( pkey_149_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_157_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8243 = ( wire8242 ) | ( (~ n_n2997)  &  (~ wire873)  &  wire7764 ) ;
 assign wire8246 = ( pksi_150_  &  pksi_71_ ) ;
 assign wire8247 = ( pkey_182_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_174_ ) ;
 assign wire8248 = ( wire8247 ) | ( (~ n_n2997)  &  (~ wire791)  &  wire7764 ) ;
 assign wire8251 = ( pksi_37_  &  pksi_124_ ) ;
 assign wire8252 = ( pstart_0_  &  pencrypt_0_  &  pkey_100_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_44_ ) ;
 assign wire8253 = ( wire8252 ) | ( (~ n_n2997)  &  (~ wire860)  &  wire7764 ) ;
 assign wire8256 = ( pksi_132_  &  pksi_42_ ) ;
 assign wire8257 = ( pkey_124_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_69_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8258 = ( wire8257 ) | ( (~ n_n2997)  &  (~ wire792)  &  wire7764 ) ;
 assign wire8261 = ( pksi_130_  &  pksi_29_ ) ;
 assign wire8262 = ( pkey_86_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_94_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8263 = ( wire8262 ) | ( (~ n_n2997)  &  (~ wire854)  &  wire7764 ) ;
 assign wire8266 = ( pksi_1_  &  pksi_105_ ) ;
 assign wire8267 = ( pstart_0_  &  pkey_52_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_60_  &  (~ pencrypt_0_) ) ;
 assign wire8268 = ( wire8267 ) | ( (~ n_n2997)  &  (~ wire804)  &  wire7764 ) ;
 assign wire8271 = ( pksi_9_  &  pksi_112_ ) ;
 assign wire8272 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_22_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_14_ ) ;
 assign wire8273 = ( wire8272 ) | ( (~ n_n2997)  &  (~ wire809)  &  wire7764 ) ;
 assign wire8276 = ( n_n2280  &  n_n2865 ) ;
 assign wire8277 = ( pkey_235_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_243_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8278 = ( wire8277 ) | ( n_n2997  &  (~ wire794)  &  wire7763 ) ;
 assign wire8281 = ( pksi_6_  &  pksi_98_ ) ;
 assign wire8282 = ( pstart_0_  &  pencrypt_0_  &  pkey_32_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_40_ ) ;
 assign wire8283 = ( wire8282 ) | ( n_n2997  &  (~ wire841)  &  wire7763 ) ;
 assign wire8286 = ( n_n2741  &  pksi_188_ ) ;
 assign wire8287 = ( pkey_212_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_204_ ) ;
 assign wire8288 = ( wire8287 ) | ( (~ wire783)  &  (~ n_n2997)  &  wire7764 ) ;
 assign wire8291 = ( pksi_152_  &  pksi_60_ ) ;
 assign wire8292 = ( pkey_132_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_140_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8293 = ( wire8292 ) | ( (~ n_n2997)  &  (~ wire868)  &  wire7764 ) ;
 assign wire8296 = ( pksi_48_  &  pksi_163_ ) ;
 assign wire8297 = ( pkey_141_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_149_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8298 = ( wire8297 ) | ( (~ n_n2997)  &  (~ wire885)  &  wire7764 ) ;
 assign wire8301 = ( pksi_166_  &  pksi_52_ ) ;
 assign wire8302 = ( pkey_182_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_190_ ) ;
 assign wire8303 = ( wire8302 ) | ( (~ n_n2997)  &  (~ wire805)  &  wire7764 ) ;
 assign wire8306 = ( pksi_131_  &  pksi_45_ ) ;
 assign wire8307 = ( pkey_92_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_100_ ) ;
 assign wire8308 = ( wire8307 ) | ( (~ n_n2997)  &  (~ wire845)  &  wire7764 ) ;
 assign wire8311 = ( n_n2943  &  pksi_32_ ) ;
 assign wire8312 = ( pkey_69_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_77_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8313 = ( wire8312 ) | ( (~ n_n2997)  &  (~ wire833)  &  wire7764 ) ;
 assign wire8316 = ( pksi_136_  &  pksi_33_ ) ;
 assign wire8317 = ( pkey_78_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_86_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8318 = ( wire8317 ) | ( (~ n_n2997)  &  (~ wire859)  &  wire7764 ) ;
 assign wire8321 = ( pksi_18_  &  pksi_108_ ) ;
 assign wire8322 = ( pstart_0_  &  pkey_60_  &  pencrypt_0_ ) | ( pkey_5_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8323 = ( wire8322 ) | ( (~ n_n2997)  &  (~ wire882)  &  wire7764 ) ;
 assign wire8326 = ( n_n2986  &  pksi_19_ ) ;
 assign wire8327 = ( pkey_6_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_14_ ) ;
 assign wire8328 = ( wire8327 ) | ( (~ n_n2997)  &  (~ wire793)  &  wire7764 ) ;
 assign wire8331 = ( n_n2737  &  pksi_185_ ) ;
 assign wire8332 = ( pkey_243_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_251_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8333 = ( wire8332 ) | ( (~ wire776)  &  n_n2997  &  wire7763 ) ;
 assign wire8336 = ( pksi_175_  &  pksi_86_ ) ;
 assign wire8337 = ( pkey_221_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_229_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8338 = ( wire8337 ) | ( (~ n_n2997)  &  (~ wire800)  &  wire7764 ) ;
 assign wire8341 = ( pksi_190_  &  pksi_76_ ) ;
 assign wire8342 = ( pkey_246_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_254_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8343 = ( wire8342 ) | ( (~ n_n2997)  &  (~ wire830)  &  wire7764 ) ;
 assign wire8346 = ( n_n2774  &  pksi_164_ ) ;
 assign wire8347 = ( pkey_140_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_148_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8348 = ( wire8347 ) | ( (~ n_n2997)  &  (~ wire864)  &  wire7764 ) ;
 assign wire8351 = ( pksi_158_  &  pksi_50_ ) ;
 assign wire8352 = ( pkey_165_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_173_ ) ;
 assign wire8353 = ( wire8352 ) | ( (~ n_n2997)  &  (~ wire831)  &  wire7764 ) ;
 assign wire8356 = ( pksi_167_  &  pksi_63_ ) ;
 assign wire8357 = ( pkey_158_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_166_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8358 = ( wire8357 ) | ( (~ n_n2997)  &  (~ wire884)  &  wire7764 ) ;
 assign wire8361 = ( pksi_133_  &  pksi_34_ ) ;
 assign wire8362 = ( pkey_92_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_84_ ) ;
 assign wire8363 = ( wire8362 ) | ( (~ n_n2997)  &  (~ wire842)  &  wire7764 ) ;
 assign wire8366 = ( n_n2945  &  pksi_24_ ) ;
 assign wire8367 = ( pkey_77_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_85_  &  (~ pencrypt_0_) ) ;
 assign wire8368 = ( wire8367 ) | ( (~ n_n2997)  &  (~ wire820)  &  wire7764 ) ;
 assign wire8371 = ( pksi_30_  &  pksi_122_ ) ;
 assign wire8372 = ( pkey_110_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_102_ ) ;
 assign wire8373 = ( wire8372 ) | ( (~ n_n2997)  &  (~ wire789)  &  wire7764 ) ;
 assign wire8376 = ( n_n2976  &  pksi_8_ ) ;
 assign wire8377 = ( pkey_5_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_13_ ) ;
 assign wire8378 = ( wire8377 ) | ( (~ n_n2997)  &  (~ wire874)  &  wire7764 ) ;
 assign wire8381 = ( pksi_169_  &  pksi_75_ ) ;
 assign wire8382 = ( pkey_251_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_194_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8383 = ( wire8382 ) | ( n_n2997  &  (~ wire822)  &  wire7763 ) ;
 assign wire8386 = ( pksi_182_  &  pksi_74_ ) ;
 assign wire8387 = ( pkey_229_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_237_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8388 = ( wire8387 ) | ( (~ n_n2997)  &  (~ wire815)  &  wire7764 ) ;
 assign wire8391 = ( pksi_174_  &  pksi_95_ ) ;
 assign wire8392 = ( pkey_238_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_246_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8393 = ( wire8392 ) | ( (~ n_n2997)  &  (~ wire785)  &  wire7764 ) ;
 assign wire8396 = ( pksi_157_  &  pksi_58_ ) ;
 assign wire8397 = ( pkey_148_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_156_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8398 = ( wire8397 ) | ( (~ n_n2997)  &  (~ wire817)  &  wire7764 ) ;
 assign wire8401 = ( pksi_151_  &  pksi_62_ ) ;
 assign wire8402 = ( pkey_157_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_165_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8403 = ( wire8402 ) | ( (~ n_n2997)  &  (~ wire880)  &  wire7764 ) ;
 assign wire8406 = ( pksi_146_  &  pksi_54_ ) ;
 assign wire8407 = ( pkey_166_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_174_ ) ;
 assign wire8408 = ( wire8407 ) | ( (~ n_n2997)  &  (~ wire881)  &  wire7764 ) ;
 assign wire8411 = ( n_n2806  &  pksi_140_ ) ;
 assign wire8412 = ( pkey_76_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_84_ ) ;
 assign wire8413 = ( wire8412 ) | ( (~ n_n2997)  &  (~ wire832)  &  wire7764 ) ;
 assign wire8416 = ( pksi_46_  &  pksi_120_ ) ;
 assign wire8417 = ( pstart_0_  &  pkey_85_  &  pencrypt_0_ ) | ( pkey_93_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8418 = ( wire8417 ) | ( (~ n_n2997)  &  (~ wire886)  &  wire7764 ) ;
 assign wire8421 = ( n_n2438  &  pksi_39_ ) ;
 assign wire8422 = ( pkey_94_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_102_ ) ;
 assign wire8423 = ( wire8422 ) | ( (~ n_n2997)  &  (~ wire803)  &  wire7764 ) ;
 assign wire8426 = ( pksi_5_  &  pksi_106_ ) ;
 assign wire8427 = ( pstart_0_  &  pencrypt_0_  &  pkey_22_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_30_ ) ;
 assign wire8428 = ( wire8427 ) | ( (~ n_n2997)  &  (~ wire821)  &  wire7764 ) ;
 assign wire8431 = ( pksi_160_  &  pksi_57_ ) ;
 assign wire8432 = ( pkey_136_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_144_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8433 = ( wire8432 ) | ( n_n2997  &  (~ wire862)  &  wire7763 ) ;
 assign wire8436 = ( pksi_36_  &  pksi_128_ ) ;
 assign wire8437 = ( pkey_66_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_74_  &  (~ pencrypt_0_) ) ;
 assign wire8438 = ( wire8437 ) | ( n_n2997  &  (~ wire818)  &  wire7763 ) ;
 assign wire8441 = ( pksi_38_  &  pksi_127_ ) ;
 assign wire8442 = ( pkey_89_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_97_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8443 = ( wire8442 ) | ( n_n2997  &  (~ wire863)  &  wire7763 ) ;
 assign wire8446 = ( pksi_28_  &  pksi_142_ ) ;
 assign wire8447 = ( pkey_112_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_120_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8448 = ( wire8447 ) | ( n_n2997  &  (~ wire819)  &  wire7763 ) ;
 assign wire8451 = ( n_n2843  &  pksi_114_ ) ;
 assign wire8452 = ( pkey_50_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_42_ ) ;
 assign wire8453 = ( wire8452 ) | ( n_n2997  &  (~ wire790)  &  wire7763 ) ;
 assign wire8456 = ( pksi_154_  &  pksi_53_ ) ;
 assign wire8457 = ( pkey_144_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_152_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8458 = ( wire8457 ) | ( n_n2997  &  (~ wire866)  &  wire7763 ) ;
 assign wire8461 = ( pksi_121_  &  pksi_27_ ) ;
 assign wire8462 = ( pkey_123_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_66_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8463 = ( wire8462 ) | ( n_n2997  &  (~ wire802)  &  wire7763 ) ;
 assign wire8466 = ( pksi_134_  &  pksi_26_ ) ;
 assign wire8467 = ( pkey_97_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_105_ ) ;
 assign wire8468 = ( wire8467 ) | ( n_n2997  &  (~ wire867)  &  wire7763 ) ;
 assign wire8471 = ( pksi_47_  &  pksi_126_ ) ;
 assign wire8472 = ( pstart_0_  &  pkey_104_  &  pencrypt_0_ ) | ( pkey_112_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8473 = ( wire8472 ) | ( n_n2997  &  (~ wire807)  &  wire7763 ) ;
 assign wire8476 = ( pksi_1_  &  pksi_105_ ) ;
 assign wire8477 = ( pkey_50_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_58_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8478 = ( wire8477 ) | ( n_n2997  &  (~ wire804)  &  wire7763 ) ;
 assign wire8481 = ( pksi_167_  &  pksi_63_ ) ;
 assign wire8482 = ( pkey_152_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_160_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8483 = ( wire8482 ) | ( n_n2997  &  (~ wire884)  &  wire7763 ) ;
 assign wire8486 = ( pksi_133_  &  pksi_34_ ) ;
 assign wire8487 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_90_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_82_ ) ;
 assign wire8488 = ( wire8487 ) | ( n_n2997  &  (~ wire842)  &  wire7763 ) ;
 assign wire8491 = ( n_n2945  &  pksi_24_ ) ;
 assign wire8492 = ( pkey_81_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_73_ ) ;
 assign wire8493 = ( wire8492 ) | ( n_n2997  &  (~ wire820)  &  wire7763 ) ;
 assign wire8496 = ( pksi_30_  &  pksi_122_ ) ;
 assign wire8497 = ( pkey_96_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_104_  &  (~ pencrypt_0_) ) ;
 assign wire8498 = ( wire8497 ) | ( n_n2997  &  (~ wire789)  &  wire7763 ) ;
 assign wire8501 = ( pksi_18_  &  pksi_108_ ) ;
 assign wire8502 = ( pkey_58_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_1_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8503 = ( wire8502 ) | ( n_n2997  &  (~ wire882)  &  wire7763 ) ;
 assign wire8506 = ( pksi_79_  &  pksi_183_ ) ;
 assign wire8507 = ( pkey_56_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_227_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8508 = ( wire8507 ) | ( n_n2997  &  (~ wire855)  &  wire7763 ) ;
 assign wire8511 = ( pksi_146_  &  pksi_54_ ) ;
 assign wire8512 = ( pkey_160_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_168_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8513 = ( wire8512 ) | ( n_n2997  &  (~ wire881)  &  wire7763 ) ;
 assign wire8516 = ( n_n2806  &  pksi_140_ ) ;
 assign wire8517 = ( pstart_0_  &  pkey_74_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_82_ ) ;
 assign wire8518 = ( wire8517 ) | ( n_n2997  &  (~ wire832)  &  wire7763 ) ;
 assign wire8521 = ( pksi_46_  &  pksi_120_ ) ;
 assign wire8522 = ( pkey_81_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_89_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8523 = ( wire8522 ) | ( n_n2997  &  (~ wire886)  &  wire7763 ) ;
 assign wire8526 = ( n_n2438  &  pksi_39_ ) ;
 assign wire8527 = ( pkey_88_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_96_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8528 = ( wire8527 ) | ( n_n2997  &  (~ wire803)  &  wire7763 ) ;
 assign wire8531 = ( n_n2976  &  pksi_8_ ) ;
 assign wire8532 = ( pkey_1_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_9_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8533 = ( wire8532 ) | ( n_n2997  &  (~ wire874)  &  wire7763 ) ;
 assign wire8536 = ( n_n2746  &  pksi_186_ ) ;
 assign wire8537 = ( pkey_234_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_242_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8538 = ( wire8537 ) | ( n_n2997  &  (~ wire836)  &  wire7763 ) ;
 assign wire8541 = ( n_n2889  &  pksi_91_ ) ;
 assign wire8542 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_200_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_192_ ) ;
 assign wire8543 = ( wire8542 ) | ( n_n2997  &  (~ wire837)  &  wire7763 ) ;
 assign wire8546 = ( pksi_145_  &  pksi_51_ ) ;
 assign wire8547 = ( pkey_130_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_187_ ) ;
 assign wire8548 = ( wire8547 ) | ( n_n2997  &  (~ wire883)  &  wire7763 ) ;
 assign wire8551 = ( pksi_144_  &  pksi_70_ ) ;
 assign wire8552 = ( pkey_145_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_153_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8553 = ( wire8552 ) | ( n_n2997  &  (~ wire873)  &  wire7763 ) ;
 assign wire8556 = ( pksi_0_  &  pksi_115_ ) ;
 assign wire8557 = ( pkey_9_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_17_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8558 = ( wire8557 ) | ( n_n2997  &  (~ wire840)  &  wire7763 ) ;
 assign wire8561 = ( pksi_177_  &  pksi_73_ ) ;
 assign wire8562 = ( pkey_242_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_250_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8563 = ( wire8562 ) | ( n_n2997  &  (~ wire847)  &  wire7763 ) ;
 assign wire8566 = ( pksi_89_  &  pksi_189_ ) ;
 assign wire8567 = ( pkey_249_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_192_ ) ;
 assign wire8568 = ( wire8567 ) | ( n_n2997  &  (~ wire848)  &  wire7763 ) ;
 assign wire8571 = ( pksi_152_  &  pksi_60_ ) ;
 assign wire8572 = ( pkey_130_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_138_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8573 = ( wire8572 ) | ( n_n2997  &  (~ wire868)  &  wire7763 ) ;
 assign wire8576 = ( pksi_48_  &  pksi_163_ ) ;
 assign wire8577 = ( pkey_137_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_145_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8578 = ( wire8577 ) | ( n_n2997  &  (~ wire885)  &  wire7763 ) ;
 assign wire8581 = ( pksi_22_  &  pksi_96_ ) ;
 assign wire8582 = ( pkey_17_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_25_ ) ;
 assign wire8583 = ( wire8582 ) | ( n_n2997  &  (~ wire857)  &  wire7763 ) ;
 assign wire8586 = ( n_n2749  &  pksi_180_ ) ;
 assign wire8587 = ( pkey_250_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_193_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8588 = ( wire8587 ) | ( n_n2997  &  (~ wire810)  &  wire7763 ) ;
 assign wire8591 = ( pksi_178_  &  pksi_77_ ) ;
 assign wire8592 = ( pstart_0_  &  pkey_208_  &  pencrypt_0_ ) | ( pkey_216_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8593 = ( wire8592 ) | ( n_n2997  &  (~ wire811)  &  wire7763 ) ;
 assign wire8596 = ( n_n2899  &  pksi_64_ ) ;
 assign wire8597 = ( pstart_0_  &  pkey_171_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_179_ ) ;
 assign wire8598 = ( wire8597 ) | ( n_n2997  &  (~ wire871)  &  wire7763 ) ;
 assign wire8601 = ( pksi_153_  &  pksi_56_ ) ;
 assign wire8602 = ( pkey_129_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_137_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8603 = ( wire8602 ) | ( n_n2997  &  (~ wire872)  &  wire7763 ) ;
 assign wire8606 = ( n_n2877  &  pksi_80_ ) ;
 assign wire8607 = ( pkey_193_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_201_ ) ;
 assign wire8608 = ( wire8607 ) | ( n_n2997  &  (~ wire823)  &  wire7763 ) ;
 assign wire8611 = ( pksi_184_  &  pksi_81_ ) ;
 assign wire8612 = ( pstart_0_  &  pkey_208_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_200_ ) ;
 assign wire8613 = ( wire8612 ) | ( n_n2997  &  (~ wire824)  &  wire7763 ) ;
 assign wire8616 = ( n_n2770  &  pksi_161_ ) ;
 assign wire8617 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_187_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_179_ ) ;
 assign wire8618 = ( wire8617 ) | ( n_n2997  &  (~ wire877)  &  wire7763 ) ;
 assign wire8621 = ( pksi_156_  &  pksi_66_ ) ;
 assign wire8622 = ( pkey_129_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_186_ ) ;
 assign wire8623 = ( wire8622 ) | ( n_n2997  &  (~ wire878)  &  wire7763 ) ;
 assign wire8626 = ( n_n2879  &  pksi_72_ ) ;
 assign wire8627 = ( pkey_209_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_201_ ) ;
 assign wire8628 = ( wire8627 ) | ( (~ wire777)  &  n_n2997  &  wire7763 ) ;
 assign wire8631 = ( pksi_78_  &  pksi_170_ ) ;
 assign wire8632 = ( pkey_224_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_232_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8633 = ( wire8632 ) | ( (~ wire778)  &  n_n2997  &  wire7763 ) ;
 assign wire8636 = ( pksi_155_  &  pksi_69_ ) ;
 assign wire8637 = ( pkey_154_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_162_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8638 = ( wire8637 ) | ( (~ wire779)  &  n_n2997  &  wire7763 ) ;
 assign wire8641 = ( n_n2789  &  pksi_147_ ) ;
 assign wire8642 = ( pstart_0_  &  pencrypt_0_  &  pkey_177_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_185_ ) ;
 assign wire8643 = ( wire8642 ) | ( (~ wire780)  &  n_n2997  &  wire7763 ) ;
 assign wire8646 = ( n_n2931  &  pksi_40_ ) ;
 assign wire8647 = ( pkey_107_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_115_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8648 = ( wire8647 ) | ( n_n2997  &  (~ wire844)  &  wire7763 ) ;
 assign wire8651 = ( n_n2943  &  pksi_32_ ) ;
 assign wire8652 = ( pstart_0_  &  pencrypt_0_  &  pkey_65_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_73_ ) ;
 assign wire8653 = ( wire8652 ) | ( n_n2997  &  (~ wire833)  &  wire7763 ) ;
 assign wire8656 = ( n_n2881  &  pksi_94_ ) ;
 assign wire8657 = ( pkey_209_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_217_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8658 = ( wire8657 ) | ( n_n2997  &  (~ wire784)  &  wire7763 ) ;
 assign wire8661 = ( n_n2391  &  pksi_87_ ) ;
 assign wire8662 = ( pkey_216_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_224_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8663 = ( wire8662 ) | ( n_n2997  &  (~ wire795)  &  wire7763 ) ;
 assign wire8666 = ( pksi_148_  &  pksi_61_ ) ;
 assign wire8667 = ( pkey_162_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_170_ ) ;
 assign wire8668 = ( wire8667 ) | ( n_n2997  &  (~ wire786)  &  wire7763 ) ;
 assign wire8671 = ( n_n2917  &  pksi_59_ ) ;
 assign wire8672 = ( pkey_169_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_177_ ) ;
 assign wire8673 = ( wire8672 ) | ( n_n2997  &  (~ wire796)  &  wire7763 ) ;
 assign wire8676 = ( n_n2802  &  pksi_137_ ) ;
 assign wire8677 = ( pkey_115_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_123_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8678 = ( wire8677 ) | ( n_n2997  &  (~ wire788)  &  wire7763 ) ;
 assign wire8681 = ( pksi_132_  &  pksi_42_ ) ;
 assign wire8682 = ( pkey_122_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_65_ ) ;
 assign wire8683 = ( wire8682 ) | ( n_n2997  &  (~ wire792)  &  wire7763 ) ;
 assign wire8686 = ( pksi_175_  &  pksi_86_ ) ;
 assign wire8687 = ( pkey_217_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_225_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8688 = ( wire8687 ) | ( n_n2997  &  (~ wire800)  &  wire7763 ) ;
 assign wire8691 = ( pksi_190_  &  pksi_76_ ) ;
 assign wire8692 = ( pkey_240_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_248_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8693 = ( wire8692 ) | ( n_n2997  &  (~ wire830)  &  wire7763 ) ;
 assign wire8696 = ( n_n2774  &  pksi_164_ ) ;
 assign wire8697 = ( pkey_138_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_146_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8698 = ( wire8697 ) | ( n_n2997  &  (~ wire864)  &  wire7763 ) ;
 assign wire8701 = ( pksi_158_  &  pksi_50_ ) ;
 assign wire8702 = ( pkey_161_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_169_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8703 = ( wire8702 ) | ( n_n2997  &  (~ wire831)  &  wire7763 ) ;
 assign wire8706 = ( pksi_136_  &  pksi_33_ ) ;
 assign wire8707 = ( pkey_80_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_72_ ) ;
 assign wire8708 = ( wire8707 ) | ( n_n2997  &  (~ wire859)  &  wire7763 ) ;
 assign wire8711 = ( pksi_104_  &  pksi_12_ ) ;
 assign wire8712 = ( pkey_2_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_10_ ) ;
 assign wire8713 = ( wire8712 ) | ( n_n2997  &  (~ wire853)  &  wire7763 ) ;
 assign wire8716 = ( pksi_182_  &  pksi_74_ ) ;
 assign wire8717 = ( pkey_225_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_233_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8718 = ( wire8717 ) | ( n_n2997  &  (~ wire815)  &  wire7763 ) ;
 assign wire8721 = ( pksi_174_  &  pksi_95_ ) ;
 assign wire8722 = ( pkey_232_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_240_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8723 = ( wire8722 ) | ( n_n2997  &  (~ wire785)  &  wire7763 ) ;
 assign wire8726 = ( pksi_157_  &  pksi_58_ ) ;
 assign wire8727 = ( pkey_146_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_154_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8728 = ( wire8727 ) | ( n_n2997  &  (~ wire817)  &  wire7763 ) ;
 assign wire8731 = ( pksi_151_  &  pksi_62_ ) ;
 assign wire8732 = ( pkey_153_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_161_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8733 = ( wire8732 ) | ( n_n2997  &  (~ wire880)  &  wire7763 ) ;
 assign wire8736 = ( pksi_130_  &  pksi_29_ ) ;
 assign wire8737 = ( pkey_80_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_88_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8738 = ( wire8737 ) | ( n_n2997  &  (~ wire854)  &  wire7763 ) ;
 assign wire8741 = ( pksi_3_  &  pksi_97_ ) ;
 assign wire8742 = ( pkey_59_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_2_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8743 = ( wire8742 ) | ( n_n2997  &  (~ wire850)  &  wire7763 ) ;
 assign wire8746 = ( n_n2885  &  pksi_83_ ) ;
 assign wire8747 = ( pkey_233_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_241_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8748 = ( wire8747 ) | ( n_n2997  &  (~ wire829)  &  wire7763 ) ;
 assign wire8751 = ( pksi_149_  &  pksi_68_ ) ;
 assign wire8752 = ( pkey_163_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_171_  &  (~ pencrypt_0_) ) ;
 assign wire8753 = ( wire8752 ) | ( n_n2997  &  (~ wire865)  &  wire7763 ) ;
 assign wire8756 = ( pksi_150_  &  pksi_71_ ) ;
 assign wire8757 = ( pkey_168_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_176_ ) ;
 assign wire8758 = ( wire8757 ) | ( n_n2997  &  (~ wire791)  &  wire7763 ) ;
 assign wire8761 = ( pksi_37_  &  pksi_124_ ) ;
 assign wire8762 = ( pkey_98_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_106_ ) ;
 assign wire8763 = ( wire8762 ) | ( n_n2997  &  (~ wire860)  &  wire7763 ) ;
 assign wire8766 = ( pksi_141_  &  pksi_41_ ) ;
 assign wire8767 = ( pkey_121_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_64_ ) ;
 assign wire8768 = ( wire8767 ) | ( n_n2997  &  (~ wire838)  &  wire7763 ) ;
 assign wire8771 = ( n_n2834  &  pksi_113_ ) ;
 assign wire8772 = ( pstart_0_  &  pkey_51_  &  pencrypt_0_ ) | ( pkey_59_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8773 = ( wire8772 ) | ( n_n2997  &  (~ wire839)  &  wire7763 ) ;
 assign wire8776 = ( n_n2838  &  pksi_116_ ) ;
 assign wire8777 = ( pkey_18_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_10_ ) ;
 assign wire8778 = ( wire8777 ) | ( n_n2997  &  (~ wire856)  &  wire7763 ) ;
 assign wire8781 = ( n_n2757  &  pksi_171_ ) ;
 assign wire8782 = ( pkey_241_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_249_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8783 = ( wire8782 ) | ( n_n2997  &  (~ wire852)  &  wire7763 ) ;
 assign wire8786 = ( pksi_159_  &  pksi_55_ ) ;
 assign wire8787 = ( pkey_248_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_163_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8788 = ( wire8787 ) | ( n_n2997  &  (~ wire816)  &  wire7763 ) ;
 assign wire8791 = ( pksi_166_  &  pksi_52_ ) ;
 assign wire8792 = ( pstart_0_  &  pencrypt_0_  &  pkey_176_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_184_ ) ;
 assign wire8793 = ( wire8792 ) | ( n_n2997  &  (~ wire805)  &  wire7763 ) ;
 assign wire8796 = ( pksi_131_  &  pksi_45_ ) ;
 assign wire8797 = ( pkey_98_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_90_ ) ;
 assign wire8798 = ( wire8797 ) | ( n_n2997  &  (~ wire845)  &  wire7763 ) ;
 assign wire8801 = ( n_n2954  &  pksi_43_ ) ;
 assign wire8802 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_72_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_64_ ) ;
 assign wire8803 = ( wire8802 ) | ( n_n2997  &  (~ wire843)  &  wire7763 ) ;
 assign wire8806 = ( n_n2964  &  pksi_16_ ) ;
 assign wire8807 = ( pstart_0_  &  pkey_51_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_43_ ) ;
 assign wire8808 = ( wire8807 ) | ( n_n2997  &  (~ wire849)  &  wire7763 ) ;
 assign wire8811 = ( pksi_10_  &  pksi_109_ ) ;
 assign wire8812 = ( pkey_18_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_26_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8813 = ( wire8812 ) | ( (~ wire781)  &  n_n2997  &  wire7763 ) ;
 assign wire8816 = ( n_n2779  &  pksi_162_ ) ;
 assign wire8817 = ( pstart_0_  &  pencrypt_0_  &  pkey_170_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_178_ ) ;
 assign wire8818 = ( wire8817 ) | ( n_n2997  &  (~ wire801)  &  wire7763 ) ;
 assign wire8821 = ( n_n2921  &  pksi_67_ ) ;
 assign wire8822 = ( pkey_128_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_136_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8823 = ( wire8822 ) | ( n_n2997  &  (~ wire879)  &  wire7763 ) ;
 assign wire8826 = ( pksi_135_  &  pksi_31_ ) ;
 assign wire8827 = ( pkey_99_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_184_ ) ;
 assign wire8828 = ( wire8827 ) | ( n_n2997  &  (~ wire812)  &  wire7763 ) ;
 assign wire8831 = ( pksi_25_  &  pksi_129_ ) ;
 assign wire8832 = ( pkey_114_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_122_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8833 = ( wire8832 ) | ( n_n2997  &  (~ wire806)  &  wire7763 ) ;
 assign wire8836 = ( n_n2950  &  pksi_35_ ) ;
 assign wire8837 = ( pkey_113_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_105_ ) ;
 assign wire8838 = ( wire8837 ) | ( n_n2997  &  (~ wire869)  &  wire7763 ) ;
 assign wire8841 = ( pksi_20_  &  pksi_101_ ) ;
 assign wire8842 = ( pstart_0_  &  pencrypt_0_  &  pkey_35_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_43_ ) ;
 assign wire8843 = ( wire8842 ) | ( n_n2997  &  (~ wire870)  &  wire7763 ) ;
 assign wire8846 = ( pksi_21_  &  pksi_107_ ) ;
 assign wire8847 = ( pkey_26_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_34_ ) ;
 assign wire8848 = ( wire8847 ) | ( n_n2997  &  (~ wire797)  &  wire7763 ) ;
 assign wire8851 = ( n_n2909  &  pksi_49_ ) ;
 assign wire8852 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_186_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_178_ ) ;
 assign wire8853 = ( wire8852 ) | ( n_n2997  &  (~ wire861)  &  wire7763 ) ;
 assign wire8856 = ( pksi_165_  &  pksi_65_ ) ;
 assign wire8857 = ( pkey_128_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_185_ ) ;
 assign wire8858 = ( wire8857 ) | ( n_n2997  &  (~ wire787)  &  wire7763 ) ;
 assign wire8861 = ( pksi_44_  &  pksi_125_ ) ;
 assign wire8862 = ( pkey_99_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_107_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8863 = ( wire8862 ) | ( n_n2997  &  (~ wire825)  &  wire7763 ) ;
 assign wire8866 = ( n_n2811  &  pksi_138_ ) ;
 assign wire8867 = ( pkey_114_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_106_ ) ;
 assign wire8868 = ( wire8867 ) | ( n_n2997  &  (~ wire826)  &  wire7763 ) ;
 assign wire8871 = ( n_n2821  &  pksi_123_ ) ;
 assign wire8872 = ( pkey_113_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_121_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire8873 = ( wire8872 ) | ( n_n2997  &  (~ wire875)  &  wire7763 ) ;
 assign wire8876 = ( pksi_7_  &  pksi_111_ ) ;
 assign wire8877 = ( pkey_120_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_35_ ) ;
 assign wire8878 = ( wire8877 ) | ( n_n2997  &  (~ wire876)  &  wire7763 ) ;
 assign wire8881 = ( pksi_13_  &  pksi_100_ ) ;
 assign wire8882 = ( pstart_0_  &  pencrypt_0_  &  pkey_34_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_42_ ) ;
 assign wire8883 = ( wire8882 ) | ( n_n2997  &  (~ wire808)  &  wire7763 ) ;
 assign wire8889 = ( pencrypt_0_  &  wire774 ) | ( (~ pcount_0_)  &  (~ pencrypt_0_)  &  wire887 ) ;


endmodule

