module s298 (
	s298_in_0_, s298_in_2_, s298_in_1_, clock, s298_out_0_, s298_out_1_, s298_out_2_, s298_out_3_, 
	s298_out_4_, s298_out_5_);

input s298_in_0_;
input s298_in_2_;
input s298_in_1_;
input clock;
output s298_out_0_;
output s298_out_1_;
output s298_out_2_;
output s298_out_3_;
output s298_out_4_;
output s298_out_5_;
wire n_n45;
wire n_n46;
wire n_n47;
wire n_n48;
wire n_n49;
wire n_n50;
wire n_n51;
wire n_n52;
wire wire24;
wire wire25;
wire wire27;
wire wire29;
wire wire30;
wire wire39;
wire wire40;
wire wire41;
wire wire42;
wire wire44;
wire wire45;
wire wire57;
wire wire58;
wire wire59;
wire wire60;
wire wire61;
wire wire62;
wire wire63;
wire wire66;
wire wire68;
wire wire69;
wire wire76;
wire wire77;
wire wire78;
wire wire79;
wire wire80;
wire wire81;
wire wire86;
wire wire87;
wire wire88;
wire wire89;
wire wire90;
wire wire91;
wire wire94;
wire wire101;
wire wire102;
wire wire103;
wire wire104;
wire wire107;
wire wire108;
wire wire109;
wire wire110;
wire wire111;
wire wire112;
wire wire113;
wire wire114;
wire wire115;
wire wire116;
wire wire117;
wire wire118;
wire wire133;
wire wire134;
wire wire135;
wire wire136;
wire wire137;
wire wire138;
wire wire139;
wire wire140;
wire wire148;
wire wire153;
wire wire154;
wire wire155;
wire wire156;
wire wire161;
wire wire179;
wire wire180;
wire wire181;
wire wire182;
wire wire202;
wire wire204;
wire wire206;
wire wire210;
wire wire214;
wire wire215;
wire wire216;
wire wire217;
wire wire218;
wire wire224;
wire wire226;
wire wire227;
wire wire228;
wire wire229;
wire wire230;
wire wire231;
wire wire232;
wire wire233;
wire wire234;
wire wire249;
wire wire250;
wire wire251;
wire wire252;
wire wire253;
wire wire254;
wire wire265;
wire wire266;
wire wire267;
wire wire269;
wire wire278;
wire wire279;
wire wire303;
wire wire304;
wire wire305;
wire wire306;
wire wire307;
wire wire308;
wire wire309;
wire wire320;
wire wire321;
wire wire322;
wire wire323;
wire wire324;
wire wire325;
wire wire334;
wire wire335;
wire wire336;
wire wire337;
wire wire338;
wire wire339;
wire wire340;
wire wire341;
wire wire342;
wire wire344;
wire wire346;
wire wire347;
wire wire351;
wire wire353;
wire wire355;
wire wire359;
wire wire360;
wire wire361;
wire wire362;
wire wire363;
wire wire364;
wire wire365;
wire wire366;
wire wire367;
wire wire368;
wire wire369;
wire wire384;
wire wire385;
wire wire386;
wire wire387;
wire wire388;
wire wire391;
wire wire397;
wire wire398;
wire wire399;
wire wire400;
wire wire401;
wire wire402;
wire wire403;
wire wire424;
wire wire425;
wire wire426;
wire wire427;
wire wire428;
wire wire429;
wire wire430;
wire wire431;
wire wire432;
wire wire436;
wire wire441;
wire wire442;
wire wire443;
wire wire444;
wire wire445;
wire wire446;
wire wire447;
wire wire448;
wire wire449;
wire wire450;
wire wire451;
wire wire452;
wire wire453;
wire wire454;
wire wire455;
wire wire457;
wire wire458;
wire wire462;
wire wire463;
wire wire464;
wire wire470;
wire wire471;
wire wire472;
wire wire473;
wire wire474;
wire wire475;
wire wire476;
wire wire477;
wire wire478;
wire wire479;
wire wire483;
wire wire484;
wire wire485;
wire wire494;
wire wire495;
wire wire496;
wire wire497;
wire wire498;
wire wire499;
wire wire500;
wire wire501;
wire wire504;
wire wire505;
wire wire506;
wire wire507;
wire wire510;
wire wire511;
wire wire513;
wire wire518;
wire wire519;
wire wire526;
wire wire531;
wire wire532;
wire wire535;
wire wire536;
wire wire542;
wire wire544;
wire wire550;
wire wire553;
wire wire556;
wire wire558;
wire wire566;
wire wire567;
wire wire568;
wire wire570;
wire wire571;
wire wire576;
wire wire577;
wire wire578;
wire wire579;
wire wire580;
wire wire581;
wire wire582;
wire wire611;
wire wire612;
wire wire613;
wire wire614;
wire wire615;
wire wire616;
wire wire619;
wire wire621;
wire wire622;
wire wire623;
wire wire624;
wire wire625;
wire wire5509;
wire wire5513;
wire wire5518;
wire wire5519;
wire wire5524;
wire wire5525;
wire wire5526;
wire wire5530;
wire wire5531;
wire wire5533;
wire wire5534;
wire wire5537;
wire wire5538;
wire wire5541;
wire wire5542;
wire wire5548;
wire wire5549;
wire wire5554;
wire wire5555;
wire wire5560;
wire wire5561;
wire wire5566;
wire wire5567;
wire wire5572;
wire wire5573;
wire wire5578;
wire wire5579;
wire wire5582;
wire wire5583;
wire wire5586;
wire wire5587;
wire wire5590;
wire wire5591;
wire wire5594;
wire wire5595;
wire wire5599;
wire wire5603;
wire wire5606;
wire wire5607;
wire wire5610;
wire wire5611;
wire wire5615;
wire wire5619;
wire wire5623;
wire wire5627;
wire wire5630;
wire wire5631;
wire wire5633;
wire wire5634;
wire wire5636;
wire wire5637;
wire wire5639;
wire wire5640;
wire wire5642;
wire wire5643;
wire wire5645;
wire wire5646;
wire wire5648;
wire wire5649;
wire wire5651;
wire wire5652;
wire wire5655;
wire wire5658;
wire wire5675;
wire wire5676;
wire wire5677;
wire wire5678;
wire wire5679;
wire wire5680;
wire wire5681;
wire wire5682;
wire wire5683;
wire wire5684;
wire wire5685;
wire wire5686;
wire wire5687;
wire wire5688;
wire wire5689;
wire wire5690;
wire wire5691;
wire wire5700;
wire wire5701;
wire wire5702;
wire wire5703;
wire wire5707;
wire wire5708;
wire wire5712;
wire wire5717;
wire wire5719;
wire wire5720;
wire wire5723;
wire wire5725;
wire wire5726;
wire wire5729;
wire wire5732;
wire wire5734;
wire wire5736;
wire wire5738;
wire wire5740;
wire wire5741;
wire wire5744;
wire wire5746;
wire wire5748;
wire wire5750;
wire wire5752;
wire wire5754;
wire wire5759;
wire wire5763;
wire wire5766;
wire wire5767;
wire wire5768;
wire wire5772;
wire wire5774;
wire wire5775;
wire wire5776;
wire wire5777;
wire wire5780;
wire wire5781;
wire wire5782;
wire wire5783;
wire wire5784;
wire wire5785;
wire wire5787;
wire wire5789;
wire wire5790;
wire wire5791;
wire wire5796;
wire wire5797;
wire wire5798;
wire wire5803;
wire wire5804;
wire wire5810;
wire wire5811;
wire wire5817;
wire wire5818;
wire wire5821;
wire wire5822;
wire wire5824;
wire wire5827;
wire wire5828;
wire wire5830;
wire wire5834;
wire wire5835;
wire wire5841;
wire wire5842;
wire wire5847;
wire wire5848;
wire wire5850;
wire wire5851;
wire wire5853;
wire wire5856;
wire wire5858;
wire wire5861;
wire wire5862;
wire wire5865;
wire wire5866;
wire wire5868;
wire wire5870;
wire wire5871;
wire wire5873;
wire wire5877;
wire wire5878;
wire wire5882;
wire wire5883;
wire wire5886;
wire wire5887;
wire wire5892;
wire wire5893;
wire wire5897;
wire wire5898;
wire wire5902;
wire wire5903;
wire wire5905;
wire wire5906;
wire wire5907;
wire wire5910;
wire wire5911;
wire wire5914;
wire wire5915;
wire wire5918;
wire wire5919;
wire wire5922;
wire wire5923;
wire wire5925;
wire wire5927;
wire wire5929;
wire wire5930;
wire wire5934;
wire wire5938;
wire wire5939;
wire wire5942;
wire wire5943;
wire wire5946;
wire wire5947;
wire wire5950;
wire wire5951;
wire wire5954;
wire wire5955;
wire wire5957;
wire wire5961;
wire wire5963;
wire wire5966;
wire wire5967;
wire wire5970;
wire wire5972;
wire wire5973;
wire wire5976;
wire wire5978;
wire wire5980;
wire wire5981;
wire wire5982;
wire wire5984;
wire wire5986;
wire wire5987;
wire wire5988;
wire wire5989;
wire wire5990;
wire wire5992;
wire wire5993;
wire wire5994;
wire wire5995;
wire wire5996;
wire wire5997;
wire wire5998;
wire wire6001;
wire wire6005;
wire wire6006;
wire wire6007;
wire wire6009;
wire wire6016;
wire wire6017;
wire wire6018;
wire wire6022;
wire wire6023;
wire wire6025;
wire wire6028;
wire wire6029;
wire wire6031;
wire wire6033;
wire wire6034;
wire wire6036;
wire wire6037;
wire wire6040;
wire wire6041;
wire wire6043;
wire wire6046;
wire wire6047;
wire wire6049;
wire wire6053;
wire wire6054;
wire wire6055;
wire wire6058;
wire wire6059;
wire wire6061;
wire wire6065;
wire wire6066;
wire wire6067;
wire wire6072;
wire wire6073;
wire wire6076;
wire wire6077;
wire wire6079;
wire wire6083;
wire wire6084;
wire wire6090;
wire wire6091;
wire wire6095;
wire wire6096;
wire wire6101;
wire wire6102;
wire wire6108;
wire wire6109;
wire wire6114;
wire wire6115;
wire wire6120;
wire wire6121;
wire wire6126;
wire wire6127;
wire wire6132;
wire wire6133;
wire wire6138;
wire wire6139;
wire wire6144;
wire wire6145;
wire wire6148;
wire wire6149;
wire wire6150;
wire wire6154;
wire wire6155;
wire wire6159;
wire wire6160;
wire wire6162;
wire wire6164;
wire wire6165;
wire wire6167;
wire wire6168;
wire wire6170;
wire wire6172;
wire wire6173;
wire wire6175;
wire wire6178;
wire wire6180;
wire wire6183;
wire wire6184;
wire wire6185;
wire wire6189;
wire wire6190;
wire wire6194;
wire wire6195;
wire wire6197;
wire wire6198;
wire wire6200;
wire wire6203;
wire wire6204;
wire wire6209;
wire wire6210;
wire wire6214;
wire wire6215;
wire wire6217;
wire wire6218;
wire wire6220;
wire wire6222;
wire wire6223;
wire wire6225;
wire wire6227;
wire wire6228;
wire wire6230;
wire wire6234;
wire wire6235;
wire wire6238;
wire wire6239;
wire wire6244;
wire wire6245;
wire wire6248;
wire wire6249;
wire wire6254;
wire wire6255;
wire wire6258;
wire wire6259;
wire wire6264;
wire wire6265;
wire wire6269;
wire wire6270;
wire wire6273;
wire wire6274;
wire wire6277;
wire wire6278;
wire wire6280;
wire wire6282;
wire wire6285;
wire wire6286;
wire wire6289;
wire wire6290;
wire wire6293;
wire wire6294;
wire wire6297;
wire wire6298;
wire wire6301;
wire wire6302;
wire wire6305;
wire wire6306;
wire wire6309;
wire wire6310;
wire wire6312;
wire wire6313;
wire wire6315;
wire wire6318;
wire wire6319;
wire wire6320;
wire wire6323;
wire wire6324;
wire wire6325;
wire wire6328;
wire wire6329;
wire wire6330;
wire wire6331;
wire wire6332;
wire wire6333;
wire wire6334;
wire wire6335;
wire wire6338;
wire wire6339;
wire wire6342;
wire wire6344;
wire wire6345;
wire wire6351;
wire wire6352;
wire wire6354;
wire wire6367;
wire wire6368;
wire wire6369;
wire wire6370;
wire wire6371;
wire wire6372;
wire wire6375;
wire wire6376;
wire wire6381;
wire wire6382;
wire wire6384;
wire wire6389;
wire wire6390;
wire wire6392;
wire wire6397;
wire wire6398;
wire wire6399;
wire wire6404;
wire wire6406;
wire wire6407;
wire wire6410;
wire wire6412;
wire wire6413;
wire wire6414;
wire wire6418;
wire wire6419;
wire wire6421;
wire wire6425;
wire wire6426;
wire wire6428;
wire wire6431;
wire wire6432;
wire wire6434;
wire wire6435;
wire wire6440;
wire wire6441;
wire wire6442;
wire wire6447;
wire wire6448;
wire wire6449;
wire wire6454;
wire wire6455;
wire wire6456;
wire wire6461;
wire wire6462;
wire wire6463;
wire wire6467;
wire wire6468;
wire wire6470;
wire wire6473;
wire wire6474;
wire wire6476;
wire wire6477;
wire wire6481;
wire wire6482;
wire wire6484;
wire wire6488;
wire wire6489;
wire wire6491;
wire wire6496;
wire wire6497;
wire wire6498;
wire wire6503;
wire wire6504;
wire wire6505;
wire wire6510;
wire wire6511;
wire wire6512;
wire wire6517;
wire wire6518;
wire wire6523;
wire wire6524;
wire wire6526;
wire wire6531;
wire wire6532;
wire wire6533;
wire wire6537;
wire wire6538;
wire wire6540;
wire wire6545;
wire wire6546;
wire wire6552;
wire wire6553;
wire wire6554;
wire wire6559;
wire wire6560;
wire wire6561;
wire wire6566;
wire wire6567;
wire wire6568;
wire wire6572;
wire wire6573;
wire wire6575;
wire wire6580;
wire wire6581;
wire wire6582;
wire wire6586;
wire wire6587;
wire wire6589;
wire wire6594;
wire wire6595;
wire wire6600;
wire wire6601;
wire wire6603;
wire wire6608;
wire wire6609;
wire wire6610;
wire wire6615;
wire wire6616;
wire wire6622;
wire wire6623;
wire wire6629;
wire wire6630;
wire wire6631;
wire wire6636;
wire wire6637;
wire wire6638;
wire wire6643;
wire wire6644;
wire wire6650;
wire wire6651;
wire wire6657;
wire wire6658;
wire wire6664;
wire wire6665;
wire wire6671;
wire wire6672;
wire wire6678;
wire wire6679;
wire wire6685;
wire wire6686;
wire wire6692;
wire wire6693;
wire wire6699;
wire wire6700;
wire wire6705;
wire wire6706;
wire wire6707;
wire wire6711;
wire wire6712;
wire wire6713;
wire wire6715;
wire wire6716;
wire wire6718;
wire wire6719;
wire wire6721;
wire wire6722;
wire wire6724;
wire wire6725;
wire wire6728;
wire wire6729;
wire wire6731;
wire wire6733;
wire wire6734;
wire wire6736;
wire wire6737;
wire wire6740;
wire wire6741;
wire wire6743;
wire wire6747;
wire wire6748;
wire wire6749;
wire wire6754;
wire wire6755;
wire wire6760;
wire wire6761;
wire wire6763;
wire wire6764;
wire wire6767;
wire wire6770;
wire wire6772;
wire wire6773;
wire wire6778;
wire wire6779;
wire wire6783;
wire wire6784;
wire wire6785;
wire wire6787;
wire wire6788;
wire wire6790;
wire wire6791;
wire wire6794;
wire wire6795;
wire wire6797;
wire wire6800;
wire wire6801;
wire wire6803;
wire wire6807;
wire wire6808;
wire wire6809;
wire wire6814;
wire wire6815;
wire wire6820;
wire wire6821;
wire wire6826;
wire wire6827;
wire wire6830;
wire wire6831;
wire wire6833;
wire wire6838;
wire wire6839;
wire wire6844;
wire wire6845;
wire wire6850;
wire wire6851;
wire wire6856;
wire wire6857;
wire wire6862;
wire wire6863;
wire wire6867;
wire wire6869;
wire wire6874;
wire wire6875;
wire wire6880;
wire wire6881;
wire wire6885;
wire wire6886;
wire wire6887;
wire wire6892;
wire wire6893;
wire wire6898;
wire wire6899;
wire wire6904;
wire wire6905;
wire wire6910;
wire wire6911;
wire wire6916;
wire wire6917;
wire wire6922;
wire wire6923;
wire wire6928;
wire wire6929;
wire wire6934;
wire wire6935;
wire wire6940;
wire wire6941;
wire wire6946;
wire wire6947;
wire wire6952;
wire wire6953;
wire wire6958;
wire wire6959;
wire wire6962;
wire wire6963;
wire wire6964;
wire wire6967;
wire wire6968;
wire wire6969;
wire wire6973;
wire wire6974;
wire wire6977;
wire wire6978;
wire wire6979;
wire wire6982;
wire wire6984;
wire wire6987;
wire wire6989;
wire wire6992;
wire wire6994;
wire wire6997;
wire wire6998;
wire wire6999;
wire wire7003;
wire wire7004;
wire wire7008;
wire wire7009;
wire wire7013;
wire wire7014;
wire wire7017;
wire wire7018;
wire wire7019;
wire wire7022;
wire wire7023;
wire wire7024;
wire wire7028;
wire wire7029;
wire wire7033;
wire wire7034;
wire wire7037;
wire wire7038;
wire wire7039;
wire wire7042;
wire wire7044;
wire wire7047;
wire wire7049;
wire wire7052;
wire wire7054;
wire wire7056;
wire wire7057;
wire wire7059;
wire wire7063;
wire wire7064;
wire wire7068;
wire wire7069;
wire wire7072;
wire wire7073;
wire wire7078;
wire wire7079;
wire wire7083;
wire wire7084;
wire wire7086;
wire wire7087;
wire wire7088;
wire wire7091;
wire wire7092;
wire wire7095;
wire wire7096;
wire wire7099;
wire wire7100;
wire wire7103;
wire wire7104;
wire wire7106;
wire wire7108;
wire wire7110;
wire wire7111;
wire wire7112;
wire wire7114;
wire wire7115;
wire wire7116;
wire wire7117;
wire wire7118;
wire wire7119;
wire wire7120;
wire wire7127;
wire wire7128;
wire wire7129;
wire wire7130;
wire wire7131;
wire wire7135;
wire wire7136;
wire wire7137;
wire wire7138;
wire wire7139;
wire wire7140;
wire wire7141;
wire wire7145;
wire wire7148;
wire wire7149;
wire wire7150;
wire wire7151;
wire wire7152;
wire wire7154;
wire wire7155;
wire wire7156;
wire wire7159;
wire wire7161;
wire wire7162;
wire wire7164;
wire wire7173;
wire wire7174;
wire wire7175;
wire wire7176;
wire wire7178;
wire wire7179;
wire wire7190;
wire wire7191;
wire wire7192;
wire wire7193;
wire wire7194;
wire wire7195;
wire wire7199;
wire wire7200;
wire wire7202;
wire wire7203;
wire wire7204;
wire wire7205;
wire wire7206;
wire wire7207;
wire wire7208;
wire wire7209;
wire wire7210;
wire wire7211;
wire wire7212;
wire wire7213;
wire wire7214;
wire wire7215;
wire wire7216;
wire wire7217;
wire wire7218;
wire wire7228;
wire wire7229;
wire wire7230;
wire wire7231;
wire wire7232;
wire wire7235;
wire wire7240;
wire wire7241;
wire wire7243;
wire wire7245;
wire wire7246;
wire wire7249;
wire wire7250;
wire wire7254;
wire wire7255;
wire wire7257;
wire wire7261;
wire wire7263;
wire wire7264;
wire wire7268;
wire wire7269;
wire wire7271;
wire wire7276;
wire wire7277;
wire wire7278;
wire wire7282;
wire wire7283;
wire wire7285;
wire wire7290;
wire wire7291;
wire wire7292;
wire wire7297;
wire wire7298;
wire wire7299;
wire wire7304;
wire wire7305;
wire wire7311;
wire wire7312;
wire wire7313;
wire wire7318;
wire wire7319;
wire wire7320;
wire wire7325;
wire wire7326;
wire wire7327;
wire wire7332;
wire wire7333;
wire wire7334;
wire wire7339;
wire wire7340;
wire wire7341;
wire wire7345;
wire wire7346;
wire wire7348;
wire wire7353;
wire wire7354;
wire wire7355;
wire wire7360;
wire wire7361;
wire wire7362;
wire wire7367;
wire wire7368;
wire wire7369;
wire wire7374;
wire wire7375;
wire wire7376;
wire wire7381;
wire wire7382;
wire wire7383;
wire wire7388;
wire wire7389;
wire wire7395;
wire wire7396;
wire wire7402;
wire wire7403;
wire wire7409;
wire wire7410;
wire wire7416;
wire wire7417;
wire wire7421;
wire wire7422;
wire wire7423;
wire wire7424;
wire wire7428;
wire wire7429;
wire wire7430;
wire wire7433;
wire wire7434;
wire wire7436;
wire wire7440;
wire wire7442;
wire wire7446;
wire wire7448;
wire wire7453;
wire wire7454;
wire wire7459;
wire wire7460;
wire wire7465;
wire wire7466;
wire wire7471;
wire wire7472;
wire wire7477;
wire wire7478;
wire wire7481;
wire wire7482;
wire wire7483;
wire wire7484;
wire wire7489;
wire wire7490;
wire wire7494;
wire wire7495;
wire wire7501;
wire wire7502;
wire wire7505;
wire wire7506;
wire wire7508;
wire wire7513;
wire wire7514;
wire wire7519;
wire wire7520;
wire wire7522;
wire wire7523;
wire wire7526;
wire wire7529;
wire wire7530;
wire wire7531;
wire wire7532;
wire wire7537;
wire wire7538;
wire wire7542;
wire wire7543;
wire wire7549;
wire wire7550;
wire wire7555;
wire wire7556;
wire wire7560;
wire wire7561;
wire wire7567;
wire wire7568;
wire wire7573;
wire wire7574;
wire wire7579;
wire wire7580;
wire wire7585;
wire wire7586;
wire wire7591;
wire wire7592;
wire wire7597;
wire wire7598;
wire wire7601;
wire wire7602;
wire wire7604;
wire wire7607;
wire wire7608;
wire wire7610;
wire wire7613;
wire wire7614;
wire wire7616;
wire wire7621;
wire wire7622;
wire wire7626;
wire wire7627;
wire wire7632;
wire wire7633;
wire wire7638;
wire wire7639;
wire wire7645;
wire wire7646;
wire wire7650;
wire wire7651;
wire wire7656;
wire wire7657;
wire wire7662;
wire wire7663;
wire wire7664;
wire wire7668;
wire wire7669;
wire wire7675;
wire wire7676;
wire wire7681;
wire wire7682;
wire wire7686;
wire wire7687;
wire wire7693;
wire wire7694;
wire wire7699;
wire wire7700;
wire wire7705;
wire wire7706;
wire wire7711;
wire wire7712;
wire wire7717;
wire wire7718;
wire wire7723;
wire wire7724;
wire wire7727;
wire wire7728;
wire wire7729;
wire wire7732;
wire wire7733;
wire wire7734;
wire wire7737;
wire wire7738;
wire wire7739;
wire wire7741;
wire wire7742;
wire wire7744;
wire wire7747;
wire wire7748;
wire wire7749;
wire wire7752;
wire wire7753;
wire wire7754;
wire wire7757;
wire wire7758;
wire wire7759;
wire wire7762;
wire wire7763;
wire wire7764;
wire wire7766;
wire wire7767;
wire wire7768;
wire wire7769;
wire wire7772;
wire wire7773;
wire wire7774;
wire wire7777;
wire wire7778;
wire wire7779;
wire wire7782;
wire wire7783;
wire wire7784;
wire wire7786;
wire wire7787;
wire wire7789;
wire wire7792;
wire wire7794;
wire wire7797;
wire wire7799;
wire wire7802;
wire wire7803;
wire wire7804;
wire wire7808;
wire wire7809;
wire wire7811;
wire wire7812;
wire wire7814;
wire wire7817;
wire wire7818;
wire wire7819;
wire wire7821;
wire wire7822;
wire wire7824;
wire wire7828;
wire wire7829;
wire wire7833;
wire wire7834;
wire wire7836;
wire wire7837;
wire wire7839;
wire wire7842;
wire wire7843;
wire wire7847;
wire wire7848;
wire wire7851;
wire wire7853;
wire wire7856;
wire wire7857;
wire wire7860;
wire wire7861;
wire wire7864;
wire wire7865;
wire wire7868;
wire wire7869;
wire wire7872;
wire wire7873;
wire wire7876;
wire wire7877;
wire wire7880;
wire wire7881;
wire wire7884;
wire wire7886;
wire wire7887;
wire wire7889;
wire wire7890;
wire wire7892;
wire wire7894;
wire wire7895;
wire wire7896;
wire wire7897;
wire wire7902;
wire wire7903;
wire wire7904;
wire wire7905;
wire wire7908;
wire wire7909;
wire wire7910;
wire wire7911;
wire wire7912;
wire wire7913;
wire wire7915;
wire wire7916;
wire wire7917;
wire wire7918;
wire wire7921;
wire wire7922;
wire wire7923;
wire wire7924;
wire wire7925;
wire wire7926;
wire wire7927;
wire wire7930;
wire wire7933;
wire wire7935;
wire wire7936;
wire wire7937;
wire wire7939;
wire wire7945;
wire wire7946;
wire wire7947;
wire wire7949;
wire wire7959;
wire wire7960;
wire wire7961;
wire wire7962;
wire wire7964;
wire wire7965;
wire wire7968;
wire wire7969;
wire wire7970;
wire wire7971;
wire wire7972;
wire wire7973;
wire wire7974;
wire wire7975;
wire wire7976;
wire wire7977;
wire wire7978;
wire wire7979;
wire wire7980;
wire wire7981;
wire wire7982;
wire wire7983;
wire wire7984;
wire wire7985;
wire wire7986;
wire wire7987;
wire wire7988;
wire wire7998;
wire wire8000;
wire wire8001;
wire wire8002;
wire wire8003;
wire wire8004;
wire wire8006;
wire wire8012;
wire wire8013;
wire wire8015;
wire wire8019;
wire wire8021;
wire wire8022;
wire wire8026;
wire wire8027;
wire wire8029;
wire wire8032;
wire wire8033;
wire wire8035;
wire wire8036;
wire wire8040;
wire wire8041;
wire wire8043;
wire wire8048;
wire wire8049;
wire wire8050;
wire wire8054;
wire wire8056;
wire wire8057;
wire wire8062;
wire wire8063;
wire wire8064;
wire wire8069;
wire wire8070;
wire wire8075;
wire wire8076;
wire wire8078;
wire wire8083;
wire wire8084;
wire wire8090;
wire wire8091;
wire wire8092;
wire wire8097;
wire wire8098;
wire wire8099;
wire wire8104;
wire wire8105;
wire wire8106;
wire wire8111;
wire wire8112;
wire wire8113;
wire wire8118;
wire wire8119;
wire wire8120;
wire wire8125;
wire wire8126;
wire wire8132;
wire wire8133;
wire wire8139;
wire wire8140;
wire wire8146;
wire wire8147;
wire wire8153;
wire wire8154;
wire wire8160;
wire wire8161;
wire wire8167;
wire wire8168;
wire wire8174;
wire wire8175;
wire wire8180;
wire wire8181;
wire wire8182;
wire wire8186;
wire wire8187;
wire wire8188;
wire wire8192;
wire wire8193;
wire wire8194;
wire wire8198;
wire wire8199;
wire wire8200;
wire wire8202;
wire wire8203;
wire wire8206;
wire wire8209;
wire wire8211;
wire wire8212;
wire wire8216;
wire wire8218;
wire wire8222;
wire wire8223;
wire wire8224;
wire wire8229;
wire wire8230;
wire wire8235;
wire wire8236;
wire wire8240;
wire wire8242;
wire wire8246;
wire wire8248;
wire wire8252;
wire wire8254;
wire wire8258;
wire wire8259;
wire wire8260;
wire wire8265;
wire wire8266;
wire wire8269;
wire wire8270;
wire wire8272;
wire wire8277;
wire wire8278;
wire wire8281;
wire wire8282;
wire wire8284;
wire wire8287;
wire wire8289;
wire wire8290;
wire wire8294;
wire wire8295;
wire wire8296;
wire wire8299;
wire wire8301;
wire wire8302;
wire wire8305;
wire wire8306;
wire wire8308;
wire wire8313;
wire wire8314;
wire wire8319;
wire wire8320;
wire wire8325;
wire wire8326;
wire wire8331;
wire wire8332;
wire wire8337;
wire wire8338;
wire wire8342;
wire wire8343;
wire wire8348;
wire wire8349;
wire wire8354;
wire wire8356;
wire wire8360;
wire wire8361;
wire wire8367;
wire wire8368;
wire wire8372;
wire wire8373;
wire wire8378;
wire wire8379;
wire wire8385;
wire wire8386;
wire wire8391;
wire wire8392;
wire wire8397;
wire wire8398;
wire wire8403;
wire wire8404;
wire wire8409;
wire wire8410;
wire wire8415;
wire wire8416;
wire wire8421;
wire wire8422;
wire wire8427;
wire wire8428;
wire wire8433;
wire wire8434;
wire wire8437;
wire wire8438;
wire wire8439;
wire wire8442;
wire wire8443;
wire wire8444;
wire wire8447;
wire wire8448;
wire wire8449;
wire wire8452;
wire wire8453;
wire wire8454;
wire wire8456;
wire wire8457;
wire wire8459;
wire wire8462;
wire wire8463;
wire wire8464;
wire wire8467;
wire wire8468;
wire wire8469;
wire wire8472;
wire wire8473;
wire wire8474;
wire wire8477;
wire wire8478;
wire wire8479;
wire wire8482;
wire wire8483;
wire wire8484;
wire wire8487;
wire wire8488;
wire wire8489;
wire wire8492;
wire wire8493;
wire wire8494;
wire wire8496;
wire wire8497;
wire wire8499;
wire wire8501;
wire wire8502;
wire wire8504;
wire wire8506;
wire wire8507;
wire wire8509;
wire wire8512;
wire wire8514;
wire wire8518;
wire wire8519;
wire wire8522;
wire wire8523;
wire wire8524;
wire wire8526;
wire wire8527;
wire wire8529;
wire wire8531;
wire wire8532;
wire wire8534;
wire wire8537;
wire wire8539;
wire wire8543;
wire wire8544;
wire wire8548;
wire wire8549;
wire wire8552;
wire wire8553;
wire wire8558;
wire wire8559;
wire wire8562;
wire wire8563;
wire wire8568;
wire wire8569;
wire wire8571;
wire wire8572;
wire wire8573;
wire wire8575;
wire wire8576;
wire wire8577;
wire wire8580;
wire wire8581;
wire wire8584;
wire wire8585;
wire wire8587;
wire wire8588;
wire wire8589;
wire wire8591;
wire wire8592;
wire wire8593;
wire wire8596;
wire wire8597;
wire wire8600;
wire wire8601;
wire wire8604;
wire wire8605;
wire wire8608;
wire wire8609;
wire wire8612;
wire wire8613;
wire wire8616;
wire wire8617;
wire wire8620;
wire wire8621;
wire wire8624;
wire wire8626;
wire wire8627;
wire wire8630;
wire wire8631;
wire wire8633;
wire wire8635;
wire wire8637;
wire wire8638;
wire wire8639;
wire wire8640;
wire wire8647;
wire wire8648;
wire wire8649;
wire wire8650;
wire wire8651;
wire wire8652;
wire wire8656;
wire wire8657;
wire wire8658;
wire wire8659;
wire wire8660;
wire wire8661;
wire wire8664;
wire wire8665;
wire wire8666;
wire wire8668;
wire wire8670;
wire wire8671;
wire wire8672;
wire wire8674;
wire wire8675;
wire wire8676;
wire wire8677;
wire wire8680;
wire wire8687;
wire wire8688;
wire wire8689;
wire wire8691;
wire wire8698;
wire wire8699;
wire wire8700;
wire wire8701;
wire wire8704;
wire wire8705;
wire wire8706;
wire wire8707;
wire wire8708;
wire wire8709;
wire wire8710;
wire wire8711;
wire wire8712;
wire wire8713;
wire wire8714;
wire wire8715;
wire wire8716;
wire wire8717;
wire wire8718;
wire wire8719;
wire wire8720;
wire wire8721;
wire wire8722;
wire wire8723;
wire wire8724;
wire wire8725;
wire wire8726;
wire wire8727;
wire wire8728;
wire wire8741;
wire wire8742;
wire wire8743;
wire wire8744;
wire wire8745;
wire wire8746;
wire wire8750;
wire wire8755;
wire wire8756;
wire wire8758;
wire wire8763;
wire wire8764;
wire wire8765;
wire wire8769;
wire wire8770;
wire wire8772;
wire wire8776;
wire wire8777;
wire wire8779;
wire wire8783;
wire wire8784;
wire wire8786;
wire wire8791;
wire wire8792;
wire wire8793;
wire wire8798;
wire wire8799;
wire wire8802;
wire wire8803;
wire wire8805;
wire wire8806;
wire wire8809;
wire wire8810;
wire wire8812;
wire wire8815;
wire wire8816;
wire wire8818;
wire wire8820;
wire wire8821;
wire wire8824;
wire wire8828;
wire wire8830;
wire wire8833;
wire wire8835;
wire wire8836;
wire wire8840;
wire wire8841;
wire wire8842;
wire wire8846;
wire wire8847;
wire wire8848;
wire wire8852;
wire wire8854;
wire wire8859;
wire wire8860;
wire wire8864;
wire wire8866;
wire wire8870;
wire wire8871;
wire wire8877;
wire wire8878;
wire wire8882;
wire wire8883;
wire wire8887;
wire wire8888;
wire wire8889;
wire wire8890;
wire wire8893;
wire wire8894;
wire wire8895;
wire wire8898;
wire wire8899;
wire wire8900;
wire wire8902;
wire wire8904;
wire wire8905;
wire wire8908;
wire wire8909;
wire wire8910;
wire wire8913;
wire wire8914;
wire wire8915;
wire wire8918;
wire wire8919;
wire wire8920;
wire wire8923;
wire wire8924;
wire wire8925;
wire wire8927;
wire wire8928;
wire wire8930;
wire wire8932;
wire wire8933;
wire wire8935;
wire wire8938;
wire wire8940;
wire wire8943;
wire wire8944;
wire wire8945;
wire wire8948;
wire wire8949;
wire wire8950;
wire wire8954;
wire wire8955;
wire wire8959;
wire wire8960;
wire wire8964;
wire wire8965;
wire wire8969;
wire wire8970;
wire wire8974;
wire wire8975;
wire wire8979;
wire wire8980;
wire wire8983;
wire wire8984;
wire wire8989;
wire wire8990;
wire wire8993;
wire wire8994;
wire wire8995;
wire wire8998;
wire wire8999;
wire wire9004;
wire wire9005;
wire wire9010;
wire wire9012;
wire wire9013;
wire wire9014;
wire wire9017;
wire wire9018;
wire wire9021;
wire wire9022;
wire wire9025;
wire wire9026;
wire wire9029;
wire wire9030;
wire wire9032;
wire wire9033;
wire wire9034;
wire wire9035;
wire wire9036;
wire wire9037;
wire wire9038;
wire wire9040;
wire wire9041;
wire wire9042;
wire wire9044;
wire wire9045;
wire wire9046;
wire wire9049;
wire wire9050;
wire wire9053;
wire wire9057;
wire wire9058;
wire wire9059;
wire wire9060;
wire wire9061;
wire wire9063;
wire wire9064;
wire wire9066;
wire wire9067;
wire wire9070;
wire wire9072;
wire wire9073;
wire wire9075;
wire wire9076;
wire wire9079;
wire wire9081;
wire wire9082;
wire wire9084;
wire wire9085;
wire wire9087;
wire wire9088;
wire wire9089;
wire wire9090;
wire wire9092;
wire wire9094;
wire wire9096;
wire wire9097;
wire wire9098;
wire wire9099;
wire wire9101;
wire wire9104;
wire wire9105;
wire wire9109;
wire wire9110;
wire wire9121;
wire wire9122;
wire wire9123;
wire wire9124;
wire wire9125;
wire wire9128;
wire wire9129;
wire wire9131;
wire wire9132;
wire wire9133;
wire wire9134;
wire wire9135;
wire wire9136;
wire wire9137;
wire wire9138;
wire wire9139;
wire wire9140;
wire wire9141;
wire wire9142;
wire wire9143;
wire wire9144;
wire wire9145;
wire wire9146;
wire wire9155;
wire wire9156;
wire wire9157;
wire wire9158;
wire wire9161;
reg n_n852;

reg n_n853;

reg n_n854;

reg n_n855;

reg n_n856;

reg n_n857;

reg n_n858;

reg n_n859;

always  @(posedge clock)
	n_n852<=n_n45;

 always  @(posedge clock)
	n_n853<=n_n46;

 always  @(posedge clock)
	n_n854<=n_n47;

 always  @(posedge clock)
	n_n855<=n_n48;

 always  @(posedge clock)
	n_n856<=n_n49;

 always  @(posedge clock)
	n_n857<=n_n50;

 always  @(posedge clock)
	n_n858<=n_n51;

 always  @(posedge clock)
	n_n859<=n_n52;

 assign s298_out_0_ = ( wire578 ) | ( wire579 ) ;
 assign s298_out_1_ = ( wire581 ) | ( wire582 ) | ( (~ s298_out_3_)  &  wire5524 ) ;
 assign s298_out_2_ = ( wire619 ) | ( wire621 ) | ( wire622 ) ;
 assign s298_out_3_ = ( (~ n_n856)  &  n_n857  &  n_n858  &  (~ n_n859) ) ;
 assign s298_out_4_ = ( wire621 ) | ( wire622 ) ;
 assign s298_out_5_ = ( wire623 ) | ( (~ n_n858)  &  n_n859 ) | ( (~ n_n857)  &  n_n858  &  (~ n_n859) ) ;
 assign n_n45 = ( wire7230 ) | ( wire7231 ) | ( wire7235 ) ;
 assign n_n46 = ( wire8000 ) | ( wire8001 ) | ( wire8004 ) | ( wire8006 ) ;
 assign n_n47 = ( wire8745 ) | ( wire8746 ) | ( wire8750 ) ;
 assign n_n48 = ( wire9156 ) | ( wire9157 ) | ( wire9161 ) ;
 assign n_n49 = ( wire6371 ) | ( wire6372 ) | ( wire6376 ) ;
 assign n_n50 = ( wire6016 ) | ( wire6017 ) | ( wire6018 ) ;
 assign n_n51 = ( wire5700 ) | ( wire5701 ) | ( wire5702 ) | ( wire5703 ) ;
 assign n_n52 = ( wire5783 ) | ( wire5784 ) | ( wire5790 ) | ( wire5791 ) ;
 assign wire24 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8758 ) ;
 assign wire25 = ( (~ wire6371)  &  (~ wire6372)  &  (~ wire6376)  &  wire8765 ) ;
 assign wire27 = ( wire5789  &  wire8779 ) | ( wire5790  &  wire8779 ) | ( wire5791  &  wire8779 ) ;
 assign wire29 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8793 ) ;
 assign wire30 = ( n_n856  &  n_n858  &  wire8798  &  wire8799 ) ;
 assign wire39 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8854 ) ;
 assign wire40 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8860 ) ;
 assign wire41 = ( wire6016  &  wire8866 ) | ( wire6017  &  wire8866 ) | ( wire6018  &  wire8866 ) ;
 assign wire42 = ( (~ wire578)  &  (~ wire579)  &  wire8870  &  wire8871 ) ;
 assign wire44 = ( wire621  &  wire8882  &  wire8883 ) | ( wire622  &  wire8882  &  wire8883 ) ;
 assign wire45 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8890 ) ;
 assign wire57 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8950 ) ;
 assign wire58 = ( wire580  &  wire8955 ) | ( wire581  &  wire8955 ) | ( wire582  &  wire8955 ) ;
 assign wire59 = ( wire580  &  wire8960 ) | ( wire581  &  wire8960 ) | ( wire582  &  wire8960 ) ;
 assign wire60 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8965 ) ;
 assign wire61 = ( wire6016  &  wire8970 ) | ( wire6017  &  wire8970 ) | ( wire6018  &  wire8970 ) ;
 assign wire62 = ( wire6016  &  wire8975 ) | ( wire6017  &  wire8975 ) | ( wire6018  &  wire8975 ) ;
 assign wire63 = ( wire6016  &  wire8980 ) | ( wire6017  &  wire8980 ) | ( wire6018  &  wire8980 ) ;
 assign wire66 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8995 ) ;
 assign wire68 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire9005 ) ;
 assign wire69 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire9010 ) ;
 assign wire76 = ( wire6016  &  wire9038 ) | ( wire6017  &  wire9038 ) | ( wire6018  &  wire9038 ) ;
 assign wire77 = ( wire6016  &  wire9042 ) | ( wire6017  &  wire9042 ) | ( wire6018  &  wire9042 ) ;
 assign wire78 = ( wire6016  &  wire9046 ) | ( wire6017  &  wire9046 ) | ( wire6018  &  wire9046 ) ;
 assign wire79 = ( wire6016  &  wire9050 ) | ( wire6017  &  wire9050 ) | ( wire6018  &  wire9050 ) ;
 assign wire80 = ( n_n51  &  wire578  &  wire9053 ) | ( n_n51  &  wire579  &  wire9053 ) ;
 assign wire81 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire9058 ) ;
 assign wire86 = ( wire6016  &  wire9073 ) | ( wire6017  &  wire9073 ) | ( wire6018  &  wire9073 ) ;
 assign wire87 = ( wire6016  &  wire9076 ) | ( wire6017  &  wire9076 ) | ( wire6018  &  wire9076 ) ;
 assign wire88 = ( wire6016  &  wire9079 ) | ( wire6017  &  wire9079 ) | ( wire6018  &  wire9079 ) ;
 assign wire89 = ( wire6016  &  wire9082 ) | ( wire6017  &  wire9082 ) | ( wire6018  &  wire9082 ) ;
 assign wire90 = ( wire6016  &  wire9085 ) | ( wire6017  &  wire9085 ) | ( wire6018  &  wire9085 ) ;
 assign wire91 = ( wire6016  &  wire9088 ) | ( wire6017  &  wire9088 ) | ( wire6018  &  wire9088 ) ;
 assign wire94 = ( s298_in_2_  &  wire6016 ) | ( s298_in_2_  &  wire6017 ) | ( s298_in_2_  &  wire6018 ) ;
 assign wire101 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8057 ) ;
 assign wire102 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8064 ) ;
 assign wire103 = ( (~ n_n51)  &  (~ wire578)  &  (~ wire579)  &  wire8070 ) ;
 assign wire104 = ( wire5789  &  wire8078 ) | ( wire5790  &  wire8078 ) | ( wire5791  &  wire8078 ) ;
 assign wire107 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8099 ) ;
 assign wire108 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8106 ) ;
 assign wire109 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8113 ) ;
 assign wire110 = ( wire5789  &  wire8120 ) | ( wire5790  &  wire8120 ) | ( wire5791  &  wire8120 ) ;
 assign wire111 = ( (~ n_n856)  &  n_n857  &  wire8125  &  wire8126 ) ;
 assign wire112 = ( (~ n_n855)  &  (~ n_n856)  &  wire8132  &  wire8133 ) ;
 assign wire113 = ( n_n855  &  (~ n_n857)  &  wire8139  &  wire8140 ) ;
 assign wire114 = ( (~ n_n855)  &  n_n858  &  wire8146  &  wire8147 ) ;
 assign wire115 = ( (~ n_n855)  &  n_n856  &  wire8153  &  wire8154 ) ;
 assign wire116 = ( n_n855  &  (~ n_n856)  &  wire8160  &  wire8161 ) ;
 assign wire117 = ( n_n855  &  n_n856  &  wire8167  &  wire8168 ) ;
 assign wire118 = ( n_n856  &  n_n857  &  wire8174  &  wire8175 ) ;
 assign wire133 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8266 ) ;
 assign wire134 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8272 ) ;
 assign wire135 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8278 ) ;
 assign wire136 = ( wire6016  &  wire8284 ) | ( wire6017  &  wire8284 ) | ( wire6018  &  wire8284 ) ;
 assign wire137 = ( wire6016  &  wire8290 ) | ( wire6017  &  wire8290 ) | ( wire6018  &  wire8290 ) ;
 assign wire138 = ( wire6016  &  wire8296 ) | ( wire6017  &  wire8296 ) | ( wire6018  &  wire8296 ) ;
 assign wire139 = ( wire5789  &  wire8302 ) | ( wire5790  &  wire8302 ) | ( wire5791  &  wire8302 ) ;
 assign wire140 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8308 ) ;
 assign wire148 = ( wire5789  &  wire8356 ) | ( wire5790  &  wire8356 ) | ( wire5791  &  wire8356 ) ;
 assign wire153 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8386 ) ;
 assign wire154 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8392 ) ;
 assign wire155 = ( wire5789  &  wire8398 ) | ( wire5790  &  wire8398 ) | ( wire5791  &  wire8398 ) ;
 assign wire156 = ( wire619  &  wire8404 ) | ( wire621  &  wire8404 ) | ( wire622  &  wire8404 ) ;
 assign wire161 = ( wire8433  &  wire8434 ) ;
 assign wire179 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8524 ) ;
 assign wire180 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8529 ) ;
 assign wire181 = ( wire6016  &  wire8534 ) | ( wire6017  &  wire8534 ) | ( wire6018  &  wire8534 ) ;
 assign wire182 = ( wire6016  &  wire8539 ) | ( wire6017  &  wire8539 ) | ( wire6018  &  wire8539 ) ;
 assign wire202 = ( (~ s298_in_1_)  &  s298_out_3_  &  (~ n_n852)  &  wire8624 ) ;
 assign wire204 = ( wire6016  &  wire8631 ) | ( wire6017  &  wire8631 ) | ( wire6018  &  wire8631 ) ;
 assign wire206 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8635 ) ;
 assign wire210 = ( (~ wire6371)  &  (~ wire6372)  &  (~ wire6376)  &  wire7250 ) ;
 assign wire214 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire7278 ) ;
 assign wire215 = ( wire6016  &  wire7285 ) | ( wire6017  &  wire7285 ) | ( wire6018  &  wire7285 ) ;
 assign wire216 = ( wire6016  &  wire7292 ) | ( wire6017  &  wire7292 ) | ( wire6018  &  wire7292 ) ;
 assign wire217 = ( wire6016  &  wire7299 ) | ( wire6017  &  wire7299 ) | ( wire6018  &  wire7299 ) ;
 assign wire218 = ( (~ wire578)  &  (~ wire579)  &  wire7304  &  wire7305 ) ;
 assign wire224 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7348 ) ;
 assign wire226 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7362 ) ;
 assign wire227 = ( wire5789  &  wire7369 ) | ( wire5790  &  wire7369 ) | ( wire5791  &  wire7369 ) ;
 assign wire228 = ( wire5789  &  wire7376 ) | ( wire5790  &  wire7376 ) | ( wire5791  &  wire7376 ) ;
 assign wire229 = ( wire5789  &  wire7383 ) | ( wire5790  &  wire7383 ) | ( wire5791  &  wire7383 ) ;
 assign wire230 = ( (~ s298_out_3_)  &  wire7388  &  wire7389 ) ;
 assign wire231 = ( n_n857  &  n_n858  &  wire7395  &  wire7396 ) ;
 assign wire232 = ( (~ n_n856)  &  (~ n_n857)  &  wire7402  &  wire7403 ) ;
 assign wire233 = ( n_n856  &  n_n857  &  wire7409  &  wire7410 ) ;
 assign wire234 = ( n_n856  &  (~ n_n857)  &  wire7416  &  wire7417 ) ;
 assign wire249 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7508 ) ;
 assign wire250 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7514 ) ;
 assign wire251 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7520 ) ;
 assign wire252 = ( wire6016  &  wire7526 ) | ( wire6017  &  wire7526 ) | ( wire6018  &  wire7526 ) ;
 assign wire253 = ( wire6016  &  wire7532 ) | ( wire6017  &  wire7532 ) | ( wire6018  &  wire7532 ) ;
 assign wire254 = ( wire6016  &  wire7538 ) | ( wire6017  &  wire7538 ) | ( wire6018  &  wire7538 ) ;
 assign wire265 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7604 ) ;
 assign wire266 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7610 ) ;
 assign wire267 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7616 ) ;
 assign wire269 = ( wire621  &  wire7626  &  wire7627 ) | ( wire622  &  wire7626  &  wire7627 ) ;
 assign wire278 = ( wire5789  &  wire7682 ) | ( wire5790  &  wire7682 ) | ( wire5791  &  wire7682 ) ;
 assign wire279 = ( (~ s298_out_3_)  &  wire7686  &  wire7687 ) ;
 assign wire303 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7814 ) ;
 assign wire304 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7819 ) ;
 assign wire305 = ( wire6016  &  wire7824 ) | ( wire6017  &  wire7824 ) | ( wire6018  &  wire7824 ) ;
 assign wire306 = ( wire6016  &  wire7829 ) | ( wire6017  &  wire7829 ) | ( wire6018  &  wire7829 ) ;
 assign wire307 = ( wire6016  &  wire7834 ) | ( wire6017  &  wire7834 ) | ( wire6018  &  wire7834 ) ;
 assign wire308 = ( wire5789  &  wire7839 ) | ( wire5790  &  wire7839 ) | ( wire5791  &  wire7839 ) ;
 assign wire309 = ( wire578  &  wire7842  &  wire7843 ) | ( wire579  &  wire7842  &  wire7843 ) ;
 assign wire320 = ( wire6016  &  wire7887 ) | ( wire6017  &  wire7887 ) | ( wire6018  &  wire7887 ) ;
 assign wire321 = ( wire6016  &  wire7890 ) | ( wire6017  &  wire7890 ) | ( wire6018  &  wire7890 ) ;
 assign wire322 = ( wire6371  &  wire7892 ) | ( wire6372  &  wire7892 ) | ( wire6376  &  wire7892 ) ;
 assign wire323 = ( wire6016  &  wire7894 ) | ( wire6017  &  wire7894 ) | ( wire6018  &  wire7894 ) ;
 assign wire324 = ( (~ wire6371)  &  (~ wire6372)  &  (~ wire6376)  &  wire6384 ) ;
 assign wire325 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6392 ) ;
 assign wire334 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire6456 ) ;
 assign wire335 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire6463 ) ;
 assign wire336 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6470 ) ;
 assign wire337 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6477 ) ;
 assign wire338 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6484 ) ;
 assign wire339 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6491 ) ;
 assign wire340 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6498 ) ;
 assign wire341 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6505 ) ;
 assign wire342 = ( wire6016  &  wire6512 ) | ( wire6017  &  wire6512 ) | ( wire6018  &  wire6512 ) ;
 assign wire344 = ( wire5789  &  wire6526 ) | ( wire5790  &  wire6526 ) | ( wire5791  &  wire6526 ) ;
 assign wire346 = ( wire5789  &  wire6540 ) | ( wire5790  &  wire6540 ) | ( wire5791  &  wire6540 ) ;
 assign wire347 = ( (~ wire621)  &  (~ wire622)  &  wire6545  &  wire6546 ) ;
 assign wire351 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6575 ) ;
 assign wire353 = ( wire5789  &  wire6589 ) | ( wire5790  &  wire6589 ) | ( wire5791  &  wire6589 ) ;
 assign wire355 = ( wire5789  &  wire6603 ) | ( wire5790  &  wire6603 ) | ( wire5791  &  wire6603 ) ;
 assign wire359 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6631 ) ;
 assign wire360 = ( wire619  &  wire6638 ) | ( wire621  &  wire6638 ) | ( wire622  &  wire6638 ) ;
 assign wire361 = ( (~ n_n856)  &  (~ n_n857)  &  wire6643  &  wire6644 ) ;
 assign wire362 = ( (~ n_n855)  &  (~ n_n856)  &  wire6650  &  wire6651 ) ;
 assign wire363 = ( n_n856  &  (~ n_n857)  &  wire6657  &  wire6658 ) ;
 assign wire364 = ( (~ n_n855)  &  (~ n_n856)  &  wire6664  &  wire6665 ) ;
 assign wire365 = ( n_n855  &  (~ n_n856)  &  wire6671  &  wire6672 ) ;
 assign wire366 = ( n_n855  &  (~ n_n856)  &  wire6678  &  wire6679 ) ;
 assign wire367 = ( (~ n_n855)  &  n_n857  &  wire6685  &  wire6686 ) ;
 assign wire368 = ( n_n856  &  n_n857  &  wire6692  &  wire6693 ) ;
 assign wire369 = ( n_n856  &  n_n857  &  wire6699  &  wire6700 ) ;
 assign wire384 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6791 ) ;
 assign wire385 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6797 ) ;
 assign wire386 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6803 ) ;
 assign wire387 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6809 ) ;
 assign wire388 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6815 ) ;
 assign wire391 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6833 ) ;
 assign wire397 = ( wire5789  &  wire6869 ) | ( wire5790  &  wire6869 ) | ( wire5791  &  wire6869 ) ;
 assign wire398 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6875 ) ;
 assign wire399 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6881 ) ;
 assign wire400 = ( wire5789  &  wire6887 ) | ( wire5790  &  wire6887 ) | ( wire5791  &  wire6887 ) ;
 assign wire401 = ( wire5789  &  wire6893 ) | ( wire5790  &  wire6893 ) | ( wire5791  &  wire6893 ) ;
 assign wire402 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire6899 ) ;
 assign wire403 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire6905 ) ;
 assign wire424 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7019 ) ;
 assign wire425 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7024 ) ;
 assign wire426 = ( wire580  &  wire7029 ) | ( wire581  &  wire7029 ) | ( wire582  &  wire7029 ) ;
 assign wire427 = ( wire580  &  wire7034 ) | ( wire581  &  wire7034 ) | ( wire582  &  wire7034 ) ;
 assign wire428 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7039 ) ;
 assign wire429 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7044 ) ;
 assign wire430 = ( wire6016  &  wire7049 ) | ( wire6017  &  wire7049 ) | ( wire6018  &  wire7049 ) ;
 assign wire431 = ( wire6016  &  wire7054 ) | ( wire6017  &  wire7054 ) | ( wire6018  &  wire7054 ) ;
 assign wire432 = ( wire5789  &  wire7059 ) | ( wire5790  &  wire7059 ) | ( wire5791  &  wire7059 ) ;
 assign wire436 = ( wire5789  &  wire7079 ) | ( wire5790  &  wire7079 ) | ( wire5791  &  wire7079 ) ;
 assign wire441 = ( wire6371  &  wire7100 ) | ( wire6372  &  wire7100 ) | ( wire6376  &  wire7100 ) ;
 assign wire442 = ( wire580  &  wire7104 ) | ( wire581  &  wire7104 ) | ( wire582  &  wire7104 ) ;
 assign wire443 = ( wire6016  &  wire7108 ) | ( wire6017  &  wire7108 ) | ( wire6018  &  wire7108 ) ;
 assign wire444 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7112 ) ;
 assign wire445 = ( wire6016  &  wire7115 ) | ( wire6017  &  wire7115 ) | ( wire6018  &  wire7115 ) ;
 assign wire446 = ( n_n855  &  (~ n_n856)  &  wire5518  &  wire5519 ) ;
 assign wire447 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5798 ) ;
 assign wire448 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6025 ) ;
 assign wire449 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6031 ) ;
 assign wire450 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6037 ) ;
 assign wire451 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6043 ) ;
 assign wire452 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6049 ) ;
 assign wire453 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6055 ) ;
 assign wire454 = ( wire6016  &  wire6061 ) | ( wire6017  &  wire6061 ) | ( wire6018  &  wire6061 ) ;
 assign wire455 = ( wire6016  &  wire6067 ) | ( wire6017  &  wire6067 ) | ( wire6018  &  wire6067 ) ;
 assign wire457 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6079 ) ;
 assign wire458 = ( wire621  &  wire6083  &  wire6084 ) | ( wire622  &  wire6083  &  wire6084 ) ;
 assign wire462 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6109 ) ;
 assign wire463 = ( wire5789  &  wire6115 ) | ( wire5790  &  wire6115 ) | ( wire5791  &  wire6115 ) ;
 assign wire464 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire6121 ) ;
 assign wire470 = ( wire580  &  wire6155 ) | ( wire581  &  wire6155 ) | ( wire582  &  wire6155 ) ;
 assign wire471 = ( wire580  &  wire6160 ) | ( wire581  &  wire6160 ) | ( wire582  &  wire6160 ) ;
 assign wire472 = ( wire6016  &  wire6165 ) | ( wire6017  &  wire6165 ) | ( wire6018  &  wire6165 ) ;
 assign wire473 = ( wire6016  &  wire6170 ) | ( wire6017  &  wire6170 ) | ( wire6018  &  wire6170 ) ;
 assign wire474 = ( wire6016  &  wire6175 ) | ( wire6017  &  wire6175 ) | ( wire6018  &  wire6175 ) ;
 assign wire475 = ( wire6016  &  wire6180 ) | ( wire6017  &  wire6180 ) | ( wire6018  &  wire6180 ) ;
 assign wire476 = ( wire6016  &  wire6185 ) | ( wire6017  &  wire6185 ) | ( wire6018  &  wire6185 ) ;
 assign wire477 = ( wire6016  &  wire6190 ) | ( wire6017  &  wire6190 ) | ( wire6018  &  wire6190 ) ;
 assign wire478 = ( wire6016  &  wire6195 ) | ( wire6017  &  wire6195 ) | ( wire6018  &  wire6195 ) ;
 assign wire479 = ( wire5789  &  wire6200 ) | ( wire5790  &  wire6200 ) | ( wire5791  &  wire6200 ) ;
 assign wire483 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6220 ) ;
 assign wire484 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6225 ) ;
 assign wire485 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6230 ) ;
 assign wire494 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6274 ) ;
 assign wire495 = ( wire580  &  wire6278 ) | ( wire581  &  wire6278 ) | ( wire582  &  wire6278 ) ;
 assign wire496 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6282 ) ;
 assign wire497 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6286 ) ;
 assign wire498 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6290 ) ;
 assign wire499 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6294 ) ;
 assign wire500 = ( wire6016  &  wire6298 ) | ( wire6017  &  wire6298 ) | ( wire6018  &  wire6298 ) ;
 assign wire501 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire6302 ) ;
 assign wire504 = ( wire6016  &  wire6313 ) | ( wire6017  &  wire6313 ) | ( wire6018  &  wire6313 ) ;
 assign wire505 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6315 ) ;
 assign wire506 = ( s298_out_0_  &  (~ n_n855)  &  (~ n_n857)  &  n_n51 ) ;
 assign wire507 = ( wire578  &  wire5803  &  wire5804 ) | ( wire579  &  wire5803  &  wire5804 ) ;
 assign wire510 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5824 ) ;
 assign wire511 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5830 ) ;
 assign wire513 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5842 ) ;
 assign wire518 = ( wire5789  &  wire5868 ) | ( wire5790  &  wire5868 ) | ( wire5791  &  wire5868 ) ;
 assign wire519 = ( wire5789  &  wire5873 ) | ( wire5790  &  wire5873 ) | ( wire5791  &  wire5873 ) ;
 assign wire526 = ( wire5789  &  wire5907 ) | ( wire5790  &  wire5907 ) | ( wire5791  &  wire5907 ) ;
 assign wire531 = ( wire5789  &  wire5927 ) | ( wire5790  &  wire5927 ) | ( wire5791  &  wire5927 ) ;
 assign wire532 = ( wire621  &  wire5929  &  wire5930 ) | ( wire622  &  wire5929  &  wire5930 ) ;
 assign wire535 = ( wire5789  &  wire5943 ) | ( wire5790  &  wire5943 ) | ( wire5791  &  wire5943 ) ;
 assign wire536 = ( wire5789  &  wire5947 ) | ( wire5790  &  wire5947 ) | ( wire5791  &  wire5947 ) ;
 assign wire542 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5967 ) ;
 assign wire544 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire5973 ) ;
 assign wire550 = ( wire621  &  wire5537  &  wire5538 ) | ( wire622  &  wire5537  &  wire5538 ) ;
 assign wire553 = ( (~ s298_out_3_)  &  n_n854  &  (~ n_n856)  &  wire5712 ) ;
 assign wire556 = ( (~ wire578)  &  (~ wire579)  &  wire5726 ) ;
 assign wire558 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire5732 ) ;
 assign wire566 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire5748 ) ;
 assign wire567 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire5750 ) ;
 assign wire568 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire5752 ) ;
 assign wire570 = ( n_n852  &  (~ n_n853)  &  (~ n_n854)  &  (~ n_n858) ) ;
 assign wire571 = ( n_n853  &  n_n855  &  n_n857  &  (~ n_n858) ) ;
 assign wire576 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire5763 ) ;
 assign wire577 = ( (~ n_n855)  &  (~ n_n857)  &  (~ n_n858) ) ;
 assign wire578 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire5723 ) ;
 assign wire579 = ( (~ n_n858)  &  n_n859 ) | ( n_n857  &  n_n859  &  wire5509 ) ;
 assign wire580 = ( (~ s298_out_3_)  &  n_n855  &  n_n858  &  (~ n_n859) ) ;
 assign wire581 = ( wire623  &  wire5525 ) | ( wire624  &  wire5525 ) | ( wire625  &  wire5525 ) ;
 assign wire582 = ( wire623  &  wire5526 ) | ( wire624  &  wire5526 ) | ( wire625  &  wire5526 ) ;
 assign wire611 = ( (~ n_n852)  &  n_n853  &  (~ n_n854)  &  (~ n_n859) ) ;
 assign wire612 = ( n_n852  &  (~ n_n854)  &  n_n857  &  (~ n_n859) ) ;
 assign wire613 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n854)  &  (~ n_n859) ) ;
 assign wire614 = ( (~ n_n854)  &  n_n856  &  (~ n_n857)  &  (~ n_n859) ) ;
 assign wire615 = ( n_n853  &  n_n855  &  n_n857  &  (~ n_n859) ) ;
 assign wire616 = ( n_n854  &  (~ n_n858)  &  (~ n_n859) ) ;
 assign wire619 = ( (~ n_n857)  &  n_n858  &  n_n859 ) | ( n_n857  &  n_n858  &  (~ n_n859) ) | ( n_n857  &  n_n858  &  (~ wire5509) ) | ( n_n858  &  n_n859  &  (~ wire5509) ) ;
 assign wire621 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire5513 ) ;
 assign wire622 = ( (~ n_n857)  &  n_n858  &  n_n859 ) | ( n_n858  &  n_n859  &  (~ wire5509) ) ;
 assign wire623 = ( (~ n_n855)  &  n_n856  &  n_n857  &  n_n859 ) ;
 assign wire624 = ( (~ n_n857)  &  n_n858  &  (~ n_n859) ) ;
 assign wire625 = ( (~ n_n858)  &  n_n859 ) ;
 assign wire5509 = ( n_n856  &  (~ n_n855) ) ;
 assign wire5513 = ( n_n857  &  n_n856 ) ;
 assign wire5518 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire5519 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire5524 = ( n_n855  &  n_n858  &  (~ n_n859) ) ;
 assign wire5525 = ( (~ n_n859)  &  (~ n_n854) ) ;
 assign wire5526 = ( (~ n_n859)  &  (~ n_n856) ) ;
 assign wire5530 = ( (~ s298_in_0_)  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire5531 = ( wire621  &  wire5530 ) | ( wire622  &  wire5530 ) ;
 assign wire5533 = ( n_n855  &  (~ n_n854) ) ;
 assign wire5534 = ( n_n852  &  n_n853  &  (~ n_n856) ) ;
 assign wire5537 = ( n_n854  &  (~ n_n853) ) ;
 assign wire5538 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n859) ) ;
 assign wire5541 = ( n_n856  &  n_n855 ) ;
 assign wire5542 = ( n_n853  &  n_n854  &  (~ n_n857) ) ;
 assign wire5548 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire5549 = ( (~ n_n853)  &  n_n854  &  n_n856  &  (~ n_n859) ) ;
 assign wire5554 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire5555 = ( (~ n_n854)  &  (~ n_n855)  &  n_n856  &  n_n857 ) ;
 assign wire5560 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire5561 = ( (~ n_n854)  &  (~ n_n855)  &  n_n856  &  n_n857 ) ;
 assign wire5566 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire5567 = ( n_n854  &  (~ n_n855)  &  n_n856  &  n_n857 ) ;
 assign wire5572 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire5573 = ( n_n854  &  (~ n_n855)  &  n_n856  &  n_n857 ) ;
 assign wire5578 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire5579 = ( n_n854  &  n_n855  &  n_n856  &  (~ n_n858) ) ;
 assign wire5582 = ( (~ n_n859)  &  (~ n_n857) ) ;
 assign wire5583 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n853)  &  n_n855 ) ;
 assign wire5586 = ( (~ n_n859)  &  (~ n_n855) ) ;
 assign wire5587 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire5590 = ( (~ n_n859)  &  n_n856 ) ;
 assign wire5591 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire5594 = ( (~ n_n858)  &  n_n857 ) ;
 assign wire5595 = ( (~ n_n852)  &  (~ n_n853)  &  (~ n_n854)  &  (~ n_n856) ) ;
 assign wire5599 = ( (~ n_n852)  &  (~ n_n853)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire5603 = ( (~ n_n852)  &  (~ n_n853)  &  n_n854  &  (~ n_n855) ) ;
 assign wire5606 = ( n_n857  &  n_n856 ) ;
 assign wire5607 = ( n_n852  &  n_n853  &  n_n854  &  (~ n_n855) ) ;
 assign wire5610 = ( (~ n_n858)  &  n_n856 ) ;
 assign wire5611 = ( (~ s298_in_2_)  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire5615 = ( n_n852  &  n_n854  &  n_n855  &  n_n856 ) ;
 assign wire5619 = ( n_n852  &  n_n854  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire5623 = ( n_n853  &  n_n854  &  n_n855  &  n_n856 ) ;
 assign wire5627 = ( (~ s298_in_2_)  &  n_n853  &  n_n854  &  n_n856 ) ;
 assign wire5630 = ( (~ n_n858)  &  n_n857 ) ;
 assign wire5631 = ( n_n853  &  n_n854  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire5633 = ( (~ n_n857)  &  n_n855 ) ;
 assign wire5634 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n859) ) ;
 assign wire5636 = ( n_n858  &  (~ n_n856) ) ;
 assign wire5637 = ( (~ n_n854)  &  (~ n_n855)  &  (~ n_n859) ) ;
 assign wire5639 = ( (~ n_n855)  &  n_n853 ) ;
 assign wire5640 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n859) ) ;
 assign wire5642 = ( (~ n_n857)  &  (~ n_n856) ) ;
 assign wire5643 = ( n_n852  &  (~ n_n855)  &  (~ n_n859) ) ;
 assign wire5645 = ( (~ n_n856)  &  (~ n_n855) ) ;
 assign wire5646 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n859) ) ;
 assign wire5648 = ( (~ n_n857)  &  (~ n_n856) ) ;
 assign wire5649 = ( n_n853  &  (~ n_n855)  &  (~ n_n859) ) ;
 assign wire5651 = ( n_n858  &  n_n857 ) ;
 assign wire5652 = ( (~ n_n855)  &  n_n856  &  n_n859 ) ;
 assign wire5655 = ( n_n852  &  (~ n_n854)  &  n_n858 ) ;
 assign wire5658 = ( n_n853  &  (~ n_n854)  &  n_n858 ) ;
 assign wire5675 = ( n_n855  &  n_n856  &  (~ n_n859) ) | ( n_n855  &  (~ n_n858)  &  (~ n_n859) ) ;
 assign wire5676 = ( wire5548  &  wire5549 ) | ( wire5554  &  wire5555 ) ;
 assign wire5677 = ( wire5560  &  wire5561 ) | ( wire5566  &  wire5567 ) ;
 assign wire5678 = ( wire5572  &  wire5573 ) | ( wire5578  &  wire5579 ) ;
 assign wire5679 = ( wire5582  &  wire5583 ) | ( wire5586  &  wire5587 ) ;
 assign wire5680 = ( wire5590  &  wire5591 ) | ( wire5594  &  wire5595 ) ;
 assign wire5681 = ( n_n857  &  (~ n_n858)  &  wire5599 ) | ( n_n857  &  n_n858  &  wire5603 ) ;
 assign wire5682 = ( wire5606  &  wire5607 ) | ( wire5610  &  wire5611 ) ;
 assign wire5683 = ( (~ n_n857)  &  (~ n_n858)  &  wire5615 ) | ( n_n857  &  (~ n_n858)  &  wire5619 ) ;
 assign wire5684 = ( (~ n_n857)  &  (~ n_n858)  &  wire5623 ) | ( (~ n_n857)  &  (~ n_n858)  &  wire5627 ) ;
 assign wire5685 = ( wire5630  &  wire5631 ) | ( wire5633  &  wire5634 ) ;
 assign wire5686 = ( wire5636  &  wire5637 ) | ( wire5639  &  wire5640 ) ;
 assign wire5687 = ( wire5642  &  wire5643 ) | ( wire5645  &  wire5646 ) ;
 assign wire5688 = ( wire5648  &  wire5649 ) | ( wire5651  &  wire5652 ) ;
 assign wire5689 = ( (~ n_n855)  &  n_n857  &  wire5655 ) | ( (~ n_n855)  &  n_n857  &  wire5658 ) ;
 assign wire5690 = ( wire611 ) | ( wire612 ) | ( wire613 ) | ( wire614 ) ;
 assign wire5691 = ( wire615 ) | ( wire616 ) | ( wire5675 ) ;
 assign wire5700 = ( wire5676 ) | ( wire5677 ) | ( wire5678 ) | ( wire5679 ) ;
 assign wire5701 = ( wire5680 ) | ( wire5681 ) | ( wire5682 ) | ( wire5683 ) ;
 assign wire5702 = ( wire5684 ) | ( wire5685 ) | ( wire5686 ) | ( wire5687 ) ;
 assign wire5703 = ( wire5688 ) | ( wire5689 ) | ( wire5690 ) | ( wire5691 ) ;
 assign wire5707 = ( (~ n_n855)  &  n_n854 ) ;
 assign wire5708 = ( (~ n_n852)  &  (~ n_n853)  &  (~ n_n856) ) ;
 assign wire5712 = ( (~ n_n852)  &  (~ n_n853)  &  n_n857 ) ;
 assign wire5717 = ( n_n852  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire5719 = ( (~ n_n854)  &  (~ n_n855)  &  n_n858 ) ;
 assign wire5720 = ( (~ wire621)  &  (~ wire622)  &  wire5719 ) ;
 assign wire5723 = ( n_n854  &  n_n856  &  n_n858  &  (~ n_n859) ) ;
 assign wire5725 = ( n_n852  &  (~ n_n855)  &  n_n857 ) ;
 assign wire5726 = ( wire619  &  wire5725 ) | ( wire621  &  wire5725 ) | ( wire622  &  wire5725 ) ;
 assign wire5729 = ( n_n853  &  (~ n_n855)  &  (~ n_n856)  &  n_n857 ) ;
 assign wire5732 = ( (~ n_n853)  &  n_n854  &  n_n855  &  (~ n_n859) ) ;
 assign wire5734 = ( (~ n_n852)  &  (~ n_n855)  &  (~ n_n858) ) ;
 assign wire5736 = ( s298_in_0_  &  (~ n_n852)  &  (~ n_n858) ) ;
 assign wire5738 = ( (~ n_n853)  &  n_n856  &  (~ n_n858) ) ;
 assign wire5740 = ( (~ s298_in_1_)  &  (~ n_n852)  &  wire621 ) | ( (~ s298_in_1_)  &  (~ n_n852)  &  wire622 ) ;
 assign wire5741 = ( (~ n_n853)  &  (~ n_n852) ) ;
 assign wire5744 = ( n_n852  &  n_n853  &  (~ n_n859) ) ;
 assign wire5746 = ( (~ n_n852)  &  (~ n_n857)  &  n_n859 ) ;
 assign wire5748 = ( s298_in_1_  &  (~ n_n857)  &  (~ n_n859) ) ;
 assign wire5750 = ( (~ s298_in_0_)  &  n_n852  &  (~ n_n858) ) ;
 assign wire5752 = ( (~ s298_in_1_)  &  (~ n_n856)  &  (~ n_n858) ) ;
 assign wire5754 = ( (~ n_n854)  &  (~ n_n856)  &  n_n857 ) ;
 assign wire5759 = ( s298_in_2_  &  wire621 ) | ( s298_in_2_  &  wire622 ) ;
 assign wire5763 = ( (~ n_n858)  &  s298_in_2_ ) ;
 assign wire5766 = ( wire577 ) | ( n_n856  &  (~ n_n857)  &  wire5717 ) ;
 assign wire5767 = ( wire553 ) | ( wire570 ) | ( wire571 ) ;
 assign wire5768 = ( wire5766 ) | ( (~ s298_out_5_)  &  wire5541  &  wire5542 ) ;
 assign wire5772 = ( wire566 ) | ( wire567 ) | ( wire568 ) | ( wire576 ) ;
 assign wire5774 = ( wire5772 ) | ( s298_out_1_  &  wire5531 ) ;
 assign wire5775 = ( (~ s298_out_1_)  &  wire5720 ) | ( s298_out_1_  &  wire5533  &  wire5534 ) ;
 assign wire5776 = ( wire550 ) | ( wire558 ) | ( wire5767 ) | ( wire5768 ) ;
 assign wire5777 = ( (~ n_n51)  &  wire5754 ) | ( (~ n_n51)  &  wire5707  &  wire5708 ) ;
 assign wire5780 = ( (~ wire578)  &  (~ wire579)  &  wire5729 ) | ( (~ wire578)  &  (~ wire579)  &  wire5734 ) ;
 assign wire5781 = ( (~ wire578)  &  (~ wire579)  &  wire5736 ) | ( (~ wire578)  &  (~ wire579)  &  wire5738 ) ;
 assign wire5782 = ( s298_out_0_  &  wire5740 ) | ( s298_out_0_  &  (~ n_n51)  &  wire5741 ) ;
 assign wire5783 = ( wire578  &  wire5744 ) | ( wire579  &  wire5744 ) | ( wire578  &  wire5746 ) | ( wire579  &  wire5746 ) ;
 assign wire5784 = ( s298_out_0_  &  wire5759 ) | ( s298_out_0_  &  (~ n_n51)  &  (~ n_n859) ) ;
 assign wire5785 = ( s298_out_0_  &  (~ n_n854)  &  (~ n_n51) ) | ( s298_out_0_  &  n_n855  &  (~ n_n51) ) ;
 assign wire5787 = ( wire556 ) | ( wire5776 ) | ( wire5780 ) ;
 assign wire5789 = ( wire5784 ) | ( wire5783 ) ;
 assign wire5790 = ( wire5774 ) | ( wire5775 ) | ( wire5777 ) | ( wire5785 ) ;
 assign wire5791 = ( wire5781 ) | ( wire5782 ) | ( wire5787 ) ;
 assign wire5796 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire5797 = ( n_n855  &  (~ n_n856)  &  wire5796 ) ;
 assign wire5798 = ( wire580  &  wire5797 ) | ( wire581  &  wire5797 ) | ( wire582  &  wire5797 ) ;
 assign wire5803 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire5804 = ( (~ n_n854)  &  n_n855  &  n_n856  &  (~ n_n857) ) ;
 assign wire5810 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire5811 = ( n_n854  &  n_n856  &  (~ n_n857)  &  (~ n_n858) ) ;
 assign wire5817 = ( s298_in_1_  &  (~ n_n852)  &  n_n854  &  n_n856 ) ;
 assign wire5818 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857  &  wire5817 ) ;
 assign wire5821 = ( n_n857  &  (~ n_n854) ) ;
 assign wire5822 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n853 ) ;
 assign wire5824 = ( wire621  &  wire5821  &  wire5822 ) | ( wire622  &  wire5821  &  wire5822 ) ;
 assign wire5827 = ( n_n856  &  n_n854 ) ;
 assign wire5828 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire5830 = ( wire621  &  wire5827  &  wire5828 ) | ( wire622  &  wire5827  &  wire5828 ) ;
 assign wire5834 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire5835 = ( s298_in_1_  &  (~ n_n853)  &  (~ n_n855)  &  n_n858 ) ;
 assign wire5841 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire5842 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire5841 ) ;
 assign wire5847 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n852  &  n_n854 ) ;
 assign wire5848 = ( (~ n_n855)  &  n_n856  &  (~ n_n857)  &  n_n858 ) ;
 assign wire5850 = ( (~ n_n855)  &  n_n854 ) ;
 assign wire5851 = ( (~ s298_in_2_)  &  n_n852  &  n_n856 ) ;
 assign wire5853 = ( wire621  &  wire5850  &  wire5851 ) | ( wire622  &  wire5850  &  wire5851 ) ;
 assign wire5856 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n857 ) ;
 assign wire5858 = ( (~ s298_out_3_)  &  n_n853  &  (~ n_n854)  &  wire5856 ) ;
 assign wire5861 = ( (~ s298_in_2_)  &  (~ n_n853)  &  n_n857 ) ;
 assign wire5862 = ( (~ n_n854)  &  (~ n_n856)  &  wire5861 ) ;
 assign wire5865 = ( (~ n_n854)  &  n_n853 ) ;
 assign wire5866 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n856 ) ;
 assign wire5868 = ( wire578  &  wire5865  &  wire5866 ) | ( wire579  &  wire5865  &  wire5866 ) ;
 assign wire5870 = ( (~ n_n856)  &  n_n854 ) ;
 assign wire5871 = ( (~ s298_in_2_)  &  n_n853  &  n_n857 ) ;
 assign wire5873 = ( wire578  &  wire5870  &  wire5871 ) | ( wire579  &  wire5870  &  wire5871 ) ;
 assign wire5877 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire5878 = ( (~ n_n856)  &  (~ n_n857)  &  wire5877 ) ;
 assign wire5882 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire5883 = ( (~ n_n857)  &  (~ n_n858)  &  wire5882 ) ;
 assign wire5886 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n856 ) ;
 assign wire5887 = ( n_n854  &  n_n855  &  wire5886 ) ;
 assign wire5892 = ( (~ n_n852)  &  (~ n_n853)  &  n_n854  &  (~ n_n855) ) ;
 assign wire5893 = ( n_n858  &  (~ n_n859)  &  wire5892 ) ;
 assign wire5897 = ( n_n852  &  n_n853  &  n_n854  &  n_n856 ) ;
 assign wire5898 = ( n_n857  &  (~ n_n858)  &  wire5897 ) ;
 assign wire5902 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire5903 = ( (~ n_n853)  &  n_n854  &  n_n855  &  n_n856 ) ;
 assign wire5905 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n855) ) ;
 assign wire5906 = ( wire619  &  wire5905 ) | ( wire621  &  wire5905 ) | ( wire622  &  wire5905 ) ;
 assign wire5907 = ( (~ wire578)  &  (~ wire579)  &  wire5906 ) ;
 assign wire5910 = ( (~ s298_in_2_)  &  (~ n_n853)  &  n_n857 ) ;
 assign wire5911 = ( n_n854  &  n_n856  &  wire5910 ) ;
 assign wire5914 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire5915 = ( (~ n_n852)  &  (~ n_n853)  &  wire5914 ) ;
 assign wire5918 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n857) ) ;
 assign wire5919 = ( (~ n_n854)  &  (~ n_n856)  &  wire5918 ) ;
 assign wire5922 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n858) ) ;
 assign wire5923 = ( n_n853  &  (~ n_n857)  &  wire5922 ) ;
 assign wire5925 = ( (~ s298_in_2_)  &  n_n852  &  n_n858 ) ;
 assign wire5927 = ( n_n51  &  (~ wire621)  &  (~ wire622)  &  wire5925 ) ;
 assign wire5929 = ( (~ n_n855)  &  (~ n_n854) ) ;
 assign wire5930 = ( (~ s298_in_2_)  &  n_n853  &  n_n856 ) ;
 assign wire5934 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire5938 = ( (~ s298_in_2_)  &  n_n852  &  n_n856 ) ;
 assign wire5939 = ( (~ n_n854)  &  n_n855  &  wire5938 ) ;
 assign wire5942 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n857 ) ;
 assign wire5943 = ( (~ n_n853)  &  n_n854  &  wire5942 ) ;
 assign wire5946 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n857) ) ;
 assign wire5947 = ( n_n855  &  n_n856  &  wire5946 ) ;
 assign wire5950 = ( n_n857  &  n_n856 ) ;
 assign wire5951 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire5954 = ( n_n858  &  n_n857 ) ;
 assign wire5955 = ( (~ s298_in_2_)  &  (~ n_n854)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire5957 = ( (~ s298_in_2_)  &  n_n855  &  n_n857 ) ;
 assign wire5961 = ( (~ s298_in_2_)  &  n_n854  &  n_n857  &  (~ n_n858) ) ;
 assign wire5963 = ( n_n852  &  n_n853  &  (~ n_n857) ) ;
 assign wire5966 = ( (~ n_n854)  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire5967 = ( wire578  &  wire5966 ) | ( wire579  &  wire5966 ) ;
 assign wire5970 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n853  &  (~ n_n859) ) ;
 assign wire5972 = ( (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire5973 = ( (~ wire621)  &  (~ wire622)  &  wire5972 ) ;
 assign wire5976 = ( n_n852  &  (~ n_n854)  &  n_n855  &  n_n857 ) ;
 assign wire5978 = ( (~ n_n854)  &  n_n855  &  wire621 ) | ( (~ n_n854)  &  n_n855  &  wire622 ) ;
 assign wire5980 = ( n_n853  &  n_n855  &  n_n857 ) ;
 assign wire5981 = ( wire5847  &  wire5848 ) | ( wire5902  &  wire5903 ) ;
 assign wire5982 = ( wire5950  &  wire5951 ) | ( wire5954  &  wire5955 ) ;
 assign wire5984 = ( (~ s298_out_5_)  &  wire5893 ) | ( (~ s298_out_5_)  &  wire5834  &  wire5835 ) ;
 assign wire5986 = ( wire532 ) | ( wire5981 ) | ( wire5982 ) | ( wire5984 ) ;
 assign wire5987 = ( wire5986 ) | ( (~ n_n51)  &  wire5810  &  wire5811 ) ;
 assign wire5988 = ( n_n51  &  wire5898 ) | ( (~ s298_out_5_)  &  n_n51  &  wire5887 ) ;
 assign wire5989 = ( n_n51  &  wire5939 ) | ( s298_out_3_  &  n_n51  &  wire5934 ) ;
 assign wire5990 = ( n_n51  &  wire5976 ) | ( n_n51  &  wire5978 ) ;
 assign wire5992 = ( (~ wire578)  &  (~ wire579)  &  wire5818 ) | ( (~ wire578)  &  (~ wire579)  &  wire5853 ) ;
 assign wire5993 = ( (~ s298_out_0_)  &  wire5858 ) | ( s298_out_0_  &  (~ n_n51)  &  wire5862 ) ;
 assign wire5994 = ( wire578  &  wire5878 ) | ( wire579  &  wire5878 ) | ( wire578  &  wire5883 ) | ( wire579  &  wire5883 ) ;
 assign wire5995 = ( wire578  &  wire5915 ) | ( wire579  &  wire5915 ) | ( (~ wire578)  &  (~ wire579)  &  wire5911 ) ;
 assign wire5996 = ( wire578  &  wire5919 ) | ( wire579  &  wire5919 ) | ( wire578  &  wire5923 ) | ( wire579  &  wire5923 ) ;
 assign wire5997 = ( (~ s298_out_0_)  &  wire5961 ) | ( (~ s298_out_0_)  &  n_n51  &  wire5957 ) ;
 assign wire5998 = ( s298_out_0_  &  wire5970 ) | ( s298_out_0_  &  n_n51  &  wire5963 ) ;
 assign wire6001 = ( wire507 ) | ( wire5992 ) | ( n_n51  &  wire5980 ) ;
 assign wire6005 = ( wire5987 ) | ( wire5988 ) | ( wire5989 ) | ( wire5990 ) ;
 assign wire6006 = ( wire5993 ) | ( wire5994 ) | ( wire6001 ) ;
 assign wire6007 = ( wire5995 ) | ( wire5996 ) | ( wire5997 ) | ( wire5998 ) ;
 assign wire6009 = ( wire6005 ) | ( wire6006 ) | ( wire6007 ) ;
 assign wire6016 = ( wire510 ) | ( wire511 ) | ( wire513 ) | ( wire518 ) ;
 assign wire6017 = ( wire519 ) | ( wire526 ) | ( wire531 ) | ( wire535 ) ;
 assign wire6018 = ( wire536 ) | ( wire542 ) | ( wire544 ) | ( wire6009 ) ;
 assign wire6022 = ( n_n855  &  (~ n_n853) ) ;
 assign wire6023 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6025 = ( wire578  &  wire6022  &  wire6023 ) | ( wire579  &  wire6022  &  wire6023 ) ;
 assign wire6028 = ( n_n858  &  (~ n_n855) ) ;
 assign wire6029 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n853  &  (~ n_n854) ) ;
 assign wire6031 = ( (~ wire621)  &  (~ wire622)  &  wire6028  &  wire6029 ) ;
 assign wire6033 = ( n_n854  &  s298_in_1_ ) ;
 assign wire6034 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856 ) ;
 assign wire6036 = ( wire621  &  wire6033  &  wire6034 ) | ( wire622  &  wire6033  &  wire6034 ) ;
 assign wire6037 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6036 ) ;
 assign wire6040 = ( n_n854  &  n_n853 ) ;
 assign wire6041 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6043 = ( wire621  &  wire6040  &  wire6041 ) | ( wire622  &  wire6040  &  wire6041 ) ;
 assign wire6046 = ( n_n856  &  n_n853 ) ;
 assign wire6047 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6049 = ( wire621  &  wire6046  &  wire6047 ) | ( wire622  &  wire6046  &  wire6047 ) ;
 assign wire6053 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6054 = ( n_n856  &  n_n857  &  n_n858 ) | ( n_n857  &  n_n858  &  n_n859 ) ;
 assign wire6055 = ( wire6054  &  wire6053 ) ;
 assign wire6058 = ( n_n857  &  (~ n_n856) ) ;
 assign wire6059 = ( s298_in_0_  &  s298_in_1_  &  n_n854  &  n_n855 ) ;
 assign wire6061 = ( wire578  &  wire6058  &  wire6059 ) | ( wire579  &  wire6058  &  wire6059 ) ;
 assign wire6065 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n853  &  n_n854 ) ;
 assign wire6066 = ( n_n856  &  n_n858  &  (~ n_n859) ) | ( (~ n_n857)  &  n_n858  &  (~ n_n859) ) ;
 assign wire6067 = ( wire6066  &  wire6065 ) ;
 assign wire6072 = ( s298_in_1_  &  n_n852  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6073 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire6072 ) ;
 assign wire6076 = ( n_n857  &  (~ n_n854) ) ;
 assign wire6077 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n852  &  (~ n_n853) ) ;
 assign wire6079 = ( wire621  &  wire6076  &  wire6077 ) | ( wire622  &  wire6076  &  wire6077 ) ;
 assign wire6083 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire6084 = ( s298_in_1_  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire6090 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n855 ) ;
 assign wire6091 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire6090 ) ;
 assign wire6095 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire6096 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n855 ) ;
 assign wire6101 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire6102 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  n_n857 ) ;
 assign wire6108 = ( n_n852  &  n_n853  &  (~ n_n854)  &  n_n856 ) ;
 assign wire6109 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire6108 ) ;
 assign wire6114 = ( (~ s298_in_1_)  &  n_n852  &  n_n854  &  (~ n_n856) ) ;
 assign wire6115 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire6114 ) ;
 assign wire6120 = ( (~ s298_in_1_)  &  n_n852  &  n_n854  &  n_n855 ) ;
 assign wire6121 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire6120 ) ;
 assign wire6126 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6127 = ( (~ n_n853)  &  (~ n_n854)  &  n_n856  &  (~ n_n858) ) ;
 assign wire6132 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6133 = ( n_n853  &  (~ n_n854)  &  n_n856  &  (~ n_n858) ) ;
 assign wire6138 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n854) ) ;
 assign wire6139 = ( (~ n_n855)  &  n_n856  &  n_n857  &  (~ n_n858) ) ;
 assign wire6144 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6145 = ( (~ n_n855)  &  n_n856  &  n_n857  &  (~ n_n858) ) ;
 assign wire6148 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n854 ) ;
 assign wire6149 = ( n_n852  &  n_n853  &  wire6148 ) ;
 assign wire6150 = ( wire580  &  wire6149 ) | ( wire581  &  wire6149 ) | ( wire582  &  wire6149 ) ;
 assign wire6154 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6155 = ( (~ n_n855)  &  (~ n_n856)  &  wire6154 ) ;
 assign wire6159 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  (~ n_n853) ) ;
 assign wire6160 = ( n_n854  &  (~ n_n855)  &  wire6159 ) ;
 assign wire6162 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n857) ) ;
 assign wire6164 = ( n_n51  &  wire578  &  wire6162 ) | ( n_n51  &  wire579  &  wire6162 ) ;
 assign wire6165 = ( wire5789  &  wire6164 ) | ( wire5790  &  wire6164 ) | ( wire5791  &  wire6164 ) ;
 assign wire6167 = ( (~ n_n854)  &  n_n852 ) ;
 assign wire6168 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n855 ) ;
 assign wire6170 = ( wire578  &  wire6167  &  wire6168 ) | ( wire579  &  wire6167  &  wire6168 ) ;
 assign wire6172 = ( n_n855  &  n_n854 ) ;
 assign wire6173 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n856) ) ;
 assign wire6175 = ( wire621  &  wire6172  &  wire6173 ) | ( wire622  &  wire6172  &  wire6173 ) ;
 assign wire6178 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n859) ) ;
 assign wire6180 = ( (~ s298_out_5_)  &  n_n852  &  (~ n_n857)  &  wire6178 ) ;
 assign wire6183 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n854 ) ;
 assign wire6184 = ( n_n852  &  (~ n_n853)  &  wire6183 ) ;
 assign wire6185 = ( wire5789  &  wire6184 ) | ( wire5790  &  wire6184 ) | ( wire5791  &  wire6184 ) ;
 assign wire6189 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n854  &  (~ n_n855) ) ;
 assign wire6190 = ( (~ n_n856)  &  (~ n_n857)  &  wire6189 ) ;
 assign wire6194 = ( (~ s298_in_2_)  &  n_n852  &  n_n855  &  n_n856 ) ;
 assign wire6195 = ( n_n857  &  (~ n_n858)  &  wire6194 ) ;
 assign wire6197 = ( (~ n_n856)  &  n_n855 ) ;
 assign wire6198 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n857) ) ;
 assign wire6200 = ( (~ wire578)  &  (~ wire579)  &  wire6197  &  wire6198 ) ;
 assign wire6203 = ( (~ s298_in_2_)  &  n_n852  &  n_n857 ) ;
 assign wire6204 = ( (~ n_n854)  &  n_n856  &  wire6203 ) ;
 assign wire6209 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire6210 = ( n_n857  &  (~ n_n858)  &  wire6209 ) ;
 assign wire6214 = ( (~ s298_in_2_)  &  n_n852  &  n_n854  &  n_n855 ) ;
 assign wire6215 = ( (~ n_n856)  &  (~ n_n857)  &  wire6214 ) ;
 assign wire6217 = ( (~ n_n854)  &  n_n852 ) ;
 assign wire6218 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n857 ) ;
 assign wire6220 = ( wire621  &  wire6217  &  wire6218 ) | ( wire622  &  wire6217  &  wire6218 ) ;
 assign wire6222 = ( n_n854  &  n_n853 ) ;
 assign wire6223 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n857 ) ;
 assign wire6225 = ( wire621  &  wire6222  &  wire6223 ) | ( wire622  &  wire6222  &  wire6223 ) ;
 assign wire6227 = ( (~ n_n855)  &  n_n854 ) ;
 assign wire6228 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n856) ) ;
 assign wire6230 = ( wire621  &  wire6227  &  wire6228 ) | ( wire622  &  wire6227  &  wire6228 ) ;
 assign wire6234 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6235 = ( (~ n_n856)  &  (~ n_n857)  &  wire6234 ) ;
 assign wire6238 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n856 ) ;
 assign wire6239 = ( (~ n_n854)  &  (~ n_n855)  &  wire6238 ) ;
 assign wire6244 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6245 = ( n_n855  &  (~ n_n858)  &  wire6244 ) ;
 assign wire6248 = ( (~ n_n858)  &  n_n856 ) ;
 assign wire6249 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n855) ) ;
 assign wire6254 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6255 = ( n_n855  &  n_n856  &  wire6254 ) ;
 assign wire6258 = ( n_n857  &  (~ n_n856) ) ;
 assign wire6259 = ( (~ s298_in_2_)  &  n_n853  &  n_n854  &  n_n855 ) ;
 assign wire6264 = ( (~ s298_in_2_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n855 ) ;
 assign wire6265 = ( (~ n_n856)  &  n_n857  &  wire6264 ) ;
 assign wire6269 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire6270 = ( s298_in_1_  &  n_n854  &  n_n857  &  (~ n_n858) ) ;
 assign wire6273 = ( (~ s298_in_2_)  &  n_n852  &  n_n854  &  n_n856 ) ;
 assign wire6274 = ( wire580  &  wire6273 ) | ( wire581  &  wire6273 ) | ( wire582  &  wire6273 ) ;
 assign wire6277 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855) ) ;
 assign wire6278 = ( (~ n_n852)  &  n_n853  &  wire6277 ) ;
 assign wire6280 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire6282 = ( n_n51  &  wire578  &  wire6280 ) | ( n_n51  &  wire579  &  wire6280 ) ;
 assign wire6285 = ( (~ s298_in_2_)  &  n_n854  &  (~ n_n855)  &  n_n856 ) ;
 assign wire6286 = ( wire621  &  wire6285 ) | ( wire622  &  wire6285 ) ;
 assign wire6289 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n855)  &  n_n856 ) ;
 assign wire6290 = ( wire621  &  wire6289 ) | ( wire622  &  wire6289 ) ;
 assign wire6293 = ( (~ s298_in_2_)  &  n_n856  &  (~ n_n857)  &  (~ n_n858) ) ;
 assign wire6294 = ( (~ n_n51)  &  wire6293 ) ;
 assign wire6297 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n859) ) ;
 assign wire6298 = ( n_n854  &  (~ n_n855)  &  wire6297 ) ;
 assign wire6301 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6302 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire6301 ) ;
 assign wire6305 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n858) ) ;
 assign wire6306 = ( n_n854  &  (~ n_n856)  &  wire6305 ) ;
 assign wire6309 = ( (~ n_n858)  &  (~ n_n857) ) ;
 assign wire6310 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6312 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire6313 = ( wire578  &  wire6312 ) | ( wire579  &  wire6312 ) ;
 assign wire6315 = ( (~ s298_in_2_)  &  s298_out_3_  &  n_n51 ) ;
 assign wire6318 = ( wire6126  &  wire6127 ) | ( wire6132  &  wire6133 ) ;
 assign wire6319 = ( wire6138  &  wire6139 ) | ( wire6144  &  wire6145 ) ;
 assign wire6320 = ( wire6269  &  wire6270 ) | ( wire6309  &  wire6310 ) ;
 assign wire6323 = ( (~ s298_out_5_)  &  wire6245 ) | ( (~ s298_out_5_)  &  wire6095  &  wire6096 ) ;
 assign wire6324 = ( (~ s298_out_5_)  &  wire6306 ) | ( (~ s298_out_5_)  &  wire6248  &  wire6249 ) ;
 assign wire6325 = ( wire446 ) | ( wire6318 ) | ( wire6319 ) | ( wire6320 ) ;
 assign wire6328 = ( wire621  &  wire6091 ) | ( wire622  &  wire6091 ) | ( wire621  &  wire6235 ) | ( wire622  &  wire6235 ) ;
 assign wire6329 = ( wire464 ) | ( wire6323 ) | ( wire6324 ) ;
 assign wire6330 = ( wire471 ) | ( wire470 ) ;
 assign wire6331 = ( wire501 ) | ( wire495 ) ;
 assign wire6332 = ( wire458 ) | ( wire6325 ) | ( wire6328 ) ;
 assign wire6333 = ( n_n51  &  wire6150 ) | ( n_n51  &  wire6101  &  wire6102 ) ;
 assign wire6334 = ( (~ n_n51)  &  wire6255 ) | ( (~ s298_out_5_)  &  n_n51  &  wire6239 ) ;
 assign wire6335 = ( n_n51  &  wire6265 ) | ( (~ n_n51)  &  wire6258  &  wire6259 ) ;
 assign wire6338 = ( s298_out_0_  &  wire6073 ) | ( s298_out_0_  &  (~ n_n51)  &  wire6204 ) ;
 assign wire6339 = ( wire578  &  wire6210 ) | ( wire579  &  wire6210 ) | ( wire578  &  wire6215 ) | ( wire579  &  wire6215 ) ;
 assign wire6342 = ( wire6329 ) | ( wire6330 ) | ( wire6331 ) | ( wire6332 ) ;
 assign wire6344 = ( wire506 ) | ( wire6333 ) | ( wire6334 ) | ( wire6335 ) ;
 assign wire6345 = ( wire6338 ) | ( wire6339 ) | ( wire6342 ) ;
 assign wire6351 = ( wire447 ) | ( wire485 ) | ( wire6344 ) | ( wire6345 ) ;
 assign wire6352 = ( wire457 ) | ( wire462 ) | ( wire463 ) | ( wire479 ) ;
 assign wire6354 = ( wire483 ) | ( wire484 ) | ( wire6351 ) | ( wire6352 ) ;
 assign wire6367 = ( wire448 ) | ( wire449 ) | ( wire450 ) | ( wire6354 ) ;
 assign wire6368 = ( wire451 ) | ( wire452 ) | ( wire453 ) | ( wire454 ) ;
 assign wire6369 = ( wire455 ) | ( wire472 ) | ( wire473 ) | ( wire474 ) ;
 assign wire6370 = ( wire475 ) | ( wire476 ) | ( wire477 ) | ( wire478 ) ;
 assign wire6371 = ( wire494 ) | ( wire496 ) | ( wire497 ) | ( wire498 ) ;
 assign wire6372 = ( wire499 ) | ( wire500 ) | ( wire504 ) | ( wire505 ) ;
 assign wire6375 = ( wire6372 ) | ( wire6371 ) ;
 assign wire6376 = ( wire6367 ) | ( wire6368 ) | ( wire6369 ) | ( wire6370 ) ;
 assign wire6381 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6382 = ( n_n853  &  (~ n_n854)  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire6384 = ( (~ wire621)  &  (~ wire622)  &  wire6381  &  wire6382 ) ;
 assign wire6389 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6390 = ( (~ n_n853)  &  n_n855  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire6392 = ( (~ wire578)  &  (~ wire579)  &  wire6389  &  wire6390 ) ;
 assign wire6397 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6398 = ( (~ n_n853)  &  (~ n_n855)  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire6399 = ( wire6398  &  wire6397 ) ;
 assign wire6404 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6406 = ( (~ s298_out_5_)  &  (~ n_n853)  &  (~ n_n859)  &  wire6404 ) ;
 assign wire6407 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6406 ) ;
 assign wire6410 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n853) ) ;
 assign wire6412 = ( (~ s298_in_1_)  &  s298_out_5_  &  (~ n_n852)  &  wire6410 ) ;
 assign wire6413 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6412 ) ;
 assign wire6414 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6413 ) ;
 assign wire6418 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire6419 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6421 = ( (~ wire578)  &  (~ wire579)  &  wire6418  &  wire6419 ) ;
 assign wire6425 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6426 = ( (~ n_n853)  &  (~ n_n855)  &  wire6425 ) ;
 assign wire6428 = ( (~ s298_out_5_)  &  (~ n_n859)  &  (~ wire5513)  &  wire6426 ) ;
 assign wire6431 = ( (~ n_n856)  &  n_n853 ) ;
 assign wire6432 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6434 = ( wire621  &  wire6431  &  wire6432 ) | ( wire622  &  wire6431  &  wire6432 ) ;
 assign wire6435 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6434 ) ;
 assign wire6440 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6441 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire6440 ) ;
 assign wire6442 = ( wire5789  &  wire6441 ) | ( wire5790  &  wire6441 ) | ( wire5791  &  wire6441 ) ;
 assign wire6447 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  (~ n_n856) ) ;
 assign wire6448 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire6447 ) ;
 assign wire6449 = ( wire5789  &  wire6448 ) | ( wire5790  &  wire6448 ) | ( wire5791  &  wire6448 ) ;
 assign wire6454 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire6455 = ( (~ n_n854)  &  n_n855  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire6456 = ( wire6455  &  wire6454 ) ;
 assign wire6461 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6462 = ( n_n853  &  n_n854  &  n_n856  &  (~ n_n857) ) ;
 assign wire6463 = ( wire6462  &  wire6461 ) ;
 assign wire6467 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire6468 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire6470 = ( (~ wire578)  &  (~ wire579)  &  wire6467  &  wire6468 ) ;
 assign wire6473 = ( (~ n_n855)  &  n_n854 ) ;
 assign wire6474 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n853) ) ;
 assign wire6476 = ( wire578  &  wire6473  &  wire6474 ) | ( wire579  &  wire6473  &  wire6474 ) ;
 assign wire6477 = ( wire5789  &  wire6476 ) | ( wire5790  &  wire6476 ) | ( wire5791  &  wire6476 ) ;
 assign wire6481 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855) ) ;
 assign wire6482 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6484 = ( wire621  &  wire6481  &  wire6482 ) | ( wire622  &  wire6481  &  wire6482 ) ;
 assign wire6488 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire6489 = ( (~ s298_in_1_)  &  (~ n_n853)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6491 = ( (~ s298_out_3_)  &  wire6488  &  wire6489 ) ;
 assign wire6496 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6497 = ( n_n853  &  (~ n_n855)  &  (~ n_n856)  &  n_n859 ) ;
 assign wire6498 = ( wire6497  &  wire6496 ) ;
 assign wire6503 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6504 = ( (~ n_n853)  &  n_n854  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire6505 = ( wire6504  &  wire6503 ) ;
 assign wire6510 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6511 = ( n_n853  &  n_n854  &  (~ n_n857)  &  n_n859 ) ;
 assign wire6512 = ( wire6511  &  wire6510 ) ;
 assign wire6517 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6518 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855)  &  wire6517 ) ;
 assign wire6523 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855) ) ;
 assign wire6524 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6526 = ( wire578  &  wire6523  &  wire6524 ) | ( wire579  &  wire6523  &  wire6524 ) ;
 assign wire6531 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6532 = ( (~ n_n853)  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire6533 = ( wire6532  &  wire6531 ) ;
 assign wire6537 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire6538 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  (~ n_n854) ) ;
 assign wire6540 = ( (~ wire621)  &  (~ wire622)  &  wire6537  &  wire6538 ) ;
 assign wire6545 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire6546 = ( (~ n_n854)  &  (~ n_n855)  &  n_n858  &  (~ n_n859) ) ;
 assign wire6552 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6553 = ( (~ n_n853)  &  (~ n_n855)  &  n_n857  &  (~ n_n859) ) ;
 assign wire6554 = ( wire6553  &  wire6552 ) ;
 assign wire6559 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6560 = ( n_n853  &  n_n854  &  (~ n_n855)  &  n_n858 ) ;
 assign wire6561 = ( wire6560  &  wire6559 ) ;
 assign wire6566 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire6567 = ( n_n854  &  (~ n_n855)  &  (~ n_n856)  &  n_n858 ) ;
 assign wire6568 = ( wire6567  &  wire6566 ) ;
 assign wire6572 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire6573 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n855) ) ;
 assign wire6575 = ( wire621  &  wire6572  &  wire6573 ) | ( wire622  &  wire6572  &  wire6573 ) ;
 assign wire6580 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6581 = ( (~ n_n853)  &  (~ n_n854)  &  n_n855  &  (~ n_n857) ) ;
 assign wire6582 = ( wire6581  &  wire6580 ) ;
 assign wire6586 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856 ) ;
 assign wire6587 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire6589 = ( (~ s298_out_5_)  &  wire6586  &  wire6587 ) ;
 assign wire6594 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6595 = ( (~ n_n853)  &  n_n854  &  n_n855  &  (~ n_n858) ) ;
 assign wire6600 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire6601 = ( s298_in_1_  &  (~ n_n852)  &  n_n855  &  n_n856 ) ;
 assign wire6603 = ( (~ n_n51)  &  wire6600  &  wire6601 ) ;
 assign wire6608 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n856) ) ;
 assign wire6609 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire6608 ) ;
 assign wire6610 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire6609 ) ;
 assign wire6615 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6616 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire6622 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6623 = ( (~ n_n853)  &  n_n854  &  (~ n_n856)  &  n_n857 ) ;
 assign wire6629 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6630 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire6631 = ( wire6630  &  wire6629 ) ;
 assign wire6636 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6637 = ( n_n853  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire6638 = ( wire6637  &  wire6636 ) ;
 assign wire6643 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire6644 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n855 ) ;
 assign wire6650 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire6651 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6657 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire6658 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  (~ n_n855) ) ;
 assign wire6664 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire6665 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6671 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire6672 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6678 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire6679 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6685 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire6686 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire6692 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire6693 = ( s298_in_1_  &  n_n852  &  n_n854  &  (~ n_n855) ) ;
 assign wire6699 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire6700 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  n_n855 ) ;
 assign wire6705 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6706 = ( n_n853  &  (~ n_n859)  &  wire6705 ) ;
 assign wire6707 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire6706 ) ;
 assign wire6711 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6712 = ( (~ n_n855)  &  (~ n_n856)  &  wire6711 ) ;
 assign wire6713 = ( wire580  &  wire6712 ) | ( wire581  &  wire6712 ) | ( wire582  &  wire6712 ) ;
 assign wire6715 = ( (~ n_n852)  &  (~ s298_in_1_) ) ;
 assign wire6716 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n854) ) ;
 assign wire6718 = ( wire578  &  wire6715  &  wire6716 ) | ( wire579  &  wire6715  &  wire6716 ) ;
 assign wire6719 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6718 ) ;
 assign wire6721 = ( (~ n_n852)  &  s298_in_1_ ) ;
 assign wire6722 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n853 ) ;
 assign wire6724 = ( wire621  &  wire6721  &  wire6722 ) | ( wire622  &  wire6721  &  wire6722 ) ;
 assign wire6725 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6724 ) ;
 assign wire6728 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire6729 = ( (~ s298_in_1_)  &  n_n852  &  wire6728 ) ;
 assign wire6731 = ( (~ n_n51)  &  (~ wire621)  &  (~ wire622)  &  wire6729 ) ;
 assign wire6733 = ( n_n854  &  s298_in_1_ ) ;
 assign wire6734 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire6736 = ( (~ wire621)  &  (~ wire622)  &  wire6733  &  wire6734 ) ;
 assign wire6737 = ( wire5789  &  wire6736 ) | ( wire5790  &  wire6736 ) | ( wire5791  &  wire6736 ) ;
 assign wire6740 = ( n_n856  &  n_n854 ) ;
 assign wire6741 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire6743 = ( wire621  &  wire6740  &  wire6741 ) | ( wire622  &  wire6740  &  wire6741 ) ;
 assign wire6747 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6748 = ( n_n853  &  (~ n_n857)  &  wire6747 ) ;
 assign wire6749 = ( wire5789  &  wire6748 ) | ( wire5790  &  wire6748 ) | ( wire5791  &  wire6748 ) ;
 assign wire6754 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n854)  &  n_n856 ) ;
 assign wire6755 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858)  &  wire6754 ) ;
 assign wire6760 = ( s298_in_1_  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire6761 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire6760 ) ;
 assign wire6763 = ( (~ n_n855)  &  n_n853 ) ;
 assign wire6764 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n856 ) ;
 assign wire6767 = ( s298_out_5_  &  (~ n_n51)  &  wire6763  &  wire6764 ) ;
 assign wire6770 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n855 ) ;
 assign wire6772 = ( n_n853  &  (~ n_n854)  &  n_n51  &  wire6770 ) ;
 assign wire6773 = ( wire5789  &  wire6772 ) | ( wire5790  &  wire6772 ) | ( wire5791  &  wire6772 ) ;
 assign wire6778 = ( (~ n_n853)  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire6779 = ( s298_in_1_  &  n_n852  &  (~ n_n857)  &  wire6778 ) ;
 assign wire6783 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6784 = ( (~ n_n855)  &  n_n856  &  wire6783 ) ;
 assign wire6785 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire6784 ) ;
 assign wire6787 = ( n_n854  &  (~ n_n852) ) ;
 assign wire6788 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n855) ) ;
 assign wire6790 = ( wire578  &  wire6787  &  wire6788 ) | ( wire579  &  wire6787  &  wire6788 ) ;
 assign wire6791 = ( wire5789  &  wire6790 ) | ( wire5790  &  wire6790 ) | ( wire5791  &  wire6790 ) ;
 assign wire6794 = ( n_n856  &  (~ n_n855) ) ;
 assign wire6795 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire6797 = ( wire578  &  wire6794  &  wire6795 ) | ( wire579  &  wire6794  &  wire6795 ) ;
 assign wire6800 = ( n_n856  &  (~ n_n855) ) ;
 assign wire6801 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n854) ) ;
 assign wire6803 = ( wire621  &  wire6800  &  wire6801 ) | ( wire622  &  wire6800  &  wire6801 ) ;
 assign wire6807 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n853  &  (~ n_n854) ) ;
 assign wire6808 = ( n_n855  &  (~ n_n856)  &  wire6807 ) ;
 assign wire6809 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire6808 ) ;
 assign wire6814 = ( n_n852  &  n_n854  &  n_n855  &  (~ n_n857) ) ;
 assign wire6815 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n859  &  wire6814 ) ;
 assign wire6820 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  (~ n_n855) ) ;
 assign wire6821 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856  &  wire6820 ) ;
 assign wire6826 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n855)  &  n_n857 ) ;
 assign wire6827 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858)  &  wire6826 ) ;
 assign wire6830 = ( n_n855  &  (~ n_n854) ) ;
 assign wire6831 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire6833 = ( wire621  &  wire6830  &  wire6831 ) | ( wire622  &  wire6830  &  wire6831 ) ;
 assign wire6838 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n854)  &  n_n855 ) ;
 assign wire6839 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856  &  wire6838 ) ;
 assign wire6844 = ( s298_in_1_  &  (~ n_n852)  &  n_n854  &  n_n855 ) ;
 assign wire6845 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire6844 ) ;
 assign wire6850 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire6851 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n855)  &  wire6850 ) ;
 assign wire6856 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n856 ) ;
 assign wire6857 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire6856 ) ;
 assign wire6862 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n854)  &  n_n856 ) ;
 assign wire6863 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire6862 ) ;
 assign wire6867 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire6869 = ( n_n855  &  n_n857  &  n_n51  &  wire6867 ) ;
 assign wire6874 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n855 ) ;
 assign wire6875 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856  &  wire6874 ) ;
 assign wire6880 = ( n_n852  &  (~ n_n853)  &  n_n855  &  n_n856 ) ;
 assign wire6881 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n857)  &  wire6880 ) ;
 assign wire6885 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n853 ) ;
 assign wire6886 = ( n_n854  &  (~ n_n859)  &  wire6885 ) ;
 assign wire6887 = ( wire619  &  wire6886 ) | ( wire621  &  wire6886 ) | ( wire622  &  wire6886 ) ;
 assign wire6892 = ( (~ s298_in_1_)  &  n_n854  &  n_n855  &  n_n856 ) ;
 assign wire6893 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire6892 ) ;
 assign wire6898 = ( s298_in_1_  &  n_n852  &  (~ n_n854)  &  (~ n_n856) ) ;
 assign wire6899 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857  &  wire6898 ) ;
 assign wire6904 = ( s298_in_1_  &  n_n854  &  n_n855  &  (~ n_n856) ) ;
 assign wire6905 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire6904 ) ;
 assign wire6910 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire6911 = ( n_n853  &  (~ n_n854)  &  n_n856  &  (~ n_n859) ) ;
 assign wire6916 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6917 = ( (~ n_n853)  &  n_n854  &  n_n856  &  (~ n_n859) ) ;
 assign wire6922 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire6923 = ( n_n853  &  n_n856  &  n_n858  &  (~ n_n859) ) ;
 assign wire6928 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6929 = ( (~ n_n855)  &  n_n856  &  n_n858  &  (~ n_n859) ) ;
 assign wire6934 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n853) ) ;
 assign wire6935 = ( (~ n_n854)  &  (~ n_n856)  &  n_n857  &  n_n859 ) ;
 assign wire6940 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire6941 = ( n_n853  &  (~ n_n854)  &  (~ n_n856)  &  n_n857 ) ;
 assign wire6946 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6947 = ( (~ n_n853)  &  n_n856  &  n_n857  &  (~ n_n858) ) ;
 assign wire6952 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire6953 = ( n_n853  &  (~ n_n855)  &  n_n857  &  n_n858 ) ;
 assign wire6958 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire6959 = ( (~ n_n855)  &  n_n856  &  n_n857  &  (~ n_n858) ) ;
 assign wire6962 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n855)  &  n_n856 ) ;
 assign wire6963 = ( wire621  &  wire6962 ) | ( wire622  &  wire6962 ) ;
 assign wire6964 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire6963 ) ;
 assign wire6967 = ( (~ s298_in_1_)  &  n_n854  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire6968 = ( wire623  &  wire6967 ) | ( wire624  &  wire6967 ) | ( wire625  &  wire6967 ) ;
 assign wire6969 = ( wire6016  &  wire6968 ) | ( wire6017  &  wire6968 ) | ( wire6018  &  wire6968 ) ;
 assign wire6973 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  (~ n_n854) ) ;
 assign wire6974 = ( n_n856  &  (~ n_n858)  &  wire6973 ) ;
 assign wire6977 = ( s298_in_1_  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire6978 = ( wire578  &  wire6977 ) | ( wire579  &  wire6977 ) ;
 assign wire6979 = ( wire6016  &  wire6978 ) | ( wire6017  &  wire6978 ) | ( wire6018  &  wire6978 ) ;
 assign wire6982 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n856) ) ;
 assign wire6984 = ( (~ s298_out_5_)  &  n_n854  &  (~ n_n855)  &  wire6982 ) ;
 assign wire6987 = ( s298_in_0_  &  s298_in_1_  &  n_n855 ) ;
 assign wire6989 = ( (~ s298_out_5_)  &  n_n852  &  n_n853  &  wire6987 ) ;
 assign wire6992 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n857) ) ;
 assign wire6994 = ( s298_out_5_  &  (~ n_n854)  &  (~ n_n856)  &  wire6992 ) ;
 assign wire6997 = ( s298_in_1_  &  (~ n_n852)  &  n_n856 ) ;
 assign wire6998 = ( (~ n_n853)  &  n_n854  &  wire6997 ) ;
 assign wire6999 = ( wire5789  &  wire6998 ) | ( wire5790  &  wire6998 ) | ( wire5791  &  wire6998 ) ;
 assign wire7003 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire7004 = ( (~ n_n855)  &  n_n859  &  wire7003 ) ;
 assign wire7008 = ( s298_in_0_  &  s298_in_1_  &  n_n853  &  n_n854 ) ;
 assign wire7009 = ( n_n855  &  (~ n_n856)  &  wire7008 ) ;
 assign wire7013 = ( (~ s298_in_1_)  &  n_n852  &  n_n855  &  n_n856 ) ;
 assign wire7014 = ( n_n857  &  (~ n_n858)  &  wire7013 ) ;
 assign wire7017 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire7018 = ( s298_in_1_  &  (~ n_n853)  &  wire7017 ) ;
 assign wire7019 = ( wire580  &  wire7018 ) | ( wire581  &  wire7018 ) | ( wire582  &  wire7018 ) ;
 assign wire7022 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7023 = ( wire580  &  wire7022 ) | ( wire581  &  wire7022 ) | ( wire582  &  wire7022 ) ;
 assign wire7024 = ( wire7023  &  (~ n_n51) ) ;
 assign wire7028 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire7029 = ( n_n855  &  n_n856  &  wire7028 ) ;
 assign wire7033 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  n_n853 ) ;
 assign wire7034 = ( n_n855  &  n_n856  &  wire7033 ) ;
 assign wire7037 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n859) ) ;
 assign wire7038 = ( (~ n_n853)  &  n_n856  &  wire7037 ) ;
 assign wire7039 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7038 ) ;
 assign wire7042 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire7044 = ( s298_in_1_  &  s298_out_3_  &  (~ n_n852)  &  wire7042 ) ;
 assign wire7047 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n855) ) ;
 assign wire7049 = ( n_n852  &  n_n853  &  (~ n_n51)  &  wire7047 ) ;
 assign wire7052 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n857) ) ;
 assign wire7054 = ( (~ n_n852)  &  n_n854  &  n_n51  &  wire7052 ) ;
 assign wire7056 = ( n_n853  &  (~ s298_in_1_) ) ;
 assign wire7057 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire7059 = ( wire621  &  wire7056  &  wire7057 ) | ( wire622  &  wire7056  &  wire7057 ) ;
 assign wire7063 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire7064 = ( (~ n_n855)  &  n_n857  &  wire7063 ) ;
 assign wire7068 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire7069 = ( n_n855  &  (~ n_n856)  &  wire7068 ) ;
 assign wire7072 = ( n_n857  &  n_n855 ) ;
 assign wire7073 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire7078 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n855) ) ;
 assign wire7079 = ( n_n856  &  n_n857  &  wire7078 ) ;
 assign wire7083 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire7084 = ( s298_in_1_  &  n_n855  &  n_n857  &  (~ n_n858) ) ;
 assign wire7086 = ( (~ s298_in_1_)  &  n_n855  &  (~ n_n856) ) ;
 assign wire7087 = ( wire621  &  wire7086 ) | ( wire622  &  wire7086 ) ;
 assign wire7088 = ( wire6016  &  wire7087 ) | ( wire6017  &  wire7087 ) | ( wire6018  &  wire7087 ) ;
 assign wire7091 = ( s298_in_1_  &  (~ n_n853)  &  n_n857  &  n_n858 ) ;
 assign wire7092 = ( wire578  &  wire7091 ) | ( wire579  &  wire7091 ) ;
 assign wire7095 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n852  &  n_n856 ) ;
 assign wire7096 = ( wire621  &  wire7095 ) | ( wire622  &  wire7095 ) ;
 assign wire7099 = ( (~ s298_in_1_)  &  n_n852  &  n_n858 ) ;
 assign wire7100 = ( (~ n_n853)  &  (~ n_n856)  &  wire7099 ) ;
 assign wire7103 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n855) ) ;
 assign wire7104 = ( s298_in_1_  &  n_n854  &  wire7103 ) ;
 assign wire7106 = ( (~ s298_in_1_)  &  n_n853  &  n_n859 ) ;
 assign wire7108 = ( n_n51  &  wire621  &  wire7106 ) | ( n_n51  &  wire622  &  wire7106 ) ;
 assign wire7110 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7111 = ( wire619  &  wire7110 ) | ( wire621  &  wire7110 ) | ( wire622  &  wire7110 ) ;
 assign wire7112 = ( wire7111  &  n_n51 ) ;
 assign wire7114 = ( (~ s298_in_1_)  &  n_n852  &  n_n858 ) ;
 assign wire7115 = ( wire578  &  wire7114 ) | ( wire579  &  wire7114 ) ;
 assign wire7116 = ( wire6910  &  wire6911 ) | ( wire6916  &  wire6917 ) ;
 assign wire7117 = ( wire6922  &  wire6923 ) | ( wire6928  &  wire6929 ) ;
 assign wire7118 = ( wire6934  &  wire6935 ) | ( wire6940  &  wire6941 ) ;
 assign wire7119 = ( wire6946  &  wire6947 ) | ( wire6952  &  wire6953 ) ;
 assign wire7120 = ( wire6958  &  wire6959 ) | ( wire7083  &  wire7084 ) ;
 assign wire7127 = ( wire7120 ) | ( wire7119 ) ;
 assign wire7128 = ( (~ s298_out_5_)  &  wire6863 ) | ( (~ s298_out_5_)  &  wire6594  &  wire6595 ) ;
 assign wire7129 = ( wire361 ) | ( wire362 ) | ( wire363 ) | ( wire364 ) ;
 assign wire7130 = ( wire365 ) | ( wire366 ) | ( wire367 ) | ( wire368 ) ;
 assign wire7131 = ( wire369 ) | ( wire7116 ) | ( wire7117 ) | ( wire7118 ) ;
 assign wire7135 = ( (~ wire621)  &  (~ wire622)  &  wire6554 ) | ( (~ wire621)  &  (~ wire622)  &  wire6561 ) ;
 assign wire7136 = ( wire621  &  wire6582 ) | ( wire622  &  wire6582 ) | ( (~ wire621)  &  (~ wire622)  &  wire6568 ) ;
 assign wire7137 = ( wire621  &  wire6839 ) | ( wire622  &  wire6839 ) | ( wire621  &  wire6845 ) | ( wire622  &  wire6845 ) ;
 assign wire7138 = ( wire621  &  wire6851 ) | ( wire622  &  wire6851 ) | ( wire621  &  wire6857 ) | ( wire622  &  wire6857 ) ;
 assign wire7139 = ( wire621  &  wire7064 ) | ( wire622  &  wire7064 ) | ( wire621  &  wire7069 ) | ( wire622  &  wire7069 ) ;
 assign wire7140 = ( wire7127 ) | ( wire7128 ) | ( wire7129 ) | ( wire7130 ) ;
 assign wire7141 = ( wire335 ) | ( wire334 ) ;
 assign wire7145 = ( wire347 ) | ( wire7131 ) | ( wire7135 ) ;
 assign wire7148 = ( wire7140 ) | ( (~ s298_out_5_)  &  n_n51  &  wire6399 ) ;
 assign wire7149 = ( n_n51  &  wire6610 ) | ( n_n51  &  wire6615  &  wire6616 ) ;
 assign wire7150 = ( n_n51  &  wire6785 ) | ( n_n51  &  wire6622  &  wire6623 ) ;
 assign wire7151 = ( wire7141 ) | ( n_n51  &  wire7072  &  wire7073 ) ;
 assign wire7152 = ( wire360 ) | ( wire402 ) | ( wire403 ) | ( wire426 ) ;
 assign wire7154 = ( wire7136 ) | ( wire7137 ) | ( wire7138 ) | ( wire7139 ) ;
 assign wire7155 = ( s298_out_0_  &  wire6533 ) | ( s298_out_0_  &  (~ n_n51)  &  wire6518 ) ;
 assign wire7156 = ( wire578  &  wire6827 ) | ( wire579  &  wire6827 ) | ( (~ wire578)  &  (~ wire579)  &  wire6821 ) ;
 assign wire7159 = ( wire427 ) | ( wire442 ) | ( wire7145 ) | ( wire7152 ) ;
 assign wire7161 = ( wire7148 ) | ( wire7149 ) | ( wire7156 ) ;
 assign wire7162 = ( wire7150 ) | ( wire7151 ) | ( wire7159 ) ;
 assign wire7164 = ( wire7154 ) | ( wire7155 ) | ( wire7161 ) | ( wire7162 ) ;
 assign wire7173 = ( wire344 ) | ( wire444 ) | ( wire7164 ) ;
 assign wire7174 = ( wire346 ) | ( wire351 ) | ( wire353 ) | ( wire355 ) ;
 assign wire7175 = ( wire359 ) | ( wire391 ) | ( wire397 ) | ( wire398 ) ;
 assign wire7176 = ( wire399 ) | ( wire400 ) | ( wire401 ) | ( wire425 ) ;
 assign wire7178 = ( wire7175 ) | ( wire7174 ) ;
 assign wire7179 = ( wire432 ) | ( wire436 ) | ( wire7173 ) | ( wire7176 ) ;
 assign wire7190 = ( wire445 ) | ( wire443 ) ;
 assign wire7191 = ( wire325 ) | ( wire336 ) | ( wire7178 ) | ( wire7179 ) ;
 assign wire7192 = ( wire337 ) | ( wire338 ) | ( wire339 ) | ( wire340 ) ;
 assign wire7193 = ( wire341 ) | ( wire342 ) | ( wire384 ) | ( wire385 ) ;
 assign wire7194 = ( wire386 ) | ( wire387 ) | ( wire388 ) | ( wire424 ) ;
 assign wire7195 = ( wire428 ) | ( wire429 ) | ( wire430 ) | ( wire431 ) ;
 assign wire7199 = ( wire7190 ) | ( wire7191 ) | ( wire7192 ) | ( wire7193 ) ;
 assign wire7200 = ( wire7194 ) | ( wire7195 ) | ( wire7199 ) ;
 assign wire7202 = ( (~ wire6375)  &  (~ wire6376)  &  wire6407 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6414 ) ;
 assign wire7203 = ( (~ wire6375)  &  (~ wire6376)  &  wire6421 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6428 ) ;
 assign wire7204 = ( (~ wire6375)  &  (~ wire6376)  &  wire6435 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6442 ) ;
 assign wire7205 = ( (~ wire6375)  &  (~ wire6376)  &  wire6449 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6707 ) ;
 assign wire7206 = ( (~ wire6375)  &  (~ wire6376)  &  wire6713 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6719 ) ;
 assign wire7207 = ( (~ wire6375)  &  (~ wire6376)  &  wire6725 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6731 ) ;
 assign wire7208 = ( (~ wire6375)  &  (~ wire6376)  &  wire6737 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6743 ) ;
 assign wire7209 = ( (~ wire6375)  &  (~ wire6376)  &  wire6749 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6755 ) ;
 assign wire7210 = ( wire6375  &  wire6767 ) | ( wire6376  &  wire6767 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6761 ) ;
 assign wire7211 = ( wire6375  &  wire6773 ) | ( wire6376  &  wire6773 ) | ( wire6375  &  wire6779 ) | ( wire6376  &  wire6779 ) ;
 assign wire7212 = ( (~ wire6375)  &  (~ wire6376)  &  wire6964 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6969 ) ;
 assign wire7213 = ( wire6375  &  wire6979 ) | ( wire6376  &  wire6979 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire6974 ) ;
 assign wire7214 = ( wire6375  &  wire6984 ) | ( wire6376  &  wire6984 ) | ( wire6375  &  wire6989 ) | ( wire6376  &  wire6989 ) ;
 assign wire7215 = ( wire6375  &  wire6994 ) | ( wire6376  &  wire6994 ) | ( wire6375  &  wire6999 ) | ( wire6376  &  wire6999 ) ;
 assign wire7216 = ( wire6375  &  wire7004 ) | ( wire6376  &  wire7004 ) | ( wire6375  &  wire7009 ) | ( wire6376  &  wire7009 ) ;
 assign wire7217 = ( wire6375  &  wire7014 ) | ( wire6376  &  wire7014 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7088 ) ;
 assign wire7218 = ( wire6375  &  wire7092 ) | ( wire6376  &  wire7092 ) | ( wire6375  &  wire7096 ) | ( wire6376  &  wire7096 ) ;
 assign wire7228 = ( wire324 ) | ( wire441 ) | ( wire7200 ) | ( wire7218 ) ;
 assign wire7229 = ( wire7202 ) | ( wire7203 ) | ( wire7204 ) | ( wire7205 ) ;
 assign wire7230 = ( wire7206 ) | ( wire7207 ) | ( wire7208 ) | ( wire7209 ) ;
 assign wire7231 = ( wire7210 ) | ( wire7211 ) | ( wire7212 ) | ( wire7213 ) ;
 assign wire7232 = ( wire7214 ) | ( wire7215 ) | ( wire7216 ) | ( wire7217 ) ;
 assign wire7235 = ( wire7228 ) | ( wire7229 ) | ( wire7232 ) ;
 assign wire7240 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire7241 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire7243 = ( (~ n_n855)  &  (~ n_n857)  &  wire7240  &  wire7241 ) ;
 assign wire7245 = ( (~ n_n854)  &  (~ n_n853) ) ;
 assign wire7246 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire7249 = ( (~ s298_out_3_)  &  n_n51  &  wire7245  &  wire7246 ) ;
 assign wire7250 = ( wire6016  &  wire7249 ) | ( wire6017  &  wire7249 ) | ( wire6018  &  wire7249 ) ;
 assign wire7254 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire7255 = ( s298_in_1_  &  n_n852  &  n_n855  &  n_n857 ) ;
 assign wire7257 = ( wire621  &  wire7254  &  wire7255 ) | ( wire622  &  wire7254  &  wire7255 ) ;
 assign wire7261 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire7263 = ( n_n855  &  (~ n_n856)  &  (~ n_n51)  &  wire7261 ) ;
 assign wire7264 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7263 ) ;
 assign wire7268 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n858) ) ;
 assign wire7269 = ( n_n852  &  n_n853  &  n_n854  &  n_n857 ) ;
 assign wire7271 = ( n_n51  &  wire7268  &  wire7269 ) ;
 assign wire7276 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7277 = ( (~ n_n853)  &  (~ n_n854)  &  n_n856  &  n_n858 ) ;
 assign wire7278 = ( wire7277  &  wire7276 ) ;
 assign wire7282 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire7283 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  (~ n_n854) ) ;
 assign wire7285 = ( n_n51  &  wire7282  &  wire7283 ) ;
 assign wire7290 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire7291 = ( n_n853  &  (~ n_n854)  &  n_n855  &  (~ n_n856) ) ;
 assign wire7292 = ( wire7291  &  wire7290 ) ;
 assign wire7297 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7298 = ( n_n853  &  n_n854  &  n_n855  &  n_n857 ) ;
 assign wire7299 = ( wire7298  &  wire7297 ) ;
 assign wire7304 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7305 = ( n_n854  &  (~ n_n855)  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire7311 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7312 = ( n_n853  &  n_n854  &  (~ n_n855)  &  (~ n_n858) ) ;
 assign wire7313 = ( wire7312  &  wire7311 ) ;
 assign wire7318 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7319 = ( n_n853  &  n_n854  &  n_n855  &  (~ n_n857) ) ;
 assign wire7320 = ( wire7319  &  wire7318 ) ;
 assign wire7325 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7326 = ( (~ n_n853)  &  (~ n_n855)  &  n_n857  &  (~ n_n858) ) ;
 assign wire7327 = ( wire7326  &  wire7325 ) ;
 assign wire7332 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7333 = ( n_n853  &  n_n854  &  (~ n_n855)  &  n_n857 ) ;
 assign wire7334 = ( wire7333  &  wire7332 ) ;
 assign wire7339 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7340 = ( n_n853  &  (~ n_n855)  &  n_n856  &  (~ n_n857) ) ;
 assign wire7341 = ( wire7340  &  wire7339 ) ;
 assign wire7345 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire7346 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n854)  &  n_n855 ) ;
 assign wire7348 = ( wire621  &  wire7345  &  wire7346 ) | ( wire622  &  wire7345  &  wire7346 ) ;
 assign wire7353 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7354 = ( n_n853  &  n_n854  &  n_n855  &  (~ n_n856) ) ;
 assign wire7355 = ( wire7354  &  wire7353 ) ;
 assign wire7360 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire7361 = ( n_n854  &  (~ n_n855)  &  n_n858  &  n_n859 ) ;
 assign wire7362 = ( wire7361  &  wire7360 ) ;
 assign wire7367 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7368 = ( (~ n_n853)  &  (~ n_n855)  &  (~ n_n856)  &  n_n859 ) ;
 assign wire7369 = ( wire7368  &  wire7367 ) ;
 assign wire7374 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7375 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire7376 = ( wire7375  &  wire7374 ) ;
 assign wire7381 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire7382 = ( (~ n_n854)  &  n_n855  &  n_n856  &  (~ n_n857) ) ;
 assign wire7383 = ( wire7382  &  wire7381 ) ;
 assign wire7388 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7389 = ( n_n853  &  (~ n_n854)  &  (~ n_n856)  &  n_n858 ) ;
 assign wire7395 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire7396 = ( s298_in_1_  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire7402 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire7403 = ( (~ s298_in_1_)  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire7409 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire7410 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire7416 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire7417 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire7421 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n855 ) ;
 assign wire7422 = ( (~ n_n852)  &  (~ n_n853)  &  wire7421 ) ;
 assign wire7423 = ( wire580  &  wire7422 ) | ( wire581  &  wire7422 ) | ( wire582  &  wire7422 ) ;
 assign wire7424 = ( wire7423  &  n_n51 ) ;
 assign wire7428 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire7429 = ( n_n856  &  (~ n_n859)  &  wire7428 ) ;
 assign wire7430 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7429 ) ;
 assign wire7433 = ( (~ n_n856)  &  (~ n_n853) ) ;
 assign wire7434 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7436 = ( wire578  &  wire7433  &  wire7434 ) | ( wire579  &  wire7433  &  wire7434 ) ;
 assign wire7440 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n854) ) ;
 assign wire7442 = ( n_n855  &  (~ n_n857)  &  (~ n_n51)  &  wire7440 ) ;
 assign wire7446 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire7448 = ( (~ n_n856)  &  (~ n_n857)  &  n_n51  &  wire7446 ) ;
 assign wire7453 = ( n_n853  &  (~ n_n854)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire7454 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n859)  &  wire7453 ) ;
 assign wire7459 = ( n_n853  &  n_n854  &  (~ n_n855)  &  n_n858 ) ;
 assign wire7460 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n859  &  wire7459 ) ;
 assign wire7465 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire7466 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858)  &  wire7465 ) ;
 assign wire7471 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n854)  &  n_n855 ) ;
 assign wire7472 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856  &  wire7471 ) ;
 assign wire7477 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n856 ) ;
 assign wire7478 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858  &  wire7477 ) ;
 assign wire7481 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n855 ) ;
 assign wire7482 = ( (~ n_n852)  &  n_n853  &  wire7481 ) ;
 assign wire7483 = ( wire5789  &  wire7482 ) | ( wire5790  &  wire7482 ) | ( wire5791  &  wire7482 ) ;
 assign wire7484 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7483 ) ;
 assign wire7489 = ( (~ n_n853)  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire7490 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n857  &  wire7489 ) ;
 assign wire7494 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7495 = ( n_n853  &  (~ n_n854)  &  wire7494 ) ;
 assign wire7501 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  n_n855 ) ;
 assign wire7502 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire7501 ) ;
 assign wire7505 = ( n_n856  &  n_n855 ) ;
 assign wire7506 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n853) ) ;
 assign wire7508 = ( wire621  &  wire7505  &  wire7506 ) | ( wire622  &  wire7505  &  wire7506 ) ;
 assign wire7513 = ( (~ n_n852)  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire7514 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n858)  &  wire7513 ) ;
 assign wire7519 = ( n_n852  &  n_n854  &  (~ n_n855)  &  n_n856 ) ;
 assign wire7520 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n858)  &  wire7519 ) ;
 assign wire7522 = ( n_n852  &  (~ s298_in_1_) ) ;
 assign wire7523 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire7526 = ( (~ s298_out_3_)  &  (~ s298_out_5_)  &  wire7522  &  wire7523 ) ;
 assign wire7529 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n853) ) ;
 assign wire7530 = ( s298_in_1_  &  (~ n_n852)  &  wire7529 ) ;
 assign wire7531 = ( wire619  &  wire7530 ) | ( wire621  &  wire7530 ) | ( wire622  &  wire7530 ) ;
 assign wire7532 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7531 ) ;
 assign wire7537 = ( (~ n_n852)  &  n_n853  &  (~ n_n854)  &  n_n858 ) ;
 assign wire7538 = ( s298_in_0_  &  s298_in_1_  &  n_n859  &  wire7537 ) ;
 assign wire7542 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire7543 = ( n_n854  &  n_n857  &  wire7542 ) ;
 assign wire7549 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire7550 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire7549 ) ;
 assign wire7555 = ( (~ s298_in_1_)  &  (~ n_n853)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire7556 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858)  &  wire7555 ) ;
 assign wire7560 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n852  &  n_n853 ) ;
 assign wire7561 = ( (~ n_n855)  &  (~ n_n858)  &  wire7560 ) ;
 assign wire7567 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire7568 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire7567 ) ;
 assign wire7573 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire7574 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire7573 ) ;
 assign wire7579 = ( n_n852  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire7580 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856  &  wire7579 ) ;
 assign wire7585 = ( s298_in_1_  &  (~ n_n853)  &  n_n854  &  (~ n_n856) ) ;
 assign wire7586 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire7585 ) ;
 assign wire7591 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n855 ) ;
 assign wire7592 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856  &  wire7591 ) ;
 assign wire7597 = ( (~ s298_in_1_)  &  n_n852  &  n_n854  &  n_n855 ) ;
 assign wire7598 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858  &  wire7597 ) ;
 assign wire7601 = ( (~ n_n856)  &  (~ n_n855) ) ;
 assign wire7602 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n854) ) ;
 assign wire7604 = ( wire621  &  wire7601  &  wire7602 ) | ( wire622  &  wire7601  &  wire7602 ) ;
 assign wire7607 = ( (~ n_n856)  &  n_n854 ) ;
 assign wire7608 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7610 = ( wire621  &  wire7607  &  wire7608 ) | ( wire622  &  wire7607  &  wire7608 ) ;
 assign wire7613 = ( (~ n_n856)  &  n_n854 ) ;
 assign wire7614 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7616 = ( wire621  &  wire7613  &  wire7614 ) | ( wire622  &  wire7613  &  wire7614 ) ;
 assign wire7621 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire7622 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857  &  wire7621 ) ;
 assign wire7626 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire7627 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n853)  &  n_n856 ) ;
 assign wire7632 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire7633 = ( n_n853  &  n_n855  &  wire7632 ) ;
 assign wire7638 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n858) ) ;
 assign wire7639 = ( n_n852  &  n_n854  &  n_n855  &  (~ n_n856) ) ;
 assign wire7645 = ( s298_in_1_  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire7646 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858)  &  wire7645 ) ;
 assign wire7650 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire7651 = ( n_n854  &  n_n855  &  wire7650 ) ;
 assign wire7656 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856 ) ;
 assign wire7657 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire7662 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire7663 = ( n_n854  &  n_n857  &  wire7662 ) ;
 assign wire7664 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire7663 ) ;
 assign wire7668 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire7669 = ( n_n852  &  n_n853  &  n_n854  &  n_n858 ) ;
 assign wire7675 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n857 ) ;
 assign wire7676 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire7675 ) ;
 assign wire7681 = ( (~ n_n852)  &  n_n853  &  n_n854  &  n_n856 ) ;
 assign wire7682 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n857  &  wire7681 ) ;
 assign wire7686 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire7687 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  (~ n_n855) ) ;
 assign wire7693 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n852  &  (~ n_n853) ) ;
 assign wire7694 = ( (~ n_n854)  &  n_n857  &  (~ n_n858)  &  (~ n_n859) ) ;
 assign wire7699 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7700 = ( n_n853  &  (~ n_n854)  &  n_n857  &  (~ n_n859) ) ;
 assign wire7705 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852  &  (~ n_n853) ) ;
 assign wire7706 = ( n_n854  &  n_n856  &  n_n858  &  (~ n_n859) ) ;
 assign wire7711 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire7712 = ( n_n853  &  (~ n_n854)  &  n_n857  &  (~ n_n858) ) ;
 assign wire7717 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7718 = ( n_n853  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire7723 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire7724 = ( n_n853  &  (~ n_n855)  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire7727 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n854  &  (~ n_n855) ) ;
 assign wire7728 = ( wire580  &  wire7727 ) | ( wire581  &  wire7727 ) | ( wire582  &  wire7727 ) ;
 assign wire7729 = ( wire7728  &  n_n51 ) ;
 assign wire7732 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  (~ n_n855) ) ;
 assign wire7733 = ( wire621  &  wire7732 ) | ( wire622  &  wire7732 ) ;
 assign wire7734 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7733 ) ;
 assign wire7737 = ( s298_in_1_  &  n_n852  &  (~ n_n859) ) ;
 assign wire7738 = ( (~ n_n855)  &  n_n858  &  wire7737 ) ;
 assign wire7739 = ( wire6016  &  wire7738 ) | ( wire6017  &  wire7738 ) | ( wire6018  &  wire7738 ) ;
 assign wire7741 = ( (~ n_n856)  &  n_n853 ) ;
 assign wire7742 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n857) ) ;
 assign wire7744 = ( wire578  &  wire7741  &  wire7742 ) | ( wire579  &  wire7741  &  wire7742 ) ;
 assign wire7747 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire7748 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire7747 ) ;
 assign wire7749 = ( n_n51  &  wire7748 ) ;
 assign wire7752 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n857 ) ;
 assign wire7753 = ( (~ wire578)  &  (~ wire579)  &  wire7752 ) ;
 assign wire7754 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7753 ) ;
 assign wire7757 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n853  &  n_n854 ) ;
 assign wire7758 = ( wire578  &  wire7757 ) | ( wire579  &  wire7757 ) ;
 assign wire7759 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7758 ) ;
 assign wire7762 = ( s298_in_1_  &  n_n853  &  (~ n_n855)  &  n_n856 ) ;
 assign wire7763 = ( wire621  &  wire7762 ) | ( wire622  &  wire7762 ) ;
 assign wire7764 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7763 ) ;
 assign wire7766 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n854) ) ;
 assign wire7767 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire7766 ) ;
 assign wire7768 = ( n_n51  &  wire7767 ) ;
 assign wire7769 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7768 ) ;
 assign wire7772 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n852  &  (~ n_n855) ) ;
 assign wire7773 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire7772 ) ;
 assign wire7774 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire7773 ) ;
 assign wire7777 = ( s298_in_0_  &  s298_in_1_  &  n_n852  &  (~ n_n856) ) ;
 assign wire7778 = ( wire578  &  wire7777 ) | ( wire579  &  wire7777 ) ;
 assign wire7779 = ( wire6016  &  wire7778 ) | ( wire6017  &  wire7778 ) | ( wire6018  &  wire7778 ) ;
 assign wire7782 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n857) ) ;
 assign wire7783 = ( (~ n_n51)  &  wire7782 ) ;
 assign wire7784 = ( wire6016  &  wire7783 ) | ( wire6017  &  wire7783 ) | ( wire6018  &  wire7783 ) ;
 assign wire7786 = ( (~ n_n854)  &  (~ n_n852) ) ;
 assign wire7787 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n857) ) ;
 assign wire7789 = ( wire621  &  wire7786  &  wire7787 ) | ( wire622  &  wire7786  &  wire7787 ) ;
 assign wire7792 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n857) ) ;
 assign wire7794 = ( (~ s298_out_5_)  &  n_n853  &  n_n856  &  wire7792 ) ;
 assign wire7797 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n857 ) ;
 assign wire7799 = ( (~ n_n852)  &  (~ n_n856)  &  n_n51  &  wire7797 ) ;
 assign wire7802 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n856) ) ;
 assign wire7803 = ( (~ n_n852)  &  (~ n_n854)  &  wire7802 ) ;
 assign wire7804 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire7803 ) ;
 assign wire7808 = ( s298_in_0_  &  s298_in_1_  &  n_n852  &  n_n855 ) ;
 assign wire7809 = ( n_n856  &  (~ n_n857)  &  wire7808 ) ;
 assign wire7811 = ( (~ n_n854)  &  n_n853 ) ;
 assign wire7812 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n856) ) ;
 assign wire7814 = ( wire578  &  wire7811  &  wire7812 ) | ( wire579  &  wire7811  &  wire7812 ) ;
 assign wire7817 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n855 ) ;
 assign wire7818 = ( wire621  &  wire7817 ) | ( wire622  &  wire7817 ) ;
 assign wire7819 = ( wire5789  &  wire7818 ) | ( wire5790  &  wire7818 ) | ( wire5791  &  wire7818 ) ;
 assign wire7821 = ( n_n855  &  n_n852 ) ;
 assign wire7822 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n856) ) ;
 assign wire7824 = ( wire578  &  wire7821  &  wire7822 ) | ( wire579  &  wire7821  &  wire7822 ) ;
 assign wire7828 = ( (~ s298_in_1_)  &  (~ n_n853)  &  n_n854  &  n_n856 ) ;
 assign wire7829 = ( n_n857  &  (~ n_n858)  &  wire7828 ) ;
 assign wire7833 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n852  &  (~ n_n853) ) ;
 assign wire7834 = ( (~ n_n855)  &  n_n856  &  wire7833 ) ;
 assign wire7836 = ( n_n855  &  n_n853 ) ;
 assign wire7837 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n856 ) ;
 assign wire7839 = ( (~ wire578)  &  (~ wire579)  &  wire7836  &  wire7837 ) ;
 assign wire7842 = ( n_n857  &  n_n855 ) ;
 assign wire7843 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire7847 = ( n_n857  &  n_n855 ) ;
 assign wire7848 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire7851 = ( (~ s298_in_0_)  &  (~ n_n853)  &  n_n858 ) ;
 assign wire7853 = ( (~ s298_out_1_)  &  (~ wire621)  &  (~ wire622)  &  wire7851 ) ;
 assign wire7856 = ( s298_in_0_  &  n_n852  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire7857 = ( wire580  &  wire7856 ) | ( wire581  &  wire7856 ) | ( wire582  &  wire7856 ) ;
 assign wire7860 = ( (~ s298_in_1_)  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n51) ) ;
 assign wire7861 = ( wire6016  &  wire7860 ) | ( wire6017  &  wire7860 ) | ( wire6018  &  wire7860 ) ;
 assign wire7864 = ( s298_in_1_  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire7865 = ( wire578  &  wire7864 ) | ( wire579  &  wire7864 ) ;
 assign wire7868 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n855 ) ;
 assign wire7869 = ( wire578  &  wire7868 ) | ( wire579  &  wire7868 ) ;
 assign wire7872 = ( (~ s298_in_1_)  &  n_n854  &  n_n855  &  n_n856 ) ;
 assign wire7873 = ( wire621  &  wire7872 ) | ( wire622  &  wire7872 ) ;
 assign wire7876 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n859) ) ;
 assign wire7877 = ( (~ n_n852)  &  (~ n_n853)  &  wire7876 ) ;
 assign wire7880 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n859) ) ;
 assign wire7881 = ( (~ wire621)  &  (~ wire622)  &  wire7880 ) ;
 assign wire7884 = ( s298_out_0_  &  (~ n_n852)  &  n_n51  &  (~ n_n859) ) ;
 assign wire7886 = ( s298_in_1_  &  (~ n_n854)  &  (~ n_n857) ) ;
 assign wire7887 = ( wire621  &  wire7886 ) | ( wire622  &  wire7886 ) ;
 assign wire7889 = ( s298_in_1_  &  n_n855  &  (~ n_n856) ) ;
 assign wire7890 = ( wire621  &  wire7889 ) | ( wire622  &  wire7889 ) ;
 assign wire7892 = ( (~ n_n856)  &  n_n51  &  wire578 ) | ( (~ n_n856)  &  n_n51  &  wire579 ) ;
 assign wire7894 = ( n_n852  &  (~ n_n51)  &  (~ n_n859) ) ;
 assign wire7895 = ( wire7693  &  wire7694 ) | ( wire7699  &  wire7700 ) ;
 assign wire7896 = ( wire7705  &  wire7706 ) | ( wire7711  &  wire7712 ) ;
 assign wire7897 = ( wire7717  &  wire7718 ) | ( wire7723  &  wire7724 ) ;
 assign wire7902 = ( wire7897 ) | ( (~ s298_out_5_)  &  wire7243 ) ;
 assign wire7903 = ( (~ s298_out_5_)  &  wire7646 ) | ( (~ s298_out_5_)  &  wire7638  &  wire7639 ) ;
 assign wire7904 = ( wire230 ) | ( wire231 ) | ( wire232 ) | ( wire233 ) ;
 assign wire7905 = ( wire234 ) | ( wire279 ) | ( wire7895 ) | ( wire7896 ) ;
 assign wire7908 = ( (~ wire621)  &  (~ wire622)  &  wire7334 ) | ( (~ wire621)  &  (~ wire622)  &  wire7341 ) ;
 assign wire7909 = ( wire621  &  wire7622 ) | ( wire622  &  wire7622 ) | ( (~ wire621)  &  (~ wire622)  &  wire7598 ) ;
 assign wire7910 = ( wire269 ) | ( wire7902 ) | ( wire7903 ) ;
 assign wire7911 = ( wire214 ) | ( wire7904 ) | ( wire7905 ) ;
 assign wire7912 = ( s298_out_1_  &  wire7502 ) | ( s298_out_1_  &  s298_out_5_  &  wire7495 ) ;
 assign wire7913 = ( wire7909 ) | ( wire7908 ) ;
 assign wire7915 = ( (~ s298_out_5_)  &  n_n51  &  wire7633 ) | ( s298_out_5_  &  n_n51  &  wire7651 ) ;
 assign wire7916 = ( n_n51  &  wire7664 ) | ( (~ n_n51)  &  wire7656  &  wire7657 ) ;
 assign wire7917 = ( n_n51  &  wire7676 ) | ( n_n51  &  wire7668  &  wire7669 ) ;
 assign wire7918 = ( (~ n_n51)  &  wire7881 ) | ( n_n51  &  wire7847  &  wire7848 ) ;
 assign wire7921 = ( wire578  &  wire7313 ) | ( wire579  &  wire7313 ) | ( wire578  &  wire7320 ) | ( wire579  &  wire7320 ) ;
 assign wire7922 = ( s298_out_0_  &  wire7327 ) | ( (~ s298_out_0_)  &  (~ n_n51)  &  wire7543 ) ;
 assign wire7923 = ( (~ wire578)  &  (~ wire579)  &  wire7550 ) | ( (~ wire578)  &  (~ wire579)  &  wire7556 ) ;
 assign wire7924 = ( s298_out_0_  &  wire7568 ) | ( s298_out_0_  &  n_n51  &  wire7561 ) ;
 assign wire7925 = ( wire578  &  wire7574 ) | ( wire579  &  wire7574 ) | ( wire578  &  wire7580 ) | ( wire579  &  wire7580 ) ;
 assign wire7926 = ( wire578  &  wire7586 ) | ( wire579  &  wire7586 ) | ( wire578  &  wire7592 ) | ( wire579  &  wire7592 ) ;
 assign wire7927 = ( wire309 ) | ( wire7910 ) | ( (~ n_n51)  &  wire7355 ) ;
 assign wire7930 = ( wire218 ) | ( wire7911 ) | ( wire7912 ) | ( wire7913 ) ;
 assign wire7933 = ( wire7926 ) | ( wire7925 ) ;
 assign wire7935 = ( wire7917 ) | ( wire7918 ) | ( wire7930 ) ;
 assign wire7936 = ( wire7921 ) | ( wire7922 ) | ( wire7923 ) | ( wire7924 ) ;
 assign wire7937 = ( wire7915 ) | ( wire7916 ) | ( wire7927 ) | ( wire7933 ) ;
 assign wire7939 = ( wire7935 ) | ( wire7936 ) | ( wire7937 ) ;
 assign wire7945 = ( wire224 ) | ( wire226 ) | ( wire7939 ) ;
 assign wire7946 = ( wire227 ) | ( wire228 ) | ( wire229 ) | ( wire265 ) ;
 assign wire7947 = ( wire266 ) | ( wire267 ) | ( wire278 ) | ( wire308 ) ;
 assign wire7949 = ( wire7945 ) | ( wire7946 ) | ( wire7947 ) ;
 assign wire7959 = ( wire215 ) | ( wire216 ) | ( wire217 ) | ( wire7949 ) ;
 assign wire7960 = ( wire249 ) | ( wire250 ) | ( wire251 ) | ( wire252 ) ;
 assign wire7961 = ( wire253 ) | ( wire254 ) | ( wire303 ) | ( wire304 ) ;
 assign wire7962 = ( wire305 ) | ( wire306 ) | ( wire307 ) | ( wire320 ) ;
 assign wire7964 = ( wire7961 ) | ( wire7960 ) ;
 assign wire7965 = ( wire321 ) | ( wire323 ) | ( wire7959 ) | ( wire7962 ) ;
 assign wire7968 = ( (~ wire6375)  &  (~ wire6376)  &  wire7257 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7264 ) ;
 assign wire7969 = ( wire6375  &  wire7271 ) | ( wire6376  &  wire7271 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7424 ) ;
 assign wire7970 = ( (~ wire6375)  &  (~ wire6376)  &  wire7430 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7436 ) ;
 assign wire7971 = ( (~ wire6375)  &  (~ wire6376)  &  wire7442 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7448 ) ;
 assign wire7972 = ( (~ wire6375)  &  (~ wire6376)  &  wire7454 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7460 ) ;
 assign wire7973 = ( (~ wire6375)  &  (~ wire6376)  &  wire7466 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7472 ) ;
 assign wire7974 = ( wire6375  &  wire7484 ) | ( wire6376  &  wire7484 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7478 ) ;
 assign wire7975 = ( wire6375  &  wire7490 ) | ( wire6376  &  wire7490 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7729 ) ;
 assign wire7976 = ( (~ wire6375)  &  (~ wire6376)  &  wire7734 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7739 ) ;
 assign wire7977 = ( (~ wire6375)  &  (~ wire6376)  &  wire7744 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire7749 ) ;
 assign wire7978 = ( wire6375  &  wire7754 ) | ( wire6376  &  wire7754 ) | ( wire6375  &  wire7759 ) | ( wire6376  &  wire7759 ) ;
 assign wire7979 = ( wire6375  &  wire7764 ) | ( wire6376  &  wire7764 ) | ( wire6375  &  wire7769 ) | ( wire6376  &  wire7769 ) ;
 assign wire7980 = ( wire6375  &  wire7774 ) | ( wire6376  &  wire7774 ) | ( wire6375  &  wire7779 ) | ( wire6376  &  wire7779 ) ;
 assign wire7981 = ( wire6375  &  wire7784 ) | ( wire6376  &  wire7784 ) | ( wire6375  &  wire7789 ) | ( wire6376  &  wire7789 ) ;
 assign wire7982 = ( wire6375  &  wire7794 ) | ( wire6376  &  wire7794 ) | ( wire6375  &  wire7799 ) | ( wire6376  &  wire7799 ) ;
 assign wire7983 = ( wire6375  &  wire7804 ) | ( wire6376  &  wire7804 ) | ( wire6375  &  wire7809 ) | ( wire6376  &  wire7809 ) ;
 assign wire7984 = ( wire6375  &  wire7853 ) | ( wire6376  &  wire7853 ) | ( wire6375  &  wire7857 ) | ( wire6376  &  wire7857 ) ;
 assign wire7985 = ( wire6375  &  wire7861 ) | ( wire6376  &  wire7861 ) | ( wire6375  &  wire7865 ) | ( wire6376  &  wire7865 ) ;
 assign wire7986 = ( wire6375  &  wire7869 ) | ( wire6376  &  wire7869 ) | ( wire6375  &  wire7873 ) | ( wire6376  &  wire7873 ) ;
 assign wire7987 = ( wire6375  &  wire7877 ) | ( wire6376  &  wire7877 ) | ( wire6375  &  wire7884 ) | ( wire6376  &  wire7884 ) ;
 assign wire7988 = ( wire210 ) | ( wire322 ) | ( wire7964 ) | ( wire7965 ) ;
 assign wire7998 = ( wire7987 ) | ( wire7986 ) ;
 assign wire8000 = ( wire7970 ) | ( wire7971 ) | ( wire7972 ) | ( wire7973 ) ;
 assign wire8001 = ( wire7974 ) | ( wire7975 ) | ( wire7976 ) | ( wire7977 ) ;
 assign wire8002 = ( wire7978 ) | ( wire7979 ) | ( wire7980 ) | ( wire7981 ) ;
 assign wire8003 = ( wire7982 ) | ( wire7983 ) | ( wire7984 ) | ( wire7985 ) ;
 assign wire8004 = ( wire7968 ) | ( wire7969 ) | ( wire7988 ) | ( wire7998 ) ;
 assign wire8006 = ( wire8003 ) | ( wire8002 ) ;
 assign wire8012 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire8013 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire8015 = ( (~ wire621)  &  (~ wire622)  &  wire8012  &  wire8013 ) ;
 assign wire8019 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8021 = ( s298_out_5_  &  (~ n_n853)  &  (~ n_n854)  &  wire8019 ) ;
 assign wire8022 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8021 ) ;
 assign wire8026 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire8027 = ( (~ n_n854)  &  n_n855  &  wire8026 ) ;
 assign wire8029 = ( (~ n_n51)  &  wire578  &  wire8027 ) | ( (~ n_n51)  &  wire579  &  wire8027 ) ;
 assign wire8032 = ( n_n856  &  (~ n_n854) ) ;
 assign wire8033 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire8035 = ( wire621  &  wire8032  &  wire8033 ) | ( wire622  &  wire8032  &  wire8033 ) ;
 assign wire8036 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8035 ) ;
 assign wire8040 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire8041 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire8043 = ( (~ n_n51)  &  wire8040  &  wire8041 ) ;
 assign wire8048 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8049 = ( n_n853  &  (~ n_n854)  &  (~ n_n857)  &  (~ n_n858) ) ;
 assign wire8050 = ( wire8049  &  wire8048 ) ;
 assign wire8054 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8056 = ( (~ s298_out_3_)  &  n_n854  &  n_n855  &  wire8054 ) ;
 assign wire8057 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8056 ) ;
 assign wire8062 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire8063 = ( (~ n_n853)  &  (~ n_n854)  &  n_n855  &  n_n856 ) ;
 assign wire8064 = ( wire8063  &  wire8062 ) ;
 assign wire8069 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire8070 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n856  &  wire8069 ) ;
 assign wire8075 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire8076 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n855) ) ;
 assign wire8078 = ( (~ wire578)  &  (~ wire579)  &  wire8075  &  wire8076 ) ;
 assign wire8083 = ( (~ s298_in_1_)  &  (~ n_n853)  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire8084 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856  &  wire8083 ) ;
 assign wire8090 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852) ) ;
 assign wire8091 = ( (~ n_n853)  &  n_n854  &  n_n856  &  (~ n_n858) ) ;
 assign wire8092 = ( wire8091  &  wire8090 ) ;
 assign wire8097 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n853) ) ;
 assign wire8098 = ( n_n854  &  (~ n_n855)  &  n_n858  &  n_n859 ) ;
 assign wire8099 = ( wire8098  &  wire8097 ) ;
 assign wire8104 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8105 = ( (~ n_n854)  &  n_n855  &  n_n857  &  n_n858 ) ;
 assign wire8106 = ( wire8105  &  wire8104 ) ;
 assign wire8111 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8112 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n856)  &  (~ n_n857) ) ;
 assign wire8113 = ( wire8112  &  wire8111 ) ;
 assign wire8118 = ( n_n852  &  (~ n_n853)  &  n_n854  &  (~ n_n856) ) ;
 assign wire8119 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n857  &  wire8118 ) ;
 assign wire8120 = ( (~ wire619)  &  (~ wire621)  &  (~ wire622)  &  wire8119 ) ;
 assign wire8125 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire8126 = ( s298_in_1_  &  n_n852  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire8132 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire8133 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire8139 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire8140 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire8146 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire8147 = ( s298_in_1_  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire8153 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire8154 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire8160 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire8161 = ( s298_in_1_  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire8167 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire8168 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire8174 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n858) ) ;
 assign wire8175 = ( s298_in_1_  &  (~ n_n853)  &  n_n854  &  (~ n_n855) ) ;
 assign wire8180 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n852)  &  n_n855 ) ;
 assign wire8181 = ( (~ n_n857)  &  n_n859  &  wire8180 ) ;
 assign wire8182 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8181 ) ;
 assign wire8186 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n852)  &  n_n854 ) ;
 assign wire8187 = ( (~ n_n856)  &  (~ n_n858)  &  wire8186 ) ;
 assign wire8188 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8187 ) ;
 assign wire8192 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire8193 = ( (~ n_n854)  &  (~ n_n856)  &  wire8192 ) ;
 assign wire8194 = ( wire6016  &  wire8193 ) | ( wire6017  &  wire8193 ) | ( wire6018  &  wire8193 ) ;
 assign wire8198 = ( s298_in_0_  &  s298_in_1_  &  n_n853  &  (~ n_n854) ) ;
 assign wire8199 = ( (~ n_n855)  &  n_n856  &  wire8198 ) ;
 assign wire8200 = ( wire6016  &  wire8199 ) | ( wire6017  &  wire8199 ) | ( wire6018  &  wire8199 ) ;
 assign wire8202 = ( (~ n_n856)  &  (~ n_n853) ) ;
 assign wire8203 = ( (~ s298_in_0_)  &  n_n852  &  (~ n_n857) ) ;
 assign wire8206 = ( (~ s298_out_5_)  &  n_n51  &  wire8202  &  wire8203 ) ;
 assign wire8209 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire8211 = ( (~ s298_out_5_)  &  n_n854  &  (~ n_n855)  &  wire8209 ) ;
 assign wire8212 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8211 ) ;
 assign wire8216 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8218 = ( n_n856  &  n_n51  &  n_n858  &  wire8216 ) ;
 assign wire8222 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n854 ) ;
 assign wire8223 = ( n_n855  &  (~ n_n856)  &  wire8222 ) ;
 assign wire8224 = ( wire5789  &  wire8223 ) | ( wire5790  &  wire8223 ) | ( wire5791  &  wire8223 ) ;
 assign wire8229 = ( n_n852  &  (~ n_n854)  &  n_n855  &  (~ n_n856) ) ;
 assign wire8230 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire8229 ) ;
 assign wire8235 = ( n_n852  &  n_n853  &  n_n854  &  (~ n_n855) ) ;
 assign wire8236 = ( (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n858  &  wire8235 ) ;
 assign wire8240 = ( (~ s298_in_0_)  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire8242 = ( (~ s298_out_5_)  &  n_n855  &  n_n856  &  wire8240 ) ;
 assign wire8246 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n852  &  n_n854 ) ;
 assign wire8248 = ( (~ s298_out_5_)  &  (~ n_n855)  &  (~ n_n857)  &  wire8246 ) ;
 assign wire8252 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n852  &  n_n853 ) ;
 assign wire8254 = ( n_n856  &  (~ n_n857)  &  (~ n_n51)  &  wire8252 ) ;
 assign wire8258 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8259 = ( (~ n_n856)  &  (~ n_n857)  &  wire8258 ) ;
 assign wire8260 = ( wire5789  &  wire8259 ) | ( wire5790  &  wire8259 ) | ( wire5791  &  wire8259 ) ;
 assign wire8265 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n854)  &  n_n858 ) ;
 assign wire8266 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire8265 ) ;
 assign wire8269 = ( (~ n_n857)  &  (~ n_n855) ) ;
 assign wire8270 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  (~ n_n854) ) ;
 assign wire8272 = ( wire578  &  wire8269  &  wire8270 ) | ( wire579  &  wire8269  &  wire8270 ) ;
 assign wire8277 = ( (~ s298_in_1_)  &  (~ n_n852)  &  n_n853  &  n_n855 ) ;
 assign wire8278 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire8277 ) ;
 assign wire8281 = ( (~ n_n857)  &  n_n856 ) ;
 assign wire8282 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n854) ) ;
 assign wire8284 = ( wire578  &  wire8281  &  wire8282 ) | ( wire579  &  wire8281  &  wire8282 ) ;
 assign wire8287 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n857 ) ;
 assign wire8289 = ( (~ s298_out_5_)  &  (~ n_n852)  &  n_n853  &  wire8287 ) ;
 assign wire8290 = ( wire5789  &  wire8289 ) | ( wire5790  &  wire8289 ) | ( wire5791  &  wire8289 ) ;
 assign wire8294 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n853)  &  n_n855 ) ;
 assign wire8295 = ( (~ n_n856)  &  n_n857  &  wire8294 ) ;
 assign wire8296 = ( wire5789  &  wire8295 ) | ( wire5790  &  wire8295 ) | ( wire5791  &  wire8295 ) ;
 assign wire8299 = ( (~ s298_in_1_)  &  (~ n_n853)  &  (~ n_n859) ) ;
 assign wire8301 = ( (~ s298_out_3_)  &  n_n854  &  n_n857  &  wire8299 ) ;
 assign wire8302 = ( (~ wire578)  &  (~ wire579)  &  wire8301 ) ;
 assign wire8305 = ( n_n857  &  n_n855 ) ;
 assign wire8306 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n854) ) ;
 assign wire8308 = ( wire621  &  wire8305  &  wire8306 ) | ( wire622  &  wire8305  &  wire8306 ) ;
 assign wire8313 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire8314 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire8313 ) ;
 assign wire8319 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n854)  &  n_n856 ) ;
 assign wire8320 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire8319 ) ;
 assign wire8325 = ( n_n852  &  (~ n_n853)  &  n_n854  &  (~ n_n856) ) ;
 assign wire8326 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857  &  wire8325 ) ;
 assign wire8331 = ( (~ n_n852)  &  n_n853  &  n_n855  &  (~ n_n856) ) ;
 assign wire8332 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857  &  wire8331 ) ;
 assign wire8337 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  n_n855 ) ;
 assign wire8338 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire8337 ) ;
 assign wire8342 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire8343 = ( (~ n_n856)  &  (~ n_n857)  &  wire8342 ) ;
 assign wire8348 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8349 = ( (~ n_n856)  &  (~ n_n857)  &  wire8348 ) ;
 assign wire8354 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8356 = ( (~ s298_out_5_)  &  (~ n_n854)  &  n_n856  &  wire8354 ) ;
 assign wire8360 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859) ) ;
 assign wire8361 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n858 ) ;
 assign wire8367 = ( n_n852  &  n_n853  &  n_n854  &  n_n855 ) ;
 assign wire8368 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n858)  &  wire8367 ) ;
 assign wire8372 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire8373 = ( (~ n_n852)  &  n_n853  &  n_n854  &  (~ n_n855) ) ;
 assign wire8378 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire8379 = ( (~ s298_in_1_)  &  (~ n_n853)  &  n_n854  &  (~ n_n855) ) ;
 assign wire8385 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  (~ n_n854) ) ;
 assign wire8386 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855)  &  wire8385 ) ;
 assign wire8391 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire8392 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855)  &  wire8391 ) ;
 assign wire8397 = ( (~ n_n852)  &  (~ n_n853)  &  (~ n_n855)  &  n_n856 ) ;
 assign wire8398 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n857  &  wire8397 ) ;
 assign wire8403 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  n_n855 ) ;
 assign wire8404 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n859)  &  wire8403 ) ;
 assign wire8409 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8410 = ( (~ n_n853)  &  n_n855  &  (~ n_n856)  &  n_n859 ) ;
 assign wire8415 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8416 = ( (~ n_n854)  &  (~ n_n855)  &  n_n857  &  (~ n_n858) ) ;
 assign wire8421 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire8422 = ( n_n853  &  (~ n_n854)  &  (~ n_n855)  &  (~ n_n858) ) ;
 assign wire8427 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire8428 = ( n_n854  &  (~ n_n855)  &  n_n856  &  n_n857 ) ;
 assign wire8433 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8434 = ( (~ n_n853)  &  n_n854  &  n_n856  &  n_n858 ) ;
 assign wire8437 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n854) ) ;
 assign wire8438 = ( (~ s298_in_1_)  &  n_n853  &  wire8437 ) ;
 assign wire8439 = ( wire580  &  wire8438 ) | ( wire581  &  wire8438 ) | ( wire582  &  wire8438 ) ;
 assign wire8442 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire8443 = ( s298_in_1_  &  n_n852  &  wire8442 ) ;
 assign wire8444 = ( wire580  &  wire8443 ) | ( wire581  &  wire8443 ) | ( wire582  &  wire8443 ) ;
 assign wire8447 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n854  &  n_n856 ) ;
 assign wire8448 = ( wire621  &  wire8447 ) | ( wire622  &  wire8447 ) ;
 assign wire8449 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8448 ) ;
 assign wire8452 = ( s298_in_1_  &  (~ s298_out_3_)  &  (~ n_n853)  &  (~ n_n856) ) ;
 assign wire8453 = ( wire5789  &  wire8452 ) | ( wire5790  &  wire8452 ) | ( wire5791  &  wire8452 ) ;
 assign wire8454 = ( wire6016  &  wire8453 ) | ( wire6017  &  wire8453 ) | ( wire6018  &  wire8453 ) ;
 assign wire8456 = ( (~ n_n855)  &  n_n854 ) ;
 assign wire8457 = ( s298_in_0_  &  (~ n_n853)  &  (~ n_n858) ) ;
 assign wire8459 = ( (~ wire578)  &  (~ wire579)  &  wire8456  &  wire8457 ) ;
 assign wire8462 = ( s298_in_0_  &  n_n852  &  (~ n_n859) ) ;
 assign wire8463 = ( (~ n_n854)  &  n_n856  &  wire8462 ) ;
 assign wire8464 = ( wire5789  &  wire8463 ) | ( wire5790  &  wire8463 ) | ( wire5791  &  wire8463 ) ;
 assign wire8467 = ( n_n852  &  (~ n_n853)  &  n_n856 ) ;
 assign wire8468 = ( n_n854  &  n_n855  &  wire8467 ) ;
 assign wire8469 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8468 ) ;
 assign wire8472 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n854) ) ;
 assign wire8473 = ( wire578  &  wire8472 ) | ( wire579  &  wire8472 ) ;
 assign wire8474 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8473 ) ;
 assign wire8477 = ( s298_in_0_  &  (~ n_n852)  &  n_n854  &  (~ n_n858) ) ;
 assign wire8478 = ( wire578  &  wire8477 ) | ( wire579  &  wire8477 ) ;
 assign wire8479 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8478 ) ;
 assign wire8482 = ( (~ s298_in_0_)  &  n_n852  &  (~ n_n857) ) ;
 assign wire8483 = ( n_n855  &  n_n856  &  wire8482 ) ;
 assign wire8484 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8483 ) ;
 assign wire8487 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n852  &  n_n857 ) ;
 assign wire8488 = ( (~ n_n51)  &  wire8487 ) ;
 assign wire8489 = ( wire6016  &  wire8488 ) | ( wire6017  &  wire8488 ) | ( wire6018  &  wire8488 ) ;
 assign wire8492 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n856 ) ;
 assign wire8493 = ( (~ n_n853)  &  (~ n_n854)  &  wire8492 ) ;
 assign wire8494 = ( wire6016  &  wire8493 ) | ( wire6017  &  wire8493 ) | ( wire6018  &  wire8493 ) ;
 assign wire8496 = ( n_n855  &  (~ n_n852) ) ;
 assign wire8497 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n857 ) ;
 assign wire8499 = ( wire578  &  wire8496  &  wire8497 ) | ( wire579  &  wire8496  &  wire8497 ) ;
 assign wire8501 = ( (~ n_n855)  &  (~ n_n853) ) ;
 assign wire8502 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n858) ) ;
 assign wire8504 = ( wire578  &  wire8501  &  wire8502 ) | ( wire579  &  wire8501  &  wire8502 ) ;
 assign wire8506 = ( n_n853  &  (~ n_n852) ) ;
 assign wire8507 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n854) ) ;
 assign wire8509 = ( wire621  &  wire8506  &  wire8507 ) | ( wire622  &  wire8506  &  wire8507 ) ;
 assign wire8512 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  (~ n_n858) ) ;
 assign wire8514 = ( (~ s298_out_5_)  &  (~ n_n853)  &  n_n854  &  wire8512 ) ;
 assign wire8518 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n853  &  (~ n_n854) ) ;
 assign wire8519 = ( n_n856  &  n_n857  &  wire8518 ) ;
 assign wire8522 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n854)  &  (~ n_n855) ) ;
 assign wire8523 = ( wire621  &  wire8522 ) | ( wire622  &  wire8522 ) ;
 assign wire8524 = ( wire5789  &  wire8523 ) | ( wire5790  &  wire8523 ) | ( wire5791  &  wire8523 ) ;
 assign wire8526 = ( n_n854  &  n_n853 ) ;
 assign wire8527 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n855 ) ;
 assign wire8529 = ( wire621  &  wire8526  &  wire8527 ) | ( wire622  &  wire8526  &  wire8527 ) ;
 assign wire8531 = ( (~ n_n853)  &  (~ n_n852) ) ;
 assign wire8532 = ( s298_in_0_  &  s298_in_1_  &  n_n859 ) ;
 assign wire8534 = ( wire621  &  wire8531  &  wire8532 ) | ( wire622  &  wire8531  &  wire8532 ) ;
 assign wire8537 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n858) ) ;
 assign wire8539 = ( (~ s298_out_5_)  &  n_n852  &  n_n853  &  wire8537 ) ;
 assign wire8543 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n853  &  n_n854 ) ;
 assign wire8544 = ( n_n856  &  (~ n_n858)  &  wire8543 ) ;
 assign wire8548 = ( s298_in_0_  &  (~ n_n852)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire8549 = ( (~ n_n856)  &  (~ n_n858)  &  wire8548 ) ;
 assign wire8552 = ( (~ n_n858)  &  n_n855 ) ;
 assign wire8553 = ( (~ s298_in_0_)  &  (~ n_n852)  &  n_n853  &  n_n854 ) ;
 assign wire8558 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8559 = ( (~ n_n854)  &  n_n855  &  wire8558 ) ;
 assign wire8562 = ( n_n857  &  n_n855 ) ;
 assign wire8563 = ( (~ s298_in_2_)  &  s298_in_1_  &  n_n852  &  (~ n_n854) ) ;
 assign wire8568 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire8569 = ( (~ n_n855)  &  (~ n_n857)  &  wire8568 ) ;
 assign wire8571 = ( (~ s298_in_1_)  &  n_n853  &  n_n856 ) ;
 assign wire8572 = ( wire580  &  wire8571 ) | ( wire581  &  wire8571 ) | ( wire582  &  wire8571 ) ;
 assign wire8573 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8572 ) ;
 assign wire8575 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n855) ) ;
 assign wire8576 = ( wire580  &  wire8575 ) | ( wire581  &  wire8575 ) | ( wire582  &  wire8575 ) ;
 assign wire8577 = ( wire8576  &  n_n51 ) ;
 assign wire8580 = ( (~ s298_in_2_)  &  n_n854  &  (~ n_n857)  &  n_n51 ) ;
 assign wire8581 = ( wire6016  &  wire8580 ) | ( wire6017  &  wire8580 ) | ( wire6018  &  wire8580 ) ;
 assign wire8584 = ( (~ s298_in_1_)  &  n_n854  &  (~ n_n855)  &  (~ n_n857) ) ;
 assign wire8585 = ( wire6016  &  wire8584 ) | ( wire6017  &  wire8584 ) | ( wire6018  &  wire8584 ) ;
 assign wire8587 = ( (~ n_n852)  &  n_n858  &  (~ n_n859) ) ;
 assign wire8588 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8587 ) ;
 assign wire8589 = ( wire8588  &  n_n51 ) ;
 assign wire8591 = ( n_n852  &  n_n855  &  n_n856 ) ;
 assign wire8592 = ( wire621  &  wire8591 ) | ( wire622  &  wire8591 ) ;
 assign wire8593 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8592 ) ;
 assign wire8596 = ( (~ s298_in_1_)  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire8597 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8596 ) ;
 assign wire8600 = ( (~ s298_in_0_)  &  n_n853  &  n_n856  &  n_n857 ) ;
 assign wire8601 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8600 ) ;
 assign wire8604 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n859) ) ;
 assign wire8605 = ( (~ n_n852)  &  (~ n_n854)  &  wire8604 ) ;
 assign wire8608 = ( (~ s298_in_1_)  &  n_n852  &  n_n857 ) ;
 assign wire8609 = ( (~ n_n854)  &  (~ n_n855)  &  wire8608 ) ;
 assign wire8612 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n858) ) ;
 assign wire8613 = ( (~ n_n855)  &  n_n856  &  wire8612 ) ;
 assign wire8616 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire8617 = ( (~ n_n852)  &  (~ n_n853)  &  wire8616 ) ;
 assign wire8620 = ( s298_in_1_  &  n_n853  &  (~ n_n858) ) ;
 assign wire8621 = ( n_n855  &  n_n856  &  wire8620 ) ;
 assign wire8624 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n855) ) ;
 assign wire8626 = ( (~ s298_out_3_)  &  s298_in_2_ ) ;
 assign wire8627 = ( (~ wire580)  &  (~ wire581)  &  (~ wire582)  &  wire8626 ) ;
 assign wire8630 = ( (~ s298_in_2_)  &  (~ n_n853)  &  (~ n_n859) ) ;
 assign wire8631 = ( wire578  &  wire8630 ) | ( wire579  &  wire8630 ) ;
 assign wire8633 = ( s298_in_2_  &  n_n854  &  wire621 ) | ( s298_in_2_  &  n_n854  &  wire622 ) ;
 assign wire8635 = ( s298_in_2_  &  n_n51  &  (~ wire621)  &  (~ wire622) ) ;
 assign wire8637 = ( (~ n_n855)  &  (~ n_n857)  &  n_n859 ) ;
 assign wire8638 = ( (~ n_n858)  &  s298_in_2_ ) ;
 assign wire8639 = ( wire8409  &  wire8410 ) | ( wire8415  &  wire8416 ) ;
 assign wire8640 = ( wire8421  &  wire8422 ) | ( wire8427  &  wire8428 ) ;
 assign wire8647 = ( (~ s298_out_5_)  &  wire8368 ) | ( (~ s298_out_5_)  &  wire8360  &  wire8361 ) ;
 assign wire8648 = ( (~ s298_out_5_)  &  wire8549 ) | ( s298_out_5_  &  wire8372  &  wire8373 ) ;
 assign wire8649 = ( (~ s298_out_5_)  &  wire8621 ) | ( (~ s298_out_5_)  &  wire8552  &  wire8553 ) ;
 assign wire8650 = ( wire111 ) | ( wire112 ) | ( wire113 ) | ( wire161 ) ;
 assign wire8651 = ( wire114 ) | ( wire115 ) | ( wire116 ) | ( wire117 ) ;
 assign wire8652 = ( wire118 ) | ( wire202 ) | ( wire8639 ) | ( wire8640 ) ;
 assign wire8656 = ( wire621  &  wire8314 ) | ( wire622  &  wire8314 ) | ( wire621  &  wire8320 ) | ( wire622  &  wire8320 ) ;
 assign wire8657 = ( wire621  &  wire8326 ) | ( wire622  &  wire8326 ) | ( wire621  &  wire8332 ) | ( wire622  &  wire8332 ) ;
 assign wire8658 = ( wire621  &  wire8338 ) | ( wire622  &  wire8338 ) | ( wire621  &  wire8638 ) | ( wire622  &  wire8638 ) ;
 assign wire8659 = ( wire8647 ) | ( wire8648 ) | ( wire8649 ) | ( wire8650 ) ;
 assign wire8660 = ( wire133 ) | ( wire8651 ) | ( wire8652 ) ;
 assign wire8661 = ( wire156 ) | ( s298_out_1_  &  wire8633 ) ;
 assign wire8664 = ( (~ s298_out_5_)  &  n_n51  &  wire8343 ) | ( (~ s298_out_5_)  &  n_n51  &  wire8349 ) ;
 assign wire8665 = ( n_n51  &  wire8559 ) | ( (~ n_n51)  &  wire8378  &  wire8379 ) ;
 assign wire8666 = ( n_n51  &  wire8569 ) | ( n_n51  &  wire8562  &  wire8563 ) ;
 assign wire8668 = ( wire8656 ) | ( wire8657 ) | ( wire8661 ) ;
 assign wire8670 = ( s298_out_0_  &  wire8092 ) | ( s298_out_0_  &  (~ n_n51)  &  wire8084 ) ;
 assign wire8671 = ( (~ wire578)  &  (~ wire579)  &  wire8544 ) | ( (~ wire578)  &  (~ wire579)  &  wire8613 ) ;
 assign wire8672 = ( s298_out_0_  &  wire8617 ) | ( (~ s298_out_0_)  &  n_n51  &  wire8627 ) ;
 assign wire8674 = ( wire8660 ) | ( wire8666 ) | ( n_n51  &  wire8637 ) ;
 assign wire8675 = ( wire103 ) | ( wire8658 ) | ( wire8659 ) | ( wire8668 ) ;
 assign wire8676 = ( wire8671 ) | ( wire8670 ) ;
 assign wire8677 = ( wire8664 ) | ( wire8665 ) | ( wire8672 ) ;
 assign wire8680 = ( wire8674 ) | ( wire8675 ) | ( wire8676 ) | ( wire8677 ) ;
 assign wire8687 = ( wire104 ) | ( wire107 ) | ( wire108 ) | ( wire8680 ) ;
 assign wire8688 = ( wire109 ) | ( wire110 ) | ( wire139 ) | ( wire140 ) ;
 assign wire8689 = ( wire148 ) | ( wire153 ) | ( wire154 ) | ( wire155 ) ;
 assign wire8691 = ( wire8687 ) | ( wire8688 ) | ( wire8689 ) ;
 assign wire8698 = ( wire206 ) | ( wire204 ) ;
 assign wire8699 = ( wire101 ) | ( wire102 ) | ( wire134 ) | ( wire8691 ) ;
 assign wire8700 = ( wire135 ) | ( wire136 ) | ( wire137 ) | ( wire138 ) ;
 assign wire8701 = ( wire179 ) | ( wire180 ) | ( wire181 ) | ( wire182 ) ;
 assign wire8704 = ( wire8698 ) | ( wire8699 ) | ( wire8700 ) | ( wire8701 ) ;
 assign wire8705 = ( wire8704 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8015 ) ;
 assign wire8706 = ( (~ wire6375)  &  (~ wire6376)  &  wire8022 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8029 ) ;
 assign wire8707 = ( (~ wire6375)  &  (~ wire6376)  &  wire8036 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8043 ) ;
 assign wire8708 = ( (~ wire6375)  &  (~ wire6376)  &  wire8050 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8182 ) ;
 assign wire8709 = ( (~ wire6375)  &  (~ wire6376)  &  wire8188 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8194 ) ;
 assign wire8710 = ( (~ wire6375)  &  (~ wire6376)  &  wire8200 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8206 ) ;
 assign wire8711 = ( (~ wire6375)  &  (~ wire6376)  &  wire8212 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8218 ) ;
 assign wire8712 = ( (~ wire6375)  &  (~ wire6376)  &  wire8224 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8230 ) ;
 assign wire8713 = ( wire6375  &  wire8242 ) | ( wire6376  &  wire8242 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8236 ) ;
 assign wire8714 = ( wire6375  &  wire8248 ) | ( wire6376  &  wire8248 ) | ( wire6375  &  wire8254 ) | ( wire6376  &  wire8254 ) ;
 assign wire8715 = ( wire6375  &  wire8260 ) | ( wire6376  &  wire8260 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8439 ) ;
 assign wire8716 = ( (~ wire6375)  &  (~ wire6376)  &  wire8444 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8449 ) ;
 assign wire8717 = ( (~ wire6375)  &  (~ wire6376)  &  wire8454 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8459 ) ;
 assign wire8718 = ( wire6375  &  wire8469 ) | ( wire6376  &  wire8469 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8464 ) ;
 assign wire8719 = ( wire6375  &  wire8474 ) | ( wire6376  &  wire8474 ) | ( wire6375  &  wire8479 ) | ( wire6376  &  wire8479 ) ;
 assign wire8720 = ( wire6375  &  wire8484 ) | ( wire6376  &  wire8484 ) | ( wire6375  &  wire8489 ) | ( wire6376  &  wire8489 ) ;
 assign wire8721 = ( wire6375  &  wire8494 ) | ( wire6376  &  wire8494 ) | ( wire6375  &  wire8499 ) | ( wire6376  &  wire8499 ) ;
 assign wire8722 = ( wire6375  &  wire8504 ) | ( wire6376  &  wire8504 ) | ( wire6375  &  wire8509 ) | ( wire6376  &  wire8509 ) ;
 assign wire8723 = ( wire6375  &  wire8514 ) | ( wire6376  &  wire8514 ) | ( wire6375  &  wire8519 ) | ( wire6376  &  wire8519 ) ;
 assign wire8724 = ( (~ wire6375)  &  (~ wire6376)  &  wire8573 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8577 ) ;
 assign wire8725 = ( (~ wire6375)  &  (~ wire6376)  &  wire8581 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8585 ) ;
 assign wire8726 = ( wire6375  &  wire8589 ) | ( wire6376  &  wire8589 ) | ( wire6375  &  wire8593 ) | ( wire6376  &  wire8593 ) ;
 assign wire8727 = ( wire6375  &  wire8597 ) | ( wire6376  &  wire8597 ) | ( wire6375  &  wire8601 ) | ( wire6376  &  wire8601 ) ;
 assign wire8728 = ( wire6375  &  wire8605 ) | ( wire6376  &  wire8605 ) | ( wire6375  &  wire8609 ) | ( wire6376  &  wire8609 ) ;
 assign wire8741 = ( wire8705 ) | ( wire8706 ) | ( wire8707 ) | ( wire8708 ) ;
 assign wire8742 = ( wire8709 ) | ( wire8710 ) | ( wire8711 ) | ( wire8712 ) ;
 assign wire8743 = ( wire8713 ) | ( wire8714 ) | ( wire8715 ) | ( wire8716 ) ;
 assign wire8744 = ( wire8717 ) | ( wire8718 ) | ( wire8719 ) | ( wire8720 ) ;
 assign wire8745 = ( wire8721 ) | ( wire8722 ) | ( wire8723 ) | ( wire8724 ) ;
 assign wire8746 = ( wire8725 ) | ( wire8726 ) | ( wire8727 ) | ( wire8728 ) ;
 assign wire8750 = ( wire8741 ) | ( wire8742 ) | ( wire8743 ) | ( wire8744 ) ;
 assign wire8755 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire8756 = ( (~ s298_in_1_)  &  n_n852  &  n_n853  &  (~ n_n854) ) ;
 assign wire8758 = ( (~ n_n855)  &  n_n856  &  wire8755  &  wire8756 ) ;
 assign wire8763 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire8764 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n857)  &  wire8763 ) ;
 assign wire8765 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8764 ) ;
 assign wire8769 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n858) ) ;
 assign wire8770 = ( (~ n_n852)  &  (~ n_n854)  &  (~ n_n855)  &  n_n857 ) ;
 assign wire8772 = ( wire578  &  wire8769  &  wire8770 ) | ( wire579  &  wire8769  &  wire8770 ) ;
 assign wire8776 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire8777 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  (~ n_n854) ) ;
 assign wire8779 = ( s298_out_5_  &  wire8776  &  wire8777 ) ;
 assign wire8783 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n858 ) ;
 assign wire8784 = ( (~ s298_in_1_)  &  n_n852  &  (~ n_n855)  &  (~ n_n856) ) ;
 assign wire8786 = ( (~ s298_out_3_)  &  wire8783  &  wire8784 ) ;
 assign wire8791 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n853) ) ;
 assign wire8792 = ( (~ n_n855)  &  n_n856  &  n_n858  &  n_n859 ) ;
 assign wire8793 = ( wire8792  &  wire8791 ) ;
 assign wire8798 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n859 ) ;
 assign wire8799 = ( s298_in_1_  &  n_n852  &  n_n853  &  n_n854 ) ;
 assign wire8802 = ( (~ n_n852)  &  (~ s298_in_1_) ) ;
 assign wire8803 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n857 ) ;
 assign wire8805 = ( wire621  &  wire8802  &  wire8803 ) | ( wire622  &  wire8802  &  wire8803 ) ;
 assign wire8806 = ( wire5789  &  wire8805 ) | ( wire5790  &  wire8805 ) | ( wire5791  &  wire8805 ) ;
 assign wire8809 = ( n_n855  &  (~ n_n854) ) ;
 assign wire8810 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n852 ) ;
 assign wire8812 = ( wire621  &  wire8809  &  wire8810 ) | ( wire622  &  wire8809  &  wire8810 ) ;
 assign wire8815 = ( (~ n_n856)  &  n_n854 ) ;
 assign wire8816 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8818 = ( wire621  &  wire8815  &  wire8816 ) | ( wire622  &  wire8815  &  wire8816 ) ;
 assign wire8820 = ( (~ n_n854)  &  (~ s298_in_1_) ) ;
 assign wire8821 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n857) ) ;
 assign wire8824 = ( (~ s298_out_5_)  &  n_n51  &  wire8820  &  wire8821 ) ;
 assign wire8828 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n852) ) ;
 assign wire8830 = ( n_n854  &  n_n51  &  (~ n_n858)  &  wire8828 ) ;
 assign wire8833 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n854 ) ;
 assign wire8835 = ( (~ n_n852)  &  n_n853  &  n_n51  &  wire8833 ) ;
 assign wire8836 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8835 ) ;
 assign wire8840 = ( s298_in_0_  &  s298_in_1_  &  n_n853  &  (~ n_n855) ) ;
 assign wire8841 = ( n_n857  &  (~ n_n858)  &  wire8840 ) ;
 assign wire8842 = ( wire6016  &  wire8841 ) | ( wire6017  &  wire8841 ) | ( wire6018  &  wire8841 ) ;
 assign wire8846 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8847 = ( (~ n_n856)  &  (~ n_n857)  &  wire8846 ) ;
 assign wire8848 = ( wire5789  &  wire8847 ) | ( wire5790  &  wire8847 ) | ( wire5791  &  wire8847 ) ;
 assign wire8852 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire8854 = ( (~ n_n854)  &  n_n856  &  n_n51  &  wire8852 ) ;
 assign wire8859 = ( s298_in_1_  &  (~ n_n852)  &  (~ n_n854)  &  n_n856 ) ;
 assign wire8860 = ( s298_in_0_  &  (~ s298_in_2_)  &  n_n858  &  wire8859 ) ;
 assign wire8864 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8866 = ( (~ n_n855)  &  (~ n_n51)  &  (~ n_n858)  &  wire8864 ) ;
 assign wire8870 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  n_n856 ) ;
 assign wire8871 = ( s298_in_1_  &  n_n852  &  (~ n_n853)  &  (~ n_n855) ) ;
 assign wire8877 = ( (~ s298_in_1_)  &  (~ n_n852)  &  (~ n_n853)  &  n_n854 ) ;
 assign wire8878 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ n_n856)  &  wire8877 ) ;
 assign wire8882 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n856) ) ;
 assign wire8883 = ( s298_in_1_  &  (~ n_n853)  &  n_n854  &  n_n855 ) ;
 assign wire8887 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n854) ) ;
 assign wire8888 = ( n_n852  &  n_n853  &  wire8887 ) ;
 assign wire8889 = ( wire619  &  wire8888 ) | ( wire621  &  wire8888 ) | ( wire622  &  wire8888 ) ;
 assign wire8890 = ( wire8889  &  n_n51 ) ;
 assign wire8893 = ( (~ s298_in_2_)  &  s298_in_1_  &  (~ n_n854)  &  n_n855 ) ;
 assign wire8894 = ( wire580  &  wire8893 ) | ( wire581  &  wire8893 ) | ( wire582  &  wire8893 ) ;
 assign wire8895 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8894 ) ;
 assign wire8898 = ( (~ s298_in_2_)  &  n_n853  &  (~ n_n854)  &  (~ n_n857) ) ;
 assign wire8899 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire8898 ) ;
 assign wire8900 = ( n_n51  &  wire8899 ) ;
 assign wire8902 = ( (~ s298_in_2_)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire8904 = ( (~ s298_out_3_)  &  (~ s298_out_5_)  &  wire8902 ) ;
 assign wire8905 = ( wire5789  &  wire8904 ) | ( wire5790  &  wire8904 ) | ( wire5791  &  wire8904 ) ;
 assign wire8908 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  n_n852 ) ;
 assign wire8909 = ( (~ n_n51)  &  wire8908 ) ;
 assign wire8910 = ( wire5789  &  wire8909 ) | ( wire5790  &  wire8909 ) | ( wire5791  &  wire8909 ) ;
 assign wire8913 = ( (~ s298_in_2_)  &  (~ n_n853)  &  n_n859 ) ;
 assign wire8914 = ( n_n855  &  (~ n_n856)  &  wire8913 ) ;
 assign wire8915 = ( wire5789  &  wire8914 ) | ( wire5790  &  wire8914 ) | ( wire5791  &  wire8914 ) ;
 assign wire8918 = ( (~ s298_in_2_)  &  n_n853  &  n_n859 ) ;
 assign wire8919 = ( (~ n_n855)  &  (~ n_n856)  &  wire8918 ) ;
 assign wire8920 = ( wire5789  &  wire8919 ) | ( wire5790  &  wire8919 ) | ( wire5791  &  wire8919 ) ;
 assign wire8923 = ( (~ s298_in_0_)  &  s298_in_1_  &  n_n857 ) ;
 assign wire8924 = ( n_n852  &  (~ n_n855)  &  wire8923 ) ;
 assign wire8925 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire8924 ) ;
 assign wire8927 = ( n_n854  &  (~ n_n852) ) ;
 assign wire8928 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n857 ) ;
 assign wire8930 = ( (~ wire578)  &  (~ wire579)  &  wire8927  &  wire8928 ) ;
 assign wire8932 = ( (~ n_n855)  &  (~ n_n852) ) ;
 assign wire8933 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n856) ) ;
 assign wire8935 = ( wire578  &  wire8932  &  wire8933 ) | ( wire579  &  wire8932  &  wire8933 ) ;
 assign wire8938 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n857) ) ;
 assign wire8940 = ( (~ n_n853)  &  (~ n_n854)  &  (~ n_n51)  &  wire8938 ) ;
 assign wire8943 = ( s298_in_0_  &  (~ s298_in_1_)  &  n_n857 ) ;
 assign wire8944 = ( n_n852  &  n_n853  &  wire8943 ) ;
 assign wire8945 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8944 ) ;
 assign wire8948 = ( s298_in_0_  &  (~ s298_in_2_)  &  (~ s298_in_1_)  &  (~ n_n853) ) ;
 assign wire8949 = ( wire580  &  wire8948 ) | ( wire581  &  wire8948 ) | ( wire582  &  wire8948 ) ;
 assign wire8950 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire8949 ) ;
 assign wire8954 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire8955 = ( (~ n_n854)  &  n_n856  &  wire8954 ) ;
 assign wire8959 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire8960 = ( n_n855  &  n_n856  &  wire8959 ) ;
 assign wire8964 = ( (~ s298_in_2_)  &  (~ n_n853)  &  (~ n_n854)  &  n_n855 ) ;
 assign wire8965 = ( n_n856  &  (~ n_n857)  &  wire8964 ) ;
 assign wire8969 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n852)  &  n_n854 ) ;
 assign wire8970 = ( (~ n_n855)  &  (~ n_n859)  &  wire8969 ) ;
 assign wire8974 = ( s298_in_0_  &  s298_in_1_  &  (~ n_n852)  &  (~ n_n853) ) ;
 assign wire8975 = ( n_n854  &  (~ n_n857)  &  wire8974 ) ;
 assign wire8979 = ( s298_in_0_  &  (~ s298_in_1_)  &  (~ n_n852)  &  n_n853 ) ;
 assign wire8980 = ( (~ n_n855)  &  n_n858  &  wire8979 ) ;
 assign wire8983 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n853  &  (~ n_n855) ) ;
 assign wire8984 = ( wire8983  &  (~ s298_out_3_) ) ;
 assign wire8989 = ( s298_in_0_  &  (~ s298_in_2_)  &  s298_in_1_  &  n_n853 ) ;
 assign wire8990 = ( n_n856  &  (~ n_n858)  &  wire8989 ) ;
 assign wire8993 = ( (~ s298_in_0_)  &  (~ s298_in_1_)  &  n_n852  &  (~ n_n853) ) ;
 assign wire8994 = ( wire619  &  wire8993 ) | ( wire621  &  wire8993 ) | ( wire622  &  wire8993 ) ;
 assign wire8995 = ( wire8994  &  n_n51 ) ;
 assign wire8998 = ( (~ n_n857)  &  (~ n_n856) ) ;
 assign wire8999 = ( (~ s298_in_2_)  &  n_n853  &  n_n854  &  (~ n_n855) ) ;
 assign wire9004 = ( (~ s298_in_2_)  &  n_n852  &  (~ n_n853)  &  n_n854 ) ;
 assign wire9005 = ( n_n855  &  (~ n_n857)  &  wire9004 ) ;
 assign wire9010 = ( s298_in_1_  &  (~ n_n852)  &  n_n853  &  (~ n_n854) ) ;
 assign wire9012 = ( (~ s298_in_2_)  &  (~ n_n852)  &  n_n856 ) ;
 assign wire9013 = ( wire621  &  wire9012 ) | ( wire622  &  wire9012 ) ;
 assign wire9014 = ( (~ wire6016)  &  (~ wire6017)  &  (~ wire6018)  &  wire9013 ) ;
 assign wire9017 = ( (~ s298_in_2_)  &  n_n853  &  n_n855  &  (~ n_n857) ) ;
 assign wire9018 = ( wire621  &  wire9017 ) | ( wire622  &  wire9017 ) ;
 assign wire9021 = ( (~ s298_in_2_)  &  n_n852  &  n_n854  &  (~ n_n856) ) ;
 assign wire9022 = ( wire5789  &  wire9021 ) | ( wire5790  &  wire9021 ) | ( wire5791  &  wire9021 ) ;
 assign wire9025 = ( s298_in_0_  &  (~ n_n854)  &  (~ n_n856)  &  (~ n_n858) ) ;
 assign wire9026 = ( wire6016  &  wire9025 ) | ( wire6017  &  wire9025 ) | ( wire6018  &  wire9025 ) ;
 assign wire9029 = ( (~ s298_in_0_)  &  s298_in_1_  &  (~ n_n853)  &  n_n856 ) ;
 assign wire9030 = ( wire6016  &  wire9029 ) | ( wire6017  &  wire9029 ) | ( wire6018  &  wire9029 ) ;
 assign wire9032 = ( (~ n_n853)  &  n_n854  &  n_n856 ) ;
 assign wire9033 = ( (~ wire621)  &  (~ wire622)  &  wire9032 ) ;
 assign wire9034 = ( wire5789  &  wire9033 ) | ( wire5790  &  wire9033 ) | ( wire5791  &  wire9033 ) ;
 assign wire9035 = ( n_n853  &  (~ s298_in_0_) ) ;
 assign wire9036 = ( wire623  &  wire9035 ) | ( wire624  &  wire9035 ) | ( wire625  &  wire9035 ) ;
 assign wire9037 = ( wire580  &  wire9036 ) | ( wire581  &  wire9036 ) | ( wire582  &  wire9036 ) ;
 assign wire9038 = ( (~ wire5789)  &  (~ wire5790)  &  (~ wire5791)  &  wire9037 ) ;
 assign wire9040 = ( (~ s298_in_1_)  &  n_n855  &  (~ n_n859) ) ;
 assign wire9041 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire9040 ) ;
 assign wire9042 = ( wire5789  &  wire9041 ) | ( wire5790  &  wire9041 ) | ( wire5791  &  wire9041 ) ;
 assign wire9044 = ( n_n855  &  n_n856  &  (~ n_n858) ) ;
 assign wire9045 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire9044 ) ;
 assign wire9046 = ( wire5789  &  wire9045 ) | ( wire5790  &  wire9045 ) | ( wire5791  &  wire9045 ) ;
 assign wire9049 = ( n_n852  &  (~ n_n854)  &  n_n856  &  n_n858 ) ;
 assign wire9050 = ( wire5789  &  wire9049 ) | ( wire5790  &  wire9049 ) | ( wire5791  &  wire9049 ) ;
 assign wire9053 = ( (~ s298_in_0_)  &  (~ s298_in_2_)  &  (~ n_n854)  &  (~ n_n856) ) ;
 assign wire9057 = ( (~ s298_in_2_)  &  n_n853  &  n_n857 ) ;
 assign wire9058 = ( n_n855  &  (~ n_n856)  &  wire9057 ) ;
 assign wire9059 = ( n_n854  &  n_n852 ) ;
 assign wire9060 = ( wire580  &  wire9059 ) | ( wire581  &  wire9059 ) | ( wire582  &  wire9059 ) ;
 assign wire9061 = ( wire6016  &  wire9060 ) | ( wire6017  &  wire9060 ) | ( wire6018  &  wire9060 ) ;
 assign wire9063 = ( n_n853  &  n_n854  &  n_n856 ) ;
 assign wire9064 = ( (~ wire578)  &  (~ wire579)  &  wire9063 ) ;
 assign wire9066 = ( n_n852  &  n_n856  &  n_n858 ) ;
 assign wire9067 = ( (~ wire578)  &  (~ wire579)  &  wire9066 ) ;
 assign wire9070 = ( (~ n_n855)  &  n_n856  &  n_n858  &  n_n859 ) ;
 assign wire9072 = ( s298_in_0_  &  (~ n_n852)  &  n_n853 ) ;
 assign wire9073 = ( wire580  &  wire9072 ) | ( wire581  &  wire9072 ) | ( wire582  &  wire9072 ) ;
 assign wire9075 = ( (~ s298_in_1_)  &  n_n854  &  (~ n_n858) ) ;
 assign wire9076 = ( (~ wire578)  &  (~ wire579)  &  wire9075 ) ;
 assign wire9079 = ( s298_out_0_  &  n_n855  &  (~ n_n857)  &  n_n51 ) ;
 assign wire9081 = ( n_n853  &  (~ n_n854)  &  (~ n_n856) ) ;
 assign wire9082 = ( wire578  &  wire9081 ) | ( wire579  &  wire9081 ) ;
 assign wire9084 = ( (~ s298_in_1_)  &  n_n853  &  (~ n_n858) ) ;
 assign wire9085 = ( wire621  &  wire9084 ) | ( wire622  &  wire9084 ) ;
 assign wire9087 = ( (~ s298_in_0_)  &  n_n854  &  (~ n_n858) ) ;
 assign wire9088 = ( (~ wire623)  &  (~ wire624)  &  (~ wire625)  &  wire9087 ) ;
 assign wire9089 = ( (~ n_n51)  &  (~ n_n859) ) ;
 assign wire9090 = ( wire6016  &  wire9089 ) | ( wire6017  &  wire9089 ) | ( wire6018  &  wire9089 ) ;
 assign wire9092 = ( (~ n_n854)  &  (~ n_n855)  &  n_n858 ) ;
 assign wire9094 = ( wire30 ) | ( wire69 ) | ( (~ s298_out_5_)  &  wire8990 ) ;
 assign wire9096 = ( wire58 ) | ( wire24 ) ;
 assign wire9097 = ( wire81 ) | ( wire59 ) ;
 assign wire9098 = ( wire44 ) | ( wire9094 ) | ( n_n51  &  wire8786 ) ;
 assign wire9099 = ( wire9096 ) | ( n_n51  &  wire8998  &  wire8999 ) ;
 assign wire9101 = ( s298_out_0_  &  wire8878 ) | ( (~ s298_out_0_)  &  n_n51  &  wire8984 ) ;
 assign wire9104 = ( wire80 ) | ( wire9098 ) | ( wire9101 ) ;
 assign wire9105 = ( wire42 ) | ( wire9097 ) | ( wire9099 ) | ( wire9104 ) ;
 assign wire9109 = ( wire27 ) | ( wire29 ) | ( wire45 ) | ( wire9105 ) ;
 assign wire9110 = ( wire66 ) | ( wire68 ) | ( wire9109 ) ;
 assign wire9121 = ( wire39 ) | ( wire40 ) | ( wire41 ) | ( wire9110 ) ;
 assign wire9122 = ( wire57 ) | ( wire60 ) | ( wire61 ) | ( wire62 ) ;
 assign wire9123 = ( wire63 ) | ( wire76 ) | ( wire77 ) | ( wire78 ) ;
 assign wire9124 = ( wire79 ) | ( wire86 ) | ( wire87 ) | ( wire88 ) ;
 assign wire9125 = ( wire89 ) | ( wire90 ) | ( wire91 ) | ( wire94 ) ;
 assign wire9128 = ( wire9121 ) | ( wire9122 ) | ( wire9125 ) ;
 assign wire9129 = ( wire9123 ) | ( wire9124 ) | ( wire9128 ) ;
 assign wire9131 = ( (~ wire6375)  &  (~ wire6376)  &  wire8772 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8806 ) ;
 assign wire9132 = ( (~ wire6375)  &  (~ wire6376)  &  wire8812 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8818 ) ;
 assign wire9133 = ( (~ wire6375)  &  (~ wire6376)  &  wire8824 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8830 ) ;
 assign wire9134 = ( wire6375  &  wire8836 ) | ( wire6376  &  wire8836 ) | ( wire6375  &  wire8842 ) | ( wire6376  &  wire8842 ) ;
 assign wire9135 = ( wire6375  &  wire8848 ) | ( wire6376  &  wire8848 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8895 ) ;
 assign wire9136 = ( (~ wire6375)  &  (~ wire6376)  &  wire8900 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8905 ) ;
 assign wire9137 = ( (~ wire6375)  &  (~ wire6376)  &  wire8910 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8915 ) ;
 assign wire9138 = ( wire6375  &  wire8925 ) | ( wire6376  &  wire8925 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire8920 ) ;
 assign wire9139 = ( wire6375  &  wire8930 ) | ( wire6376  &  wire8930 ) | ( wire6375  &  wire8935 ) | ( wire6376  &  wire8935 ) ;
 assign wire9140 = ( wire6375  &  wire8940 ) | ( wire6376  &  wire8940 ) | ( wire6375  &  wire8945 ) | ( wire6376  &  wire8945 ) ;
 assign wire9141 = ( (~ wire6375)  &  (~ wire6376)  &  wire9014 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire9018 ) ;
 assign wire9142 = ( wire6375  &  wire9026 ) | ( wire6376  &  wire9026 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire9022 ) ;
 assign wire9143 = ( wire6375  &  wire9030 ) | ( wire6376  &  wire9030 ) | ( wire6375  &  wire9034 ) | ( wire6376  &  wire9034 ) ;
 assign wire9144 = ( wire6375  &  wire9064 ) | ( wire6376  &  wire9064 ) | ( (~ wire6375)  &  (~ wire6376)  &  wire9061 ) ;
 assign wire9145 = ( wire6375  &  wire9067 ) | ( wire6376  &  wire9067 ) | ( wire6375  &  wire9070 ) | ( wire6376  &  wire9070 ) ;
 assign wire9146 = ( wire6375  &  wire9090 ) | ( wire6376  &  wire9090 ) | ( wire6375  &  wire9092 ) | ( wire6376  &  wire9092 ) ;
 assign wire9155 = ( wire25 ) | ( wire9129 ) | ( wire9131 ) | ( wire9146 ) ;
 assign wire9156 = ( wire9132 ) | ( wire9133 ) | ( wire9134 ) | ( wire9135 ) ;
 assign wire9157 = ( wire9136 ) | ( wire9137 ) | ( wire9138 ) | ( wire9139 ) ;
 assign wire9158 = ( wire9140 ) | ( wire9141 ) | ( wire9142 ) | ( wire9143 ) ;
 assign wire9161 = ( wire9144 ) | ( wire9145 ) | ( wire9155 ) | ( wire9158 ) ;


endmodule

