module diffeq (
	tin_puport_10_10_, tin_puport_0_0_, tin_pxport_10_10_, tin_pxport_0_0_, pdxport_4_4_, tin_puport_1_1_, tin_pxport_1_1_, tin_puport_2_2_, 
	tin_pyport_10_10_, tin_pyport_0_0_, tin_pxport_2_2_, preset_0_0_, pdxport_5_5_, tin_puport_3_3_, tin_pyport_1_1_, paport_11_11_, pready_0_0_, paport_6_6_, 
	pdxport_6_6_, paport_7_7_, paport_8_8_, pdxport_7_7_, paport_9_9_, tin_pxport_7_7_, tin_puport_8_8_, tin_pyport_6_6_, paport_2_2_, tin_pxport_8_8_, 
	pdxport_8_8_, pdxport_0_0_, pclk, tin_puport_9_9_, tin_pyport_7_7_, paport_3_3_, tin_pxport_9_9_, tin_pyport_8_8_, paport_4_4_, pdxport_9_9_, 
	pdxport_1_1_, tin_pyport_9_9_, paport_5_5_, tin_pxport_3_3_, tin_puport_4_4_, tin_pyport_2_2_, tin_pxport_4_4_, pdxport_2_2_, tin_puport_11_11_, tin_puport_5_5_, 
	tin_pyport_3_3_, tin_pxport_5_5_, pdxport_11_11_, pdxport_10_10_, tin_puport_6_6_, tin_pyport_4_4_, paport_10_10_, paport_0_0_, preset, tin_pxport_11_11_, 
	tin_pxport_6_6_, pdxport_3_3_, tin_puport_7_7_, tin_pyport_11_11_, tin_pyport_5_5_, paport_1_1_, puport_10_10_, puport_0_0_, pxport_10_10_, pxport_0_0_, 
	puport_1_1_, pxport_1_1_, puport_2_2_, pyport_10_10_, pyport_0_0_, pxport_2_2_, puport_3_3_, pyport_1_1_, pnext_0_0_, pxport_7_7_, 
	puport_8_8_, pyport_6_6_, pxport_8_8_, puport_9_9_, pyport_7_7_, pxport_9_9_, pover_0_0_, pyport_8_8_, pyport_9_9_, pxport_3_3_, 
	puport_4_4_, pyport_2_2_, pdn, pxport_4_4_, puport_11_11_, puport_5_5_, pyport_3_3_, pxport_5_5_, puport_6_6_, pyport_4_4_, 
	pxport_11_11_, pxport_6_6_, puport_7_7_, pyport_11_11_, pyport_5_5_);

input tin_puport_10_10_;
input tin_puport_0_0_;
input tin_pxport_10_10_;
input tin_pxport_0_0_;
input pdxport_4_4_;
input tin_puport_1_1_;
input tin_pxport_1_1_;
input tin_puport_2_2_;
input tin_pyport_10_10_;
input tin_pyport_0_0_;
input tin_pxport_2_2_;
input preset_0_0_;
input pdxport_5_5_;
input tin_puport_3_3_;
input tin_pyport_1_1_;
input paport_11_11_;
input pready_0_0_;
input paport_6_6_;
input pdxport_6_6_;
input paport_7_7_;
input paport_8_8_;
input pdxport_7_7_;
input paport_9_9_;
input tin_pxport_7_7_;
input tin_puport_8_8_;
input tin_pyport_6_6_;
input paport_2_2_;
input tin_pxport_8_8_;
input pdxport_8_8_;
input pdxport_0_0_;
input pclk;
input tin_puport_9_9_;
input tin_pyport_7_7_;
input paport_3_3_;
input tin_pxport_9_9_;
input tin_pyport_8_8_;
input paport_4_4_;
input pdxport_9_9_;
input pdxport_1_1_;
input tin_pyport_9_9_;
input paport_5_5_;
input tin_pxport_3_3_;
input tin_puport_4_4_;
input tin_pyport_2_2_;
input tin_pxport_4_4_;
input pdxport_2_2_;
input tin_puport_11_11_;
input tin_puport_5_5_;
input tin_pyport_3_3_;
input tin_pxport_5_5_;
input pdxport_11_11_;
input pdxport_10_10_;
input tin_puport_6_6_;
input tin_pyport_4_4_;
input paport_10_10_;
input paport_0_0_;
input preset;
input tin_pxport_11_11_;
input tin_pxport_6_6_;
input pdxport_3_3_;
input tin_puport_7_7_;
input tin_pyport_11_11_;
input tin_pyport_5_5_;
input paport_1_1_;
output puport_10_10_;
output puport_0_0_;
output pxport_10_10_;
output pxport_0_0_;
output puport_1_1_;
output pxport_1_1_;
output puport_2_2_;
output pyport_10_10_;
output pyport_0_0_;
output pxport_2_2_;
output puport_3_3_;
output pyport_1_1_;
output pnext_0_0_;
output pxport_7_7_;
output puport_8_8_;
output pyport_6_6_;
output pxport_8_8_;
output puport_9_9_;
output pyport_7_7_;
output pxport_9_9_;
output pover_0_0_;
output pyport_8_8_;
output pyport_9_9_;
output pxport_3_3_;
output puport_4_4_;
output pyport_2_2_;
output pdn;
output pxport_4_4_;
output puport_11_11_;
output puport_5_5_;
output pyport_3_3_;
output pxport_5_5_;
output puport_6_6_;
output pyport_4_4_;
output pxport_11_11_;
output pxport_6_6_;
output puport_7_7_;
output pyport_11_11_;
output pyport_5_5_;
wire n_n3032;
wire n_n2959;
wire n_n3174;
wire n_n2952;
wire n_n2973;
wire n_n3488;
wire n_n3596;
wire n_n3969;
wire n_n2970;
wire n_n3259;
wire n_n4007;
wire n_n3483;
wire n_n3073;
wire n_n3653;
wire n_n3051;
wire n_n3137;
wire n_n4098;
wire n_n3007;
wire n_n3086;
wire n_n3602;
wire n_n3499;
wire n_n3956;
wire n_n3752;
wire n_n3941;
wire n_n3299;
wire n_n3284;
wire n_n3618;
wire n_n3353;
wire n_n2972;
wire n_n3070;
wire n_n3454;
wire n_n3640;
wire n_n2992;
wire n_n3063;
wire n_n4147;
wire n_n3772;
wire n_n3132;
wire n_n2969;
wire n_n3616;
wire n_n3183;
wire n_n3523;
wire n_n3004;
wire n_n3206;
wire n_n2984;
wire n_n4038;
wire n_n3481;
wire n_n3322;
wire n_n3144;
wire n_n3401;
wire n_n3584;
wire n_n3926;
wire n_n2958;
wire n_n3739;
wire n_n2990;
wire n_n3744;
wire n_n3690;
wire n_n3018;
wire n_n3334;
wire n_n2997;
wire n_n3566;
wire n_n3798;
wire n_n2974;
wire n_n3115;
wire n_n3811;
wire n_n3059;
wire n_n3325;
wire n_n3052;
wire n_n3030;
wire n_n3153;
wire n_n3705;
wire n_n3432;
wire n_n2983;
wire n_n3040;
wire n_n3209;
wire n_n3165;
wire n_n3057;
wire n_n3127;
wire n_n4254;
wire n_n3163;
wire n_n3041;
wire n_n3972;
wire n_n3150;
wire n_n3814;
wire n_n3349;
wire n_n3247;
wire n_n3661;
wire n_n3652;
wire n_n3315;
wire n_n3316;
wire n_n3456;
wire n_n3168;
wire n_n3037;
wire n_n3119;
wire n_n2966;
wire n_n3795;
wire n_n4113;
wire n_n3014;
wire n_n3103;
wire n_n4238;
wire n_n3210;
wire n_n3113;
wire n_n3740;
wire n_n3202;
wire n_n3720;
wire n_n3314;
wire n_n3650;
wire n_n3046;
wire n_n3458;
wire n_n3409;
wire n_n3227;
wire n_n2963;
wire n_n3005;
wire n_n2998;
wire n_n3638;
wire n_n4063;
wire n_n3240;
wire n_n3987;
wire n_n3177;
wire n_n2996;
wire n_n3061;
wire n_n3091;
wire n_n3178;
wire n_n3193;
wire n_n3016;
wire n_n3712;
wire n_n4053;
wire n_n3310;
wire n_n3431;
wire n_n3599;
wire n_n3146;
wire n_n3058;
wire n_n3914;
wire n_n3389;
wire n_n3379;
wire n_n3633;
wire n_n3147;
wire n_n3586;
wire n_n4089;
wire n_n3963;
wire n_n3213;
wire n_n3538;
wire n_n4055;
wire n_n3009;
wire n_n3050;
wire n_n4229;
wire n_n3595;
wire n_n3245;
wire n_n2955;
wire n_n3172;
wire n_n3710;
wire n_n2979;
wire n_n3012;
wire n_n3397;
wire n_n3211;
wire n_n3863;
wire n_n4029;
wire n_n3487;
wire n_n4085;
wire n_n3664;
wire n_n3609;
wire n_n3266;
wire n_n3658;
wire n_n3244;
wire n_n3200;
wire n_n2985;
wire n_n2957;
wire n_n3348;
wire n_n3683;
wire n_n3615;
wire n_n4231;
wire n_n3287;
wire n_n3049;
wire n_n3558;
wire n_n3263;
wire n_n3946;
wire n_n3614;
wire n_n3437;
wire n_n3180;
wire n_n2978;
wire n_n4256;
wire n_n4139;
wire n_n3853;
wire n_n3530;
wire n_n4011;
wire n_n3648;
wire n_n3064;
wire n_n3276;
wire n_n3570;
wire n_n3339;
wire n_n3524;
wire n_n3241;
wire n_n2956;
wire n_n3145;
wire n_n3592;
wire n_n3102;
wire n_n3093;
wire n_n3191;
wire n_n3476;
wire n_n4041;
wire n_n3479;
wire n_n3895;
wire n_n3158;
wire n_n3249;
wire n_n3717;
wire n_n3106;
wire n_n4020;
wire n_n3765;
wire n_n2999;
wire n_n3909;
wire n_n3726;
wire n_n4110;
wire n_n3620;
wire n_n2980;
wire n_n3696;
wire n_n4105;
wire n_n4094;
wire n_n3497;
wire n_n3692;
wire n_n3308;
wire n_n3847;
wire n_n3801;
wire n_n3162;
wire n_n3189;
wire n_n3465;
wire n_n3043;
wire n_n4174;
wire n_n2976;
wire n_n3008;
wire n_n4032;
wire n_n3305;
wire n_n3204;
wire n_n3028;
wire n_n3075;
wire n_n3087;
wire n_n3326;
wire n_n3817;
wire n_n3136;
wire n_n3668;
wire n_n3068;
wire n_n3413;
wire n_n3222;
wire n_n3627;
wire n_n3399;
wire n_n2994;
wire n_n2987;
wire n_n3429;
wire n_n3372;
wire n_n3915;
wire n_n3452;
wire n_n3447;
wire n_n3156;
wire n_n3201;
wire n_n3472;
wire n_n3611;
wire n_n4074;
wire n_n3449;
wire n_n3904;
wire n_n3542;
wire n_n2964;
wire n_n4028;
wire n_n3423;
wire n_n2977;
wire n_n3130;
wire n_n3042;
wire n_n3338;
wire n_n3078;
wire n_n3374;
wire n_n3425;
wire n_n3486;
wire n_n3104;
wire n_n3129;
wire n_n3152;
wire n_n3053;
wire n_n3133;
wire n_n3770;
wire n_n3003;
wire n_n3010;
wire n_n3666;
wire n_n3605;
wire n_n3899;
wire n_n2961;
wire n_n4166;
wire n_n3511;
wire n_n3022;
wire n_n3155;
wire n_n3117;
wire n_n3027;
wire n_n3885;
wire n_n3335;
wire n_n3197;
wire n_n3034;
wire n_n2962;
wire n_n3823;
wire n_n3160;
wire n_n3029;
wire n_n3406;
wire n_n3787;
wire n_n3506;
wire n_n3216;
wire n_n3215;
wire n_n3721;
wire n_n3173;
wire n_n3785;
wire n_n3277;
wire n_n3562;
wire n_n4023;
wire n_n3015;
wire n_n3120;
wire n_n3621;
wire n_n3645;
wire n_n2965;
wire n_n3913;
wire n_n3695;
wire n_n4217;
wire n_n3416;
wire n_n3687;
wire n_n3320;
wire n_n3559;
wire n_n4044;
wire n_n3435;
wire n_n3967;
wire n_n3352;
wire n_n3321;
wire n_n3318;
wire n_n3066;
wire n_n2967;
wire n_n3707;
wire n_n3194;
wire n_n3825;
wire n_n3123;
wire n_n3579;
wire n_n3491;
wire n_n3980;
wire n_n3859;
wire n_n3723;
wire n_n3231;
wire n_n3400;
wire n_n3048;
wire n_n3804;
wire n_n3001;
wire n_n2953;
wire n_n2981;
wire n_n3850;
wire n_n3332;
wire n_n2988;
wire n_n3390;
wire n_n3589;
wire n_n3192;
wire n_n3273;
wire n_n2975;
wire n_n3662;
wire n_n3038;
wire n_n3671;
wire n_n3190;
wire n_n3101;
wire n_n3366;
wire n_n3958;
wire n_n4046;
wire n_n3503;
wire n_n4065;
wire n_n3474;
wire n_n47;
wire n_n36;
wire n_n41;
wire n_n3828;
wire n_n3553;
wire n_n40;
wire n_n3754;
wire n_n3555;
wire n_n39;
wire n_n44;
wire n_n45;
wire n_n38;
wire n_n43;
wire n_n46;
wire n_n37;
wire n_n42;
wire wire806;
wire n_n3827;
wire wire802;
wire wire811;
wire n_n4170;
wire wire797;
wire wire918;
wire wire799;
wire wire857;
wire n_n4008;
wire n_n4144;
wire n_n3948;
wire n_n4131;
wire wire813;
wire wire875;
wire wire860;
wire wire862;
wire n_n4000;
wire wire796;
wire n_n3944;
wire n_n3301;
wire wire839;
wire wire816;
wire n_n3975;
wire n_n4168;
wire n_n4084;
wire n_n4082;
wire n_n3099;
wire n_n3920;
wire n_n4211;
wire wire838;
wire wire940;
wire n_n4151;
wire wire869;
wire n_n4017;
wire n_n4219;
wire n_n3888;
wire wire870;
wire n_n3746;
wire n_n4245;
wire n_n3643;
wire n_n3142;
wire n_n3869;
wire wire917;
wire n_n3925;
wire n_n4019;
wire wire907;
wire n_n3966;
wire n_n3837;
wire n_n3991;
wire n_n4196;
wire n_n4198;
wire nak3_9;
wire n_n4146;
wire n_n3403;
wire n_n4253;
wire n_n4069;
wire n_n4115;
wire n_n3565;
wire n_n4178;
wire n_n4125;
wire wire841;
wire n_n3993;
wire n_n3833;
wire n_n3549;
wire n_n3903;
wire n_n3439;
wire nrq5_5;
wire nrq5_2;
wire n_n4228;
wire n_n3359;
wire wire945;
wire n_n3404;
wire n_n3779;
wire wire877;
wire n_n4129;
wire wire878;
wire n_n4189;
wire nrq5_9;
wire wire809;
wire wire879;
wire wire923;
wire n_n4184;
wire n_n3118;
wire n_n3857;
wire n_n3135;
wire wire880;
wire wire916;
wire wire955;
wire wire926;
wire ndn_latch5_5;
wire nrq5_6;
wire wire844;
wire n_n4052;
wire n_n3363;
wire wire845;
wire n_n3729;
wire nrq2_2;
wire ndn_latch5_3;
wire ndn_latch5_8;
wire wire946;
wire wire947;
wire ndn_latch5_2;
wire wire883;
wire n_n3892;
wire nrq5_10;
wire ndn_latch5_4;
wire ndn_latch5_7;
wire n_n4123;
wire wire914;
wire n_n4160;
wire n_n3532;
wire wire846;
wire n_n3236;
wire n_n3434;
wire wire948;
wire n_n3281;
wire wire886;
wire n_n4202;
wire n_n3897;
wire n_n3883;
wire wire818;
wire wire989;
wire n_n3762;
wire n_n3396;
wire wire939;
wire wire975;
wire n_n3581;
wire wire843;
wire wire929;
wire n_n3950;
wire n_n3976;
wire wire949;
wire wire950;
wire wire951;
wire n_n3521;
wire n_n4200;
wire n_n3569;
wire n_n3111;
wire wire849;
wire n_n3025;
wire wire850;
wire n_n3955;
wire n_n4248;
wire wire890;
wire wire930;
wire n_n3484;
wire wire931;
wire wire952;
wire wire932;
wire n_n4062;
wire n_n3512;
wire wire953;
wire wire933;
wire n_n3543;
wire wire851;
wire n_n4051;
wire wire934;
wire n_n4153;
wire wire852;
wire n_n3035;
wire n_n3635;
wire n_n3748;
wire wire935;
wire wire817;
wire wire936;
wire wire835;
wire wire876;
wire wire938;
wire wire954;
wire wire963;
wire wire964;
wire wire970;
wire wire971;
wire wire972;
wire wire973;
wire wire976;
wire wire977;
wire wire979;
wire wire980;
wire wire983;
wire wire985;
wire wire987;
wire wire988;
wire wire991;
wire wire992;
wire wire993;
wire wire996;
wire wire998;
wire wire999;
wire wire1000;
wire wire1002;
wire wire1003;
wire wire1007;
wire wire1008;
wire wire1017;
wire wire1018;
wire wire1020;
wire wire1023;
wire wire1026;
wire wire1032;
wire wire1034;
wire wire1037;
wire wire1041;
wire wire1042;
wire wire1043;
wire wire1044;
wire wire1045;
wire wire1049;
wire wire1050;
wire wire1052;
wire wire1056;
wire wire1057;
wire wire1058;
wire wire1060;
wire wire1061;
wire wire1062;
wire wire1063;
wire wire1064;
wire wire1065;
wire wire1067;
wire wire1071;
wire wire1073;
wire wire1076;
wire wire1078;
wire wire1081;
wire wire1084;
wire wire1086;
wire wire1087;
wire wire1089;
wire wire1093;
wire wire1097;
wire wire1098;
wire wire1099;
wire wire1104;
wire wire1105;
wire wire1106;
wire wire1108;
wire wire1110;
wire wire1111;
wire wire1114;
wire wire1115;
wire wire1117;
wire wire1120;
wire wire1124;
wire wire1125;
wire wire1129;
wire wire1131;
wire wire1132;
wire wire1133;
wire wire1134;
wire wire1136;
wire wire1137;
wire wire1138;
wire wire1141;
wire wire1145;
wire wire1146;
wire wire1147;
wire wire1148;
wire wire1151;
wire wire1152;
wire wire1153;
wire wire1154;
wire wire1155;
wire wire1156;
wire wire1157;
wire wire1159;
wire wire1160;
wire wire1161;
wire wire1162;
wire wire1163;
wire wire1166;
wire wire1169;
wire wire1170;
wire wire1174;
wire wire1176;
wire wire1179;
wire wire1180;
wire wire1184;
wire wire1187;
wire wire1188;
wire wire1190;
wire wire1194;
wire wire1195;
wire wire1197;
wire wire1200;
wire wire1203;
wire wire1204;
wire wire1205;
wire wire1208;
wire wire1210;
wire wire1213;
wire wire1214;
wire wire1215;
wire wire1216;
wire wire1217;
wire wire1218;
wire wire1219;
wire wire1221;
wire wire1223;
wire wire1226;
wire wire1227;
wire wire1232;
wire wire1233;
wire wire1235;
wire wire1240;
wire wire1241;
wire wire1243;
wire wire1246;
wire wire1247;
wire wire1248;
wire wire1249;
wire wire1250;
wire wire1251;
wire wire1253;
wire wire1254;
wire wire1256;
wire wire1258;
wire wire1259;
wire wire1261;
wire wire1262;
wire wire1263;
wire wire1264;
wire wire1265;
wire wire1267;
wire wire1268;
wire wire1270;
wire wire1271;
wire wire1273;
wire wire1276;
wire wire1279;
wire wire1282;
wire wire1286;
wire wire1297;
wire wire1302;
wire wire1303;
wire wire1304;
wire wire1308;
wire wire1312;
wire wire1313;
wire wire1314;
wire wire1315;
wire wire1316;
wire wire1317;
wire wire1319;
wire wire1320;
wire wire1321;
wire wire1322;
wire wire1323;
wire wire1324;
wire wire1327;
wire wire1328;
wire wire1338;
wire wire1341;
wire wire1344;
wire wire1345;
wire wire1346;
wire wire1347;
wire wire1348;
wire wire1349;
wire wire1352;
wire wire1353;
wire wire1354;
wire wire1355;
wire wire1356;
wire wire1361;
wire wire1362;
wire wire1363;
wire wire1364;
wire wire1365;
wire wire1366;
wire wire1367;
wire wire1368;
wire wire1369;
wire wire1370;
wire wire1371;
wire wire1372;
wire wire1373;
wire wire1374;
wire wire1375;
wire wire1376;
wire wire1378;
wire wire1379;
wire wire1381;
wire wire1384;
wire wire1385;
wire wire1386;
wire wire1387;
wire wire1388;
wire wire1390;
wire wire1391;
wire wire1393;
wire wire1395;
wire wire1396;
wire wire1398;
wire wire1401;
wire wire1402;
wire wire1403;
wire wire1405;
wire wire1406;
wire wire1407;
wire wire1408;
wire wire1411;
wire wire1413;
wire wire1418;
wire wire1419;
wire wire1421;
wire wire1422;
wire wire1423;
wire wire1426;
wire wire1427;
wire wire1430;
wire wire1431;
wire wire1432;
wire wire1435;
wire wire1436;
wire wire1437;
wire wire1440;
wire wire1441;
wire wire1443;
wire wire1445;
wire wire1446;
wire wire1447;
wire wire1448;
wire wire1450;
wire wire1451;
wire wire1453;
wire wire1454;
wire wire1456;
wire wire1457;
wire wire1460;
wire wire1461;
wire wire1464;
wire wire1465;
wire wire1467;
wire wire1468;
wire wire1469;
wire wire1470;
wire wire1472;
wire wire1475;
wire wire1476;
wire wire1477;
wire wire1495;
wire wire1500;
wire wire1503;
wire wire1505;
wire wire1507;
wire wire1508;
wire wire1509;
wire wire1511;
wire wire1514;
wire wire1517;
wire wire1520;
wire wire1526;
wire wire1528;
wire wire1530;
wire wire1534;
wire wire1535;
wire wire1539;
wire wire1540;
wire wire1544;
wire wire1545;
wire wire1546;
wire wire1548;
wire wire1553;
wire wire1559;
wire wire1562;
wire wire1564;
wire wire1567;
wire wire1568;
wire wire1571;
wire wire1572;
wire wire1574;
wire wire1577;
wire wire1578;
wire wire1582;
wire wire1585;
wire wire1586;
wire wire1588;
wire wire1589;
wire wire1590;
wire wire1592;
wire wire1596;
wire wire1597;
wire wire1598;
wire wire1599;
wire wire1600;
wire wire1602;
wire wire1605;
wire wire1606;
wire wire1607;
wire wire1608;
wire wire1610;
wire wire1613;
wire wire1614;
wire wire1617;
wire wire1618;
wire wire1619;
wire wire1622;
wire wire1623;
wire wire1624;
wire wire1625;
wire wire1626;
wire wire1631;
wire wire1636;
wire wire1638;
wire wire1639;
wire wire1642;
wire wire1643;
wire wire1645;
wire wire1646;
wire wire1647;
wire wire1649;
wire wire1650;
wire wire1652;
wire wire1654;
wire wire1656;
wire wire1657;
wire wire1660;
wire wire1666;
wire wire1667;
wire wire1669;
wire wire1670;
wire wire1671;
wire wire1672;
wire wire1674;
wire wire1675;
wire wire1677;
wire wire1678;
wire wire1686;
wire wire1687;
wire wire1690;
wire wire1693;
wire wire1694;
wire wire1697;
wire wire1700;
wire wire1701;
wire wire1702;
wire wire1705;
wire wire1708;
wire wire1721;
wire wire1722;
wire wire1723;
wire wire1729;
wire wire1730;
wire wire1733;
wire wire1734;
wire wire1735;
wire wire1736;
wire wire1737;
wire wire1745;
wire wire1751;
wire wire1752;
wire wire1754;
wire wire1769;
wire wire1775;
wire wire1776;
wire wire1777;
wire wire1780;
wire wire1781;
wire wire1783;
wire wire1784;
wire wire1785;
wire wire1787;
wire wire1790;
wire wire1794;
wire wire1795;
wire wire1797;
wire wire1802;
wire wire1803;
wire wire1804;
wire wire1805;
wire wire1806;
wire wire1807;
wire wire1809;
wire wire1814;
wire wire1815;
wire wire1816;
wire wire1819;
wire wire1823;
wire wire1826;
wire wire1827;
wire wire1828;
wire wire1829;
wire wire1831;
wire wire1832;
wire wire1835;
wire wire1836;
wire wire1841;
wire wire1842;
wire wire1844;
wire wire1848;
wire wire1851;
wire wire1855;
wire wire1857;
wire wire1859;
wire wire1860;
wire wire1865;
wire wire1866;
wire wire1867;
wire wire1870;
wire wire1873;
wire wire1877;
wire wire1879;
wire wire1882;
wire wire1886;
wire wire1889;
wire wire1890;
wire wire1894;
wire wire1898;
wire wire1902;
wire wire1904;
wire wire1905;
wire wire1906;
wire wire1908;
wire wire1915;
wire wire1929;
wire wire1937;
wire wire1938;
wire wire1944;
wire wire1948;
wire wire1950;
wire wire1955;
wire wire1956;
wire wire1959;
wire wire1960;
wire wire1963;
wire wire1966;
wire wire1967;
wire wire1968;
wire wire1969;
wire wire1970;
wire wire1971;
wire wire1974;
wire wire1975;
wire wire1976;
wire wire1977;
wire wire1978;
wire wire1983;
wire wire1984;
wire wire1985;
wire wire1986;
wire wire1987;
wire wire1990;
wire wire1991;
wire wire1992;
wire wire1993;
wire wire1994;
wire wire1999;
wire wire2000;
wire wire2001;
wire wire2002;
wire wire2003;
wire wire2007;
wire wire2008;
wire wire2009;
wire wire2010;
wire wire2011;
wire wire2012;
wire wire2013;
wire wire2014;
wire wire2015;
wire wire2016;
wire wire2017;
wire wire2018;
wire wire2019;
wire wire2020;
wire wire2021;
wire wire2022;
wire wire2023;
wire wire2024;
wire wire2025;
wire wire2026;
wire wire2028;
wire wire2031;
wire wire2034;
wire wire2035;
wire wire2036;
wire wire2037;
wire wire2038;
wire wire2039;
wire wire2041;
wire wire2046;
wire wire2051;
wire wire2057;
wire wire2058;
wire wire2059;
wire wire2060;
wire wire2061;
wire wire2063;
wire wire2064;
wire wire2066;
wire wire2068;
wire wire2069;
wire wire2071;
wire wire2073;
wire wire2074;
wire wire2075;
wire wire2080;
wire wire2085;
wire wire2090;
wire wire2096;
wire wire2101;
wire wire2103;
wire wire2104;
wire wire2107;
wire wire2112;
wire wire2118;
wire wire2123;
wire wire2129;
wire wire2134;
wire wire2136;
wire wire2137;
wire wire2140;
wire wire2145;
wire wire2151;
wire wire2156;
wire wire2160;
wire wire2162;
wire wire2172;
wire wire2181;
wire wire2185;
wire wire2186;
wire wire2189;
wire wire2190;
wire wire2195;
wire wire2196;
wire wire2197;
wire wire2200;
wire wire2201;
wire wire2202;
wire wire2203;
wire wire2204;
wire wire2207;
wire wire2208;
wire wire2209;
wire wire2210;
wire wire2211;
wire wire2235;
wire wire2236;
wire wire2238;
wire wire2239;
wire wire2244;
wire wire2247;
wire wire2248;
wire wire2249;
wire wire2250;
wire wire2251;
wire wire2252;
wire wire2253;
wire wire2254;
wire wire2255;
wire wire2256;
wire wire2257;
wire wire2258;
wire wire2259;
wire wire2260;
wire wire2261;
wire wire2262;
wire wire2263;
wire wire2264;
wire wire2265;
wire wire2266;
wire wire2267;
wire wire2268;
wire wire2269;
wire wire2270;
wire wire2271;
wire wire2272;
wire wire2273;
wire wire2274;
wire wire2275;
wire wire2276;
wire wire2277;
wire wire2278;
wire wire2279;
wire wire2280;
wire wire2281;
wire wire2282;
wire wire2283;
wire wire2284;
wire wire2285;
wire wire2286;
wire wire2287;
wire wire2288;
wire wire2289;
wire wire2290;
wire wire2291;
wire wire2292;
wire wire2293;
wire wire2294;
wire wire2295;
wire wire2296;
wire wire2297;
wire wire2298;
wire wire2299;
wire wire2300;
wire wire2301;
wire wire2302;
wire wire2303;
wire wire2304;
wire wire2305;
wire wire2306;
wire wire2307;
wire wire2308;
wire wire2309;
wire wire6930;
wire wire6933;
wire wire6936;
wire wire6939;
wire wire6942;
wire wire6945;
wire wire6948;
wire wire6951;
wire wire6954;
wire wire6957;
wire wire6960;
wire wire6963;
wire wire6964;
wire wire6965;
wire wire6966;
wire wire6967;
wire wire6968;
wire wire6969;
wire wire6973;
wire wire6974;
wire wire6975;
wire wire6976;
wire wire6977;
wire wire6989;
wire wire6990;
wire wire6993;
wire wire6994;
wire wire6995;
wire wire6996;
wire wire6997;
wire wire6999;
wire wire7000;
wire wire7002;
wire wire7003;
wire wire7004;
wire wire7005;
wire wire7007;
wire wire7008;
wire wire7009;
wire wire7010;
wire wire7011;
wire wire7012;
wire wire7013;
wire wire7017;
wire wire7018;
wire wire7020;
wire wire7021;
wire wire7026;
wire wire7027;
wire wire7028;
wire wire7031;
wire wire7032;
wire wire7034;
wire wire7035;
wire wire7040;
wire wire7041;
wire wire7042;
wire wire7045;
wire wire7046;
wire wire7048;
wire wire7049;
wire wire7054;
wire wire7055;
wire wire7056;
wire wire7059;
wire wire7060;
wire wire7062;
wire wire7063;
wire wire7068;
wire wire7069;
wire wire7070;
wire wire7073;
wire wire7074;
wire wire7076;
wire wire7077;
wire wire7082;
wire wire7083;
wire wire7084;
wire wire7087;
wire wire7088;
wire wire7090;
wire wire7091;
wire wire7096;
wire wire7097;
wire wire7098;
wire wire7102;
wire wire7104;
wire wire7107;
wire wire7108;
wire wire7109;
wire wire7110;
wire wire7112;
wire wire7113;
wire wire7118;
wire wire7119;
wire wire7120;
wire wire7125;
wire wire7126;
wire wire7128;
wire wire7129;
wire wire7130;
wire wire7132;
wire wire7133;
wire wire7135;
wire wire7136;
wire wire7141;
wire wire7142;
wire wire7143;
wire wire7149;
wire wire7152;
wire wire7155;
wire wire7158;
wire wire7164;
wire wire7167;
wire wire7170;
wire wire7173;
wire wire7175;
wire wire7183;
wire wire7184;
wire wire7186;
wire wire7189;
wire wire7190;
wire wire7191;
wire wire7192;
wire wire7196;
wire wire7197;
wire wire7198;
wire wire7201;
wire wire7203;
wire wire7205;
wire wire7207;
wire wire7209;
wire wire7219;
wire wire7220;
wire wire7221;
wire wire7223;
wire wire7224;
wire wire7225;
wire wire7226;
wire wire7227;
wire wire7228;
wire wire7229;
wire wire7230;
wire wire7231;
wire wire7232;
wire wire7233;
wire wire7234;
wire wire7236;
wire wire7239;
wire wire7240;
wire wire7241;
wire wire7243;
wire wire7244;
wire wire7245;
wire wire7246;
wire wire7247;
wire wire7248;
wire wire7250;
wire wire7251;
wire wire7252;
wire wire7257;
wire wire7263;
wire wire7270;
wire wire7271;
wire wire7272;
wire wire7273;
wire wire7274;
wire wire7275;
wire wire7279;
wire wire7280;
wire wire7282;
wire wire7283;
wire wire7288;
wire wire7289;
wire wire7290;
wire wire7294;
wire wire7302;
wire wire7304;
wire wire7307;
wire wire7308;
wire wire7310;
wire wire7311;
wire wire7316;
wire wire7317;
wire wire7318;
wire wire7322;
wire wire7324;
wire wire7326;
wire wire7328;
wire wire7333;
wire wire7334;
wire wire7335;
wire wire7336;
wire wire7347;
wire wire7354;
wire wire7360;
wire wire7361;
wire wire7364;
wire wire7365;
wire wire7368;
wire wire7370;
wire wire7372;
wire wire7373;
wire wire7375;
wire wire7381;
wire wire7384;
wire wire7387;
wire wire7389;
wire wire7405;
wire wire7407;
wire wire7408;
wire wire7409;
wire wire7410;
wire wire7411;
wire wire7412;
wire wire7414;
wire wire7415;
wire wire7416;
wire wire7417;
wire wire7418;
wire wire7419;
wire wire7423;
wire wire7424;
wire wire7425;
wire wire7426;
wire wire7427;
wire wire7428;
wire wire7429;
wire wire7430;
wire wire7431;
wire wire7432;
wire wire7433;
wire wire7436;
wire wire7437;
wire wire7438;
wire wire7439;
wire wire7440;
wire wire7441;
wire wire7442;
wire wire7443;
wire wire7447;
wire wire7449;
wire wire7451;
wire wire7454;
wire wire7455;
wire wire7456;
wire wire7462;
wire wire7467;
wire wire7468;
wire wire7472;
wire wire7478;
wire wire7483;
wire wire7486;
wire wire7495;
wire wire7500;
wire wire7501;
wire wire7502;
wire wire7506;
wire wire7508;
wire wire7511;
wire wire7512;
wire wire7518;
wire wire7520;
wire wire7521;
wire wire7524;
wire wire7525;
wire wire7526;
wire wire7527;
wire wire7529;
wire wire7532;
wire wire7533;
wire wire7534;
wire wire7535;
wire wire7537;
wire wire7539;
reg n_n3033;

reg n_n2960;

reg n_n3175;

reg n_n3871;

reg n_n3420;

reg n_n3489;

reg n_n4171;

reg n_n4116;

reg n_n2971;

reg n_n3700;

reg n_n4057;

reg n_n4206;

reg n_n3074;

reg n_n3791;

reg n_n4194;

reg n_n3139;

reg n_n4099;

reg n_n3715;

reg n_n3832;

reg n_n3949;

reg n_n3500;

reg n_n3957;

reg ndn3_8;

reg n_n4220;

reg n_n3300;

reg n_n3778;

reg nen5_9;

reg n_n3354;

reg n_n3157;

reg n_n3071;

reg n_n3535;

reg n_n3761;

reg n_n3516;

reg ndn5_16;

reg n_n4149;

reg n_n3870;

reg n_n3805;

reg n_n3011;

reg n_n3709;

reg n_n3184;

reg n_n3574;

reg n_n3822;

reg n_n4072;

reg n_n3262;

reg n_n4039;

reg n_n3482;

reg n_n3908;

reg n_n3164;

reg n_n3517;

reg n_n3585;

reg n_n3928;

reg n_n4182;

reg ndn5_4;

reg n_n2991;

reg n_n3745;

reg n_n3691;

reg n_n3019;

reg n_n4180;

reg n_n4133;

reg n_n3567;

reg n_n3799;

reg n_n3235;

reg n_n3751;

reg nlc1_2;

reg n_n3060;

reg n_n3575;

reg n_n4242;

reg n_n3031;

reg n_n3813;

reg n_n3882;

reg n_n3838;

reg n_n3280;

reg n_n3750;

reg n_n3221;

reg n_n3369;

reg n_n3331;

reg n_n3128;

reg n_n3999;

reg n_n3797;

reg ndn5_3;

reg n_n3973;

reg n_n3151;

reg n_n3815;

reg n_n3808;

reg n_n3248;

reg n_n4117;

reg n_n3922;

reg n_n3844;

reg n_n3810;

reg n_n3736;

reg n_n3170;

reg n_n3346;

reg n_n3324;

reg n_n3312;

reg n_n3796;

reg n_n4114;

reg n_n3821;

reg n_n3344;

reg n_n4239;

reg n_n3304;

reg n_n3875;

reg n_n3741;

reg n_n3203;

reg n_n4193;

reg n_n4223;

reg n_n3651;

reg n_n3047;

reg ndn5_9;

reg n_n3924;

reg n_n3923;

reg n_n4083;

reg pnext_0_0_;

reg n_n3677;

reg nak5_2;

reg n_n4064;

reg n_n3529;

reg n_n3988;

reg n_n3293;

reg n_n3469;

reg pover_0_0_;

reg n_n4004;

reg n_n3179;

reg n_n4070;

reg ndn5_6;

reg n_n3713;

reg n_n4054;

reg n_n3311;

reg n_n3841;

reg n_n4212;

reg n_n4165;

reg n_n4159;

reg n_n4243;

reg n_n3578;

reg n_n3381;

reg n_n3634;

reg n_n4093;

reg n_n4224;

reg n_n4090;

reg n_n4179;

reg n_n3214;

reg ndn5_7;

reg n_n4056;

reg n_n3062;

reg n_n3540;

reg n_n4230;

reg n_n3733;

reg n_n3246;

reg n_n3919;

reg n_n3433;

reg n_n3711;

reg n_n3356;

reg n_n3013;

reg n_n3398;

reg n_n3212;

reg n_n3864;

reg n_n4030;

reg n_n3513;

reg n_n4086;

reg n_n3774;

reg n_n3610;

reg n_n3480;

reg n_n3659;

reg n_n3931;

reg n_n3996;

reg n_n2986;

reg n_n4135;

reg ndn5_5;

reg n_n3684;

reg n_n4071;

reg n_n4232;

reg ndn3_11;

reg n_n3679;

reg n_n3625;

reg n_n3940;

reg n_n3947;

reg n_n3776;

reg n_n4158;

reg n_n3182;

reg n_n3384;

reg n_n4259;

reg n_n4140;

reg n_n3855;

reg ndn3_3;

reg n_n4014;

reg n_n3649;

reg n_n3065;

reg n_n4246;

reg n_n3890;

reg n_n3340;

reg n_n3921;

reg n_n3509;

reg n_n3868;

reg n_n3387;

reg n_n3918;

reg n_n3457;

reg n_n4036;

reg n_n4136;

reg ndn2_2;

reg n_n4042;

reg n_n4176;

reg n_n4120;

reg n_n3159;

reg n_n3250;

reg n_n4018;

reg n_n3965;

reg n_n4021;

reg n_n3767;

reg n_n3000;

reg n_n3910;

reg n_n3728;

reg n_n4111;

reg pdn;

reg n_n4027;

reg n_n3698;

reg n_n4106;

reg n_n4095;

reg n_n3498;

reg n_n3694;

reg n_n3309;

reg n_n4197;

reg n_n3971;

reg n_n3626;

reg n_n3932;

reg nlak3_9;

reg n_n3044;

reg n_n4222;

reg n_n3630;

reg n_n3680;

reg n_n4079;

reg ndn1_4;

reg n_n3205;

reg n_n3100;

reg n_n3188;

reg n_n4177;

reg n_n3327;

reg n_n3818;

reg n_n3143;

reg n_n3843;

reg n_n3069;

reg n_n3842;

reg n_n4145;

reg n_n3628;

reg n_n3716;

reg n_n2995;

reg nlak3_2;

reg n_n3430;

reg n_n3373;

reg n_n3916;

reg n_n3453;

reg n_n3448;

reg n_n4134;

reg n_n3800;

reg n_n3473;

reg n_n3612;

reg n_n4075;

reg n_n3912;

reg n_n3905;

reg ngfdn_3;

reg n_n3961;

reg n_n4236;

reg n_n3424;

reg n_n3081;

reg n_n4208;

reg nld3_9;

reg n_n4073;

reg n_n3345;

reg n_n3375;

reg n_n3426;

reg n_n4221;

reg n_n3105;

reg n_n3807;

reg n_n3196;

reg n_n3283;

reg n_n3840;

reg n_n3771;

reg n_n3906;

reg n_n4080;

reg n_n3743;

reg n_n3606;

reg n_n3901;

reg n_n3866;

reg n_n4167;

reg n_n4205;

reg n_n3024;

reg n_n3445;

reg n_n3862;

reg n_n3974;

reg n_n3887;

reg n_n3336;

reg n_n3199;

reg n_n3470;

reg n_n3541;

reg n_n3824;

reg ndn5_2;

reg ndn5_8;

reg n_n4119;

reg n_n3788;

reg n_n4118;

reg n_n3464;

reg n_n3442;

reg n_n3722;

reg n_n3806;

reg n_n3786;

reg n_n4126;

reg n_n3563;

reg n_n4024;

reg n_n3735;

reg n_n3122;

reg n_n3622;

reg n_n3646;

reg n_n3294;

reg n_n4015;

reg n_n3793;

reg n_n4218;

reg n_n3417;

reg n_n3689;

reg n_n3323;

reg n_n3794;

reg n_n4045;

reg n_n3436;

reg n_n3968;

reg n_n3533;

reg n_n3884;

reg n_n3393;

reg n_n3067;

reg n_n2968;

reg n_n3708;

reg n_n4132;

reg n_n3826;

reg n_n3872;

reg n_n3580;

reg n_n3493;

reg n_n3981;

reg n_n4227;

reg n_n3992;

reg ndn5_10;

reg n_n3681;

reg n_n3701;

reg n_n3876;

reg n_n3002;

reg n_n3388;

reg n_n2982;

reg n_n3851;

reg n_n4214;

reg n_n2989;

reg n_n4181;

reg n_n3939;

reg n_n4237;

reg n_n3274;

reg n_n3607;

reg n_n3663;

reg n_n3468;

reg n_n4252;

reg n_n4183;

reg n_n3303;

reg n_n3367;

reg n_n3959;

reg n_n4047;

reg n_n4209;

reg n_n4068;

reg n_n3475;

reg n_n4060;

reg n_n3998;

reg nsr5_4;

reg n_n3829;

reg n_n3554;

reg nsr3_9;

reg n_n3755;

reg n_n3556;

reg nsr5_5;

reg nsr5_3;

reg nsr5_2;

reg nsr5_7;

reg n_n3462;

reg nsr3_2;

reg nsr5_8;

reg n_n3460;

always  @(posedge pclk)
	n_n3033<=n_n3032;

 always  @(posedge pclk)
	n_n2960<=n_n2959;

 always  @(posedge pclk)
	n_n3175<=n_n3174;

 always  @(posedge pclk)
	n_n3871<=n_n2952;

 always  @(posedge pclk)
	n_n3420<=n_n2973;

 always  @(posedge pclk)
	n_n3489<=n_n3488;

 always  @(posedge pclk)
	n_n4171<=n_n3596;

 always  @(posedge pclk)
	n_n4116<=n_n3969;

 always  @(posedge pclk)
	n_n2971<=n_n2970;

 always  @(posedge pclk)
	n_n3700<=n_n3259;

 always  @(posedge pclk)
	n_n4057<=n_n4007;

 always  @(posedge pclk)
	n_n4206<=n_n3483;

 always  @(posedge pclk)
	n_n3074<=n_n3073;

 always  @(posedge pclk)
	n_n3791<=n_n3653;

 always  @(posedge pclk)
	n_n4194<=n_n3051;

 always  @(posedge pclk)
	n_n3139<=n_n3137;

 always  @(posedge pclk)
	n_n4099<=n_n4098;

 always  @(posedge pclk)
	n_n3715<=n_n3007;

 always  @(posedge pclk)
	n_n3832<=n_n3086;

 always  @(posedge pclk)
	n_n3949<=n_n3602;

 always  @(posedge pclk)
	n_n3500<=n_n3499;

 always  @(posedge pclk)
	n_n3957<=n_n3956;

 always  @(posedge pclk)
	ndn3_8<=n_n3752;

 always  @(posedge pclk)
	n_n4220<=n_n3941;

 always  @(posedge pclk)
	n_n3300<=n_n3299;

 always  @(posedge pclk)
	n_n3778<=n_n3284;

 always  @(posedge pclk)
	nen5_9<=n_n3618;

 always  @(posedge pclk)
	n_n3354<=n_n3353;

 always  @(posedge pclk)
	n_n3157<=n_n2972;

 always  @(posedge pclk)
	n_n3071<=n_n3070;

 always  @(posedge pclk)
	n_n3535<=n_n3454;

 always  @(posedge pclk)
	n_n3761<=n_n3640;

 always  @(posedge pclk)
	n_n3516<=n_n2992;

 always  @(posedge pclk)
	ndn5_16<=n_n3063;

 always  @(posedge pclk)
	n_n4149<=n_n4147;

 always  @(posedge pclk)
	n_n3870<=n_n3772;

 always  @(posedge pclk)
	n_n3805<=n_n3132;

 always  @(posedge pclk)
	n_n3011<=n_n2969;

 always  @(posedge pclk)
	n_n3709<=n_n3616;

 always  @(posedge pclk)
	n_n3184<=n_n3183;

 always  @(posedge pclk)
	n_n3574<=n_n3523;

 always  @(posedge pclk)
	n_n3822<=n_n3004;

 always  @(posedge pclk)
	n_n4072<=n_n3206;

 always  @(posedge pclk)
	n_n3262<=n_n2984;

 always  @(posedge pclk)
	n_n4039<=n_n4038;

 always  @(posedge pclk)
	n_n3482<=n_n3481;

 always  @(posedge pclk)
	n_n3908<=n_n3322;

 always  @(posedge pclk)
	n_n3164<=n_n3144;

 always  @(posedge pclk)
	n_n3517<=n_n3401;

 always  @(posedge pclk)
	n_n3585<=n_n3584;

 always  @(posedge pclk)
	n_n3928<=n_n3926;

 always  @(posedge pclk)
	n_n4182<=n_n2958;

 always  @(posedge pclk)
	ndn5_4<=n_n3739;

 always  @(posedge pclk)
	n_n2991<=n_n2990;

 always  @(posedge pclk)
	n_n3745<=n_n3744;

 always  @(posedge pclk)
	n_n3691<=n_n3690;

 always  @(posedge pclk)
	n_n3019<=n_n3018;

 always  @(posedge pclk)
	n_n4180<=n_n3334;

 always  @(posedge pclk)
	n_n4133<=n_n2997;

 always  @(posedge pclk)
	n_n3567<=n_n3566;

 always  @(posedge pclk)
	n_n3799<=n_n3798;

 always  @(posedge pclk)
	n_n3235<=n_n2974;

 always  @(posedge pclk)
	n_n3751<=n_n3115;

 always  @(posedge pclk)
	nlc1_2<=n_n3811;

 always  @(posedge pclk)
	n_n3060<=n_n3059;

 always  @(posedge pclk)
	n_n3575<=n_n3325;

 always  @(posedge pclk)
	n_n4242<=n_n3052;

 always  @(posedge pclk)
	n_n3031<=n_n3030;

 always  @(posedge pclk)
	n_n3813<=n_n3153;

 always  @(posedge pclk)
	n_n3882<=n_n3705;

 always  @(posedge pclk)
	n_n3838<=n_n3432;

 always  @(posedge pclk)
	n_n3280<=n_n2983;

 always  @(posedge pclk)
	n_n3750<=n_n3040;

 always  @(posedge pclk)
	n_n3221<=n_n3209;

 always  @(posedge pclk)
	n_n3369<=n_n3165;

 always  @(posedge pclk)
	n_n3331<=n_n3057;

 always  @(posedge pclk)
	n_n3128<=n_n3127;

 always  @(posedge pclk)
	n_n3999<=n_n4254;

 always  @(posedge pclk)
	n_n3797<=n_n3163;

 always  @(posedge pclk)
	ndn5_3<=n_n3041;

 always  @(posedge pclk)
	n_n3973<=n_n3972;

 always  @(posedge pclk)
	n_n3151<=n_n3150;

 always  @(posedge pclk)
	n_n3815<=n_n3814;

 always  @(posedge pclk)
	n_n3808<=n_n3349;

 always  @(posedge pclk)
	n_n3248<=n_n3247;

 always  @(posedge pclk)
	n_n4117<=n_n3661;

 always  @(posedge pclk)
	n_n3922<=n_n3652;

 always  @(posedge pclk)
	n_n3844<=n_n3315;

 always  @(posedge pclk)
	n_n3810<=n_n3316;

 always  @(posedge pclk)
	n_n3736<=n_n3456;

 always  @(posedge pclk)
	n_n3170<=n_n3168;

 always  @(posedge pclk)
	n_n3346<=n_n3037;

 always  @(posedge pclk)
	n_n3324<=n_n3119;

 always  @(posedge pclk)
	n_n3312<=n_n2966;

 always  @(posedge pclk)
	n_n3796<=n_n3795;

 always  @(posedge pclk)
	n_n4114<=n_n4113;

 always  @(posedge pclk)
	n_n3821<=n_n3014;

 always  @(posedge pclk)
	n_n3344<=n_n3103;

 always  @(posedge pclk)
	n_n4239<=n_n4238;

 always  @(posedge pclk)
	n_n3304<=n_n3210;

 always  @(posedge pclk)
	n_n3875<=n_n3113;

 always  @(posedge pclk)
	n_n3741<=n_n3740;

 always  @(posedge pclk)
	n_n3203<=n_n3202;

 always  @(posedge pclk)
	n_n4193<=n_n3720;

 always  @(posedge pclk)
	n_n4223<=n_n3314;

 always  @(posedge pclk)
	n_n3651<=n_n3650;

 always  @(posedge pclk)
	n_n3047<=n_n3046;

 always  @(posedge pclk)
	ndn5_9<=n_n3458;

 always  @(posedge pclk)
	n_n3924<=n_n3409;

 always  @(posedge pclk)
	n_n3923<=n_n3227;

 always  @(posedge pclk)
	n_n4083<=n_n2963;

 always  @(posedge pclk)
	pnext_0_0_<=n_n3005;

 always  @(posedge pclk)
	n_n3677<=n_n2998;

 always  @(posedge pclk)
	nak5_2<=n_n3638;

 always  @(posedge pclk)
	n_n4064<=n_n4063;

 always  @(posedge pclk)
	n_n3529<=n_n3240;

 always  @(posedge pclk)
	n_n3988<=n_n3987;

 always  @(posedge pclk)
	n_n3293<=n_n3177;

 always  @(posedge pclk)
	n_n3469<=n_n2996;

 always  @(posedge pclk)
	pover_0_0_<=n_n3061;

 always  @(posedge pclk)
	n_n4004<=n_n3091;

 always  @(posedge pclk)
	n_n3179<=n_n3178;

 always  @(posedge pclk)
	n_n4070<=n_n3193;

 always  @(posedge pclk)
	ndn5_6<=n_n3016;

 always  @(posedge pclk)
	n_n3713<=n_n3712;

 always  @(posedge pclk)
	n_n4054<=n_n4053;

 always  @(posedge pclk)
	n_n3311<=n_n3310;

 always  @(posedge pclk)
	n_n3841<=n_n3431;

 always  @(posedge pclk)
	n_n4212<=n_n3599;

 always  @(posedge pclk)
	n_n4165<=n_n3146;

 always  @(posedge pclk)
	n_n4159<=n_n3058;

 always  @(posedge pclk)
	n_n4243<=n_n3914;

 always  @(posedge pclk)
	n_n3578<=n_n3389;

 always  @(posedge pclk)
	n_n3381<=n_n3379;

 always  @(posedge pclk)
	n_n3634<=n_n3633;

 always  @(posedge pclk)
	n_n4093<=n_n3147;

 always  @(posedge pclk)
	n_n4224<=n_n3586;

 always  @(posedge pclk)
	n_n4090<=n_n4089;

 always  @(posedge pclk)
	n_n4179<=n_n3963;

 always  @(posedge pclk)
	n_n3214<=n_n3213;

 always  @(posedge pclk)
	ndn5_7<=n_n3538;

 always  @(posedge pclk)
	n_n4056<=n_n4055;

 always  @(posedge pclk)
	n_n3062<=n_n3009;

 always  @(posedge pclk)
	n_n3540<=n_n3050;

 always  @(posedge pclk)
	n_n4230<=n_n4229;

 always  @(posedge pclk)
	n_n3733<=n_n3595;

 always  @(posedge pclk)
	n_n3246<=n_n3245;

 always  @(posedge pclk)
	n_n3919<=n_n2955;

 always  @(posedge pclk)
	n_n3433<=n_n3172;

 always  @(posedge pclk)
	n_n3711<=n_n3710;

 always  @(posedge pclk)
	n_n3356<=n_n2979;

 always  @(posedge pclk)
	n_n3013<=n_n3012;

 always  @(posedge pclk)
	n_n3398<=n_n3397;

 always  @(posedge pclk)
	n_n3212<=n_n3211;

 always  @(posedge pclk)
	n_n3864<=n_n3863;

 always  @(posedge pclk)
	n_n4030<=n_n4029;

 always  @(posedge pclk)
	n_n3513<=n_n3487;

 always  @(posedge pclk)
	n_n4086<=n_n4085;

 always  @(posedge pclk)
	n_n3774<=n_n3664;

 always  @(posedge pclk)
	n_n3610<=n_n3609;

 always  @(posedge pclk)
	n_n3480<=n_n3266;

 always  @(posedge pclk)
	n_n3659<=n_n3658;

 always  @(posedge pclk)
	n_n3931<=n_n3244;

 always  @(posedge pclk)
	n_n3996<=n_n3200;

 always  @(posedge pclk)
	n_n2986<=n_n2985;

 always  @(posedge pclk)
	n_n4135<=n_n2957;

 always  @(posedge pclk)
	ndn5_5<=n_n3348;

 always  @(posedge pclk)
	n_n3684<=n_n3683;

 always  @(posedge pclk)
	n_n4071<=n_n3615;

 always  @(posedge pclk)
	n_n4232<=n_n4231;

 always  @(posedge pclk)
	ndn3_11<=n_n3287;

 always  @(posedge pclk)
	n_n3679<=n_n3049;

 always  @(posedge pclk)
	n_n3625<=n_n3558;

 always  @(posedge pclk)
	n_n3940<=n_n3263;

 always  @(posedge pclk)
	n_n3947<=n_n3946;

 always  @(posedge pclk)
	n_n3776<=n_n3614;

 always  @(posedge pclk)
	n_n4158<=n_n3437;

 always  @(posedge pclk)
	n_n3182<=n_n3180;

 always  @(posedge pclk)
	n_n3384<=n_n2978;

 always  @(posedge pclk)
	n_n4259<=n_n4256;

 always  @(posedge pclk)
	n_n4140<=n_n4139;

 always  @(posedge pclk)
	n_n3855<=n_n3853;

 always  @(posedge pclk)
	ndn3_3<=n_n3530;

 always  @(posedge pclk)
	n_n4014<=n_n4011;

 always  @(posedge pclk)
	n_n3649<=n_n3648;

 always  @(posedge pclk)
	n_n3065<=n_n3064;

 always  @(posedge pclk)
	n_n4246<=n_n3276;

 always  @(posedge pclk)
	n_n3890<=n_n3570;

 always  @(posedge pclk)
	n_n3340<=n_n3339;

 always  @(posedge pclk)
	n_n3921<=n_n3524;

 always  @(posedge pclk)
	n_n3509<=n_n3241;

 always  @(posedge pclk)
	n_n3868<=n_n2956;

 always  @(posedge pclk)
	n_n3387<=n_n3145;

 always  @(posedge pclk)
	n_n3918<=n_n3592;

 always  @(posedge pclk)
	n_n3457<=n_n3102;

 always  @(posedge pclk)
	n_n4036<=n_n3093;

 always  @(posedge pclk)
	n_n4136<=n_n3191;

 always  @(posedge pclk)
	ndn2_2<=n_n3476;

 always  @(posedge pclk)
	n_n4042<=n_n4041;

 always  @(posedge pclk)
	n_n4176<=n_n3479;

 always  @(posedge pclk)
	n_n4120<=n_n3895;

 always  @(posedge pclk)
	n_n3159<=n_n3158;

 always  @(posedge pclk)
	n_n3250<=n_n3249;

 always  @(posedge pclk)
	n_n4018<=n_n3717;

 always  @(posedge pclk)
	n_n3965<=n_n3106;

 always  @(posedge pclk)
	n_n4021<=n_n4020;

 always  @(posedge pclk)
	n_n3767<=n_n3765;

 always  @(posedge pclk)
	n_n3000<=n_n2999;

 always  @(posedge pclk)
	n_n3910<=n_n3909;

 always  @(posedge pclk)
	n_n3728<=n_n3726;

 always  @(posedge pclk)
	n_n4111<=n_n4110;

 always  @(posedge pclk)
	pdn<=n_n3620;

 always  @(posedge pclk)
	n_n4027<=n_n2980;

 always  @(posedge pclk)
	n_n3698<=n_n3696;

 always  @(posedge pclk)
	n_n4106<=n_n4105;

 always  @(posedge pclk)
	n_n4095<=n_n4094;

 always  @(posedge pclk)
	n_n3498<=n_n3497;

 always  @(posedge pclk)
	n_n3694<=n_n3692;

 always  @(posedge pclk)
	n_n3309<=n_n3308;

 always  @(posedge pclk)
	n_n4197<=n_n3847;

 always  @(posedge pclk)
	n_n3971<=n_n3801;

 always  @(posedge pclk)
	n_n3626<=n_n3162;

 always  @(posedge pclk)
	n_n3932<=n_n3189;

 always  @(posedge pclk)
	nlak3_9<=n_n3465;

 always  @(posedge pclk)
	n_n3044<=n_n3043;

 always  @(posedge pclk)
	n_n4222<=n_n4174;

 always  @(posedge pclk)
	n_n3630<=n_n2976;

 always  @(posedge pclk)
	n_n3680<=n_n3008;

 always  @(posedge pclk)
	n_n4079<=n_n4032;

 always  @(posedge pclk)
	ndn1_4<=n_n3305;

 always  @(posedge pclk)
	n_n3205<=n_n3204;

 always  @(posedge pclk)
	n_n3100<=n_n3028;

 always  @(posedge pclk)
	n_n3188<=n_n3075;

 always  @(posedge pclk)
	n_n4177<=n_n3087;

 always  @(posedge pclk)
	n_n3327<=n_n3326;

 always  @(posedge pclk)
	n_n3818<=n_n3817;

 always  @(posedge pclk)
	n_n3143<=n_n3136;

 always  @(posedge pclk)
	n_n3843<=n_n3668;

 always  @(posedge pclk)
	n_n3069<=n_n3068;

 always  @(posedge pclk)
	n_n3842<=n_n3413;

 always  @(posedge pclk)
	n_n4145<=n_n3222;

 always  @(posedge pclk)
	n_n3628<=n_n3627;

 always  @(posedge pclk)
	n_n3716<=n_n3399;

 always  @(posedge pclk)
	n_n2995<=n_n2994;

 always  @(posedge pclk)
	nlak3_2<=n_n2987;

 always  @(posedge pclk)
	n_n3430<=n_n3429;

 always  @(posedge pclk)
	n_n3373<=n_n3372;

 always  @(posedge pclk)
	n_n3916<=n_n3915;

 always  @(posedge pclk)
	n_n3453<=n_n3452;

 always  @(posedge pclk)
	n_n3448<=n_n3447;

 always  @(posedge pclk)
	n_n4134<=n_n3156;

 always  @(posedge pclk)
	n_n3800<=n_n3201;

 always  @(posedge pclk)
	n_n3473<=n_n3472;

 always  @(posedge pclk)
	n_n3612<=n_n3611;

 always  @(posedge pclk)
	n_n4075<=n_n4074;

 always  @(posedge pclk)
	n_n3912<=n_n3449;

 always  @(posedge pclk)
	n_n3905<=n_n3904;

 always  @(posedge pclk)
	ngfdn_3<=n_n3542;

 always  @(posedge pclk)
	n_n3961<=n_n2964;

 always  @(posedge pclk)
	n_n4236<=n_n4028;

 always  @(posedge pclk)
	n_n3424<=n_n3423;

 always  @(posedge pclk)
	n_n3081<=n_n2977;

 always  @(posedge pclk)
	n_n4208<=n_n3130;

 always  @(posedge pclk)
	nld3_9<=n_n3042;

 always  @(posedge pclk)
	n_n4073<=n_n3338;

 always  @(posedge pclk)
	n_n3345<=n_n3078;

 always  @(posedge pclk)
	n_n3375<=n_n3374;

 always  @(posedge pclk)
	n_n3426<=n_n3425;

 always  @(posedge pclk)
	n_n4221<=n_n3486;

 always  @(posedge pclk)
	n_n3105<=n_n3104;

 always  @(posedge pclk)
	n_n3807<=n_n3129;

 always  @(posedge pclk)
	n_n3196<=n_n3152;

 always  @(posedge pclk)
	n_n3283<=n_n3053;

 always  @(posedge pclk)
	n_n3840<=n_n3133;

 always  @(posedge pclk)
	n_n3771<=n_n3770;

 always  @(posedge pclk)
	n_n3906<=n_n3003;

 always  @(posedge pclk)
	n_n4080<=n_n3010;

 always  @(posedge pclk)
	n_n3743<=n_n3666;

 always  @(posedge pclk)
	n_n3606<=n_n3605;

 always  @(posedge pclk)
	n_n3901<=n_n3899;

 always  @(posedge pclk)
	n_n3866<=n_n2961;

 always  @(posedge pclk)
	n_n4167<=n_n4166;

 always  @(posedge pclk)
	n_n4205<=n_n3511;

 always  @(posedge pclk)
	n_n3024<=n_n3022;

 always  @(posedge pclk)
	n_n3445<=n_n3155;

 always  @(posedge pclk)
	n_n3862<=n_n3117;

 always  @(posedge pclk)
	n_n3974<=n_n3027;

 always  @(posedge pclk)
	n_n3887<=n_n3885;

 always  @(posedge pclk)
	n_n3336<=n_n3335;

 always  @(posedge pclk)
	n_n3199<=n_n3197;

 always  @(posedge pclk)
	n_n3470<=n_n3034;

 always  @(posedge pclk)
	n_n3541<=n_n2962;

 always  @(posedge pclk)
	n_n3824<=n_n3823;

 always  @(posedge pclk)
	ndn5_2<=n_n3160;

 always  @(posedge pclk)
	ndn5_8<=n_n3029;

 always  @(posedge pclk)
	n_n4119<=n_n3406;

 always  @(posedge pclk)
	n_n3788<=n_n3787;

 always  @(posedge pclk)
	n_n4118<=n_n3506;

 always  @(posedge pclk)
	n_n3464<=n_n3216;

 always  @(posedge pclk)
	n_n3442<=n_n3215;

 always  @(posedge pclk)
	n_n3722<=n_n3721;

 always  @(posedge pclk)
	n_n3806<=n_n3173;

 always  @(posedge pclk)
	n_n3786<=n_n3785;

 always  @(posedge pclk)
	n_n4126<=n_n3277;

 always  @(posedge pclk)
	n_n3563<=n_n3562;

 always  @(posedge pclk)
	n_n4024<=n_n4023;

 always  @(posedge pclk)
	n_n3735<=n_n3015;

 always  @(posedge pclk)
	n_n3122<=n_n3120;

 always  @(posedge pclk)
	n_n3622<=n_n3621;

 always  @(posedge pclk)
	n_n3646<=n_n3645;

 always  @(posedge pclk)
	n_n3294<=n_n2965;

 always  @(posedge pclk)
	n_n4015<=n_n3913;

 always  @(posedge pclk)
	n_n3793<=n_n3695;

 always  @(posedge pclk)
	n_n4218<=n_n4217;

 always  @(posedge pclk)
	n_n3417<=n_n3416;

 always  @(posedge pclk)
	n_n3689<=n_n3687;

 always  @(posedge pclk)
	n_n3323<=n_n3320;

 always  @(posedge pclk)
	n_n3794<=n_n3559;

 always  @(posedge pclk)
	n_n4045<=n_n4044;

 always  @(posedge pclk)
	n_n3436<=n_n3435;

 always  @(posedge pclk)
	n_n3968<=n_n3967;

 always  @(posedge pclk)
	n_n3533<=n_n3352;

 always  @(posedge pclk)
	n_n3884<=n_n3321;

 always  @(posedge pclk)
	n_n3393<=n_n3318;

 always  @(posedge pclk)
	n_n3067<=n_n3066;

 always  @(posedge pclk)
	n_n2968<=n_n2967;

 always  @(posedge pclk)
	n_n3708<=n_n3707;

 always  @(posedge pclk)
	n_n4132<=n_n3194;

 always  @(posedge pclk)
	n_n3826<=n_n3825;

 always  @(posedge pclk)
	n_n3872<=n_n3123;

 always  @(posedge pclk)
	n_n3580<=n_n3579;

 always  @(posedge pclk)
	n_n3493<=n_n3491;

 always  @(posedge pclk)
	n_n3981<=n_n3980;

 always  @(posedge pclk)
	n_n4227<=n_n3859;

 always  @(posedge pclk)
	n_n3992<=n_n3723;

 always  @(posedge pclk)
	ndn5_10<=n_n3231;

 always  @(posedge pclk)
	n_n3681<=n_n3400;

 always  @(posedge pclk)
	n_n3701<=n_n3048;

 always  @(posedge pclk)
	n_n3876<=n_n3804;

 always  @(posedge pclk)
	n_n3002<=n_n3001;

 always  @(posedge pclk)
	n_n3388<=n_n2953;

 always  @(posedge pclk)
	n_n2982<=n_n2981;

 always  @(posedge pclk)
	n_n3851<=n_n3850;

 always  @(posedge pclk)
	n_n4214<=n_n3332;

 always  @(posedge pclk)
	n_n2989<=n_n2988;

 always  @(posedge pclk)
	n_n4181<=n_n3390;

 always  @(posedge pclk)
	n_n3939<=n_n3589;

 always  @(posedge pclk)
	n_n4237<=n_n3192;

 always  @(posedge pclk)
	n_n3274<=n_n3273;

 always  @(posedge pclk)
	n_n3607<=n_n2975;

 always  @(posedge pclk)
	n_n3663<=n_n3662;

 always  @(posedge pclk)
	n_n3468<=n_n3038;

 always  @(posedge pclk)
	n_n4252<=n_n3671;

 always  @(posedge pclk)
	n_n4183<=n_n3190;

 always  @(posedge pclk)
	n_n3303<=n_n3101;

 always  @(posedge pclk)
	n_n3367<=n_n3366;

 always  @(posedge pclk)
	n_n3959<=n_n3958;

 always  @(posedge pclk)
	n_n4047<=n_n4046;

 always  @(posedge pclk)
	n_n4209<=n_n3503;

 always  @(posedge pclk)
	n_n4068<=n_n4065;

 always  @(posedge pclk)
	n_n3475<=n_n3474;

 always  @(posedge pclk)
	n_n4060<=n_n47;

 always  @(posedge pclk)
	n_n3998<=n_n36;

 always  @(posedge pclk)
	nsr5_4<=n_n41;

 always  @(posedge pclk)
	n_n3829<=n_n3828;

 always  @(posedge pclk)
	n_n3554<=n_n3553;

 always  @(posedge pclk)
	nsr3_9<=n_n40;

 always  @(posedge pclk)
	n_n3755<=n_n3754;

 always  @(posedge pclk)
	n_n3556<=n_n3555;

 always  @(posedge pclk)
	nsr5_5<=n_n39;

 always  @(posedge pclk)
	nsr5_3<=n_n44;

 always  @(posedge pclk)
	nsr5_2<=n_n45;

 always  @(posedge pclk)
	nsr5_7<=n_n38;

 always  @(posedge pclk)
	n_n3462<=n_n43;

 always  @(posedge pclk)
	nsr3_2<=n_n46;

 always  @(posedge pclk)
	nsr5_8<=n_n37;

 always  @(posedge pclk)
	n_n3460<=n_n42;

 assign puport_10_10_ = ( tin_puport_10_10_  &  (~ n_n3430) ) | ( n_n3430  &  n_n4068 ) ;
 assign puport_0_0_ = ( n_n3381  &  n_n2982 ) | ( tin_puport_0_0_  &  (~ n_n2982) ) ;
 assign pxport_10_10_ = ( n_n3887  &  n_n3556 ) | ( tin_pxport_10_10_  &  (~ n_n3556) ) ;
 assign pxport_0_0_ = ( tin_pxport_0_0_  &  (~ n_n3074) ) | ( n_n3074  &  n_n3628 ) ;
 assign puport_1_1_ = ( tin_puport_1_1_  &  (~ n_n3013) ) | ( n_n3013  &  n_n3065 ) ;
 assign pxport_1_1_ = ( tin_pxport_1_1_  &  (~ n_n3398) ) | ( n_n3398  &  n_n4259 ) ;
 assign puport_2_2_ = ( n_n3024  &  n_n3851 ) | ( tin_puport_2_2_  &  (~ n_n3851) ) ;
 assign pyport_10_10_ = ( tin_pyport_10_10_  &  (~ n_n3567) ) | ( n_n3567  &  n_n3182 ) ;
 assign pyport_0_0_ = ( tin_pyport_0_0_  &  (~ n_n3033) ) | ( n_n3033  &  n_n3928 ) ;
 assign pxport_2_2_ = ( n_n4149  &  n_n3453 ) | ( tin_pxport_2_2_  &  (~ n_n3453) ) ;
 assign puport_3_3_ = ( tin_puport_3_3_  &  (~ n_n3651) ) | ( n_n3651  &  n_n3493 ) ;
 assign pyport_1_1_ = ( n_n3060  &  n_n3000 ) | ( tin_pyport_1_1_  &  (~ n_n3000) ) ;
 assign pxport_7_7_ = ( tin_pxport_7_7_  &  (~ n_n3151) ) | ( n_n3151  &  n_n3855 ) ;
 assign puport_8_8_ = ( tin_puport_8_8_  &  (~ n_n4064) ) | ( n_n4064  &  n_n3901 ) ;
 assign pyport_6_6_ = ( tin_pyport_6_6_  &  (~ n_n3300) ) | ( n_n3300  &  n_n2968 ) ;
 assign pxport_8_8_ = ( n_n2995  &  n_n3448 ) | ( tin_pxport_8_8_  &  (~ n_n3448) ) ;
 assign puport_9_9_ = ( n_n2960  &  n_n3649 ) | ( tin_puport_9_9_  &  (~ n_n3649) ) ;
 assign pyport_7_7_ = ( tin_pyport_7_7_  &  (~ n_n3646) ) | ( n_n3646  &  n_n3002 ) ;
 assign pxport_9_9_ = ( tin_pxport_9_9_  &  (~ n_n3159) ) | ( n_n3159  &  n_n3067 ) ;
 assign pyport_8_8_ = ( tin_pyport_8_8_  &  (~ n_n2986) ) | ( n_n2986  &  n_n3498 ) ;
 assign pyport_9_9_ = ( n_n3170  &  n_n3622 ) | ( tin_pyport_9_9_  &  (~ n_n3622) ) ;
 assign pxport_3_3_ = ( tin_pxport_3_3_  &  (~ n_n3973) ) | ( n_n3973  &  n_n3199 ) ;
 assign puport_4_4_ = ( n_n3139  &  n_n3184 ) | ( tin_puport_4_4_  &  (~ n_n3184) ) ;
 assign pyport_2_2_ = ( n_n4014  &  n_n3554 ) | ( tin_pyport_2_2_  &  (~ n_n3554) ) ;
 assign pxport_4_4_ = ( tin_pxport_4_4_  &  (~ n_n3246) ) | ( n_n3246  &  n_n3563 ) ;
 assign puport_11_11_ = ( n_n3694  &  n_n3771 ) | ( tin_puport_11_11_  &  (~ n_n3771) ) ;
 assign puport_5_5_ = ( n_n3019  &  n_n3047 ) | ( tin_puport_5_5_  &  (~ n_n3047) ) ;
 assign pyport_3_3_ = ( tin_pyport_3_3_  &  (~ n_n3610) ) | ( n_n3610  &  n_n3122 ) ;
 assign pxport_5_5_ = ( n_n3128  &  n_n3755 ) | ( tin_pxport_5_5_  &  (~ n_n3755) ) ;
 assign puport_6_6_ = ( tin_puport_6_6_  &  (~ n_n3031) ) | ( n_n3031  &  n_n3728 ) ;
 assign pyport_4_4_ = ( tin_pyport_4_4_  &  (~ n_n2991) ) | ( n_n2991  &  n_n3327 ) ;
 assign pxport_11_11_ = ( tin_pxport_11_11_  &  (~ n_n3354) ) | ( n_n3354  &  n_n3698 ) ;
 assign pxport_6_6_ = ( n_n2971  &  n_n3044 ) | ( tin_pxport_6_6_  &  (~ n_n3044) ) ;
 assign puport_7_7_ = ( tin_puport_7_7_  &  (~ n_n3864) ) | ( n_n3864  &  n_n3309 ) ;
 assign pyport_11_11_ = ( tin_pyport_11_11_  &  (~ n_n3722) ) | ( n_n3722  &  n_n3689 ) ;
 assign pyport_5_5_ = ( n_n3767  &  n_n3606 ) | ( tin_pyport_5_5_  &  (~ n_n3606) ) ;
 assign n_n3032 = ( (~ preset)  &  n_n3033 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n2959 = ( wire2308 ) | ( wire2309 ) ;
 assign n_n3174 = ( wire2244 ) | ( n_n4027  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n2952 = ( wire2238 ) | ( wire2239 ) | ( n_n3871  &  wire806 ) ;
 assign n_n2973 = ( wire2162 ) | ( n_n3827  &  wire802 ) ;
 assign n_n3488 = ( wire2080 ) | ( wire811  &  (~ n_n3236)  &  n_n3111 ) | ( wire811  &  n_n3236  &  (~ n_n3111) ) ;
 assign n_n3596 = ( wire2068 ) | ( wire2069 ) | ( wire7130 ) ;
 assign n_n3969 = ( wire2066 ) | ( n_n4027  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n2970 = ( wire2063 ) | ( wire2064 ) ;
 assign n_n3259 = ( wire2061 ) | ( n_n4083  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n4007 = ( wire2059 ) | ( wire2060 ) ;
 assign n_n3483 = ( wire2057 ) | ( wire2058 ) ;
 assign n_n3073 = ( (~ preset)  &  n_n3074 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3653 = ( wire2041 ) | ( wire802  &  wire857 ) ;
 assign n_n3051 = ( wire2038 ) | ( wire2039 ) ;
 assign n_n3137 = ( wire2036 ) | ( wire2037 ) ;
 assign n_n4098 = ( wire2034 ) | ( wire2035 ) | ( n_n4099  &  wire806 ) ;
 assign n_n3007 = ( wire2031 ) | ( wire802  &  n_n4008 ) ;
 assign n_n3086 = ( wire2028 ) | ( wire811  &  (~ n_n3955)  &  n_n3543 ) | ( wire811  &  n_n3955  &  (~ n_n3543) ) ;
 assign n_n3602 = ( wire1968 ) | ( wire1969 ) | ( wire1970 ) | ( wire1971 ) ;
 assign n_n3499 = ( wire1966 ) | ( wire1967 ) | ( n_n3500  &  wire806 ) ;
 assign n_n3956 = ( wire1963 ) | ( n_n3996  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3752 = ( (~ preset)  &  ndn3_8  &  (~ ngfdn_3) ) | ( (~ preset)  &  ndn3_3  &  (~ ngfdn_3) ) ;
 assign n_n3941 = ( wire1959 ) | ( wire1960 ) ;
 assign n_n3299 = ( (~ preset)  &  n_n3300 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3284 = ( wire1955 ) | ( wire1956 ) ;
 assign n_n3618 = ( (~ preset)  &  nen5_9  &  (~ nld3_9) ) | ( (~ preset)  &  (~ nld3_9)  &  (~ nsr5_8) ) ;
 assign n_n3353 = ( (~ preset)  &  n_n3354 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n2972 = ( wire1950 ) | ( n_n4027  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3070 = ( wire1948 ) | ( n_n3974  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3454 = ( wire1944 ) | ( wire811  &  (~ n_n4153)  &  n_n3035 ) | ( wire811  &  n_n4153  &  (~ n_n3035) ) ;
 assign n_n3640 = ( (~ preset)  &  wire860  &  nrq5_6 ) | ( (~ preset)  &  n_n3761  &  (~ nrq5_6) ) ;
 assign n_n2992 = ( wire1908 ) | ( wire802  &  (~ n_n4189)  &  n_n3892 ) | ( wire802  &  n_n4189  &  (~ n_n3892) ) ;
 assign n_n3063 = ( (~ preset)  &  ndn5_16  &  (~ nld3_9) ) ;
 assign n_n4147 = ( wire1905 ) | ( wire1906 ) ;
 assign n_n3772 = ( wire1904 ) | ( n_n3974  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3132 = ( wire1902 ) | ( n_n3912  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n2969 = ( wire1898 ) | ( pxport_10_10_  &  wire799 ) ;
 assign n_n3616 = ( wire1894 ) | ( wire802  &  wire862 ) ;
 assign n_n3183 = ( (~ preset)  &  n_n3184 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3523 = ( wire1889 ) | ( wire1890 ) ;
 assign n_n3004 = ( wire1886 ) | ( puport_10_10_  &  wire799 ) ;
 assign n_n3206 = ( (~ preset)  &  n_n4072  &  (~ nrq2_2) ) ;
 assign n_n2984 = ( wire1882 ) | ( pxport_4_4_  &  wire799 ) ;
 assign n_n4038 = ( wire1879 ) | ( n_n4227  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3481 = ( wire1877 ) | ( n_n4197  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3322 = ( (~ preset)  &  wire857  &  nrq5_6 ) | ( (~ preset)  &  n_n3908  &  (~ nrq5_6) ) ;
 assign n_n3144 = ( wire1873 ) | ( n_n4145  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3401 = ( wire1870 ) | ( puport_7_7_  &  wire799 ) ;
 assign n_n3584 = ( wire1867 ) | ( n_n3949  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3926 = ( wire1865 ) | ( wire1866 ) ;
 assign n_n2958 = ( (~ preset)  &  n_n4182  &  (~ nrq2_2) ) ;
 assign n_n3739 = ( (~ preset)  &  (~ nsr5_4) ) ;
 assign n_n2990 = ( (~ preset)  &  n_n2991 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3744 = ( (~ preset)  &  n_n3745 ) | ( (~ preset)  &  nrq2_2 ) ;
 assign n_n3690 = ( (~ preset)  &  n_n3691  &  (~ nrq2_2) ) ;
 assign n_n3018 = ( wire1859 ) | ( wire1860 ) ;
 assign n_n3334 = ( wire1857 ) | ( n_n3974  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n2997 = ( wire1855 ) | ( n_n3949  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3566 = ( (~ preset)  &  n_n3567 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3798 = ( wire1851 ) | ( n_n3992  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n2974 = ( wire1848 ) | ( pyport_9_9_  &  wire799 ) ;
 assign n_n3115 = ( wire1844 ) | ( puport_4_4_  &  wire799 ) ;
 assign n_n3811 = ( (~ preset)  &  (~ pdn) ) ;
 assign n_n3059 = ( wire1841 ) | ( wire1842 ) ;
 assign n_n3325 = ( (~ preset)  &  (~ n_n3142)  &  wire7205 ) ;
 assign n_n3052 = ( wire1835 ) | ( wire1836 ) ;
 assign n_n3030 = ( (~ preset)  &  n_n3031 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3153 = ( wire1831 ) | ( wire1832 ) | ( n_n3813  &  wire806 ) ;
 assign n_n3705 = ( wire1828 ) | ( wire1829 ) ;
 assign n_n3432 = ( wire1826 ) | ( wire1827 ) ;
 assign n_n2983 = ( wire1823 ) | ( pxport_6_6_  &  wire799 ) ;
 assign n_n3040 = ( wire1819 ) | ( wire802  &  (~ n_n4202)  &  n_n4062 ) | ( wire802  &  n_n4202  &  (~ n_n4062) ) ;
 assign n_n3209 = ( wire1816 ) | ( n_n3992  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3165 = ( wire1814 ) | ( wire1815 ) | ( wire7209 ) ;
 assign n_n3057 = ( wire1809 ) | ( puport_1_1_  &  wire799 ) ;
 assign n_n3127 = ( wire1806 ) | ( wire1807 ) ;
 assign n_n4254 = ( wire1804 ) | ( wire1805 ) ;
 assign n_n3163 = ( wire1802 ) | ( wire1803 ) ;
 assign n_n3041 = ( (~ preset)  &  (~ nsr5_3) ) ;
 assign n_n3972 = ( (~ preset)  &  n_n3973 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3150 = ( (~ preset)  &  n_n3151 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3814 = ( wire1797 ) | ( wire816  &  (~ n_n4189)  &  n_n3892 ) | ( wire816  &  n_n4189  &  (~ n_n3892) ) ;
 assign n_n3349 = ( wire1794 ) | ( wire1795 ) | ( n_n3808  &  wire806 ) ;
 assign n_n3247 = ( wire1790 ) | ( pxport_5_5_  &  wire799 ) ;
 assign n_n3661 = ( wire1787 ) | ( n_n4027  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3652 = ( wire1785 ) | ( n_n3996  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3315 = ( wire1783 ) | ( wire1784 ) | ( n_n3844  &  wire806 ) ;
 assign n_n3316 = ( wire1780 ) | ( wire1781 ) | ( n_n3810  &  wire806 ) ;
 assign n_n3456 = ( wire1777 ) | ( n_n4145  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3168 = ( wire1775 ) | ( wire1776 ) ;
 assign n_n3037 = ( (~ preset)  &  n_n3346 ) | ( (~ preset)  &  nrq2_2 ) ;
 assign n_n3119 = ( (~ preset)  &  n_n3324  &  (~ nrq2_2) ) ;
 assign n_n2966 = ( (~ preset)  &  n_n3312  &  (~ nrq2_2) ) ;
 assign n_n3795 = ( wire1769 ) | ( wire816  &  n_n3975 ) ;
 assign n_n4113 = ( wire1708 ) | ( wire802  &  n_n4168 ) ;
 assign n_n3014 = ( wire1705 ) | ( wire802  &  (~ n_n3118)  &  n_n3857 ) | ( wire802  &  n_n3118  &  (~ n_n3857) ) ;
 assign n_n3103 = ( wire1702 ) | ( n_n3992  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n4238 = ( wire1700 ) | ( wire1701 ) | ( n_n4239  &  wire806 ) ;
 assign n_n3210 = ( wire1697 ) | ( n_n3965  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3113 = ( wire1693 ) | ( wire1694 ) ;
 assign n_n3740 = ( wire1690 ) | ( pyport_0_0_  &  wire799 ) ;
 assign n_n3202 = ( wire1687 ) | ( n_n3974  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3720 = ( wire1686 ) | ( n_n4197  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3314 = ( (~ preset)  &  n_n4223  &  (~ nrq2_2) ) ;
 assign n_n3650 = ( (~ preset)  &  n_n3651 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3046 = ( (~ preset)  &  n_n3047 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3458 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) | ( (~ preset)  &  nen5_9  &  (~ ndn5_9)  &  (~ nld3_9) ) ;
 assign n_n3409 = ( wire1677 ) | ( wire1678 ) | ( n_n3924  &  wire806 ) ;
 assign n_n3227 = ( wire1674 ) | ( wire1675 ) | ( n_n3923  &  wire806 ) ;
 assign n_n2963 = ( wire1669 ) | ( wire1670 ) | ( wire1671 ) | ( wire1672 ) ;
 assign n_n3005 = ( n_n3042 ) | ( wire1666 ) | ( wire1667 ) ;
 assign n_n2998 = ( wire1660 ) | ( wire802  &  wire7274 ) | ( wire802  &  wire7275 ) ;
 assign n_n3638 = ( (~ preset)  &  (~ n_n3460) ) | ( (~ preset)  &  wire2075 ) ;
 assign n_n4063 = ( (~ preset)  &  n_n4064 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3240 = ( wire1656 ) | ( wire1657 ) ;
 assign n_n3987 = ( wire1654 ) | ( n_n4083  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3177 = ( wire1652 ) | ( n_n4145  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n2996 = ( (~ preset)  &  n_n3469  &  (~ nrq2_2) ) ;
 assign n_n3061 = ( n_n3542 ) | ( wire1649 ) | ( wire1650 ) ;
 assign n_n3091 = ( wire1646 ) | ( wire1647 ) | ( wire797  &  n_n3099 ) ;
 assign n_n3178 = ( wire1645 ) | ( wire802  &  (~ n_n4153)  &  n_n3035 ) | ( wire802  &  n_n4153  &  (~ n_n3035) ) ;
 assign n_n3193 = ( wire1642 ) | ( wire1643 ) ;
 assign n_n3016 = ( (~ preset)  &  ndn5_6  &  (~ nld3_9) ) | ( (~ preset)  &  (~ nld3_9)  &  nrq5_6 ) ;
 assign n_n3712 = ( wire1625 ) | ( wire1626 ) ;
 assign n_n4053 = ( wire1623 ) | ( wire1624 ) ;
 assign n_n3310 = ( wire1622 ) | ( n_n3912  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3431 = ( wire1619 ) | ( n_n3949  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3599 = ( wire1617 ) | ( wire1618 ) | ( wire7294 ) ;
 assign n_n3146 = ( wire1613 ) | ( wire1614 ) ;
 assign n_n3058 = ( wire1610 ) | ( pyport_11_11_  &  wire799 ) ;
 assign n_n3914 = ( wire1607 ) | ( wire1608 ) ;
 assign n_n3389 = ( (~ preset)  &  n_n3578  &  n_n3460  &  (~ wire2075) ) ;
 assign n_n3379 = ( wire1605 ) | ( wire1606 ) ;
 assign n_n3633 = ( wire1602 ) | ( pxport_8_8_  &  wire799 ) ;
 assign n_n3147 = ( wire1598 ) | ( wire1599 ) | ( wire1600 ) ;
 assign n_n3586 = ( wire1596 ) | ( wire1597 ) | ( n_n4224  &  wire806 ) ;
 assign n_n4089 = ( wire1592 ) | ( pyport_6_6_  &  wire799 ) ;
 assign n_n3963 = ( wire1589 ) | ( wire1590 ) ;
 assign n_n3213 = ( wire1588 ) | ( wire802  &  wire860 ) ;
 assign n_n3538 = ( (~ preset)  &  (~ nsr5_7) ) ;
 assign n_n4055 = ( wire1585 ) | ( wire1586 ) ;
 assign n_n3009 = ( wire1582 ) | ( pxport_9_9_  &  wire799 ) ;
 assign n_n3050 = ( wire1577 ) | ( wire1578 ) ;
 assign n_n4229 = ( wire1574 ) | ( pyport_3_3_  &  wire799 ) ;
 assign n_n3595 = ( wire1571 ) | ( wire1572 ) ;
 assign n_n3245 = ( (~ preset)  &  n_n3246 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n2955 = ( wire1567 ) | ( wire1568 ) | ( n_n3919  &  wire806 ) ;
 assign n_n3172 = ( wire1564 ) | ( n_n4227  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3710 = ( wire1562 ) | ( n_n4018  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n2979 = ( wire1559 ) | ( pyport_2_2_  &  wire799 ) ;
 assign n_n3012 = ( (~ preset)  &  n_n3013 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3397 = ( (~ preset)  &  n_n3398 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3211 = ( wire1553 ) | ( wire802  &  (~ n_n3236)  &  n_n3111 ) | ( wire802  &  n_n3236  &  (~ n_n3111) ) ;
 assign n_n3863 = ( (~ preset)  &  n_n3864 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n4029 = ( wire1548 ) | ( n_n3974  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3487 = ( wire1546 ) | ( (~ preset)  &  n_n3513  &  (~ nrq5_6) ) ;
 assign n_n4085 = ( wire1544 ) | ( wire1545 ) | ( n_n4086  &  wire806 ) ;
 assign n_n3664 = ( wire1539 ) | ( wire1540 ) ;
 assign n_n3609 = ( (~ preset)  &  n_n3610 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3266 = ( wire1535 ) | ( n_n4008  &  wire816 ) ;
 assign n_n3658 = ( wire1534 ) | ( n_n4227  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3244 = ( wire1530 ) | ( wire802  &  wire869 ) ;
 assign n_n3200 = ( wire1526 ) | ( wire1528 ) | ( wire7304 ) ;
 assign n_n2985 = ( (~ preset)  &  n_n2986 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n2957 = ( (~ preset)  &  n_n4135  &  (~ nrq2_2) ) ;
 assign n_n3348 = ( (~ preset)  &  (~ nsr5_5) ) ;
 assign n_n3683 = ( wire1520 ) | ( wire816  &  wire870 ) ;
 assign n_n3615 = ( wire1517 ) | ( n_n3912  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n4231 = ( wire1514 ) | ( pyport_1_1_  &  wire799 ) ;
 assign n_n3287 = ( (~ preset)  &  ndn3_11  &  (~ ngfdn_3) ) ;
 assign n_n3049 = ( wire1511 ) | ( n_n4018  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3558 = ( wire1509 ) | ( n_n3965  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3263 = ( wire1507 ) | ( wire1508 ) | ( n_n3940  &  wire806 ) ;
 assign n_n3946 = ( wire1505 ) | ( wire816  &  wire869 ) ;
 assign n_n3614 = ( wire1503 ) | ( n_n4018  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3437 = ( wire1477 ) | ( wire802  &  n_n3746 ) ;
 assign n_n3180 = ( wire1475 ) | ( wire1476 ) ;
 assign n_n2978 = ( wire1472 ) | ( pyport_4_4_  &  wire799 ) ;
 assign n_n4256 = ( wire1469 ) | ( wire1470 ) ;
 assign n_n4139 = ( wire1467 ) | ( wire1468 ) | ( n_n4140  &  wire806 ) ;
 assign n_n3853 = ( wire1464 ) | ( wire1465 ) ;
 assign n_n3530 = ( (~ preset)  &  ndn3_3  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_2) ) ;
 assign n_n4011 = ( wire1460 ) | ( wire1461 ) ;
 assign n_n3648 = ( (~ preset)  &  n_n3649 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3064 = ( wire1456 ) | ( wire1457 ) ;
 assign n_n3276 = ( wire1453 ) | ( wire1454 ) | ( wire7347 ) ;
 assign n_n3570 = ( wire1450 ) | ( wire1451 ) | ( n_n3890  &  wire806 ) ;
 assign n_n3339 = ( wire1446 ) | ( wire1447 ) | ( wire1448 ) ;
 assign n_n3524 = ( wire1445 ) | ( n_n3996  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3241 = ( wire1443 ) | ( wire816  &  (~ n_n4202)  &  n_n4062 ) | ( wire816  &  n_n4202  &  (~ n_n4062) ) ;
 assign n_n2956 = ( wire1440 ) | ( wire1441 ) | ( n_n3868  &  wire806 ) ;
 assign n_n3145 = ( wire1437 ) | ( n_n3965  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3592 = ( wire1435 ) | ( wire1436 ) | ( n_n3918  &  wire806 ) ;
 assign n_n3102 = ( wire1432 ) | ( n_n4197  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3093 = ( wire1430 ) | ( wire1431 ) | ( wire7354 ) ;
 assign n_n3191 = ( wire1426 ) | ( wire1427 ) | ( n_n4136  &  wire806 ) ;
 assign n_n3476 = ( (~ preset)  &  ndn2_2  &  wire917 ) ;
 assign n_n4041 = ( wire1423 ) | ( n_n3912  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3479 = ( wire1421 ) | ( wire1422 ) | ( n_n4176  &  wire806 ) ;
 assign n_n3895 = ( wire1418 ) | ( wire1419 ) ;
 assign n_n3158 = ( (~ preset)  &  n_n3159 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3249 = ( wire1413 ) | ( pxport_3_3_  &  wire799 ) ;
 assign n_n3717 = ( wire1408 ) | ( wire1411 ) | ( wire7364 ) ;
 assign n_n3106 = ( wire1405 ) | ( wire1406 ) | ( wire1407 ) ;
 assign n_n4020 = ( wire1403 ) | ( n_n4018  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3765 = ( wire1401 ) | ( wire1402 ) ;
 assign n_n2999 = ( (~ preset)  &  n_n3000 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3909 = ( wire1398 ) | ( n_n3965  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3726 = ( wire1395 ) | ( wire1396 ) ;
 assign n_n4110 = ( wire1393 ) | ( wire811  &  wire7274 ) | ( wire811  &  wire7275 ) ;
 assign n_n3620 = ( wire1391 ) | ( (~ preset)  &  (~ pdn)  &  ngfdn_3 ) ;
 assign n_n2980 = ( wire1387 ) | ( wire1388 ) | ( wire1390 ) | ( wire7375 ) ;
 assign n_n3696 = ( wire1384 ) | ( wire1385 ) ;
 assign n_n4105 = ( wire1381 ) | ( puport_3_3_  &  wire799 ) ;
 assign n_n4094 = ( wire1378 ) | ( wire1379 ) | ( n_n4095  &  wire806 ) ;
 assign n_n3497 = ( wire1375 ) | ( wire1376 ) ;
 assign n_n3692 = ( wire1373 ) | ( wire1374 ) ;
 assign n_n3308 = ( wire1371 ) | ( wire1372 ) ;
 assign n_n3847 = ( wire1346 ) | ( wire1347 ) | ( wire1348 ) | ( wire1349 ) ;
 assign n_n3801 = ( wire1344 ) | ( wire1345 ) | ( n_n3971  &  wire806 ) ;
 assign n_n3162 = ( wire1341 ) | ( n_n3965  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3189 = ( wire1338 ) | ( puport_8_8_  &  wire799 ) ;
 assign n_n3465 = ( (~ preset)  &  nak3_9 ) ;
 assign n_n3043 = ( (~ preset)  &  n_n3044 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n4174 = ( (~ preset)  &  n_n4222  &  (~ nrq2_2) ) ;
 assign n_n2976 = ( wire1282 ) | ( n_n4083  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3008 = ( wire1279 ) | ( wire802  &  n_n3975 ) ;
 assign n_n4032 = ( wire1276 ) | ( wire802  &  (~ n_n4052)  &  n_n3729 ) | ( wire802  &  n_n4052  &  (~ n_n3729) ) ;
 assign n_n3305 = ( (~ preset)  &  (~ pdn)  &  ndn1_4 ) ;
 assign n_n3204 = ( wire1273 ) | ( n_n3996  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3028 = ( wire1271 ) | ( n_n3949  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3075 = ( wire1270 ) | ( n_n4083  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3087 = ( wire1267 ) | ( wire1268 ) | ( n_n4177  &  wire806 ) ;
 assign n_n3326 = ( wire1264 ) | ( wire1265 ) ;
 assign n_n3817 = ( wire1262 ) | ( wire1263 ) ;
 assign n_n3136 = ( wire1261 ) | ( n_n3996  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3668 = ( wire1258 ) | ( wire1259 ) | ( n_n3843  &  wire806 ) ;
 assign n_n3068 = ( wire1256 ) | ( n_n3949  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3413 = ( wire1253 ) | ( wire1254 ) | ( n_n3842  &  wire806 ) ;
 assign n_n3222 = ( wire1248 ) | ( wire1249 ) | ( wire1250 ) | ( wire1251 ) ;
 assign n_n3627 = ( wire1246 ) | ( wire1247 ) ;
 assign n_n3399 = ( wire1243 ) | ( puport_2_2_  &  wire799 ) ;
 assign n_n2994 = ( wire1240 ) | ( wire1241 ) ;
 assign n_n2987 = ( pready_0_0_  &  (~ nlak3_2)  &  (~ n_n4253)  &  wire7468 ) ;
 assign n_n3429 = ( (~ preset)  &  n_n3430 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3372 = ( wire1235 ) | ( pxport_11_11_  &  wire799 ) ;
 assign n_n3915 = ( wire1232 ) | ( wire1233 ) ;
 assign n_n3452 = ( (~ preset)  &  n_n3453 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3447 = ( (~ preset)  &  n_n3448 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3156 = ( (~ preset)  &  n_n4134  &  (~ nrq2_2) ) ;
 assign n_n3201 = ( wire1226 ) | ( wire1227 ) | ( n_n3800  &  wire806 ) ;
 assign n_n3472 = ( wire1223 ) | ( n_n4197  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3611 = ( wire1221 ) | ( n_n4227  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n4074 = ( wire1219 ) | ( n_n4197  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3449 = ( wire1215 ) | ( wire1216 ) | ( wire1217 ) | ( wire1218 ) ;
 assign n_n3904 = ( (~ preset)  &  n_n3905  &  (~ nrq2_2) ) ;
 assign n_n3542 = ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_9) ) ;
 assign n_n2964 = ( wire1213 ) | ( wire1214 ) | ( wire7478 ) ;
 assign n_n4028 = ( wire1210 ) | ( n_n4227  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3423 = ( wire1208 ) | ( n_n4018  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n2977 = ( wire1205 ) | ( n_n3974  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3130 = ( wire1203 ) | ( wire1204 ) | ( n_n4208  &  wire806 ) ;
 assign n_n3042 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3338 = ( (~ preset)  &  n_n4073  &  (~ nrq2_2) ) ;
 assign n_n3078 = ( (~ preset)  &  n_n3345  &  (~ nrq2_2) ) ;
 assign n_n3374 = ( (~ preset)  &  n_n3375  &  (~ nrq2_2) ) ;
 assign n_n3425 = ( (~ preset)  &  n_n3426  &  (~ nrq2_2) ) ;
 assign n_n3486 = ( wire1200 ) | ( n_n3996  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3104 = ( wire1197 ) | ( pxport_7_7_  &  wire799 ) ;
 assign n_n3129 = ( wire1194 ) | ( wire1195 ) | ( n_n3807  &  wire806 ) ;
 assign n_n3152 = ( wire1190 ) | ( pyport_7_7_  &  wire799 ) ;
 assign n_n3053 = ( wire1187 ) | ( wire1188 ) | ( wire7483 ) ;
 assign n_n3133 = ( wire1184 ) | ( n_n3949  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3770 = ( (~ preset)  &  n_n3771 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3003 = ( wire1179 ) | ( wire1180 ) ;
 assign n_n3010 = ( wire1176 ) | ( pyport_10_10_  &  wire799 ) ;
 assign n_n3666 = ( wire1174 ) | ( wire802  &  (~ n_n3955)  &  n_n3543 ) | ( wire802  &  n_n3955  &  (~ n_n3543) ) ;
 assign n_n3605 = ( (~ preset)  &  n_n3606 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3899 = ( wire1169 ) | ( wire1170 ) ;
 assign n_n2961 = ( wire1166 ) | ( puport_11_11_  &  wire799 ) ;
 assign n_n4166 = ( wire1163 ) | ( wire816  &  n_n4168 ) ;
 assign n_n3511 = ( wire1161 ) | ( wire1162 ) ;
 assign n_n3022 = ( wire1159 ) | ( wire1160 ) ;
 assign n_n3155 = ( (~ preset)  &  n_n3445  &  (~ nrq2_2) ) ;
 assign n_n3117 = ( wire1157 ) | ( (~ preset)  &  n_n3862  &  (~ nrq5_6) ) ;
 assign n_n3027 = ( wire1153 ) | ( wire1154 ) | ( wire1155 ) | ( wire1156 ) ;
 assign n_n3885 = ( wire1151 ) | ( wire1152 ) ;
 assign n_n3335 = ( (~ preset)  &  n_n3746  &  nrq5_6 ) | ( (~ preset)  &  n_n3336  &  (~ nrq5_6) ) ;
 assign n_n3197 = ( wire1147 ) | ( wire1148 ) ;
 assign n_n3034 = ( wire1145 ) | ( wire1146 ) | ( n_n3470  &  wire806 ) ;
 assign n_n2962 = ( wire1141 ) | ( puport_9_9_  &  wire799 ) ;
 assign n_n3823 = ( wire1138 ) | ( n_n3912  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3160 = ( (~ preset)  &  (~ nsr5_2) ) ;
 assign n_n3029 = ( (~ preset)  &  (~ nsr5_8) ) ;
 assign n_n3406 = ( wire1136 ) | ( wire1137 ) | ( n_n4119  &  wire806 ) ;
 assign n_n3787 = ( wire1133 ) | ( wire1134 ) ;
 assign n_n3506 = ( wire1131 ) | ( wire1132 ) | ( n_n4118  &  wire806 ) ;
 assign n_n3216 = ( wire1129 ) | ( wire802  &  wire870 ) ;
 assign n_n3215 = ( wire1124 ) | ( wire1125 ) ;
 assign n_n3721 = ( (~ preset)  &  n_n3722 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3173 = ( wire1120 ) | ( n_n3912  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3785 = ( wire1117 ) | ( pyport_5_5_  &  wire799 ) ;
 assign n_n3277 = ( wire1114 ) | ( wire1115 ) | ( wire7495 ) ;
 assign n_n3562 = ( wire1110 ) | ( wire1111 ) ;
 assign n_n4023 = ( wire1108 ) | ( n_n3992  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3015 = ( wire1106 ) | ( n_n4145  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n3120 = ( wire1104 ) | ( wire1105 ) ;
 assign n_n3621 = ( (~ preset)  &  n_n3622 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3645 = ( (~ preset)  &  n_n3646 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n2965 = ( (~ preset)  &  n_n3294  &  (~ nrq2_2) ) ;
 assign n_n3913 = ( wire1098 ) | ( wire1099 ) ;
 assign n_n3695 = ( wire1097 ) | ( n_n3992  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n4217 = ( wire1093 ) | ( pxport_0_0_  &  wire799 ) ;
 assign n_n3416 = ( wire1089 ) | ( pxport_2_2_  &  wire799 ) ;
 assign n_n3687 = ( wire1086 ) | ( wire1087 ) ;
 assign n_n3320 = ( wire1084 ) | ( n_n4018  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3559 = ( (~ preset)  &  wire862  &  nrq5_6 ) | ( (~ preset)  &  n_n3794  &  (~ nrq5_6) ) ;
 assign n_n4044 = ( wire1081 ) | ( n_n4197  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3435 = ( wire1078 ) | ( n_n4083  &  wire796  &  ndn_latch5_3 ) ;
 assign n_n3967 = ( wire1076 ) | ( n_n4027  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3352 = ( wire1073 ) | ( pyport_8_8_  &  wire799 ) ;
 assign n_n3321 = ( wire1071 ) | ( wire811  &  (~ n_n4052)  &  n_n3729 ) | ( wire811  &  n_n4052  &  (~ n_n3729) ) ;
 assign n_n3318 = ( wire1067 ) | ( puport_5_5_  &  wire799 ) ;
 assign n_n3066 = ( wire1064 ) | ( wire1065 ) ;
 assign n_n2967 = ( wire1062 ) | ( wire1063 ) ;
 assign n_n3707 = ( (~ preset)  &  n_n3708  &  (~ nrq2_2) ) ;
 assign n_n3194 = ( wire1060 ) | ( wire1061 ) ;
 assign n_n3825 = ( wire1058 ) | ( n_n3827  &  wire816 ) ;
 assign n_n3123 = ( wire1056 ) | ( wire1057 ) | ( n_n3872  &  wire806 ) ;
 assign n_n3579 = ( wire1052 ) | ( pxport_1_1_  &  wire799 ) ;
 assign n_n3491 = ( wire1049 ) | ( wire1050 ) ;
 assign n_n3980 = ( wire1045 ) | ( (~ preset)  &  n_n3981  &  (~ nrq5_6) ) ;
 assign n_n3859 = ( wire1037 ) | ( (~ wire841)  &  wire7501 ) | ( wire841  &  wire7502 ) ;
 assign n_n3723 = ( wire1032 ) | ( wire1034 ) | ( wire7508 ) ;
 assign n_n3231 = ( (~ preset)  &  (~ nld3_9)  &  ndn5_10 ) | ( (~ preset)  &  (~ nld3_9)  &  (~ nsr5_7) ) ;
 assign n_n3400 = ( wire1026 ) | ( puport_0_0_  &  wire799 ) ;
 assign n_n3048 = ( wire1023 ) | ( n_n4083  &  wire796  &  ndn_latch5_7 ) ;
 assign n_n3804 = ( wire1020 ) | ( puport_6_6_  &  wire799 ) ;
 assign n_n3001 = ( wire1017 ) | ( wire1018 ) ;
 assign n_n2953 = ( (~ preset)  &  n_n3388 ) | ( (~ preset)  &  nrq2_2 ) ;
 assign n_n2981 = ( (~ preset)  &  n_n2982 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3850 = ( (~ preset)  &  n_n3851 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3332 = ( wire1007 ) | ( n_n3142  &  wire7511 ) | ( (~ wire7205)  &  wire7511 ) ;
 assign n_n2988 = ( (~ preset)  &  n_n2989 ) | ( (~ preset)  &  nrq2_2 ) ;
 assign n_n3390 = ( (~ preset)  &  n_n4181  &  (~ nrq2_2) ) ;
 assign n_n3589 = ( wire1002 ) | ( wire1003 ) | ( n_n3939  &  wire806 ) ;
 assign n_n3192 = ( wire999 ) | ( wire1000 ) ;
 assign n_n3273 = ( wire998 ) | ( wire816  &  (~ n_n3118)  &  n_n3857 ) | ( wire816  &  n_n3118  &  (~ n_n3857) ) ;
 assign n_n2975 = ( wire996 ) | ( n_n4145  &  wire796  &  ndn_latch5_5 ) ;
 assign n_n3662 = ( wire993 ) | ( n_n4227  &  wire796  &  ndn_latch5_2 ) ;
 assign n_n3038 = ( (~ preset)  &  n_n3468  &  (~ nrq2_2) ) ;
 assign n_n3671 = ( wire991 ) | ( wire992 ) | ( n_n4252  &  wire806 ) ;
 assign n_n3190 = ( wire987 ) | ( wire988 ) | ( n_n4183  &  wire806 ) ;
 assign n_n3101 = ( wire985 ) | ( n_n3965  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3366 = ( wire983 ) | ( n_n3992  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3958 = ( wire980 ) | ( n_n4027  &  wire796  &  ndn_latch5_8 ) ;
 assign n_n4046 = ( wire979 ) | ( n_n4145  &  wire796  &  ndn_latch5_4 ) ;
 assign n_n3503 = ( wire976 ) | ( wire977 ) | ( n_n4209  &  wire806 ) ;
 assign n_n4065 = ( wire972 ) | ( wire973 ) ;
 assign n_n3474 = ( wire970 ) | ( wire971 ) ;
 assign n_n47 = ( wire963 ) | ( wire964 ) | ( wire7527 ) | ( wire7529 ) ;
 assign n_n36 = ( preset ) | ( pdn  &  n_n3998 ) | ( (~ preset)  &  (~ pdn)  &  (~ n_n4253) ) ;
 assign n_n41 = ( preset ) | ( wire7532 ) | ( nsr5_4  &  nsr5_3 ) ;
 assign n_n3828 = ( wire938 ) | ( wire954 ) ;
 assign n_n3553 = ( (~ preset)  &  n_n3554 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n40 = ( wire7533 ) | ( nsr3_9  &  (~ nak3_9) ) ;
 assign n_n3754 = ( (~ preset)  &  n_n3755 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n3555 = ( (~ preset)  &  n_n3556 ) | ( (~ preset)  &  ndn5_9  &  (~ nld3_9) ) ;
 assign n_n39 = ( preset ) | ( wire7534 ) | ( nsr5_4  &  nsr5_5 ) ;
 assign n_n44 = ( preset ) | ( wire7535 ) | ( nsr5_3  &  nsr5_2 ) ;
 assign n_n45 = ( wire875 ) | ( (~ nak5_2)  &  nrq5_2 ) | ( nsr5_2  &  (~ nrq5_2) ) ;
 assign n_n38 = ( preset ) | ( wire7537 ) | ( nsr5_5  &  nsr5_7 ) ;
 assign n_n43 = ( preset ) | ( (~ n_n3460) ) | ( wire876 ) | ( wire2075 ) ;
 assign n_n46 = ( preset ) | ( pdn ) | ( wire835 ) ;
 assign n_n37 = ( preset ) | ( wire7539 ) | ( nsr5_7  &  nsr5_8 ) ;
 assign n_n42 = ( wire1008 ) | ( wire7512 ) ;
 assign wire806 = ( wire6975  &  wire6976 ) | ( (~ n_n4253)  &  wire6977 ) ;
 assign n_n3827 = ( (~ n_n3779)  &  n_n4202  &  n_n3897 ) | ( (~ n_n3779)  &  n_n4202  &  n_n4062 ) | ( n_n3779  &  (~ n_n4202)  &  n_n4062 ) | ( (~ n_n3779)  &  n_n3897  &  (~ n_n4062) ) | ( n_n3779  &  (~ n_n3897)  &  (~ n_n4062) ) ;
 assign wire802 = ( (~ preset)  &  nen5_9  &  (~ ndn5_9) ) ;
 assign wire811 = ( (~ preset)  &  nrq5_6 ) ;
 assign n_n4170 = ( wire6930 ) | ( n_n4165  &  nrq5_5 ) | ( n_n4165  &  nrq5_2 ) ;
 assign wire797 = ( (~ preset)  &  (~ n_n3575)  &  n_n4214  &  n_n3462 ) ;
 assign wire918 = ( n_n4004 ) | ( (~ n_n4004)  &  n_n3961 ) | ( (~ n_n4004)  &  n_n4126 ) | ( (~ n_n4004)  &  (~ n_n4060) ) ;
 assign wire799 = ( (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire857 = ( (~ n_n3236)  &  n_n3950  &  n_n3111 ) | ( n_n3236  &  (~ n_n3950)  &  n_n3111 ) | ( (~ n_n3950)  &  (~ n_n3111)  &  wire849 ) | ( (~ n_n3236)  &  n_n3950  &  (~ wire849) ) | ( n_n3950  &  (~ n_n3111)  &  (~ wire849) ) ;
 assign n_n4008 = ( wire2189  &  wire7007 ) | ( wire2190  &  wire7007 ) | ( wire2189  &  wire7008 ) | ( wire2190  &  wire7008 ) | ( (~ wire2189)  &  (~ wire2190)  &  (~ wire7007)  &  (~ wire7008) ) ;
 assign n_n4144 = ( n_n3949  &  n_n3948 ) | ( n_n3949  &  wire1974 ) | ( n_n3948  &  wire1974 ) | ( n_n3949  &  wire7173 ) | ( n_n3948  &  wire7173 ) ;
 assign n_n3948 = ( n_n4083  &  n_n4082 ) | ( n_n4083  &  wire2022 ) | ( n_n4082  &  wire2022 ) | ( n_n4083  &  wire7149 ) | ( n_n4082  &  wire7149 ) ;
 assign n_n4131 = ( wire7173 ) | ( n_n4136  &  nrq5_5 ) | ( n_n4136  &  nrq5_2 ) ;
 assign wire813 = ( (~ preset)  &  (~ n_n3575)  &  n_n4214  &  n_n3462 ) ;
 assign wire875 = ( preset ) | ( nld3_9 ) ;
 assign wire860 = ( (~ n_n3955)  &  n_n3543  &  n_n3635 ) | ( (~ n_n3955)  &  (~ wire851)  &  n_n3635 ) | ( (~ n_n3543)  &  (~ wire851)  &  n_n3635 ) | ( n_n3955  &  n_n3543  &  (~ n_n3635) ) | ( (~ n_n3543)  &  wire851  &  (~ n_n3635) ) ;
 assign wire862 = ( n_n3569  &  (~ n_n4153)  &  (~ wire852) ) | ( (~ n_n3569)  &  n_n4153  &  n_n3035 ) | ( n_n3569  &  (~ n_n4153)  &  n_n3035 ) | ( (~ n_n3569)  &  wire852  &  (~ n_n3035) ) | ( n_n3569  &  (~ wire852)  &  (~ n_n3035) ) ;
 assign n_n4000 = ( n_n3460  &  (~ n_n3549)  &  wire955 ) ;
 assign wire796 = ( (~ preset)  &  (~ wire2247)  &  (~ wire6973) ) | ( (~ preset)  &  (~ wire2247)  &  (~ wire6974) ) ;
 assign n_n3944 = ( wire6933 ) | ( n_n4070  &  nrq5_5 ) | ( n_n4070  &  nrq5_2 ) ;
 assign n_n3301 = ( n_n4093 ) | ( n_n4246 ) | ( (~ n_n4093)  &  wire940 ) ;
 assign wire839 = ( n_n3369 ) | ( n_n4093 ) | ( n_n4246 ) | ( (~ n_n4093)  &  wire940 ) ;
 assign wire816 = ( (~ preset)  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign n_n3975 = ( (~ wire2196)  &  (~ wire2197)  &  wire2235 ) | ( (~ wire2196)  &  (~ wire2197)  &  wire2236 ) | ( wire2196  &  (~ wire2235)  &  (~ wire2236) ) | ( wire2197  &  (~ wire2235)  &  (~ wire2236) ) ;
 assign n_n4168 = ( wire7257 ) | ( n_n3118  &  (~ n_n3857)  &  n_n3135 ) | ( n_n3118  &  n_n3857  &  (~ n_n3135) ) ;
 assign n_n4084 = ( wire7149 ) | ( n_n3844  &  nrq5_5 ) | ( n_n3844  &  nrq5_2 ) ;
 assign n_n4082 = ( n_n3974  &  n_n3925 ) | ( n_n3974  &  wire1983 ) | ( n_n3925  &  wire1983 ) | ( n_n3974  &  wire7170 ) | ( n_n3925  &  wire7170 ) ;
 assign n_n3099 = ( n_n4004  &  n_n3961 ) | ( n_n4004  &  n_n4126 ) | ( n_n4004  &  (~ n_n4060) ) | ( (~ n_n4004)  &  (~ n_n3961)  &  (~ n_n4126)  &  n_n4060 ) ;
 assign n_n3920 = ( wire6936 ) | ( n_n4220  &  nrq5_5 ) | ( n_n4220  &  nrq5_2 ) ;
 assign n_n4211 = ( wire6939 ) | ( n_n4206  &  nrq5_5 ) | ( n_n4206  &  nrq5_2 ) ;
 assign wire838 = ( n_n4171 ) | ( n_n4036 ) | ( wire918 ) ;
 assign wire940 = ( n_n4171 ) | ( n_n4212 ) | ( n_n4036 ) | ( wire918 ) ;
 assign n_n4151 = ( wire6942 ) | ( n_n4132  &  nrq5_5 ) | ( n_n4132  &  nrq5_2 ) ;
 assign wire869 = ( (~ n_n4189)  &  n_n4184  &  (~ wire883) ) | ( (~ n_n4189)  &  n_n4184  &  n_n3892 ) | ( n_n4189  &  (~ n_n4184)  &  n_n3892 ) | ( (~ n_n4184)  &  wire883  &  (~ n_n3892) ) | ( n_n4184  &  (~ wire883)  &  (~ n_n3892) ) ;
 assign n_n4017 = ( n_n3996  &  n_n3888 ) | ( n_n3996  &  wire2017 ) | ( n_n3888  &  wire2017 ) | ( n_n3996  &  wire7152 ) | ( n_n3888  &  wire7152 ) ;
 assign n_n4219 = ( wire7152 ) | ( n_n4224  &  nrq5_5 ) | ( n_n4224  &  nrq5_2 ) ;
 assign n_n3888 = ( n_n3992  &  n_n3991 ) | ( n_n3992  &  wire1999 ) | ( n_n3991  &  wire1999 ) | ( n_n3992  &  wire7164 ) | ( n_n3991  &  wire7164 ) ;
 assign wire870 = ( (~ n_n4051)  &  wire2195 ) | ( (~ n_n4051)  &  wire7012 ) | ( (~ n_n4051)  &  wire7013 ) | ( n_n4051  &  (~ wire2195)  &  (~ wire7012)  &  (~ wire7013) ) ;
 assign n_n3746 = ( (~ wire844)  &  (~ n_n4052)  &  n_n3748 ) | ( n_n4052  &  (~ n_n3729)  &  n_n3748 ) | ( wire844  &  (~ n_n4052)  &  (~ n_n3748) ) | ( n_n4052  &  n_n3729  &  (~ n_n3748) ) ;
 assign n_n4245 = ( wire6945 ) | ( n_n4242  &  nrq5_5 ) | ( n_n4242  &  nrq5_2 ) ;
 assign n_n3643 = ( wire6948 ) | ( n_n4237  &  nrq5_5 ) | ( n_n4237  &  nrq5_2 ) ;
 assign n_n3142 = ( n_n3340  &  n_n3283 ) | ( n_n3340  &  wire839 ) | ( (~ n_n3340)  &  (~ n_n3283)  &  (~ wire839) ) ;
 assign n_n3869 = ( wire6951 ) | ( n_n4179  &  nrq5_5 ) | ( n_n4179  &  nrq5_2 ) ;
 assign wire917 = ( (~ preset_0_0_) ) | ( pdn ) | ( nlc1_2 ) ;
 assign n_n3925 = ( n_n4018  &  n_n4017 ) | ( n_n4018  &  wire1990 ) | ( n_n4017  &  wire1990 ) | ( n_n4018  &  wire7167 ) | ( n_n4017  &  wire7167 ) ;
 assign n_n4019 = ( wire7167 ) | ( n_n3890  &  nrq5_5 ) | ( n_n3890  &  nrq5_2 ) ;
 assign wire907 = ( n_n4019 ) | ( n_n3996  &  n_n4219 ) | ( n_n3996  &  n_n3888 ) | ( n_n4219  &  n_n3888 ) ;
 assign n_n3966 = ( wire7155 ) | ( n_n3971  &  nrq5_5 ) | ( n_n3971  &  nrq5_2 ) ;
 assign n_n3837 = ( wire7158 ) | ( n_n3500  &  nrq5_5 ) | ( n_n3500  &  nrq5_2 ) ;
 assign n_n3991 = ( n_n4027  &  n_n3837 ) | ( n_n3965  &  n_n4027  &  n_n3966 ) | ( n_n3965  &  n_n3966  &  n_n3837 ) ;
 assign n_n4196 = ( n_n3912  &  n_n3403 ) | ( n_n3912  &  wire1366 ) | ( n_n3403  &  wire1366 ) | ( n_n3912  &  wire7384 ) | ( n_n3403  &  wire7384 ) ;
 assign n_n4198 = ( wire7387 ) | ( n_n3470  &  nrq5_5 ) | ( n_n3470  &  nrq5_2 ) ;
 assign nak3_9 = ( wire7456 ) | ( wire989  &  wire7454 ) | ( wire989  &  wire7455 ) ;
 assign n_n4146 = ( wire7381 ) | ( n_n3810  &  nrq5_5 ) | ( n_n3810  &  nrq5_2 ) ;
 assign n_n3403 = ( n_n4145  &  n_n4144 ) | ( n_n4145  &  wire1361 ) | ( n_n4144  &  wire1361 ) | ( n_n4145  &  wire7381 ) | ( n_n4144  &  wire7381 ) ;
 assign n_n4253 = ( preset_0_0_  &  (~ nlc1_2) ) | ( nlc1_2  &  (~ n_n3998) ) ;
 assign n_n4069 = ( wire7384 ) | ( n_n4140  &  nrq5_5 ) | ( n_n4140  &  nrq5_2 ) ;
 assign n_n4115 = ( wire6954 ) | ( n_n4120  &  nrq5_5 ) | ( n_n4120  &  nrq5_2 ) ;
 assign n_n3565 = ( wire6957 ) | ( n_n4194  &  nrq5_5 ) | ( n_n4194  &  nrq5_2 ) ;
 assign n_n4178 = ( wire7170 ) | ( n_n4183  &  nrq5_5 ) | ( n_n4183  &  nrq5_2 ) ;
 assign n_n4125 = ( wire6960 ) | ( n_n4057  &  nrq5_5 ) | ( n_n4057  &  nrq5_2 ) ;
 assign wire841 = ( n_n4197  &  n_n4196  &  n_n4228 ) | ( n_n4197  &  n_n4198  &  n_n4228 ) | ( n_n4196  &  n_n4198  &  n_n4228 ) | ( (~ n_n4197)  &  (~ n_n4196)  &  (~ n_n4228) ) | ( (~ n_n4197)  &  (~ n_n4198)  &  (~ n_n4228) ) | ( (~ n_n4196)  &  (~ n_n4198)  &  (~ n_n4228) ) ;
 assign n_n3993 = ( wire7164 ) | ( n_n4086  &  nrq5_5 ) | ( n_n4086  &  nrq5_2 ) ;
 assign n_n3833 = ( (~ n_n4214)  &  n_n3460  &  (~ n_n3549)  &  wire955 ) ;
 assign n_n3549 = ( (~ n_n3838)  &  n_n3999 ) | ( wire6973  &  wire6974 ) ;
 assign n_n3903 = ( (~ n_n3575)  &  n_n4214  &  n_n3462 ) ;
 assign n_n3439 = ( (~ n_n3578)  &  (~ n_n3460) ) | ( (~ n_n3578)  &  wire2075 ) ;
 assign nrq5_5 = ( (~ nsr5_4)  &  nsr5_5 ) ;
 assign nrq5_2 = ( ndn3_8  &  (~ nlak3_9)  &  nsr3_9  &  nsr5_2 ) ;
 assign n_n4228 = ( wire7500 ) | ( n_n4095  &  nrq5_5 ) | ( n_n4095  &  nrq5_2 ) ;
 assign n_n3359 = ( wire945  &  n_n3434  &  wire948  &  wire952 ) ;
 assign wire945 = ( (~ n_n3700)  &  (~ n_n3701) ) | ( (~ n_n3701)  &  (~ nrq5_9) ) | ( (~ n_n3700)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign n_n3404 = ( wire945  &  (~ n_n3434) ) | ( wire945  &  (~ wire948) ) | ( wire945  &  (~ wire952) ) | ( (~ wire945)  &  n_n3434  &  wire948  &  wire952 ) ;
 assign n_n3779 = ( wire2207 ) | ( wire2208 ) | ( wire2209 ) | ( wire2210 ) ;
 assign wire877 = ( wire2211 ) | ( (~ ndn5_10)  &  n_n4183  &  (~ nsr5_7) ) ;
 assign n_n4129 = ( wire7186 ) | ( n_n3404  &  wire7183 ) | ( n_n3404  &  wire7184 ) ;
 assign wire878 = ( wire1929 ) | ( n_n3844  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign n_n4189 = ( (~ n_n4129)  &  wire878 ) | ( n_n4129  &  wire1937 ) | ( n_n4129  &  wire1938 ) ;
 assign nrq5_9 = ( nen5_9  &  (~ ndn5_9) ) ;
 assign wire809 = ( (~ nen5_9)  &  ndn5_10 ) | ( ndn5_9  &  ndn5_10 ) | ( (~ nen5_9)  &  nsr5_7 ) | ( ndn5_9  &  nsr5_7 ) ;
 assign wire879 = ( wire1737 ) | ( n_n3810  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire923 = ( (~ n_n3810) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n4184 = ( wire1733 ) | ( wire1734 ) | ( wire1735 ) | ( wire1736 ) ;
 assign n_n3118 = ( wire916  &  wire7223 ) | ( wire916  &  wire7224 ) | ( wire880  &  (~ wire7223)  &  (~ wire7224) ) ;
 assign n_n3857 = ( wire890  &  (~ n_n3484) ) | ( n_n3484  &  wire1729 ) | ( n_n3484  &  wire1730 ) ;
 assign n_n3135 = ( wire7244 ) | ( (~ n_n4160)  &  (~ wire934) ) | ( (~ n_n4160)  &  wire7241 ) ;
 assign wire880 = ( wire1754 ) | ( n_n3470  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire916 = ( wire809 ) | ( wire1751 ) | ( wire1752 ) ;
 assign wire955 = ( nrq5_5 ) | ( nrq5_2 ) | ( wire7125 ) | ( wire7126 ) ;
 assign wire926 = ( (~ n_n3844) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign ndn_latch5_5 = ( (~ ndn5_5)  &  (~ nsr5_5) ) ;
 assign nrq5_6 = ( ndn3_8  &  (~ ndn5_6)  &  (~ nlak3_9)  &  nsr3_9 ) ;
 assign wire844 = ( wire1500 ) | ( n_n4194  &  nrq5_6 ) ;
 assign n_n4052 = ( wire1495 ) | ( wire7316 ) | ( wire7317 ) | ( wire7318 ) ;
 assign n_n3363 = ( wire1631 ) | ( wire7288 ) | ( wire7289 ) | ( wire7290 ) ;
 assign wire845 = ( wire1636 ) | ( n_n4070  &  nrq5_6 ) ;
 assign n_n3729 = ( (~ n_n3363)  &  wire845 ) | ( n_n3363  &  wire1638 ) | ( n_n3363  &  wire1639 ) ;
 assign nrq2_2 = ( preset_0_0_  &  (~ pdn)  &  (~ nlc1_2)  &  (~ ndn2_2) ) ;
 assign ndn_latch5_3 = ( (~ ndn5_3)  &  (~ nsr5_3) ) ;
 assign ndn_latch5_8 = ( (~ ndn5_8)  &  (~ nsr5_8) ) ;
 assign wire946 = ( (~ n_n3585)  &  (~ n_n3100) ) | ( (~ n_n3100)  &  (~ nrq5_9) ) | ( (~ n_n3585)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign wire947 = ( (~ n_n3736)  &  (~ n_n3735) ) | ( (~ n_n3736)  &  (~ nrq5_9) ) | ( (~ n_n3735)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign ndn_latch5_2 = ( (~ ndn5_2)  &  (~ nsr5_2) ) ;
 assign wire883 = ( wire1915 ) | ( n_n4136  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign n_n3892 = ( wire7191 ) | ( wire7192 ) ;
 assign nrq5_10 = ( (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign ndn_latch5_4 = ( (~ ndn5_4)  &  (~ nsr5_4) ) ;
 assign ndn_latch5_7 = ( (~ ndn5_7)  &  (~ nsr5_7) ) ;
 assign n_n4123 = ( n_n3359  &  wire946  &  wire947  &  wire953 ) ;
 assign wire914 = ( (~ n_n3482) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n4160 = ( wire1721 ) | ( wire1722 ) | ( wire1723 ) | ( wire7236 ) ;
 assign n_n3532 = ( wire2096 ) | ( wire7026 ) | ( wire7027 ) | ( wire7028 ) ;
 assign wire846 = ( wire2101 ) | ( n_n3813  &  nrq5_6 ) ;
 assign n_n3236 = ( (~ n_n3532)  &  wire846 ) | ( n_n3532  &  wire2103 ) | ( n_n3532  &  wire2104 ) ;
 assign n_n3434 = ( (~ n_n3976)  &  wire949  &  wire950  &  wire951 ) ;
 assign wire948 = ( (~ n_n3679)  &  (~ n_n4021) ) | ( (~ n_n3679)  &  (~ nrq5_9) ) | ( (~ n_n4021)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign n_n3281 = ( wire7002 ) | ( n_n4200  &  wire6999 ) | ( n_n4200  &  wire7000 ) ;
 assign wire886 = ( wire2181 ) | ( n_n4224  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign n_n4202 = ( (~ n_n3281)  &  wire886 ) | ( n_n3281  &  wire2185 ) | ( n_n3281  &  wire2186 ) ;
 assign n_n3897 = ( (~ n_n3434)  &  wire948 ) | ( n_n3434  &  (~ wire948) ) ;
 assign n_n3883 = ( (~ n_n3513)  &  n_n3581 ) | ( n_n3818  &  n_n3581 ) | ( (~ n_n3513)  &  n_n3818  &  n_n3512 ) ;
 assign wire818 = ( n_n3513  &  n_n3512 ) | ( (~ n_n3818)  &  n_n3512 ) | ( n_n3513  &  (~ n_n3818)  &  n_n3581 ) ;
 assign wire989 = ( (~ n_n3882)  &  wire818 ) | ( n_n3884  &  wire818 ) | ( (~ n_n3882)  &  n_n3884  &  n_n3883 ) ;
 assign n_n3762 = ( wire1316 ) | ( wire7433 ) | ( wire7437 ) ;
 assign n_n3396 = ( wire1308 ) | ( wire929  &  (~ wire7436)  &  (~ wire7437) ) ;
 assign wire939 = ( (~ n_n3489) ) | ( n_n4054 ) ;
 assign wire975 = ( n_n3908 ) | ( (~ n_n4015) ) ;
 assign n_n3581 = ( wire1302 ) | ( wire1303 ) | ( wire1304 ) | ( wire7443 ) ;
 assign wire843 = ( n_n4243 ) | ( (~ n_n3862) ) ;
 assign wire929 = ( wire1317 ) | ( wire7423 ) | ( wire7424 ) | ( (~ wire7423)  &  (~ wire7424) ) ;
 assign n_n3950 = ( wire2046 ) | ( wire7141 ) | ( wire7142 ) | ( wire7143 ) ;
 assign n_n3976 = ( wire2236 ) | ( nen5_9  &  (~ ndn5_9)  &  n_n3625 ) ;
 assign wire949 = ( (~ n_n3968)  &  (~ n_n3959) ) | ( (~ n_n3968)  &  (~ nrq5_9) ) | ( (~ n_n3959)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign wire950 = ( (~ n_n3799)  &  (~ n_n4024) ) | ( (~ n_n3799)  &  (~ nrq5_9) ) | ( (~ n_n4024)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign wire951 = ( (~ n_n3957)  &  (~ n_n3205) ) | ( (~ n_n3205)  &  (~ nrq5_9) ) | ( (~ n_n3957)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign n_n3521 = ( (~ wire949)  &  wire950 ) | ( wire950  &  wire2235 ) | ( wire950  &  wire2236 ) | ( wire949  &  (~ wire950)  &  (~ wire2235)  &  (~ wire2236) ) ;
 assign n_n4200 = ( n_n3976  &  wire951 ) | ( (~ wire949)  &  wire951 ) | ( (~ wire950)  &  wire951 ) | ( (~ n_n3976)  &  wire949  &  wire950  &  (~ wire951) ) ;
 assign n_n3569 = ( wire2140 ) | ( wire7082 ) | ( wire7083 ) | ( wire7084 ) ;
 assign n_n3111 = ( wire2085 ) | ( wire7118 ) | ( wire7119 ) | ( wire7120 ) ;
 assign wire849 = ( wire2090 ) | ( n_n4132  &  nrq5_6 ) ;
 assign n_n3025 = ( wire2129 ) | ( wire7068 ) | ( wire7069 ) | ( wire7070 ) ;
 assign wire850 = ( wire2134 ) | ( n_n3924  &  nrq5_6 ) ;
 assign n_n3955 = ( (~ n_n3025)  &  wire850 ) | ( n_n3025  &  wire2136 ) | ( n_n3025  &  wire2137 ) ;
 assign n_n4248 = ( (~ n_n3359)  &  wire953 ) | ( (~ wire946)  &  wire953 ) | ( (~ wire947)  &  wire953 ) | ( n_n3359  &  wire946  &  wire947  &  (~ wire953) ) ;
 assign wire890 = ( wire1745 ) | ( n_n4140  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire930 = ( (~ n_n4140) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n3484 = ( wire7250 ) | ( n_n4248  &  wire7247 ) | ( n_n4248  &  wire7248 ) ;
 assign wire931 = ( ndn5_10 ) | ( (~ n_n4183) ) | ( nsr5_7 ) ;
 assign wire952 = ( (~ n_n3203)  &  (~ n_n3081) ) | ( (~ n_n3203)  &  (~ nrq5_9) ) | ( (~ n_n3081)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign wire932 = ( (~ n_n3890) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n4062 = ( wire2172 ) | ( wire6996 ) | ( wire6997 ) ;
 assign n_n3512 = ( wire1297 ) | ( n_n3762  &  (~ n_n3581) ) | ( n_n3396  &  (~ n_n3581) ) ;
 assign wire953 = ( (~ n_n4042)  &  (~ n_n3824) ) | ( (~ n_n4042)  &  (~ nrq5_9) ) | ( (~ n_n3824)  &  (~ nrq5_10) ) | ( (~ nrq5_9)  &  (~ nrq5_10) ) ;
 assign wire933 = ( (~ n_n4224) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n3543 = ( wire2118 ) | ( wire7054 ) | ( wire7055 ) | ( wire7056 ) ;
 assign wire851 = ( wire2123 ) | ( n_n3868  &  nrq5_6 ) ;
 assign n_n4051 = ( wire2196  &  wire2235 ) | ( wire2197  &  wire2235 ) | ( wire2196  &  wire2236 ) | ( wire2197  &  wire2236 ) ;
 assign wire934 = ( (~ n_n4095) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign n_n4153 = ( wire2160 ) | ( wire7108 ) | ( nrq5_6  &  wire7102 ) ;
 assign wire852 = ( wire2156 ) | ( n_n4120  &  nrq5_6 ) ;
 assign n_n3035 = ( wire2151 ) | ( wire7096 ) | ( wire7097 ) | ( wire7098 ) ;
 assign n_n3635 = ( wire2107 ) | ( wire7040 ) | ( wire7041 ) | ( wire7042 ) ;
 assign n_n3748 = ( wire7333 ) | ( wire7334 ) | ( wire7335 ) | ( wire7336 ) ;
 assign wire935 = ( (~ n_n4086) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign wire817 = ( n_n3513 ) | ( (~ n_n3818) ) ;
 assign wire936 = ( (~ n_n3500) ) | ( ndn5_10 ) | ( nsr5_7 ) ;
 assign wire835 = ( (~ n_n3811)  &  nsr3_2 ) | ( nsr3_2  &  n_n4253 ) | ( nsr3_2  &  (~ wire7467) ) ;
 assign wire876 = ( (~ n_n4214)  &  n_n3462 ) | ( n_n3462  &  n_n3142 ) | ( n_n3462  &  (~ wire7205) ) ;
 assign wire938 = ( wire816  &  (~ n_n3281)  &  wire2185 ) | ( wire816  &  (~ n_n3281)  &  wire2186 ) | ( wire816  &  n_n3281  &  (~ wire2185)  &  (~ wire2186) ) ;
 assign wire954 = ( (~ preset)  &  ndn5_10  &  n_n3829 ) | ( (~ preset)  &  n_n3829  &  nsr5_7 ) ;
 assign wire963 = ( n_n3833  &  (~ n_n3439)  &  wire7518 ) | ( n_n3903  &  (~ n_n3439)  &  wire7518 ) ;
 assign wire964 = ( n_n3833  &  wire7521 ) | ( n_n3903  &  wire7521 ) | ( n_n3439  &  wire7521 ) ;
 assign wire970 = ( wire802  &  (~ n_n3025)  &  wire2136 ) | ( wire802  &  (~ n_n3025)  &  wire2137 ) | ( wire802  &  n_n3025  &  (~ wire2136)  &  (~ wire2137) ) ;
 assign wire971 = ( (~ preset)  &  (~ nen5_9)  &  n_n3475 ) | ( (~ preset)  &  ndn5_9  &  n_n3475 ) ;
 assign wire972 = ( (~ preset)  &  (~ ndn5_9)  &  n_n4068 ) | ( (~ preset)  &  nld3_9  &  n_n4068 ) ;
 assign wire973 = ( (~ preset)  &  n_n3821  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire976 = ( (~ preset)  &  nld3_9  &  n_n3336 ) ;
 assign wire977 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3373 ) ;
 assign wire979 = ( (~ preset)  &  ndn5_4  &  n_n4047 ) | ( (~ preset)  &  n_n4047  &  nsr5_4 ) ;
 assign wire980 = ( (~ preset)  &  ndn5_8  &  n_n3959 ) | ( (~ preset)  &  n_n3959  &  nsr5_8 ) ;
 assign wire983 = ( (~ preset)  &  ndn5_4  &  n_n3367 ) | ( (~ preset)  &  n_n3367  &  nsr5_4 ) ;
 assign wire985 = ( (~ preset)  &  ndn5_4  &  n_n3303 ) | ( (~ preset)  &  n_n3303  &  nsr5_4 ) ;
 assign wire987 = ( (~ preset)  &  n_n3420  &  nld3_9 ) ;
 assign wire988 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3393 ) ;
 assign wire991 = ( (~ preset)  &  n_n3791  &  nld3_9 ) ;
 assign wire992 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3533 ) ;
 assign wire993 = ( (~ preset)  &  ndn5_2  &  n_n3663 ) | ( (~ preset)  &  n_n3663  &  nsr5_2 ) ;
 assign wire996 = ( (~ preset)  &  ndn5_5  &  n_n3607 ) | ( (~ preset)  &  n_n3607  &  nsr5_5 ) ;
 assign wire998 = ( (~ preset)  &  ndn5_10  &  n_n3274 ) | ( (~ preset)  &  n_n3274  &  nsr5_7 ) ;
 assign wire999 = ( pdxport_11_11_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1000 = ( (~ preset)  &  ndn3_3  &  n_n4237 ) | ( (~ preset)  &  n_n4237  &  nsr3_2 ) ;
 assign wire1002 = ( (~ preset)  &  n_n3677  &  nld3_9 ) ;
 assign wire1003 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3741  &  ndn3_3 ) ;
 assign wire1007 = ( (~ preset)  &  n_n4000  &  wire1008  &  wire7129 ) ;
 assign wire1008 = ( (~ n_n4214)  &  n_n3462 ) | ( n_n3462  &  n_n3142 ) | ( n_n3462  &  (~ wire7205) ) ;
 assign wire1017 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3002 ) | ( (~ preset)  &  nld3_9  &  n_n3002 ) ;
 assign wire1018 = ( (~ preset)  &  ndn5_9  &  n_n3212  &  (~ nld3_9) ) ;
 assign wire1020 = ( (~ preset)  &  ndn3_3  &  n_n3876 ) | ( (~ preset)  &  n_n3876  &  nsr3_2 ) ;
 assign wire1023 = ( (~ preset)  &  ndn5_7  &  n_n3701 ) | ( (~ preset)  &  n_n3701  &  nsr5_7 ) ;
 assign wire1026 = ( (~ preset)  &  ndn3_3  &  n_n3681 ) | ( (~ preset)  &  n_n3681  &  nsr3_2 ) ;
 assign wire1032 = ( (~ preset)  &  n_n3903  &  wire7506 ) ;
 assign wire1034 = ( (~ preset)  &  n_n3992  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1037 = ( (~ preset)  &  n_n4227  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1041 = ( n_n4237  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1042 = ( n_n3445  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1043 = ( n_n3905  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1044 = ( n_n3663  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1045 = ( wire811  &  (~ n_n3025)  &  wire2136 ) | ( wire811  &  (~ n_n3025)  &  wire2137 ) | ( wire811  &  n_n3025  &  (~ wire2136)  &  (~ wire2137) ) ;
 assign wire1049 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3493 ) | ( (~ preset)  &  nld3_9  &  n_n3493 ) ;
 assign wire1050 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3442 ) ;
 assign wire1052 = ( (~ preset)  &  ndn3_3  &  n_n3580 ) | ( (~ preset)  &  n_n3580  &  nsr3_2 ) ;
 assign wire1056 = ( (~ preset)  &  n_n3761  &  nld3_9 ) ;
 assign wire1057 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3248  &  ndn3_3 ) ;
 assign wire1058 = ( (~ preset)  &  n_n3826  &  ndn5_10 ) | ( (~ preset)  &  n_n3826  &  nsr5_7 ) ;
 assign wire1060 = ( pdxport_7_7_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1061 = ( (~ preset)  &  ndn3_3  &  n_n4132 ) | ( (~ preset)  &  n_n4132  &  nsr3_2 ) ;
 assign wire1062 = ( (~ preset)  &  (~ ndn5_9)  &  n_n2968 ) | ( (~ preset)  &  nld3_9  &  n_n2968 ) ;
 assign wire1063 = ( (~ preset)  &  ndn5_9  &  n_n3774  &  (~ nld3_9) ) ;
 assign wire1064 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3067 ) | ( (~ preset)  &  nld3_9  &  n_n3067 ) ;
 assign wire1065 = ( (~ preset)  &  ndn5_9  &  n_n3513  &  (~ nld3_9) ) ;
 assign wire1067 = ( (~ preset)  &  ndn3_3  &  n_n3393 ) | ( (~ preset)  &  n_n3393  &  nsr3_2 ) ;
 assign wire1071 = ( (~ preset)  &  n_n3884  &  (~ nrq5_6) ) ;
 assign wire1073 = ( (~ preset)  &  ndn3_3  &  n_n3533 ) | ( (~ preset)  &  n_n3533  &  nsr3_2 ) ;
 assign wire1076 = ( (~ preset)  &  ndn5_7  &  n_n3968 ) | ( (~ preset)  &  n_n3968  &  nsr5_7 ) ;
 assign wire1078 = ( (~ preset)  &  ndn5_3  &  n_n3436 ) | ( (~ preset)  &  n_n3436  &  nsr5_3 ) ;
 assign wire1081 = ( (~ preset)  &  ndn5_4  &  n_n4045 ) | ( (~ preset)  &  n_n4045  &  nsr5_4 ) ;
 assign wire1084 = ( (~ preset)  &  ndn5_2  &  n_n3323 ) | ( (~ preset)  &  n_n3323  &  nsr5_2 ) ;
 assign wire1086 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3689 ) | ( (~ preset)  &  nld3_9  &  n_n3689 ) ;
 assign wire1087 = ( (~ preset)  &  ndn5_9  &  n_n4158  &  (~ nld3_9) ) ;
 assign wire1089 = ( (~ preset)  &  ndn3_3  &  n_n3417 ) | ( (~ preset)  &  n_n3417  &  nsr3_2 ) ;
 assign wire1093 = ( (~ preset)  &  ndn3_3  &  n_n4218 ) | ( (~ preset)  &  n_n4218  &  nsr3_2 ) ;
 assign wire1097 = ( (~ preset)  &  ndn5_5  &  n_n3793 ) | ( (~ preset)  &  n_n3793  &  nsr5_5 ) ;
 assign wire1098 = ( paport_8_8_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1099 = ( (~ preset)  &  ndn3_3  &  n_n4015 ) | ( (~ preset)  &  n_n4015  &  nsr3_2 ) ;
 assign wire1104 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3122 ) | ( (~ preset)  &  nld3_9  &  n_n3122 ) ;
 assign wire1105 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3475 ) ;
 assign wire1106 = ( (~ preset)  &  ndn5_8  &  n_n3735 ) | ( (~ preset)  &  n_n3735  &  nsr5_8 ) ;
 assign wire1108 = ( (~ preset)  &  ndn5_8  &  n_n4024 ) | ( (~ preset)  &  n_n4024  &  nsr5_8 ) ;
 assign wire1110 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3563 ) | ( (~ preset)  &  nld3_9  &  n_n3563 ) ;
 assign wire1111 = ( (~ preset)  &  n_n3832  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1114 = ( n_n4125  &  wire2071 ) | ( (~ preset)  &  n_n4125  &  n_n3833 ) ;
 assign wire1115 = ( n_n4126  &  wire2073 ) | ( n_n4126  &  wire2074 ) ;
 assign wire1117 = ( (~ preset)  &  ndn3_3  &  n_n3786 ) | ( (~ preset)  &  n_n3786  &  nsr3_2 ) ;
 assign wire1120 = ( (~ preset)  &  ndn5_3  &  n_n3806 ) | ( (~ preset)  &  n_n3806  &  nsr5_3 ) ;
 assign wire1124 = ( wire802  &  (~ n_n3281)  &  wire2185 ) | ( wire802  &  (~ n_n3281)  &  wire2186 ) | ( wire802  &  n_n3281  &  (~ wire2185)  &  (~ wire2186) ) ;
 assign wire1125 = ( (~ preset)  &  (~ nen5_9)  &  n_n3442 ) | ( (~ preset)  &  ndn5_9  &  n_n3442 ) ;
 assign wire1129 = ( (~ preset)  &  (~ nen5_9)  &  n_n3464 ) | ( (~ preset)  &  ndn5_9  &  n_n3464 ) ;
 assign wire1131 = ( (~ preset)  &  n_n3179  &  nld3_9 ) ;
 assign wire1132 = ( (~ preset)  &  (~ ndn3_8)  &  n_n4232  &  ndn3_3 ) ;
 assign wire1133 = ( wire816  &  (~ n_n3484)  &  wire1729 ) | ( wire816  &  (~ n_n3484)  &  wire1730 ) | ( wire816  &  n_n3484  &  (~ wire1729)  &  (~ wire1730) ) ;
 assign wire1134 = ( (~ preset)  &  n_n3788  &  ndn5_10 ) | ( (~ preset)  &  n_n3788  &  nsr5_7 ) ;
 assign wire1136 = ( (~ preset)  &  n_n3535  &  nld3_9 ) ;
 assign wire1137 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3580 ) ;
 assign wire1138 = ( (~ preset)  &  n_n3824  &  ndn5_8 ) | ( (~ preset)  &  n_n3824  &  nsr5_8 ) ;
 assign wire1141 = ( (~ preset)  &  ndn3_3  &  n_n3541 ) | ( (~ preset)  &  n_n3541  &  nsr3_2 ) ;
 assign wire1145 = ( (~ preset)  &  n_n3821  &  nld3_9 ) ;
 assign wire1146 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3822  &  ndn3_3 ) ;
 assign wire1147 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3199 ) | ( (~ preset)  &  nld3_9  &  n_n3199 ) ;
 assign wire1148 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3981 ) ;
 assign wire1151 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3887 ) | ( (~ preset)  &  nld3_9  &  n_n3887 ) ;
 assign wire1152 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3884 ) ;
 assign wire1153 = ( n_n4018  &  n_n4017  &  wire7486 ) | ( n_n4018  &  n_n4019  &  wire7486 ) | ( n_n4017  &  n_n4019  &  wire7486 ) ;
 assign wire1154 = ( (~ n_n3974)  &  wire813  &  (~ n_n3925)  &  n_n4178 ) | ( (~ n_n3974)  &  wire813  &  n_n3925  &  (~ n_n4178) ) ;
 assign wire1155 = ( n_n3974  &  wire797  &  (~ n_n3925)  &  (~ n_n4178) ) ;
 assign wire1156 = ( (~ preset)  &  n_n3974  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1157 = ( wire811  &  (~ n_n3532)  &  wire2103 ) | ( wire811  &  (~ n_n3532)  &  wire2104 ) | ( wire811  &  n_n3532  &  (~ wire2103)  &  (~ wire2104) ) ;
 assign wire1159 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3024 ) | ( (~ preset)  &  nld3_9  &  n_n3024 ) ;
 assign wire1160 = ( (~ preset)  &  n_n3715  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1161 = ( paport_11_11_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1162 = ( (~ preset)  &  ndn3_3  &  n_n4205 ) | ( (~ preset)  &  n_n4205  &  nsr3_2 ) ;
 assign wire1163 = ( (~ preset)  &  n_n4167  &  ndn5_10 ) | ( (~ preset)  &  n_n4167  &  nsr5_7 ) ;
 assign wire1166 = ( (~ preset)  &  ndn3_3  &  n_n3866 ) | ( (~ preset)  &  n_n3866  &  nsr3_2 ) ;
 assign wire1169 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3901 ) | ( (~ preset)  &  nld3_9  &  n_n3901 ) ;
 assign wire1170 = ( (~ preset)  &  ndn5_9  &  n_n3931  &  (~ nld3_9) ) ;
 assign wire1174 = ( (~ preset)  &  (~ nen5_9)  &  n_n3743 ) | ( (~ preset)  &  ndn5_9  &  n_n3743 ) ;
 assign wire1176 = ( (~ preset)  &  ndn3_3  &  n_n4080 ) | ( (~ preset)  &  n_n4080  &  nsr3_2 ) ;
 assign wire1179 = ( pdxport_0_0_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1180 = ( (~ preset)  &  ndn3_3  &  n_n3906 ) | ( (~ preset)  &  n_n3906  &  nsr3_2 ) ;
 assign wire1184 = ( (~ preset)  &  ndn5_4  &  n_n3840 ) | ( (~ preset)  &  n_n3840  &  nsr5_4 ) ;
 assign wire1187 = ( n_n3565  &  wire2071 ) | ( (~ preset)  &  n_n3565  &  n_n3833 ) ;
 assign wire1188 = ( n_n3283  &  wire2073 ) | ( n_n3283  &  wire2074 ) ;
 assign wire1190 = ( (~ preset)  &  ndn3_3  &  n_n3196 ) | ( (~ preset)  &  n_n3196  &  nsr3_2 ) ;
 assign wire1194 = ( (~ preset)  &  n_n3713  &  nld3_9 ) ;
 assign wire1195 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3235  &  ndn3_3 ) ;
 assign wire1197 = ( (~ preset)  &  ndn3_3  &  n_n3105 ) | ( (~ preset)  &  n_n3105  &  nsr3_2 ) ;
 assign wire1200 = ( (~ preset)  &  n_n4221  &  ndn5_2 ) | ( (~ preset)  &  n_n4221  &  nsr5_2 ) ;
 assign wire1203 = ( (~ preset)  &  n_n4158  &  nld3_9 ) ;
 assign wire1204 = ( (~ preset)  &  (~ ndn3_8)  &  n_n4159  &  ndn3_3 ) ;
 assign wire1205 = ( (~ preset)  &  n_n3081  &  ndn5_8 ) | ( (~ preset)  &  n_n3081  &  nsr5_8 ) ;
 assign wire1208 = ( (~ preset)  &  ndn5_4  &  n_n3424 ) | ( (~ preset)  &  n_n3424  &  nsr5_4 ) ;
 assign wire1210 = ( (~ preset)  &  ndn5_5  &  n_n4236 ) | ( (~ preset)  &  n_n4236  &  nsr5_5 ) ;
 assign wire1213 = ( n_n4115  &  wire2071 ) | ( (~ preset)  &  n_n4115  &  n_n3833 ) ;
 assign wire1214 = ( n_n3961  &  wire2073 ) | ( n_n3961  &  wire2074 ) ;
 assign wire1215 = ( n_n4145  &  n_n4144  &  wire7472 ) | ( n_n4145  &  n_n4146  &  wire7472 ) | ( n_n4144  &  n_n4146  &  wire7472 ) ;
 assign wire1216 = ( (~ n_n3912)  &  wire813  &  (~ n_n3403)  &  n_n4069 ) | ( (~ n_n3912)  &  wire813  &  n_n3403  &  (~ n_n4069) ) ;
 assign wire1217 = ( n_n3912  &  wire797  &  (~ n_n3403)  &  (~ n_n4069) ) ;
 assign wire1218 = ( (~ preset)  &  n_n3912  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1219 = ( (~ preset)  &  n_n4075  &  ndn5_8 ) | ( (~ preset)  &  n_n4075  &  nsr5_8 ) ;
 assign wire1221 = ( (~ preset)  &  n_n3612  &  ndn5_8 ) | ( (~ preset)  &  n_n3612  &  nsr5_8 ) ;
 assign wire1223 = ( (~ preset)  &  n_n3473  &  ndn5_2 ) | ( (~ preset)  &  n_n3473  &  nsr5_2 ) ;
 assign wire1226 = ( (~ preset)  &  n_n3908  &  nld3_9 ) ;
 assign wire1227 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3634  &  ndn3_3 ) ;
 assign wire1232 = ( paport_0_0_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1233 = ( (~ preset)  &  ndn3_3  &  n_n3916 ) | ( (~ preset)  &  n_n3916  &  nsr3_2 ) ;
 assign wire1235 = ( (~ preset)  &  ndn3_3  &  n_n3373 ) | ( (~ preset)  &  n_n3373  &  nsr3_2 ) ;
 assign wire1240 = ( (~ preset)  &  (~ ndn5_9)  &  n_n2995 ) | ( (~ preset)  &  n_n2995  &  nld3_9 ) ;
 assign wire1241 = ( (~ preset)  &  n_n3908  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1243 = ( (~ preset)  &  ndn3_3  &  n_n3716 ) | ( (~ preset)  &  n_n3716  &  nsr3_2 ) ;
 assign wire1246 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3628 ) | ( (~ preset)  &  n_n3628  &  nld3_9 ) ;
 assign wire1247 = ( (~ preset)  &  ndn5_9  &  n_n4111  &  (~ nld3_9) ) ;
 assign wire1248 = ( n_n3949  &  n_n3948  &  wire7462 ) | ( n_n3949  &  n_n4131  &  wire7462 ) | ( n_n3948  &  n_n4131  &  wire7462 ) ;
 assign wire1249 = ( (~ n_n4145)  &  (~ n_n4144)  &  wire813  &  n_n4146 ) | ( (~ n_n4145)  &  n_n4144  &  wire813  &  (~ n_n4146) ) ;
 assign wire1250 = ( n_n4145  &  wire797  &  (~ n_n4144)  &  (~ n_n4146) ) ;
 assign wire1251 = ( (~ preset)  &  n_n4145  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1253 = ( (~ preset)  &  n_n3212  &  nld3_9 ) ;
 assign wire1254 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3196 ) ;
 assign wire1256 = ( (~ preset)  &  ndn5_5  &  n_n3069 ) | ( (~ preset)  &  n_n3069  &  nsr5_5 ) ;
 assign wire1258 = ( (~ preset)  &  n_n3489  &  nld3_9 ) ;
 assign wire1259 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3105 ) ;
 assign wire1261 = ( (~ preset)  &  ndn5_5  &  n_n3143 ) | ( (~ preset)  &  n_n3143  &  nsr5_5 ) ;
 assign wire1262 = ( paport_9_9_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1263 = ( (~ preset)  &  ndn3_3  &  n_n3818 ) | ( (~ preset)  &  n_n3818  &  nsr3_2 ) ;
 assign wire1264 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3327 ) | ( (~ preset)  &  n_n3327  &  nld3_9 ) ;
 assign wire1265 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3743 ) ;
 assign wire1267 = ( (~ preset)  &  nld3_9  &  n_n3884 ) ;
 assign wire1268 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3011  &  ndn3_3 ) ;
 assign wire1270 = ( (~ preset)  &  ndn5_4  &  n_n3188 ) | ( (~ preset)  &  n_n3188  &  nsr5_4 ) ;
 assign wire1271 = ( (~ preset)  &  ndn5_7  &  n_n3100 ) | ( (~ preset)  &  n_n3100  &  nsr5_7 ) ;
 assign wire1273 = ( (~ preset)  &  ndn5_7  &  n_n3205 ) | ( (~ preset)  &  n_n3205  &  nsr5_7 ) ;
 assign wire1276 = ( (~ preset)  &  (~ nen5_9)  &  n_n4079 ) | ( (~ preset)  &  ndn5_9  &  n_n4079 ) ;
 assign wire1279 = ( (~ preset)  &  (~ nen5_9)  &  n_n3680 ) | ( (~ preset)  &  ndn5_9  &  n_n3680 ) ;
 assign wire1282 = ( (~ preset)  &  ndn5_5  &  n_n3630 ) | ( (~ preset)  &  n_n3630  &  nsr5_5 ) ;
 assign wire1286 = ( wire7447  &  wire7451 ) | ( n_n3512  &  (~ wire817)  &  wire7451 ) ;
 assign wire1297 = ( wire975  &  wire7438 ) | ( n_n3396  &  (~ wire939)  &  wire975 ) ;
 assign wire1302 = ( (~ n_n3396)  &  (~ wire7438)  &  wire7441 ) | ( wire939  &  (~ wire7438)  &  wire7441 ) ;
 assign wire1303 = ( (~ n_n3396)  &  (~ wire7438)  &  wire7442 ) | ( wire939  &  (~ wire7438)  &  wire7442 ) ;
 assign wire1304 = ( (~ wire975)  &  wire7438 ) | ( n_n3396  &  (~ wire939)  &  (~ wire975) ) ;
 assign wire1308 = ( wire7423  &  wire7425 ) | ( wire7424  &  wire7425 ) ;
 assign wire1312 = ( wire1317  &  wire7429 ) | ( (~ wire7423)  &  (~ wire7424)  &  wire7429 ) ;
 assign wire1313 = ( wire1317  &  wire7430 ) | ( (~ wire7423)  &  (~ wire7424)  &  wire7430 ) ;
 assign wire1314 = ( wire1317  &  wire7431 ) | ( (~ wire7423)  &  (~ wire7424)  &  wire7431 ) ;
 assign wire1315 = ( wire1317  &  wire7432 ) | ( (~ wire7423)  &  (~ wire7424)  &  wire7432 ) ;
 assign wire1316 = ( (~ wire843)  &  wire1317 ) | ( (~ wire843)  &  wire7423 ) | ( (~ wire843)  &  wire7424 ) | ( (~ wire843)  &  (~ wire7423)  &  (~ wire7424) ) ;
 assign wire1317 = ( wire7410  &  wire7428 ) | ( wire7411  &  wire7428 ) | ( wire7412  &  wire7428 ) ;
 assign wire1319 = ( wire7410  &  wire7414 ) | ( wire7411  &  wire7414 ) | ( wire7412  &  wire7414 ) ;
 assign wire1320 = ( wire7410  &  wire7415 ) | ( wire7411  &  wire7415 ) | ( wire7412  &  wire7415 ) ;
 assign wire1321 = ( (~ wire7410)  &  (~ wire7411)  &  (~ wire7412)  &  wire7416 ) ;
 assign wire1322 = ( (~ wire7410)  &  (~ wire7411)  &  (~ wire7412)  &  wire7417 ) ;
 assign wire1323 = ( (~ wire7410)  &  (~ wire7411)  &  (~ wire7412)  &  wire7418 ) ;
 assign wire1324 = ( (~ wire7410)  &  (~ wire7411)  &  (~ wire7412)  &  wire7419 ) ;
 assign wire1327 = ( n_n3535  &  (~ n_n3916)  &  n_n3794 ) ;
 assign wire1328 = ( (~ n_n3797)  &  n_n4111  &  n_n3794 ) ;
 assign wire1338 = ( (~ preset)  &  ndn3_3  &  n_n3932 ) | ( (~ preset)  &  n_n3932  &  nsr3_2 ) ;
 assign wire1341 = ( (~ preset)  &  ndn5_7  &  n_n3626 ) | ( (~ preset)  &  n_n3626  &  nsr5_7 ) ;
 assign wire1344 = ( (~ preset)  &  n_n3680  &  nld3_9 ) ;
 assign wire1345 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3681 ) ;
 assign wire1346 = ( n_n3912  &  n_n3403  &  wire7389 ) | ( n_n3912  &  n_n4069  &  wire7389 ) | ( n_n3403  &  n_n4069  &  wire7389 ) ;
 assign wire1347 = ( (~ n_n4197)  &  wire813  &  (~ n_n4196)  &  n_n4198 ) | ( (~ n_n4197)  &  wire813  &  n_n4196  &  (~ n_n4198) ) ;
 assign wire1348 = ( n_n4197  &  wire797  &  (~ n_n4196)  &  (~ n_n4198) ) ;
 assign wire1349 = ( (~ preset)  &  n_n4197  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1352 = ( n_n3470  &  nrq5_2 ) | ( n_n3470  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1353 = ( n_n4194  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1354 = ( n_n3468  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1355 = ( n_n3469  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1356 = ( n_n3473  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1361 = ( n_n3810  &  nrq5_2 ) | ( n_n3810  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1362 = ( n_n4242  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1363 = ( n_n3426  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1364 = ( n_n3294  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1365 = ( n_n3293  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1366 = ( n_n4140  &  nrq5_2 ) | ( n_n4140  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1367 = ( n_n4070  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1368 = ( n_n4072  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1369 = ( n_n4073  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1370 = ( n_n4071  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1371 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3309 ) | ( (~ preset)  &  n_n3309  &  nld3_9 ) ;
 assign wire1372 = ( (~ preset)  &  n_n3516  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1373 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3694 ) | ( (~ preset)  &  n_n3694  &  nld3_9 ) ;
 assign wire1374 = ( (~ preset)  &  n_n4114  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1375 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3498 ) | ( (~ preset)  &  n_n3498  &  nld3_9 ) ;
 assign wire1376 = ( (~ preset)  &  n_n3791  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1378 = ( (~ preset)  &  n_n4114  &  nld3_9 ) ;
 assign wire1379 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3866 ) ;
 assign wire1381 = ( (~ preset)  &  ndn3_3  &  n_n4106 ) | ( (~ preset)  &  n_n4106  &  nsr3_2 ) ;
 assign wire1384 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3698 ) | ( (~ preset)  &  n_n3698  &  nld3_9 ) ;
 assign wire1385 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3336 ) ;
 assign wire1386 = ( wire2012  &  wire7370 ) | ( wire7158  &  wire7370 ) ;
 assign wire1387 = ( (~ wire1405)  &  (~ wire1406)  &  (~ wire1407)  &  wire7372 ) ;
 assign wire1388 = ( (~ preset)  &  n_n3903  &  wire7373 ) ;
 assign wire1390 = ( (~ preset)  &  n_n4027  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1391 = ( preset_0_0_  &  (~ preset)  &  (~ pdn)  &  (~ nlc1_2) ) ;
 assign wire1393 = ( (~ preset)  &  n_n4111  &  (~ nrq5_6) ) ;
 assign wire1395 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3728 ) | ( (~ preset)  &  n_n3728  &  nld3_9 ) ;
 assign wire1396 = ( (~ preset)  &  n_n3875  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1398 = ( (~ preset)  &  ndn5_5  &  n_n3910 ) | ( (~ preset)  &  n_n3910  &  nsr5_5 ) ;
 assign wire1401 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3767 ) | ( (~ preset)  &  n_n3767  &  nld3_9 ) ;
 assign wire1402 = ( (~ preset)  &  ndn5_9  &  n_n3214  &  (~ nld3_9) ) ;
 assign wire1403 = ( (~ preset)  &  n_n4021  &  ndn5_8 ) | ( (~ preset)  &  n_n4021  &  nsr5_8 ) ;
 assign wire1405 = ( (~ preset)  &  n_n3903  &  wire7365 ) ;
 assign wire1406 = ( n_n3965  &  wire797  &  (~ wire2007)  &  (~ wire7155) ) ;
 assign wire1407 = ( (~ preset)  &  n_n3965  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1408 = ( n_n3996  &  n_n4219  &  wire7360 ) | ( n_n3996  &  n_n3888  &  wire7360 ) | ( n_n4219  &  n_n3888  &  wire7360 ) ;
 assign wire1411 = ( (~ preset)  &  n_n4018  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1413 = ( (~ preset)  &  ndn3_3  &  n_n3250 ) | ( (~ preset)  &  n_n3250  &  nsr3_2 ) ;
 assign wire1418 = ( pdxport_1_1_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1419 = ( (~ preset)  &  ndn3_3  &  n_n4120 ) | ( (~ preset)  &  n_n4120  &  nsr3_2 ) ;
 assign wire1421 = ( (~ preset)  &  n_n4079  &  nld3_9 ) ;
 assign wire1422 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n4080 ) ;
 assign wire1423 = ( (~ preset)  &  ndn5_7  &  n_n4042 ) | ( (~ preset)  &  n_n4042  &  nsr5_7 ) ;
 assign wire1426 = ( (~ preset)  &  n_n3516  &  nld3_9 ) ;
 assign wire1427 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3517  &  ndn3_3 ) ;
 assign wire1430 = ( n_n3869  &  wire2071 ) | ( (~ preset)  &  n_n3869  &  n_n3833 ) ;
 assign wire1431 = ( n_n4036  &  wire2073 ) | ( n_n4036  &  wire2074 ) ;
 assign wire1432 = ( (~ preset)  &  ndn5_3  &  n_n3457 ) | ( (~ preset)  &  n_n3457  &  nsr5_3 ) ;
 assign wire1435 = ( (~ preset)  &  n_n3709  &  nld3_9 ) ;
 assign wire1436 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3356  &  ndn3_3 ) ;
 assign wire1437 = ( (~ preset)  &  n_n3387  &  ndn5_2 ) | ( (~ preset)  &  n_n3387  &  nsr5_2 ) ;
 assign wire1440 = ( (~ preset)  &  n_n3832  &  nld3_9 ) ;
 assign wire1441 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3262  &  ndn3_3 ) ;
 assign wire1443 = ( (~ preset)  &  n_n3509  &  ndn5_10 ) | ( (~ preset)  &  n_n3509  &  nsr5_7 ) ;
 assign wire1445 = ( (~ preset)  &  ndn5_4  &  n_n3921 ) | ( (~ preset)  &  n_n3921  &  nsr5_4 ) ;
 assign wire1446 = ( n_n3643  &  wire2071 ) | ( (~ preset)  &  n_n3643  &  n_n3833 ) ;
 assign wire1447 = ( n_n3340  &  wire2073 ) | ( n_n3340  &  wire2074 ) ;
 assign wire1448 = ( n_n3340  &  n_n3283  &  wire797 ) | ( n_n3340  &  wire797  &  wire839 ) | ( (~ n_n3340)  &  (~ n_n3283)  &  wire797  &  (~ wire839) ) ;
 assign wire1450 = ( (~ preset)  &  n_n3750  &  nld3_9 ) ;
 assign wire1451 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3751  &  ndn3_3 ) ;
 assign wire1453 = ( n_n4245  &  wire2071 ) | ( (~ preset)  &  n_n4245  &  n_n3833 ) ;
 assign wire1454 = ( n_n4246  &  wire2073 ) | ( n_n4246  &  wire2074 ) ;
 assign wire1456 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3065 ) | ( (~ preset)  &  n_n3065  &  nld3_9 ) ;
 assign wire1457 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3464 ) ;
 assign wire1460 = ( (~ preset)  &  (~ ndn5_9)  &  n_n4014 ) | ( (~ preset)  &  n_n4014  &  nld3_9 ) ;
 assign wire1461 = ( (~ preset)  &  n_n3709  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1464 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3855 ) | ( (~ preset)  &  n_n3855  &  nld3_9 ) ;
 assign wire1465 = ( (~ preset)  &  n_n3489  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1467 = ( (~ preset)  &  n_n3540  &  nld3_9 ) ;
 assign wire1468 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3541 ) ;
 assign wire1469 = ( (~ preset)  &  (~ ndn5_9)  &  n_n4259 ) | ( (~ preset)  &  n_n4259  &  nld3_9 ) ;
 assign wire1470 = ( (~ preset)  &  n_n3535  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1472 = ( (~ preset)  &  n_n3384  &  ndn3_3 ) | ( (~ preset)  &  n_n3384  &  nsr3_2 ) ;
 assign wire1475 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3182 ) | ( (~ preset)  &  n_n3182  &  nld3_9 ) ;
 assign wire1476 = ( (~ preset)  &  ndn5_9  &  n_n4079  &  (~ nld3_9) ) ;
 assign wire1477 = ( (~ preset)  &  (~ nen5_9)  &  n_n4158 ) | ( (~ preset)  &  ndn5_9  &  n_n4158 ) ;
 assign wire1495 = ( wire1500  &  wire7311 ) | ( n_n4194  &  nrq5_6  &  wire7311 ) ;
 assign wire1500 = ( nen5_9  &  n_n4193  &  (~ ndn5_9) ) ;
 assign wire1503 = ( (~ preset)  &  ndn5_5  &  n_n3776 ) | ( (~ preset)  &  n_n3776  &  nsr5_5 ) ;
 assign wire1505 = ( (~ preset)  &  n_n3947  &  ndn5_10 ) | ( (~ preset)  &  n_n3947  &  nsr5_7 ) ;
 assign wire1507 = ( (~ preset)  &  n_n4111  &  nld3_9 ) ;
 assign wire1508 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n4218 ) ;
 assign wire1509 = ( (~ preset)  &  n_n3625  &  ndn5_8 ) | ( (~ preset)  &  n_n3625  &  nsr5_8 ) ;
 assign wire1511 = ( (~ preset)  &  ndn5_7  &  n_n3679 ) | ( (~ preset)  &  n_n3679  &  nsr5_7 ) ;
 assign wire1514 = ( (~ preset)  &  n_n4232  &  ndn3_3 ) | ( (~ preset)  &  n_n4232  &  nsr3_2 ) ;
 assign wire1517 = ( (~ preset)  &  n_n4071  &  ndn5_2 ) | ( (~ preset)  &  n_n4071  &  nsr5_2 ) ;
 assign wire1520 = ( (~ preset)  &  n_n3684  &  ndn5_10 ) | ( (~ preset)  &  n_n3684  &  nsr5_7 ) ;
 assign wire1526 = ( (~ preset)  &  n_n3903  &  wire7302 ) ;
 assign wire1528 = ( (~ preset)  &  n_n3996  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1530 = ( (~ preset)  &  (~ nen5_9)  &  n_n3931 ) | ( (~ preset)  &  ndn5_9  &  n_n3931 ) ;
 assign wire1534 = ( (~ preset)  &  ndn5_4  &  n_n3659 ) | ( (~ preset)  &  n_n3659  &  nsr5_4 ) ;
 assign wire1535 = ( (~ preset)  &  n_n3480  &  ndn5_10 ) | ( (~ preset)  &  n_n3480  &  nsr5_7 ) ;
 assign wire1539 = ( wire802  &  (~ n_n3532)  &  wire2103 ) | ( wire802  &  (~ n_n3532)  &  wire2104 ) | ( wire802  &  n_n3532  &  (~ wire2103)  &  (~ wire2104) ) ;
 assign wire1540 = ( (~ preset)  &  (~ nen5_9)  &  n_n3774 ) | ( (~ preset)  &  ndn5_9  &  n_n3774 ) ;
 assign wire1544 = ( (~ preset)  &  n_n3715  &  nld3_9 ) ;
 assign wire1545 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3716 ) ;
 assign wire1546 = ( wire811  &  (~ n_n3363)  &  wire1638 ) | ( wire811  &  (~ n_n3363)  &  wire1639 ) | ( wire811  &  n_n3363  &  (~ wire1638)  &  (~ wire1639) ) ;
 assign wire1548 = ( (~ preset)  &  ndn5_3  &  n_n4030 ) | ( (~ preset)  &  n_n4030  &  nsr5_3 ) ;
 assign wire1553 = ( (~ preset)  &  (~ nen5_9)  &  n_n3212 ) | ( (~ preset)  &  ndn5_9  &  n_n3212 ) ;
 assign wire1559 = ( (~ preset)  &  n_n3356  &  ndn3_3 ) | ( (~ preset)  &  n_n3356  &  nsr3_2 ) ;
 assign wire1562 = ( (~ preset)  &  ndn5_3  &  n_n3711 ) | ( (~ preset)  &  n_n3711  &  nsr5_3 ) ;
 assign wire1564 = ( (~ preset)  &  ndn5_3  &  n_n3433 ) | ( (~ preset)  &  n_n3433  &  nsr5_3 ) ;
 assign wire1567 = ( (~ preset)  &  nld3_9  &  n_n3794 ) ;
 assign wire1568 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3417 ) ;
 assign wire1571 = ( paport_2_2_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1572 = ( (~ preset)  &  n_n3733  &  ndn3_3 ) | ( (~ preset)  &  n_n3733  &  nsr3_2 ) ;
 assign wire1574 = ( (~ preset)  &  n_n4230  &  ndn3_3 ) | ( (~ preset)  &  n_n4230  &  nsr3_2 ) ;
 assign wire1577 = ( wire802  &  (~ n_n3484)  &  wire1729 ) | ( wire802  &  (~ n_n3484)  &  wire1730 ) | ( wire802  &  n_n3484  &  (~ wire1729)  &  (~ wire1730) ) ;
 assign wire1578 = ( (~ preset)  &  (~ nen5_9)  &  n_n3540 ) | ( (~ preset)  &  ndn5_9  &  n_n3540 ) ;
 assign wire1582 = ( (~ preset)  &  n_n3062  &  ndn3_3 ) | ( (~ preset)  &  n_n3062  &  nsr3_2 ) ;
 assign wire1585 = ( paport_5_5_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1586 = ( (~ preset)  &  n_n4056  &  ndn3_3 ) | ( (~ preset)  &  n_n4056  &  nsr3_2 ) ;
 assign wire1588 = ( (~ preset)  &  (~ nen5_9)  &  n_n3214 ) | ( (~ preset)  &  ndn5_9  &  n_n3214 ) ;
 assign wire1589 = ( pdxport_5_5_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1590 = ( (~ preset)  &  n_n4179  &  ndn3_3 ) | ( (~ preset)  &  n_n4179  &  nsr3_2 ) ;
 assign wire1592 = ( (~ preset)  &  n_n4090  &  ndn3_3 ) | ( (~ preset)  &  n_n4090  &  nsr3_2 ) ;
 assign wire1596 = ( (~ preset)  &  nld3_9  &  n_n3442 ) ;
 assign wire1597 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n4106 ) ;
 assign wire1598 = ( n_n4151  &  wire2071 ) | ( (~ preset)  &  n_n4151  &  n_n3833 ) ;
 assign wire1599 = ( n_n4093  &  wire2073 ) | ( n_n4093  &  wire2074 ) ;
 assign wire1600 = ( n_n4093  &  wire797  &  wire940 ) | ( (~ n_n4093)  &  wire797  &  (~ wire940) ) ;
 assign wire1602 = ( (~ preset)  &  n_n3634  &  ndn3_3 ) | ( (~ preset)  &  n_n3634  &  nsr3_2 ) ;
 assign wire1605 = ( (~ preset)  &  (~ ndn5_9)  &  n_n3381 ) | ( (~ preset)  &  n_n3381  &  nld3_9 ) ;
 assign wire1606 = ( (~ preset)  &  ndn5_9  &  n_n3680  &  (~ nld3_9) ) ;
 assign wire1607 = ( paport_6_6_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1608 = ( (~ preset)  &  n_n4243  &  ndn3_3 ) | ( (~ preset)  &  n_n4243  &  nsr3_2 ) ;
 assign wire1610 = ( (~ preset)  &  n_n4159  &  ndn3_3 ) | ( (~ preset)  &  n_n4159  &  nsr3_2 ) ;
 assign wire1613 = ( pdxport_4_4_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1614 = ( (~ preset)  &  n_n4165  &  ndn3_3 ) | ( (~ preset)  &  n_n4165  &  nsr3_2 ) ;
 assign wire1617 = ( n_n4211  &  wire2071 ) | ( (~ preset)  &  n_n4211  &  n_n3833 ) ;
 assign wire1618 = ( n_n4212  &  wire2073 ) | ( n_n4212  &  wire2074 ) ;
 assign wire1619 = ( (~ preset)  &  ndn5_3  &  n_n3841 ) | ( (~ preset)  &  n_n3841  &  nsr5_3 ) ;
 assign wire1622 = ( (~ preset)  &  n_n3311  &  ndn5_5 ) | ( (~ preset)  &  n_n3311  &  nsr5_5 ) ;
 assign wire1623 = ( paport_7_7_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1624 = ( (~ preset)  &  n_n4054  &  ndn3_3 ) | ( (~ preset)  &  n_n4054  &  nsr3_2 ) ;
 assign wire1625 = ( wire802  &  (~ n_n3363)  &  wire1638 ) | ( wire802  &  (~ n_n3363)  &  wire1639 ) | ( wire802  &  n_n3363  &  (~ wire1638)  &  (~ wire1639) ) ;
 assign wire1626 = ( (~ preset)  &  (~ nen5_9)  &  n_n3713 ) | ( (~ preset)  &  ndn5_9  &  n_n3713 ) ;
 assign wire1631 = ( wire1636  &  wire7283 ) | ( n_n4070  &  nrq5_6  &  wire7283 ) ;
 assign wire1636 = ( nen5_9  &  (~ ndn5_9)  &  n_n3311 ) ;
 assign wire1638 = ( (~ n_n3950)  &  wire2051 ) | ( n_n3800  &  nrq5_6  &  (~ n_n3950) ) ;
 assign wire1639 = ( n_n3236  &  n_n3950  &  n_n3111 ) | ( n_n3950  &  (~ n_n3111)  &  wire849 ) ;
 assign wire1642 = ( pdxport_9_9_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1643 = ( (~ preset)  &  n_n4070  &  ndn3_3 ) | ( (~ preset)  &  n_n4070  &  nsr3_2 ) ;
 assign wire1645 = ( (~ preset)  &  (~ nen5_9)  &  n_n3179 ) | ( (~ preset)  &  ndn5_9  &  n_n3179 ) ;
 assign wire1646 = ( n_n3920  &  wire2071 ) | ( (~ preset)  &  n_n3920  &  n_n3833 ) ;
 assign wire1647 = ( n_n4004  &  wire2073 ) | ( n_n4004  &  wire2074 ) ;
 assign wire1649 = ( (~ preset)  &  pover_0_0_  &  ndn3_11 ) ;
 assign wire1650 = ( (~ preset)  &  pover_0_0_  &  (~ ngfdn_3) ) ;
 assign wire1652 = ( (~ preset)  &  n_n3293  &  ndn5_2 ) | ( (~ preset)  &  n_n3293  &  nsr5_2 ) ;
 assign wire1654 = ( (~ preset)  &  n_n3988  &  ndn5_2 ) | ( (~ preset)  &  n_n3988  &  nsr5_2 ) ;
 assign wire1656 = ( wire816  &  (~ n_n4129)  &  wire1937 ) | ( wire816  &  (~ n_n4129)  &  wire1938 ) | ( wire816  &  n_n4129  &  (~ wire1937)  &  (~ wire1938) ) ;
 assign wire1657 = ( (~ preset)  &  n_n3529  &  ndn5_10 ) | ( (~ preset)  &  n_n3529  &  nsr5_7 ) ;
 assign wire1660 = ( (~ preset)  &  (~ nen5_9)  &  n_n3677 ) | ( (~ preset)  &  ndn5_9  &  n_n3677 ) ;
 assign wire1666 = ( (~ preset)  &  pnext_0_0_  &  ndn5_16 ) ;
 assign wire1667 = ( (~ preset)  &  pnext_0_0_  &  (~ nld3_9) ) ;
 assign wire1669 = ( n_n3974  &  n_n3925  &  wire7263 ) | ( n_n3974  &  n_n4178  &  wire7263 ) | ( n_n3925  &  n_n4178  &  wire7263 ) ;
 assign wire1670 = ( (~ n_n4083)  &  wire813  &  (~ n_n4084)  &  n_n4082 ) | ( (~ n_n4083)  &  wire813  &  n_n4084  &  (~ n_n4082) ) ;
 assign wire1671 = ( n_n4083  &  wire797  &  (~ n_n4084)  &  (~ n_n4082) ) ;
 assign wire1672 = ( (~ preset)  &  n_n4083  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1674 = ( (~ preset)  &  nld3_9  &  n_n3475 ) ;
 assign wire1675 = ( (~ preset)  &  (~ ndn3_8)  &  n_n4230  &  ndn3_3 ) ;
 assign wire1677 = ( (~ preset)  &  nld3_9  &  n_n3981 ) ;
 assign wire1678 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3250 ) ;
 assign wire1686 = ( (~ preset)  &  n_n4193  &  ndn5_5 ) | ( (~ preset)  &  n_n4193  &  nsr5_5 ) ;
 assign wire1687 = ( (~ preset)  &  n_n3203  &  ndn5_7 ) | ( (~ preset)  &  n_n3203  &  nsr5_7 ) ;
 assign wire1690 = ( (~ preset)  &  n_n3741  &  ndn3_3 ) | ( (~ preset)  &  n_n3741  &  nsr3_2 ) ;
 assign wire1693 = ( wire802  &  (~ n_n4129)  &  wire1937 ) | ( wire802  &  (~ n_n4129)  &  wire1938 ) | ( wire802  &  n_n4129  &  (~ wire1937)  &  (~ wire1938) ) ;
 assign wire1694 = ( (~ preset)  &  (~ nen5_9)  &  n_n3875 ) | ( (~ preset)  &  n_n3875  &  ndn5_9 ) ;
 assign wire1697 = ( (~ preset)  &  ndn5_3  &  n_n3304 ) | ( (~ preset)  &  n_n3304  &  nsr5_3 ) ;
 assign wire1700 = ( (~ preset)  &  n_n3774  &  nld3_9 ) ;
 assign wire1701 = ( (~ preset)  &  (~ ndn3_8)  &  n_n4090  &  ndn3_3 ) ;
 assign wire1702 = ( (~ preset)  &  n_n3344  &  ndn5_2 ) | ( (~ preset)  &  n_n3344  &  nsr5_2 ) ;
 assign wire1705 = ( (~ preset)  &  (~ nen5_9)  &  n_n3821 ) | ( (~ preset)  &  n_n3821  &  ndn5_9 ) ;
 assign wire1708 = ( (~ preset)  &  (~ nen5_9)  &  n_n4114 ) | ( (~ preset)  &  n_n4114  &  ndn5_9 ) ;
 assign wire1721 = ( n_n4123  &  (~ wire7223)  &  (~ wire7224)  &  wire7228 ) ;
 assign wire1722 = ( n_n4123  &  (~ wire7223)  &  (~ wire7224)  &  wire7229 ) ;
 assign wire1723 = ( (~ n_n4123)  &  wire7230 ) | ( wire7223  &  wire7230 ) | ( wire7224  &  wire7230 ) ;
 assign wire1729 = ( (~ wire923)  &  (~ n_n4184) ) | ( (~ n_n4184)  &  wire1737 ) ;
 assign wire1730 = ( n_n4189  &  n_n4184  &  n_n3892 ) | ( n_n4184  &  wire883  &  (~ n_n3892) ) ;
 assign wire1733 = ( (~ n_n3359)  &  wire947  &  wire7251 ) | ( (~ wire946)  &  wire947  &  wire7251 ) | ( n_n3359  &  wire946  &  (~ wire947)  &  wire7251 ) ;
 assign wire1734 = ( (~ n_n3359)  &  wire947  &  wire7252 ) | ( (~ wire946)  &  wire947  &  wire7252 ) | ( n_n3359  &  wire946  &  (~ wire947)  &  wire7252 ) ;
 assign wire1735 = ( (~ n_n3359)  &  wire879  &  (~ wire947) ) | ( wire879  &  (~ wire946)  &  (~ wire947) ) | ( n_n3359  &  wire879  &  wire946  &  wire947 ) ;
 assign wire1736 = ( (~ n_n3359)  &  wire809  &  wire947 ) | ( wire809  &  (~ wire946)  &  wire947 ) | ( n_n3359  &  wire809  &  wire946  &  (~ wire947) ) ;
 assign wire1737 = ( nen5_9  &  (~ ndn5_9)  &  n_n3947 ) ;
 assign wire1745 = ( nen5_9  &  (~ ndn5_9)  &  n_n3788 ) ;
 assign wire1751 = ( (~ n_n3470)  &  (~ n_n3274) ) | ( ndn5_10  &  (~ n_n3274) ) | ( (~ n_n3274)  &  nsr5_7 ) ;
 assign wire1752 = ( (~ nen5_9)  &  (~ n_n3470) ) | ( ndn5_9  &  (~ n_n3470) ) ;
 assign wire1754 = ( nen5_9  &  (~ ndn5_9)  &  n_n3274 ) ;
 assign wire1769 = ( (~ preset)  &  n_n3796  &  ndn5_10 ) | ( (~ preset)  &  n_n3796  &  nsr5_7 ) ;
 assign wire1775 = ( (~ preset)  &  n_n3170  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3170  &  nld3_9 ) ;
 assign wire1776 = ( (~ preset)  &  ndn5_9  &  n_n3713  &  (~ nld3_9) ) ;
 assign wire1777 = ( (~ preset)  &  n_n3736  &  ndn5_7 ) | ( (~ preset)  &  n_n3736  &  nsr5_7 ) ;
 assign wire1780 = ( (~ preset)  &  n_n3931  &  nld3_9 ) ;
 assign wire1781 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3932 ) ;
 assign wire1783 = ( (~ preset)  &  n_n3875  &  nld3_9 ) ;
 assign wire1784 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3876 ) ;
 assign wire1785 = ( (~ preset)  &  ndn5_3  &  n_n3922 ) | ( (~ preset)  &  n_n3922  &  nsr5_3 ) ;
 assign wire1787 = ( (~ preset)  &  ndn5_3  &  n_n4117 ) | ( (~ preset)  &  n_n4117  &  nsr5_3 ) ;
 assign wire1790 = ( (~ preset)  &  n_n3248  &  ndn3_3 ) | ( (~ preset)  &  n_n3248  &  nsr3_2 ) ;
 assign wire1794 = ( (~ preset)  &  n_n3513  &  nld3_9 ) ;
 assign wire1795 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3062  &  ndn3_3 ) ;
 assign wire1797 = ( (~ preset)  &  n_n3815  &  ndn5_10 ) | ( (~ preset)  &  n_n3815  &  nsr5_7 ) ;
 assign wire1802 = ( (~ preset)  &  paport_1_1_  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1803 = ( (~ preset)  &  n_n3797  &  ndn3_3 ) | ( (~ preset)  &  n_n3797  &  nsr3_2 ) ;
 assign wire1804 = ( (~ preset)  &  n_n3460  &  (~ n_n3549)  &  wire955 ) ;
 assign wire1805 = ( (~ preset)  &  n_n3999  &  n_n3460  &  (~ wire2075) ) ;
 assign wire1806 = ( (~ preset)  &  n_n3128  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3128  &  nld3_9 ) ;
 assign wire1807 = ( (~ preset)  &  n_n3761  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1809 = ( (~ preset)  &  n_n3331  &  ndn3_3 ) | ( (~ preset)  &  n_n3331  &  nsr3_2 ) ;
 assign wire1814 = ( n_n3944  &  wire2071 ) | ( (~ preset)  &  n_n3944  &  n_n3833 ) ;
 assign wire1815 = ( n_n3369  &  wire2073 ) | ( n_n3369  &  wire2074 ) ;
 assign wire1816 = ( (~ preset)  &  n_n3221  &  ndn5_3 ) | ( (~ preset)  &  n_n3221  &  nsr5_3 ) ;
 assign wire1819 = ( (~ preset)  &  (~ nen5_9)  &  n_n3750 ) | ( (~ preset)  &  n_n3750  &  ndn5_9 ) ;
 assign wire1823 = ( (~ preset)  &  n_n3280  &  ndn3_3 ) | ( (~ preset)  &  n_n3280  &  nsr3_2 ) ;
 assign wire1826 = ( (~ n_n3460)  &  wire7207 ) | ( (~ wire955)  &  wire7207 ) | ( n_n3549  &  wire955  &  wire7207 ) ;
 assign wire1827 = ( (~ preset)  &  n_n3460  &  (~ n_n3549)  &  wire955 ) ;
 assign wire1828 = ( paport_10_10_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1829 = ( (~ preset)  &  n_n3882  &  ndn3_3 ) | ( (~ preset)  &  n_n3882  &  nsr3_2 ) ;
 assign wire1831 = ( (~ preset)  &  nld3_9  &  n_n3862 ) ;
 assign wire1832 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3280  &  ndn3_3 ) ;
 assign wire1835 = ( pdxport_8_8_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1836 = ( (~ preset)  &  n_n4242  &  ndn3_3 ) | ( (~ preset)  &  n_n4242  &  nsr3_2 ) ;
 assign wire1841 = ( (~ preset)  &  n_n3060  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3060  &  nld3_9 ) ;
 assign wire1842 = ( (~ preset)  &  ndn5_9  &  n_n3179  &  (~ nld3_9) ) ;
 assign wire1844 = ( (~ preset)  &  n_n3751  &  ndn3_3 ) | ( (~ preset)  &  n_n3751  &  nsr3_2 ) ;
 assign wire1848 = ( (~ preset)  &  n_n3235  &  ndn3_3 ) | ( (~ preset)  &  n_n3235  &  nsr3_2 ) ;
 assign wire1851 = ( (~ preset)  &  n_n3799  &  ndn5_7 ) | ( (~ preset)  &  n_n3799  &  nsr5_7 ) ;
 assign wire1855 = ( (~ preset)  &  n_n4133  &  ndn5_2 ) | ( (~ preset)  &  n_n4133  &  nsr5_2 ) ;
 assign wire1857 = ( (~ preset)  &  n_n4180  &  ndn5_2 ) | ( (~ preset)  &  n_n4180  &  nsr5_2 ) ;
 assign wire1859 = ( (~ preset)  &  n_n3019  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3019  &  nld3_9 ) ;
 assign wire1860 = ( (~ preset)  &  n_n3420  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire1865 = ( (~ preset)  &  n_n3928  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3928  &  nld3_9 ) ;
 assign wire1866 = ( (~ preset)  &  ndn5_9  &  n_n3677  &  (~ nld3_9) ) ;
 assign wire1867 = ( (~ preset)  &  n_n3585  &  ndn5_8 ) | ( (~ preset)  &  n_n3585  &  nsr5_8 ) ;
 assign wire1870 = ( (~ preset)  &  n_n3517  &  ndn3_3 ) | ( (~ preset)  &  n_n3517  &  nsr3_2 ) ;
 assign wire1873 = ( (~ preset)  &  n_n3164  &  ndn5_3 ) | ( (~ preset)  &  n_n3164  &  nsr5_3 ) ;
 assign wire1877 = ( (~ preset)  &  n_n3482  &  ndn5_7 ) | ( (~ preset)  &  n_n3482  &  nsr5_7 ) ;
 assign wire1879 = ( (~ preset)  &  n_n4039  &  ndn5_7 ) | ( (~ preset)  &  n_n4039  &  nsr5_7 ) ;
 assign wire1882 = ( (~ preset)  &  n_n3262  &  ndn3_3 ) | ( (~ preset)  &  n_n3262  &  nsr3_2 ) ;
 assign wire1886 = ( (~ preset)  &  n_n3822  &  ndn3_3 ) | ( (~ preset)  &  n_n3822  &  nsr3_2 ) ;
 assign wire1889 = ( paport_4_4_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1890 = ( (~ preset)  &  n_n3574  &  ndn3_3 ) | ( (~ preset)  &  n_n3574  &  nsr3_2 ) ;
 assign wire1894 = ( (~ preset)  &  (~ nen5_9)  &  n_n3709 ) | ( (~ preset)  &  n_n3709  &  ndn5_9 ) ;
 assign wire1898 = ( (~ preset)  &  n_n3011  &  ndn3_3 ) | ( (~ preset)  &  n_n3011  &  nsr3_2 ) ;
 assign wire1902 = ( (~ preset)  &  n_n3805  &  ndn5_4 ) | ( (~ preset)  &  n_n3805  &  nsr5_4 ) ;
 assign wire1904 = ( (~ preset)  &  n_n3870  &  ndn5_4 ) | ( (~ preset)  &  n_n3870  &  nsr5_4 ) ;
 assign wire1905 = ( (~ preset)  &  n_n4149  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n4149  &  nld3_9 ) ;
 assign wire1906 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3794 ) ;
 assign wire1908 = ( (~ preset)  &  (~ nen5_9)  &  n_n3516 ) | ( (~ preset)  &  n_n3516  &  ndn5_9 ) ;
 assign wire1915 = ( nen5_9  &  n_n3815  &  (~ ndn5_9) ) ;
 assign wire1929 = ( nen5_9  &  (~ ndn5_9)  &  n_n3529 ) ;
 assign wire1937 = ( (~ n_n3779)  &  (~ wire931) ) | ( (~ n_n3779)  &  wire2211 ) ;
 assign wire1938 = ( n_n3779  &  n_n4202  &  n_n3897 ) | ( n_n3779  &  n_n4202  &  n_n4062 ) | ( n_n3779  &  n_n3897  &  (~ n_n4062) ) ;
 assign wire1944 = ( (~ preset)  &  n_n3535  &  (~ nrq5_6) ) ;
 assign wire1948 = ( (~ preset)  &  n_n3071  &  ndn5_5 ) | ( (~ preset)  &  n_n3071  &  nsr5_5 ) ;
 assign wire1950 = ( (~ preset)  &  n_n3157  &  ndn5_5 ) | ( (~ preset)  &  n_n3157  &  nsr5_5 ) ;
 assign wire1955 = ( paport_3_3_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1956 = ( (~ preset)  &  n_n3778  &  ndn3_3 ) | ( (~ preset)  &  n_n3778  &  nsr3_2 ) ;
 assign wire1959 = ( (~ preset)  &  pdxport_3_3_  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire1960 = ( (~ preset)  &  n_n4220  &  ndn3_3 ) | ( (~ preset)  &  n_n4220  &  nsr3_2 ) ;
 assign wire1963 = ( (~ preset)  &  n_n3957  &  ndn5_8 ) | ( (~ preset)  &  n_n3957  &  nsr5_8 ) ;
 assign wire1966 = ( (~ preset)  &  nld3_9  &  n_n3464 ) ;
 assign wire1967 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3331  &  ndn3_3 ) ;
 assign wire1968 = ( n_n4083  &  n_n4084  &  wire7175 ) | ( n_n4083  &  n_n4082  &  wire7175 ) | ( n_n4084  &  n_n4082  &  wire7175 ) ;
 assign wire1969 = ( (~ n_n3949)  &  (~ n_n3948)  &  n_n4131  &  wire813 ) | ( (~ n_n3949)  &  n_n3948  &  (~ n_n4131)  &  wire813 ) ;
 assign wire1970 = ( n_n3949  &  wire797  &  (~ n_n3948)  &  (~ n_n4131) ) ;
 assign wire1971 = ( (~ preset)  &  n_n3949  &  (~ n_n3833)  &  (~ n_n3903) ) ;
 assign wire1974 = ( n_n4136  &  nrq5_2 ) | ( n_n4136  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1975 = ( n_n4132  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1976 = ( n_n4134  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1977 = ( n_n4135  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1978 = ( n_n4133  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1983 = ( n_n4183  &  nrq5_2 ) | ( n_n4183  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1984 = ( n_n4179  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1985 = ( n_n4181  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1986 = ( n_n4182  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1987 = ( n_n4180  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1990 = ( n_n3890  &  nrq5_2 ) | ( n_n3890  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire1991 = ( n_n4165  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire1992 = ( n_n3691  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire1993 = ( n_n3324  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire1994 = ( n_n3323  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire1999 = ( n_n4086  &  nrq5_2 ) | ( n_n4086  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2000 = ( n_n4057  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2001 = ( n_n3345  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2002 = ( n_n3346  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2003 = ( n_n3344  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2007 = ( n_n3971  &  nrq5_2 ) | ( n_n3971  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2008 = ( n_n3906  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2009 = ( n_n3745  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2010 = ( n_n3388  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2011 = ( n_n3387  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2012 = ( n_n3500  &  nrq5_2 ) | ( n_n3500  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2013 = ( n_n4120  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2014 = ( n_n2989  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2015 = ( n_n3708  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2016 = ( n_n3175  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2017 = ( n_n4224  &  nrq5_2 ) | ( n_n4224  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2018 = ( n_n4220  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2019 = ( n_n4222  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2020 = ( n_n4223  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2021 = ( n_n4221  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2022 = ( n_n3844  &  nrq5_2 ) | ( n_n3844  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2023 = ( n_n4206  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2024 = ( n_n3375  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2025 = ( n_n3312  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2026 = ( n_n3988  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2028 = ( (~ preset)  &  n_n3832  &  (~ nrq5_6) ) ;
 assign wire2031 = ( (~ preset)  &  n_n3715  &  (~ nen5_9) ) | ( (~ preset)  &  n_n3715  &  ndn5_9 ) ;
 assign wire2034 = ( (~ preset)  &  nld3_9  &  n_n3743 ) ;
 assign wire2035 = ( (~ preset)  &  (~ ndn3_8)  &  n_n3384  &  ndn3_3 ) ;
 assign wire2036 = ( (~ preset)  &  n_n3139  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n3139  &  nld3_9 ) ;
 assign wire2037 = ( (~ preset)  &  n_n3750  &  ndn5_9  &  (~ nld3_9) ) ;
 assign wire2038 = ( pdxport_10_10_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire2039 = ( (~ preset)  &  n_n4194  &  ndn3_3 ) | ( (~ preset)  &  n_n4194  &  nsr3_2 ) ;
 assign wire2041 = ( (~ preset)  &  n_n3791  &  (~ nen5_9) ) | ( (~ preset)  &  n_n3791  &  ndn5_9 ) ;
 assign wire2046 = ( wire2051  &  wire7136 ) | ( n_n3800  &  nrq5_6  &  wire7136 ) ;
 assign wire2051 = ( nen5_9  &  (~ ndn5_9)  &  n_n4252 ) ;
 assign wire2057 = ( pdxport_6_6_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire2058 = ( (~ preset)  &  n_n4206  &  ndn3_3 ) | ( (~ preset)  &  n_n4206  &  nsr3_2 ) ;
 assign wire2059 = ( pdxport_2_2_  &  (~ preset)  &  (~ ndn3_3)  &  (~ nsr3_2) ) ;
 assign wire2060 = ( (~ preset)  &  n_n4057  &  ndn3_3 ) | ( (~ preset)  &  n_n4057  &  nsr3_2 ) ;
 assign wire2061 = ( (~ preset)  &  n_n3700  &  ndn5_8 ) | ( (~ preset)  &  n_n3700  &  nsr5_8 ) ;
 assign wire2063 = ( (~ preset)  &  n_n2971  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n2971  &  nld3_9 ) ;
 assign wire2064 = ( (~ preset)  &  ndn5_9  &  (~ nld3_9)  &  n_n3862 ) ;
 assign wire2066 = ( (~ preset)  &  n_n4116  &  ndn5_4 ) | ( (~ preset)  &  n_n4116  &  nsr5_4 ) ;
 assign wire2068 = ( n_n4170  &  wire2071 ) | ( (~ preset)  &  n_n4170  &  n_n3833 ) ;
 assign wire2069 = ( n_n4171  &  wire2073 ) | ( n_n4171  &  wire2074 ) ;
 assign wire2071 = ( (~ n_n3578)  &  (~ n_n3460)  &  wire7128 ) | ( (~ n_n3578)  &  wire2075  &  wire7128 ) ;
 assign wire2073 = ( (~ n_n3578)  &  (~ n_n3460)  &  wire796 ) | ( (~ n_n3578)  &  wire796  &  wire2075 ) ;
 assign wire2074 = ( (~ preset)  &  (~ n_n3833)  &  (~ n_n3903)  &  (~ n_n3439) ) ;
 assign wire2075 = ( wire955  &  wire2247 ) | ( wire955  &  wire6973  &  wire6974 ) ;
 assign wire2080 = ( (~ preset)  &  n_n3489  &  (~ nrq5_6) ) ;
 assign wire2085 = ( wire2090  &  wire7113 ) | ( n_n4132  &  nrq5_6  &  wire7113 ) ;
 assign wire2090 = ( nen5_9  &  (~ ndn5_9)  &  n_n3069 ) ;
 assign wire2096 = ( wire2101  &  wire7021 ) | ( n_n3813  &  nrq5_6  &  wire7021 ) ;
 assign wire2101 = ( nen5_9  &  n_n4239  &  (~ ndn5_9) ) ;
 assign wire2103 = ( (~ n_n3635)  &  wire2112 ) | ( n_n3872  &  nrq5_6  &  (~ n_n3635) ) ;
 assign wire2104 = ( n_n3955  &  n_n3543  &  n_n3635 ) | ( (~ n_n3543)  &  wire851  &  n_n3635 ) ;
 assign wire2107 = ( wire2112  &  wire7035 ) | ( n_n3872  &  nrq5_6  &  wire7035 ) ;
 assign wire2112 = ( n_n3871  &  nen5_9  &  (~ ndn5_9) ) ;
 assign wire2118 = ( wire2123  &  wire7049 ) | ( n_n3868  &  nrq5_6  &  wire7049 ) ;
 assign wire2123 = ( n_n4099  &  nen5_9  &  (~ ndn5_9) ) ;
 assign wire2129 = ( wire2134  &  wire7063 ) | ( n_n3924  &  nrq5_6  &  wire7063 ) ;
 assign wire2134 = ( nen5_9  &  (~ ndn5_9)  &  n_n3923 ) ;
 assign wire2136 = ( (~ n_n3569)  &  wire2145 ) | ( n_n3919  &  nrq5_6  &  (~ n_n3569) ) ;
 assign wire2137 = ( n_n3569  &  n_n4153  &  n_n3035 ) | ( n_n3569  &  wire852  &  (~ n_n3035) ) ;
 assign wire2140 = ( wire2145  &  wire7077 ) | ( n_n3919  &  nrq5_6  &  wire7077 ) ;
 assign wire2145 = ( nen5_9  &  (~ ndn5_9)  &  n_n3918 ) ;
 assign wire2151 = ( wire2156  &  wire7091 ) | ( n_n4120  &  nrq5_6  &  wire7091 ) ;
 assign wire2156 = ( nen5_9  &  n_n3157  &  (~ ndn5_9) ) ;
 assign wire2160 = ( nen5_9  &  (~ ndn5_9)  &  n_n3910  &  n_n3939 ) ;
 assign wire2162 = ( (~ preset)  &  n_n3420  &  (~ nen5_9) ) | ( (~ preset)  &  n_n3420  &  ndn5_9 ) ;
 assign wire2172 = ( wire809  &  (~ n_n3434)  &  wire948 ) | ( wire809  &  n_n3434  &  (~ wire948) ) ;
 assign wire2181 = ( nen5_9  &  (~ ndn5_9)  &  n_n3829 ) ;
 assign wire2185 = ( n_n3521  &  (~ wire2202)  &  (~ wire2203)  &  (~ wire7008) ) ;
 assign wire2186 = ( (~ wire2189)  &  (~ wire2190)  &  wire7007 ) | ( (~ wire2189)  &  (~ wire2190)  &  wire7008 ) ;
 assign wire2189 = ( (~ n_n3976)  &  wire949  &  (~ wire7012)  &  (~ wire7013) ) | ( n_n3976  &  (~ wire949)  &  (~ wire7012)  &  (~ wire7013) ) ;
 assign wire2190 = ( (~ n_n4051)  &  wire2195 ) | ( (~ n_n4051)  &  wire7012 ) | ( (~ n_n4051)  &  wire7013 ) ;
 assign wire2195 = ( wire809  &  wire949  &  wire2235 ) | ( wire809  &  wire949  &  wire2236 ) | ( wire809  &  (~ wire949)  &  (~ wire2235)  &  (~ wire2236) ) ;
 assign wire2196 = ( nen5_9  &  n_n3796  &  (~ ndn5_9) ) ;
 assign wire2197 = ( n_n3971  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire2200 = ( n_n3976  &  wire950  &  wire7003 ) | ( (~ wire949)  &  wire950  &  wire7003 ) | ( (~ n_n3976)  &  wire949  &  (~ wire950)  &  wire7003 ) ;
 assign wire2201 = ( n_n3976  &  (~ wire950)  &  wire7004 ) | ( (~ wire949)  &  (~ wire950)  &  wire7004 ) | ( (~ n_n3976)  &  wire949  &  wire950  &  wire7004 ) ;
 assign wire2202 = ( n_n3976  &  wire950  &  wire7005 ) | ( (~ wire949)  &  wire950  &  wire7005 ) | ( (~ n_n3976)  &  wire949  &  (~ wire950)  &  wire7005 ) ;
 assign wire2203 = ( n_n3976  &  (~ wire950)  &  (~ wire935) ) | ( (~ wire949)  &  (~ wire950)  &  (~ wire935) ) | ( (~ n_n3976)  &  wire949  &  wire950  &  (~ wire935) ) ;
 assign wire2204 = ( wire809  &  n_n3976  &  wire950 ) | ( wire809  &  (~ wire949)  &  wire950 ) | ( wire809  &  (~ n_n3976)  &  wire949  &  (~ wire950) ) ;
 assign wire2207 = ( (~ n_n3434)  &  wire952  &  wire6989 ) | ( (~ wire948)  &  wire952  &  wire6989 ) | ( n_n3434  &  wire948  &  (~ wire952)  &  wire6989 ) ;
 assign wire2208 = ( (~ n_n3434)  &  wire952  &  wire6990 ) | ( (~ wire948)  &  wire952  &  wire6990 ) | ( n_n3434  &  wire948  &  (~ wire952)  &  wire6990 ) ;
 assign wire2209 = ( wire877  &  (~ n_n3434)  &  (~ wire952) ) | ( wire877  &  (~ wire948)  &  (~ wire952) ) | ( wire877  &  n_n3434  &  wire948  &  wire952 ) ;
 assign wire2210 = ( wire809  &  (~ n_n3434)  &  wire952 ) | ( wire809  &  (~ wire948)  &  wire952 ) | ( wire809  &  n_n3434  &  wire948  &  (~ wire952) ) ;
 assign wire2211 = ( nen5_9  &  (~ ndn5_9)  &  n_n3826 ) ;
 assign wire2235 = ( nen5_9  &  (~ ndn5_9)  &  n_n3625 ) ;
 assign wire2236 = ( n_n3626  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire2238 = ( (~ preset)  &  n_n3214  &  nld3_9 ) ;
 assign wire2239 = ( (~ preset)  &  (~ ndn3_8)  &  ndn3_3  &  n_n3786 ) ;
 assign wire2244 = ( (~ preset)  &  n_n3175  &  ndn5_2 ) | ( (~ preset)  &  n_n3175  &  nsr5_2 ) ;
 assign wire2247 = ( (~ n_n3838)  &  n_n3999 ) ;
 assign wire2248 = ( n_n4165  &  nrq5_2 ) | ( n_n4165  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2249 = ( n_n3424  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2250 = ( n_n4099  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2251 = ( n_n3868  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2252 = ( n_n3711  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2253 = ( n_n4132  &  nrq5_2 ) | ( n_n4132  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2254 = ( n_n3840  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2255 = ( n_n3842  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2256 = ( n_n3843  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2257 = ( n_n3841  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2258 = ( n_n4057  &  nrq5_2 ) | ( n_n4057  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2259 = ( n_n3367  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2260 = ( n_n3918  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2261 = ( n_n3919  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2262 = ( n_n3221  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2263 = ( n_n4220  &  nrq5_2 ) | ( n_n4220  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2264 = ( n_n3921  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2265 = ( n_n3923  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2266 = ( n_n3924  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2267 = ( n_n3922  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2268 = ( n_n3906  &  nrq5_2 ) | ( n_n3906  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2269 = ( n_n3303  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2270 = ( n_n3939  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2271 = ( n_n3940  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2272 = ( n_n3304  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2273 = ( n_n4120  &  nrq5_2 ) | ( n_n4120  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2274 = ( n_n4116  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2275 = ( n_n4118  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2276 = ( n_n4119  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2277 = ( n_n4117  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2278 = ( n_n4206  &  nrq5_2 ) | ( n_n4206  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2279 = ( n_n3188  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2280 = ( n_n4239  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2281 = ( n_n3813  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2282 = ( n_n3436  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2283 = ( n_n4194  &  nrq5_2 ) | ( n_n4194  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2284 = ( n_n4045  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2285 = ( n_n4176  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2286 = ( n_n4177  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2287 = ( n_n3457  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2288 = ( n_n4237  &  nrq5_2 ) | ( n_n4237  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2289 = ( n_n3659  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2290 = ( n_n4208  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2291 = ( n_n4209  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2292 = ( n_n3433  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2293 = ( n_n4179  &  nrq5_2 ) | ( n_n4179  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2294 = ( n_n3870  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2295 = ( n_n3871  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2296 = ( n_n3872  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2297 = ( n_n4030  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2298 = ( n_n4070  &  nrq5_2 ) | ( n_n4070  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2299 = ( n_n3805  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2300 = ( n_n3807  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2301 = ( n_n3808  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2302 = ( n_n3806  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2303 = ( n_n4242  &  nrq5_2 ) | ( n_n4242  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire2304 = ( n_n4047  &  (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire2305 = ( n_n4252  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire2306 = ( n_n3800  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire2307 = ( n_n3164  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire2308 = ( (~ preset)  &  n_n2960  &  (~ ndn5_9) ) | ( (~ preset)  &  n_n2960  &  nld3_9 ) ;
 assign wire2309 = ( (~ preset)  &  ndn5_9  &  n_n3540  &  (~ nld3_9) ) ;
 assign wire6930 = ( wire2249 ) | ( wire2250 ) | ( wire2251 ) | ( wire2252 ) ;
 assign wire6933 = ( wire2299 ) | ( wire2300 ) | ( wire2301 ) | ( wire2302 ) ;
 assign wire6936 = ( wire2264 ) | ( wire2265 ) | ( wire2266 ) | ( wire2267 ) ;
 assign wire6939 = ( wire2279 ) | ( wire2280 ) | ( wire2281 ) | ( wire2282 ) ;
 assign wire6942 = ( wire2254 ) | ( wire2255 ) | ( wire2256 ) | ( wire2257 ) ;
 assign wire6945 = ( wire2304 ) | ( wire2305 ) | ( wire2306 ) | ( wire2307 ) ;
 assign wire6948 = ( wire2289 ) | ( wire2290 ) | ( wire2291 ) | ( wire2292 ) ;
 assign wire6951 = ( wire2294 ) | ( wire2295 ) | ( wire2296 ) | ( wire2297 ) ;
 assign wire6954 = ( wire2274 ) | ( wire2275 ) | ( wire2276 ) | ( wire2277 ) ;
 assign wire6957 = ( wire2284 ) | ( wire2285 ) | ( wire2286 ) | ( wire2287 ) ;
 assign wire6960 = ( wire2259 ) | ( wire2260 ) | ( wire2261 ) | ( wire2262 ) ;
 assign wire6963 = ( wire2269 ) | ( wire2270 ) | ( wire2271 ) | ( wire2272 ) ;
 assign wire6964 = ( (~ n_n3999)  &  (~ wire2248)  &  (~ wire6930) ) ;
 assign wire6965 = ( (~ wire2263)  &  (~ wire2298)  &  (~ wire6933)  &  (~ wire6936) ) ;
 assign wire6966 = ( (~ wire2253)  &  (~ wire2278)  &  (~ wire6939)  &  (~ wire6942) ) ;
 assign wire6967 = ( (~ wire2288)  &  (~ wire2303)  &  (~ wire6945)  &  (~ wire6948) ) ;
 assign wire6968 = ( (~ wire2273)  &  (~ wire2293)  &  (~ wire6951)  &  (~ wire6954) ) ;
 assign wire6969 = ( (~ wire2258)  &  (~ wire2283)  &  (~ wire6957)  &  (~ wire6960) ) ;
 assign wire6973 = ( (~ wire2268)  &  (~ wire6963)  &  wire6964  &  wire6969 ) ;
 assign wire6974 = ( wire6965  &  wire6966  &  wire6967  &  wire6968 ) ;
 assign wire6975 = ( (~ nld3_9)  &  (~ preset) ) ;
 assign wire6976 = ( (~ pdn)  &  ndn3_8 ) | ( (~ pdn)  &  (~ ndn3_3) ) | ( ndn3_8  &  ndn1_4 ) | ( (~ ndn3_3)  &  ndn1_4 ) ;
 assign wire6977 = ( (~ preset)  &  pdn  &  (~ ndn1_4) ) ;
 assign wire6989 = ( (~ n_n3826)  &  ndn5_10 ) | ( (~ n_n3826)  &  (~ n_n4183) ) | ( (~ n_n3826)  &  nsr5_7 ) ;
 assign wire6990 = ( (~ nen5_9)  &  (~ n_n4183) ) | ( ndn5_9  &  (~ n_n4183) ) ;
 assign wire6993 = ( (~ n_n3890)  &  (~ n_n3509) ) | ( (~ n_n3509)  &  ndn5_10 ) | ( (~ n_n3509)  &  nsr5_7 ) ;
 assign wire6994 = ( nen5_9  &  (~ ndn5_9)  &  n_n3509 ) ;
 assign wire6995 = ( (~ nen5_9)  &  (~ n_n3890) ) | ( ndn5_9  &  (~ n_n3890) ) ;
 assign wire6996 = ( (~ n_n3434)  &  wire948  &  wire6993 ) | ( n_n3434  &  (~ wire948)  &  wire6993 ) | ( n_n3434  &  wire948  &  wire6994 ) | ( (~ n_n3434)  &  (~ wire948)  &  wire6994 ) ;
 assign wire6997 = ( n_n3434  &  wire948  &  (~ wire932) ) | ( (~ n_n3434)  &  (~ wire948)  &  (~ wire932) ) | ( (~ n_n3434)  &  wire948  &  wire6995 ) | ( n_n3434  &  (~ wire948)  &  wire6995 ) ;
 assign wire6999 = ( (~ n_n4224)  &  (~ n_n3829) ) | ( ndn5_10  &  (~ n_n3829) ) | ( (~ n_n3829)  &  nsr5_7 ) ;
 assign wire7000 = ( (~ nen5_9)  &  (~ n_n4224) ) | ( ndn5_9  &  (~ n_n4224) ) ;
 assign wire7002 = ( wire809  &  n_n4200 ) | ( (~ n_n4200)  &  (~ wire933) ) | ( (~ n_n4200)  &  wire2181 ) ;
 assign wire7003 = ( (~ n_n4086)  &  (~ n_n3480) ) | ( (~ n_n3480)  &  ndn5_10 ) | ( (~ n_n3480)  &  nsr5_7 ) ;
 assign wire7004 = ( nen5_9  &  (~ ndn5_9)  &  n_n3480 ) ;
 assign wire7005 = ( (~ nen5_9)  &  (~ n_n4086) ) | ( ndn5_9  &  (~ n_n4086) ) ;
 assign wire7007 = ( wire2203 ) | ( wire2202 ) ;
 assign wire7008 = ( wire2200 ) | ( wire2201 ) | ( wire2204 ) ;
 assign wire7009 = ( (~ n_n3500)  &  (~ n_n3684) ) | ( (~ n_n3684)  &  ndn5_10 ) | ( (~ n_n3684)  &  nsr5_7 ) ;
 assign wire7010 = ( nen5_9  &  (~ ndn5_9)  &  n_n3684 ) ;
 assign wire7011 = ( (~ n_n3500)  &  (~ nen5_9) ) | ( (~ n_n3500)  &  ndn5_9 ) ;
 assign wire7012 = ( n_n3976  &  wire949  &  wire7009 ) | ( (~ n_n3976)  &  (~ wire949)  &  wire7009 ) | ( (~ n_n3976)  &  wire949  &  wire7010 ) | ( n_n3976  &  (~ wire949)  &  wire7010 ) ;
 assign wire7013 = ( (~ n_n3976)  &  wire949  &  (~ wire936) ) | ( n_n3976  &  (~ wire949)  &  (~ wire936) ) | ( n_n3976  &  wire949  &  wire7011 ) | ( (~ n_n3976)  &  (~ wire949)  &  wire7011 ) ;
 assign wire7017 = ( (~ n_n4239)  &  (~ n_n3813) ) ;
 assign wire7018 = ( nen5_9  &  (~ ndn5_9)  &  n_n3630 ) ;
 assign wire7020 = ( n_n4206  &  (~ n_n3813)  &  (~ n_n4239) ) ;
 assign wire7021 = ( (~ n_n3630)  &  (~ n_n4206) ) ;
 assign wire7026 = ( wire7017  &  wire7018 ) | ( nrq5_6  &  wire7020 ) ;
 assign wire7027 = ( (~ n_n4239)  &  n_n3630  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n4239  &  (~ n_n3630)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7028 = ( (~ n_n4206)  &  n_n3813  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4206  &  (~ n_n3813)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7031 = ( n_n3071  &  (~ n_n3871) ) ;
 assign wire7032 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n3872) ) ;
 assign wire7034 = ( (~ n_n3871)  &  n_n4179  &  (~ n_n3872) ) ;
 assign wire7035 = ( (~ n_n4179)  &  (~ n_n3071) ) ;
 assign wire7040 = ( wire7031  &  wire7032 ) | ( nrq5_6  &  wire7034 ) ;
 assign wire7041 = ( (~ n_n3871)  &  n_n3071  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3871  &  (~ n_n3071)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7042 = ( (~ n_n4179)  &  n_n3872  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4179  &  (~ n_n3872)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7045 = ( n_n3776  &  (~ n_n4099) ) ;
 assign wire7046 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n3868) ) ;
 assign wire7048 = ( (~ n_n4099)  &  n_n4165  &  (~ n_n3868) ) ;
 assign wire7049 = ( (~ n_n3776)  &  (~ n_n4165) ) ;
 assign wire7054 = ( wire7045  &  wire7046 ) | ( nrq5_6  &  wire7048 ) ;
 assign wire7055 = ( (~ n_n4099)  &  n_n3776  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n4099  &  (~ n_n3776)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7056 = ( (~ n_n4165)  &  n_n3868  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4165  &  (~ n_n3868)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7059 = ( (~ n_n3923)  &  (~ n_n3924) ) ;
 assign wire7060 = ( nen5_9  &  (~ ndn5_9)  &  n_n3143 ) ;
 assign wire7062 = ( n_n4220  &  (~ n_n3924)  &  (~ n_n3923) ) ;
 assign wire7063 = ( (~ n_n3143)  &  (~ n_n4220) ) ;
 assign wire7068 = ( wire7059  &  wire7060 ) | ( nrq5_6  &  wire7062 ) ;
 assign wire7069 = ( (~ n_n3923)  &  n_n3143  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3923  &  (~ n_n3143)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7070 = ( (~ n_n4220)  &  n_n3924  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4220  &  (~ n_n3924)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7073 = ( (~ n_n3918)  &  (~ n_n3919) ) ;
 assign wire7074 = ( nen5_9  &  (~ ndn5_9)  &  n_n3793 ) ;
 assign wire7076 = ( n_n4057  &  (~ n_n3919)  &  (~ n_n3918) ) ;
 assign wire7077 = ( (~ n_n3793)  &  (~ n_n4057) ) ;
 assign wire7082 = ( wire7073  &  wire7074 ) | ( nrq5_6  &  wire7076 ) ;
 assign wire7083 = ( (~ n_n3918)  &  n_n3793  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3918  &  (~ n_n3793)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7084 = ( (~ n_n4057)  &  n_n3919  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4057  &  (~ n_n3919)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7087 = ( (~ n_n4120)  &  (~ n_n3157) ) ;
 assign wire7088 = ( nen5_9  &  (~ ndn5_9)  &  n_n4118 ) ;
 assign wire7090 = ( (~ n_n3157)  &  (~ n_n4120)  &  n_n4119 ) ;
 assign wire7091 = ( (~ n_n4118)  &  (~ n_n4119) ) ;
 assign wire7096 = ( wire7087  &  wire7088 ) | ( nrq5_6  &  wire7090 ) ;
 assign wire7097 = ( (~ n_n3157)  &  n_n4118  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3157  &  (~ n_n4118)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7098 = ( (~ n_n4120)  &  n_n4119  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4120  &  (~ n_n4119)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7102 = ( nen5_9  &  (~ ndn5_9)  &  n_n3906  &  n_n3939 ) ;
 assign wire7104 = ( nen5_9  &  (~ ndn5_9)  &  n_n3940  &  n_n3910 ) ;
 assign wire7107 = ( wire2160 ) | ( nrq5_6  &  wire7102 ) ;
 assign wire7108 = ( nrq5_6  &  wire7104 ) | ( n_n3940  &  n_n3906  &  nrq5_6 ) ;
 assign wire7109 = ( n_n3842  &  (~ n_n3069) ) ;
 assign wire7110 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n4132) ) ;
 assign wire7112 = ( n_n3843  &  (~ n_n3069)  &  (~ n_n4132) ) ;
 assign wire7113 = ( (~ n_n3842)  &  (~ n_n3843) ) ;
 assign wire7118 = ( wire7109  &  wire7110 ) | ( nrq5_6  &  wire7112 ) ;
 assign wire7119 = ( (~ n_n3069)  &  n_n3842  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3069  &  (~ n_n3842)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7120 = ( (~ n_n3843)  &  n_n4132  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n3843  &  (~ n_n4132)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7125 = ( nsr5_4  &  (~ nsr5_3) ) | ( nsr5_3  &  (~ nsr5_2) ) ;
 assign wire7126 = ( (~ nsr5_5)  &  nsr5_7 ) | ( (~ nsr5_7)  &  nsr5_8 ) ;
 assign wire7128 = ( (~ preset)  &  wire2247 ) | ( (~ preset)  &  wire6973  &  wire6974 ) ;
 assign wire7129 = ( (~ n_n4214)  &  (~ wire2247)  &  (~ wire6973) ) | ( (~ n_n4214)  &  (~ wire2247)  &  (~ wire6974) ) ;
 assign wire7130 = ( n_n4171  &  wire797  &  wire918 ) | ( (~ n_n4171)  &  wire797  &  (~ wire918) ) ;
 assign wire7132 = ( n_n3607  &  (~ n_n3800) ) ;
 assign wire7133 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n4252) ) ;
 assign wire7135 = ( n_n4242  &  (~ n_n3800)  &  (~ n_n4252) ) ;
 assign wire7136 = ( (~ n_n3607)  &  (~ n_n4242) ) ;
 assign wire7141 = ( wire7132  &  wire7133 ) | ( nrq5_6  &  wire7135 ) ;
 assign wire7142 = ( (~ n_n3607)  &  n_n4252  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3607  &  (~ n_n4252)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7143 = ( (~ n_n4242)  &  n_n3800  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4242  &  (~ n_n3800)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7149 = ( wire2023 ) | ( wire2024 ) | ( wire2025 ) | ( wire2026 ) ;
 assign wire7152 = ( wire2018 ) | ( wire2019 ) | ( wire2020 ) | ( wire2021 ) ;
 assign wire7155 = ( wire2008 ) | ( wire2009 ) | ( wire2010 ) | ( wire2011 ) ;
 assign wire7158 = ( wire2013 ) | ( wire2014 ) | ( wire2015 ) | ( wire2016 ) ;
 assign wire7164 = ( wire2000 ) | ( wire2001 ) | ( wire2002 ) | ( wire2003 ) ;
 assign wire7167 = ( wire1991 ) | ( wire1992 ) | ( wire1993 ) | ( wire1994 ) ;
 assign wire7170 = ( wire1984 ) | ( wire1985 ) | ( wire1986 ) | ( wire1987 ) ;
 assign wire7173 = ( wire1975 ) | ( wire1976 ) | ( wire1977 ) | ( wire1978 ) ;
 assign wire7175 = ( n_n3949  &  wire797  &  wire1974 ) | ( n_n3949  &  wire797  &  wire7173 ) ;
 assign wire7183 = ( (~ n_n3844)  &  (~ n_n3529) ) | ( (~ n_n3529)  &  ndn5_10 ) | ( (~ n_n3529)  &  nsr5_7 ) ;
 assign wire7184 = ( (~ nen5_9)  &  (~ n_n3844) ) | ( (~ n_n3844)  &  ndn5_9 ) ;
 assign wire7186 = ( n_n3404  &  wire809 ) | ( (~ n_n3404)  &  (~ wire926) ) | ( (~ n_n3404)  &  wire1929 ) ;
 assign wire7189 = ( (~ n_n3815)  &  (~ n_n4136) ) | ( (~ n_n3815)  &  ndn5_10 ) | ( (~ n_n3815)  &  nsr5_7 ) ;
 assign wire7190 = ( (~ nen5_9)  &  (~ n_n4136) ) | ( ndn5_9  &  (~ n_n4136) ) ;
 assign wire7191 = ( (~ n_n3359)  &  wire946  &  wire7189 ) | ( n_n3359  &  (~ wire946)  &  wire7189 ) | ( (~ n_n3359)  &  wire946  &  wire7190 ) | ( n_n3359  &  (~ wire946)  &  wire7190 ) ;
 assign wire7192 = ( (~ n_n3359)  &  wire809  &  wire946 ) | ( n_n3359  &  wire809  &  (~ wire946) ) | ( n_n3359  &  wire946  &  wire883 ) | ( (~ n_n3359)  &  (~ wire946)  &  wire883 ) ;
 assign wire7196 = ( (~ n_n4126)  &  (~ n_n3283) ) ;
 assign wire7197 = ( (~ n_n4171)  &  (~ n_n3369)  &  (~ n_n4060) ) ;
 assign wire7198 = ( (~ n_n4212)  &  (~ n_n4246)  &  (~ n_n4036)  &  (~ n_n3961) ) ;
 assign wire7201 = ( n_n3903  &  wire7196  &  wire7197  &  wire7198 ) ;
 assign wire7203 = ( n_n4171  &  (~ n_n3099)  &  wire7201 ) | ( wire918  &  (~ n_n3099)  &  wire7201 ) ;
 assign wire7205 = ( (~ n_n4093)  &  wire940  &  wire7203 ) | ( n_n4093  &  (~ wire940)  &  wire7203 ) ;
 assign wire7207 = ( n_n3838  &  (~ preset) ) ;
 assign wire7209 = ( n_n3369  &  wire797  &  n_n3301 ) | ( (~ n_n3369)  &  wire797  &  (~ n_n3301) ) ;
 assign wire7219 = ( (~ n_n3482)  &  (~ n_n4075) ) | ( (~ n_n4075)  &  ndn5_10 ) | ( (~ n_n4075)  &  nsr5_7 ) ;
 assign wire7220 = ( (~ nen5_9)  &  (~ n_n3482) ) | ( (~ n_n3482)  &  ndn5_9 ) ;
 assign wire7221 = ( nen5_9  &  (~ ndn5_9)  &  n_n4075 ) ;
 assign wire7223 = ( n_n4123  &  (~ wire914) ) | ( n_n4123  &  wire7221 ) ;
 assign wire7224 = ( wire809  &  (~ n_n4123) ) | ( (~ n_n4123)  &  wire7219 ) | ( (~ n_n4123)  &  wire7220 ) ;
 assign wire7225 = ( n_n4075  &  (~ n_n3612) ) ;
 assign wire7226 = ( nen5_9  &  (~ ndn5_9)  &  ndn5_10 ) | ( nen5_9  &  (~ ndn5_9)  &  nsr5_7 ) ;
 assign wire7227 = ( (~ nen5_9)  &  (~ n_n4039) ) | ( (~ n_n4039)  &  ndn5_9 ) ;
 assign wire7228 = ( nen5_9  &  (~ ndn5_9)  &  n_n3612 ) ;
 assign wire7229 = ( n_n4039  &  (~ ndn5_10)  &  (~ nsr5_7) ) ;
 assign wire7230 = ( (~ n_n3612)  &  (~ n_n4039) ) ;
 assign wire7231 = ( (~ nen5_9)  &  (~ n_n4039) ) | ( (~ n_n4039)  &  ndn5_9 ) ;
 assign wire7232 = ( (~ n_n3612)  &  ndn5_10 ) | ( (~ n_n3612)  &  nsr5_7 ) ;
 assign wire7233 = ( wire7225  &  wire7226 ) | ( (~ wire914)  &  wire7227 ) ;
 assign wire7234 = ( wire7233 ) | ( (~ n_n4123)  &  wire7231 ) ;
 assign wire7236 = ( wire7234 ) | ( wire809  &  (~ n_n4123) ) | ( (~ n_n4123)  &  wire7232 ) ;
 assign wire7239 = ( (~ n_n4095)  &  (~ n_n4167) ) | ( (~ n_n4167)  &  ndn5_10 ) | ( (~ n_n4167)  &  nsr5_7 ) ;
 assign wire7240 = ( (~ nen5_9)  &  (~ n_n4095) ) | ( ndn5_9  &  (~ n_n4095) ) ;
 assign wire7241 = ( nen5_9  &  (~ ndn5_9)  &  n_n4167 ) ;
 assign wire7243 = ( (~ n_n4160)  &  (~ wire934) ) | ( (~ n_n4160)  &  wire7241 ) ;
 assign wire7244 = ( wire809  &  n_n4160 ) | ( n_n4160  &  wire7239 ) | ( n_n4160  &  wire7240 ) ;
 assign wire7245 = ( (~ wire880)  &  wire916  &  (~ wire7223)  &  (~ wire7224) ) ;
 assign wire7246 = ( wire880  &  (~ wire916)  &  wire7223 ) | ( wire880  &  (~ wire916)  &  wire7224 ) ;
 assign wire7247 = ( (~ n_n4140)  &  (~ n_n3788) ) | ( (~ n_n3788)  &  ndn5_10 ) | ( (~ n_n3788)  &  nsr5_7 ) ;
 assign wire7248 = ( (~ nen5_9)  &  (~ n_n4140) ) | ( ndn5_9  &  (~ n_n4140) ) ;
 assign wire7250 = ( wire809  &  n_n4248 ) | ( (~ n_n4248)  &  (~ wire930) ) | ( (~ n_n4248)  &  wire1745 ) ;
 assign wire7251 = ( (~ n_n3810)  &  (~ n_n3947) ) | ( (~ n_n3947)  &  ndn5_10 ) | ( (~ n_n3947)  &  nsr5_7 ) ;
 assign wire7252 = ( (~ nen5_9)  &  (~ n_n3810) ) | ( (~ n_n3810)  &  ndn5_9 ) ;
 assign wire7257 = ( wire7243  &  wire7245 ) | ( wire7244  &  wire7245 ) | ( (~ wire7243)  &  (~ wire7244)  &  wire7246 ) ;
 assign wire7263 = ( n_n4083  &  wire797  &  wire2022 ) | ( n_n4083  &  wire797  &  wire7149 ) ;
 assign wire7270 = ( nen5_9  &  (~ ndn5_9)  &  n_n3939 ) ;
 assign wire7271 = ( nen5_9  &  (~ ndn5_9)  &  n_n3910 ) ;
 assign wire7272 = ( nrq5_6  &  n_n3906 ) ;
 assign wire7273 = ( nrq5_6  &  n_n3940 ) ;
 assign wire7274 = ( (~ wire7107)  &  (~ wire7108)  &  wire7270 ) | ( (~ wire7107)  &  (~ wire7108)  &  wire7271 ) ;
 assign wire7275 = ( (~ wire7107)  &  (~ wire7108)  &  wire7272 ) | ( (~ wire7107)  &  (~ wire7108)  &  wire7273 ) ;
 assign wire7279 = ( (~ n_n3311)  &  (~ n_n4070) ) ;
 assign wire7280 = ( nen5_9  &  (~ ndn5_9)  &  n_n3807 ) ;
 assign wire7282 = ( n_n3808  &  (~ n_n4070)  &  (~ n_n3311) ) ;
 assign wire7283 = ( (~ n_n3807)  &  (~ n_n3808) ) ;
 assign wire7288 = ( wire7279  &  wire7280 ) | ( nrq5_6  &  wire7282 ) ;
 assign wire7289 = ( (~ n_n3311)  &  n_n3807  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n3311  &  (~ n_n3807)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7290 = ( (~ n_n3808)  &  n_n4070  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n3808  &  (~ n_n4070)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7294 = ( n_n4212  &  wire797  &  wire838 ) | ( (~ n_n4212)  &  wire797  &  (~ wire838) ) ;
 assign wire7302 = ( (~ n_n3996)  &  (~ n_n3888)  &  wire2017 ) | ( (~ n_n3996)  &  (~ n_n3888)  &  wire7152 ) | ( (~ n_n3996)  &  n_n3888  &  (~ wire2017)  &  (~ wire7152) ) ;
 assign wire7304 = ( n_n3996  &  wire797  &  n_n4219  &  n_n3888 ) | ( n_n3996  &  wire797  &  (~ n_n4219)  &  (~ n_n3888) ) ;
 assign wire7307 = ( (~ n_n4193)  &  (~ n_n4194) ) ;
 assign wire7308 = ( nen5_9  &  (~ ndn5_9)  &  n_n4176 ) ;
 assign wire7310 = ( (~ n_n4194)  &  (~ n_n4193)  &  n_n4177 ) ;
 assign wire7311 = ( (~ n_n4177)  &  (~ n_n4176) ) ;
 assign wire7316 = ( wire7307  &  wire7308 ) | ( nrq5_6  &  wire7310 ) ;
 assign wire7317 = ( (~ n_n4193)  &  n_n4176  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n4193  &  (~ n_n4176)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7318 = ( (~ n_n4194)  &  n_n4177  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4194  &  (~ n_n4177)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7322 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n4209) ) ;
 assign wire7324 = ( nen5_9  &  (~ ndn5_9)  &  (~ n_n4237) ) ;
 assign wire7326 = ( (~ n_n4208)  &  n_n4237  &  (~ n_n4209) ) ;
 assign wire7328 = ( (~ n_n4236)  &  (~ n_n4237)  &  n_n4209 ) ;
 assign wire7333 = ( n_n4236  &  (~ n_n4208)  &  wire7322 ) | ( (~ n_n4236)  &  n_n4208  &  wire7324 ) ;
 assign wire7334 = ( nrq5_6  &  wire7326 ) | ( nrq5_6  &  wire7328 ) ;
 assign wire7335 = ( (~ n_n4236)  &  n_n4208  &  nrq5_9  &  (~ nrq5_6) ) | ( n_n4236  &  (~ n_n4208)  &  nrq5_9  &  (~ nrq5_6) ) ;
 assign wire7336 = ( (~ n_n4237)  &  n_n4209  &  (~ nrq5_9)  &  nrq5_6 ) | ( n_n4237  &  (~ n_n4209)  &  (~ nrq5_9)  &  nrq5_6 ) ;
 assign wire7347 = ( n_n4093  &  n_n4246  &  wire797 ) | ( (~ n_n4093)  &  n_n4246  &  wire797  &  wire940 ) | ( (~ n_n4093)  &  (~ n_n4246)  &  wire797  &  (~ wire940) ) ;
 assign wire7354 = ( n_n4171  &  n_n4036  &  wire797 ) | ( n_n4036  &  wire797  &  wire918 ) | ( (~ n_n4171)  &  (~ n_n4036)  &  wire797  &  (~ wire918) ) ;
 assign wire7360 = ( n_n4018  &  wire797  &  wire1990 ) | ( n_n4018  &  wire797  &  wire7167 ) ;
 assign wire7361 = ( (~ preset)  &  wire907  &  n_n3903 ) ;
 assign wire7364 = ( (~ n_n3925)  &  wire7361 ) | ( n_n4018  &  wire797  &  (~ n_n3925) ) ;
 assign wire7365 = ( (~ n_n3965)  &  wire2007 ) | ( (~ n_n3965)  &  wire7155 ) ;
 assign wire7368 = ( n_n4027  &  n_n3965 ) ;
 assign wire7370 = ( wire797  &  wire2007  &  wire7368 ) | ( wire797  &  wire7155  &  wire7368 ) ;
 assign wire7372 = ( n_n3965  &  wire797  &  (~ n_n3991) ) ;
 assign wire7373 = ( (~ n_n3965)  &  (~ n_n4027)  &  n_n3837 ) | ( (~ n_n4027)  &  (~ n_n3966)  &  n_n3837 ) ;
 assign wire7375 = ( wire1386 ) | ( n_n4027  &  wire797  &  (~ n_n3991) ) ;
 assign wire7381 = ( wire1362 ) | ( wire1363 ) | ( wire1364 ) | ( wire1365 ) ;
 assign wire7384 = ( wire1367 ) | ( wire1368 ) | ( wire1369 ) | ( wire1370 ) ;
 assign wire7387 = ( wire1353 ) | ( wire1354 ) | ( wire1355 ) | ( wire1356 ) ;
 assign wire7389 = ( n_n4197  &  wire797  &  wire1352 ) | ( n_n4197  &  wire797  &  wire7387 ) ;
 assign wire7405 = ( (~ n_n3733)  &  n_n3794 ) | ( (~ n_n3797)  &  (~ n_n3916)  &  n_n3794 ) ;
 assign wire7407 = ( n_n3535  &  (~ n_n3797)  &  n_n3794 ) | ( n_n3535  &  n_n4111  &  n_n3794 ) ;
 assign wire7408 = ( n_n3535  &  (~ n_n3733)  &  (~ n_n3916) ) | ( (~ n_n3797)  &  (~ n_n3733)  &  (~ n_n3916) ) ;
 assign wire7409 = ( n_n3535  &  (~ n_n3733)  &  n_n4111 ) | ( (~ n_n3797)  &  (~ n_n3733)  &  n_n4111 ) ;
 assign wire7410 = ( wire7405 ) | ( n_n3535  &  (~ n_n3797)  &  (~ n_n3733) ) ;
 assign wire7411 = ( wire1327 ) | ( wire1328 ) | ( wire7407 ) ;
 assign wire7412 = ( wire7409 ) | ( wire7408 ) ;
 assign wire7414 = ( n_n3778  &  n_n3574  &  (~ n_n3981) ) ;
 assign wire7415 = ( (~ n_n3832)  &  n_n3778  &  (~ n_n3981) ) ;
 assign wire7416 = ( (~ n_n3981)  &  n_n3574 ) ;
 assign wire7417 = ( (~ n_n3981)  &  (~ n_n3832) ) ;
 assign wire7418 = ( n_n3574  &  n_n3778 ) ;
 assign wire7419 = ( n_n3778  &  (~ n_n3832) ) ;
 assign wire7423 = ( wire1319 ) | ( wire1324 ) | ( (~ n_n3832)  &  n_n3574 ) ;
 assign wire7424 = ( wire1320 ) | ( wire1321 ) | ( wire1322 ) | ( wire1323 ) ;
 assign wire7425 = ( (~ n_n3761)  &  n_n4243 ) | ( n_n4243  &  n_n4056 ) | ( (~ n_n3761)  &  (~ n_n3862) ) | ( n_n4056  &  (~ n_n3862) ) ;
 assign wire7426 = ( n_n3761  &  (~ n_n4056)  &  n_n3862 ) ;
 assign wire7427 = ( n_n3761  &  (~ n_n4243)  &  (~ n_n4056) ) ;
 assign wire7428 = ( n_n3832  &  (~ n_n3778) ) | ( (~ n_n3778)  &  (~ n_n3574) ) | ( n_n3832  &  n_n3981 ) | ( (~ n_n3574)  &  n_n3981 ) ;
 assign wire7429 = ( n_n3862  &  (~ n_n4056) ) ;
 assign wire7430 = ( n_n3862  &  n_n3761 ) ;
 assign wire7431 = ( (~ n_n4056)  &  (~ n_n4243) ) ;
 assign wire7432 = ( (~ n_n4243)  &  n_n3761 ) ;
 assign wire7433 = ( wire7423  &  wire7426 ) | ( wire7424  &  wire7426 ) | ( wire7423  &  wire7427 ) | ( wire7424  &  wire7427 ) ;
 assign wire7436 = ( wire1316 ) | ( wire7433 ) ;
 assign wire7437 = ( wire1312 ) | ( wire1313 ) | ( wire1314 ) | ( wire1315 ) ;
 assign wire7438 = ( n_n3489  &  wire7436 ) | ( (~ n_n4054)  &  wire7436 ) | ( n_n3489  &  wire7437 ) | ( (~ n_n4054)  &  wire7437 ) ;
 assign wire7439 = ( (~ n_n3489)  &  n_n4015 ) | ( n_n4054  &  n_n4015 ) ;
 assign wire7440 = ( (~ n_n3489)  &  (~ n_n3908) ) | ( (~ n_n3908)  &  n_n4054 ) ;
 assign wire7441 = ( n_n4015  &  wire1316 ) | ( n_n4015  &  wire7433 ) | ( n_n4015  &  wire7437 ) ;
 assign wire7442 = ( (~ n_n3908)  &  wire1316 ) | ( (~ n_n3908)  &  wire7433 ) | ( (~ n_n3908)  &  wire7437 ) ;
 assign wire7443 = ( n_n3396  &  wire7439 ) | ( n_n3396  &  wire7440 ) ;
 assign wire7447 = ( (~ n_n3513)  &  n_n3581 ) | ( n_n3818  &  n_n3581 ) ;
 assign wire7449 = ( nld3_9  &  (~ n_n4205)  &  n_n3336 ) ;
 assign wire7451 = ( nld3_9  &  (~ n_n4205)  &  n_n3336 ) ;
 assign wire7454 = ( n_n3336  &  nld3_9 ) ;
 assign wire7455 = ( (~ n_n4205)  &  nld3_9 ) ;
 assign wire7456 = ( wire1286 ) | ( wire818  &  wire7449 ) ;
 assign wire7462 = ( n_n4145  &  wire797  &  wire1361 ) | ( n_n4145  &  wire797  &  wire7381 ) ;
 assign wire7467 = ( (~ nlak3_2)  &  pready_0_0_ ) ;
 assign wire7468 = ( (~ preset)  &  (~ pdn)  &  nsr3_2 ) ;
 assign wire7472 = ( n_n3912  &  wire797  &  wire1366 ) | ( n_n3912  &  wire797  &  wire7384 ) ;
 assign wire7478 = ( (~ n_n3961)  &  n_n4060  &  wire797 ) | ( n_n3961  &  (~ n_n4060)  &  wire797 ) ;
 assign wire7483 = ( n_n3283  &  wire797  &  wire839 ) | ( (~ n_n3283)  &  wire797  &  (~ wire839) ) ;
 assign wire7486 = ( n_n3974  &  wire797  &  wire1983 ) | ( n_n3974  &  wire797  &  wire7170 ) ;
 assign wire7495 = ( n_n3961  &  n_n4126  &  wire797 ) | ( n_n4126  &  (~ n_n4060)  &  wire797 ) | ( (~ n_n3961)  &  (~ n_n4126)  &  n_n4060  &  wire797 ) ;
 assign wire7500 = ( wire1041 ) | ( wire1042 ) | ( wire1043 ) | ( wire1044 ) ;
 assign wire7501 = ( (~ preset)  &  (~ n_n4227)  &  n_n3903 ) ;
 assign wire7502 = ( wire797  &  n_n4227 ) ;
 assign wire7506 = ( (~ n_n3992)  &  (~ n_n3991)  &  wire1999 ) | ( (~ n_n3992)  &  (~ n_n3991)  &  wire7164 ) | ( (~ n_n3992)  &  n_n3991  &  (~ wire1999)  &  (~ wire7164) ) ;
 assign wire7508 = ( n_n3992  &  wire797  &  n_n3991  &  n_n3993 ) | ( n_n3992  &  wire797  &  (~ n_n3991)  &  (~ n_n3993) ) ;
 assign wire7511 = ( (~ preset)  &  n_n4214  &  n_n3462 ) ;
 assign wire7512 = ( preset ) | ( (~ n_n3460) ) | ( (~ wire955) ) | ( n_n3549  &  wire955 ) ;
 assign wire7518 = ( (~ n_n4060)  &  (~ wire2268)  &  (~ wire6963) ) ;
 assign wire7520 = ( (~ n_n4060)  &  (~ wire2268)  &  (~ wire6963) ) ;
 assign wire7521 = ( wire2247  &  wire7520 ) | ( wire6973  &  wire6974  &  wire7520 ) ;
 assign wire7524 = ( n_n3575  &  n_n4060 ) | ( (~ n_n4214)  &  n_n4060 ) | ( n_n4060  &  (~ n_n3462) ) ;
 assign wire7525 = ( n_n4060  &  (~ wire2247)  &  (~ wire6973) ) | ( n_n4060  &  (~ wire2247)  &  (~ wire6974) ) ;
 assign wire7526 = ( preset ) | ( (~ wire2268)  &  (~ wire6963)  &  wire7524 ) ;
 assign wire7527 = ( wire7526 ) | ( (~ n_n3833)  &  (~ n_n3903)  &  wire7525 ) ;
 assign wire7529 = ( (~ n_n4060)  &  (~ n_n3833)  &  n_n3903  &  (~ n_n3439) ) | ( n_n4060  &  (~ n_n3833)  &  (~ n_n3903)  &  (~ n_n3439) ) ;
 assign wire7532 = ( nld3_9 ) | ( (~ nak5_2)  &  nsr5_4  &  (~ nsr5_3) ) ;
 assign wire7533 = ( preset ) | ( pdn ) | ( (~ ndn3_8)  &  nsr3_9 ) ;
 assign wire7534 = ( nld3_9 ) | ( (~ nak5_2)  &  (~ nsr5_4)  &  nsr5_5 ) ;
 assign wire7535 = ( nld3_9 ) | ( (~ nak5_2)  &  nsr5_3  &  (~ nsr5_2) ) ;
 assign wire7537 = ( nld3_9 ) | ( (~ nak5_2)  &  (~ nsr5_5)  &  nsr5_7 ) ;
 assign wire7539 = ( nld3_9 ) | ( (~ nak5_2)  &  (~ nsr5_7)  &  nsr5_8 ) ;


endmodule

