module elliptic (
	tin_psv39_8_8_, tin_psv39_0_0_, tin_psv13_5_5_, tin_psv2_13_13_, tin_psv2_8_8_, pinp_2_2_, tin_psv38_2_2_, tin_psv33_5_5_, 
	tin_psv26_6_6_, tin_psv2_9_9_, pinp_3_3_, tin_psv18_2_2_, tin_psv39_9_9_, tin_psv39_1_1_, tin_psv13_6_6_, tin_psv2_6_6_, pinp_0_0_, tin_psv38_3_3_, 
	tin_psv33_6_6_, tin_psv26_13_13_, tin_psv26_12_12_, tin_psv26_7_7_, tin_psv2_7_7_, pinp_1_1_, preset_0_0_, tin_psv18_3_3_, tin_psv39_2_2_, tin_psv33_12_12_, 
	tin_psv33_11_11_, tin_psv33_10_10_, tin_psv13_7_7_, tin_psv2_10_10_, tin_psv38_4_4_, tin_psv39_10_10_, tin_psv33_7_7_, tin_psv26_15_15_, tin_psv26_14_14_, tin_psv26_8_8_, 
	tin_psv26_0_0_, tin_psv13_12_12_, tin_psv13_11_11_, tin_psv18_4_4_, tin_psv39_3_3_, tin_psv13_8_8_, tin_psv13_0_0_, pinp_15_15_, pinp_12_12_, tin_psv38_5_5_, 
	tin_psv33_8_8_, tin_psv33_0_0_, tin_psv26_9_9_, tin_psv26_1_1_, tin_psv13_10_10_, tin_psv18_5_5_, tin_psv39_4_4_, tin_psv13_9_9_, tin_psv13_1_1_, tin_psv2_15_15_, 
	tin_psv2_11_11_, tin_psv2_0_0_, tin_psv38_14_14_, tin_psv38_12_12_, tin_psv38_10_10_, tin_psv38_6_6_, tin_psv18_15_15_, tin_psv18_13_13_, tin_psv18_11_11_, tin_psv33_9_9_, 
	tin_psv33_1_1_, tin_psv26_2_2_, tin_psv2_1_1_, pclk, tin_psv38_15_15_, tin_psv38_11_11_, tin_psv18_12_12_, tin_psv18_6_6_, tin_psv39_5_5_, tin_psv13_2_2_, 
	pinp_14_14_, pinp_11_11_, pinp_8_8_, tin_psv38_7_7_, tin_psv39_12_12_, tin_psv39_11_11_, tin_psv33_2_2_, tin_psv26_3_3_, tin_psv13_14_14_, tin_psv13_13_13_, 
	pinp_9_9_, tin_psv18_10_10_, tin_psv18_7_7_, tin_psv39_6_6_, tin_psv33_15_15_, tin_psv33_14_14_, tin_psv33_13_13_, tin_psv13_3_3_, tin_psv2_14_14_, tin_psv2_12_12_, 
	tin_psv2_4_4_, pinp_6_6_, tin_psv38_8_8_, tin_psv38_0_0_, tin_psv39_14_14_, tin_psv39_13_13_, tin_psv33_3_3_, tin_psv26_11_11_, tin_psv26_10_10_, tin_psv26_4_4_, 
	tin_psv13_15_15_, tin_psv2_5_5_, pinp_7_7_, tin_psv18_8_8_, tin_psv18_0_0_, tin_psv39_7_7_, tin_psv13_4_4_, tin_psv2_2_2_, pinp_13_13_, pinp_10_10_, 
	pinp_4_4_, tin_psv38_9_9_, tin_psv38_1_1_, preset, tin_psv39_15_15_, tin_psv33_4_4_, tin_psv26_5_5_, tin_psv2_3_3_, pinp_5_5_, tin_psv38_13_13_, 
	tin_psv18_14_14_, tin_psv18_9_9_, tin_psv18_1_1_, psv39_8_8_, psv39_0_0_, psv13_5_5_, psv2_13_13_, psv2_8_8_, psv38_2_2_, psv33_5_5_, 
	psv26_6_6_, psv2_9_9_, psv18_2_2_, psv39_9_9_, psv39_1_1_, psv13_6_6_, psv2_6_6_, psv38_3_3_, psv33_6_6_, psv26_13_13_, 
	psv26_12_12_, psv26_7_7_, psv2_7_7_, psv18_3_3_, psv39_2_2_, psv33_12_12_, psv33_11_11_, psv33_10_10_, psv13_7_7_, psv2_10_10_, 
	psv38_4_4_, psv39_10_10_, psv33_7_7_, psv26_15_15_, psv26_14_14_, psv26_8_8_, psv26_0_0_, psv13_12_12_, psv13_11_11_, psv18_4_4_, 
	psv39_3_3_, psv13_8_8_, psv13_0_0_, psv38_5_5_, psv33_8_8_, psv33_0_0_, psv26_9_9_, psv26_1_1_, psv13_10_10_, psv18_5_5_, 
	psv39_4_4_, psv13_9_9_, psv13_1_1_, psv2_15_15_, psv2_11_11_, psv2_0_0_, psv38_14_14_, psv38_12_12_, psv38_10_10_, psv38_6_6_, 
	psv18_15_15_, psv18_13_13_, psv18_11_11_, psv33_9_9_, psv33_1_1_, psv26_2_2_, psv2_1_1_, psv38_15_15_, psv38_11_11_, psv18_12_12_, 
	psv18_6_6_, psv39_5_5_, psv13_2_2_, pover_0_0_, psv38_7_7_, psv39_12_12_, psv39_11_11_, psv33_2_2_, psv26_3_3_, psv13_14_14_, 
	psv13_13_13_, psv18_10_10_, psv18_7_7_, psv39_6_6_, psv33_15_15_, psv33_14_14_, psv33_13_13_, psv13_3_3_, psv2_14_14_, psv2_12_12_, 
	psv2_4_4_, psv38_8_8_, psv38_0_0_, pdn, psv39_14_14_, psv39_13_13_, psv33_3_3_, psv26_11_11_, psv26_10_10_, psv26_4_4_, 
	psv13_15_15_, psv2_5_5_, psv18_8_8_, psv18_0_0_, psv39_7_7_, psv13_4_4_, psv2_2_2_, psv38_9_9_, psv38_1_1_, psv39_15_15_, 
	psv33_4_4_, psv26_5_5_, psv2_3_3_, psv38_13_13_, psv18_14_14_, psv18_9_9_, psv18_1_1_);

input tin_psv39_8_8_;
input tin_psv39_0_0_;
input tin_psv13_5_5_;
input tin_psv2_13_13_;
input tin_psv2_8_8_;
input pinp_2_2_;
input tin_psv38_2_2_;
input tin_psv33_5_5_;
input tin_psv26_6_6_;
input tin_psv2_9_9_;
input pinp_3_3_;
input tin_psv18_2_2_;
input tin_psv39_9_9_;
input tin_psv39_1_1_;
input tin_psv13_6_6_;
input tin_psv2_6_6_;
input pinp_0_0_;
input tin_psv38_3_3_;
input tin_psv33_6_6_;
input tin_psv26_13_13_;
input tin_psv26_12_12_;
input tin_psv26_7_7_;
input tin_psv2_7_7_;
input pinp_1_1_;
input preset_0_0_;
input tin_psv18_3_3_;
input tin_psv39_2_2_;
input tin_psv33_12_12_;
input tin_psv33_11_11_;
input tin_psv33_10_10_;
input tin_psv13_7_7_;
input tin_psv2_10_10_;
input tin_psv38_4_4_;
input tin_psv39_10_10_;
input tin_psv33_7_7_;
input tin_psv26_15_15_;
input tin_psv26_14_14_;
input tin_psv26_8_8_;
input tin_psv26_0_0_;
input tin_psv13_12_12_;
input tin_psv13_11_11_;
input tin_psv18_4_4_;
input tin_psv39_3_3_;
input tin_psv13_8_8_;
input tin_psv13_0_0_;
input pinp_15_15_;
input pinp_12_12_;
input tin_psv38_5_5_;
input tin_psv33_8_8_;
input tin_psv33_0_0_;
input tin_psv26_9_9_;
input tin_psv26_1_1_;
input tin_psv13_10_10_;
input tin_psv18_5_5_;
input tin_psv39_4_4_;
input tin_psv13_9_9_;
input tin_psv13_1_1_;
input tin_psv2_15_15_;
input tin_psv2_11_11_;
input tin_psv2_0_0_;
input tin_psv38_14_14_;
input tin_psv38_12_12_;
input tin_psv38_10_10_;
input tin_psv38_6_6_;
input tin_psv18_15_15_;
input tin_psv18_13_13_;
input tin_psv18_11_11_;
input tin_psv33_9_9_;
input tin_psv33_1_1_;
input tin_psv26_2_2_;
input tin_psv2_1_1_;
input pclk;
input tin_psv38_15_15_;
input tin_psv38_11_11_;
input tin_psv18_12_12_;
input tin_psv18_6_6_;
input tin_psv39_5_5_;
input tin_psv13_2_2_;
input pinp_14_14_;
input pinp_11_11_;
input pinp_8_8_;
input tin_psv38_7_7_;
input tin_psv39_12_12_;
input tin_psv39_11_11_;
input tin_psv33_2_2_;
input tin_psv26_3_3_;
input tin_psv13_14_14_;
input tin_psv13_13_13_;
input pinp_9_9_;
input tin_psv18_10_10_;
input tin_psv18_7_7_;
input tin_psv39_6_6_;
input tin_psv33_15_15_;
input tin_psv33_14_14_;
input tin_psv33_13_13_;
input tin_psv13_3_3_;
input tin_psv2_14_14_;
input tin_psv2_12_12_;
input tin_psv2_4_4_;
input pinp_6_6_;
input tin_psv38_8_8_;
input tin_psv38_0_0_;
input tin_psv39_14_14_;
input tin_psv39_13_13_;
input tin_psv33_3_3_;
input tin_psv26_11_11_;
input tin_psv26_10_10_;
input tin_psv26_4_4_;
input tin_psv13_15_15_;
input tin_psv2_5_5_;
input pinp_7_7_;
input tin_psv18_8_8_;
input tin_psv18_0_0_;
input tin_psv39_7_7_;
input tin_psv13_4_4_;
input tin_psv2_2_2_;
input pinp_13_13_;
input pinp_10_10_;
input pinp_4_4_;
input tin_psv38_9_9_;
input tin_psv38_1_1_;
input preset;
input tin_psv39_15_15_;
input tin_psv33_4_4_;
input tin_psv26_5_5_;
input tin_psv2_3_3_;
input pinp_5_5_;
input tin_psv38_13_13_;
input tin_psv18_14_14_;
input tin_psv18_9_9_;
input tin_psv18_1_1_;
output psv39_8_8_;
output psv39_0_0_;
output psv13_5_5_;
output psv2_13_13_;
output psv2_8_8_;
output psv38_2_2_;
output psv33_5_5_;
output psv26_6_6_;
output psv2_9_9_;
output psv18_2_2_;
output psv39_9_9_;
output psv39_1_1_;
output psv13_6_6_;
output psv2_6_6_;
output psv38_3_3_;
output psv33_6_6_;
output psv26_13_13_;
output psv26_12_12_;
output psv26_7_7_;
output psv2_7_7_;
output psv18_3_3_;
output psv39_2_2_;
output psv33_12_12_;
output psv33_11_11_;
output psv33_10_10_;
output psv13_7_7_;
output psv2_10_10_;
output psv38_4_4_;
output psv39_10_10_;
output psv33_7_7_;
output psv26_15_15_;
output psv26_14_14_;
output psv26_8_8_;
output psv26_0_0_;
output psv13_12_12_;
output psv13_11_11_;
output psv18_4_4_;
output psv39_3_3_;
output psv13_8_8_;
output psv13_0_0_;
output psv38_5_5_;
output psv33_8_8_;
output psv33_0_0_;
output psv26_9_9_;
output psv26_1_1_;
output psv13_10_10_;
output psv18_5_5_;
output psv39_4_4_;
output psv13_9_9_;
output psv13_1_1_;
output psv2_15_15_;
output psv2_11_11_;
output psv2_0_0_;
output psv38_14_14_;
output psv38_12_12_;
output psv38_10_10_;
output psv38_6_6_;
output psv18_15_15_;
output psv18_13_13_;
output psv18_11_11_;
output psv33_9_9_;
output psv33_1_1_;
output psv26_2_2_;
output psv2_1_1_;
output psv38_15_15_;
output psv38_11_11_;
output psv18_12_12_;
output psv18_6_6_;
output psv39_5_5_;
output psv13_2_2_;
output pover_0_0_;
output psv38_7_7_;
output psv39_12_12_;
output psv39_11_11_;
output psv33_2_2_;
output psv26_3_3_;
output psv13_14_14_;
output psv13_13_13_;
output psv18_10_10_;
output psv18_7_7_;
output psv39_6_6_;
output psv33_15_15_;
output psv33_14_14_;
output psv33_13_13_;
output psv13_3_3_;
output psv2_14_14_;
output psv2_12_12_;
output psv2_4_4_;
output psv38_8_8_;
output psv38_0_0_;
output pdn;
output psv39_14_14_;
output psv39_13_13_;
output psv33_3_3_;
output psv26_11_11_;
output psv26_10_10_;
output psv26_4_4_;
output psv13_15_15_;
output psv2_5_5_;
output psv18_8_8_;
output psv18_0_0_;
output psv39_7_7_;
output psv13_4_4_;
output psv2_2_2_;
output psv38_9_9_;
output psv38_1_1_;
output psv39_15_15_;
output psv33_4_4_;
output psv26_5_5_;
output psv2_3_3_;
output psv38_13_13_;
output psv18_14_14_;
output psv18_9_9_;
output psv18_1_1_;
wire n_n9279;
wire n_n8265;
wire n_n8264;
wire n_n7724;
wire n_n8190;
wire n_n7893;
wire n_n9149;
wire n_n7216;
wire n_n7778;
wire n_n8834;
wire n_n8149;
wire n_n7034;
wire n_n7166;
wire n_n7868;
wire n_n8590;
wire n_n8870;
wire n_n7251;
wire n_n7269;
wire n_n6990;
wire n_n7671;
wire n_n7412;
wire n_n7201;
wire n_n7524;
wire n_n9545;
wire n_n9466;
wire n_n7205;
wire n_n6949;
wire n_n7077;
wire n_n7243;
wire n_n7369;
wire n_n8189;
wire n_n7123;
wire n_n9579;
wire n_n6944;
wire n_n6994;
wire n_n9234;
wire n_n7521;
wire n_n7229;
wire n_n9084;
wire n_n7416;
wire n_n7066;
wire n_n8774;
wire n_n7438;
wire n_n8409;
wire n_n8207;
wire n_n8376;
wire n_n7028;
wire n_n7421;
wire n_n7753;
wire n_n7680;
wire n_n7669;
wire n_n7455;
wire n_n6989;
wire n_n8596;
wire n_n7472;
wire n_n8393;
wire n_n7591;
wire n_n7481;
wire n_n9140;
wire n_n7331;
wire n_n8757;
wire n_n7422;
wire n_n7040;
wire n_n7277;
wire n_n9007;
wire n_n7580;
wire n_n7067;
wire n_n7092;
wire n_n7199;
wire n_n8598;
wire n_n7240;
wire n_n7382;
wire n_n8411;
wire n_n7147;
wire n_n7517;
wire n_n9250;
wire n_n7188;
wire n_n8612;
wire n_n8532;
wire n_n8698;
wire n_n8608;
wire n_n8307;
wire n_n8654;
wire n_n7125;
wire n_n7357;
wire n_n7;
wire n_n8787;
wire n_n8785;
wire n_n7473;
wire n_n7214;
wire n_n7063;
wire n_n9472;
wire n_n8999;
wire n_n7495;
wire n_n7266;
wire n_n8507;
wire n_n9634;
wire n_n7189;
wire n_n8700;
wire n_n9105;
wire n_n7408;
wire n_n7137;
wire n_n7504;
wire n_n8527;
wire n_n9208;
wire n_n7177;
wire n_n7615;
wire n_n7087;
wire n_n8293;
wire n_n8217;
wire n_n9538;
wire n_n7091;
wire n_n8487;
wire n_n8299;
wire n_n7796;
wire n_n8130;
wire n_n8660;
wire n_n7325;
wire n_n8332;
wire n_n7037;
wire n_n7797;
wire n_n7005;
wire n_n7200;
wire n_n9527;
wire n_n7523;
wire n_n8250;
wire n_n7483;
wire n_n8481;
wire n_n7451;
wire n_n7055;
wire n_n7555;
wire n_n9063;
wire n_n7207;
wire n_n7100;
wire n_n7799;
wire n_n7471;
wire n_n7219;
wire n_n7614;
wire n_n7250;
wire n_n7590;
wire n_n6915;
wire n_n8052;
wire n_n9014;
wire n_n8065;
wire n_n9517;
wire n_n8089;
wire n_n9256;
wire n_n8174;
wire n_n8490;
wire n_n8113;
wire n_n7039;
wire n_n7095;
wire n_n8034;
wire n_n7094;
wire n_n8242;
wire n_n7855;
wire n_n7098;
wire n_n7632;
wire n_n9079;
wire n_n7090;
wire n_n7299;
wire n_n9480;
wire n_n9409;
wire n_n7385;
wire n_n7406;
wire n_n7405;
wire n_n7782;
wire n_n7372;
wire n_n7053;
wire n_n7086;
wire n_n8730;
wire n_n1;
wire n_n9090;
wire n_n7547;
wire n_n8335;
wire n_n7323;
wire n_n9610;
wire n_n8111;
wire n_n8039;
wire n_n9617;
wire n_n9612;
wire n_n9241;
wire n_n7383;
wire n_n6933;
wire n_n7461;
wire n_n7613;
wire n_n8764;
wire n_n7014;
wire n_n7897;
wire n_n8379;
wire n_n8861;
wire n_n8036;
wire n_n8026;
wire n_n7883;
wire n_n8973;
wire n_n7285;
wire n_n9222;
wire n_n8147;
wire n_n9167;
wire n_n8310;
wire n_n8317;
wire n_n7168;
wire n_n7397;
wire n_n7165;
wire n_n7070;
wire n_n8109;
wire n_n7268;
wire n_n8567;
wire n_n7228;
wire n_n7718;
wire n_n7494;
wire n_n7235;
wire n_n8218;
wire n_n9567;
wire n_n9199;
wire n_n8544;
wire n_n6934;
wire n_n6914;
wire n_n8735;
wire n_n8474;
wire n_n8498;
wire n_n8085;
wire n_n7802;
wire n_n7061;
wire n_n9097;
wire n_n7159;
wire n_n7303;
wire n_n9565;
wire n_n7833;
wire n_n8413;
wire n_n6969;
wire n_n8345;
wire n_n7800;
wire n_n7172;
wire n_n7212;
wire n_n7545;
wire n_n7099;
wire n_n8997;
wire n_n7479;
wire n_n9463;
wire n_n8346;
wire n_n8874;
wire n_n7354;
wire n_n8958;
wire n_n8956;
wire n_n8246;
wire n_n8257;
wire n_n7404;
wire n_n8842;
wire n_n8443;
wire n_n7163;
wire n_n6;
wire n_n8025;
wire n_n7982;
wire n_n7186;
wire n_n7248;
wire n_n7639;
wire n_n8347;
wire n_n8835;
wire n_n8444;
wire n_n7425;
wire n_n7830;
wire n_n7618;
wire n_n9062;
wire n_n9430;
wire n_n8676;
wire n_n8023;
wire n_n7141;
wire n_n8995;
wire n_n7917;
wire n_n8259;
wire n_n9207;
wire n_n9188;
wire n_n9094;
wire n_n8179;
wire n_n7773;
wire n_n7647;
wire n_n7038;
wire n_n7157;
wire n_n8940;
wire n_n8041;
wire n_n8679;
wire n_n8658;
wire n_n9109;
wire n_n9572;
wire n_n8950;
wire n_n9240;
wire n_n9386;
wire n_n7594;
wire n_n7210;
wire n_n8405;
wire n_n7892;
wire n_n7221;
wire n_n7350;
wire n_n8465;
wire n_n6983;
wire n_n7719;
wire n_n7551;
wire n_n8737;
wire n_n7361;
wire n_n9299;
wire n_n9549;
wire n_n9287;
wire n_n8776;
wire n_n7009;
wire n_n7355;
wire n_n7776;
wire n_n7550;
wire n_n8172;
wire n_n7497;
wire n_n9146;
wire n_n8752;
wire n_n8771;
wire n_n8048;
wire n_n7870;
wire n_n7015;
wire n_n7470;
wire n_n9002;
wire n_n7532;
wire n_n7442;
wire n_n9078;
wire n_n8367;
wire n_n9330;
wire n_n7103;
wire n_n8399;
wire n_n7526;
wire n_n9035;
wire n_n7264;
wire n_n8696;
wire n_n7080;
wire n_n7290;
wire n_n11;
wire n_n2;
wire n_n7548;
wire n_n7294;
wire n_n8949;
wire n_n7633;
wire n_n8934;
wire n_n9243;
wire n_n7194;
wire n_n7465;
wire n_n8610;
wire n_n7746;
wire n_n7349;
wire n_n8169;
wire n_n7316;
wire n_n8495;
wire n_n6995;
wire n_n7468;
wire n_n7049;
wire n_n7304;
wire n_n7139;
wire n_n7142;
wire n_n6947;
wire n_n8548;
wire n_n9543;
wire n_n9620;
wire n_n7101;
wire n_n8092;
wire n_n8624;
wire n_n8380;
wire n_n6965;
wire n_n7891;
wire n_n8907;
wire n_n7571;
wire n_n7559;
wire n_n7612;
wire n_n8985;
wire n_n8890;
wire n_n7999;
wire n_n7220;
wire n_n8748;
wire n_n6942;
wire n_n9367;
wire n_n8518;
wire n_n6955;
wire n_n8297;
wire n_n6922;
wire n_n7016;
wire n_n8637;
wire n_n9551;
wire n_n8286;
wire n_n8015;
wire n_n7345;
wire n_n7010;
wire n_n8587;
wire n_n7097;
wire n_n6953;
wire n_n8457;
wire n_n7940;
wire n_n8163;
wire n_n8860;
wire n_n7319;
wire n_n5;
wire n_n6924;
wire n_n8614;
wire n_n6941;
wire n_n7000;
wire n_n7280;
wire n_n8137;
wire n_n7313;
wire n_n7832;
wire n_n8021;
wire n_n8517;
wire n_n8136;
wire n_n7122;
wire n_n7616;
wire n_n8684;
wire n_n9529;
wire n_n9509;
wire n_n7042;
wire n_n8479;
wire n_n8542;
wire n_n7088;
wire n_n7096;
wire n_n8878;
wire n_n8331;
wire n_n7301;
wire n_n7972;
wire n_n6951;
wire n_n8863;
wire n_n6993;
wire n_n7057;
wire n_n7143;
wire n_n6945;
wire n_n9101;
wire n_n7307;
wire n_n7300;
wire n_n7036;
wire n_n8759;
wire n_n6911;
wire n_n7352;
wire n_n7535;
wire n_n7457;
wire n_n8703;
wire n_n7520;
wire n_n8475;
wire n_n8429;
wire n_n9018;
wire n_n7698;
wire n_n6972;
wire n_n7480;
wire n_n8338;
wire n_n7213;
wire n_n6960;
wire n_n9427;
wire n_n7478;
wire n_n7060;
wire n_n7318;
wire n_n8967;
wire n_n9369;
wire n_n7320;
wire n_n7867;
wire n_n9372;
wire n_n10;
wire n_n6940;
wire n_n6925;
wire n_n7007;
wire n_n6936;
wire n_n7198;
wire n_n8547;
wire n_n6954;
wire n_n9622;
wire n_n9469;
wire n_n7569;
wire n_n7339;
wire n_n9364;
wire n_n7180;
wire n_n8738;
wire n_n6932;
wire n_n7255;
wire n_n7519;
wire n_n7486;
wire n_n7259;
wire n_n8460;
wire n_n7987;
wire n_n8378;
wire n_n8724;
wire n_n8625;
wire n_n9082;
wire n_n8209;
wire n_n7414;
wire n_n8899;
wire n_n7477;
wire n_n8761;
wire n_n7996;
wire n_n8094;
wire n_n7112;
wire n_n7386;
wire n_n8768;
wire n_n7611;
wire n_n7834;
wire n_n9156;
wire n_n8551;
wire n_n7380;
wire n_n9445;
wire n_n8632;
wire n_n7353;
wire n_n7309;
wire n_n8401;
wire n_n7488;
wire n_n7733;
wire n_n8503;
wire n_n8455;
wire n_n7512;
wire n_n7314;
wire n_n9474;
wire n_n8275;
wire n_n8832;
wire n_n7921;
wire n_n7105;
wire n_n9511;
wire n_n8763;
wire n_n4;
wire n_n7153;
wire n_n8754;
wire n_n7592;
wire n_n8853;
wire n_n8620;
wire n_n9214;
wire n_n8987;
wire n_n7895;
wire n_n8071;
wire n_n8969;
wire n_n8714;
wire n_n8485;
wire n_n7245;
wire n_n7865;
wire n_n8336;
wire n_n7634;
wire n_n7508;
wire n_n7359;
wire n_n8559;
wire n_n9107;
wire n_n9285;
wire n_n7460;
wire n_n8540;
wire n_n7296;
wire n_n7192;
wire n_n7058;
wire n_n7297;
wire n_n9213;
wire n_n7370;
wire n_n8463;
wire n_n7658;
wire n_n7238;
wire n_n7109;
wire n_n8690;
wire n_n6943;
wire n_n9326;
wire n_n7994;
wire n_n7394;
wire n_n7589;
wire n_n7506;
wire n_n7958;
wire n_n7503;
wire n_n8008;
wire n_n7562;
wire n_n7223;
wire n_n8105;
wire n_n7456;
wire n_n7043;
wire n_n7279;
wire n_n8960;
wire n_n8013;
wire n_n9276;
wire n_n9086;
wire n_n7542;
wire n_n7448;
wire n_n8164;
wire n_n8478;
wire n_n9415;
wire n_n9;
wire n_n0;
wire n_n7025;
wire n_n8855;
wire n_n7894;
wire n_n7249;
wire n_n7984;
wire n_n8311;
wire n_n7230;
wire n_n7317;
wire n_n8799;
wire n_n8682;
wire n_n9425;
wire n_n8244;
wire n_n9457;
wire n_n9301;
wire n_n7391;
wire n_n6962;
wire n_n6916;
wire n_n7224;
wire n_n7505;
wire n_n7169;
wire n_n6970;
wire n_n8176;
wire n_n8388;
wire n_n7998;
wire n_n7595;
wire n_n6996;
wire n_n7263;
wire n_n7979;
wire n_n6992;
wire n_n7675;
wire n_n8395;
wire n_n9532;
wire n_n7208;
wire n_n7002;
wire n_n7004;
wire n_n7623;
wire n_n8790;
wire n_n7253;
wire n_n7161;
wire n_n7943;
wire n_n6997;
wire n_n8098;
wire n_n6987;
wire n_n6985;
wire n_n8926;
wire n_n7116;
wire n_n8372;
wire n_n7379;
wire n_n9218;
wire n_n7048;
wire n_n8080;
wire n_n7131;
wire n_n8709;
wire n_n7621;
wire n_n7340;
wire n_n7114;
wire n_n7032;
wire n_n9088;
wire n_n9185;
wire n_n8129;
wire n_n7564;
wire n_n7018;
wire n_n8309;
wire n_n7260;
wire n_n7839;
wire n_n7619;
wire n_n7992;
wire n_n7138;
wire n_n8252;
wire n_n8888;
wire n_n7234;
wire n_n8917;
wire n_n7501;
wire n_n7084;
wire n_n8074;
wire n_n7337;
wire n_n8103;
wire n_n8170;
wire n_n9058;
wire n_n9022;
wire n_n7152;
wire n_n8952;
wire n_n6919;
wire n_n8830;
wire n_n8440;
wire n_n8231;
wire n_n9251;
wire n_n7981;
wire n_n8565;
wire n_n9461;
wire n_n7560;
wire n_n8922;
wire n_n7977;
wire n_n7828;
wire n_n7170;
wire n_n8712;
wire n_n8943;
wire n_n7371;
wire n_n7215;
wire n_n7027;
wire n_n6982;
wire n_n7115;
wire n_n7072;
wire n_n7445;
wire n_n7963;
wire n_n7348;
wire n_n8897;
wire n_n7974;
wire n_n7648;
wire n_n7035;
wire n_n7960;
wire n_n7423;
wire n_n7475;
wire n_n8766;
wire n_n9032;
wire n_n8829;
wire n_n8186;
wire n_n9120;
wire n_n8059;
wire n_n7801;
wire n_n7450;
wire n_n9204;
wire n_n8391;
wire n_n7538;
wire n_n8374;
wire n_n8327;
wire n_n9297;
wire n_n7062;
wire n_n8505;
wire n_n7729;
wire n_n7226;
wire n_n7419;
wire n_n7957;
wire n_n7945;
wire n_n7662;
wire n_n8254;
wire n_n9037;
wire n_n7282;
wire n_n7082;
wire n_n7388;
wire n_n9001;
wire n_n6967;
wire n_n8451;
wire n_n7044;
wire n_n7012;
wire n_n9625;
wire n_n7132;
wire n_n8645;
wire n_n8802;
wire n_n9569;
wire n_n8365;
wire n_n7104;
wire n_n7785;
wire n_n7006;
wire n_n7275;
wire n_n9211;
wire n_n8382;
wire n_n9453;
wire n_n8434;
wire n_n7574;
wire n_n6981;
wire n_n6966;
wire n_n7700;
wire n_n7126;
wire n_n8424;
wire n_n9103;
wire n_n9220;
wire n_n9447;
wire n_n8593;
wire n_n7233;
wire n_n7466;
wire n_n8232;
wire n_n7167;
wire n_n8063;
wire n_n9039;
wire n_n7916;
wire n_n8054;
wire n_n7267;
wire n_n8255;
wire n_n7924;
wire n_n7502;
wire n_n7258;
wire n_n7262;
wire n_n7705;
wire n_n7293;
wire n_n9419;
wire n_n7625;
wire n_n7093;
wire n_n8261;
wire n_n8442;
wire n_n7516;
wire n_n6923;
wire n_n7587;
wire n_n9122;
wire n_n9158;
wire n_n8859;
wire n_n8043;
wire n_n7727;
wire n_n8722;
wire n_n7399;
wire n_n9354;
wire n_n7211;
wire n_n8469;
wire n_n7312;
wire n_n8795;
wire n_n9116;
wire n_n7989;
wire n_n8780;
wire n_n8816;
wire n_n9111;
wire n_n9091;
wire n_n6938;
wire n_n8212;
wire n_n7593;
wire n_n8686;
wire n_n7836;
wire n_n6939;
wire n_n9202;
wire n_n7113;
wire n_n8945;
wire n_n7051;
wire n_n9614;
wire n_n8472;
wire n_n6935;
wire n_n7237;
wire n_n7204;
wire n_n7525;
wire n_n9020;
wire n_n7780;
wire n_n6931;
wire n_n7107;
wire n_n7489;
wire n_n7265;
wire n_n8546;
wire n_n7046;
wire n_n8220;
wire n_n7396;
wire n_n7899;
wire n_n9229;
wire n_n7515;
wire n_n6929;
wire n_n6917;
wire n_n8501;
wire n_n8432;
wire n_n7631;
wire n_n9038;
wire n_n7410;
wire n_n7326;
wire n_n7134;
wire n_n7068;
wire n_n8616;
wire n_n7241;
wire n_n8229;
wire n_n9293;
wire n_n8248;
wire n_n8971;
wire n_n7073;
wire n_n7492;
wire n_n8289;
wire n_n7184;
wire n_n7162;
wire n_n7490;
wire n_n8291;
wire n_n8731;
wire n_n8046;
wire n_n9628;
wire n_n6918;
wire n_n9507;
wire n_n9154;
wire n_n7377;
wire n_n8994;
wire n_n7690;
wire n_n7608;
wire n_n8184;
wire n_n7529;
wire n_n8838;
wire n_n7902;
wire n_n9138;
wire n_n9074;
wire n_n7449;
wire n_n6977;
wire n_n7151;
wire n_n7747;
wire n_n7145;
wire n_n7056;
wire n_n7175;
wire n_n8476;
wire n_n8412;
wire n_n8635;
wire n_n7182;
wire n_n8656;
wire n_n8483;
wire n_n6946;
wire n_n7530;
wire n_n8534;
wire n_n8618;
wire n_n8908;
wire n_n7596;
wire n_n9118;
wire n_n7534;
wire n_n8914;
wire n_n8728;
wire n_n8385;
wire n_n8778;
wire n_n6979;
wire n_n7714;
wire n_n9066;
wire n_n7059;
wire n_n7400;
wire n_n7247;
wire n_n8689;
wire n_n8788;
wire n_n8553;
wire n_n7528;
wire n_n7292;
wire n_n8669;
wire n_n8642;
wire n_n6998;
wire n_n8187;
wire n_n7029;
wire n_n9065;
wire n_n7364;
wire n_n8359;
wire n_n9227;
wire n_n8919;
wire n_n8509;
wire n_n8837;
wire n_n8639;
wire n_n9422;
wire n_n8356;
wire n_n3;
wire n_n7447;
wire n_n8467;
wire n_n7120;
wire n_n7482;
wire n_n7232;
wire n_n8500;
wire n_n7351;
wire n_n8038;
wire n_n8814;
wire n_n8407;
wire n_n8576;
wire n_n7078;
wire n_n8827;
wire n_n8767;
wire n_n8585;
wire n_n7900;
wire n_n8627;
wire n_n7750;
wire n_n7118;
wire n_n8181;
wire n_n8062;
wire n_n8851;
wire n_n6930;
wire n_n8010;
wire n_n7716;
wire n_n8325;
wire n_n7193;
wire n_n8343;
wire n_n8295;
wire n_n8115;
wire n_n8266;
wire n_n7563;
wire n_n9060;
wire n_n9206;
wire n_n7278;
wire n_n9080;
wire n_n6909;
wire n_n8726;
wire n_n7672;
wire n_n7329;
wire n_n8965;
wire n_n7841;
wire n_n8283;
wire n_n9374;
wire n_n7171;
wire n_n6927;
wire n_n7071;
wire n_n8144;
wire n_n8437;
wire n_n6999;
wire n_n8117;
wire n_n7610;
wire n_n9238;
wire n_n9236;
wire n_n6913;
wire n_n9443;
wire n_n9521;
wire n_n7518;
wire n_n7433;
wire n_n8664;
wire n_n8318;
wire n_n8301;
wire n_n7020;
wire n_n8133;
wire n_n8896;
wire n_n7149;
wire n_n9454;
wire n_n8370;
wire n_n8;
wire n_n7047;
wire n_n8836;
wire n_n7443;
wire n_n7158;
wire n_n7128;
wire n_n7676;
wire n_n8101;
wire n_n9224;
wire n_n8461;
wire n_n8087;
wire n_n9024;
wire n_n8178;
wire n_n7660;
wire n_n8107;
wire n_n8920;
wire n_n7858;
wire n_n7731;
wire n_n7427;
wire n_n9519;
wire n_n6964;
wire n_n7677;
wire n_n7222;
wire n_n7679;
wire n_n8840;
wire n_n7335;
wire n_n7197;
wire n_n7754;
wire n_n7195;
wire n_n8769;
wire n_n8422;
wire n_n7085;
wire n_n9524;
wire n_n8032;
wire n_n7533;
wire n_n7426;
wire n_n9231;
wire n_n7257;
wire n_n9562;
wire n_n8671;
wire n_n7106;
wire n_n7008;
wire n_n8755;
wire n_n8640;
wire n_n8191;
wire n_n8057;
wire n_n7439;
wire n_n9305;
wire n_n6928;
wire n_n8848;
wire n_n9209;
wire n_n8122;
wire n_n7254;
wire n_n8050;
wire n_n7135;
wire n_n7081;
wire n_n9005;
wire n_n7407;
wire n_n7904;
wire n_n7030;
wire n_n7064;
wire n_n8211;
wire n_n7023;
wire n_n7585;
wire n_n8415;
wire n_n8166;
wire n_n8140;
wire n_n7446;
wire n_n8120;
wire n_n8162;
wire n_n8337;
wire n_n8194;
wire n_n9515;
wire n_n9076;
wire n_n8363;
wire n_n8773;
wire n_n7089;
wire n_n7840;
wire n_n7321;
wire n_n8873;
wire n_n7745;
wire n_n7001;
wire n_n6959;
wire n_n7196;
wire n_n8205;
wire n_n7367;
wire n_n8818;
wire n_n7110;
wire n_n7804;
wire n_n8494;
wire n_n7206;
wire n_n8872;
wire n_n8364;
wire n_n8496;
wire n_n6971;
wire n_n8453;
wire n_n7413;
wire n_n9504;
wire n_n8825;
wire n_n9631;
wire n_n7075;
wire n_n7469;
wire n_n8634;
wire n_n9577;
wire n_n8134;
wire n_n9328;
wire n_n7499;
wire n_n6973;
wire n_n8604;
wire n_n9295;
wire n_n7155;
wire n_n7919;
wire n_n8893;
wire n_n7620;
wire n_n8138;
wire n_n9274;
wire n_n7202;
wire n_n7805;
wire n_n7343;
wire n_n6975;
wire n_n6958;
wire n_n7617;
wire n_n7646;
wire n_n9012;
wire n_n7287;
wire n_n8077;
wire n_n7333;
wire n_n6957;
wire n_n7496;
wire n_n8525;
wire n_n7795;
wire n_n7851;
wire n_n8446;
wire n_n7484;
wire n_n7305;
wire n_n6921;
wire n_n7191;
wire n_n6926;
wire n_n8489;
wire n_n8947;
wire n_n8471;
wire n_n8215;
wire n_n8180;
wire n_n7295;
wire n_n7437;
wire n_n9143;
wire n_n8426;
wire n_n8558;
wire n_n7838;
wire wire2421;
wire wire2371;
wire nrq3_11;
wire n_n9616;
wire ndn_latch3_12;
wire wire2405;
wire ndn_latch3_26;
wire nrq3_9;
wire wire2370;
wire nrq3_39;
wire wire2408;
wire wire2363;
wire wire2395;
wire wire2453;
wire ndn_latch3_27;
wire nrq3_34;
wire wire2369;
wire wire2469;
wire wire2368;
wire wire2436;
wire nrq3_19;
wire wire2367;
wire wire2447;
wire n_n9581;
wire ndn_latch3_29;
wire n_n8979;
wire n_n7432;
wire n_n8323;
wire wire2402;
wire nrq3_4;
wire nrq3_16;
wire nrq3_36;
wire nrq3_18;
wire wire2404;
wire ndn_latch3_7;
wire ndn_latch3_32;
wire nrq3_15;
wire nrq3_17;
wire wire2431;
wire n_n7378;
wire nrq3_21;
wire wire2418;
wire n_n9619;
wire wire2406;
wire ndn_latch3_25;
wire wire2423;
wire wire2427;
wire ndn_latch3_28;
wire n_n8880;
wire n_n8431;
wire n_n8783;
wire wire2429;
wire n_n9056;
wire wire2451;
wire n_n8403;
wire n_n8630;
wire ngfdn_2;
wire n_n9246;
wire n_n9564;
wire n_n9633;
wire n_n8522;
wire n_n8521;
wire n_n8538;
wire n_n8963;
wire n_n8537;
wire n_n8653;
wire n_n8706;
wire n_n8484;
wire n_n8708;
wire n_n8418;
wire n_n8353;
wire n_n8355;
wire n_n9356;
wire n_n8734;
wire n_n8733;
wire wire2460;
wire n_n8784;
wire n_n8373;
wire n_n7864;
wire n_n8876;
wire n_n9072;
wire n_n7787;
wire n_n8976;
wire n_n7637;
wire n_n9553;
wire n_n9627;
wire n_n8450;
wire n_n8448;
wire n_n8324;
wire n_n8820;
wire n_n8936;
wire n_n8740;
wire n_n8822;
wire n_n8807;
wire n_n9216;
wire n_n8606;
wire n_n9010;
wire n_n8823;
wire n_n9029;
wire n_n9288;
wire n_n9114;
wire n_n9435;
wire n_n9152;
wire n_n8846;
wire nen3_2;
wire n_n8806;
wire n_n8420;
wire n_n7543;
wire n_n8694;
wire n_n9385;
wire n_n9384;
wire nrq2_9;
wire wire2372;
wire wire2373;
wire wire2374;
wire wire2375;
wire wire2377;
wire wire2380;
wire wire2381;
wire wire2383;
wire n_n9583;
wire n_n7997;
wire n_n9639;
wire n_n8493;
wire n_n8019;
wire n_n7573;
wire n_n7869;
wire n_n8028;
wire n_n8953;
wire n_n9197;
wire n_n8667;
wire n_n7566;
wire n_n8154;
wire n_n7818;
wire n_n7597;
wire n_n8314;
wire n_n9040;
wire n_n9307;
wire n_n9332;
wire n_n8321;
wire n_n7311;
wire n_n7544;
wire n_n8320;
wire n_n8156;
wire n_n8155;
wire n_n9124;
wire n_n9389;
wire n_n7784;
wire n_n7872;
wire n_n8126;
wire n_n8125;
wire n_n9478;
wire n_n8865;
wire n_n8579;
wire n_n8342;
wire n_n8932;
wire n_n7274;
wire n_n7218;
wire n_n8315;
wire n_n7939;
wire n_n8204;
wire n_n8316;
wire n_n9258;
wire n_n9587;
wire wire2364;
wire wire2379;
wire wire2382;
wire wire2470;
wire wire2471;
wire wire2472;
wire wire2474;
wire wire2475;
wire wire2480;
wire wire2482;
wire wire2484;
wire wire2485;
wire wire2488;
wire wire2490;
wire wire2492;
wire wire2493;
wire wire2494;
wire wire2498;
wire wire2502;
wire wire2504;
wire wire2505;
wire wire2506;
wire wire2508;
wire wire2509;
wire wire2512;
wire wire2513;
wire wire2514;
wire wire2516;
wire wire2517;
wire wire2518;
wire wire2519;
wire wire2522;
wire wire2524;
wire wire2525;
wire wire2526;
wire wire2528;
wire wire2529;
wire wire2532;
wire wire2534;
wire wire2535;
wire wire2542;
wire wire2543;
wire wire2544;
wire wire2545;
wire wire2548;
wire wire2549;
wire wire2550;
wire wire2554;
wire wire2558;
wire wire2559;
wire wire2564;
wire wire2565;
wire wire2568;
wire wire2569;
wire wire2570;
wire wire2571;
wire wire2572;
wire wire2573;
wire wire2576;
wire wire2578;
wire wire2580;
wire wire2581;
wire wire2584;
wire wire2586;
wire wire2588;
wire wire2590;
wire wire2591;
wire wire2592;
wire wire2593;
wire wire2594;
wire wire2595;
wire wire2596;
wire wire2597;
wire wire2598;
wire wire2606;
wire wire2607;
wire wire2612;
wire wire2613;
wire wire2614;
wire wire2615;
wire wire2630;
wire wire2634;
wire wire2635;
wire wire2638;
wire wire2640;
wire wire2641;
wire wire2648;
wire wire2649;
wire wire2655;
wire wire2656;
wire wire2657;
wire wire2659;
wire wire2660;
wire wire2665;
wire wire2673;
wire wire2675;
wire wire2676;
wire wire2679;
wire wire2680;
wire wire2683;
wire wire2684;
wire wire2687;
wire wire2688;
wire wire2691;
wire wire2697;
wire wire2698;
wire wire2701;
wire wire2702;
wire wire2703;
wire wire2704;
wire wire2705;
wire wire2709;
wire wire2711;
wire wire2712;
wire wire2713;
wire wire2715;
wire wire2716;
wire wire2717;
wire wire2718;
wire wire2719;
wire wire2721;
wire wire2722;
wire wire2725;
wire wire2727;
wire wire2731;
wire wire2732;
wire wire2735;
wire wire2736;
wire wire2737;
wire wire2738;
wire wire2743;
wire wire2744;
wire wire2747;
wire wire2748;
wire wire2749;
wire wire2751;
wire wire2752;
wire wire2755;
wire wire2757;
wire wire2758;
wire wire2762;
wire wire2763;
wire wire2764;
wire wire2768;
wire wire2769;
wire wire2772;
wire wire2773;
wire wire2774;
wire wire2775;
wire wire2776;
wire wire2777;
wire wire2780;
wire wire2781;
wire wire2782;
wire wire2783;
wire wire2784;
wire wire2788;
wire wire2790;
wire wire2792;
wire wire2794;
wire wire2796;
wire wire2798;
wire wire2799;
wire wire2800;
wire wire2801;
wire wire2806;
wire wire2807;
wire wire2809;
wire wire2810;
wire wire2811;
wire wire2812;
wire wire2813;
wire wire2814;
wire wire2819;
wire wire2820;
wire wire2821;
wire wire2823;
wire wire2824;
wire wire2825;
wire wire2827;
wire wire2828;
wire wire2831;
wire wire2833;
wire wire2835;
wire wire2836;
wire wire2837;
wire wire2838;
wire wire2841;
wire wire2842;
wire wire2845;
wire wire2846;
wire wire2847;
wire wire2851;
wire wire2855;
wire wire2856;
wire wire2857;
wire wire2864;
wire wire2865;
wire wire2869;
wire wire2870;
wire wire2871;
wire wire2872;
wire wire2875;
wire wire2876;
wire wire2879;
wire wire2885;
wire wire2886;
wire wire2891;
wire wire2892;
wire wire2895;
wire wire2897;
wire wire2898;
wire wire2903;
wire wire2904;
wire wire2907;
wire wire2908;
wire wire2909;
wire wire2910;
wire wire2915;
wire wire2916;
wire wire2917;
wire wire2918;
wire wire2919;
wire wire2925;
wire wire2929;
wire wire2930;
wire wire2931;
wire wire2932;
wire wire2933;
wire wire2935;
wire wire2937;
wire wire2938;
wire wire2939;
wire wire2941;
wire wire2942;
wire wire2943;
wire wire2945;
wire wire2946;
wire wire2949;
wire wire2951;
wire wire2953;
wire wire2954;
wire wire2955;
wire wire2956;
wire wire2957;
wire wire2958;
wire wire2961;
wire wire2962;
wire wire2965;
wire wire2966;
wire wire2967;
wire wire2968;
wire wire2969;
wire wire2970;
wire wire2974;
wire wire2975;
wire wire2976;
wire wire2977;
wire wire2978;
wire wire2979;
wire wire2980;
wire wire2981;
wire wire2984;
wire wire2985;
wire wire2988;
wire wire2989;
wire wire2992;
wire wire2994;
wire wire2995;
wire wire2998;
wire wire3000;
wire wire3001;
wire wire3002;
wire wire3004;
wire wire3006;
wire wire3010;
wire wire3014;
wire wire3018;
wire wire3019;
wire wire3025;
wire wire3026;
wire wire3027;
wire wire3028;
wire wire3032;
wire wire3034;
wire wire3037;
wire wire3038;
wire wire3041;
wire wire3045;
wire wire3046;
wire wire3049;
wire wire3051;
wire wire3052;
wire wire3053;
wire wire3055;
wire wire3056;
wire wire3059;
wire wire3060;
wire wire3061;
wire wire3062;
wire wire3065;
wire wire3066;
wire wire3067;
wire wire3068;
wire wire3073;
wire wire3074;
wire wire3075;
wire wire3081;
wire wire3082;
wire wire3085;
wire wire3086;
wire wire3087;
wire wire3088;
wire wire3091;
wire wire3095;
wire wire3101;
wire wire3102;
wire wire3107;
wire wire3108;
wire wire3113;
wire wire3114;
wire wire3117;
wire wire3121;
wire wire3122;
wire wire3123;
wire wire3125;
wire wire3126;
wire wire3127;
wire wire3128;
wire wire3129;
wire wire3131;
wire wire3132;
wire wire3135;
wire wire3139;
wire wire3140;
wire wire3143;
wire wire3155;
wire wire3157;
wire wire3158;
wire wire3165;
wire wire3167;
wire wire3168;
wire wire3171;
wire wire3177;
wire wire3178;
wire wire3179;
wire wire3183;
wire wire3185;
wire wire3187;
wire wire3188;
wire wire3189;
wire wire3191;
wire wire3192;
wire wire3193;
wire wire3195;
wire wire3196;
wire wire3197;
wire wire3199;
wire wire3205;
wire wire3207;
wire wire3211;
wire wire3212;
wire wire3213;
wire wire3214;
wire wire3215;
wire wire3216;
wire wire3217;
wire wire3218;
wire wire3219;
wire wire3220;
wire wire3221;
wire wire3223;
wire wire3224;
wire wire3227;
wire wire3228;
wire wire3231;
wire wire3233;
wire wire3235;
wire wire3239;
wire wire3243;
wire wire3245;
wire wire3247;
wire wire3248;
wire wire3251;
wire wire3253;
wire wire3254;
wire wire3255;
wire wire3256;
wire wire3257;
wire wire3258;
wire wire3259;
wire wire3260;
wire wire3261;
wire wire3263;
wire wire3267;
wire wire3268;
wire wire3269;
wire wire3270;
wire wire3271;
wire wire3272;
wire wire3277;
wire wire3278;
wire wire3279;
wire wire3280;
wire wire3281;
wire wire3282;
wire wire3283;
wire wire3284;
wire wire3289;
wire wire3290;
wire wire3291;
wire wire3292;
wire wire3293;
wire wire3295;
wire wire3299;
wire wire3300;
wire wire3303;
wire wire3307;
wire wire3308;
wire wire3309;
wire wire3310;
wire wire3313;
wire wire3314;
wire wire3315;
wire wire3317;
wire wire3318;
wire wire3319;
wire wire3321;
wire wire3322;
wire wire3325;
wire wire3326;
wire wire3327;
wire wire3328;
wire wire3331;
wire wire3332;
wire wire3335;
wire wire3336;
wire wire3337;
wire wire3342;
wire wire3343;
wire wire3346;
wire wire3348;
wire wire3349;
wire wire3350;
wire wire3351;
wire wire3352;
wire wire3353;
wire wire3356;
wire wire3357;
wire wire3360;
wire wire3362;
wire wire3364;
wire wire3365;
wire wire3366;
wire wire3367;
wire wire3370;
wire wire3371;
wire wire3374;
wire wire3376;
wire wire3377;
wire wire3378;
wire wire3379;
wire wire3380;
wire wire3382;
wire wire3383;
wire wire3384;
wire wire3386;
wire wire3387;
wire wire3388;
wire wire3389;
wire wire3390;
wire wire3391;
wire wire3401;
wire wire3402;
wire wire3406;
wire wire3407;
wire wire3410;
wire wire3411;
wire wire3414;
wire wire3415;
wire wire3416;
wire wire3422;
wire wire3423;
wire wire3424;
wire wire3425;
wire wire3428;
wire wire3429;
wire wire3432;
wire wire3446;
wire wire3447;
wire wire3448;
wire wire3449;
wire wire3450;
wire wire3451;
wire wire3452;
wire wire3453;
wire wire3456;
wire wire3457;
wire wire3458;
wire wire3462;
wire wire3466;
wire wire3468;
wire wire3474;
wire wire3476;
wire wire3480;
wire wire3481;
wire wire3482;
wire wire3484;
wire wire3489;
wire wire3490;
wire wire3495;
wire wire3496;
wire wire3497;
wire wire3501;
wire wire3502;
wire wire3505;
wire wire3506;
wire wire3507;
wire wire3515;
wire wire3516;
wire wire3517;
wire wire3519;
wire wire3521;
wire wire3522;
wire wire3525;
wire wire3527;
wire wire3529;
wire wire3531;
wire wire3532;
wire wire3535;
wire wire3536;
wire wire3537;
wire wire3541;
wire wire3542;
wire wire3545;
wire wire3547;
wire wire3549;
wire wire3550;
wire wire3551;
wire wire3552;
wire wire3553;
wire wire3554;
wire wire3557;
wire wire3565;
wire wire3566;
wire wire3567;
wire wire3568;
wire wire3571;
wire wire3572;
wire wire3573;
wire wire3575;
wire wire3576;
wire wire3581;
wire wire3582;
wire wire3586;
wire wire3587;
wire wire3588;
wire wire3589;
wire wire3590;
wire wire3591;
wire wire3594;
wire wire3595;
wire wire3600;
wire wire3601;
wire wire3602;
wire wire3604;
wire wire3606;
wire wire3607;
wire wire3610;
wire wire3611;
wire wire3614;
wire wire3615;
wire wire3618;
wire wire3620;
wire wire3621;
wire wire3622;
wire wire3623;
wire wire3624;
wire wire3625;
wire wire3630;
wire wire3632;
wire wire3633;
wire wire3636;
wire wire3638;
wire wire3640;
wire wire3644;
wire wire3646;
wire wire3648;
wire wire3649;
wire wire3654;
wire wire3656;
wire wire3668;
wire wire3670;
wire wire3671;
wire wire3672;
wire wire3676;
wire wire3677;
wire wire3678;
wire wire3679;
wire wire3684;
wire wire3685;
wire wire3686;
wire wire3687;
wire wire3690;
wire wire3691;
wire wire3692;
wire wire3694;
wire wire3695;
wire wire3696;
wire wire3697;
wire wire3700;
wire wire3701;
wire wire3702;
wire wire3704;
wire wire3705;
wire wire3713;
wire wire3714;
wire wire3715;
wire wire3719;
wire wire3721;
wire wire3722;
wire wire3723;
wire wire3725;
wire wire3726;
wire wire3731;
wire wire3732;
wire wire3733;
wire wire3734;
wire wire3737;
wire wire3738;
wire wire3741;
wire wire3743;
wire wire3744;
wire wire3745;
wire wire3749;
wire wire3757;
wire wire3761;
wire wire3762;
wire wire3765;
wire wire3766;
wire wire3769;
wire wire3773;
wire wire3775;
wire wire3783;
wire wire3787;
wire wire3791;
wire wire3792;
wire wire3797;
wire wire3799;
wire wire3800;
wire wire3801;
wire wire3802;
wire wire3805;
wire wire3807;
wire wire3808;
wire wire3809;
wire wire3810;
wire wire3811;
wire wire3812;
wire wire3817;
wire wire3818;
wire wire3819;
wire wire3821;
wire wire3822;
wire wire3823;
wire wire3824;
wire wire3825;
wire wire3827;
wire wire3829;
wire wire3830;
wire wire3833;
wire wire3837;
wire wire3838;
wire wire3839;
wire wire3843;
wire wire3844;
wire wire3847;
wire wire3848;
wire wire3849;
wire wire3850;
wire wire3851;
wire wire3853;
wire wire3854;
wire wire3857;
wire wire3858;
wire wire3859;
wire wire3860;
wire wire3861;
wire wire3863;
wire wire3864;
wire wire3865;
wire wire3866;
wire wire3875;
wire wire3876;
wire wire3877;
wire wire3879;
wire wire3886;
wire wire3887;
wire wire3888;
wire wire3889;
wire wire3892;
wire wire3893;
wire wire3894;
wire wire3896;
wire wire3897;
wire wire3902;
wire wire3903;
wire wire3904;
wire wire3906;
wire wire3908;
wire wire3909;
wire wire3910;
wire wire3911;
wire wire3914;
wire wire3918;
wire wire3919;
wire wire3920;
wire wire3921;
wire wire3928;
wire wire3930;
wire wire3931;
wire wire3932;
wire wire3936;
wire wire3938;
wire wire3940;
wire wire3941;
wire wire3942;
wire wire3943;
wire wire3944;
wire wire3949;
wire wire3951;
wire wire3952;
wire wire3953;
wire wire3954;
wire wire3964;
wire wire3966;
wire wire3968;
wire wire3969;
wire wire3972;
wire wire3973;
wire wire3975;
wire wire3976;
wire wire3977;
wire wire3978;
wire wire3981;
wire wire3982;
wire wire3983;
wire wire3989;
wire wire3991;
wire wire3993;
wire wire3994;
wire wire3995;
wire wire3997;
wire wire3998;
wire wire4001;
wire wire4002;
wire wire4003;
wire wire4004;
wire wire4007;
wire wire4008;
wire wire4009;
wire wire4013;
wire wire4015;
wire wire4017;
wire wire4019;
wire wire4020;
wire wire4021;
wire wire4022;
wire wire4027;
wire wire4028;
wire wire4029;
wire wire4030;
wire wire4033;
wire wire4037;
wire wire4041;
wire wire4042;
wire wire4045;
wire wire4047;
wire wire4048;
wire wire4051;
wire wire4053;
wire wire4054;
wire wire4059;
wire wire4071;
wire wire4073;
wire wire4075;
wire wire4077;
wire wire4081;
wire wire4083;
wire wire4084;
wire wire4085;
wire wire4086;
wire wire4087;
wire wire4088;
wire wire4091;
wire wire4092;
wire wire4093;
wire wire4094;
wire wire4099;
wire wire4100;
wire wire4101;
wire wire4102;
wire wire4103;
wire wire4104;
wire wire4105;
wire wire4106;
wire wire4107;
wire wire4108;
wire wire4113;
wire wire4114;
wire wire4117;
wire wire4118;
wire wire4123;
wire wire4124;
wire wire4125;
wire wire4129;
wire wire4133;
wire wire4135;
wire wire4139;
wire wire4141;
wire wire4142;
wire wire4143;
wire wire4144;
wire wire4147;
wire wire4149;
wire wire4151;
wire wire4152;
wire wire4155;
wire wire4157;
wire wire4158;
wire wire4159;
wire wire4161;
wire wire4163;
wire wire4164;
wire wire4171;
wire wire4172;
wire wire4173;
wire wire4174;
wire wire4175;
wire wire4177;
wire wire4179;
wire wire4181;
wire wire4183;
wire wire4185;
wire wire4187;
wire wire4189;
wire wire4190;
wire wire4191;
wire wire4192;
wire wire4193;
wire wire4194;
wire wire4197;
wire wire4199;
wire wire4201;
wire wire4202;
wire wire4205;
wire wire4207;
wire wire4208;
wire wire4211;
wire wire4213;
wire wire4214;
wire wire4215;
wire wire4220;
wire wire4221;
wire wire4222;
wire wire4224;
wire wire4226;
wire wire4228;
wire wire4230;
wire wire4232;
wire wire4233;
wire wire4234;
wire wire4235;
wire wire4238;
wire wire4240;
wire wire4241;
wire wire4242;
wire wire4243;
wire wire4246;
wire wire4248;
wire wire4249;
wire wire4250;
wire wire4251;
wire wire4254;
wire wire4255;
wire wire4256;
wire wire4257;
wire wire4258;
wire wire4260;
wire wire4261;
wire wire4264;
wire wire4265;
wire wire4272;
wire wire4273;
wire wire4274;
wire wire4275;
wire wire4278;
wire wire4280;
wire wire4281;
wire wire4282;
wire wire4283;
wire wire4288;
wire wire4289;
wire wire4290;
wire wire4291;
wire wire4292;
wire wire4294;
wire wire4295;
wire wire4296;
wire wire4297;
wire wire4302;
wire wire4304;
wire wire4310;
wire wire4311;
wire wire4314;
wire wire4316;
wire wire4317;
wire wire4318;
wire wire4319;
wire wire4320;
wire wire4322;
wire wire4323;
wire wire4326;
wire wire4327;
wire wire4328;
wire wire4329;
wire wire4330;
wire wire4331;
wire wire4344;
wire wire4346;
wire wire4350;
wire wire4352;
wire wire4354;
wire wire4355;
wire wire4358;
wire wire4360;
wire wire4361;
wire wire4364;
wire wire4365;
wire wire4370;
wire wire4372;
wire wire4374;
wire wire4376;
wire wire4378;
wire wire4380;
wire wire4382;
wire wire4384;
wire wire4385;
wire wire4386;
wire wire4388;
wire wire4389;
wire wire4390;
wire wire4392;
wire wire4394;
wire wire4396;
wire wire4397;
wire wire4398;
wire wire4400;
wire wire4401;
wire wire4404;
wire wire4406;
wire wire4407;
wire wire4411;
wire wire4412;
wire wire4416;
wire wire4417;
wire wire4421;
wire wire4424;
wire wire4425;
wire wire4428;
wire wire4429;
wire wire4432;
wire wire4433;
wire wire4434;
wire wire4436;
wire wire4437;
wire wire4440;
wire wire4444;
wire wire4445;
wire wire4448;
wire wire4450;
wire wire4452;
wire wire4456;
wire wire4460;
wire wire4462;
wire wire4463;
wire wire4464;
wire wire4468;
wire wire4469;
wire wire4472;
wire wire4473;
wire wire4474;
wire wire4475;
wire wire4480;
wire wire4481;
wire wire4488;
wire wire4489;
wire wire4490;
wire wire4491;
wire wire4494;
wire wire4496;
wire wire4497;
wire wire4498;
wire wire4499;
wire wire4502;
wire wire4504;
wire wire4505;
wire wire4508;
wire wire4509;
wire wire4510;
wire wire4518;
wire wire4519;
wire wire4520;
wire wire4521;
wire wire4522;
wire wire4523;
wire wire4526;
wire wire4527;
wire wire4530;
wire wire4531;
wire wire4532;
wire wire4533;
wire wire4534;
wire wire4535;
wire wire4536;
wire wire4538;
wire wire4544;
wire wire4545;
wire wire4546;
wire wire4548;
wire wire4549;
wire wire4582;
wire wire4588;
wire wire4590;
wire wire4591;
wire wire4592;
wire wire4594;
wire wire4598;
wire wire4600;
wire wire4602;
wire wire4603;
wire wire4606;
wire wire4614;
wire wire4618;
wire wire4619;
wire wire4620;
wire wire4621;
wire wire4624;
wire wire4625;
wire wire4628;
wire wire4630;
wire wire4631;
wire wire4634;
wire wire4635;
wire wire4636;
wire wire4637;
wire wire4640;
wire wire4641;
wire wire4644;
wire wire4646;
wire wire4648;
wire wire4649;
wire wire4650;
wire wire4651;
wire wire4652;
wire wire4653;
wire wire4654;
wire wire4655;
wire wire4660;
wire wire4662;
wire wire4664;
wire wire4665;
wire wire4666;
wire wire4668;
wire wire4672;
wire wire4673;
wire wire4678;
wire wire4679;
wire wire4684;
wire wire4685;
wire wire4686;
wire wire4687;
wire wire4688;
wire wire4689;
wire wire4690;
wire wire4691;
wire wire4692;
wire wire4693;
wire wire4694;
wire wire4695;
wire wire4696;
wire wire4697;
wire wire4701;
wire wire4702;
wire wire4703;
wire wire4704;
wire wire4705;
wire wire4706;
wire wire4707;
wire wire4708;
wire wire4709;
wire wire4710;
wire wire4711;
wire wire4712;
wire wire4713;
wire wire4714;
wire wire4717;
wire wire4718;
wire wire4723;
wire wire4724;
wire wire4725;
wire wire4726;
wire wire4727;
wire wire4728;
wire wire4729;
wire wire4730;
wire wire4731;
wire wire4732;
wire wire4733;
wire wire4734;
wire wire4735;
wire wire4736;
wire wire4740;
wire wire4741;
wire wire4742;
wire wire4743;
wire wire4744;
wire wire4745;
wire wire4746;
wire wire4747;
wire wire4748;
wire wire4749;
wire wire4750;
wire wire4751;
wire wire4752;
wire wire4753;
wire wire4760;
wire wire4761;
wire wire4768;
wire wire4769;
wire wire4773;
wire wire4774;
wire wire4775;
wire wire4776;
wire wire4777;
wire wire4778;
wire wire4779;
wire wire4780;
wire wire4781;
wire wire4782;
wire wire4783;
wire wire4784;
wire wire4785;
wire wire4786;
wire wire4787;
wire wire4788;
wire wire4793;
wire wire4794;
wire wire4795;
wire wire4796;
wire wire4797;
wire wire4798;
wire wire4799;
wire wire4800;
wire wire4801;
wire wire4802;
wire wire4803;
wire wire4804;
wire wire4805;
wire wire4809;
wire wire4810;
wire wire4811;
wire wire4812;
wire wire4817;
wire wire4818;
wire wire4819;
wire wire4821;
wire wire4823;
wire wire4827;
wire wire4828;
wire wire4833;
wire wire4843;
wire wire4844;
wire wire4847;
wire wire4848;
wire wire4851;
wire wire4852;
wire wire4857;
wire wire4861;
wire wire4864;
wire wire4865;
wire wire4866;
wire wire4867;
wire wire4868;
wire wire4869;
wire wire4870;
wire wire4877;
wire wire4878;
wire wire4879;
wire wire4880;
wire wire4881;
wire wire4882;
wire wire4883;
wire wire4886;
wire wire4887;
wire wire4888;
wire wire4889;
wire wire4890;
wire wire4891;
wire wire4892;
wire wire4899;
wire wire4900;
wire wire4901;
wire wire4902;
wire wire4903;
wire wire4904;
wire wire4905;
wire wire4918;
wire wire4919;
wire wire4920;
wire wire4921;
wire wire4922;
wire wire4923;
wire wire4924;
wire wire4927;
wire wire4928;
wire wire4929;
wire wire4930;
wire wire4931;
wire wire4932;
wire wire4933;
wire wire4934;
wire wire4935;
wire wire4936;
wire wire4937;
wire wire4938;
wire wire4939;
wire wire4940;
wire wire4941;
wire wire4942;
wire wire4943;
wire wire4944;
wire wire4945;
wire wire4946;
wire wire4947;
wire wire4948;
wire wire4949;
wire wire4950;
wire wire4951;
wire wire4952;
wire wire4953;
wire wire4954;
wire wire4955;
wire wire4956;
wire wire4957;
wire wire4958;
wire wire4959;
wire wire4960;
wire wire4961;
wire wire4962;
wire wire4963;
wire wire4964;
wire wire4965;
wire wire4966;
wire wire4967;
wire wire4968;
wire wire4969;
wire wire4970;
wire wire4971;
wire wire4972;
wire wire4973;
wire wire4974;
wire wire4975;
wire wire4976;
wire wire4977;
wire wire4978;
wire wire4979;
wire wire4980;
wire wire4981;
wire wire4982;
wire wire4983;
wire wire4984;
wire wire4985;
wire wire4986;
wire wire4987;
wire wire4988;
wire wire4989;
wire wire4990;
wire wire4991;
wire wire4992;
wire wire4993;
wire wire4994;
wire wire4995;
wire wire4996;
wire wire4997;
wire wire4998;
wire wire4999;
wire wire5000;
wire wire5001;
wire wire5002;
wire wire5003;
wire wire5004;
wire wire5005;
wire wire5006;
wire wire5007;
wire wire5008;
wire wire5009;
wire wire5010;
wire wire5012;
wire wire5013;
wire wire5022;
wire wire5026;
wire wire5027;
wire wire5032;
wire wire5033;
wire wire5037;
wire wire5038;
wire wire5039;
wire wire5040;
wire wire5041;
wire wire5042;
wire wire5043;
wire wire5044;
wire wire5045;
wire wire5046;
wire wire5047;
wire wire5048;
wire wire5049;
wire wire5050;
wire wire5051;
wire wire5052;
wire wire5057;
wire wire5058;
wire wire5059;
wire wire5060;
wire wire5061;
wire wire5062;
wire wire5063;
wire wire5064;
wire wire5065;
wire wire5066;
wire wire5067;
wire wire5068;
wire wire5069;
wire wire5070;
wire wire5071;
wire wire5072;
wire wire5077;
wire wire5083;
wire wire5084;
wire wire5088;
wire wire5089;
wire wire5090;
wire wire5091;
wire wire5092;
wire wire5093;
wire wire5094;
wire wire5095;
wire wire5096;
wire wire5097;
wire wire5098;
wire wire5099;
wire wire5100;
wire wire5101;
wire wire5102;
wire wire5103;
wire wire5108;
wire wire5109;
wire wire5110;
wire wire5111;
wire wire5112;
wire wire5113;
wire wire5114;
wire wire5115;
wire wire5116;
wire wire5117;
wire wire5118;
wire wire5119;
wire wire5124;
wire wire5125;
wire wire5130;
wire wire5131;
wire wire5132;
wire wire5133;
wire wire5134;
wire wire5135;
wire wire5136;
wire wire5137;
wire wire5138;
wire wire5139;
wire wire5140;
wire wire5141;
wire wire5142;
wire wire5143;
wire wire5147;
wire wire5148;
wire wire5149;
wire wire5150;
wire wire5151;
wire wire5152;
wire wire5153;
wire wire5154;
wire wire5155;
wire wire5156;
wire wire5157;
wire wire5158;
wire wire5159;
wire wire5160;
wire wire5165;
wire wire5166;
wire wire5170;
wire wire5171;
wire wire5172;
wire wire5173;
wire wire5174;
wire wire5175;
wire wire5176;
wire wire5177;
wire wire5178;
wire wire5179;
wire wire5180;
wire wire5181;
wire wire5182;
wire wire5183;
wire wire5184;
wire wire5185;
wire wire5188;
wire wire5189;
wire wire5193;
wire wire5194;
wire wire5195;
wire wire5196;
wire wire5197;
wire wire5198;
wire wire5199;
wire wire5200;
wire wire5201;
wire wire5202;
wire wire5203;
wire wire5204;
wire wire5205;
wire wire5206;
wire wire5209;
wire wire5210;
wire wire5215;
wire wire5216;
wire wire5217;
wire wire5218;
wire wire5219;
wire wire5220;
wire wire5221;
wire wire5222;
wire wire5223;
wire wire5224;
wire wire5225;
wire wire5226;
wire wire5227;
wire wire5228;
wire wire5233;
wire wire5234;
wire wire5235;
wire wire5236;
wire wire5237;
wire wire5238;
wire wire5239;
wire wire5240;
wire wire5241;
wire wire5242;
wire wire5243;
wire wire5244;
wire wire5245;
wire wire5246;
wire wire5251;
wire wire5252;
wire wire5256;
wire wire5257;
wire wire5258;
wire wire5259;
wire wire5260;
wire wire5261;
wire wire5262;
wire wire5263;
wire wire5264;
wire wire5265;
wire wire5266;
wire wire5267;
wire wire5268;
wire wire5269;
wire wire5270;
wire wire5271;
wire wire5276;
wire wire5277;
wire wire5278;
wire wire5279;
wire wire5280;
wire wire5281;
wire wire5282;
wire wire5283;
wire wire5284;
wire wire5285;
wire wire5286;
wire wire5287;
wire wire5292;
wire wire5293;
wire wire5297;
wire wire5298;
wire wire5299;
wire wire5300;
wire wire5301;
wire wire5302;
wire wire5303;
wire wire5304;
wire wire5305;
wire wire5306;
wire wire5307;
wire wire5308;
wire wire5309;
wire wire5310;
wire wire5311;
wire wire5312;
wire wire5319;
wire wire5320;
wire wire5324;
wire wire5325;
wire wire5326;
wire wire5327;
wire wire5328;
wire wire5329;
wire wire5330;
wire wire5331;
wire wire5332;
wire wire5333;
wire wire5334;
wire wire5335;
wire wire5336;
wire wire5337;
wire wire5338;
wire wire5339;
wire wire5342;
wire wire5343;
wire wire5347;
wire wire5348;
wire wire5349;
wire wire5350;
wire wire5351;
wire wire5352;
wire wire5353;
wire wire5354;
wire wire5355;
wire wire5356;
wire wire5357;
wire wire5358;
wire wire5359;
wire wire5360;
wire wire5363;
wire wire5364;
wire wire5368;
wire wire5369;
wire wire5370;
wire wire5371;
wire wire5372;
wire wire5373;
wire wire5374;
wire wire5375;
wire wire5376;
wire wire5377;
wire wire5378;
wire wire5379;
wire wire5380;
wire wire5381;
wire wire5382;
wire wire5383;
wire wire5388;
wire wire5389;
wire wire5390;
wire wire5391;
wire wire5392;
wire wire5393;
wire wire5394;
wire wire5395;
wire wire5396;
wire wire5397;
wire wire5398;
wire wire5399;
wire wire5402;
wire wire5403;
wire wire5408;
wire wire5409;
wire wire5410;
wire wire5411;
wire wire5412;
wire wire5413;
wire wire5414;
wire wire5415;
wire wire5416;
wire wire5417;
wire wire5418;
wire wire5419;
wire wire5420;
wire wire5421;
wire wire5425;
wire wire5426;
wire wire5427;
wire wire5428;
wire wire5429;
wire wire5430;
wire wire5431;
wire wire5432;
wire wire5433;
wire wire5434;
wire wire5435;
wire wire5436;
wire wire5437;
wire wire5438;
wire wire5439;
wire wire5440;
wire wire5445;
wire wire5446;
wire wire5447;
wire wire5448;
wire wire5449;
wire wire5450;
wire wire5451;
wire wire5452;
wire wire5453;
wire wire5454;
wire wire5455;
wire wire5456;
wire wire5457;
wire wire5458;
wire wire5463;
wire wire5464;
wire wire5465;
wire wire5466;
wire wire5467;
wire wire5468;
wire wire5469;
wire wire5470;
wire wire5471;
wire wire5472;
wire wire5473;
wire wire5474;
wire wire5477;
wire wire5478;
wire wire5483;
wire wire5484;
wire wire5485;
wire wire5486;
wire wire5487;
wire wire5488;
wire wire5489;
wire wire5490;
wire wire5491;
wire wire5492;
wire wire5493;
wire wire5494;
wire wire5495;
wire wire5496;
wire wire5500;
wire wire5501;
wire wire5502;
wire wire5503;
wire wire5504;
wire wire5505;
wire wire5506;
wire wire5507;
wire wire5508;
wire wire5509;
wire wire5510;
wire wire5511;
wire wire5512;
wire wire5513;
wire wire5516;
wire wire5517;
wire wire5521;
wire wire5522;
wire wire5523;
wire wire5524;
wire wire5525;
wire wire5526;
wire wire5527;
wire wire5528;
wire wire5529;
wire wire5530;
wire wire5531;
wire wire5532;
wire wire5533;
wire wire5534;
wire wire5535;
wire wire5536;
wire wire5541;
wire wire5542;
wire wire5543;
wire wire5544;
wire wire5545;
wire wire5546;
wire wire5547;
wire wire5548;
wire wire5549;
wire wire5550;
wire wire5551;
wire wire5552;
wire wire5553;
wire wire5554;
wire wire5559;
wire wire5560;
wire wire5561;
wire wire5562;
wire wire5563;
wire wire5564;
wire wire5565;
wire wire5566;
wire wire5567;
wire wire5568;
wire wire5569;
wire wire5570;
wire wire5571;
wire wire5572;
wire wire5573;
wire wire5575;
wire wire5579;
wire wire5580;
wire wire5581;
wire wire5582;
wire wire5583;
wire wire5584;
wire wire5585;
wire wire5586;
wire wire5587;
wire wire5588;
wire wire5589;
wire wire5590;
wire wire5591;
wire wire5592;
wire wire5593;
wire wire5594;
wire wire5595;
wire wire5596;
wire wire5597;
wire wire5598;
wire wire5599;
wire wire5600;
wire wire5601;
wire wire5602;
wire wire5603;
wire wire5604;
wire wire5605;
wire wire5606;
wire wire5607;
wire wire5608;
wire wire5609;
wire wire5610;
wire wire5611;
wire wire5612;
wire wire5613;
wire wire5614;
wire wire5615;
wire wire5616;
wire wire5617;
wire wire5618;
wire wire5619;
wire wire5620;
wire wire5621;
wire wire5622;
wire wire5623;
wire wire5624;
wire wire5625;
wire wire5626;
wire wire5627;
wire wire5628;
wire wire5629;
wire wire5630;
wire wire5631;
wire wire5632;
wire wire5633;
wire wire5634;
wire wire5635;
wire wire5636;
wire wire5637;
wire wire5638;
wire wire5639;
wire wire5640;
wire wire5641;
wire wire5642;
wire wire5643;
wire wire5644;
wire wire5645;
wire wire5646;
wire wire5647;
wire wire5648;
wire wire5649;
wire wire5650;
wire wire5651;
wire wire5652;
wire wire5653;
wire wire5654;
wire wire5655;
wire wire5656;
wire wire5657;
wire wire5658;
wire wire5659;
wire wire5660;
wire wire5661;
wire wire5662;
wire wire5663;
wire wire5664;
wire wire5665;
wire wire5666;
wire wire5667;
wire wire5668;
wire wire5669;
wire wire5670;
wire wire5671;
wire wire5672;
wire wire5673;
wire wire5674;
wire wire5675;
wire wire5676;
wire wire5677;
wire wire5678;
wire wire5679;
wire wire5680;
wire wire5681;
wire wire5682;
wire wire5683;
wire wire5684;
wire wire5685;
wire wire5686;
wire wire5687;
wire wire5688;
wire wire5689;
wire wire5690;
wire wire5691;
wire wire5692;
wire wire5693;
wire wire5694;
wire wire5695;
wire wire5696;
wire wire5697;
wire wire5698;
wire wire5699;
wire wire5700;
wire wire5701;
wire wire5702;
wire wire5703;
wire wire5704;
wire wire5705;
wire wire5706;
wire wire15923;
wire wire15924;
wire wire15929;
wire wire15930;
wire wire15935;
wire wire15936;
wire wire15941;
wire wire15942;
wire wire15947;
wire wire15948;
wire wire15953;
wire wire15954;
wire wire15959;
wire wire15960;
wire wire15965;
wire wire15966;
wire wire15971;
wire wire15972;
wire wire15977;
wire wire15978;
wire wire15983;
wire wire15984;
wire wire15989;
wire wire15990;
wire wire15995;
wire wire15996;
wire wire16001;
wire wire16002;
wire wire16007;
wire wire16008;
wire wire16013;
wire wire16014;
wire wire16015;
wire wire16016;
wire wire16017;
wire wire16018;
wire wire16019;
wire wire16020;
wire wire16021;
wire wire16022;
wire wire16027;
wire wire16028;
wire wire16029;
wire wire16030;
wire wire16037;
wire wire16038;
wire wire16039;
wire wire16040;
wire wire16041;
wire wire16045;
wire wire16046;
wire wire16047;
wire wire16048;
wire wire16056;
wire wire16057;
wire wire16058;
wire wire16059;
wire wire16060;
wire wire16064;
wire wire16065;
wire wire16073;
wire wire16074;
wire wire16075;
wire wire16076;
wire wire16077;
wire wire16081;
wire wire16082;
wire wire16089;
wire wire16090;
wire wire16091;
wire wire16092;
wire wire16093;
wire wire16097;
wire wire16098;
wire wire16106;
wire wire16107;
wire wire16108;
wire wire16109;
wire wire16110;
wire wire16114;
wire wire16115;
wire wire16122;
wire wire16123;
wire wire16124;
wire wire16125;
wire wire16126;
wire wire16130;
wire wire16131;
wire wire16138;
wire wire16139;
wire wire16140;
wire wire16141;
wire wire16142;
wire wire16146;
wire wire16147;
wire wire16155;
wire wire16156;
wire wire16157;
wire wire16158;
wire wire16159;
wire wire16163;
wire wire16164;
wire wire16171;
wire wire16172;
wire wire16173;
wire wire16174;
wire wire16175;
wire wire16179;
wire wire16180;
wire wire16188;
wire wire16189;
wire wire16190;
wire wire16191;
wire wire16192;
wire wire16196;
wire wire16197;
wire wire16204;
wire wire16205;
wire wire16206;
wire wire16207;
wire wire16208;
wire wire16212;
wire wire16213;
wire wire16221;
wire wire16222;
wire wire16223;
wire wire16224;
wire wire16225;
wire wire16229;
wire wire16230;
wire wire16237;
wire wire16238;
wire wire16239;
wire wire16240;
wire wire16241;
wire wire16245;
wire wire16246;
wire wire16254;
wire wire16255;
wire wire16256;
wire wire16257;
wire wire16258;
wire wire16262;
wire wire16263;
wire wire16270;
wire wire16271;
wire wire16272;
wire wire16273;
wire wire16274;
wire wire16278;
wire wire16279;
wire wire16287;
wire wire16288;
wire wire16289;
wire wire16290;
wire wire16291;
wire wire16295;
wire wire16296;
wire wire16303;
wire wire16304;
wire wire16305;
wire wire16306;
wire wire16307;
wire wire16311;
wire wire16312;
wire wire16320;
wire wire16321;
wire wire16322;
wire wire16323;
wire wire16324;
wire wire16328;
wire wire16329;
wire wire16336;
wire wire16337;
wire wire16338;
wire wire16339;
wire wire16340;
wire wire16344;
wire wire16345;
wire wire16353;
wire wire16354;
wire wire16355;
wire wire16356;
wire wire16357;
wire wire16361;
wire wire16362;
wire wire16369;
wire wire16370;
wire wire16371;
wire wire16372;
wire wire16373;
wire wire16377;
wire wire16378;
wire wire16386;
wire wire16387;
wire wire16388;
wire wire16389;
wire wire16390;
wire wire16394;
wire wire16395;
wire wire16402;
wire wire16403;
wire wire16404;
wire wire16405;
wire wire16406;
wire wire16410;
wire wire16411;
wire wire16419;
wire wire16420;
wire wire16421;
wire wire16422;
wire wire16423;
wire wire16427;
wire wire16428;
wire wire16437;
wire wire16438;
wire wire16439;
wire wire16440;
wire wire16441;
wire wire16445;
wire wire16446;
wire wire16453;
wire wire16454;
wire wire16455;
wire wire16456;
wire wire16457;
wire wire16461;
wire wire16462;
wire wire16463;
wire wire16464;
wire wire16465;
wire wire16466;
wire wire16469;
wire wire16473;
wire wire16474;
wire wire16478;
wire wire16479;
wire wire16483;
wire wire16484;
wire wire16488;
wire wire16489;
wire wire16493;
wire wire16494;
wire wire16498;
wire wire16499;
wire wire16503;
wire wire16504;
wire wire16508;
wire wire16509;
wire wire16513;
wire wire16514;
wire wire16518;
wire wire16519;
wire wire16523;
wire wire16524;
wire wire16528;
wire wire16529;
wire wire16533;
wire wire16534;
wire wire16538;
wire wire16539;
wire wire16543;
wire wire16544;
wire wire16549;
wire wire16550;
wire wire16551;
wire wire16554;
wire wire16565;
wire wire16566;
wire wire16567;
wire wire16568;
wire wire16569;
wire wire16573;
wire wire16574;
wire wire16582;
wire wire16583;
wire wire16584;
wire wire16585;
wire wire16586;
wire wire16590;
wire wire16591;
wire wire16599;
wire wire16600;
wire wire16601;
wire wire16602;
wire wire16603;
wire wire16607;
wire wire16608;
wire wire16615;
wire wire16616;
wire wire16617;
wire wire16618;
wire wire16619;
wire wire16623;
wire wire16624;
wire wire16631;
wire wire16632;
wire wire16633;
wire wire16634;
wire wire16635;
wire wire16639;
wire wire16640;
wire wire16648;
wire wire16649;
wire wire16650;
wire wire16651;
wire wire16652;
wire wire16656;
wire wire16657;
wire wire16661;
wire wire16662;
wire wire16663;
wire wire16664;
wire wire16667;
wire wire16668;
wire wire16670;
wire wire16671;
wire wire16674;
wire wire16676;
wire wire16682;
wire wire16686;
wire wire16687;
wire wire16688;
wire wire16690;
wire wire16698;
wire wire16701;
wire wire16703;
wire wire16704;
wire wire16705;
wire wire16707;
wire wire16714;
wire wire16715;
wire wire16716;
wire wire16717;
wire wire16719;
wire wire16721;
wire wire16726;
wire wire16727;
wire wire16728;
wire wire16729;
wire wire16732;
wire wire16734;
wire wire16742;
wire wire16748;
wire wire16754;
wire wire16759;
wire wire16760;
wire wire16763;
wire wire16765;
wire wire16766;
wire wire16768;
wire wire16775;
wire wire16777;
wire wire16782;
wire wire16786;
wire wire16790;
reg n_n9280;

reg n_n9172;

reg n_n9260;

reg n_n7726;

reg n_n8270;

reg n_n8196;

reg n_n9150;

reg n_n9267;

reg n_n7779;

reg n_n9503;

reg n_n8150;

reg n_n9401;

reg n_n7341;

reg n_n9180;

reg n_n8592;

reg n_n8871;

reg n_n7252;

reg n_n7271;

reg n_n6991;

reg n_n8557;

reg n_n7707;

reg n_n7552;

reg ndn3_23;

reg n_n9548;

reg n_n9467;

reg n_n8002;

reg n_n6950;

reg n_n8930;

reg n_n7244;

reg n_n7819;

reg n_n8883;

reg n_n7709;

reg n_n9580;

reg n_n9130;

reg n_n9486;

reg n_n9235;

reg n_n7522;

reg n_n7373;

reg n_n9085;

reg n_n9638;

reg n_n7452;

reg n_n8775;

reg n_n7654;

reg n_n8410;

reg n_n8208;

reg n_n8377;

reg n_n7558;

reg n_n7599;

reg n_n8225;

reg n_n8202;

reg n_n7670;

reg n_n7888;

reg n_n7889;

reg n_n8597;

reg n_n8152;

reg n_n8394;

reg n_n7812;

reg n_n7816;

reg n_n9141;

reg n_n7332;

reg n_n8758;

reg n_n7765;

reg n_n7877;

reg n_n7814;

reg n_n9008;

reg n_n7581;

reg n_n7376;

reg n_n7970;

reg pover_0_0_;

reg n_n8599;

reg n_n8227;

reg n_n9442;

reg n_n9485;

reg n_n7148;

reg n_n9311;

reg n_n9273;

reg ndn3_9;

reg n_n8613;

reg n_n8533;

reg n_n8699;

reg n_n8609;

reg n_n8308;

reg n_n8655;

reg n_n8981;

reg n_n7583;

reg n_n9198;

reg n_n9602;

reg n_n8786;

reg n_n9598;

reg n_n7738;

reg n_n8573;

reg n_n9473;

reg n_n9000;

reg n_n8001;

reg n_n9554;

reg n_n8508;

reg n_n9635;

reg n_n7190;

reg n_n8702;

reg n_n9106;

reg n_n7409;

reg n_n9437;

reg n_n9052;

reg n_n8647;

reg n_n9265;

reg n_n7179;

reg ndn3_13;

reg ndn3_17;

reg ndn3_25;

reg ndn3_29;

reg n_n9539;

reg n_n7953;

reg n_n8488;

reg nen3_22;

reg n_n9438;

reg n_n8132;

reg n_n8661;

reg n_n7759;

reg n_n8333;

reg n_n9399;

reg n_n7798;

reg n_n9434;

reg n_n7910;

reg n_n9528;

reg n_n7850;

reg n_n8251;

reg n_n7937;

reg n_n8482;

reg n_n9290;

reg n_n8007;

reg n_n7556;

reg n_n9064;

reg n_n9398;

reg n_n9412;

reg n_n9361;

reg n_n9304;

reg n_n7651;

reg n_n7712;

reg n_n7735;

reg n_n7934;

reg n_n7811;

reg n_n8053;

reg n_n9015;

reg n_n8066;

reg n_n9518;

reg n_n8091;

reg n_n9257;

reg n_n8175;

reg n_n8491;

reg n_n8114;

reg n_n7951;

reg n_n8913;

reg n_n8035;

reg n_n8631;

reg n_n8243;

reg n_n7857;

reg ngfdn_3;

reg n_n7791;

reg n_n9175;

reg n_n9588;

reg n_n9049;

reg n_n9483;

reg n_n9410;

reg n_n7691;

reg n_n7740;

reg n_n7602;

reg n_n7783;

reg n_n7948;

reg n_n7054;

reg n_n9343;

reg n_n9400;

reg nsr1_2;

reg n_n9127;

reg n_n8531;

reg n_n9335;

reg n_n7324;

reg n_n9611;

reg n_n8112;

reg n_n9406;

reg n_n9618;

reg n_n9613;

reg n_n9242;

reg n_n7384;

reg n_n8884;

reg n_n7462;

reg n_n7908;

reg n_n8765;

reg n_n7909;

reg n_n7898;

reg n_n9135;

reg n_n8862;

reg n_n8037;

reg ndn3_18;

reg ndn3_22;

reg n_n8974;

reg n_n7286;

reg n_n9223;

reg n_n7306;

reg n_n9169;

reg n_n9125;

reg nen3_39;

reg n_n8278;

reg n_n9557;

reg n_n7758;

reg n_n9391;

reg n_n8110;

reg n_n9597;

reg n_n8568;

reg n_n7428;

reg n_n7931;

reg n_n7742;

reg n_n7236;

reg n_n8219;

reg n_n9568;

reg n_n9200;

reg n_n8545;

reg n_n7823;

reg n_n8005;

reg n_n8736;

reg n_n9339;

reg n_n8499;

reg n_n8086;

reg n_n7803;

reg n_n7640;

reg n_n9098;

reg n_n7160;

reg n_n7713;

reg n_n9566;

reg n_n7955;

reg n_n8414;

reg n_n8006;

reg n_n9560;

reg n_n8742;

reg n_n7174;

reg n_n8882;

reg n_n7546;

reg n_n8282;

reg n_n8998;

reg n_n7656;

reg n_n9465;

reg n_n9601;

reg n_n8875;

reg n_n7954;

reg n_n8959;

reg n_n8957;

reg n_n8247;

reg n_n8258;

reg n_n7641;

reg n_n8843;

reg n_n9321;

reg n_n7702;

reg nsr3_23;

reg n_n8199;

reg n_n7983;

reg n_n7217;

reg n_n7821;

reg n_n9489;

reg n_n8348;

reg n_n9408;

reg n_n8445;

reg n_n9501;

reg n_n7831;

reg n_n7757;

reg n_n9174;

reg n_n9432;

reg n_n8678;

reg n_n8024;

reg n_n7806;

reg n_n8996;

reg n_n7918;

reg n_n8260;

reg n_n9341;

reg n_n9189;

reg n_n9096;

reg ndn3_30;

reg n_n7775;

reg n_n7693;

reg nen3_16;

reg n_n7643;

reg n_n8941;

reg n_n8042;

reg n_n8681;

reg n_n8659;

reg n_n9110;

reg n_n9573;

reg n_n8951;

reg n_n9589;

reg n_n9387;

reg n_n8279;

reg n_n7790;

reg n_n8406;

reg n_n8582;

reg n_n7911;

reg n_n7474;

reg n_n8466;

reg n_n6984;

reg n_n7760;

reg n_n7847;

reg n_n9559;

reg n_n7362;

reg n_n9300;

reg n_n9550;

reg n_n9492;

reg n_n8777;

reg n_n7764;

reg n_n7826;

reg n_n7777;

reg n_n7824;

reg n_n8173;

reg n_n7498;

reg n_n9148;

reg n_n8753;

reg n_n8772;

reg n_n8049;

reg n_n9362;

reg ndn1_4;

reg n_n9561;

reg n_n9004;

reg n_n8203;

reg n_n8153;

reg n_n9263;

reg n_n8369;

reg n_n9331;

reg n_n7454;

reg ndn3_7;

reg n_n7527;

reg n_n9036;

reg n_n7875;

reg n_n8697;

reg n_n9497;

reg n_n7291;

reg nsr3_13;

reg nsr3_38;

reg n_n8240;

reg n_n7703;

reg n_n9282;

reg n_n8237;

reg n_n8935;

reg n_n9244;

reg n_n8648;

reg n_n8235;

reg n_n8611;

reg n_n9045;

reg n_n9334;

reg n_n8572;

reg n_n9491;

reg n_n9134;

reg n_n9555;

reg n_n9336;

reg n_n7050;

reg n_n9346;

reg n_n7140;

reg n_n7681;

reg n_n6948;

reg n_n8549;

reg ndn3_19;

reg ndn3_28;

reg n_n7102;

reg n_n8093;

reg n_n9041;

reg n_n8381;

reg n_n8810;

reg nen3_36;

reg n_n9047;

reg n_n9333;

reg n_n7736;

reg n_n7820;

reg n_n8986;

reg n_n8891;

reg n_n8000;

reg n_n7968;

reg n_n8750;

reg n_n9558;

reg n_n9368;

reg n_n8519;

reg n_n6956;

reg n_n8298;

reg n_n9397;

reg n_n7017;

reg n_n8638;

reg n_n9552;

reg n_n8964;

reg n_n8016;

reg n_n7603;

reg n_n7696;

reg n_n8589;

reg n_n9337;

reg n_n9132;

reg n_n8652;

reg n_n8707;

reg n_n9407;

reg n_n9044;

reg n_n8808;

reg nsr3_30;

reg n_n8274;

reg n_n8615;

reg n_n8238;

reg n_n7854;

reg n_n8649;

reg n_n8236;

reg n_n8269;

reg n_n9592;

reg n_n8022;

reg n_n8744;

reg n_n8529;

reg n_n7967;

reg n_n9487;

reg n_n8685;

reg n_n9531;

reg n_n9510;

reg n_n7771;

reg n_n8480;

reg n_n8543;

reg n_n7789;

reg ndn3_11;

reg ndn3_15;

reg ndn3_21;

reg n_n7584;

reg n_n8354;

reg n_n6952;

reg n_n8864;

reg n_n7930;

reg n_n7962;

reg n_n7929;

reg n_n9316;

reg n_n9102;

reg n_n7308;

reg n_n7657;

reg n_n9264;

reg n_n8760;

reg n_n6912;

reg n_n7887;

reg n_n8911;

reg n_n7952;

reg n_n8704;

reg n_n7876;

reg n_n9596;

reg n_n8430;

reg n_n9019;

reg n_n7699;

reg n_n7375;

reg n_n7936;

reg n_n8340;

reg n_n8809;

reg n_n6961;

reg n_n9429;

reg n_n7743;

reg n_n8980;

reg n_n7582;

reg n_n8968;

reg n_n9371;

reg n_n8741;

reg n_n9502;

reg n_n9373;

reg n_n9248;

reg n_n7822;

reg n_n9054;

reg n_n8273;

reg n_n6937;

reg n_n9342;

reg n_n9325;

reg n_n9609;

reg n_n9623;

reg n_n9470;

reg n_n7570;

reg n_n9310;

reg n_n9366;

reg n_n7181;

reg n_n8739;

reg n_n8939;

reg n_n7256;

reg n_n8983;

reg n_n7487;

reg n_n9268;

reg n_n8906;

reg n_n7988;

reg n_n9181;

reg n_n8725;

reg n_n8626;

reg ndn3_27;

reg n_n8210;

reg n_n7415;

reg n_n8900;

reg nen3_19;

reg n_n8762;

reg n_n8512;

reg n_n8095;

reg n_n8982;

reg n_n7387;

reg n_n9494;

reg n_n7689;

reg n_n7835;

reg n_n9157;

reg n_n8552;

reg n_n7381;

reg n_n9446;

reg n_n8633;

reg n_n7684;

reg n_n7310;

reg n_n8402;

reg n_n9315;

reg n_n7950;

reg n_n8504;

reg n_n8456;

reg n_n7514;

reg n_n7315;

reg n_n9476;

reg n_n8276;

reg n_n8833;

reg n_n7923;

reg n_n9395;

reg n_n9512;

reg n_n9319;

reg nsr3_35;

reg n_n7154;

reg n_n9495;

reg n_n9137;

reg n_n8854;

reg n_n9183;

reg n_n9323;

reg n_n9349;

reg n_n7896;

reg n_n8073;

reg n_n8970;

reg n_n9314;

reg n_n8486;

reg n_n7246;

reg n_n7866;

reg n_n9599;

reg n_n7635;

reg n_n8984;

reg n_n7360;

reg n_n8794;

reg n_n9108;

reg n_n9286;

reg ndn3_12;

reg ndn3_16;

reg n_n7708;

reg n_n7807;

reg n_n7650;

reg n_n7947;

reg n_n9500;

reg n_n7734;

reg n_n8464;

reg n_n7659;

reg n_n7630;

reg n_n7756;

reg n_n8691;

reg n_n9176;

reg n_n9327;

reg n_n7995;

reg n_n7395;

reg n_n7878;

reg n_n7507;

reg n_n7959;

reg n_n7825;

reg n_n8009;

reg n_n8281;

reg n_n7685;

reg n_n8106;

reg n_n7687;

reg n_n7766;

reg n_n7880;

reg n_n8961;

reg n_n8014;

reg n_n9278;

reg n_n9087;

reg n_n9182;

reg n_n7852;

reg n_n9324;

reg nak3_13;

reg n_n9416;

reg nsr3_14;

reg n_n8603;

reg n_n7026;

reg n_n8856;

reg n_n8272;

reg n_n9312;

reg n_n7985;

reg n_n8312;

reg n_n7231;

reg n_n9396;

reg n_n8801;

reg n_n8683;

reg ndn3_39;

reg n_n8245;

reg n_n9458;

reg n_n9302;

reg n_n7392;

reg n_n6963;

reg n_n7808;

reg n_n7225;

reg n_n7817;

reg n_n8201;

reg n_n7793;

reg n_n8177;

reg n_n8389;

reg n_n9440;

reg n_n7683;

reg n_n7761;

reg n_n7667;

reg n_n7980;

reg n_n7509;

reg n_n7813;

reg n_n8396;

reg n_n9535;

reg n_n7209;

reg n_n7003;

reg n_n7695;

reg n_n7624;

reg n_n8791;

reg n_n7374;

reg n_n7429;

reg n_n7944;

reg n_n9266;

reg n_n8100;

reg n_n6988;

reg n_n6986;

reg n_n8933;

reg n_n7117;

reg n_n9043;

reg n_n8241;

reg n_n9219;

reg n_n8198;

reg n_n8081;

reg n_n8575;

reg n_n8710;

reg n_n7622;

reg n_n7966;

reg n_n7885;

reg n_n7033;

reg ndn3_34;

reg n_n9186;

reg ndn3_50;

reg n_n7879;

reg n_n7019;

reg n_n9171;

reg n_n7261;

reg n_n8223;

reg n_n8989;

reg n_n7993;

reg n_n7845;

reg n_n8253;

reg n_n8889;

reg n_n7809;

reg n_n8918;

reg n_n8515;

reg n_n7933;

reg n_n8075;

reg n_n7338;

reg n_n8104;

reg n_n8171;

reg n_n9059;

reg n_n9023;

reg n_n7692;

reg n_n9441;

reg n_n6920;

reg n_n8831;

reg n_n8441;

reg n_n9576;

reg n_n9252;

reg n_n9363;

reg ndn3_4;

reg n_n9247;

reg n_n7561;

reg n_n8923;

reg n_n7978;

reg n_n8978;

reg n_n9499;

reg n_n8713;

reg n_n8944;

reg n_n8239;

reg n_n7652;

reg n_n9042;

reg n_n8530;

reg n_n9271;

reg n_n9318;

reg n_n7706;

reg n_n7964;

reg n_n8222;

reg n_n8898;

reg n_n7976;

reg n_n7649;

reg n_n7604;

reg n_n7961;

reg n_n7424;

reg n_n7476;

reg n_n9259;

reg n_n9309;

reg n_n9161;

reg n_n8436;

reg n_n9121;

reg n_n8061;

reg n_n8004;

reg n_n9360;

reg n_n9205;

reg n_n8392;

reg n_n9034;

reg n_n8375;

reg n_n8328;

reg n_n9298;

reg n_n7598;

reg n_n8506;

reg pdn;

reg n_n7737;

reg n_n7420;

reg n_n9291;

reg n_n7946;

reg n_n8584;

reg n_n9308;

reg n_n9403;

reg n_n7284;

reg n_n9270;

reg n_n7390;

reg n_n9351;

reg n_n6968;

reg n_n8668;

reg n_n9605;

reg n_n7013;

reg n_n9626;

reg n_n8200;

reg n_n9028;

reg n_n8803;

reg n_n9570;

reg n_n8366;

reg n_n9050;

reg n_n8650;

reg n_n8574;

reg n_n7276;

reg n_n9212;

reg n_n8384;

reg ndn3_35;

reg n_n8449;

reg ndn3_46;

reg n_n7554;

reg n_n8743;

reg n_n8277;

reg n_n9359;

reg n_n8425;

reg n_n9104;

reg n_n9221;

reg n_n9448;

reg n_n9537;

reg n_n8003;

reg n_n7467;

reg n_n8233;

reg n_n7932;

reg n_n8064;

reg n_n9162;

reg n_n7971;

reg n_n8055;

reg n_n7711;

reg n_n8256;

reg n_n7925;

reg n_n7762;

reg n_n7668;

reg n_n7914;

reg n_n7873;

reg n_n7849;

reg n_n9421;

reg n_n7626;

reg n_n7848;

reg n_n8263;

reg n_n9100;

reg n_n9393;

reg n_n9591;

reg n_n7588;

reg n_n9123;

reg n_n9159;

reg n_n9128;

reg n_n8045;

reg n_n7728;

reg n_n8929;

reg n_n7739;

reg n_n9355;

reg n_n9394;

reg n_n8470;

reg n_n8571;

reg n_n8796;

reg ndn3_36;

reg n_n7990;

reg n_n8781;

reg n_n8817;

reg n_n9160;

reg n_n9092;

reg n_n8513;

reg n_n8213;

reg n_n8581;

reg n_n9284;

reg n_n7837;

reg n_n8224;

reg n_n9203;

reg n_n7655;

reg n_n8946;

reg n_n7052;

reg n_n9615;

reg n_n8473;

reg n_n7741;

reg n_n9460;

reg n_n7912;

reg n_n7606;

reg n_n9021;

reg n_n7781;

reg n_n7810;

reg n_n7108;

reg n_n7697;

reg n_n7642;

reg n_n9595;

reg n_n7694;

reg n_n8221;

reg n_n7600;

reg n_n7935;

reg n_n9230;

reg n_n7701;

reg n_n7510;

reg n_n7627;

reg n_n8502;

reg n_n8516;

reg n_n7913;

reg n_n9320;

reg n_n7411;

reg n_n9129;

reg n_n9053;

reg n_n7069;

reg n_n8617;

reg n_n7242;

reg n_n8230;

reg n_n9294;

reg n_n8249;

reg n_n8972;

reg n_n7074;

reg n_n7493;

reg n_n8290;

reg n_n8821;

reg n_n7769;

reg n_n7491;

reg n_n9600;

reg n_n9317;

reg n_n8047;

reg n_n9629;

reg n_n9126;

reg n_n9508;

reg n_n9155;

reg n_n8528;

reg ndn3_37;

reg ndn3_42;

reg n_n9358;

reg n_n8185;

reg nen3_28;

reg n_n8839;

reg n_n7903;

reg n_n9139;

reg n_n9075;

reg n_n9439;

reg n_n9353;

reg n_n7665;

reg n_n8798;

reg n_n7146;

reg n_n7890;

reg n_n7176;

reg n_n8477;

reg n_n8514;

reg n_n8636;

reg n_n7183;

reg n_n8657;

reg n_n9493;

reg n_n7969;

reg n_n9255;

reg n_n8535;

reg n_n8619;

reg n_n8909;

reg n_n7744;

reg n_n9119;

reg n_n7827;

reg n_n8916;

reg n_n8729;

reg n_n9011;

reg n_n8779;

reg n_n6980;

reg n_n7715;

reg n_n9067;

reg n_n9164;

reg n_n7402;

reg n_n8938;

reg n_n9046;

reg n_n8789;

reg n_n9390;

reg n_n7768;

reg n_n9136;

reg n_n8670;

reg n_n8644;

reg n_n9178;

reg n_n8188;

reg n_n7083;

reg n_n9344;

reg n_n7366;

reg n_n8361;

reg n_n9228;

reg n_n9402;

reg n_n8510;

reg n_n8881;

reg n_n9404;

reg n_n9424;

reg n_n9031;

reg nsr3_37;

reg n_n8197;

reg n_n8468;

reg n_n7121;

reg n_n7511;

reg ndn3_44;

reg n_n9322;

reg n_n7682;

reg n_n9603;

reg nlc1_2;

reg n_n8408;

reg n_n8577;

reg n_n7079;

reg n_n8828;

reg n_n9340;

reg n_n8586;

reg n_n7901;

reg n_n8628;

reg n_n8869;

reg n_n7710;

reg n_n8993;

reg n_n9586;

reg n_n8852;

reg n_n8583;

reg n_n8011;

reg n_n7717;

reg n_n8326;

reg n_n9163;

reg n_n8344;

reg n_n8296;

reg n_n8116;

reg n_n8267;

reg n_n7686;

reg n_n9061;

reg n_n9338;

reg n_n7688;

reg n_n9081;

reg n_n6910;

reg n_n8727;

reg n_n7674;

reg n_n7330;

reg n_n8966;

reg n_n7843;

reg n_n8847;

reg n_n9376;

reg n_n7553;

reg n_n9292;

reg n_n7464;

reg n_n8146;

reg n_n8439;

reg n_n9498;

reg n_n8118;

reg n_n9452;

reg n_n9239;

reg n_n9237;

reg n_n9488;

reg ndn3_2;

reg n_n9522;

reg n_n9313;

reg n_n7435;

reg n_n8665;

reg n_n9593;

reg n_n8303;

reg n_n7022;

reg n_n9173;

reg n_n9261;

reg n_n7150;

reg n_n9455;

reg n_n8371;

reg nsr3_20;

reg n_n8271;

reg n_n9542;

reg n_n7444;

reg ndn3_40;

reg n_n7130;

reg n_n9347;

reg n_n8102;

reg n_n9225;

reg n_n8462;

reg n_n8088;

reg n_n9026;

reg n_n9289;

reg n_n7661;

reg n_n8108;

reg n_n8921;

reg n_n7859;

reg n_n7732;

reg n_n7956;

reg n_n9520;

reg n_n7666;

reg n_n7678;

reg n_n7846;

reg n_n8280;

reg n_n8841;

reg n_n7336;

reg n_n8226;

reg n_n8151;

reg n_n7644;

reg n_n8770;

reg n_n8423;

reg n_n7763;

reg n_n9525;

reg n_n8033;

reg n_n7881;

reg n_n7815;

reg n_n9232;

reg n_n7792;

reg n_n9563;

reg n_n8672;

reg n_n7346;

reg n_n7949;

reg n_n8756;

reg n_n8641;

reg n_n8192;

reg n_n8058;

reg n_n8561;

reg n_n9306;

reg n_n9165;

reg n_n8850;

reg n_n9210;

reg ndn2_2;

reg n_n7342;

reg n_n8051;

reg n_n7136;

reg n_n9348;

reg n_n9006;

reg n_n7653;

reg n_n7905;

reg n_n9166;

reg n_n7065;

reg n_n9490;

reg n_n7024;

reg n_n7586;

reg n_n8416;

reg n_n8937;

reg n_n8141;

reg n_n7853;

reg n_n8121;

reg n_n9604;

reg n_n9496;

reg n_n8195;

reg n_n9516;

reg n_n9077;

reg n_n9436;

reg n_n9051;

reg n_n7664;

reg n_n8419;

reg n_n7874;

reg n_n9133;

reg n_n9392;

reg n_n7770;

reg ndn3_32;

reg n_n7601;

reg n_n8206;

reg n_n7927;

reg n_n9606;

reg n_n7111;

reg n_n9269;

reg ndn3_38;

reg n_n7886;

reg n_n9179;

reg n_n9357;

reg n_n9594;

reg n_n7628;

reg n_n8454;

reg ndn3_20;

reg n_n9505;

reg nen3_34;

reg n_n9632;

reg n_n7076;

reg n_n9262;

reg n_n9048;

reg n_n9578;

reg n_n8135;

reg ndn3_26;

reg n_n7500;

reg n_n6974;

reg n_n8605;

reg n_n9296;

reg n_n7156;

reg n_n7920;

reg n_n8895;

reg n_n8991;

reg n_n8139;

reg n_n9275;

reg n_n7203;

reg n_n9590;

reg n_n7344;

reg n_n6976;

reg n_n7629;

reg ndn3_14;

reg n_n7862;

reg n_n9013;

reg n_n7288;

reg n_n8078;

reg n_n7334;

reg n_n7704;

reg n_n7788;

reg n_n8526;

reg n_n9556;

reg n_n9345;

reg n_n8447;

reg n_n7485;

reg n_n8570;

reg n_n7453;

reg n_n7928;

reg n_n8646;

reg n_n9405;

reg n_n8948;

reg n_n9131;

reg n_n8216;

reg n_n9177;

reg n_n7844;

reg n_n8811;

reg n_n9145;

reg n_n8428;

reg n_n8858;

reg n_n8580;

always  @(posedge pclk)
	n_n9280<=n_n9279;

 always  @(posedge pclk)
	n_n9172<=n_n8265;

 always  @(posedge pclk)
	n_n9260<=n_n8264;

 always  @(posedge pclk)
	n_n7726<=n_n7724;

 always  @(posedge pclk)
	n_n8270<=n_n8190;

 always  @(posedge pclk)
	n_n8196<=n_n7893;

 always  @(posedge pclk)
	n_n9150<=n_n9149;

 always  @(posedge pclk)
	n_n9267<=n_n7216;

 always  @(posedge pclk)
	n_n7779<=n_n7778;

 always  @(posedge pclk)
	n_n9503<=n_n8834;

 always  @(posedge pclk)
	n_n8150<=n_n8149;

 always  @(posedge pclk)
	n_n9401<=n_n7034;

 always  @(posedge pclk)
	n_n7341<=n_n7166;

 always  @(posedge pclk)
	n_n9180<=n_n7868;

 always  @(posedge pclk)
	n_n8592<=n_n8590;

 always  @(posedge pclk)
	n_n8871<=n_n8870;

 always  @(posedge pclk)
	n_n7252<=n_n7251;

 always  @(posedge pclk)
	n_n7271<=n_n7269;

 always  @(posedge pclk)
	n_n6991<=n_n6990;

 always  @(posedge pclk)
	n_n8557<=n_n7671;

 always  @(posedge pclk)
	n_n7707<=n_n7412;

 always  @(posedge pclk)
	n_n7552<=n_n7201;

 always  @(posedge pclk)
	ndn3_23<=n_n7524;

 always  @(posedge pclk)
	n_n9548<=n_n9545;

 always  @(posedge pclk)
	n_n9467<=n_n9466;

 always  @(posedge pclk)
	n_n8002<=n_n7205;

 always  @(posedge pclk)
	n_n6950<=n_n6949;

 always  @(posedge pclk)
	n_n8930<=n_n7077;

 always  @(posedge pclk)
	n_n7244<=n_n7243;

 always  @(posedge pclk)
	n_n7819<=n_n7369;

 always  @(posedge pclk)
	n_n8883<=n_n8189;

 always  @(posedge pclk)
	n_n7709<=n_n7123;

 always  @(posedge pclk)
	n_n9580<=n_n9579;

 always  @(posedge pclk)
	n_n9130<=n_n6944;

 always  @(posedge pclk)
	n_n9486<=n_n6994;

 always  @(posedge pclk)
	n_n9235<=n_n9234;

 always  @(posedge pclk)
	n_n7522<=n_n7521;

 always  @(posedge pclk)
	n_n7373<=n_n7229;

 always  @(posedge pclk)
	n_n9085<=n_n9084;

 always  @(posedge pclk)
	n_n9638<=n_n7416;

 always  @(posedge pclk)
	n_n7452<=n_n7066;

 always  @(posedge pclk)
	n_n8775<=n_n8774;

 always  @(posedge pclk)
	n_n7654<=n_n7438;

 always  @(posedge pclk)
	n_n8410<=n_n8409;

 always  @(posedge pclk)
	n_n8208<=n_n8207;

 always  @(posedge pclk)
	n_n8377<=n_n8376;

 always  @(posedge pclk)
	n_n7558<=n_n7028;

 always  @(posedge pclk)
	n_n7599<=n_n7421;

 always  @(posedge pclk)
	n_n8225<=n_n7753;

 always  @(posedge pclk)
	n_n8202<=n_n7680;

 always  @(posedge pclk)
	n_n7670<=n_n7669;

 always  @(posedge pclk)
	n_n7888<=n_n7455;

 always  @(posedge pclk)
	n_n7889<=n_n6989;

 always  @(posedge pclk)
	n_n8597<=n_n8596;

 always  @(posedge pclk)
	n_n8152<=n_n7472;

 always  @(posedge pclk)
	n_n8394<=n_n8393;

 always  @(posedge pclk)
	n_n7812<=n_n7591;

 always  @(posedge pclk)
	n_n7816<=n_n7481;

 always  @(posedge pclk)
	n_n9141<=n_n9140;

 always  @(posedge pclk)
	n_n7332<=n_n7331;

 always  @(posedge pclk)
	n_n8758<=n_n8757;

 always  @(posedge pclk)
	n_n7765<=n_n7422;

 always  @(posedge pclk)
	n_n7877<=n_n7040;

 always  @(posedge pclk)
	n_n7814<=n_n7277;

 always  @(posedge pclk)
	n_n9008<=n_n9007;

 always  @(posedge pclk)
	n_n7581<=n_n7580;

 always  @(posedge pclk)
	n_n7376<=n_n7067;

 always  @(posedge pclk)
	n_n7970<=n_n7092;

 always  @(posedge pclk)
	pover_0_0_<=n_n7199;

 always  @(posedge pclk)
	n_n8599<=n_n8598;

 always  @(posedge pclk)
	n_n8227<=n_n7240;

 always  @(posedge pclk)
	n_n9442<=n_n7382;

 always  @(posedge pclk)
	n_n9485<=n_n8411;

 always  @(posedge pclk)
	n_n7148<=n_n7147;

 always  @(posedge pclk)
	n_n9311<=n_n7517;

 always  @(posedge pclk)
	n_n9273<=n_n9250;

 always  @(posedge pclk)
	ndn3_9<=n_n7188;

 always  @(posedge pclk)
	n_n8613<=n_n8612;

 always  @(posedge pclk)
	n_n8533<=n_n8532;

 always  @(posedge pclk)
	n_n8699<=n_n8698;

 always  @(posedge pclk)
	n_n8609<=n_n8608;

 always  @(posedge pclk)
	n_n8308<=n_n8307;

 always  @(posedge pclk)
	n_n8655<=n_n8654;

 always  @(posedge pclk)
	n_n8981<=n_n7125;

 always  @(posedge pclk)
	n_n7583<=n_n7357;

 always  @(posedge pclk)
	n_n9198<=n_n7;

 always  @(posedge pclk)
	n_n9602<=n_n8787;

 always  @(posedge pclk)
	n_n8786<=n_n8785;

 always  @(posedge pclk)
	n_n9598<=n_n7473;

 always  @(posedge pclk)
	n_n7738<=n_n7214;

 always  @(posedge pclk)
	n_n8573<=n_n7063;

 always  @(posedge pclk)
	n_n9473<=n_n9472;

 always  @(posedge pclk)
	n_n9000<=n_n8999;

 always  @(posedge pclk)
	n_n8001<=n_n7495;

 always  @(posedge pclk)
	n_n9554<=n_n7266;

 always  @(posedge pclk)
	n_n8508<=n_n8507;

 always  @(posedge pclk)
	n_n9635<=n_n9634;

 always  @(posedge pclk)
	n_n7190<=n_n7189;

 always  @(posedge pclk)
	n_n8702<=n_n8700;

 always  @(posedge pclk)
	n_n9106<=n_n9105;

 always  @(posedge pclk)
	n_n7409<=n_n7408;

 always  @(posedge pclk)
	n_n9437<=n_n7137;

 always  @(posedge pclk)
	n_n9052<=n_n7504;

 always  @(posedge pclk)
	n_n8647<=n_n8527;

 always  @(posedge pclk)
	n_n9265<=n_n9208;

 always  @(posedge pclk)
	n_n7179<=n_n7177;

 always  @(posedge pclk)
	ndn3_13<=n_n7615;

 always  @(posedge pclk)
	ndn3_17<=n_n7087;

 always  @(posedge pclk)
	ndn3_25<=n_n8293;

 always  @(posedge pclk)
	ndn3_29<=n_n8217;

 always  @(posedge pclk)
	n_n9539<=n_n9538;

 always  @(posedge pclk)
	n_n7953<=n_n7091;

 always  @(posedge pclk)
	n_n8488<=n_n8487;

 always  @(posedge pclk)
	nen3_22<=n_n8299;

 always  @(posedge pclk)
	n_n9438<=n_n7796;

 always  @(posedge pclk)
	n_n8132<=n_n8130;

 always  @(posedge pclk)
	n_n8661<=n_n8660;

 always  @(posedge pclk)
	n_n7759<=n_n7325;

 always  @(posedge pclk)
	n_n8333<=n_n8332;

 always  @(posedge pclk)
	n_n9399<=n_n7037;

 always  @(posedge pclk)
	n_n7798<=n_n7797;

 always  @(posedge pclk)
	n_n9434<=n_n7005;

 always  @(posedge pclk)
	n_n7910<=n_n7200;

 always  @(posedge pclk)
	n_n9528<=n_n9527;

 always  @(posedge pclk)
	n_n7850<=n_n7523;

 always  @(posedge pclk)
	n_n8251<=n_n8250;

 always  @(posedge pclk)
	n_n7937<=n_n7483;

 always  @(posedge pclk)
	n_n8482<=n_n8481;

 always  @(posedge pclk)
	n_n9290<=n_n7451;

 always  @(posedge pclk)
	n_n8007<=n_n7055;

 always  @(posedge pclk)
	n_n7556<=n_n7555;

 always  @(posedge pclk)
	n_n9064<=n_n9063;

 always  @(posedge pclk)
	n_n9398<=n_n7207;

 always  @(posedge pclk)
	n_n9412<=n_n7100;

 always  @(posedge pclk)
	n_n9361<=n_n7799;

 always  @(posedge pclk)
	n_n9304<=n_n7471;

 always  @(posedge pclk)
	n_n7651<=n_n7219;

 always  @(posedge pclk)
	n_n7712<=n_n7614;

 always  @(posedge pclk)
	n_n7735<=n_n7250;

 always  @(posedge pclk)
	n_n7934<=n_n7590;

 always  @(posedge pclk)
	n_n7811<=n_n6915;

 always  @(posedge pclk)
	n_n8053<=n_n8052;

 always  @(posedge pclk)
	n_n9015<=n_n9014;

 always  @(posedge pclk)
	n_n8066<=n_n8065;

 always  @(posedge pclk)
	n_n9518<=n_n9517;

 always  @(posedge pclk)
	n_n8091<=n_n8089;

 always  @(posedge pclk)
	n_n9257<=n_n9256;

 always  @(posedge pclk)
	n_n8175<=n_n8174;

 always  @(posedge pclk)
	n_n8491<=n_n8490;

 always  @(posedge pclk)
	n_n8114<=n_n8113;

 always  @(posedge pclk)
	n_n7951<=n_n7039;

 always  @(posedge pclk)
	n_n8913<=n_n7095;

 always  @(posedge pclk)
	n_n8035<=n_n8034;

 always  @(posedge pclk)
	n_n8631<=n_n7094;

 always  @(posedge pclk)
	n_n8243<=n_n8242;

 always  @(posedge pclk)
	n_n7857<=n_n7855;

 always  @(posedge pclk)
	ngfdn_3<=n_n7098;

 always  @(posedge pclk)
	n_n7791<=n_n7632;

 always  @(posedge pclk)
	n_n9175<=n_n9079;

 always  @(posedge pclk)
	n_n9588<=n_n7090;

 always  @(posedge pclk)
	n_n9049<=n_n7299;

 always  @(posedge pclk)
	n_n9483<=n_n9480;

 always  @(posedge pclk)
	n_n9410<=n_n9409;

 always  @(posedge pclk)
	n_n7691<=n_n7385;

 always  @(posedge pclk)
	n_n7740<=n_n7406;

 always  @(posedge pclk)
	n_n7602<=n_n7405;

 always  @(posedge pclk)
	n_n7783<=n_n7782;

 always  @(posedge pclk)
	n_n7948<=n_n7372;

 always  @(posedge pclk)
	n_n7054<=n_n7053;

 always  @(posedge pclk)
	n_n9343<=n_n7086;

 always  @(posedge pclk)
	n_n9400<=n_n8730;

 always  @(posedge pclk)
	nsr1_2<=n_n1;

 always  @(posedge pclk)
	n_n9127<=n_n9090;

 always  @(posedge pclk)
	n_n8531<=n_n7547;

 always  @(posedge pclk)
	n_n9335<=n_n8335;

 always  @(posedge pclk)
	n_n7324<=n_n7323;

 always  @(posedge pclk)
	n_n9611<=n_n9610;

 always  @(posedge pclk)
	n_n8112<=n_n8111;

 always  @(posedge pclk)
	n_n9406<=n_n8039;

 always  @(posedge pclk)
	n_n9618<=n_n9617;

 always  @(posedge pclk)
	n_n9613<=n_n9612;

 always  @(posedge pclk)
	n_n9242<=n_n9241;

 always  @(posedge pclk)
	n_n7384<=n_n7383;

 always  @(posedge pclk)
	n_n8884<=n_n6933;

 always  @(posedge pclk)
	n_n7462<=n_n7461;

 always  @(posedge pclk)
	n_n7908<=n_n7613;

 always  @(posedge pclk)
	n_n8765<=n_n8764;

 always  @(posedge pclk)
	n_n7909<=n_n7014;

 always  @(posedge pclk)
	n_n7898<=n_n7897;

 always  @(posedge pclk)
	n_n9135<=n_n8379;

 always  @(posedge pclk)
	n_n8862<=n_n8861;

 always  @(posedge pclk)
	n_n8037<=n_n8036;

 always  @(posedge pclk)
	ndn3_18<=n_n8026;

 always  @(posedge pclk)
	ndn3_22<=n_n7883;

 always  @(posedge pclk)
	n_n8974<=n_n8973;

 always  @(posedge pclk)
	n_n7286<=n_n7285;

 always  @(posedge pclk)
	n_n9223<=n_n9222;

 always  @(posedge pclk)
	n_n7306<=n_n8147;

 always  @(posedge pclk)
	n_n9169<=n_n9167;

 always  @(posedge pclk)
	n_n9125<=n_n8310;

 always  @(posedge pclk)
	nen3_39<=n_n8317;

 always  @(posedge pclk)
	n_n8278<=n_n7168;

 always  @(posedge pclk)
	n_n9557<=n_n7397;

 always  @(posedge pclk)
	n_n7758<=n_n7165;

 always  @(posedge pclk)
	n_n9391<=n_n7070;

 always  @(posedge pclk)
	n_n8110<=n_n8109;

 always  @(posedge pclk)
	n_n9597<=n_n7268;

 always  @(posedge pclk)
	n_n8568<=n_n8567;

 always  @(posedge pclk)
	n_n7428<=n_n7228;

 always  @(posedge pclk)
	n_n7931<=n_n7718;

 always  @(posedge pclk)
	n_n7742<=n_n7494;

 always  @(posedge pclk)
	n_n7236<=n_n7235;

 always  @(posedge pclk)
	n_n8219<=n_n8218;

 always  @(posedge pclk)
	n_n9568<=n_n9567;

 always  @(posedge pclk)
	n_n9200<=n_n9199;

 always  @(posedge pclk)
	n_n8545<=n_n8544;

 always  @(posedge pclk)
	n_n7823<=n_n6934;

 always  @(posedge pclk)
	n_n8005<=n_n6914;

 always  @(posedge pclk)
	n_n8736<=n_n8735;

 always  @(posedge pclk)
	n_n9339<=n_n8474;

 always  @(posedge pclk)
	n_n8499<=n_n8498;

 always  @(posedge pclk)
	n_n8086<=n_n8085;

 always  @(posedge pclk)
	n_n7803<=n_n7802;

 always  @(posedge pclk)
	n_n7640<=n_n7061;

 always  @(posedge pclk)
	n_n9098<=n_n9097;

 always  @(posedge pclk)
	n_n7160<=n_n7159;

 always  @(posedge pclk)
	n_n7713<=n_n7303;

 always  @(posedge pclk)
	n_n9566<=n_n9565;

 always  @(posedge pclk)
	n_n7955<=n_n7833;

 always  @(posedge pclk)
	n_n8414<=n_n8413;

 always  @(posedge pclk)
	n_n8006<=n_n6969;

 always  @(posedge pclk)
	n_n9560<=n_n8345;

 always  @(posedge pclk)
	n_n8742<=n_n7800;

 always  @(posedge pclk)
	n_n7174<=n_n7172;

 always  @(posedge pclk)
	n_n8882<=n_n7212;

 always  @(posedge pclk)
	n_n7546<=n_n7545;

 always  @(posedge pclk)
	n_n8282<=n_n7099;

 always  @(posedge pclk)
	n_n8998<=n_n8997;

 always  @(posedge pclk)
	n_n7656<=n_n7479;

 always  @(posedge pclk)
	n_n9465<=n_n9463;

 always  @(posedge pclk)
	n_n9601<=n_n8346;

 always  @(posedge pclk)
	n_n8875<=n_n8874;

 always  @(posedge pclk)
	n_n7954<=n_n7354;

 always  @(posedge pclk)
	n_n8959<=n_n8958;

 always  @(posedge pclk)
	n_n8957<=n_n8956;

 always  @(posedge pclk)
	n_n8247<=n_n8246;

 always  @(posedge pclk)
	n_n8258<=n_n8257;

 always  @(posedge pclk)
	n_n7641<=n_n7404;

 always  @(posedge pclk)
	n_n8843<=n_n8842;

 always  @(posedge pclk)
	n_n9321<=n_n8443;

 always  @(posedge pclk)
	n_n7702<=n_n7163;

 always  @(posedge pclk)
	nsr3_23<=n_n6;

 always  @(posedge pclk)
	n_n8199<=n_n8025;

 always  @(posedge pclk)
	n_n7983<=n_n7982;

 always  @(posedge pclk)
	n_n7217<=n_n7186;

 always  @(posedge pclk)
	n_n7821<=n_n7248;

 always  @(posedge pclk)
	n_n9489<=n_n7639;

 always  @(posedge pclk)
	n_n8348<=n_n8347;

 always  @(posedge pclk)
	n_n9408<=n_n8835;

 always  @(posedge pclk)
	n_n8445<=n_n8444;

 always  @(posedge pclk)
	n_n9501<=n_n7425;

 always  @(posedge pclk)
	n_n7831<=n_n7830;

 always  @(posedge pclk)
	n_n7757<=n_n7618;

 always  @(posedge pclk)
	n_n9174<=n_n9062;

 always  @(posedge pclk)
	n_n9432<=n_n9430;

 always  @(posedge pclk)
	n_n8678<=n_n8676;

 always  @(posedge pclk)
	n_n8024<=n_n8023;

 always  @(posedge pclk)
	n_n7806<=n_n7141;

 always  @(posedge pclk)
	n_n8996<=n_n8995;

 always  @(posedge pclk)
	n_n7918<=n_n7917;

 always  @(posedge pclk)
	n_n8260<=n_n8259;

 always  @(posedge pclk)
	n_n9341<=n_n9207;

 always  @(posedge pclk)
	n_n9189<=n_n9188;

 always  @(posedge pclk)
	n_n9096<=n_n9094;

 always  @(posedge pclk)
	ndn3_30<=n_n8179;

 always  @(posedge pclk)
	n_n7775<=n_n7773;

 always  @(posedge pclk)
	n_n7693<=n_n7647;

 always  @(posedge pclk)
	nen3_16<=n_n7038;

 always  @(posedge pclk)
	n_n7643<=n_n7157;

 always  @(posedge pclk)
	n_n8941<=n_n8940;

 always  @(posedge pclk)
	n_n8042<=n_n8041;

 always  @(posedge pclk)
	n_n8681<=n_n8679;

 always  @(posedge pclk)
	n_n8659<=n_n8658;

 always  @(posedge pclk)
	n_n9110<=n_n9109;

 always  @(posedge pclk)
	n_n9573<=n_n9572;

 always  @(posedge pclk)
	n_n8951<=n_n8950;

 always  @(posedge pclk)
	n_n9589<=n_n9240;

 always  @(posedge pclk)
	n_n9387<=n_n9386;

 always  @(posedge pclk)
	n_n8279<=n_n7594;

 always  @(posedge pclk)
	n_n7790<=n_n7210;

 always  @(posedge pclk)
	n_n8406<=n_n8405;

 always  @(posedge pclk)
	n_n8582<=n_n7892;

 always  @(posedge pclk)
	n_n7911<=n_n7221;

 always  @(posedge pclk)
	n_n7474<=n_n7350;

 always  @(posedge pclk)
	n_n8466<=n_n8465;

 always  @(posedge pclk)
	n_n6984<=n_n6983;

 always  @(posedge pclk)
	n_n7760<=n_n7719;

 always  @(posedge pclk)
	n_n7847<=n_n7551;

 always  @(posedge pclk)
	n_n9559<=n_n8737;

 always  @(posedge pclk)
	n_n7362<=n_n7361;

 always  @(posedge pclk)
	n_n9300<=n_n9299;

 always  @(posedge pclk)
	n_n9550<=n_n9549;

 always  @(posedge pclk)
	n_n9492<=n_n9287;

 always  @(posedge pclk)
	n_n8777<=n_n8776;

 always  @(posedge pclk)
	n_n7764<=n_n7009;

 always  @(posedge pclk)
	n_n7826<=n_n7355;

 always  @(posedge pclk)
	n_n7777<=n_n7776;

 always  @(posedge pclk)
	n_n7824<=n_n7550;

 always  @(posedge pclk)
	n_n8173<=n_n8172;

 always  @(posedge pclk)
	n_n7498<=n_n7497;

 always  @(posedge pclk)
	n_n9148<=n_n9146;

 always  @(posedge pclk)
	n_n8753<=n_n8752;

 always  @(posedge pclk)
	n_n8772<=n_n8771;

 always  @(posedge pclk)
	n_n8049<=n_n8048;

 always  @(posedge pclk)
	n_n9362<=n_n7870;

 always  @(posedge pclk)
	ndn1_4<=n_n7015;

 always  @(posedge pclk)
	n_n9561<=n_n7470;

 always  @(posedge pclk)
	n_n9004<=n_n9002;

 always  @(posedge pclk)
	n_n8203<=n_n7532;

 always  @(posedge pclk)
	n_n8153<=n_n7442;

 always  @(posedge pclk)
	n_n9263<=n_n9078;

 always  @(posedge pclk)
	n_n8369<=n_n8367;

 always  @(posedge pclk)
	n_n9331<=n_n9330;

 always  @(posedge pclk)
	n_n7454<=n_n7103;

 always  @(posedge pclk)
	ndn3_7<=n_n8399;

 always  @(posedge pclk)
	n_n7527<=n_n7526;

 always  @(posedge pclk)
	n_n9036<=n_n9035;

 always  @(posedge pclk)
	n_n7875<=n_n7264;

 always  @(posedge pclk)
	n_n8697<=n_n8696;

 always  @(posedge pclk)
	n_n9497<=n_n7080;

 always  @(posedge pclk)
	n_n7291<=n_n7290;

 always  @(posedge pclk)
	nsr3_13<=n_n11;

 always  @(posedge pclk)
	nsr3_38<=n_n2;

 always  @(posedge pclk)
	n_n8240<=n_n7548;

 always  @(posedge pclk)
	n_n7703<=n_n7294;

 always  @(posedge pclk)
	n_n9282<=n_n8949;

 always  @(posedge pclk)
	n_n8237<=n_n7633;

 always  @(posedge pclk)
	n_n8935<=n_n8934;

 always  @(posedge pclk)
	n_n9244<=n_n9243;

 always  @(posedge pclk)
	n_n8648<=n_n7194;

 always  @(posedge pclk)
	n_n8235<=n_n7465;

 always  @(posedge pclk)
	n_n8611<=n_n8610;

 always  @(posedge pclk)
	n_n9045<=n_n7746;

 always  @(posedge pclk)
	n_n9334<=n_n7349;

 always  @(posedge pclk)
	n_n8572<=n_n8169;

 always  @(posedge pclk)
	n_n9491<=n_n7316;

 always  @(posedge pclk)
	n_n9134<=n_n8495;

 always  @(posedge pclk)
	n_n9555<=n_n6995;

 always  @(posedge pclk)
	n_n9336<=n_n7468;

 always  @(posedge pclk)
	n_n7050<=n_n7049;

 always  @(posedge pclk)
	n_n9346<=n_n7304;

 always  @(posedge pclk)
	n_n7140<=n_n7139;

 always  @(posedge pclk)
	n_n7681<=n_n7142;

 always  @(posedge pclk)
	n_n6948<=n_n6947;

 always  @(posedge pclk)
	n_n8549<=n_n8548;

 always  @(posedge pclk)
	ndn3_19<=n_n9543;

 always  @(posedge pclk)
	ndn3_28<=n_n9620;

 always  @(posedge pclk)
	n_n7102<=n_n7101;

 always  @(posedge pclk)
	n_n8093<=n_n8092;

 always  @(posedge pclk)
	n_n9041<=n_n8624;

 always  @(posedge pclk)
	n_n8381<=n_n8380;

 always  @(posedge pclk)
	n_n8810<=n_n6965;

 always  @(posedge pclk)
	nen3_36<=n_n7891;

 always  @(posedge pclk)
	n_n9047<=n_n8907;

 always  @(posedge pclk)
	n_n9333<=n_n7571;

 always  @(posedge pclk)
	n_n7736<=n_n7559;

 always  @(posedge pclk)
	n_n7820<=n_n7612;

 always  @(posedge pclk)
	n_n8986<=n_n8985;

 always  @(posedge pclk)
	n_n8891<=n_n8890;

 always  @(posedge pclk)
	n_n8000<=n_n7999;

 always  @(posedge pclk)
	n_n7968<=n_n7220;

 always  @(posedge pclk)
	n_n8750<=n_n8748;

 always  @(posedge pclk)
	n_n9558<=n_n6942;

 always  @(posedge pclk)
	n_n9368<=n_n9367;

 always  @(posedge pclk)
	n_n8519<=n_n8518;

 always  @(posedge pclk)
	n_n6956<=n_n6955;

 always  @(posedge pclk)
	n_n8298<=n_n8297;

 always  @(posedge pclk)
	n_n9397<=n_n6922;

 always  @(posedge pclk)
	n_n7017<=n_n7016;

 always  @(posedge pclk)
	n_n8638<=n_n8637;

 always  @(posedge pclk)
	n_n9552<=n_n9551;

 always  @(posedge pclk)
	n_n8964<=n_n8286;

 always  @(posedge pclk)
	n_n8016<=n_n8015;

 always  @(posedge pclk)
	n_n7603<=n_n7345;

 always  @(posedge pclk)
	n_n7696<=n_n7010;

 always  @(posedge pclk)
	n_n8589<=n_n8587;

 always  @(posedge pclk)
	n_n9337<=n_n7097;

 always  @(posedge pclk)
	n_n9132<=n_n6953;

 always  @(posedge pclk)
	n_n8652<=n_n8457;

 always  @(posedge pclk)
	n_n8707<=n_n7940;

 always  @(posedge pclk)
	n_n9407<=n_n8163;

 always  @(posedge pclk)
	n_n9044<=n_n8860;

 always  @(posedge pclk)
	n_n8808<=n_n7319;

 always  @(posedge pclk)
	nsr3_30<=n_n5;

 always  @(posedge pclk)
	n_n8274<=n_n6924;

 always  @(posedge pclk)
	n_n8615<=n_n8614;

 always  @(posedge pclk)
	n_n8238<=n_n6941;

 always  @(posedge pclk)
	n_n7854<=n_n7000;

 always  @(posedge pclk)
	n_n8649<=n_n7280;

 always  @(posedge pclk)
	n_n8236<=n_n8137;

 always  @(posedge pclk)
	n_n8269<=n_n7313;

 always  @(posedge pclk)
	n_n9592<=n_n7832;

 always  @(posedge pclk)
	n_n8022<=n_n8021;

 always  @(posedge pclk)
	n_n8744<=n_n8517;

 always  @(posedge pclk)
	n_n8529<=n_n8136;

 always  @(posedge pclk)
	n_n7967<=n_n7122;

 always  @(posedge pclk)
	n_n9487<=n_n7616;

 always  @(posedge pclk)
	n_n8685<=n_n8684;

 always  @(posedge pclk)
	n_n9531<=n_n9529;

 always  @(posedge pclk)
	n_n9510<=n_n9509;

 always  @(posedge pclk)
	n_n7771<=n_n7042;

 always  @(posedge pclk)
	n_n8480<=n_n8479;

 always  @(posedge pclk)
	n_n8543<=n_n8542;

 always  @(posedge pclk)
	n_n7789<=n_n7088;

 always  @(posedge pclk)
	ndn3_11<=n_n7096;

 always  @(posedge pclk)
	ndn3_15<=n_n8878;

 always  @(posedge pclk)
	ndn3_21<=n_n8331;

 always  @(posedge pclk)
	n_n7584<=n_n7301;

 always  @(posedge pclk)
	n_n8354<=n_n7972;

 always  @(posedge pclk)
	n_n6952<=n_n6951;

 always  @(posedge pclk)
	n_n8864<=n_n8863;

 always  @(posedge pclk)
	n_n7930<=n_n6993;

 always  @(posedge pclk)
	n_n7962<=n_n7057;

 always  @(posedge pclk)
	n_n7929<=n_n7143;

 always  @(posedge pclk)
	n_n9316<=n_n6945;

 always  @(posedge pclk)
	n_n9102<=n_n9101;

 always  @(posedge pclk)
	n_n7308<=n_n7307;

 always  @(posedge pclk)
	n_n7657<=n_n7300;

 always  @(posedge pclk)
	n_n9264<=n_n7036;

 always  @(posedge pclk)
	n_n8760<=n_n8759;

 always  @(posedge pclk)
	n_n6912<=n_n6911;

 always  @(posedge pclk)
	n_n7887<=n_n7352;

 always  @(posedge pclk)
	n_n8911<=n_n7535;

 always  @(posedge pclk)
	n_n7952<=n_n7457;

 always  @(posedge pclk)
	n_n8704<=n_n8703;

 always  @(posedge pclk)
	n_n7876<=n_n7520;

 always  @(posedge pclk)
	n_n9596<=n_n8475;

 always  @(posedge pclk)
	n_n8430<=n_n8429;

 always  @(posedge pclk)
	n_n9019<=n_n9018;

 always  @(posedge pclk)
	n_n7699<=n_n7698;

 always  @(posedge pclk)
	n_n7375<=n_n6972;

 always  @(posedge pclk)
	n_n7936<=n_n7480;

 always  @(posedge pclk)
	n_n8340<=n_n8338;

 always  @(posedge pclk)
	n_n8809<=n_n7213;

 always  @(posedge pclk)
	n_n6961<=n_n6960;

 always  @(posedge pclk)
	n_n9429<=n_n9427;

 always  @(posedge pclk)
	n_n7743<=n_n7478;

 always  @(posedge pclk)
	n_n8980<=n_n7060;

 always  @(posedge pclk)
	n_n7582<=n_n7318;

 always  @(posedge pclk)
	n_n8968<=n_n8967;

 always  @(posedge pclk)
	n_n9371<=n_n9369;

 always  @(posedge pclk)
	n_n8741<=n_n7320;

 always  @(posedge pclk)
	n_n9502<=n_n7867;

 always  @(posedge pclk)
	n_n9373<=n_n9372;

 always  @(posedge pclk)
	n_n9248<=n_n10;

 always  @(posedge pclk)
	n_n7822<=n_n6940;

 always  @(posedge pclk)
	n_n9054<=n_n6925;

 always  @(posedge pclk)
	n_n8273<=n_n7007;

 always  @(posedge pclk)
	n_n6937<=n_n6936;

 always  @(posedge pclk)
	n_n9342<=n_n7198;

 always  @(posedge pclk)
	n_n9325<=n_n8547;

 always  @(posedge pclk)
	n_n9609<=n_n6954;

 always  @(posedge pclk)
	n_n9623<=n_n9622;

 always  @(posedge pclk)
	n_n9470<=n_n9469;

 always  @(posedge pclk)
	n_n7570<=n_n7569;

 always  @(posedge pclk)
	n_n9310<=n_n7339;

 always  @(posedge pclk)
	n_n9366<=n_n9364;

 always  @(posedge pclk)
	n_n7181<=n_n7180;

 always  @(posedge pclk)
	n_n8739<=n_n8738;

 always  @(posedge pclk)
	n_n8939<=n_n6932;

 always  @(posedge pclk)
	n_n7256<=n_n7255;

 always  @(posedge pclk)
	n_n8983<=n_n7519;

 always  @(posedge pclk)
	n_n7487<=n_n7486;

 always  @(posedge pclk)
	n_n9268<=n_n7259;

 always  @(posedge pclk)
	n_n8906<=n_n8460;

 always  @(posedge pclk)
	n_n7988<=n_n7987;

 always  @(posedge pclk)
	n_n9181<=n_n8378;

 always  @(posedge pclk)
	n_n8725<=n_n8724;

 always  @(posedge pclk)
	n_n8626<=n_n8625;

 always  @(posedge pclk)
	ndn3_27<=n_n9082;

 always  @(posedge pclk)
	n_n8210<=n_n8209;

 always  @(posedge pclk)
	n_n7415<=n_n7414;

 always  @(posedge pclk)
	n_n8900<=n_n8899;

 always  @(posedge pclk)
	nen3_19<=n_n7477;

 always  @(posedge pclk)
	n_n8762<=n_n8761;

 always  @(posedge pclk)
	n_n8512<=n_n7996;

 always  @(posedge pclk)
	n_n8095<=n_n8094;

 always  @(posedge pclk)
	n_n8982<=n_n7112;

 always  @(posedge pclk)
	n_n7387<=n_n7386;

 always  @(posedge pclk)
	n_n9494<=n_n8768;

 always  @(posedge pclk)
	n_n7689<=n_n7611;

 always  @(posedge pclk)
	n_n7835<=n_n7834;

 always  @(posedge pclk)
	n_n9157<=n_n9156;

 always  @(posedge pclk)
	n_n8552<=n_n8551;

 always  @(posedge pclk)
	n_n7381<=n_n7380;

 always  @(posedge pclk)
	n_n9446<=n_n9445;

 always  @(posedge pclk)
	n_n8633<=n_n8632;

 always  @(posedge pclk)
	n_n7684<=n_n7353;

 always  @(posedge pclk)
	n_n7310<=n_n7309;

 always  @(posedge pclk)
	n_n8402<=n_n8401;

 always  @(posedge pclk)
	n_n9315<=n_n7488;

 always  @(posedge pclk)
	n_n7950<=n_n7733;

 always  @(posedge pclk)
	n_n8504<=n_n8503;

 always  @(posedge pclk)
	n_n8456<=n_n8455;

 always  @(posedge pclk)
	n_n7514<=n_n7512;

 always  @(posedge pclk)
	n_n7315<=n_n7314;

 always  @(posedge pclk)
	n_n9476<=n_n9474;

 always  @(posedge pclk)
	n_n8276<=n_n8275;

 always  @(posedge pclk)
	n_n8833<=n_n8832;

 always  @(posedge pclk)
	n_n7923<=n_n7921;

 always  @(posedge pclk)
	n_n9395<=n_n7105;

 always  @(posedge pclk)
	n_n9512<=n_n9511;

 always  @(posedge pclk)
	n_n9319<=n_n8763;

 always  @(posedge pclk)
	nsr3_35<=n_n4;

 always  @(posedge pclk)
	n_n7154<=n_n7153;

 always  @(posedge pclk)
	n_n9495<=n_n8754;

 always  @(posedge pclk)
	n_n9137<=n_n7592;

 always  @(posedge pclk)
	n_n8854<=n_n8853;

 always  @(posedge pclk)
	n_n9183<=n_n8620;

 always  @(posedge pclk)
	n_n9323<=n_n9214;

 always  @(posedge pclk)
	n_n9349<=n_n8987;

 always  @(posedge pclk)
	n_n7896<=n_n7895;

 always  @(posedge pclk)
	n_n8073<=n_n8071;

 always  @(posedge pclk)
	n_n8970<=n_n8969;

 always  @(posedge pclk)
	n_n9314<=n_n8714;

 always  @(posedge pclk)
	n_n8486<=n_n8485;

 always  @(posedge pclk)
	n_n7246<=n_n7245;

 always  @(posedge pclk)
	n_n7866<=n_n7865;

 always  @(posedge pclk)
	n_n9599<=n_n8336;

 always  @(posedge pclk)
	n_n7635<=n_n7634;

 always  @(posedge pclk)
	n_n8984<=n_n7508;

 always  @(posedge pclk)
	n_n7360<=n_n7359;

 always  @(posedge pclk)
	n_n8794<=n_n8559;

 always  @(posedge pclk)
	n_n9108<=n_n9107;

 always  @(posedge pclk)
	n_n9286<=n_n9285;

 always  @(posedge pclk)
	ndn3_12<=n_n7460;

 always  @(posedge pclk)
	ndn3_16<=n_n8540;

 always  @(posedge pclk)
	n_n7708<=n_n7296;

 always  @(posedge pclk)
	n_n7807<=n_n7192;

 always  @(posedge pclk)
	n_n7650<=n_n7058;

 always  @(posedge pclk)
	n_n7947<=n_n7297;

 always  @(posedge pclk)
	n_n9500<=n_n9213;

 always  @(posedge pclk)
	n_n7734<=n_n7370;

 always  @(posedge pclk)
	n_n8464<=n_n8463;

 always  @(posedge pclk)
	n_n7659<=n_n7658;

 always  @(posedge pclk)
	n_n7630<=n_n7238;

 always  @(posedge pclk)
	n_n7756<=n_n7109;

 always  @(posedge pclk)
	n_n8691<=n_n8690;

 always  @(posedge pclk)
	n_n9176<=n_n6943;

 always  @(posedge pclk)
	n_n9327<=n_n9326;

 always  @(posedge pclk)
	n_n7995<=n_n7994;

 always  @(posedge pclk)
	n_n7395<=n_n7394;

 always  @(posedge pclk)
	n_n7878<=n_n7589;

 always  @(posedge pclk)
	n_n7507<=n_n7506;

 always  @(posedge pclk)
	n_n7959<=n_n7958;

 always  @(posedge pclk)
	n_n7825<=n_n7503;

 always  @(posedge pclk)
	n_n8009<=n_n8008;

 always  @(posedge pclk)
	n_n8281<=n_n7562;

 always  @(posedge pclk)
	n_n7685<=n_n7223;

 always  @(posedge pclk)
	n_n8106<=n_n8105;

 always  @(posedge pclk)
	n_n7687<=n_n7456;

 always  @(posedge pclk)
	n_n7766<=n_n7043;

 always  @(posedge pclk)
	n_n7880<=n_n7279;

 always  @(posedge pclk)
	n_n8961<=n_n8960;

 always  @(posedge pclk)
	n_n8014<=n_n8013;

 always  @(posedge pclk)
	n_n9278<=n_n9276;

 always  @(posedge pclk)
	n_n9087<=n_n9086;

 always  @(posedge pclk)
	n_n9182<=n_n7542;

 always  @(posedge pclk)
	n_n7852<=n_n7448;

 always  @(posedge pclk)
	n_n9324<=n_n8164;

 always  @(posedge pclk)
	nak3_13<=n_n8478;

 always  @(posedge pclk)
	n_n9416<=n_n9415;

 always  @(posedge pclk)
	nsr3_14<=n_n9;

 always  @(posedge pclk)
	n_n8603<=n_n0;

 always  @(posedge pclk)
	n_n7026<=n_n7025;

 always  @(posedge pclk)
	n_n8856<=n_n8855;

 always  @(posedge pclk)
	n_n8272<=n_n7894;

 always  @(posedge pclk)
	n_n9312<=n_n7249;

 always  @(posedge pclk)
	n_n7985<=n_n7984;

 always  @(posedge pclk)
	n_n8312<=n_n8311;

 always  @(posedge pclk)
	n_n7231<=n_n7230;

 always  @(posedge pclk)
	n_n9396<=n_n7317;

 always  @(posedge pclk)
	n_n8801<=n_n8799;

 always  @(posedge pclk)
	n_n8683<=n_n8682;

 always  @(posedge pclk)
	ndn3_39<=n_n9425;

 always  @(posedge pclk)
	n_n8245<=n_n8244;

 always  @(posedge pclk)
	n_n9458<=n_n9457;

 always  @(posedge pclk)
	n_n9302<=n_n9301;

 always  @(posedge pclk)
	n_n7392<=n_n7391;

 always  @(posedge pclk)
	n_n6963<=n_n6962;

 always  @(posedge pclk)
	n_n7808<=n_n6916;

 always  @(posedge pclk)
	n_n7225<=n_n7224;

 always  @(posedge pclk)
	n_n7817<=n_n7505;

 always  @(posedge pclk)
	n_n8201<=n_n7169;

 always  @(posedge pclk)
	n_n7793<=n_n6970;

 always  @(posedge pclk)
	n_n8177<=n_n8176;

 always  @(posedge pclk)
	n_n8389<=n_n8388;

 always  @(posedge pclk)
	n_n9440<=n_n7998;

 always  @(posedge pclk)
	n_n7683<=n_n7595;

 always  @(posedge pclk)
	n_n7761<=n_n6996;

 always  @(posedge pclk)
	n_n7667<=n_n7263;

 always  @(posedge pclk)
	n_n7980<=n_n7979;

 always  @(posedge pclk)
	n_n7509<=n_n6992;

 always  @(posedge pclk)
	n_n7813<=n_n7675;

 always  @(posedge pclk)
	n_n8396<=n_n8395;

 always  @(posedge pclk)
	n_n9535<=n_n9532;

 always  @(posedge pclk)
	n_n7209<=n_n7208;

 always  @(posedge pclk)
	n_n7003<=n_n7002;

 always  @(posedge pclk)
	n_n7695<=n_n7004;

 always  @(posedge pclk)
	n_n7624<=n_n7623;

 always  @(posedge pclk)
	n_n8791<=n_n8790;

 always  @(posedge pclk)
	n_n7374<=n_n7253;

 always  @(posedge pclk)
	n_n7429<=n_n7161;

 always  @(posedge pclk)
	n_n7944<=n_n7943;

 always  @(posedge pclk)
	n_n9266<=n_n6997;

 always  @(posedge pclk)
	n_n8100<=n_n8098;

 always  @(posedge pclk)
	n_n6988<=n_n6987;

 always  @(posedge pclk)
	n_n6986<=n_n6985;

 always  @(posedge pclk)
	n_n8933<=n_n8926;

 always  @(posedge pclk)
	n_n7117<=n_n7116;

 always  @(posedge pclk)
	n_n9043<=n_n8372;

 always  @(posedge pclk)
	n_n8241<=n_n7379;

 always  @(posedge pclk)
	n_n9219<=n_n9218;

 always  @(posedge pclk)
	n_n8198<=n_n7048;

 always  @(posedge pclk)
	n_n8081<=n_n8080;

 always  @(posedge pclk)
	n_n8575<=n_n7131;

 always  @(posedge pclk)
	n_n8710<=n_n8709;

 always  @(posedge pclk)
	n_n7622<=n_n7621;

 always  @(posedge pclk)
	n_n7966<=n_n7340;

 always  @(posedge pclk)
	n_n7885<=n_n7114;

 always  @(posedge pclk)
	n_n7033<=n_n7032;

 always  @(posedge pclk)
	ndn3_34<=n_n9088;

 always  @(posedge pclk)
	n_n9186<=n_n9185;

 always  @(posedge pclk)
	ndn3_50<=n_n8129;

 always  @(posedge pclk)
	n_n7879<=n_n7564;

 always  @(posedge pclk)
	n_n7019<=n_n7018;

 always  @(posedge pclk)
	n_n9171<=n_n8309;

 always  @(posedge pclk)
	n_n7261<=n_n7260;

 always  @(posedge pclk)
	n_n8223<=n_n7839;

 always  @(posedge pclk)
	n_n8989<=n_n7619;

 always  @(posedge pclk)
	n_n7993<=n_n7992;

 always  @(posedge pclk)
	n_n7845<=n_n7138;

 always  @(posedge pclk)
	n_n8253<=n_n8252;

 always  @(posedge pclk)
	n_n8889<=n_n8888;

 always  @(posedge pclk)
	n_n7809<=n_n7234;

 always  @(posedge pclk)
	n_n8918<=n_n8917;

 always  @(posedge pclk)
	n_n8515<=n_n7501;

 always  @(posedge pclk)
	n_n7933<=n_n7084;

 always  @(posedge pclk)
	n_n8075<=n_n8074;

 always  @(posedge pclk)
	n_n7338<=n_n7337;

 always  @(posedge pclk)
	n_n8104<=n_n8103;

 always  @(posedge pclk)
	n_n8171<=n_n8170;

 always  @(posedge pclk)
	n_n9059<=n_n9058;

 always  @(posedge pclk)
	n_n9023<=n_n9022;

 always  @(posedge pclk)
	n_n7692<=n_n7152;

 always  @(posedge pclk)
	n_n9441<=n_n8952;

 always  @(posedge pclk)
	n_n6920<=n_n6919;

 always  @(posedge pclk)
	n_n8831<=n_n8830;

 always  @(posedge pclk)
	n_n8441<=n_n8440;

 always  @(posedge pclk)
	n_n9576<=n_n8231;

 always  @(posedge pclk)
	n_n9252<=n_n9251;

 always  @(posedge pclk)
	n_n9363<=n_n7981;

 always  @(posedge pclk)
	ndn3_4<=n_n8565;

 always  @(posedge pclk)
	n_n9247<=n_n9461;

 always  @(posedge pclk)
	n_n7561<=n_n7560;

 always  @(posedge pclk)
	n_n8923<=n_n8922;

 always  @(posedge pclk)
	n_n7978<=n_n7977;

 always  @(posedge pclk)
	n_n8978<=n_n7828;

 always  @(posedge pclk)
	n_n9499<=n_n7170;

 always  @(posedge pclk)
	n_n8713<=n_n8712;

 always  @(posedge pclk)
	n_n8944<=n_n8943;

 always  @(posedge pclk)
	n_n8239<=n_n7371;

 always  @(posedge pclk)
	n_n7652<=n_n7215;

 always  @(posedge pclk)
	n_n9042<=n_n7027;

 always  @(posedge pclk)
	n_n8530<=n_n6982;

 always  @(posedge pclk)
	n_n9271<=n_n7115;

 always  @(posedge pclk)
	n_n9318<=n_n7072;

 always  @(posedge pclk)
	n_n7706<=n_n7445;

 always  @(posedge pclk)
	n_n7964<=n_n7963;

 always  @(posedge pclk)
	n_n8222<=n_n7348;

 always  @(posedge pclk)
	n_n8898<=n_n8897;

 always  @(posedge pclk)
	n_n7976<=n_n7974;

 always  @(posedge pclk)
	n_n7649<=n_n7648;

 always  @(posedge pclk)
	n_n7604<=n_n7035;

 always  @(posedge pclk)
	n_n7961<=n_n7960;

 always  @(posedge pclk)
	n_n7424<=n_n7423;

 always  @(posedge pclk)
	n_n7476<=n_n7475;

 always  @(posedge pclk)
	n_n9259<=n_n8766;

 always  @(posedge pclk)
	n_n9309<=n_n9032;

 always  @(posedge pclk)
	n_n9161<=n_n8829;

 always  @(posedge pclk)
	n_n8436<=n_n8186;

 always  @(posedge pclk)
	n_n9121<=n_n9120;

 always  @(posedge pclk)
	n_n8061<=n_n8059;

 always  @(posedge pclk)
	n_n8004<=n_n7801;

 always  @(posedge pclk)
	n_n9360<=n_n7450;

 always  @(posedge pclk)
	n_n9205<=n_n9204;

 always  @(posedge pclk)
	n_n8392<=n_n8391;

 always  @(posedge pclk)
	n_n9034<=n_n7538;

 always  @(posedge pclk)
	n_n8375<=n_n8374;

 always  @(posedge pclk)
	n_n8328<=n_n8327;

 always  @(posedge pclk)
	n_n9298<=n_n9297;

 always  @(posedge pclk)
	n_n7598<=n_n7062;

 always  @(posedge pclk)
	n_n8506<=n_n8505;

 always  @(posedge pclk)
	pdn<=n_n7729;

 always  @(posedge pclk)
	n_n7737<=n_n7226;

 always  @(posedge pclk)
	n_n7420<=n_n7419;

 always  @(posedge pclk)
	n_n9291<=n_n7957;

 always  @(posedge pclk)
	n_n7946<=n_n7945;

 always  @(posedge pclk)
	n_n8584<=n_n7662;

 always  @(posedge pclk)
	n_n9308<=n_n8254;

 always  @(posedge pclk)
	n_n9403<=n_n9037;

 always  @(posedge pclk)
	n_n7284<=n_n7282;

 always  @(posedge pclk)
	n_n9270<=n_n7082;

 always  @(posedge pclk)
	n_n7390<=n_n7388;

 always  @(posedge pclk)
	n_n9351<=n_n9001;

 always  @(posedge pclk)
	n_n6968<=n_n6967;

 always  @(posedge pclk)
	n_n8668<=n_n8451;

 always  @(posedge pclk)
	n_n9605<=n_n7044;

 always  @(posedge pclk)
	n_n7013<=n_n7012;

 always  @(posedge pclk)
	n_n9626<=n_n9625;

 always  @(posedge pclk)
	n_n8200<=n_n7132;

 always  @(posedge pclk)
	n_n9028<=n_n8645;

 always  @(posedge pclk)
	n_n8803<=n_n8802;

 always  @(posedge pclk)
	n_n9570<=n_n9569;

 always  @(posedge pclk)
	n_n8366<=n_n8365;

 always  @(posedge pclk)
	n_n9050<=n_n7104;

 always  @(posedge pclk)
	n_n8650<=n_n7785;

 always  @(posedge pclk)
	n_n8574<=n_n7006;

 always  @(posedge pclk)
	n_n7276<=n_n7275;

 always  @(posedge pclk)
	n_n9212<=n_n9211;

 always  @(posedge pclk)
	n_n8384<=n_n8382;

 always  @(posedge pclk)
	ndn3_35<=n_n9453;

 always  @(posedge pclk)
	n_n8449<=n_n8434;

 always  @(posedge pclk)
	ndn3_46<=n_n7574;

 always  @(posedge pclk)
	n_n7554<=n_n6981;

 always  @(posedge pclk)
	n_n8743<=n_n6966;

 always  @(posedge pclk)
	n_n8277<=n_n7700;

 always  @(posedge pclk)
	n_n9359<=n_n7126;

 always  @(posedge pclk)
	n_n8425<=n_n8424;

 always  @(posedge pclk)
	n_n9104<=n_n9103;

 always  @(posedge pclk)
	n_n9221<=n_n9220;

 always  @(posedge pclk)
	n_n9448<=n_n9447;

 always  @(posedge pclk)
	n_n9537<=n_n8593;

 always  @(posedge pclk)
	n_n8003<=n_n7233;

 always  @(posedge pclk)
	n_n7467<=n_n7466;

 always  @(posedge pclk)
	n_n8233<=n_n8232;

 always  @(posedge pclk)
	n_n7932<=n_n7167;

 always  @(posedge pclk)
	n_n8064<=n_n8063;

 always  @(posedge pclk)
	n_n9162<=n_n9039;

 always  @(posedge pclk)
	n_n7971<=n_n7916;

 always  @(posedge pclk)
	n_n8055<=n_n8054;

 always  @(posedge pclk)
	n_n7711<=n_n7267;

 always  @(posedge pclk)
	n_n8256<=n_n8255;

 always  @(posedge pclk)
	n_n7925<=n_n7924;

 always  @(posedge pclk)
	n_n7762<=n_n7502;

 always  @(posedge pclk)
	n_n7668<=n_n7258;

 always  @(posedge pclk)
	n_n7914<=n_n7262;

 always  @(posedge pclk)
	n_n7873<=n_n7705;

 always  @(posedge pclk)
	n_n7849<=n_n7293;

 always  @(posedge pclk)
	n_n9421<=n_n9419;

 always  @(posedge pclk)
	n_n7626<=n_n7625;

 always  @(posedge pclk)
	n_n7848<=n_n7093;

 always  @(posedge pclk)
	n_n8263<=n_n8261;

 always  @(posedge pclk)
	n_n9100<=n_n8442;

 always  @(posedge pclk)
	n_n9393<=n_n7516;

 always  @(posedge pclk)
	n_n9591<=n_n6923;

 always  @(posedge pclk)
	n_n7588<=n_n7587;

 always  @(posedge pclk)
	n_n9123<=n_n9122;

 always  @(posedge pclk)
	n_n9159<=n_n9158;

 always  @(posedge pclk)
	n_n9128<=n_n8859;

 always  @(posedge pclk)
	n_n8045<=n_n8043;

 always  @(posedge pclk)
	n_n7728<=n_n7727;

 always  @(posedge pclk)
	n_n8929<=n_n8722;

 always  @(posedge pclk)
	n_n7739<=n_n7399;

 always  @(posedge pclk)
	n_n9355<=n_n9354;

 always  @(posedge pclk)
	n_n9394<=n_n7211;

 always  @(posedge pclk)
	n_n8470<=n_n8469;

 always  @(posedge pclk)
	n_n8571<=n_n7312;

 always  @(posedge pclk)
	n_n8796<=n_n8795;

 always  @(posedge pclk)
	ndn3_36<=n_n9116;

 always  @(posedge pclk)
	n_n7990<=n_n7989;

 always  @(posedge pclk)
	n_n8781<=n_n8780;

 always  @(posedge pclk)
	n_n8817<=n_n8816;

 always  @(posedge pclk)
	n_n9160<=n_n9111;

 always  @(posedge pclk)
	n_n9092<=n_n9091;

 always  @(posedge pclk)
	n_n8513<=n_n6938;

 always  @(posedge pclk)
	n_n8213<=n_n8212;

 always  @(posedge pclk)
	n_n8581<=n_n7593;

 always  @(posedge pclk)
	n_n9284<=n_n8686;

 always  @(posedge pclk)
	n_n7837<=n_n7836;

 always  @(posedge pclk)
	n_n8224<=n_n6939;

 always  @(posedge pclk)
	n_n9203<=n_n9202;

 always  @(posedge pclk)
	n_n7655<=n_n7113;

 always  @(posedge pclk)
	n_n8946<=n_n8945;

 always  @(posedge pclk)
	n_n7052<=n_n7051;

 always  @(posedge pclk)
	n_n9615<=n_n9614;

 always  @(posedge pclk)
	n_n8473<=n_n8472;

 always  @(posedge pclk)
	n_n7741<=n_n6935;

 always  @(posedge pclk)
	n_n9460<=n_n7237;

 always  @(posedge pclk)
	n_n7912<=n_n7204;

 always  @(posedge pclk)
	n_n7606<=n_n7525;

 always  @(posedge pclk)
	n_n9021<=n_n9020;

 always  @(posedge pclk)
	n_n7781<=n_n7780;

 always  @(posedge pclk)
	n_n7810<=n_n6931;

 always  @(posedge pclk)
	n_n7108<=n_n7107;

 always  @(posedge pclk)
	n_n7697<=n_n7489;

 always  @(posedge pclk)
	n_n7642<=n_n7265;

 always  @(posedge pclk)
	n_n9595<=n_n8546;

 always  @(posedge pclk)
	n_n7694<=n_n7046;

 always  @(posedge pclk)
	n_n8221<=n_n8220;

 always  @(posedge pclk)
	n_n7600<=n_n7396;

 always  @(posedge pclk)
	n_n7935<=n_n7899;

 always  @(posedge pclk)
	n_n9230<=n_n9229;

 always  @(posedge pclk)
	n_n7701<=n_n7515;

 always  @(posedge pclk)
	n_n7510<=n_n6929;

 always  @(posedge pclk)
	n_n7627<=n_n6917;

 always  @(posedge pclk)
	n_n8502<=n_n8501;

 always  @(posedge pclk)
	n_n8516<=n_n8432;

 always  @(posedge pclk)
	n_n7913<=n_n7631;

 always  @(posedge pclk)
	n_n9320<=n_n9038;

 always  @(posedge pclk)
	n_n7411<=n_n7410;

 always  @(posedge pclk)
	n_n9129<=n_n7326;

 always  @(posedge pclk)
	n_n9053<=n_n7134;

 always  @(posedge pclk)
	n_n7069<=n_n7068;

 always  @(posedge pclk)
	n_n8617<=n_n8616;

 always  @(posedge pclk)
	n_n7242<=n_n7241;

 always  @(posedge pclk)
	n_n8230<=n_n8229;

 always  @(posedge pclk)
	n_n9294<=n_n9293;

 always  @(posedge pclk)
	n_n8249<=n_n8248;

 always  @(posedge pclk)
	n_n8972<=n_n8971;

 always  @(posedge pclk)
	n_n7074<=n_n7073;

 always  @(posedge pclk)
	n_n7493<=n_n7492;

 always  @(posedge pclk)
	n_n8290<=n_n8289;

 always  @(posedge pclk)
	n_n8821<=n_n7184;

 always  @(posedge pclk)
	n_n7769<=n_n7162;

 always  @(posedge pclk)
	n_n7491<=n_n7490;

 always  @(posedge pclk)
	n_n9600<=n_n8291;

 always  @(posedge pclk)
	n_n9317<=n_n8731;

 always  @(posedge pclk)
	n_n8047<=n_n8046;

 always  @(posedge pclk)
	n_n9629<=n_n9628;

 always  @(posedge pclk)
	n_n9126<=n_n6918;

 always  @(posedge pclk)
	n_n9508<=n_n9507;

 always  @(posedge pclk)
	n_n9155<=n_n9154;

 always  @(posedge pclk)
	n_n8528<=n_n7377;

 always  @(posedge pclk)
	ndn3_37<=n_n8994;

 always  @(posedge pclk)
	ndn3_42<=n_n7690;

 always  @(posedge pclk)
	n_n9358<=n_n7608;

 always  @(posedge pclk)
	n_n8185<=n_n8184;

 always  @(posedge pclk)
	nen3_28<=n_n7529;

 always  @(posedge pclk)
	n_n8839<=n_n8838;

 always  @(posedge pclk)
	n_n7903<=n_n7902;

 always  @(posedge pclk)
	n_n9139<=n_n9138;

 always  @(posedge pclk)
	n_n9075<=n_n9074;

 always  @(posedge pclk)
	n_n9439<=n_n7449;

 always  @(posedge pclk)
	n_n9353<=n_n6977;

 always  @(posedge pclk)
	n_n7665<=n_n7151;

 always  @(posedge pclk)
	n_n8798<=n_n7747;

 always  @(posedge pclk)
	n_n7146<=n_n7145;

 always  @(posedge pclk)
	n_n7890<=n_n7056;

 always  @(posedge pclk)
	n_n7176<=n_n7175;

 always  @(posedge pclk)
	n_n8477<=n_n8476;

 always  @(posedge pclk)
	n_n8514<=n_n8412;

 always  @(posedge pclk)
	n_n8636<=n_n8635;

 always  @(posedge pclk)
	n_n7183<=n_n7182;

 always  @(posedge pclk)
	n_n8657<=n_n8656;

 always  @(posedge pclk)
	n_n9493<=n_n8483;

 always  @(posedge pclk)
	n_n7969<=n_n6946;

 always  @(posedge pclk)
	n_n9255<=n_n7530;

 always  @(posedge pclk)
	n_n8535<=n_n8534;

 always  @(posedge pclk)
	n_n8619<=n_n8618;

 always  @(posedge pclk)
	n_n8909<=n_n8908;

 always  @(posedge pclk)
	n_n7744<=n_n7596;

 always  @(posedge pclk)
	n_n9119<=n_n9118;

 always  @(posedge pclk)
	n_n7827<=n_n7534;

 always  @(posedge pclk)
	n_n8916<=n_n8914;

 always  @(posedge pclk)
	n_n8729<=n_n8728;

 always  @(posedge pclk)
	n_n9011<=n_n8385;

 always  @(posedge pclk)
	n_n8779<=n_n8778;

 always  @(posedge pclk)
	n_n6980<=n_n6979;

 always  @(posedge pclk)
	n_n7715<=n_n7714;

 always  @(posedge pclk)
	n_n9067<=n_n9066;

 always  @(posedge pclk)
	n_n9164<=n_n7059;

 always  @(posedge pclk)
	n_n7402<=n_n7400;

 always  @(posedge pclk)
	n_n8938<=n_n7247;

 always  @(posedge pclk)
	n_n9046<=n_n8689;

 always  @(posedge pclk)
	n_n8789<=n_n8788;

 always  @(posedge pclk)
	n_n9390<=n_n8553;

 always  @(posedge pclk)
	n_n7768<=n_n7528;

 always  @(posedge pclk)
	n_n9136<=n_n7292;

 always  @(posedge pclk)
	n_n8670<=n_n8669;

 always  @(posedge pclk)
	n_n8644<=n_n8642;

 always  @(posedge pclk)
	n_n9178<=n_n6998;

 always  @(posedge pclk)
	n_n8188<=n_n8187;

 always  @(posedge pclk)
	n_n7083<=n_n7029;

 always  @(posedge pclk)
	n_n9344<=n_n9065;

 always  @(posedge pclk)
	n_n7366<=n_n7364;

 always  @(posedge pclk)
	n_n8361<=n_n8359;

 always  @(posedge pclk)
	n_n9228<=n_n9227;

 always  @(posedge pclk)
	n_n9402<=n_n8919;

 always  @(posedge pclk)
	n_n8510<=n_n8509;

 always  @(posedge pclk)
	n_n8881<=n_n8837;

 always  @(posedge pclk)
	n_n9404<=n_n8639;

 always  @(posedge pclk)
	n_n9424<=n_n9422;

 always  @(posedge pclk)
	n_n9031<=n_n8356;

 always  @(posedge pclk)
	nsr3_37<=n_n3;

 always  @(posedge pclk)
	n_n8197<=n_n7447;

 always  @(posedge pclk)
	n_n8468<=n_n8467;

 always  @(posedge pclk)
	n_n7121<=n_n7120;

 always  @(posedge pclk)
	n_n7511<=n_n7482;

 always  @(posedge pclk)
	ndn3_44<=n_n7232;

 always  @(posedge pclk)
	n_n9322<=n_n8500;

 always  @(posedge pclk)
	n_n7682<=n_n7351;

 always  @(posedge pclk)
	n_n9603<=n_n8038;

 always  @(posedge pclk)
	nlc1_2<=n_n8814;

 always  @(posedge pclk)
	n_n8408<=n_n8407;

 always  @(posedge pclk)
	n_n8577<=n_n8576;

 always  @(posedge pclk)
	n_n7079<=n_n7078;

 always  @(posedge pclk)
	n_n8828<=n_n8827;

 always  @(posedge pclk)
	n_n9340<=n_n8767;

 always  @(posedge pclk)
	n_n8586<=n_n8585;

 always  @(posedge pclk)
	n_n7901<=n_n7900;

 always  @(posedge pclk)
	n_n8628<=n_n8627;

 always  @(posedge pclk)
	n_n8869<=n_n7750;

 always  @(posedge pclk)
	n_n7710<=n_n7118;

 always  @(posedge pclk)
	n_n8993<=n_n8181;

 always  @(posedge pclk)
	n_n9586<=n_n8062;

 always  @(posedge pclk)
	n_n8852<=n_n8851;

 always  @(posedge pclk)
	n_n8583<=n_n6930;

 always  @(posedge pclk)
	n_n8011<=n_n8010;

 always  @(posedge pclk)
	n_n7717<=n_n7716;

 always  @(posedge pclk)
	n_n8326<=n_n8325;

 always  @(posedge pclk)
	n_n9163<=n_n7193;

 always  @(posedge pclk)
	n_n8344<=n_n8343;

 always  @(posedge pclk)
	n_n8296<=n_n8295;

 always  @(posedge pclk)
	n_n8116<=n_n8115;

 always  @(posedge pclk)
	n_n8267<=n_n8266;

 always  @(posedge pclk)
	n_n7686<=n_n7563;

 always  @(posedge pclk)
	n_n9061<=n_n9060;

 always  @(posedge pclk)
	n_n9338<=n_n9206;

 always  @(posedge pclk)
	n_n7688<=n_n7278;

 always  @(posedge pclk)
	n_n9081<=n_n9080;

 always  @(posedge pclk)
	n_n6910<=n_n6909;

 always  @(posedge pclk)
	n_n8727<=n_n8726;

 always  @(posedge pclk)
	n_n7674<=n_n7672;

 always  @(posedge pclk)
	n_n7330<=n_n7329;

 always  @(posedge pclk)
	n_n8966<=n_n8965;

 always  @(posedge pclk)
	n_n7843<=n_n7841;

 always  @(posedge pclk)
	n_n8847<=n_n8283;

 always  @(posedge pclk)
	n_n9376<=n_n9374;

 always  @(posedge pclk)
	n_n7553<=n_n7171;

 always  @(posedge pclk)
	n_n9292<=n_n6927;

 always  @(posedge pclk)
	n_n7464<=n_n7071;

 always  @(posedge pclk)
	n_n8146<=n_n8144;

 always  @(posedge pclk)
	n_n8439<=n_n8437;

 always  @(posedge pclk)
	n_n9498<=n_n6999;

 always  @(posedge pclk)
	n_n8118<=n_n8117;

 always  @(posedge pclk)
	n_n9452<=n_n7610;

 always  @(posedge pclk)
	n_n9239<=n_n9238;

 always  @(posedge pclk)
	n_n9237<=n_n9236;

 always  @(posedge pclk)
	n_n9488<=n_n6913;

 always  @(posedge pclk)
	ndn3_2<=n_n9443;

 always  @(posedge pclk)
	n_n9522<=n_n9521;

 always  @(posedge pclk)
	n_n9313<=n_n7518;

 always  @(posedge pclk)
	n_n7435<=n_n7433;

 always  @(posedge pclk)
	n_n8665<=n_n8664;

 always  @(posedge pclk)
	n_n9593<=n_n8318;

 always  @(posedge pclk)
	n_n8303<=n_n8301;

 always  @(posedge pclk)
	n_n7022<=n_n7020;

 always  @(posedge pclk)
	n_n9173<=n_n8133;

 always  @(posedge pclk)
	n_n9261<=n_n8896;

 always  @(posedge pclk)
	n_n7150<=n_n7149;

 always  @(posedge pclk)
	n_n9455<=n_n9454;

 always  @(posedge pclk)
	n_n8371<=n_n8370;

 always  @(posedge pclk)
	nsr3_20<=n_n8;

 always  @(posedge pclk)
	n_n8271<=n_n7047;

 always  @(posedge pclk)
	n_n9542<=n_n8836;

 always  @(posedge pclk)
	n_n7444<=n_n7443;

 always  @(posedge pclk)
	ndn3_40<=n_n7158;

 always  @(posedge pclk)
	n_n7130<=n_n7128;

 always  @(posedge pclk)
	n_n9347<=n_n7676;

 always  @(posedge pclk)
	n_n8102<=n_n8101;

 always  @(posedge pclk)
	n_n9225<=n_n9224;

 always  @(posedge pclk)
	n_n8462<=n_n8461;

 always  @(posedge pclk)
	n_n8088<=n_n8087;

 always  @(posedge pclk)
	n_n9026<=n_n9024;

 always  @(posedge pclk)
	n_n9289<=n_n8178;

 always  @(posedge pclk)
	n_n7661<=n_n7660;

 always  @(posedge pclk)
	n_n8108<=n_n8107;

 always  @(posedge pclk)
	n_n8921<=n_n8920;

 always  @(posedge pclk)
	n_n7859<=n_n7858;

 always  @(posedge pclk)
	n_n7732<=n_n7731;

 always  @(posedge pclk)
	n_n7956<=n_n7427;

 always  @(posedge pclk)
	n_n9520<=n_n9519;

 always  @(posedge pclk)
	n_n7666<=n_n6964;

 always  @(posedge pclk)
	n_n7678<=n_n7677;

 always  @(posedge pclk)
	n_n7846<=n_n7222;

 always  @(posedge pclk)
	n_n8280<=n_n7679;

 always  @(posedge pclk)
	n_n8841<=n_n8840;

 always  @(posedge pclk)
	n_n7336<=n_n7335;

 always  @(posedge pclk)
	n_n8226<=n_n7197;

 always  @(posedge pclk)
	n_n8151<=n_n7754;

 always  @(posedge pclk)
	n_n7644<=n_n7195;

 always  @(posedge pclk)
	n_n8770<=n_n8769;

 always  @(posedge pclk)
	n_n8423<=n_n8422;

 always  @(posedge pclk)
	n_n7763<=n_n7085;

 always  @(posedge pclk)
	n_n9525<=n_n9524;

 always  @(posedge pclk)
	n_n8033<=n_n8032;

 always  @(posedge pclk)
	n_n7881<=n_n7533;

 always  @(posedge pclk)
	n_n7815<=n_n7426;

 always  @(posedge pclk)
	n_n9232<=n_n9231;

 always  @(posedge pclk)
	n_n7792<=n_n7257;

 always  @(posedge pclk)
	n_n9563<=n_n9562;

 always  @(posedge pclk)
	n_n8672<=n_n8671;

 always  @(posedge pclk)
	n_n7346<=n_n7106;

 always  @(posedge pclk)
	n_n7949<=n_n7008;

 always  @(posedge pclk)
	n_n8756<=n_n8755;

 always  @(posedge pclk)
	n_n8641<=n_n8640;

 always  @(posedge pclk)
	n_n8192<=n_n8191;

 always  @(posedge pclk)
	n_n8058<=n_n8057;

 always  @(posedge pclk)
	n_n8561<=n_n7439;

 always  @(posedge pclk)
	n_n9306<=n_n9305;

 always  @(posedge pclk)
	n_n9165<=n_n6928;

 always  @(posedge pclk)
	n_n8850<=n_n8848;

 always  @(posedge pclk)
	n_n9210<=n_n9209;

 always  @(posedge pclk)
	ndn2_2<=n_n8122;

 always  @(posedge pclk)
	n_n7342<=n_n7254;

 always  @(posedge pclk)
	n_n8051<=n_n8050;

 always  @(posedge pclk)
	n_n7136<=n_n7135;

 always  @(posedge pclk)
	n_n9348<=n_n7081;

 always  @(posedge pclk)
	n_n9006<=n_n9005;

 always  @(posedge pclk)
	n_n7653<=n_n7407;

 always  @(posedge pclk)
	n_n7905<=n_n7904;

 always  @(posedge pclk)
	n_n9166<=n_n7030;

 always  @(posedge pclk)
	n_n7065<=n_n7064;

 always  @(posedge pclk)
	n_n9490<=n_n8211;

 always  @(posedge pclk)
	n_n7024<=n_n7023;

 always  @(posedge pclk)
	n_n7586<=n_n7585;

 always  @(posedge pclk)
	n_n8416<=n_n8415;

 always  @(posedge pclk)
	n_n8937<=n_n8166;

 always  @(posedge pclk)
	n_n8141<=n_n8140;

 always  @(posedge pclk)
	n_n7853<=n_n7446;

 always  @(posedge pclk)
	n_n8121<=n_n8120;

 always  @(posedge pclk)
	n_n9604<=n_n8162;

 always  @(posedge pclk)
	n_n9496<=n_n8337;

 always  @(posedge pclk)
	n_n8195<=n_n8194;

 always  @(posedge pclk)
	n_n9516<=n_n9515;

 always  @(posedge pclk)
	n_n9077<=n_n9076;

 always  @(posedge pclk)
	n_n9436<=n_n8363;

 always  @(posedge pclk)
	n_n9051<=n_n8773;

 always  @(posedge pclk)
	n_n7664<=n_n7089;

 always  @(posedge pclk)
	n_n8419<=n_n7840;

 always  @(posedge pclk)
	n_n7874<=n_n7321;

 always  @(posedge pclk)
	n_n9133<=n_n8873;

 always  @(posedge pclk)
	n_n9392<=n_n7745;

 always  @(posedge pclk)
	n_n7770<=n_n7001;

 always  @(posedge pclk)
	ndn3_32<=n_n6959;

 always  @(posedge pclk)
	n_n7601<=n_n7196;

 always  @(posedge pclk)
	n_n8206<=n_n8205;

 always  @(posedge pclk)
	n_n7927<=n_n7367;

 always  @(posedge pclk)
	n_n9606<=n_n8818;

 always  @(posedge pclk)
	n_n7111<=n_n7110;

 always  @(posedge pclk)
	n_n9269<=n_n7804;

 always  @(posedge pclk)
	ndn3_38<=n_n8494;

 always  @(posedge pclk)
	n_n7886<=n_n7206;

 always  @(posedge pclk)
	n_n9179<=n_n8872;

 always  @(posedge pclk)
	n_n9357<=n_n8364;

 always  @(posedge pclk)
	n_n9594<=n_n8496;

 always  @(posedge pclk)
	n_n7628<=n_n6971;

 always  @(posedge pclk)
	n_n8454<=n_n8453;

 always  @(posedge pclk)
	ndn3_20<=n_n7413;

 always  @(posedge pclk)
	n_n9505<=n_n9504;

 always  @(posedge pclk)
	nen3_34<=n_n8825;

 always  @(posedge pclk)
	n_n9632<=n_n9631;

 always  @(posedge pclk)
	n_n7076<=n_n7075;

 always  @(posedge pclk)
	n_n9262<=n_n7469;

 always  @(posedge pclk)
	n_n9048<=n_n8634;

 always  @(posedge pclk)
	n_n9578<=n_n9577;

 always  @(posedge pclk)
	n_n8135<=n_n8134;

 always  @(posedge pclk)
	ndn3_26<=n_n9328;

 always  @(posedge pclk)
	n_n7500<=n_n7499;

 always  @(posedge pclk)
	n_n6974<=n_n6973;

 always  @(posedge pclk)
	n_n8605<=n_n8604;

 always  @(posedge pclk)
	n_n9296<=n_n9295;

 always  @(posedge pclk)
	n_n7156<=n_n7155;

 always  @(posedge pclk)
	n_n7920<=n_n7919;

 always  @(posedge pclk)
	n_n8895<=n_n8893;

 always  @(posedge pclk)
	n_n8991<=n_n7620;

 always  @(posedge pclk)
	n_n8139<=n_n8138;

 always  @(posedge pclk)
	n_n9275<=n_n9274;

 always  @(posedge pclk)
	n_n7203<=n_n7202;

 always  @(posedge pclk)
	n_n9590<=n_n7805;

 always  @(posedge pclk)
	n_n7344<=n_n7343;

 always  @(posedge pclk)
	n_n6976<=n_n6975;

 always  @(posedge pclk)
	n_n7629<=n_n6958;

 always  @(posedge pclk)
	ndn3_14<=n_n7617;

 always  @(posedge pclk)
	n_n7862<=n_n7646;

 always  @(posedge pclk)
	n_n9013<=n_n9012;

 always  @(posedge pclk)
	n_n7288<=n_n7287;

 always  @(posedge pclk)
	n_n8078<=n_n8077;

 always  @(posedge pclk)
	n_n7334<=n_n7333;

 always  @(posedge pclk)
	n_n7704<=n_n6957;

 always  @(posedge pclk)
	n_n7788<=n_n7496;

 always  @(posedge pclk)
	n_n8526<=n_n8525;

 always  @(posedge pclk)
	n_n9556<=n_n7795;

 always  @(posedge pclk)
	n_n9345<=n_n7851;

 always  @(posedge pclk)
	n_n8447<=n_n8446;

 always  @(posedge pclk)
	n_n7485<=n_n7484;

 always  @(posedge pclk)
	n_n8570<=n_n7305;

 always  @(posedge pclk)
	n_n7453<=n_n6921;

 always  @(posedge pclk)
	n_n7928<=n_n7191;

 always  @(posedge pclk)
	n_n8646<=n_n6926;

 always  @(posedge pclk)
	n_n9405<=n_n8489;

 always  @(posedge pclk)
	n_n8948<=n_n8947;

 always  @(posedge pclk)
	n_n9131<=n_n8471;

 always  @(posedge pclk)
	n_n8216<=n_n8215;

 always  @(posedge pclk)
	n_n9177<=n_n8180;

 always  @(posedge pclk)
	n_n7844<=n_n7295;

 always  @(posedge pclk)
	n_n8811<=n_n7437;

 always  @(posedge pclk)
	n_n9145<=n_n9143;

 always  @(posedge pclk)
	n_n8428<=n_n8426;

 always  @(posedge pclk)
	n_n8858<=n_n8558;

 always  @(posedge pclk)
	n_n8580<=n_n7838;

 assign psv39_8_8_ = ( n_n9366  &  n_n7154 ) | ( tin_psv39_8_8_  &  (~ n_n7154) ) ;
 assign psv39_0_0_ = ( tin_psv39_0_0_  &  (~ n_n6986) ) | ( n_n6986  &  n_n9424 ) ;
 assign psv13_5_5_ = ( n_n9004  &  n_n7561 ) | ( tin_psv13_5_5_  &  (~ n_n7561) ) ;
 assign psv2_13_13_ = ( n_n9169  &  n_n8245 ) | ( tin_psv2_13_13_  &  (~ n_n8245) ) ;
 assign psv2_8_8_ = ( n_n8303  &  n_n8121 ) | ( tin_psv2_8_8_  &  (~ n_n8121) ) ;
 assign psv38_2_2_ = ( tin_psv38_2_2_  &  (~ n_n7146) ) | ( n_n7146  &  n_n6910 ) ;
 assign psv33_5_5_ = ( n_n9148  &  n_n7050 ) | ( tin_psv33_5_5_  &  (~ n_n7050) ) ;
 assign psv26_6_6_ = ( tin_psv26_6_6_  &  (~ n_n7622) ) | ( n_n7622  &  n_n6980 ) ;
 assign psv2_9_9_ = ( n_n7522  &  n_n8918 ) | ( tin_psv2_9_9_  &  (~ n_n8918) ) ;
 assign psv18_2_2_ = ( n_n8801  &  n_n7905 ) | ( tin_psv18_2_2_  &  (~ n_n7905) ) ;
 assign psv39_9_9_ = ( n_n7332  &  n_n7717 ) | ( tin_psv39_9_9_  &  (~ n_n7717) ) ;
 assign psv39_1_1_ = ( n_n8430  &  n_n8946 ) | ( tin_psv39_1_1_  &  (~ n_n8946) ) ;
 assign psv13_6_6_ = ( n_n7179  &  n_n8568 ) | ( tin_psv13_6_6_  &  (~ n_n8568) ) ;
 assign psv2_6_6_ = ( n_n7022  &  n_n7150 ) | ( tin_psv2_6_6_  &  (~ n_n7150) ) ;
 assign psv38_3_3_ = ( tin_psv38_3_3_  &  (~ n_n7491) ) | ( n_n7491  &  n_n7203 ) ;
 assign psv33_6_6_ = ( tin_psv33_6_6_  &  (~ n_n8243) ) | ( n_n8243  &  n_n7344 ) ;
 assign psv26_13_13_ = ( tin_psv26_13_13_  &  (~ n_n7381) ) | ( n_n7381  &  n_n7500 ) ;
 assign psv26_12_12_ = ( n_n8488  &  n_n7798 ) | ( tin_psv26_12_12_  &  (~ n_n7798) ) ;
 assign psv26_7_7_ = ( n_n8702  &  n_n7362 ) | ( tin_psv26_7_7_  &  (~ n_n7362) ) ;
 assign psv2_7_7_ = ( n_n8061  &  n_n8392 ) | ( tin_psv2_7_7_  &  (~ n_n8392) ) ;
 assign psv18_3_3_ = ( n_n7498  &  n_n7079 ) | ( tin_psv18_3_3_  &  (~ n_n7079) ) ;
 assign psv39_2_2_ = ( n_n7726  &  n_n7978 ) | ( tin_psv39_2_2_  &  (~ n_n7978) ) ;
 assign psv33_12_12_ = ( n_n8369  &  n_n7493 ) | ( tin_psv33_12_12_  &  (~ n_n7493) ) ;
 assign psv33_11_11_ = ( n_n7923  &  n_n8665 ) | ( tin_psv33_11_11_  &  (~ n_n8665) ) ;
 assign psv33_10_10_ = ( n_n9483  &  n_n9123 ) | ( tin_psv33_10_10_  &  (~ n_n9123) ) ;
 assign psv13_7_7_ = ( n_n7546  &  n_n9228 ) | ( tin_psv13_7_7_  &  (~ n_n9228) ) ;
 assign psv2_10_10_ = ( tin_psv2_10_10_  &  (~ n_n7244) ) | ( n_n7244  &  n_n8681 ) ;
 assign psv38_4_4_ = ( tin_psv38_4_4_  &  (~ n_n7052) ) | ( n_n7052  &  n_n7674 ) ;
 assign psv39_10_10_ = ( n_n8644  &  n_n7330 ) | ( tin_psv39_10_10_  &  (~ n_n7330) ) ;
 assign psv33_7_7_ = ( tin_psv33_7_7_  &  (~ n_n7140) ) | ( n_n7140  &  n_n7843 ) ;
 assign psv26_15_15_ = ( tin_psv26_15_15_  &  (~ n_n8389) ) | ( n_n8389  &  n_n9026 ) ;
 assign psv26_14_14_ = ( tin_psv26_14_14_  &  (~ n_n9200) ) | ( n_n9200  &  n_n7392 ) ;
 assign psv26_8_8_ = ( n_n7581  &  n_n6937 ) | ( tin_psv26_8_8_  &  (~ n_n6937) ) ;
 assign psv26_0_0_ = ( n_n7017  &  n_n7246 ) | ( tin_psv26_0_0_  &  (~ n_n7246) ) ;
 assign psv13_12_12_ = ( tin_psv13_12_12_  &  (~ n_n8055) ) | ( n_n8055  &  n_n8895 ) ;
 assign psv13_11_11_ = ( n_n9548  &  n_n7336 ) | ( tin_psv13_11_11_  &  (~ n_n7336) ) ;
 assign psv18_4_4_ = ( n_n9432  &  n_n9006 ) | ( tin_psv18_4_4_  &  (~ n_n9006) ) ;
 assign psv39_3_3_ = ( tin_psv39_3_3_  &  (~ n_n7507) ) | ( n_n7507  &  n_n7108 ) ;
 assign psv13_8_8_ = ( n_n7271  &  n_n7261 ) | ( tin_psv13_8_8_  &  (~ n_n7261) ) ;
 assign psv13_0_0_ = ( n_n7775  &  n_n7176 ) | ( tin_psv13_0_0_  &  (~ n_n7176) ) ;
 assign psv38_5_5_ = ( tin_psv38_5_5_  &  (~ n_n8655) ) | ( n_n8655  &  n_n7256 ) ;
 assign psv33_8_8_ = ( tin_psv33_8_8_  &  (~ n_n9306) ) | ( n_n9306  &  n_n7288 ) ;
 assign psv33_0_0_ = ( n_n8486  &  n_n8672 ) | ( tin_psv33_0_0_  &  (~ n_n8672) ) ;
 assign psv26_9_9_ = ( tin_psv26_9_9_  &  (~ n_n7310) ) | ( n_n7310  &  n_n7360 ) ;
 assign psv26_1_1_ = ( tin_psv26_1_1_  &  (~ n_n7699) ) | ( n_n7699  &  n_n7231 ) ;
 assign psv13_10_10_ = ( tin_psv13_10_10_  &  (~ n_n6956) ) | ( n_n6956  &  n_n7976 ) ;
 assign psv18_5_5_ = ( tin_psv18_5_5_  &  (~ n_n7903) ) | ( n_n7903  &  n_n7715 ) ;
 assign psv39_4_4_ = ( tin_psv39_4_4_  &  (~ n_n7117) ) | ( n_n7117  &  n_n7121 ) ;
 assign psv13_9_9_ = ( tin_psv13_9_9_  &  (~ n_n7944) ) | ( n_n7944  &  n_n9376 ) ;
 assign psv13_1_1_ = ( n_n8589  &  n_n7013 ) | ( tin_psv13_1_1_  &  (~ n_n7013) ) ;
 assign psv2_15_15_ = ( tin_psv2_15_15_  &  (~ n_n6948) ) | ( n_n6948  &  n_n8102 ) ;
 assign psv2_11_11_ = ( tin_psv2_11_11_  &  (~ n_n6952) ) | ( n_n6952  &  n_n6963 ) ;
 assign psv2_0_0_ = ( n_n8371  &  n_n7024 ) | ( tin_psv2_0_0_  &  (~ n_n7024) ) ;
 assign psv38_14_14_ = ( n_n7174  &  n_n8454 ) | ( tin_psv38_14_14_  &  (~ n_n8454) ) ;
 assign psv38_12_12_ = ( n_n7402  &  n_n8605 ) | ( tin_psv38_12_12_  &  (~ n_n8605) ) ;
 assign psv38_10_10_ = ( tin_psv38_10_10_  &  (~ n_n7181) ) | ( n_n7181  &  n_n7284 ) ;
 assign psv38_6_6_ = ( tin_psv38_6_6_  &  (~ n_n7556) ) | ( n_n7556  &  n_n7514 ) ;
 assign psv18_15_15_ = ( tin_psv18_15_15_  &  (~ n_n7019) ) | ( n_n7019  &  n_n7074 ) ;
 assign psv18_13_13_ = ( n_n7148  &  n_n7415 ) | ( tin_psv18_13_13_  &  (~ n_n7415) ) ;
 assign psv18_11_11_ = ( n_n8439  &  n_n8195 ) | ( tin_psv18_11_11_  &  (~ n_n8195) ) ;
 assign psv33_9_9_ = ( tin_psv33_9_9_  &  (~ n_n8725) ) | ( n_n8725  &  n_n9278 ) ;
 assign psv33_1_1_ = ( n_n8091  &  n_n7635 ) | ( tin_psv33_1_1_  &  (~ n_n7635) ) ;
 assign psv26_2_2_ = ( n_n7777  &  n_n7276 ) | ( tin_psv26_2_2_  &  (~ n_n7276) ) ;
 assign psv2_1_1_ = ( tin_psv2_1_1_  &  (~ n_n7467) ) | ( n_n7467  &  n_n7678 ) ;
 assign psv38_15_15_ = ( n_n8340  &  n_n8216 ) | ( tin_psv38_15_15_  &  (~ n_n8216) ) ;
 assign psv38_11_11_ = ( n_n7857  &  n_n7033 ) | ( tin_psv38_11_11_  &  (~ n_n7033) ) ;
 assign psv18_12_12_ = ( n_n9465  &  n_n8817 ) | ( tin_psv18_12_12_  &  (~ n_n8817) ) ;
 assign psv18_6_6_ = ( tin_psv18_6_6_  &  (~ n_n8230) ) | ( n_n8230  &  n_n7156 ) ;
 assign psv39_5_5_ = ( n_n8777  &  n_n8633 ) | ( tin_psv39_5_5_  &  (~ n_n8633) ) ;
 assign psv13_2_2_ = ( tin_psv13_2_2_  &  (~ n_n8251) ) | ( n_n8251  &  n_n7130 ) ;
 assign psv38_7_7_ = ( n_n8592  &  n_n8713 ) | ( tin_psv38_7_7_  &  (~ n_n8713) ) ;
 assign psv39_12_12_ = ( tin_psv39_12_12_  &  (~ n_n9476) ) | ( n_n9476  &  n_n8100 ) ;
 assign psv39_11_11_ = ( tin_psv39_11_11_  &  (~ n_n7315) ) | ( n_n7315  &  n_n7390 ) ;
 assign psv33_2_2_ = ( tin_psv33_2_2_  &  (~ n_n7209) ) | ( n_n7209  &  n_n7111 ) ;
 assign psv26_3_3_ = ( tin_psv26_3_3_  &  (~ n_n7338) ) | ( n_n7338  &  n_n8384 ) ;
 assign psv13_14_14_ = ( n_n7252  &  n_n7959 ) | ( tin_psv13_14_14_  &  (~ n_n7959) ) ;
 assign psv13_13_13_ = ( n_n6991  &  n_n8704 ) | ( tin_psv13_13_13_  &  (~ n_n8704) ) ;
 assign psv18_10_10_ = ( tin_psv18_10_10_  &  (~ n_n8974) ) | ( n_n8974  &  n_n8146 ) ;
 assign psv18_7_7_ = ( n_n8049  &  n_n7659 ) | ( tin_psv18_7_7_  &  (~ n_n7659) ) ;
 assign psv39_6_6_ = ( n_n8073  &  n_n8047 ) | ( tin_psv39_6_6_  &  (~ n_n8047) ) ;
 assign psv33_15_15_ = ( tin_psv33_15_15_  &  (~ n_n7026) ) | ( n_n7026  &  n_n8263 ) ;
 assign psv33_14_14_ = ( n_n9429  &  n_n6988 ) | ( tin_psv33_14_14_  &  (~ n_n6988) ) ;
 assign psv33_13_13_ = ( n_n7069  &  n_n8290 ) | ( tin_psv33_13_13_  &  (~ n_n8290) ) ;
 assign psv13_3_3_ = ( n_n8850  &  n_n7586 ) | ( tin_psv13_3_3_  &  (~ n_n7586) ) ;
 assign psv2_14_14_ = ( n_n7102  &  n_n8683 ) | ( tin_psv2_14_14_  &  (~ n_n8683) ) ;
 assign psv2_12_12_ = ( n_n8132  &  n_n7286 ) | ( tin_psv2_12_12_  &  (~ n_n7286) ) ;
 assign psv2_4_4_ = ( tin_psv2_4_4_  &  (~ n_n7291) ) | ( n_n7291  &  n_n8045 ) ;
 assign psv38_8_8_ = ( tin_psv38_8_8_  &  (~ n_n6984) ) | ( n_n6984  &  n_n9421 ) ;
 assign psv38_0_0_ = ( n_n8916  &  n_n8921 ) | ( tin_psv38_0_0_  &  (~ n_n8921) ) ;
 assign psv39_14_14_ = ( n_n9371  &  n_n8441 ) | ( tin_psv39_14_14_  &  (~ n_n8441) ) ;
 assign psv39_13_13_ = ( tin_psv39_13_13_  &  (~ n_n8831) ) | ( n_n8831  &  n_n7366 ) ;
 assign psv33_3_3_ = ( tin_psv33_3_3_  &  (~ n_n7409) ) | ( n_n7409  &  n_n7420 ) ;
 assign psv26_11_11_ = ( tin_psv26_11_11_  &  (~ n_n7308) ) | ( n_n7308  &  n_n8185 ) ;
 assign psv26_10_10_ = ( tin_psv26_10_10_  &  (~ n_n9580) ) | ( n_n9580  &  n_n8781 ) ;
 assign psv26_4_4_ = ( n_n8175  &  n_n8112 ) | ( tin_psv26_4_4_  &  (~ n_n8112) ) ;
 assign psv13_15_15_ = ( tin_psv13_15_15_  &  (~ n_n8406) ) | ( n_n8406  &  n_n9145 ) ;
 assign psv2_5_5_ = ( tin_psv2_5_5_  &  (~ n_n9446) ) | ( n_n9446  &  n_n7395 ) ;
 assign psv18_8_8_ = ( n_n8678  &  n_n7242 ) | ( tin_psv18_8_8_  &  (~ n_n7242) ) ;
 assign psv18_0_0_ = ( n_n7190  &  n_n7065 ) | ( tin_psv18_0_0_  &  (~ n_n7065) ) ;
 assign psv39_7_7_ = ( n_n7160  &  n_n7183 ) | ( tin_psv39_7_7_  &  (~ n_n7183) ) ;
 assign psv13_4_4_ = ( tin_psv13_4_4_  &  (~ n_n9085) ) | ( n_n9085  &  n_n9096 ) ;
 assign psv2_2_2_ = ( n_n7054  &  n_n8510 ) | ( tin_psv2_2_2_  &  (~ n_n8510) ) ;
 assign psv38_9_9_ = ( tin_psv38_9_9_  &  (~ n_n8944) ) | ( n_n8944  &  n_n8428 ) ;
 assign psv38_1_1_ = ( tin_psv38_1_1_  &  (~ n_n9373) ) | ( n_n9373  &  n_n7964 ) ;
 assign psv39_15_15_ = ( tin_psv39_15_15_  &  (~ n_n7411) ) | ( n_n7411  &  n_n8361 ) ;
 assign psv33_4_4_ = ( n_n7462  &  n_n7003 ) | ( tin_psv33_4_4_  &  (~ n_n7003) ) ;
 assign psv26_5_5_ = ( tin_psv26_5_5_  &  (~ n_n8423) ) | ( n_n8423  &  n_n7076 ) ;
 assign psv2_3_3_ = ( n_n8750  &  n_n6912 ) | ( tin_psv2_3_3_  &  (~ n_n6912) ) ;
 assign psv38_13_13_ = ( tin_psv38_13_13_  &  (~ n_n9531) ) | ( n_n9531  &  n_n6920 ) ;
 assign psv18_14_14_ = ( tin_psv18_14_14_  &  (~ n_n8762) ) | ( n_n8762  &  n_n7435 ) ;
 assign psv18_9_9_ = ( tin_psv18_9_9_  &  (~ n_n6950) ) | ( n_n6950  &  n_n6961 ) ;
 assign psv18_1_1_ = ( tin_psv18_1_1_  &  (~ n_n7387) ) | ( n_n7387  &  n_n9535 ) ;
 assign n_n9279 = ( (~ preset)  &  n_n9280  &  (~ nrq2_9) ) ;
 assign n_n8265 = ( wire5575 ) | ( n_n9434  &  wire2421  &  n_n9639 ) ;
 assign n_n8264 = ( wire5573 ) | ( n_n9537  &  wire2421  &  n_n9639 ) ;
 assign n_n7724 = ( wire5571 ) | ( wire5572 ) ;
 assign n_n8190 = ( (~ preset)  &  n_n8270  &  (~ nrq2_9) ) ;
 assign n_n7893 = ( (~ preset)  &  n_n8196  &  (~ nrq2_9) ) ;
 assign n_n9149 = ( (~ preset)  &  n_n9150  &  (~ nrq2_9) ) ;
 assign n_n7216 = ( wire5245 ) | ( wire5246 ) ;
 assign n_n7778 = ( wire5077 ) | ( n_n7098  &  n_n9616 ) ;
 assign n_n8834 = ( wire5071 ) | ( wire5072 ) ;
 assign n_n8149 = ( wire5026 ) | ( wire5027 ) ;
 assign n_n7034 = ( wire5022 ) | ( ndn3_11  &  (~ ndn3_12)  &  wire2405 ) ;
 assign n_n7166 = ( (~ preset)  &  n_n7341  &  (~ ndn_latch3_26) ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9627 ) ;
 assign n_n7868 = ( (~ preset)  &  n_n9180  &  (~ nrq3_9) ) | ( (~ preset)  &  nrq3_9  &  n_n9581 ) ;
 assign n_n8590 = ( wire5012 ) | ( wire5013 ) ;
 assign n_n8870 = ( wire5010 ) | ( nen3_39  &  (~ ndn3_39)  &  wire2408 ) ;
 assign n_n7251 = ( wire5008 ) | ( wire5009 ) ;
 assign n_n7269 = ( wire5006 ) | ( wire5007 ) ;
 assign n_n6990 = ( wire5004 ) | ( wire5005 ) ;
 assign n_n7671 = ( wire4861 ) | ( (~ wire2453)  &  wire16550 ) | ( wire2453  &  wire16551 ) ;
 assign n_n7412 = ( wire4857 ) | ( n_n8354  &  wire2421  &  n_n9639 ) ;
 assign n_n7201 = ( (~ preset)  &  n_n7552  &  (~ ndn_latch3_27) ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9564 ) ;
 assign n_n7524 = ( (~ preset)  &  (~ nsr3_23) ) ;
 assign n_n9545 = ( wire4851 ) | ( wire4852 ) ;
 assign n_n9466 = ( wire4847 ) | ( wire4848 ) ;
 assign n_n7205 = ( wire4843 ) | ( wire4844 ) ;
 assign n_n6949 = ( (~ preset)  &  n_n6950 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7077 = ( n_n8930  &  (~ wire2469) ) | ( (~ wire2469)  &  n_n9639  &  wire16469 ) ;
 assign n_n7243 = ( (~ preset)  &  n_n7244 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n7369 = ( wire4833 ) | ( n_n9512  &  wire2436  &  n_n9639 ) ;
 assign n_n8189 = ( (~ preset)  &  n_n8883  &  (~ nrq3_19) ) | ( (~ preset)  &  nrq3_19  &  n_n9581 ) ;
 assign n_n7123 = ( wire4827 ) | ( wire4828 ) ;
 assign n_n9579 = ( (~ preset)  &  n_n9580 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n6944 = ( wire4823 ) | ( n_n9353  &  wire2447  &  n_n9639 ) ;
 assign n_n6994 = ( wire4821 ) | ( wire2368  &  n_n9581 ) ;
 assign n_n9234 = ( wire4819 ) | ( wire2370  &  (~ n_n8019)  &  n_n7573 ) | ( wire2370  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n7521 = ( wire4817 ) | ( wire4818 ) ;
 assign n_n7229 = ( (~ preset)  &  n_n7373  &  (~ ndn_latch3_29) ) | ( (~ preset)  &  ndn_latch3_29  &  n_n9564 ) ;
 assign n_n9084 = ( (~ preset)  &  n_n9085 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7416 = ( wire4809 ) | ( wire4810 ) | ( wire4811 ) | ( wire4812 ) ;
 assign n_n7066 = ( wire4805 ) | ( (~ ndn3_29)  &  ndn3_28  &  wire2402 ) ;
 assign n_n8774 = ( wire4760 ) | ( wire4761 ) ;
 assign n_n7438 = ( (~ preset)  &  n_n7654  &  (~ nrq3_16) ) | ( (~ preset)  &  nrq3_16  &  n_n9627 ) ;
 assign n_n8409 = ( (~ preset)  &  n_n8410  &  (~ nrq3_36) ) | ( (~ preset)  &  nrq3_36  &  n_n9619 ) ;
 assign n_n8207 = ( wire4668 ) | ( ndn3_17  &  (~ ndn3_18)  &  wire2404 ) ;
 assign n_n8376 = ( wire4666 ) | ( (~ ndn3_7)  &  ndn3_4  &  wire2402 ) ;
 assign n_n7028 = ( wire4664 ) | ( wire4665 ) ;
 assign n_n7421 = ( wire4662 ) | ( n_n9512  &  wire2421  &  n_n9639 ) ;
 assign n_n7753 = ( wire4660 ) | ( (~ ndn3_19)  &  nen3_19  &  wire2408 ) ;
 assign n_n7680 = ( (~ preset)  &  n_n9616  &  nrq3_19 ) | ( (~ preset)  &  n_n8202  &  (~ nrq3_19) ) ;
 assign n_n7669 = ( (~ preset)  &  n_n7670  &  (~ ndn_latch3_32) ) | ( (~ preset)  &  ndn_latch3_32  &  n_n9627 ) ;
 assign n_n7455 = ( wire4654 ) | ( wire4655 ) ;
 assign n_n6989 = ( wire4652 ) | ( wire4653 ) ;
 assign n_n8596 = ( wire4650 ) | ( wire4651 ) ;
 assign n_n7472 = ( wire4648 ) | ( wire4649 ) ;
 assign n_n8393 = ( wire4646 ) | ( n_n8449  &  wire2431  &  n_n9639 ) ;
 assign n_n7591 = ( wire4644 ) | ( n_n8419  &  wire2431  &  n_n9639 ) ;
 assign n_n7481 = ( wire4640 ) | ( wire4641 ) ;
 assign n_n9140 = ( (~ preset)  &  n_n9141  &  (~ ndn_latch3_12) ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9564 ) ;
 assign n_n7331 = ( wire4636 ) | ( wire4637 ) ;
 assign n_n8757 = ( wire4634 ) | ( wire4635 ) ;
 assign n_n7422 = ( wire4630 ) | ( wire4631 ) ;
 assign n_n7040 = ( wire4628 ) | ( ndn3_11  &  (~ ndn3_12)  &  wire2402 ) ;
 assign n_n7277 = ( wire4624 ) | ( wire4625 ) ;
 assign n_n9007 = ( wire4620 ) | ( wire4621 ) ;
 assign n_n7580 = ( wire4618 ) | ( wire4619 ) ;
 assign n_n7067 = ( (~ preset)  &  n_n7376  &  (~ nrq3_39) ) | ( (~ preset)  &  nrq3_39  &  n_n9564 ) ;
 assign n_n7092 = ( wire4614 ) | ( ndn3_9  &  (~ ndn3_11)  &  wire2404 ) ;
 assign n_n7199 = ( n_n7729  &  n_n7378 ) | ( (~ preset)  &  pover_0_0_  &  (~ n_n7378) ) ;
 assign n_n8598 = ( (~ preset)  &  n_n8599  &  (~ nrq3_18) ) | ( (~ preset)  &  nrq3_18  &  n_n9619 ) ;
 assign n_n7240 = ( wire4606 ) | ( ndn3_11  &  (~ ndn3_12)  &  wire2408 ) ;
 assign n_n7382 = ( (~ preset)  &  n_n9442  &  (~ nrq2_9) ) ;
 assign n_n8411 = ( (~ preset)  &  n_n9485  &  (~ nrq3_34) ) | ( (~ preset)  &  nrq3_34  &  n_n9581 ) ;
 assign n_n7147 = ( wire4602 ) | ( wire4603 ) ;
 assign n_n7517 = ( wire4600 ) | ( n_n9284  &  wire2436  &  n_n9639 ) ;
 assign n_n9250 = ( wire4598 ) | ( ndn3_19  &  (~ ndn3_21)  &  wire2402 ) ;
 assign n_n7188 = ( (~ preset)  &  ndn3_9  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_7 ) ;
 assign n_n8612 = ( (~ preset)  &  n_n8613  &  (~ nrq2_9) ) ;
 assign n_n8532 = ( wire4594 ) | ( n_n8707  &  wire2447  &  n_n9639 ) ;
 assign n_n8698 = ( wire4592 ) | ( n_n9512  &  wire2418  &  n_n9639 ) ;
 assign n_n8608 = ( wire4590 ) | ( wire4591 ) ;
 assign n_n8307 = ( wire4588 ) | ( wire2370  &  n_n9619 ) ;
 assign n_n8654 = ( (~ preset)  &  n_n8655 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7125 = ( wire4582 ) | ( (~ ndn3_29)  &  ndn3_28  &  wire2406 ) ;
 assign n_n7357 = ( (~ preset)  &  n_n7583  &  (~ nrq2_9) ) ;
 assign n_n7 = ( wire16674 ) | ( n_n9248  &  (~ n_n9247) ) | ( n_n9248  &  (~ n_n9246) ) ;
 assign n_n8787 = ( wire4548 ) | ( wire4549 ) ;
 assign n_n8785 = ( wire4546 ) | ( (~ ndn3_7)  &  ndn3_4  &  wire2406 ) ;
 assign n_n7473 = ( wire4544 ) | ( wire4545 ) ;
 assign n_n7214 = ( (~ preset)  &  n_n7738  &  (~ ndn_latch3_25) ) | ( (~ preset)  &  ndn_latch3_25  &  n_n9564 ) ;
 assign n_n7063 = ( (~ preset)  &  n_n8573  &  (~ nrq2_9) ) ;
 assign n_n9472 = ( (~ preset)  &  n_n9581  &  ndn_latch3_32 ) | ( (~ preset)  &  n_n9473  &  (~ ndn_latch3_32) ) ;
 assign n_n8999 = ( wire4538 ) | ( (~ ndn3_25)  &  ndn3_22  &  wire2402 ) ;
 assign n_n7495 = ( wire4536 ) | ( n_n8557  &  wire2423  &  n_n9639 ) ;
 assign n_n7266 = ( (~ preset)  &  n_n9554  &  (~ nrq2_9) ) ;
 assign n_n8507 = ( (~ preset)  &  n_n8508  &  (~ nrq2_9) ) ;
 assign n_n9634 = ( wire4534 ) | ( wire4535 ) ;
 assign n_n7189 = ( wire4532 ) | ( wire4533 ) ;
 assign n_n8700 = ( wire4530 ) | ( wire4531 ) ;
 assign n_n9105 = ( wire4526 ) | ( wire4527 ) ;
 assign n_n7408 = ( (~ preset)  &  n_n7409 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7137 = ( (~ preset)  &  n_n9437  &  (~ nrq2_9) ) ;
 assign n_n7504 = ( wire4522 ) | ( wire4523 ) ;
 assign n_n8527 = ( (~ preset)  &  n_n8647  &  (~ nrq2_9) ) ;
 assign n_n9208 = ( wire4520 ) | ( wire4521 ) ;
 assign n_n7177 = ( wire4518 ) | ( wire4519 ) ;
 assign n_n7615 = ( (~ preset)  &  (~ nsr3_13) ) ;
 assign n_n7087 = ( (~ preset)  &  ndn3_17  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_16 ) ;
 assign n_n8293 = ( (~ preset)  &  ndn3_25  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_22 ) ;
 assign n_n8217 = ( (~ preset)  &  ndn3_29  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_28 ) ;
 assign n_n9538 = ( (~ preset)  &  n_n9539  &  (~ nrq2_9) ) ;
 assign n_n7091 = ( wire4510 ) | ( n_n8821  &  wire2431  &  n_n9639 ) ;
 assign n_n8487 = ( wire4508 ) | ( wire4509 ) ;
 assign n_n8299 = ( (~ preset)  &  nen3_22  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_23) ) ;
 assign n_n7796 = ( (~ preset)  &  n_n9438  &  (~ nrq2_9) ) ;
 assign n_n8130 = ( wire4504 ) | ( wire4505 ) ;
 assign n_n8660 = ( wire4502 ) | ( n_n9416  &  wire2427  &  n_n9639 ) ;
 assign n_n7325 = ( wire4498 ) | ( wire4499 ) ;
 assign n_n8332 = ( wire4496 ) | ( wire4497 ) ;
 assign n_n7037 = ( wire4494 ) | ( n_n9353  &  wire2418  &  n_n9639 ) ;
 assign n_n7797 = ( (~ preset)  &  n_n7798 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7005 = ( wire4488 ) | ( wire4489 ) | ( wire4490 ) | ( wire4491 ) ;
 assign n_n7200 = ( (~ preset)  &  n_n7910  &  (~ ndn_latch3_27) ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9633 ) ;
 assign n_n9527 = ( (~ preset)  &  n_n9528  &  (~ nrq3_15) ) | ( (~ preset)  &  nrq3_15  &  n_n9564 ) ;
 assign n_n7523 = ( wire4480 ) | ( wire4481 ) ;
 assign n_n8250 = ( (~ preset)  &  n_n8251 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7483 = ( wire4474 ) | ( wire4475 ) ;
 assign n_n8481 = ( wire4472 ) | ( wire4473 ) ;
 assign n_n7451 = ( (~ preset)  &  n_n9290  &  (~ nrq2_9) ) ;
 assign n_n7055 = ( wire4468 ) | ( wire4469 ) ;
 assign n_n7555 = ( (~ preset)  &  n_n7556 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n9063 = ( wire4464 ) | ( n_n8449  &  wire2418  &  n_n9639 ) ;
 assign n_n7207 = ( wire4462 ) | ( wire4463 ) ;
 assign n_n7100 = ( wire4460 ) | ( ndn3_19  &  (~ ndn3_21)  &  wire2408 ) ;
 assign n_n7799 = ( (~ preset)  &  n_n9361  &  (~ nrq2_9) ) ;
 assign n_n7471 = ( (~ preset)  &  n_n9616  &  nrq3_21 ) | ( (~ preset)  &  n_n9304  &  (~ nrq3_21) ) ;
 assign n_n7219 = ( wire4456 ) | ( n_n8652  &  wire2429  &  n_n9639 ) ;
 assign n_n7614 = ( (~ preset)  &  n_n9616  &  nrq3_18 ) | ( (~ preset)  &  n_n7712  &  (~ nrq3_18) ) ;
 assign n_n7250 = ( wire4452 ) | ( n_n8707  &  wire2429  &  n_n9639 ) ;
 assign n_n7590 = ( wire4450 ) | ( n_n8549  &  wire2431  &  n_n9639 ) ;
 assign n_n6915 = ( wire4448 ) | ( (~ nsr3_13)  &  (~ ndn3_15)  &  wire2408 ) ;
 assign n_n8052 = ( wire4444 ) | ( wire4445 ) ;
 assign n_n9014 = ( (~ preset)  &  n_n9015  &  (~ ndn_latch3_12) ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9627 ) ;
 assign n_n8065 = ( wire4440 ) | ( n_n8354  &  wire2427  &  n_n9639 ) ;
 assign n_n9517 = ( (~ preset)  &  n_n9518  &  (~ ndn_latch3_32) ) | ( (~ preset)  &  ndn_latch3_32  &  n_n9619 ) ;
 assign n_n8089 = ( wire4436 ) | ( wire4437 ) ;
 assign n_n9256 = ( wire4434 ) | ( n_n9448  &  wire2431  &  n_n9639 ) ;
 assign n_n8174 = ( wire4432 ) | ( wire4433 ) ;
 assign n_n8490 = ( wire4428 ) | ( wire4429 ) ;
 assign n_n8113 = ( wire4424 ) | ( wire4425 ) ;
 assign n_n7039 = ( (~ preset)  &  n_n7951  &  (~ ndn_latch3_12) ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9619 ) ;
 assign n_n7095 = ( wire4416 ) | ( wire4417 ) | ( n_n8913  &  wire2451 ) ;
 assign n_n8034 = ( (~ preset)  &  n_n8035  &  (~ nrq3_18) ) | ( (~ preset)  &  nrq3_18  &  n_n9564 ) ;
 assign n_n7094 = ( wire4411 ) | ( wire4412 ) | ( n_n8631  &  wire2451 ) ;
 assign n_n8242 = ( (~ preset)  &  n_n8243 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7855 = ( wire4406 ) | ( wire4407 ) ;
 assign n_n7098 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7632 = ( wire4404 ) | ( ndn3_9  &  (~ ndn3_11)  &  wire2408 ) ;
 assign n_n9079 = ( (~ preset)  &  n_n9175  &  (~ ndn_latch3_27) ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9581 ) ;
 assign n_n7090 = ( wire4400 ) | ( wire4401 ) ;
 assign n_n7299 = ( wire4398 ) | ( n_n9284  &  wire2427  &  n_n9639 ) ;
 assign n_n9480 = ( wire4396 ) | ( wire4397 ) ;
 assign n_n9409 = ( (~ preset)  &  n_n9410  &  (~ nrq2_9) ) ;
 assign n_n7385 = ( wire4394 ) | ( wire2369  &  n_n9619 ) ;
 assign n_n7406 = ( wire4392 ) | ( n_n8707  &  wire2418  &  n_n9639 ) ;
 assign n_n7405 = ( wire4390 ) | ( n_n9512  &  wire2447  &  n_n9639 ) ;
 assign n_n7782 = ( wire4388 ) | ( wire4389 ) ;
 assign n_n7372 = ( wire4386 ) | ( wire2368  &  n_n9619 ) ;
 assign n_n7053 = ( wire4384 ) | ( wire4385 ) ;
 assign n_n7086 = ( wire4382 ) | ( (~ nsr3_13)  &  (~ ndn3_15)  &  wire2406 ) ;
 assign n_n8730 = ( wire4380 ) | ( nen3_16  &  (~ ndn3_16)  &  wire2405 ) ;
 assign n_n1 = ( preset ) | ( pdn ) | ( wire4378 ) ;
 assign n_n9090 = ( wire4376 ) | ( n_n9353  &  wire2421  &  n_n9639 ) ;
 assign n_n7547 = ( (~ preset)  &  n_n8531  &  (~ nrq2_9) ) ;
 assign n_n8335 = ( wire4374 ) | ( n_n9638  &  wire2421  &  n_n9639 ) ;
 assign n_n7323 = ( wire4372 ) | ( n_n7098  &  (~ n_n7311)  &  n_n7544 ) | ( n_n7098  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n9610 = ( wire4370 ) | ( nen3_39  &  (~ ndn3_39)  &  wire2404 ) ;
 assign n_n8111 = ( (~ preset)  &  n_n8112 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n8039 = ( wire4364 ) | ( wire4365 ) ;
 assign n_n9617 = ( (~ preset)  &  n_n9619  &  ndn_latch3_25 ) | ( (~ preset)  &  n_n9618  &  (~ ndn_latch3_25) ) ;
 assign n_n9612 = ( wire4360 ) | ( wire4361 ) ;
 assign n_n9241 = ( (~ preset)  &  n_n9242  &  (~ nrq2_9) ) ;
 assign n_n7383 = ( wire4358 ) | ( n_n9616  &  wire2370 ) ;
 assign n_n6933 = ( (~ preset)  &  n_n9581  &  nrq3_17 ) | ( (~ preset)  &  n_n8884  &  (~ nrq3_17) ) ;
 assign n_n7461 = ( wire4354 ) | ( wire4355 ) ;
 assign n_n7613 = ( wire4352 ) | ( n_n8549  &  wire2421  &  n_n9639 ) ;
 assign n_n8764 = ( wire4350 ) | ( wire2370  &  (~ n_n7566)  &  n_n8154 ) | ( wire2370  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n7014 = ( (~ preset)  &  n_n7909  &  (~ nrq3_36) ) | ( (~ preset)  &  nrq3_36  &  n_n9633 ) ;
 assign n_n7897 = ( wire4346 ) | ( wire2369  &  (~ n_n7566)  &  n_n8154 ) | ( wire2369  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n8379 = ( wire4344 ) | ( (~ ndn3_4)  &  ndn3_2  &  wire2405 ) ;
 assign n_n8861 = ( (~ preset)  &  n_n8862  &  (~ nrq3_34) ) | ( (~ preset)  &  nrq3_34  &  n_n9627 ) ;
 assign n_n8036 = ( (~ preset)  &  n_n8037  &  (~ nrq2_9) ) ;
 assign n_n8026 = ( (~ preset)  &  ndn3_17  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_18 ) ;
 assign n_n7883 = ( (~ preset)  &  nen3_22  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_22 ) ;
 assign n_n8973 = ( (~ preset)  &  n_n8974 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7285 = ( (~ preset)  &  n_n7286 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n9222 = ( wire4330 ) | ( wire4331 ) ;
 assign n_n8147 = ( (~ preset)  &  n_n9246 ) ;
 assign n_n9167 = ( wire4328 ) | ( wire4329 ) ;
 assign n_n8310 = ( wire4326 ) | ( wire4327 ) ;
 assign n_n8317 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_39 ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_38) ) ;
 assign n_n7168 = ( wire4322 ) | ( wire4323 ) ;
 assign n_n7397 = ( (~ preset)  &  n_n9557  &  (~ nrq2_9) ) ;
 assign n_n7165 = ( wire4320 ) | ( n_n8354  &  wire2429  &  n_n9639 ) ;
 assign n_n7070 = ( wire4318 ) | ( wire4319 ) ;
 assign n_n8109 = ( wire4316 ) | ( wire4317 ) ;
 assign n_n7268 = ( wire4314 ) | ( n_n9537  &  wire2418  &  n_n9639 ) ;
 assign n_n8567 = ( (~ preset)  &  n_n8568 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7228 = ( wire4310 ) | ( wire4311 ) ;
 assign n_n7718 = ( (~ preset)  &  n_n7931  &  (~ ndn_latch3_25) ) | ( (~ preset)  &  ndn_latch3_25  &  n_n9633 ) ;
 assign n_n7494 = ( (~ preset)  &  n_n7742  &  (~ ndn_latch3_7) ) | ( (~ preset)  &  ndn_latch3_7  &  n_n9564 ) ;
 assign n_n7235 = ( wire4304 ) | ( ndn3_19  &  (~ ndn3_21)  &  wire2404 ) ;
 assign n_n8218 = ( wire4302 ) | ( n_n8549  &  wire2418  &  n_n9639 ) ;
 assign n_n9567 = ( (~ preset)  &  n_n9568  &  (~ nrq3_4) ) | ( (~ preset)  &  nrq3_4  &  n_n9633 ) ;
 assign n_n9199 = ( (~ preset)  &  n_n9200 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n8544 = ( wire4296 ) | ( wire4297 ) ;
 assign n_n6934 = ( wire4294 ) | ( wire4295 ) ;
 assign n_n6914 = ( wire4292 ) | ( nen3_16  &  (~ ndn3_16)  &  wire2404 ) ;
 assign n_n8735 = ( wire4290 ) | ( wire4291 ) ;
 assign n_n8474 = ( wire4288 ) | ( wire4289 ) ;
 assign n_n8498 = ( (~ preset)  &  n_n8499  &  (~ ndn_latch3_32) ) | ( (~ preset)  &  ndn_latch3_32  &  n_n9564 ) ;
 assign n_n8085 = ( wire4282 ) | ( wire4283 ) ;
 assign n_n7802 = ( wire4280 ) | ( wire4281 ) ;
 assign n_n7061 = ( wire4278 ) | ( ndn3_29  &  (~ ndn3_32)  &  wire2402 ) ;
 assign n_n9097 = ( wire4274 ) | ( wire4275 ) ;
 assign n_n7159 = ( wire4272 ) | ( wire4273 ) ;
 assign n_n7303 = ( (~ preset)  &  n_n9616  &  nrq3_9 ) | ( (~ preset)  &  n_n7713  &  (~ nrq3_9) ) ;
 assign n_n9565 = ( (~ preset)  &  n_n9566  &  (~ nrq3_9) ) | ( (~ preset)  &  nrq3_9  &  n_n9627 ) ;
 assign n_n7833 = ( wire4264 ) | ( wire4265 ) ;
 assign n_n8413 = ( wire4260 ) | ( wire4261 ) ;
 assign n_n6969 = ( wire4258 ) | ( (~ ndn3_7)  &  ndn3_4  &  wire2404 ) ;
 assign n_n8345 = ( (~ preset)  &  n_n9560  &  (~ nrq2_9) ) ;
 assign n_n7800 = ( wire4256 ) | ( wire4257 ) ;
 assign n_n7172 = ( wire4254 ) | ( wire4255 ) ;
 assign n_n7212 = ( (~ preset)  &  n_n8882  &  (~ ndn_latch3_26) ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9581 ) ;
 assign n_n7545 = ( wire4250 ) | ( wire4251 ) ;
 assign n_n7099 = ( wire4248 ) | ( wire4249 ) ;
 assign n_n8997 = ( wire4246 ) | ( ndn3_25  &  (~ ndn3_26)  &  wire2406 ) ;
 assign n_n7479 = ( wire4242 ) | ( wire4243 ) ;
 assign n_n9463 = ( wire4240 ) | ( wire4241 ) ;
 assign n_n8346 = ( wire4238 ) | ( n_n9537  &  wire2431  &  n_n9639 ) ;
 assign n_n8874 = ( (~ preset)  &  n_n8875  &  (~ nrq2_9) ) ;
 assign n_n7354 = ( wire4234 ) | ( wire4235 ) ;
 assign n_n8958 = ( wire4232 ) | ( wire4233 ) ;
 assign n_n8956 = ( wire4230 ) | ( wire2371  &  n_n9619 ) ;
 assign n_n8246 = ( wire4228 ) | ( wire2368  &  n_n9564 ) ;
 assign n_n8257 = ( wire4226 ) | ( wire2370  &  (~ n_n7869)  &  n_n8028 ) | ( wire2370  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n7404 = ( wire4224 ) | ( n_n9416  &  wire2447  &  n_n9639 ) ;
 assign n_n8842 = ( wire4222 ) | ( n_n8821  &  wire2418  &  n_n9639 ) ;
 assign n_n8443 = ( wire4220 ) | ( wire4221 ) ;
 assign n_n7163 = ( (~ preset)  &  n_n7702  &  (~ nrq2_9) ) ;
 assign n_n6 = ( wire16686 ) | ( nsr3_23  &  (~ ndn3_19) ) ;
 assign n_n8025 = ( (~ preset)  &  n_n8199  &  (~ nrq2_9) ) ;
 assign n_n7982 = ( (~ preset)  &  n_n7983  &  (~ nrq2_9) ) ;
 assign n_n7186 = ( wire4215 ) | ( n_n7098  &  n_n9633 ) ;
 assign n_n7248 = ( wire4213 ) | ( wire4214 ) ;
 assign n_n7639 = ( wire4211 ) | ( n_n9434  &  wire2429  &  n_n9639 ) ;
 assign n_n8347 = ( (~ preset)  &  n_n8348  &  (~ nrq2_9) ) ;
 assign n_n8835 = ( wire4207 ) | ( wire4208 ) ;
 assign n_n8444 = ( wire4205 ) | ( n_n8549  &  wire2423  &  n_n9639 ) ;
 assign n_n7425 = ( wire4201 ) | ( wire4202 ) ;
 assign n_n7830 = ( wire4199 ) | ( n_n9638  &  wire2429  &  n_n9639 ) ;
 assign n_n7618 = ( wire4197 ) | ( n_n9616  &  wire2368 ) ;
 assign n_n9062 = ( wire4193 ) | ( wire4194 ) ;
 assign n_n9430 = ( wire4191 ) | ( wire4192 ) ;
 assign n_n8676 = ( wire4189 ) | ( wire4190 ) ;
 assign n_n8023 = ( wire4187 ) | ( wire2368  &  (~ n_n7566)  &  n_n8154 ) | ( wire2368  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n7141 = ( wire4185 ) | ( n_n8419  &  wire2423  &  n_n9639 ) ;
 assign n_n8995 = ( wire4183 ) | ( wire2371  &  (~ n_n7566)  &  n_n8154 ) | ( wire2371  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n7917 = ( wire4181 ) | ( n_n8354  &  wire2423  &  n_n9639 ) ;
 assign n_n8259 = ( wire4179 ) | ( n_n8652  &  wire2431  &  n_n9639 ) ;
 assign n_n9207 = ( wire4177 ) | ( ndn3_17  &  (~ ndn3_18)  &  wire2406 ) ;
 assign n_n9188 = ( wire4175 ) | ( n_n8707  &  wire2431  &  n_n9639 ) ;
 assign n_n9094 = ( wire4173 ) | ( wire4174 ) ;
 assign n_n8179 = ( (~ preset)  &  (~ nsr3_30) ) ;
 assign n_n7773 = ( wire4171 ) | ( wire4172 ) ;
 assign n_n7647 = ( (~ preset)  &  n_n7693  &  (~ ndn_latch3_27) ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9619 ) ;
 assign n_n7038 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_16 ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_14) ) ;
 assign n_n7157 = ( wire4163 ) | ( wire4164 ) ;
 assign n_n8940 = ( wire4161 ) | ( (~ ndn3_29)  &  ndn3_28  &  wire2404 ) ;
 assign n_n8041 = ( wire4159 ) | ( n_n9512  &  wire2427  &  n_n9639 ) ;
 assign n_n8679 = ( wire4157 ) | ( wire4158 ) ;
 assign n_n8658 = ( wire4155 ) | ( n_n8821  &  wire2427  &  n_n9639 ) ;
 assign n_n9109 = ( (~ preset)  &  n_n9616  &  ndn_latch3_32 ) | ( (~ preset)  &  n_n9110  &  (~ ndn_latch3_32) ) ;
 assign n_n9572 = ( wire4151 ) | ( wire4152 ) ;
 assign n_n8950 = ( wire4149 ) | ( wire2370  &  n_n9581 ) ;
 assign n_n9240 = ( wire4147 ) | ( wire2368  &  (~ n_n8019)  &  n_n7573 ) | ( wire2368  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n9386 = ( wire4143 ) | ( wire4144 ) ;
 assign n_n7594 = ( wire4141 ) | ( wire4142 ) ;
 assign n_n7210 = ( wire4139 ) | ( (~ ndn3_27)  &  ndn3_26  &  wire2408 ) ;
 assign n_n8405 = ( (~ preset)  &  n_n8406 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7892 = ( wire4135 ) | ( (~ ndn3_19)  &  nen3_19  &  wire2404 ) ;
 assign n_n7221 = ( wire4133 ) | ( n_n8549  &  wire2447  &  n_n9639 ) ;
 assign n_n7350 = ( (~ preset)  &  n_n7474  &  (~ ndn_latch3_29) ) | ( (~ preset)  &  ndn_latch3_29  &  n_n9619 ) ;
 assign n_n8465 = ( wire4129 ) | ( n_n7098  &  (~ n_n9385)  &  n_n9384 ) | ( n_n7098  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n6983 = ( (~ preset)  &  n_n6984 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7719 = ( wire4125 ) | ( n_n9616  &  wire2367 ) ;
 assign n_n7551 = ( wire4123 ) | ( wire4124 ) ;
 assign n_n8737 = ( (~ preset)  &  n_n9559  &  (~ nrq2_9) ) ;
 assign n_n7361 = ( (~ preset)  &  n_n7362 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n9299 = ( wire4117 ) | ( wire4118 ) ;
 assign n_n9549 = ( (~ preset)  &  n_n9550  &  (~ nrq2_9) ) ;
 assign n_n9287 = ( (~ preset)  &  n_n9581  &  ndn_latch3_25 ) | ( (~ preset)  &  n_n9492  &  (~ ndn_latch3_25) ) ;
 assign n_n8776 = ( wire4113 ) | ( wire4114 ) ;
 assign n_n7009 = ( (~ preset)  &  n_n9616  &  ndn_latch3_7 ) | ( (~ preset)  &  n_n7764  &  (~ ndn_latch3_7) ) ;
 assign n_n7355 = ( wire4107 ) | ( wire4108 ) ;
 assign n_n7776 = ( wire4105 ) | ( wire4106 ) ;
 assign n_n7550 = ( wire4103 ) | ( wire4104 ) ;
 assign n_n8172 = ( (~ preset)  &  n_n8173  &  (~ nrq2_9) ) ;
 assign n_n7497 = ( wire4101 ) | ( wire4102 ) ;
 assign n_n9146 = ( wire4099 ) | ( wire4100 ) ;
 assign n_n8752 = ( (~ preset)  &  n_n8753  &  (~ nrq3_17) ) | ( (~ preset)  &  nrq3_17  &  n_n9619 ) ;
 assign n_n8771 = ( (~ preset)  &  n_n8772  &  (~ nrq3_9) ) | ( (~ preset)  &  nrq3_9  &  n_n9633 ) ;
 assign n_n8048 = ( wire4093 ) | ( wire4094 ) ;
 assign n_n7870 = ( (~ preset)  &  n_n9362  &  (~ nrq2_9) ) ;
 assign n_n7015 = ( (~ preset)  &  (~ pdn)  &  ndn1_4 ) ;
 assign n_n7470 = ( (~ preset)  &  n_n9561  &  (~ nrq2_9) ) ;
 assign n_n9002 = ( wire4091 ) | ( wire4092 ) ;
 assign n_n7532 = ( (~ preset)  &  n_n9616  &  ndn_latch3_12 ) | ( (~ preset)  &  n_n8203  &  (~ ndn_latch3_12) ) ;
 assign n_n7442 = ( wire4087 ) | ( wire4088 ) ;
 assign n_n9078 = ( wire4085 ) | ( wire4086 ) ;
 assign n_n8367 = ( wire4083 ) | ( wire4084 ) ;
 assign n_n9330 = ( (~ preset)  &  n_n9331  &  (~ nrq2_9) ) ;
 assign n_n7103 = ( wire4081 ) | ( (~ ndn3_19)  &  nen3_19  &  wire2402 ) ;
 assign n_n8399 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_7 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_4 ) ;
 assign n_n7526 = ( wire4077 ) | ( wire2370  &  n_n9564 ) ;
 assign n_n9035 = ( wire4075 ) | ( wire2368  &  (~ n_n7869)  &  n_n8028 ) | ( wire2368  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n7264 = ( wire4073 ) | ( n_n9416  &  wire2418  &  n_n9639 ) ;
 assign n_n8696 = ( wire4071 ) | ( n_n8821  &  wire2447  &  n_n9639 ) ;
 assign n_n7080 = ( (~ preset)  &  n_n9581  &  nrq3_15 ) | ( (~ preset)  &  n_n9497  &  (~ nrq3_15) ) ;
 assign n_n7290 = ( (~ preset)  &  n_n7291 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n11 = ( wire16687 ) | ( nsr3_13  &  (~ ndn3_12) ) ;
 assign n_n2 = ( wire16688 ) | ( nsr3_38  &  (~ nen3_36) ) ;
 assign n_n7548 = ( (~ preset)  &  n_n8240  &  (~ nrq2_9) ) ;
 assign n_n7294 = ( (~ preset)  &  n_n7703  &  (~ nrq2_9) ) ;
 assign n_n8949 = ( wire4059 ) | ( n_n7098  &  n_n9619 ) ;
 assign n_n7633 = ( (~ preset)  &  n_n8237  &  (~ nrq2_9) ) ;
 assign n_n8934 = ( (~ preset)  &  n_n8935  &  (~ nrq2_9) ) ;
 assign n_n9243 = ( (~ preset)  &  n_n9244  &  (~ nrq2_9) ) ;
 assign n_n7194 = ( (~ preset)  &  n_n8648  &  (~ nrq2_9) ) ;
 assign n_n7465 = ( (~ preset)  &  n_n8235  &  (~ nrq2_9) ) ;
 assign n_n8610 = ( (~ preset)  &  n_n8611  &  (~ nrq3_39) ) | ( (~ preset)  &  nrq3_39  &  n_n9633 ) ;
 assign n_n7746 = ( wire4053 ) | ( wire4054 ) ;
 assign n_n7349 = ( wire4051 ) | ( ndn3_29  &  (~ ndn3_32)  &  wire2406 ) ;
 assign n_n8169 = ( (~ preset)  &  n_n8572  &  (~ nrq2_9) ) ;
 assign n_n7316 = ( wire4047 ) | ( wire4048 ) ;
 assign n_n8495 = ( wire4045 ) | ( (~ ndn3_9)  &  ndn3_7  &  wire2405 ) ;
 assign n_n6995 = ( (~ preset)  &  n_n9555  &  (~ nrq2_9) ) ;
 assign n_n7468 = ( wire4041 ) | ( wire4042 ) ;
 assign n_n7049 = ( (~ preset)  &  n_n7050 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7304 = ( wire4037 ) | ( (~ ndn3_9)  &  ndn3_7  &  wire2406 ) ;
 assign n_n7139 = ( (~ preset)  &  n_n7140 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7142 = ( wire4033 ) | ( n_n9448  &  wire2423  &  n_n9639 ) ;
 assign n_n6947 = ( (~ preset)  &  n_n6948 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8548 = ( wire4027 ) | ( wire4028 ) | ( wire4029 ) | ( wire4030 ) ;
 assign n_n9543 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_19 ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_19 ) ;
 assign n_n9620 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_28 ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_28 ) ;
 assign n_n7101 = ( wire4021 ) | ( wire4022 ) ;
 assign n_n8092 = ( wire4019 ) | ( wire4020 ) ;
 assign n_n8624 = ( wire4017 ) | ( wire2369  &  (~ n_n9385)  &  n_n9384 ) | ( wire2369  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n8380 = ( wire4015 ) | ( n_n8707  &  wire2427  &  n_n9639 ) ;
 assign n_n6965 = ( wire4013 ) | ( (~ ndn3_19)  &  nen3_19  &  wire2405 ) ;
 assign n_n7891 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_36 ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_37) ) ;
 assign n_n8907 = ( wire4009 ) | ( n_n9284  &  wire2447  &  n_n9639 ) ;
 assign n_n7571 = ( wire4007 ) | ( wire4008 ) ;
 assign n_n7559 = ( (~ preset)  &  n_n7736  &  (~ ndn_latch3_28) ) | ( (~ preset)  &  ndn_latch3_28  &  n_n9564 ) ;
 assign n_n7612 = ( wire4003 ) | ( wire4004 ) ;
 assign n_n8985 = ( wire4001 ) | ( wire4002 ) ;
 assign n_n8890 = ( (~ preset)  &  n_n9619  &  ndn_latch3_28 ) | ( (~ preset)  &  n_n8891  &  (~ ndn_latch3_28) ) ;
 assign n_n7999 = ( wire3997 ) | ( wire3998 ) ;
 assign n_n7220 = ( wire3995 ) | ( n_n8557  &  wire2447  &  n_n9639 ) ;
 assign n_n8748 = ( wire3993 ) | ( wire3994 ) ;
 assign n_n6942 = ( (~ preset)  &  n_n9558  &  (~ nrq2_9) ) ;
 assign n_n9367 = ( wire3991 ) | ( wire2367  &  (~ n_n9385)  &  n_n9384 ) | ( wire2367  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n8518 = ( wire3989 ) | ( (~ nsr3_13)  &  (~ ndn3_15)  &  wire2404 ) ;
 assign n_n6955 = ( (~ preset)  &  n_n6956 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n8297 = ( (~ preset)  &  n_n8298  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9564 ) ;
 assign n_n6922 = ( wire3983 ) | ( (~ ndn3_25)  &  ndn3_22  &  wire2405 ) ;
 assign n_n7016 = ( wire3981 ) | ( wire3982 ) ;
 assign n_n8637 = ( wire3977 ) | ( wire3978 ) ;
 assign n_n9551 = ( (~ preset)  &  n_n9552  &  (~ nrq2_9) ) ;
 assign n_n8286 = ( wire3975 ) | ( wire3976 ) | ( n_n8964  &  wire2451 ) ;
 assign n_n8015 = ( (~ preset)  &  n_n8016  &  (~ nrq2_9) ) ;
 assign n_n7345 = ( wire3972 ) | ( wire3973 ) ;
 assign n_n7010 = ( (~ preset)  &  n_n7696  &  (~ nrq3_4) ) | ( (~ preset)  &  nrq3_4  &  n_n9619 ) ;
 assign n_n8587 = ( wire3968 ) | ( wire3969 ) ;
 assign n_n7097 = ( wire3966 ) | ( (~ ndn3_27)  &  ndn3_26  &  wire2406 ) ;
 assign n_n6953 = ( wire3964 ) | ( n_n9353  &  wire2427  &  n_n9639 ) ;
 assign n_n8457 = ( wire16698 ) | ( (~ preset)  &  n_n8652  &  (~ n_n7274) ) ;
 assign n_n7940 = ( wire16704 ) | ( (~ preset)  &  n_n8707  &  (~ n_n7274) ) ;
 assign n_n8163 = ( wire3953 ) | ( wire3954 ) ;
 assign n_n8860 = ( wire3951 ) | ( wire3952 ) ;
 assign n_n7319 = ( wire3949 ) | ( (~ ndn3_29)  &  ndn3_28  &  wire2405 ) ;
 assign n_n5 = ( wire16705 ) | ( nsr3_30  &  (~ nak3_13) ) ;
 assign n_n6924 = ( (~ preset)  &  n_n8274  &  (~ nrq2_9) ) ;
 assign n_n8614 = ( (~ preset)  &  n_n8615  &  (~ nrq2_9) ) ;
 assign n_n6941 = ( (~ preset)  &  n_n8238  &  (~ nrq2_9) ) ;
 assign n_n7000 = ( (~ preset)  &  n_n7854  &  (~ nrq2_9) ) ;
 assign n_n7280 = ( (~ preset)  &  n_n8649  &  (~ nrq2_9) ) ;
 assign n_n8137 = ( (~ preset)  &  n_n8236  &  (~ nrq2_9) ) ;
 assign n_n7313 = ( (~ preset)  &  n_n8269  &  (~ nrq2_9) ) ;
 assign n_n7832 = ( wire3944 ) | ( n_n9537  &  wire2429  &  n_n9639 ) ;
 assign n_n8021 = ( wire3942 ) | ( wire3943 ) ;
 assign n_n8517 = ( wire3940 ) | ( wire3941 ) ;
 assign n_n8136 = ( (~ preset)  &  n_n8529  &  (~ nrq2_9) ) ;
 assign n_n7122 = ( wire3938 ) | ( nen3_36  &  (~ ndn3_36)  &  wire2404 ) ;
 assign n_n7616 = ( wire3936 ) | ( n_n9434  &  wire2423  &  n_n9639 ) ;
 assign n_n8684 = ( (~ preset)  &  n_n8685  &  (~ nrq2_9) ) ;
 assign n_n9529 = ( (~ preset)  &  n_n9531 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n9509 = ( (~ preset)  &  n_n9510  &  (~ nrq2_9) ) ;
 assign n_n7042 = ( (~ preset)  &  n_n7771  &  (~ nrq2_9) ) ;
 assign n_n8479 = ( wire3932 ) | ( n_n8449  &  wire2421  &  n_n9639 ) ;
 assign n_n8542 = ( wire3930 ) | ( wire3931 ) ;
 assign n_n7088 = ( wire3928 ) | ( nen3_36  &  (~ ndn3_36)  &  wire2408 ) ;
 assign n_n7096 = ( (~ preset)  &  ndn3_9  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_11 ) ;
 assign n_n8878 = ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_13) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_15 ) ;
 assign n_n8331 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_19 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_21 ) ;
 assign n_n7301 = ( (~ preset)  &  n_n7584  &  (~ nrq2_9) ) ;
 assign n_n7972 = ( wire3918 ) | ( wire3919 ) | ( wire3920 ) | ( wire3921 ) ;
 assign n_n6951 = ( (~ preset)  &  n_n6952 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8863 = ( wire3914 ) | ( ndn3_29  &  (~ ndn3_32)  &  wire2404 ) ;
 assign n_n6993 = ( wire3910 ) | ( wire3911 ) ;
 assign n_n7057 = ( wire3908 ) | ( wire3909 ) ;
 assign n_n7143 = ( wire3906 ) | ( n_n8549  &  wire2429  &  n_n9639 ) ;
 assign n_n6945 = ( wire3904 ) | ( n_n9284  &  wire2418  &  n_n9639 ) ;
 assign n_n9101 = ( wire3902 ) | ( wire3903 ) ;
 assign n_n7307 = ( (~ preset)  &  n_n7308 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7300 = ( wire3896 ) | ( wire3897 ) ;
 assign n_n7036 = ( wire3894 ) | ( n_n9537  &  wire2447  &  n_n9639 ) ;
 assign n_n8759 = ( wire3892 ) | ( wire3893 ) ;
 assign n_n6911 = ( (~ preset)  &  n_n6912 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n7352 = ( wire3888 ) | ( wire3889 ) ;
 assign n_n7535 = ( wire3886 ) | ( wire3887 ) | ( n_n8911  &  wire2451 ) ;
 assign n_n7457 = ( (~ preset)  &  n_n7952  &  (~ nrq3_15) ) | ( (~ preset)  &  nrq3_15  &  n_n9619 ) ;
 assign n_n8703 = ( (~ preset)  &  n_n8704 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7520 = ( wire3879 ) | ( nen3_16  &  (~ ndn3_16)  &  wire2402 ) ;
 assign n_n8475 = ( wire3877 ) | ( wire2367  &  (~ n_n8019)  &  n_n7573 ) | ( wire2367  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n8429 = ( wire3875 ) | ( wire3876 ) ;
 assign n_n9018 = ( (~ preset)  &  n_n9616  &  nrq3_17 ) | ( (~ preset)  &  n_n9019  &  (~ nrq3_17) ) ;
 assign n_n7698 = ( (~ preset)  &  n_n7699 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n6972 = ( (~ preset)  &  n_n7375  &  (~ nrq3_17) ) | ( (~ preset)  &  nrq3_17  &  n_n9564 ) ;
 assign n_n7480 = ( wire3865 ) | ( wire3866 ) ;
 assign n_n8338 = ( wire3863 ) | ( wire3864 ) ;
 assign n_n7213 = ( wire3861 ) | ( ndn3_25  &  (~ ndn3_26)  &  wire2405 ) ;
 assign n_n6960 = ( wire3859 ) | ( wire3860 ) ;
 assign n_n9427 = ( wire3857 ) | ( wire3858 ) ;
 assign n_n7478 = ( wire3853 ) | ( wire3854 ) ;
 assign n_n7060 = ( wire3851 ) | ( (~ ndn3_34)  &  nen3_34  &  wire2406 ) ;
 assign n_n7318 = ( (~ preset)  &  n_n7582  &  (~ nrq2_9) ) ;
 assign n_n8967 = ( (~ preset)  &  n_n8968  &  (~ nrq2_9) ) ;
 assign n_n9369 = ( wire3849 ) | ( wire3850 ) ;
 assign n_n7320 = ( wire3847 ) | ( wire3848 ) ;
 assign n_n7867 = ( wire3843 ) | ( wire3844 ) ;
 assign n_n9372 = ( (~ preset)  &  n_n9373 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n10 = ( wire2469 ) | ( n_n9248  &  (~ n_n9247) ) | ( n_n9248  &  (~ n_n9246) ) ;
 assign n_n6940 = ( wire3839 ) | ( wire2367  &  (~ n_n7869)  &  n_n8028 ) | ( wire2367  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n6925 = ( wire3837 ) | ( wire3838 ) ;
 assign n_n7007 = ( (~ preset)  &  n_n8273  &  (~ nrq2_9) ) ;
 assign n_n6936 = ( (~ preset)  &  n_n6937 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7198 = ( wire3833 ) | ( nen3_16  &  (~ ndn3_16)  &  wire2406 ) ;
 assign n_n8547 = ( wire3829 ) | ( wire3830 ) ;
 assign n_n6954 = ( wire3827 ) | ( wire2371  &  n_n9633 ) ;
 assign n_n9622 = ( wire3825 ) | ( wire2368  &  (~ n_n7311)  &  n_n7544 ) | ( wire2368  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n9469 = ( wire3823 ) | ( wire3824 ) ;
 assign n_n7569 = ( wire3821 ) | ( wire3822 ) ;
 assign n_n7339 = ( wire3819 ) | ( n_n9284  &  wire2423  &  n_n9639 ) ;
 assign n_n9364 = ( wire3817 ) | ( wire3818 ) ;
 assign n_n7180 = ( (~ preset)  &  n_n7181 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n8738 = ( wire3811 ) | ( wire3812 ) ;
 assign n_n6932 = ( wire3809 ) | ( wire3810 ) ;
 assign n_n7255 = ( wire3807 ) | ( wire3808 ) ;
 assign n_n7519 = ( wire3805 ) | ( (~ ndn3_17)  &  ndn3_16  &  wire2406 ) ;
 assign n_n7486 = ( (~ preset)  &  n_n7487  &  (~ ndn_latch3_26) ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9564 ) ;
 assign n_n7259 = ( wire3801 ) | ( wire3802 ) ;
 assign n_n8460 = ( wire3799 ) | ( wire3800 ) ;
 assign n_n7987 = ( wire3797 ) | ( n_n8449  &  wire2436  &  n_n9639 ) ;
 assign n_n8378 = ( (~ preset)  &  n_n9581  &  nrq3_4 ) | ( (~ preset)  &  n_n9181  &  (~ nrq3_4) ) ;
 assign n_n8724 = ( (~ preset)  &  n_n8725 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n8625 = ( wire3791 ) | ( wire3792 ) ;
 assign n_n9082 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_27 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_26 ) ;
 assign n_n8209 = ( wire3787 ) | ( n_n8652  &  wire2427  &  n_n9639 ) ;
 assign n_n7414 = ( (~ preset)  &  n_n7415 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8899 = ( wire3783 ) | ( n_n8557  &  wire2429  &  n_n9639 ) ;
 assign n_n7477 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_19 ) | ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_20) ) ;
 assign n_n8761 = ( (~ preset)  &  n_n8762 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7996 = ( (~ preset)  &  n_n8512  &  (~ ndn_latch3_32) ) | ( (~ preset)  &  ndn_latch3_32  &  n_n9633 ) ;
 assign n_n8094 = ( wire3775 ) | ( n_n8821  &  wire2436  &  n_n9639 ) ;
 assign n_n7112 = ( wire3773 ) | ( (~ ndn3_19)  &  nen3_19  &  wire2406 ) ;
 assign n_n7386 = ( (~ preset)  &  n_n7387 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8768 = ( wire3769 ) | ( n_n9434  &  wire2418  &  n_n9639 ) ;
 assign n_n7611 = ( wire3765 ) | ( wire3766 ) ;
 assign n_n7834 = ( wire3761 ) | ( wire3762 ) ;
 assign n_n9156 = ( (~ preset)  &  n_n9616  &  ndn_latch3_28 ) | ( (~ preset)  &  n_n9157  &  (~ ndn_latch3_28) ) ;
 assign n_n8551 = ( wire3757 ) | ( nen3_36  &  (~ ndn3_36)  &  wire2402 ) ;
 assign n_n7380 = ( (~ preset)  &  n_n7381 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n9445 = ( (~ preset)  &  n_n9446 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8632 = ( (~ preset)  &  n_n8633 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n7353 = ( wire3749 ) | ( wire2367  &  (~ n_n7566)  &  n_n8154 ) | ( wire2367  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n7309 = ( (~ preset)  &  n_n7310 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n8401 = ( wire3745 ) | ( ndn3_17  &  (~ ndn3_18)  &  wire2408 ) ;
 assign n_n7488 = ( wire3743 ) | ( wire3744 ) ;
 assign n_n7733 = ( wire3741 ) | ( n_n8821  &  wire2429  &  n_n9639 ) ;
 assign n_n8503 = ( wire3737 ) | ( wire3738 ) ;
 assign n_n8455 = ( wire3733 ) | ( wire3734 ) ;
 assign n_n7512 = ( wire3731 ) | ( wire3732 ) ;
 assign n_n7314 = ( (~ preset)  &  n_n7315 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n9474 = ( (~ preset)  &  n_n9476 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8275 = ( wire3725 ) | ( wire3726 ) ;
 assign n_n8832 = ( wire3723 ) | ( n_n9638  &  wire2431  &  n_n9639 ) ;
 assign n_n7921 = ( wire3721 ) | ( wire3722 ) ;
 assign n_n7105 = ( wire3719 ) | ( (~ ndn3_28)  &  nen3_28  &  wire2405 ) ;
 assign n_n9511 = ( wire16717 ) | ( (~ n_n8431)  &  wire16715 ) | ( (~ n_n8431)  &  wire16716 ) ;
 assign n_n8763 = ( wire3713 ) | ( wire3714 ) ;
 assign n_n4 = ( wire16719 ) | ( (~ ndn3_29)  &  nsr3_35 ) ;
 assign n_n7153 = ( (~ preset)  &  n_n7154 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8754 = ( (~ preset)  &  n_n9581  &  nrq3_16 ) | ( (~ preset)  &  n_n9495  &  (~ nrq3_16) ) ;
 assign n_n7592 = ( wire3704 ) | ( wire3705 ) ;
 assign n_n8853 = ( wire3702 ) | ( wire2367  &  n_n9619 ) ;
 assign n_n8620 = ( wire3700 ) | ( wire3701 ) ;
 assign n_n9214 = ( wire3696 ) | ( wire3697 ) ;
 assign n_n8987 = ( wire3694 ) | ( wire3695 ) ;
 assign n_n7895 = ( wire3692 ) | ( wire2370  &  (~ n_n7311)  &  n_n7544 ) | ( wire2370  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n8071 = ( wire3690 ) | ( wire3691 ) ;
 assign n_n8969 = ( (~ preset)  &  n_n8970  &  (~ nrq2_9) ) ;
 assign n_n8714 = ( wire3686 ) | ( wire3687 ) ;
 assign n_n8485 = ( wire3684 ) | ( wire3685 ) ;
 assign n_n7245 = ( (~ preset)  &  n_n7246 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7865 = ( wire3678 ) | ( wire3679 ) ;
 assign n_n8336 = ( wire3676 ) | ( wire3677 ) ;
 assign n_n7634 = ( (~ preset)  &  n_n7635 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7508 = ( wire3672 ) | ( ndn3_11  &  (~ ndn3_12)  &  wire2406 ) ;
 assign n_n7359 = ( wire3670 ) | ( wire3671 ) ;
 assign n_n8559 = ( wire3668 ) | ( nen3_39  &  (~ ndn3_39)  &  wire2405 ) ;
 assign n_n9107 = ( (~ preset)  &  n_n9108  &  (~ nrq3_34) ) | ( (~ preset)  &  nrq3_34  &  n_n9633 ) ;
 assign n_n9285 = ( (~ preset)  &  n_n9286  &  (~ ndn_latch3_26) ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9619 ) ;
 assign n_n7460 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_11 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_12 ) ;
 assign n_n8540 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_16 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_16 ) ;
 assign n_n7296 = ( (~ preset)  &  n_n9616  &  nrq3_36 ) | ( (~ preset)  &  n_n7708  &  (~ nrq3_36) ) ;
 assign n_n7192 = ( wire3656 ) | ( n_n8419  &  wire2436  &  n_n9639 ) ;
 assign n_n7058 = ( wire3654 ) | ( n_n8652  &  wire2436  &  n_n9639 ) ;
 assign n_n7297 = ( (~ preset)  &  n_n7947  &  (~ nrq3_34) ) | ( (~ preset)  &  nrq3_34  &  n_n9619 ) ;
 assign n_n9213 = ( wire3648 ) | ( wire3649 ) ;
 assign n_n7370 = ( wire3646 ) | ( n_n8707  &  wire2436  &  n_n9639 ) ;
 assign n_n8463 = ( wire3644 ) | ( ndn3_19  &  (~ ndn3_21)  &  wire2405 ) ;
 assign n_n7658 = ( (~ preset)  &  n_n7659 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7238 = ( (~ preset)  &  n_n7630  &  (~ nrq2_9) ) ;
 assign n_n7109 = ( wire3640 ) | ( ndn3_19  &  (~ ndn3_21)  &  wire2406 ) ;
 assign n_n8690 = ( (~ preset)  &  n_n8691  &  (~ nrq2_9) ) ;
 assign n_n6943 = ( wire3638 ) | ( n_n9434  &  wire2447  &  n_n9639 ) ;
 assign n_n9326 = ( wire3636 ) | ( (~ ndn3_28)  &  nen3_28  &  wire2402 ) ;
 assign n_n7994 = ( (~ preset)  &  n_n7995  &  (~ nrq3_36) ) | ( (~ preset)  &  nrq3_36  &  n_n9627 ) ;
 assign n_n7394 = ( wire3632 ) | ( wire3633 ) ;
 assign n_n7589 = ( wire3630 ) | ( (~ nsr3_13)  &  (~ ndn3_15)  &  wire2402 ) ;
 assign n_n7506 = ( (~ preset)  &  n_n7507 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n7958 = ( (~ preset)  &  n_n7959 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7503 = ( wire3624 ) | ( wire3625 ) ;
 assign n_n8008 = ( wire3622 ) | ( wire3623 ) ;
 assign n_n7562 = ( wire3620 ) | ( wire3621 ) ;
 assign n_n7223 = ( wire3618 ) | ( n_n9448  &  wire2418  &  n_n9639 ) ;
 assign n_n8105 = ( (~ preset)  &  n_n8106  &  (~ nrq3_15) ) | ( (~ preset)  &  nrq3_15  &  n_n9633 ) ;
 assign n_n7456 = ( wire3614 ) | ( wire3615 ) ;
 assign n_n7043 = ( wire3610 ) | ( wire3611 ) ;
 assign n_n7279 = ( wire3606 ) | ( wire3607 ) ;
 assign n_n8960 = ( wire3604 ) | ( (~ ndn3_9)  &  ndn3_7  &  wire2402 ) ;
 assign n_n8013 = ( wire3602 ) | ( (~ ndn3_9)  &  ndn3_7  &  wire2404 ) ;
 assign n_n9276 = ( wire3600 ) | ( wire3601 ) ;
 assign n_n9086 = ( (~ preset)  &  n_n9087  &  (~ nrq3_21) ) | ( (~ preset)  &  nrq3_21  &  n_n9627 ) ;
 assign n_n7542 = ( wire3594 ) | ( wire3595 ) ;
 assign n_n7448 = ( (~ preset)  &  n_n7852  &  (~ nrq2_9) ) ;
 assign n_n8164 = ( wire3590 ) | ( wire3591 ) ;
 assign n_n8478 = ( (~ preset)  &  (~ n_n9198) ) | ( (~ preset)  &  (~ n_n9639)  &  n_n9197 ) ;
 assign n_n9415 = ( wire3586 ) | ( wire3587 ) | ( wire3588 ) | ( wire3589 ) ;
 assign n_n9 = ( preset ) | ( wire16726 ) | ( nsr3_13  &  nsr3_14 ) ;
 assign n_n0 = ( wire3581 ) | ( wire3582 ) | ( wire16732 ) ;
 assign n_n7025 = ( (~ preset)  &  n_n7026 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n8855 = ( wire3575 ) | ( wire3576 ) ;
 assign n_n7894 = ( (~ preset)  &  n_n8272  &  (~ nrq2_9) ) ;
 assign n_n7249 = ( wire3573 ) | ( n_n9284  &  wire2429  &  n_n9639 ) ;
 assign n_n7984 = ( (~ preset)  &  n_n7985  &  (~ nrq2_9) ) ;
 assign n_n8311 = ( (~ preset)  &  n_n8312  &  (~ nrq2_9) ) ;
 assign n_n7230 = ( wire3571 ) | ( wire3572 ) ;
 assign n_n7317 = ( wire3567 ) | ( wire3568 ) ;
 assign n_n8799 = ( wire3565 ) | ( wire3566 ) ;
 assign n_n8682 = ( (~ preset)  &  n_n8683 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n9425 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_39 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_39 ) ;
 assign n_n8244 = ( (~ preset)  &  n_n8245 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n9457 = ( wire3557 ) | ( (~ ndn3_34)  &  nen3_34  &  wire2402 ) ;
 assign n_n9301 = ( wire3553 ) | ( wire3554 ) ;
 assign n_n7391 = ( wire3551 ) | ( wire3552 ) ;
 assign n_n6962 = ( wire3549 ) | ( wire3550 ) ;
 assign n_n6916 = ( wire3547 ) | ( n_n8419  &  wire2429  &  n_n9639 ) ;
 assign n_n7224 = ( wire3545 ) | ( n_n9638  &  wire2418  &  n_n9639 ) ;
 assign n_n7505 = ( wire3541 ) | ( wire3542 ) ;
 assign n_n7169 = ( (~ preset)  &  n_n9616  &  ndn_latch3_29 ) | ( (~ preset)  &  n_n8201  &  (~ ndn_latch3_29) ) ;
 assign n_n6970 = ( wire3537 ) | ( (~ ndn3_4)  &  ndn3_2  &  wire2408 ) ;
 assign n_n8176 = ( wire3535 ) | ( wire3536 ) ;
 assign n_n8388 = ( (~ preset)  &  n_n8389 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7998 = ( (~ preset)  &  n_n9440  &  (~ nrq2_9) ) ;
 assign n_n7595 = ( wire3531 ) | ( wire3532 ) ;
 assign n_n6996 = ( wire3529 ) | ( n_n8354  &  wire2418  &  n_n9639 ) ;
 assign n_n7263 = ( wire3527 ) | ( n_n9448  &  wire2447  &  n_n9639 ) ;
 assign n_n7979 = ( wire3525 ) | ( n_n9416  &  wire2429  &  n_n9639 ) ;
 assign n_n6992 = ( wire3521 ) | ( wire3522 ) ;
 assign n_n7675 = ( wire3519 ) | ( (~ ndn3_7)  &  ndn3_4  &  wire2408 ) ;
 assign n_n8395 = ( wire3517 ) | ( n_n8354  &  wire2431  &  n_n9639 ) ;
 assign n_n9532 = ( wire3515 ) | ( wire3516 ) ;
 assign n_n7208 = ( (~ preset)  &  n_n7209 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7002 = ( (~ preset)  &  n_n7003 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7004 = ( (~ preset)  &  n_n7695  &  (~ nrq3_9) ) | ( (~ preset)  &  nrq3_9  &  n_n9619 ) ;
 assign n_n7623 = ( wire3507 ) | ( nen3_39  &  (~ ndn3_39)  &  wire2402 ) ;
 assign n_n8790 = ( wire3505 ) | ( wire3506 ) ;
 assign n_n7253 = ( (~ preset)  &  n_n7374  &  (~ nrq3_19) ) | ( (~ preset)  &  nrq3_19  &  n_n9564 ) ;
 assign n_n7161 = ( wire3501 ) | ( wire3502 ) ;
 assign n_n7943 = ( (~ preset)  &  n_n7944 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n6997 = ( wire3497 ) | ( n_n9537  &  wire2427  &  n_n9639 ) ;
 assign n_n8098 = ( wire3495 ) | ( wire3496 ) ;
 assign n_n6987 = ( (~ preset)  &  n_n6988 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n6985 = ( (~ preset)  &  n_n6986 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8926 = ( wire3489 ) | ( wire3490 ) | ( n_n8933  &  wire2451 ) ;
 assign n_n7116 = ( (~ preset)  &  n_n7117 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8372 = ( wire3484 ) | ( n_n9284  &  wire2421  &  n_n9639 ) ;
 assign n_n7379 = ( (~ preset)  &  n_n8241  &  (~ nrq2_9) ) ;
 assign n_n9218 = ( wire3482 ) | ( n_n7098  &  (~ n_n7869)  &  n_n8028 ) | ( n_n7098  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n7048 = ( (~ preset)  &  n_n8198  &  (~ nrq2_9) ) ;
 assign n_n8080 = ( wire3480 ) | ( wire3481 ) ;
 assign n_n7131 = ( (~ preset)  &  n_n8575  &  (~ nrq2_9) ) ;
 assign n_n8709 = ( (~ preset)  &  n_n8710  &  (~ nrq2_9) ) ;
 assign n_n7621 = ( (~ preset)  &  n_n7622 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7340 = ( wire3476 ) | ( n_n8557  &  wire2421  &  n_n9639 ) ;
 assign n_n7114 = ( wire3474 ) | ( n_n8449  &  wire2423  &  n_n9639 ) ;
 assign n_n7032 = ( (~ preset)  &  n_n7033 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n9088 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_34 ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_34 ) ;
 assign n_n9185 = ( wire3468 ) | ( n_n9512  &  wire2431  &  n_n9639 ) ;
 assign n_n8129 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_50 ) ;
 assign n_n7564 = ( wire3466 ) | ( n_n9416  &  wire2431  &  n_n9639 ) ;
 assign n_n7018 = ( (~ preset)  &  n_n7019 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8309 = ( wire3462 ) | ( wire2369  &  n_n9581 ) ;
 assign n_n7260 = ( (~ preset)  &  n_n7261 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7839 = ( wire3458 ) | ( ndn3_29  &  (~ ndn3_32)  &  wire2408 ) ;
 assign n_n7619 = ( wire3456 ) | ( wire3457 ) ;
 assign n_n7992 = ( (~ preset)  &  n_n7993  &  (~ nrq3_36) ) | ( (~ preset)  &  nrq3_36  &  n_n9564 ) ;
 assign n_n7138 = ( wire3452 ) | ( wire3453 ) ;
 assign n_n8252 = ( wire3450 ) | ( wire3451 ) ;
 assign n_n8888 = ( wire3448 ) | ( wire3449 ) ;
 assign n_n7234 = ( wire3446 ) | ( wire3447 ) ;
 assign n_n8917 = ( (~ preset)  &  n_n8918 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n7501 = ( (~ preset)  &  n_n8515  &  (~ nrq3_17) ) | ( (~ preset)  &  nrq3_17  &  n_n9633 ) ;
 assign n_n7084 = ( (~ preset)  &  n_n7933  &  (~ nrq3_16) ) | ( (~ preset)  &  nrq3_16  &  n_n9633 ) ;
 assign n_n8074 = ( (~ preset)  &  n_n8075  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9627 ) ;
 assign n_n7337 = ( (~ preset)  &  n_n7338 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n8103 = ( (~ preset)  &  n_n8104  &  (~ nrq3_17) ) | ( (~ preset)  &  nrq3_17  &  n_n9627 ) ;
 assign n_n8170 = ( (~ preset)  &  n_n8171  &  (~ nrq2_9) ) ;
 assign n_n9058 = ( wire3432 ) | ( n_n8707  &  wire2423  &  n_n9639 ) ;
 assign n_n9022 = ( wire3428 ) | ( wire3429 ) ;
 assign n_n7152 = ( wire3424 ) | ( wire3425 ) ;
 assign n_n8952 = ( (~ preset)  &  n_n9441  &  (~ nrq2_9) ) ;
 assign n_n6919 = ( wire3422 ) | ( wire3423 ) ;
 assign n_n8830 = ( (~ preset)  &  n_n8831 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8440 = ( (~ preset)  &  n_n8441 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8231 = ( wire3416 ) | ( wire2371  &  n_n9564 ) ;
 assign n_n9251 = ( wire3414 ) | ( wire3415 ) ;
 assign n_n7981 = ( (~ preset)  &  n_n9363  &  (~ nrq2_9) ) ;
 assign n_n8565 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_4 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_2 ) ;
 assign n_n9461 = ( wire3410 ) | ( wire3411 ) ;
 assign n_n7560 = ( (~ preset)  &  n_n7561 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n8922 = ( wire3406 ) | ( wire3407 ) | ( n_n8923  &  wire2451 ) ;
 assign n_n7977 = ( (~ preset)  &  n_n7978 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n7828 = ( wire3401 ) | ( wire3402 ) | ( n_n8978  &  wire2451 ) ;
 assign n_n7170 = ( (~ preset)  &  n_n9581  &  ndn_latch3_7 ) | ( (~ preset)  &  n_n9499  &  (~ ndn_latch3_7) ) ;
 assign n_n8712 = ( (~ preset)  &  n_n8713 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n8943 = ( (~ preset)  &  n_n8944 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7371 = ( (~ preset)  &  n_n8239  &  (~ nrq2_9) ) ;
 assign n_n7215 = ( (~ preset)  &  n_n7652  &  (~ ndn_latch3_25) ) | ( (~ preset)  &  ndn_latch3_25  &  n_n9627 ) ;
 assign n_n7027 = ( wire3390 ) | ( wire3391 ) ;
 assign n_n6982 = ( (~ preset)  &  n_n8530  &  (~ nrq2_9) ) ;
 assign n_n7115 = ( wire3388 ) | ( wire3389 ) ;
 assign n_n7072 = ( wire3386 ) | ( wire3387 ) ;
 assign n_n7445 = ( wire3384 ) | ( n_n9616  &  wire2369 ) ;
 assign n_n7963 = ( wire3382 ) | ( wire3383 ) ;
 assign n_n7348 = ( wire3380 ) | ( (~ ndn3_34)  &  nen3_34  &  wire2408 ) ;
 assign n_n8897 = ( wire3378 ) | ( wire3379 ) ;
 assign n_n7974 = ( wire3376 ) | ( wire3377 ) ;
 assign n_n7648 = ( wire3374 ) | ( (~ ndn3_27)  &  ndn3_26  &  wire2402 ) ;
 assign n_n7035 = ( wire3370 ) | ( wire3371 ) ;
 assign n_n7960 = ( (~ preset)  &  n_n7961  &  (~ nrq2_9) ) ;
 assign n_n7423 = ( wire3366 ) | ( wire3367 ) ;
 assign n_n7475 = ( wire3364 ) | ( wire3365 ) ;
 assign n_n8766 = ( wire3362 ) | ( wire2369  &  (~ n_n8019)  &  n_n7573 ) | ( wire2369  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n9032 = ( wire3360 ) | ( wire2368  &  (~ n_n9385)  &  n_n9384 ) | ( wire2368  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n8829 = ( (~ preset)  &  n_n9161 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n8186 = ( wire3356 ) | ( wire3357 ) ;
 assign n_n9120 = ( wire3352 ) | ( wire3353 ) ;
 assign n_n8059 = ( wire3350 ) | ( wire3351 ) ;
 assign n_n7801 = ( wire3348 ) | ( wire3349 ) ;
 assign n_n7450 = ( (~ preset)  &  n_n9360  &  (~ nrq2_9) ) ;
 assign n_n9204 = ( wire3346 ) | ( ndn3_25  &  (~ ndn3_26)  &  wire2408 ) ;
 assign n_n8391 = ( (~ preset)  &  n_n8392 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n7538 = ( wire3342 ) | ( wire3343 ) | ( n_n9034  &  wire2451 ) ;
 assign n_n8374 = ( (~ preset)  &  n_n8375  &  (~ ndn_latch3_7) ) | ( (~ preset)  &  ndn_latch3_7  &  n_n9619 ) ;
 assign n_n8327 = ( wire3337 ) | ( n_n9416  &  wire2421  &  n_n9639 ) ;
 assign n_n9297 = ( (~ preset)  &  n_n9298  &  (~ nrq2_9) ) ;
 assign n_n7062 = ( wire3335 ) | ( wire3336 ) ;
 assign n_n8505 = ( wire3331 ) | ( wire3332 ) ;
 assign n_n7729 = ( (~ preset)  &  (~ pdn)  &  (~ nsr1_2) ) ;
 assign n_n7226 = ( wire3327 ) | ( wire3328 ) ;
 assign n_n7419 = ( wire3325 ) | ( wire3326 ) ;
 assign n_n7957 = ( (~ preset)  &  n_n9291  &  (~ nrq2_9) ) ;
 assign n_n7945 = ( wire3321 ) | ( wire3322 ) ;
 assign n_n7662 = ( wire3319 ) | ( ndn3_11  &  (~ ndn3_12)  &  wire2404 ) ;
 assign n_n8254 = ( wire3317 ) | ( wire3318 ) ;
 assign n_n9037 = ( wire3315 ) | ( n_n9353  &  wire2431  &  n_n9639 ) ;
 assign n_n7282 = ( wire3313 ) | ( wire3314 ) ;
 assign n_n7082 = ( wire3309 ) | ( wire3310 ) ;
 assign n_n7388 = ( wire3307 ) | ( wire3308 ) ;
 assign n_n9001 = ( (~ preset)  &  n_n9351  &  (~ nrq3_21) ) | ( (~ preset)  &  nrq3_21  &  n_n9619 ) ;
 assign n_n6967 = ( wire3303 ) | ( n_n9638  &  wire2436  &  n_n9639 ) ;
 assign n_n8451 = ( n_n8668  &  (~ wire2469) ) ;
 assign n_n7044 = ( wire3299 ) | ( wire3300 ) ;
 assign n_n7012 = ( (~ preset)  &  n_n7013 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n9625 = ( wire3295 ) | ( n_n7098  &  n_n9627 ) ;
 assign n_n7132 = ( (~ preset)  &  n_n8200  &  (~ nrq2_9) ) ;
 assign n_n8645 = ( wire3293 ) | ( n_n7098  &  n_n9564 ) ;
 assign n_n8802 = ( (~ preset)  &  n_n8803  &  (~ nrq2_9) ) ;
 assign n_n9569 = ( wire3291 ) | ( wire3292 ) ;
 assign n_n8365 = ( (~ preset)  &  n_n8366  &  (~ nrq2_9) ) ;
 assign n_n7104 = ( wire3289 ) | ( wire3290 ) ;
 assign n_n7785 = ( (~ preset)  &  n_n8650  &  (~ nrq2_9) ) ;
 assign n_n7006 = ( (~ preset)  &  n_n8574  &  (~ nrq2_9) ) ;
 assign n_n7275 = ( (~ preset)  &  n_n7276 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n9211 = ( wire3283 ) | ( wire3284 ) ;
 assign n_n8382 = ( wire3281 ) | ( wire3282 ) ;
 assign n_n9453 = ( (~ preset)  &  (~ nsr3_35) ) ;
 assign n_n8434 = ( wire3277 ) | ( wire3278 ) | ( wire3279 ) | ( wire3280 ) ;
 assign n_n7574 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_44 ) ;
 assign n_n6981 = ( wire3271 ) | ( wire3272 ) ;
 assign n_n6966 = ( wire3269 ) | ( wire3270 ) ;
 assign n_n7700 = ( wire3267 ) | ( wire3268 ) ;
 assign n_n7126 = ( (~ preset)  &  n_n9359  &  (~ nrq2_9) ) ;
 assign n_n8424 = ( (~ preset)  &  n_n8425  &  (~ ndn_latch3_28) ) | ( (~ preset)  &  ndn_latch3_28  &  n_n9633 ) ;
 assign n_n9103 = ( wire3263 ) | ( wire2371  &  (~ n_n8019)  &  n_n7573 ) | ( wire2371  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n9220 = ( wire3261 ) | ( wire2370  &  (~ n_n9385)  &  n_n9384 ) | ( wire2370  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n9447 = ( wire3257 ) | ( wire3258 ) | ( wire3259 ) | ( wire3260 ) ;
 assign n_n8593 = ( wire3253 ) | ( wire3254 ) | ( wire3255 ) | ( wire3256 ) ;
 assign n_n7233 = ( wire3251 ) | ( (~ ndn3_25)  &  ndn3_22  &  wire2404 ) ;
 assign n_n7466 = ( (~ preset)  &  n_n7467 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8232 = ( wire3247 ) | ( wire3248 ) ;
 assign n_n7167 = ( wire3245 ) | ( wire2367  &  n_n9633 ) ;
 assign n_n8063 = ( wire3243 ) | ( n_n8557  &  wire2418  &  n_n9639 ) ;
 assign n_n9039 = ( (~ preset)  &  n_n9162 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n7916 = ( wire3239 ) | ( (~ ndn3_4)  &  ndn3_2  &  wire2404 ) ;
 assign n_n8054 = ( (~ preset)  &  n_n8055 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7267 = ( wire3235 ) | ( n_n8354  &  wire2447  &  n_n9639 ) ;
 assign n_n8255 = ( wire3233 ) | ( n_n7098  &  (~ n_n8019)  &  n_n7573 ) | ( n_n7098  &  n_n8019  &  (~ n_n7573) ) ;
 assign n_n7924 = ( wire3231 ) | ( n_n9512  &  wire2429  &  n_n9639 ) ;
 assign n_n7502 = ( (~ preset)  &  n_n9616  &  nrq3_16 ) | ( (~ preset)  &  n_n7762  &  (~ nrq3_16) ) ;
 assign n_n7258 = ( wire3227 ) | ( wire3228 ) ;
 assign n_n7262 = ( wire3223 ) | ( wire3224 ) ;
 assign n_n7705 = ( wire3221 ) | ( n_n9416  &  wire2423  &  n_n9639 ) ;
 assign n_n7293 = ( wire3219 ) | ( wire3220 ) ;
 assign n_n9419 = ( wire3217 ) | ( wire3218 ) ;
 assign n_n7625 = ( wire3215 ) | ( wire3216 ) ;
 assign n_n7093 = ( wire3213 ) | ( wire3214 ) ;
 assign n_n8261 = ( wire3211 ) | ( wire3212 ) ;
 assign n_n8442 = ( (~ preset)  &  n_n9100  &  (~ nrq3_21) ) | ( (~ preset)  &  nrq3_21  &  n_n9564 ) ;
 assign n_n7516 = ( wire3207 ) | ( n_n9353  &  wire2436  &  n_n9639 ) ;
 assign n_n6923 = ( wire3205 ) | ( n_n9537  &  wire2436  &  n_n9639 ) ;
 assign n_n7587 = ( (~ preset)  &  n_n7588  &  (~ nrq3_19) ) | ( (~ preset)  &  nrq3_19  &  n_n9619 ) ;
 assign n_n9122 = ( (~ preset)  &  n_n9123 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n9158 = ( wire3199 ) | ( (~ ndn3_28)  &  nen3_28  &  wire2406 ) ;
 assign n_n8859 = ( wire3197 ) | ( nen3_36  &  (~ ndn3_36)  &  wire2405 ) ;
 assign n_n8043 = ( wire3195 ) | ( wire3196 ) ;
 assign n_n7727 = ( wire3193 ) | ( wire2367  &  n_n9627 ) ;
 assign n_n8722 = ( wire3191 ) | ( wire3192 ) ;
 assign n_n7399 = ( wire3189 ) | ( wire2367  &  n_n9564 ) ;
 assign n_n9354 = ( wire3187 ) | ( wire3188 ) ;
 assign n_n7211 = ( wire3185 ) | ( n_n9353  &  wire2429  &  n_n9639 ) ;
 assign n_n8469 = ( wire3183 ) | ( wire2369  &  (~ n_n7311)  &  n_n7544 ) | ( wire2369  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n7312 = ( (~ preset)  &  n_n8571  &  (~ nrq2_9) ) ;
 assign n_n8795 = ( (~ preset)  &  n_n8796  &  (~ nrq2_9) ) ;
 assign n_n9116 = ( (~ preset)  &  (~ ngfdn_3)  &  nen3_36 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_36 ) ;
 assign n_n7989 = ( wire3179 ) | ( n_n8354  &  wire2436  &  n_n9639 ) ;
 assign n_n8780 = ( wire3177 ) | ( wire3178 ) ;
 assign n_n8816 = ( (~ preset)  &  n_n8817 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n9111 = ( (~ preset)  &  n_n9160 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n9091 = ( wire3171 ) | ( n_n8449  &  wire2429  &  n_n9639 ) ;
 assign n_n6938 = ( (~ preset)  &  n_n8513  &  (~ ndn_latch3_29) ) | ( (~ preset)  &  ndn_latch3_29  &  n_n9633 ) ;
 assign n_n8212 = ( wire3167 ) | ( wire3168 ) ;
 assign n_n7593 = ( wire3165 ) | ( ndn3_25  &  (~ ndn3_26)  &  wire2404 ) ;
 assign n_n8686 = ( wire16766 ) | ( (~ preset)  &  n_n9284  &  (~ n_n7274) ) ;
 assign n_n7836 = ( wire3157 ) | ( wire3158 ) ;
 assign n_n6939 = ( wire3155 ) | ( (~ ndn3_29)  &  ndn3_28  &  wire2408 ) ;
 assign n_n9202 = ( (~ preset)  &  n_n9203  &  (~ ndn_latch3_26) ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9633 ) ;
 assign n_n7113 = ( (~ preset)  &  n_n7655  &  (~ ndn_latch3_7) ) | ( (~ preset)  &  ndn_latch3_7  &  n_n9627 ) ;
 assign n_n8945 = ( (~ preset)  &  n_n8946 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n7051 = ( (~ preset)  &  n_n7052 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n9614 = ( (~ preset)  &  n_n9616  &  ndn_latch3_26 ) | ( (~ preset)  &  n_n9615  &  (~ ndn_latch3_26) ) ;
 assign n_n8472 = ( wire3143 ) | ( (~ ndn3_25)  &  ndn3_22  &  wire2408 ) ;
 assign n_n6935 = ( (~ preset)  &  n_n7741  &  (~ nrq3_16) ) | ( (~ preset)  &  nrq3_16  &  n_n9564 ) ;
 assign n_n7237 = ( wire3139 ) | ( wire3140 ) ;
 assign n_n7204 = ( (~ preset)  &  n_n7912  &  (~ nrq3_18) ) | ( (~ preset)  &  nrq3_18  &  n_n9633 ) ;
 assign n_n7525 = ( wire3135 ) | ( n_n7098  &  n_n9581 ) ;
 assign n_n9020 = ( (~ preset)  &  n_n9021  &  (~ nrq3_16) ) | ( (~ preset)  &  nrq3_16  &  n_n9619 ) ;
 assign n_n7780 = ( wire3131 ) | ( wire3132 ) ;
 assign n_n6931 = ( wire3129 ) | ( nen3_16  &  (~ ndn3_16)  &  wire2408 ) ;
 assign n_n7107 = ( wire3127 ) | ( wire3128 ) ;
 assign n_n7489 = ( wire3125 ) | ( wire3126 ) ;
 assign n_n7265 = ( wire3123 ) | ( ndn3_9  &  (~ ndn3_11)  &  wire2402 ) ;
 assign n_n8546 = ( wire3121 ) | ( wire3122 ) ;
 assign n_n7046 = ( (~ preset)  &  n_n7694  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9619 ) ;
 assign n_n8220 = ( wire3117 ) | ( n_n9448  &  wire2427  &  n_n9639 ) ;
 assign n_n7396 = ( wire3113 ) | ( wire3114 ) ;
 assign n_n7899 = ( (~ preset)  &  n_n7935  &  (~ ndn_latch3_7) ) | ( (~ preset)  &  ndn_latch3_7  &  n_n9633 ) ;
 assign n_n9229 = ( wire3107 ) | ( wire3108 ) ;
 assign n_n7515 = ( (~ preset)  &  n_n7701  &  (~ nrq2_9) ) ;
 assign n_n6929 = ( (~ preset)  &  n_n7510  &  (~ nrq3_18) ) | ( (~ preset)  &  nrq3_18  &  n_n9627 ) ;
 assign n_n6917 = ( (~ preset)  &  n_n7627  &  (~ nrq2_9) ) ;
 assign n_n8501 = ( wire3101 ) | ( wire3102 ) ;
 assign n_n8432 = ( (~ preset)  &  n_n8516  &  (~ ndn_latch3_12) ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9633 ) ;
 assign n_n7631 = ( (~ preset)  &  n_n7913  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9633 ) ;
 assign n_n9038 = ( wire3095 ) | ( n_n9284  &  wire2431  &  n_n9639 ) ;
 assign n_n7410 = ( (~ preset)  &  n_n7411 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n7326 = ( wire3091 ) | ( (~ ndn3_27)  &  ndn3_26  &  wire2405 ) ;
 assign n_n7134 = ( wire3087 ) | ( wire3088 ) ;
 assign n_n7068 = ( wire3085 ) | ( wire3086 ) ;
 assign n_n8616 = ( wire3081 ) | ( wire3082 ) ;
 assign n_n7241 = ( (~ preset)  &  n_n7242 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8229 = ( (~ preset)  &  n_n8230 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n9293 = ( (~ preset)  &  n_n9294  &  (~ nrq2_9) ) ;
 assign n_n8248 = ( wire3075 ) | ( wire2368  &  n_n9627 ) ;
 assign n_n8971 = ( (~ preset)  &  n_n8972  &  (~ nrq2_9) ) ;
 assign n_n7073 = ( wire3073 ) | ( wire3074 ) ;
 assign n_n7492 = ( (~ preset)  &  n_n7493 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n8289 = ( (~ preset)  &  n_n8290 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7184 = ( wire3065 ) | ( wire3066 ) | ( wire3067 ) | ( wire3068 ) ;
 assign n_n7162 = ( (~ preset)  &  n_n7769  &  (~ nrq2_9) ) ;
 assign n_n7490 = ( (~ preset)  &  n_n7491 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n8291 = ( wire3061 ) | ( wire3062 ) ;
 assign n_n8731 = ( wire3059 ) | ( wire3060 ) ;
 assign n_n8046 = ( (~ preset)  &  n_n8047 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n9628 = ( wire3055 ) | ( wire3056 ) ;
 assign n_n6918 = ( wire3053 ) | ( ndn3_29  &  (~ ndn3_32)  &  wire2405 ) ;
 assign n_n9507 = ( wire3051 ) | ( wire3052 ) ;
 assign n_n9154 = ( wire3049 ) | ( wire2371  &  n_n9616 ) ;
 assign n_n7377 = ( (~ preset)  &  n_n8528  &  (~ nrq2_9) ) ;
 assign n_n8994 = ( (~ preset)  &  (~ nsr3_37) ) ;
 assign n_n7690 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_42 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_40 ) ;
 assign n_n7608 = ( (~ preset)  &  n_n9358  &  (~ nrq2_9) ) ;
 assign n_n8184 = ( wire3045 ) | ( wire3046 ) ;
 assign n_n7529 = ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_30) ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_28 ) ;
 assign n_n8838 = ( wire3041 ) | ( (~ ndn3_28)  &  nen3_28  &  wire2404 ) ;
 assign n_n7902 = ( (~ preset)  &  n_n7903 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n9138 = ( wire3037 ) | ( wire3038 ) ;
 assign n_n9074 = ( (~ preset)  &  n_n9075  &  (~ ndn_latch3_28) ) | ( (~ preset)  &  ndn_latch3_28  &  n_n9627 ) ;
 assign n_n7449 = ( (~ preset)  &  n_n9439  &  (~ nrq2_9) ) ;
 assign n_n6977 = ( wire3032 ) | ( wire3034 ) | ( wire16777 ) ;
 assign n_n7151 = ( wire3027 ) | ( wire3028 ) ;
 assign n_n7747 = ( wire3025 ) | ( wire3026 ) | ( n_n8798  &  wire2451 ) ;
 assign n_n7145 = ( (~ preset)  &  n_n7146 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7056 = ( wire3018 ) | ( wire3019 ) ;
 assign n_n7175 = ( (~ preset)  &  n_n7176 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n8476 = ( wire3014 ) | ( n_n8652  &  wire2421  &  n_n9639 ) ;
 assign n_n8412 = ( (~ preset)  &  n_n8514  &  (~ nrq3_19) ) | ( (~ preset)  &  nrq3_19  &  n_n9633 ) ;
 assign n_n8635 = ( wire3010 ) | ( n_n8707  &  wire2421  &  n_n9639 ) ;
 assign n_n7182 = ( (~ preset)  &  n_n7183 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8656 = ( wire3006 ) | ( n_n8419  &  wire2418  &  n_n9639 ) ;
 assign n_n8483 = ( wire3004 ) | ( wire2367  &  n_n9581 ) ;
 assign n_n6946 = ( wire3002 ) | ( n_n8557  &  wire2427  &  n_n9639 ) ;
 assign n_n7530 = ( wire3000 ) | ( wire3001 ) ;
 assign n_n8534 = ( wire2998 ) | ( n_n8549  &  wire2427  &  n_n9639 ) ;
 assign n_n8618 = ( wire2994 ) | ( wire2995 ) ;
 assign n_n8908 = ( wire2992 ) | ( n_n8449  &  wire2427  &  n_n9639 ) ;
 assign n_n7596 = ( wire2988 ) | ( wire2989 ) ;
 assign n_n9118 = ( wire2984 ) | ( wire2985 ) ;
 assign n_n7534 = ( wire2980 ) | ( wire2981 ) ;
 assign n_n8914 = ( wire2978 ) | ( wire2979 ) ;
 assign n_n8728 = ( wire2976 ) | ( wire2977 ) ;
 assign n_n8385 = ( wire2974 ) | ( wire2975 ) | ( n_n9011  &  wire2451 ) ;
 assign n_n8778 = ( wire2969 ) | ( wire2970 ) ;
 assign n_n6979 = ( wire2967 ) | ( wire2968 ) ;
 assign n_n7714 = ( wire2965 ) | ( wire2966 ) ;
 assign n_n9066 = ( wire2961 ) | ( wire2962 ) ;
 assign n_n7059 = ( (~ preset)  &  n_n9164 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n7400 = ( wire2957 ) | ( wire2958 ) ;
 assign n_n7247 = ( wire2955 ) | ( wire2956 ) ;
 assign n_n8689 = ( wire2953 ) | ( wire2954 ) ;
 assign n_n8788 = ( wire2951 ) | ( (~ ndn3_4)  &  ndn3_2  &  wire2402 ) ;
 assign n_n8553 = ( wire2949 ) | ( (~ ndn3_34)  &  nen3_34  &  wire2405 ) ;
 assign n_n7528 = ( (~ preset)  &  n_n7768  &  (~ nrq2_9) ) ;
 assign n_n7292 = ( wire2945 ) | ( wire2946 ) ;
 assign n_n8669 = ( wire2943 ) | ( wire2369  &  n_n9627 ) ;
 assign n_n8642 = ( wire2941 ) | ( wire2942 ) ;
 assign n_n6998 = ( wire2939 ) | ( n_n9434  &  wire2427  &  n_n9639 ) ;
 assign n_n8187 = ( wire2937 ) | ( wire2938 ) ;
 assign n_n7029 = ( wire2935 ) | ( wire2370  &  n_n9627 ) ;
 assign n_n9065 = ( wire2933 ) | ( n_n9638  &  wire2427  &  n_n9639 ) ;
 assign n_n7364 = ( wire2931 ) | ( wire2932 ) ;
 assign n_n8359 = ( wire2929 ) | ( wire2930 ) ;
 assign n_n9227 = ( (~ preset)  &  n_n9228 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n8919 = ( wire2925 ) | ( (~ nsr3_13)  &  (~ ndn3_15)  &  wire2405 ) ;
 assign n_n8509 = ( (~ preset)  &  n_n8510 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8837 = ( (~ preset)  &  n_n9581  &  ndn_latch3_29 ) | ( (~ preset)  &  n_n8881  &  (~ ndn_latch3_29) ) ;
 assign n_n8639 = ( wire2919 ) | ( (~ ndn3_7)  &  ndn3_4  &  wire2405 ) ;
 assign n_n9422 = ( wire2917 ) | ( wire2918 ) ;
 assign n_n8356 = ( wire2915 ) | ( wire2916 ) | ( n_n9031  &  wire2451 ) ;
 assign n_n3 = ( wire16782 ) | ( (~ nak3_13)  &  nsr3_37 ) ;
 assign n_n7447 = ( (~ preset)  &  n_n8197  &  (~ nrq2_9) ) ;
 assign n_n8467 = ( wire2909 ) | ( wire2910 ) ;
 assign n_n7120 = ( wire2907 ) | ( wire2908 ) ;
 assign n_n7482 = ( wire2903 ) | ( wire2904 ) ;
 assign n_n7232 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_42 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_44 ) ;
 assign n_n8500 = ( wire2897 ) | ( wire2898 ) ;
 assign n_n7351 = ( wire2895 ) | ( n_n9448  &  wire2436  &  n_n9639 ) ;
 assign n_n8038 = ( wire2891 ) | ( wire2892 ) ;
 assign n_n8814 = ( (~ preset)  &  (~ pdn)  &  nsr1_2 ) | ( (~ preset)  &  (~ pdn)  &  nlc1_2 ) ;
 assign n_n8407 = ( wire2885 ) | ( wire2886 ) ;
 assign n_n8576 = ( (~ preset)  &  n_n8577  &  (~ nrq2_9) ) ;
 assign n_n7078 = ( (~ preset)  &  n_n7079 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8827 = ( (~ preset)  &  n_n8828  &  (~ ndn_latch3_29) ) | ( (~ preset)  &  ndn_latch3_29  &  n_n9627 ) ;
 assign n_n8767 = ( wire2879 ) | ( n_n9638  &  wire2447  &  n_n9639 ) ;
 assign n_n8585 = ( wire2875 ) | ( wire2876 ) ;
 assign n_n7900 = ( (~ preset)  &  n_n9616  &  nrq3_4 ) | ( (~ preset)  &  n_n7901  &  (~ nrq3_4) ) ;
 assign n_n8627 = ( wire2871 ) | ( wire2872 ) ;
 assign n_n7750 = ( wire2869 ) | ( wire2870 ) | ( n_n8869  &  wire2451 ) ;
 assign n_n7118 = ( (~ preset)  &  n_n9616  &  ndn_latch3_27 ) | ( (~ preset)  &  n_n7710  &  (~ ndn_latch3_27) ) ;
 assign n_n8181 = ( wire2864 ) | ( wire2865 ) | ( n_n8993  &  wire2451 ) ;
 assign n_n8062 = ( (~ preset)  &  n_n9586  &  (~ nrq3_21) ) | ( (~ preset)  &  nrq3_21  &  n_n9633 ) ;
 assign n_n8851 = ( (~ preset)  &  n_n9616  &  ndn_latch3_25 ) | ( (~ preset)  &  n_n8852  &  (~ ndn_latch3_25) ) ;
 assign n_n6930 = ( wire2857 ) | ( (~ ndn3_17)  &  ndn3_16  &  wire2404 ) ;
 assign n_n8010 = ( wire2855 ) | ( wire2856 ) ;
 assign n_n7716 = ( (~ preset)  &  n_n7717 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8325 = ( wire2851 ) | ( n_n8821  &  wire2421  &  n_n9639 ) ;
 assign n_n7193 = ( (~ preset)  &  n_n9163 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n8343 = ( wire2847 ) | ( n_n8557  &  wire2431  &  n_n9639 ) ;
 assign n_n8295 = ( wire2845 ) | ( wire2846 ) ;
 assign n_n8115 = ( wire2841 ) | ( wire2842 ) ;
 assign n_n8266 = ( wire2837 ) | ( wire2838 ) ;
 assign n_n7563 = ( wire2835 ) | ( wire2836 ) ;
 assign n_n9060 = ( wire2833 ) | ( n_n8652  &  wire2423  &  n_n9639 ) ;
 assign n_n9206 = ( wire2831 ) | ( (~ ndn3_25)  &  ndn3_22  &  wire2406 ) ;
 assign n_n7278 = ( wire2827 ) | ( wire2828 ) ;
 assign n_n9080 = ( wire2825 ) | ( n_n9512  &  wire2423  &  n_n9639 ) ;
 assign n_n6909 = ( wire2823 ) | ( wire2824 ) ;
 assign n_n8726 = ( wire2821 ) | ( (~ ndn3_17)  &  ndn3_16  &  wire2402 ) ;
 assign n_n7672 = ( wire2819 ) | ( wire2820 ) ;
 assign n_n7329 = ( (~ preset)  &  n_n7330 ) | ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign n_n8965 = ( wire2813 ) | ( wire2814 ) ;
 assign n_n7841 = ( wire2811 ) | ( wire2812 ) ;
 assign n_n8283 = ( wire2809 ) | ( wire2810 ) | ( n_n8847  &  wire2451 ) ;
 assign n_n9374 = ( wire2806 ) | ( wire2807 ) ;
 assign n_n7171 = ( (~ preset)  &  n_n7553  &  (~ nrq3_4) ) | ( (~ preset)  &  nrq3_4  &  n_n9564 ) ;
 assign n_n6927 = ( (~ preset)  &  n_n9292  &  (~ nrq2_9) ) ;
 assign n_n7071 = ( (~ preset)  &  n_n7464  &  (~ nrq3_39) ) | ( (~ preset)  &  nrq3_39  &  n_n9619 ) ;
 assign n_n8144 = ( wire2800 ) | ( wire2801 ) ;
 assign n_n8437 = ( wire2798 ) | ( wire2799 ) ;
 assign n_n6999 = ( wire2796 ) | ( n_n9434  &  wire2431  &  n_n9639 ) ;
 assign n_n8117 = ( (~ preset)  &  n_n8118  &  (~ nrq2_9) ) ;
 assign n_n7610 = ( wire2794 ) | ( wire2371  &  n_n9627 ) ;
 assign n_n9238 = ( wire2792 ) | ( wire2369  &  n_n9564 ) ;
 assign n_n9236 = ( wire2790 ) | ( wire2369  &  (~ n_n7869)  &  n_n8028 ) | ( wire2369  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n6913 = ( wire2788 ) | ( n_n9434  &  wire2436  &  n_n9639 ) ;
 assign n_n9443 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_2 ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_2 ) ;
 assign n_n9521 = ( wire2784 ) | ( n_n8652  &  wire2447  &  n_n9639 ) ;
 assign n_n7518 = ( wire2782 ) | ( wire2783 ) ;
 assign n_n7433 = ( wire2780 ) | ( wire2781 ) ;
 assign n_n8664 = ( (~ preset)  &  n_n8665 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n8318 = ( wire2776 ) | ( wire2777 ) ;
 assign n_n8301 = ( wire2774 ) | ( wire2775 ) ;
 assign n_n7020 = ( wire2772 ) | ( wire2773 ) ;
 assign n_n8133 = ( (~ preset)  &  n_n9581  &  nrq3_36 ) | ( (~ preset)  &  n_n9173  &  (~ nrq3_36) ) ;
 assign n_n8896 = ( wire2768 ) | ( wire2769 ) ;
 assign n_n7149 = ( (~ preset)  &  n_n7150 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n9454 = ( wire2764 ) | ( nen3_36  &  (~ ndn3_36)  &  wire2406 ) ;
 assign n_n8370 = ( wire2762 ) | ( wire2763 ) ;
 assign n_n8 = ( wire16786 ) | ( (~ ndn3_17)  &  nsr3_20 ) ;
 assign n_n7047 = ( (~ preset)  &  n_n8271  &  (~ nrq2_9) ) ;
 assign n_n8836 = ( wire2757 ) | ( wire2758 ) ;
 assign n_n7443 = ( wire2755 ) | ( wire2370  &  n_n9633 ) ;
 assign n_n7158 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_39 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_40 ) ;
 assign n_n7128 = ( wire2751 ) | ( wire2752 ) ;
 assign n_n7676 = ( wire2749 ) | ( (~ ndn3_4)  &  ndn3_2  &  wire2406 ) ;
 assign n_n8101 = ( wire2747 ) | ( wire2748 ) ;
 assign n_n9224 = ( wire2743 ) | ( wire2744 ) ;
 assign n_n8461 = ( (~ preset)  &  n_n9581  &  nrq3_21 ) | ( (~ preset)  &  n_n8462  &  (~ nrq3_21) ) ;
 assign n_n8087 = ( wire2737 ) | ( wire2738 ) ;
 assign n_n9024 = ( wire2735 ) | ( wire2736 ) ;
 assign n_n8178 = ( (~ preset)  &  n_n9289  &  (~ nrq2_9) ) ;
 assign n_n7660 = ( (~ preset)  &  n_n7661  &  (~ nrq3_15) ) | ( (~ preset)  &  nrq3_15  &  n_n9627 ) ;
 assign n_n8107 = ( wire2731 ) | ( wire2732 ) ;
 assign n_n8920 = ( (~ preset)  &  n_n8921 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7858 = ( wire2727 ) | ( (~ ndn3_28)  &  nen3_28  &  wire2408 ) ;
 assign n_n7731 = ( wire2725 ) | ( n_n9448  &  wire2429  &  n_n9639 ) ;
 assign n_n7427 = ( wire2721 ) | ( wire2722 ) ;
 assign n_n9519 = ( wire2719 ) | ( wire2367  &  (~ n_n7311)  &  n_n7544 ) | ( wire2367  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n6964 = ( wire2717 ) | ( wire2718 ) ;
 assign n_n7677 = ( wire2715 ) | ( wire2716 ) ;
 assign n_n7222 = ( wire2713 ) | ( n_n8449  &  wire2447  &  n_n9639 ) ;
 assign n_n7679 = ( wire2711 ) | ( wire2712 ) ;
 assign n_n8840 = ( wire2709 ) | ( n_n8419  &  wire2447  &  n_n9639 ) ;
 assign n_n7335 = ( (~ preset)  &  n_n7336 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n7197 = ( wire2705 ) | ( (~ ndn3_17)  &  ndn3_16  &  wire2408 ) ;
 assign n_n7754 = ( wire2703 ) | ( wire2704 ) ;
 assign n_n7195 = ( wire2701 ) | ( wire2702 ) ;
 assign n_n8769 = ( wire2697 ) | ( wire2698 ) ;
 assign n_n8422 = ( (~ preset)  &  n_n8423 ) | ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign n_n7085 = ( (~ preset)  &  n_n9616  &  nrq3_15 ) | ( (~ preset)  &  n_n7763  &  (~ nrq3_15) ) ;
 assign n_n9524 = ( wire2691 ) | ( n_n8419  &  wire2427  &  n_n9639 ) ;
 assign n_n8032 = ( wire2687 ) | ( wire2688 ) ;
 assign n_n7533 = ( wire2683 ) | ( wire2684 ) ;
 assign n_n7426 = ( wire2679 ) | ( wire2680 ) ;
 assign n_n9231 = ( wire2675 ) | ( wire2676 ) ;
 assign n_n7257 = ( wire2673 ) | ( (~ ndn3_9)  &  ndn3_7  &  wire2408 ) ;
 assign n_n9562 = ( (~ preset)  &  n_n9563  &  (~ nrq3_9) ) | ( (~ preset)  &  nrq3_9  &  n_n9564 ) ;
 assign n_n8671 = ( (~ preset)  &  n_n8672 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n7106 = ( (~ preset)  &  n_n7346  &  (~ nrq3_39) ) | ( (~ preset)  &  nrq3_39  &  n_n9627 ) ;
 assign n_n7008 = ( wire2665 ) | ( n_n8821  &  wire2423  &  n_n9639 ) ;
 assign n_n8755 = ( (~ preset)  &  n_n8756  &  (~ nrq2_9) ) ;
 assign n_n8640 = ( (~ preset)  &  n_n8641  &  (~ nrq3_4) ) | ( (~ preset)  &  nrq3_4  &  n_n9627 ) ;
 assign n_n8191 = ( wire2659 ) | ( wire2660 ) ;
 assign n_n8057 = ( wire2657 ) | ( ndn3_17  &  (~ ndn3_18)  &  wire2402 ) ;
 assign n_n7439 = ( wire2655 ) | ( wire2656 ) | ( n_n8561  &  wire2451 ) ;
 assign n_n9305 = ( (~ preset)  &  n_n9306 ) | ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign n_n6928 = ( (~ preset)  &  n_n9165 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n8848 = ( wire2648 ) | ( wire2649 ) ;
 assign n_n9209 = ( (~ preset)  &  n_n9210  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9616 ) ;
 assign n_n8122 = ( (~ preset)  &  ndn2_2  &  (~ ngfdn_2) ) ;
 assign n_n7254 = ( (~ preset)  &  n_n7342  &  (~ nrq3_19) ) | ( (~ preset)  &  nrq3_19  &  n_n9627 ) ;
 assign n_n8050 = ( wire2640 ) | ( wire2641 ) ;
 assign n_n7135 = ( wire2638 ) | ( wire2371  &  (~ n_n7869)  &  n_n8028 ) | ( wire2371  &  n_n7869  &  (~ n_n8028) ) ;
 assign n_n7081 = ( wire2634 ) | ( wire2635 ) ;
 assign n_n9005 = ( (~ preset)  &  n_n9006 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7407 = ( wire2630 ) | ( n_n8652  &  wire2418  &  n_n9639 ) ;
 assign n_n7904 = ( (~ preset)  &  n_n7905 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n7030 = ( (~ preset)  &  n_n9166 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n7064 = ( (~ preset)  &  n_n7065 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n8211 = ( (~ preset)  &  n_n9581  &  ndn_latch3_28 ) | ( (~ preset)  &  n_n9490  &  (~ ndn_latch3_28) ) ;
 assign n_n7023 = ( (~ preset)  &  n_n7024 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n7585 = ( (~ preset)  &  n_n7586 ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign n_n8415 = ( wire2614 ) | ( wire2615 ) ;
 assign n_n8166 = ( wire2612 ) | ( wire2613 ) ;
 assign n_n8140 = ( (~ preset)  &  n_n8141  &  (~ nrq2_9) ) ;
 assign n_n7446 = ( (~ preset)  &  n_n7853  &  (~ nrq2_9) ) ;
 assign n_n8120 = ( (~ preset)  &  n_n8121 ) | ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign n_n8162 = ( wire2606 ) | ( wire2607 ) ;
 assign n_n8337 = ( (~ preset)  &  n_n9496  &  (~ ndn_latch3_12) ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9581 ) ;
 assign n_n8194 = ( (~ preset)  &  n_n8195 ) | ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign n_n9515 = ( (~ preset)  &  n_n9616  &  nrq3_34 ) | ( (~ preset)  &  n_n9516  &  (~ nrq3_34) ) ;
 assign n_n9076 = ( wire2598 ) | ( (~ ndn3_27)  &  ndn3_26  &  wire2404 ) ;
 assign n_n8363 = ( (~ preset)  &  n_n9436  &  (~ nrq2_9) ) ;
 assign n_n8773 = ( wire2596 ) | ( wire2597 ) ;
 assign n_n7089 = ( wire2594 ) | ( wire2595 ) ;
 assign n_n7840 = ( wire2590 ) | ( wire2591 ) | ( wire2592 ) | ( wire2593 ) ;
 assign n_n7321 = ( wire2588 ) | ( n_n9416  &  wire2436  &  n_n9639 ) ;
 assign n_n8873 = ( wire2586 ) | ( ndn3_9  &  (~ ndn3_11)  &  wire2405 ) ;
 assign n_n7745 = ( wire2584 ) | ( n_n9353  &  wire2423  &  n_n9639 ) ;
 assign n_n7001 = ( (~ preset)  &  n_n7770  &  (~ nrq2_9) ) ;
 assign n_n6959 = ( (~ preset)  &  ndn3_29  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_32 ) ;
 assign n_n7196 = ( wire2580 ) | ( wire2581 ) ;
 assign n_n8205 = ( wire2578 ) | ( wire2371  &  n_n9581 ) ;
 assign n_n7367 = ( wire2576 ) | ( wire2368  &  n_n9633 ) ;
 assign n_n8818 = ( wire2572 ) | ( wire2573 ) ;
 assign n_n7110 = ( wire2570 ) | ( wire2571 ) ;
 assign n_n7804 = ( wire2568 ) | ( wire2569 ) ;
 assign n_n8494 = ( (~ preset)  &  (~ nsr3_38) ) ;
 assign n_n7206 = ( wire2564 ) | ( wire2565 ) ;
 assign n_n8872 = ( (~ preset)  &  n_n9179  &  (~ nrq3_11) ) | ( (~ preset)  &  nrq3_11  &  n_n9581 ) ;
 assign n_n8364 = ( (~ preset)  &  n_n9357  &  (~ nrq2_9) ) ;
 assign n_n8496 = ( wire2558 ) | ( wire2559 ) ;
 assign n_n6971 = ( (~ preset)  &  n_n7628  &  (~ nrq2_9) ) ;
 assign n_n8453 = ( (~ preset)  &  n_n8454 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n7413 = ( (~ preset)  &  (~ nsr3_20) ) ;
 assign n_n9504 = ( wire2554 ) | ( n_n9448  &  wire2421  &  n_n9639 ) ;
 assign n_n8825 = ( (~ preset)  &  (~ ngfdn_3)  &  (~ nsr3_35) ) | ( (~ preset)  &  (~ ngfdn_3)  &  nen3_34 ) ;
 assign n_n9631 = ( wire2550 ) | ( wire2369  &  n_n9633 ) ;
 assign n_n7075 = ( wire2548 ) | ( wire2549 ) ;
 assign n_n7469 = ( wire2544 ) | ( wire2545 ) ;
 assign n_n8634 = ( wire2542 ) | ( wire2543 ) ;
 assign n_n9577 = ( (~ preset)  &  n_n9578 ) | ( (~ preset)  &  nrq2_9 ) ;
 assign n_n8134 = ( (~ preset)  &  n_n8135  &  (~ nrq3_34) ) | ( (~ preset)  &  nrq3_34  &  n_n9564 ) ;
 assign n_n9328 = ( (~ preset)  &  ndn3_25  &  (~ ngfdn_3) ) | ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_26 ) ;
 assign n_n7499 = ( wire2534 ) | ( wire2535 ) ;
 assign n_n6973 = ( wire2532 ) | ( wire2371  &  (~ n_n7311)  &  n_n7544 ) | ( wire2371  &  n_n7311  &  (~ n_n7544) ) ;
 assign n_n8604 = ( (~ preset)  &  n_n8605 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n9295 = ( (~ preset)  &  n_n9296  &  (~ nrq2_9) ) ;
 assign n_n7155 = ( wire2528 ) | ( wire2529 ) ;
 assign n_n7919 = ( wire2526 ) | ( n_n9638  &  wire2423  &  n_n9639 ) ;
 assign n_n8893 = ( wire2524 ) | ( wire2525 ) ;
 assign n_n7620 = ( wire2522 ) | ( nen3_39  &  (~ ndn3_39)  &  wire2406 ) ;
 assign n_n8138 = ( wire2518 ) | ( wire2519 ) ;
 assign n_n9274 = ( (~ preset)  &  n_n9275  &  (~ nrq2_9) ) ;
 assign n_n7202 = ( wire2516 ) | ( wire2517 ) ;
 assign n_n7805 = ( wire2514 ) | ( n_n9537  &  wire2423  &  n_n9639 ) ;
 assign n_n7343 = ( wire2512 ) | ( wire2513 ) ;
 assign n_n6975 = ( wire2508 ) | ( wire2509 ) ;
 assign n_n6958 = ( (~ preset)  &  n_n7629  &  (~ nrq2_9) ) ;
 assign n_n7617 = ( (~ preset)  &  (~ nsr3_14) ) ;
 assign n_n7646 = ( wire2506 ) | ( wire2371  &  (~ n_n9385)  &  n_n9384 ) | ( wire2371  &  n_n9385  &  (~ n_n9384) ) ;
 assign n_n9012 = ( (~ preset)  &  n_n9013  &  (~ nrq2_9) ) ;
 assign n_n7287 = ( wire2504 ) | ( wire2505 ) ;
 assign n_n8077 = ( wire2502 ) | ( n_n8557  &  wire2436  &  n_n9639 ) ;
 assign n_n7333 = ( (~ preset)  &  n_n9616  &  nrq3_39 ) | ( (~ preset)  &  n_n7334  &  (~ nrq3_39) ) ;
 assign n_n6957 = ( (~ preset)  &  n_n7704  &  (~ nrq2_9) ) ;
 assign n_n7496 = ( wire2498 ) | ( n_n8419  &  wire2421  &  n_n9639 ) ;
 assign n_n8525 = ( (~ preset)  &  n_n8526  &  (~ ndn_latch3_27) ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9627 ) ;
 assign n_n7795 = ( (~ preset)  &  n_n9556  &  (~ nrq2_9) ) ;
 assign n_n7851 = ( wire2494 ) | ( ndn3_9  &  (~ ndn3_11)  &  wire2406 ) ;
 assign n_n8446 = ( (~ preset)  &  n_n8447  &  (~ nrq2_9) ) ;
 assign n_n7484 = ( wire2492 ) | ( wire2493 ) ;
 assign n_n7305 = ( (~ preset)  &  n_n8570  &  (~ nrq2_9) ) ;
 assign n_n6921 = ( wire2490 ) | ( ndn3_25  &  (~ ndn3_26)  &  wire2402 ) ;
 assign n_n7191 = ( wire2488 ) | ( n_n8549  &  wire2436  &  n_n9639 ) ;
 assign n_n6926 = ( (~ preset)  &  n_n8646  &  (~ nrq2_9) ) ;
 assign n_n8489 = ( wire2484 ) | ( wire2485 ) ;
 assign n_n8947 = ( wire2482 ) | ( n_n7098  &  (~ n_n7566)  &  n_n8154 ) | ( n_n7098  &  n_n7566  &  (~ n_n8154) ) ;
 assign n_n8471 = ( wire2480 ) | ( ndn3_17  &  (~ ndn3_18)  &  wire2405 ) ;
 assign n_n8215 = ( (~ preset)  &  n_n8216 ) | ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign n_n8180 = ( (~ preset)  &  n_n9581  &  nrq3_18 ) | ( (~ preset)  &  n_n9177  &  (~ nrq3_18) ) ;
 assign n_n7295 = ( wire2474 ) | ( wire2475 ) ;
 assign n_n7437 = ( wire2472 ) | ( (~ ndn3_17)  &  ndn3_16  &  wire2405 ) ;
 assign n_n9143 = ( wire2470 ) | ( wire2471 ) ;
 assign n_n8426 = ( wire2379 ) | ( wire2382 ) ;
 assign n_n8558 = ( (~ preset)  &  n_n8858  &  (~ nrq3_39) ) | ( (~ preset)  &  nrq3_39  &  n_n9581 ) ;
 assign n_n7838 = ( wire2364 ) | ( (~ ndn3_34)  &  nen3_34  &  wire2404 ) ;
 assign wire2421 = ( (~ preset)  &  (~ ndn3_37)  &  (~ nsr3_37) ) ;
 assign wire2371 = ( (~ preset)  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign nrq3_11 = ( ndn3_9  &  (~ ndn3_11) ) ;
 assign n_n9616 = ( (~ n_n7566)  &  (~ n_n8155)  &  n_n7218 ) | ( (~ n_n8156)  &  (~ n_n8155)  &  n_n7218 ) | ( n_n8156  &  n_n8155  &  (~ n_n7218) ) | ( (~ n_n7566)  &  (~ n_n8156)  &  n_n8155  &  n_n7218 ) | ( n_n7566  &  (~ n_n8156)  &  n_n8155  &  (~ n_n7218) ) | ( n_n7566  &  n_n8156  &  (~ n_n8155)  &  (~ n_n7218) ) ;
 assign ndn_latch3_12 = ( ndn3_11  &  (~ ndn3_12) ) ;
 assign wire2405 = ( (~ preset)  &  (~ n_n9478)  &  wire5338 ) | ( (~ preset)  &  (~ n_n9478)  &  wire5339 ) | ( (~ preset)  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign ndn_latch3_26 = ( ndn3_25  &  (~ ndn3_26) ) ;
 assign nrq3_9 = ( (~ ndn3_9)  &  ndn3_7 ) ;
 assign wire2370 = ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign nrq3_39 = ( nen3_39  &  (~ ndn3_39) ) ;
 assign wire2408 = ( (~ preset)  &  (~ n_n8314)  &  wire5069 ) | ( (~ preset)  &  (~ n_n8314)  &  wire5070 ) | ( (~ preset)  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire2363 = ( (~ preset)  &  (~ n_n7306)  &  n_n9248  &  n_n9247 ) ;
 assign wire2395 = ( wire2363  &  n_n7274 ) ;
 assign wire2453 = ( n_n8549  &  n_n8522  &  n_n8579 ) | ( n_n8549  &  n_n8521  &  n_n8579 ) | ( n_n8522  &  n_n8521  &  n_n8579 ) | ( (~ n_n8549)  &  (~ n_n8522)  &  (~ n_n8579) ) | ( (~ n_n8549)  &  (~ n_n8521)  &  (~ n_n8579) ) | ( (~ n_n8522)  &  (~ n_n8521)  &  (~ n_n8579) ) ;
 assign ndn_latch3_27 = ( (~ ndn3_27)  &  ndn3_26 ) ;
 assign nrq3_34 = ( (~ ndn3_34)  &  nen3_34 ) ;
 assign wire2369 = ( (~ preset)  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire2469 = ( preset ) | ( (~ n_n9198) ) | ( (~ n_n9639)  &  n_n9197 ) ;
 assign wire2368 = ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire2436 = ( (~ preset)  &  (~ nsr3_35)  &  (~ ndn3_35) ) ;
 assign nrq3_19 = ( (~ ndn3_19)  &  nen3_19 ) ;
 assign wire2367 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22) ) ;
 assign wire2447 = ( (~ preset)  &  (~ ndn3_23)  &  (~ nsr3_23) ) ;
 assign n_n9581 = ( (~ n_n9583)  &  n_n7818  &  n_n7597 ) | ( n_n9583  &  (~ n_n8028)  &  (~ n_n7597) ) | ( n_n9583  &  (~ n_n7818)  &  (~ n_n7597) ) | ( (~ n_n9583)  &  n_n8028  &  (~ n_n7818)  &  n_n7597 ) | ( n_n9583  &  (~ n_n8028)  &  (~ n_n7818)  &  n_n7597 ) | ( (~ n_n9583)  &  n_n8028  &  n_n7818  &  (~ n_n7597) ) ;
 assign ndn_latch3_29 = ( (~ ndn3_29)  &  ndn3_28 ) ;
 assign n_n8979 = ( wire4976 ) | ( wire4977 ) | ( wire4978 ) | ( wire16484 ) ;
 assign n_n7432 = ( n_n8821  &  n_n8820 ) | ( n_n8821  &  wire16528 ) | ( n_n8820  &  wire16528 ) | ( n_n8821  &  wire16529 ) | ( n_n8820  &  wire16529 ) ;
 assign n_n8323 = ( n_n9638  &  n_n7432 ) | ( n_n9638  &  wire16483 ) | ( n_n7432  &  wire16483 ) | ( n_n9638  &  wire16484 ) | ( n_n7432  &  wire16484 ) ;
 assign wire2402 = ( (~ preset)  &  (~ n_n7939)  &  wire5311 ) | ( (~ preset)  &  (~ n_n7939)  &  wire5312 ) | ( (~ preset)  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign nrq3_4 = ( (~ ndn3_4)  &  ndn3_2 ) ;
 assign nrq3_16 = ( nen3_16  &  (~ ndn3_16) ) ;
 assign nrq3_36 = ( nen3_36  &  (~ ndn3_36) ) ;
 assign nrq3_18 = ( ndn3_17  &  (~ ndn3_18) ) ;
 assign wire2404 = ( (~ preset)  &  (~ n_n8865)  &  wire4672 ) | ( (~ preset)  &  (~ n_n8865)  &  wire4673 ) | ( (~ preset)  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign ndn_latch3_7 = ( (~ ndn3_7)  &  ndn3_4 ) ;
 assign ndn_latch3_32 = ( ndn3_29  &  (~ ndn3_32) ) ;
 assign nrq3_15 = ( (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign nrq3_17 = ( (~ ndn3_17)  &  ndn3_16 ) ;
 assign wire2431 = ( (~ preset)  &  (~ ndn3_13)  &  (~ nsr3_13) ) ;
 assign n_n7378 = ( (~ pdn)  &  (~ nsr1_2) ) | ( pdn  &  (~ ndn1_4) ) ;
 assign nrq3_21 = ( ndn3_19  &  (~ ndn3_21) ) ;
 assign wire2418 = ( (~ preset)  &  (~ nsr3_20)  &  (~ ndn3_20) ) ;
 assign n_n9619 = ( (~ n_n7997)  &  n_n9258  &  n_n9587 ) | ( n_n7997  &  (~ n_n8019)  &  (~ n_n9587) ) | ( n_n7997  &  (~ n_n9258)  &  (~ n_n9587) ) | ( (~ n_n7997)  &  n_n8019  &  (~ n_n9258)  &  n_n9587 ) | ( n_n7997  &  (~ n_n8019)  &  (~ n_n9258)  &  n_n9587 ) | ( (~ n_n7997)  &  n_n8019  &  n_n9258  &  (~ n_n9587) ) ;
 assign wire2406 = ( (~ preset)  &  (~ n_n8320)  &  wire5184 ) | ( (~ preset)  &  (~ n_n8320)  &  wire5185 ) | ( (~ preset)  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign ndn_latch3_25 = ( (~ ndn3_25)  &  ndn3_22 ) ;
 assign wire2423 = ( (~ preset)  &  (~ nsr3_38)  &  (~ ndn3_38) ) ;
 assign wire2427 = ( (~ preset)  &  (~ nsr3_14)  &  (~ ndn3_14) ) ;
 assign ndn_latch3_28 = ( (~ ndn3_28)  &  nen3_28 ) ;
 assign n_n8880 = ( wire4955 ) | ( wire4956 ) | ( wire4957 ) | ( wire16489 ) ;
 assign n_n8431 = ( n_n9512  &  n_n8733 ) | ( n_n9512  &  wire16493 ) | ( n_n8733  &  wire16493 ) | ( n_n9512  &  wire16494 ) | ( n_n8733  &  wire16494 ) ;
 assign n_n8783 = ( n_n9434  &  n_n8431 ) | ( n_n9434  &  wire16488 ) | ( n_n8431  &  wire16488 ) | ( n_n9434  &  wire16489 ) | ( n_n8431  &  wire16489 ) ;
 assign wire2429 = ( (~ preset)  &  (~ ndn3_30)  &  (~ nsr3_30) ) ;
 assign n_n9056 = ( wire15923 ) | ( wire15924 ) ;
 assign wire2451 = ( (~ preset)  &  n_n9639  &  n_n8667 ) | ( (~ preset)  &  (~ n_n8667)  &  (~ n_n7274) ) ;
 assign n_n8403 = ( n_n8631  &  n_n8561 ) | ( n_n8631  &  n_n8342 ) | ( (~ n_n8631)  &  (~ n_n8561)  &  (~ n_n8342) ) ;
 assign n_n8630 = ( wire15929 ) | ( wire15930 ) ;
 assign ngfdn_2 = ( preset_0_0_  &  nsr1_2  &  (~ nlc1_2) ) ;
 assign n_n9246 = ( (~ n_n8538)  &  (~ n_n8606)  &  wire16670  &  wire16671 ) ;
 assign n_n9564 = ( (~ n_n8953)  &  n_n9040  &  n_n9307 ) | ( (~ n_n9384)  &  n_n8953  &  (~ n_n9307) ) | ( n_n8953  &  (~ n_n9040)  &  (~ n_n9307) ) | ( (~ n_n9384)  &  n_n8953  &  (~ n_n9040)  &  n_n9307 ) | ( n_n9384  &  (~ n_n8953)  &  (~ n_n9040)  &  n_n9307 ) | ( n_n9384  &  (~ n_n8953)  &  n_n9040  &  (~ n_n9307) ) ;
 assign n_n9633 = ( (~ n_n7543)  &  n_n8126  &  n_n8125 ) | ( n_n7543  &  (~ n_n7544)  &  (~ n_n8125) ) | ( n_n7543  &  (~ n_n8126)  &  (~ n_n8125) ) | ( (~ n_n7543)  &  n_n7544  &  (~ n_n8126)  &  n_n8125 ) | ( n_n7543  &  (~ n_n7544)  &  (~ n_n8126)  &  n_n8125 ) | ( (~ n_n7543)  &  n_n7544  &  n_n8126  &  (~ n_n8125) ) ;
 assign n_n8522 = ( wire4997 ) | ( wire4998 ) | ( wire4999 ) | ( wire16474 ) ;
 assign n_n8521 = ( n_n8449  &  n_n8448 ) | ( n_n8449  &  wire16478 ) | ( n_n8448  &  wire16478 ) | ( n_n8449  &  wire16479 ) | ( n_n8448  &  wire16479 ) ;
 assign n_n8538 = ( n_n8913  &  n_n8964 ) | ( n_n8964  &  n_n8493 ) | ( (~ n_n8913)  &  (~ n_n8964)  &  (~ n_n8493) ) ;
 assign n_n8963 = ( wire15935 ) | ( wire15936 ) ;
 assign n_n8537 = ( n_n8652  &  wire16498 ) | ( n_n8652  &  wire16499 ) ;
 assign n_n8653 = ( wire4927 ) | ( wire4928 ) | ( wire4929 ) | ( wire16499 ) ;
 assign n_n8706 = ( n_n9284  &  n_n8537 ) | ( n_n9284  &  wire16503 ) | ( n_n8537  &  wire16503 ) | ( n_n9284  &  wire16504 ) | ( n_n8537  &  wire16504 ) ;
 assign n_n8484 = ( n_n8707  &  n_n8706 ) | ( n_n8707  &  wire16508 ) | ( n_n8706  &  wire16508 ) | ( n_n8707  &  wire16509 ) | ( n_n8706  &  wire16509 ) ;
 assign n_n8708 = ( wire4918 ) | ( wire4919 ) | ( wire4920 ) | ( wire16509 ) ;
 assign n_n8418 = ( n_n8354  &  n_n8353 ) | ( n_n8354  &  wire16538 ) | ( n_n8353  &  wire16538 ) | ( n_n8354  &  wire16539 ) | ( n_n8353  &  wire16539 ) ;
 assign n_n8353 = ( n_n9448  &  n_n8323 ) | ( n_n9448  &  wire16533 ) | ( n_n8323  &  wire16533 ) | ( n_n9448  &  wire16534 ) | ( n_n8323  &  wire16534 ) ;
 assign n_n8355 = ( wire4886 ) | ( wire4887 ) | ( wire4888 ) | ( wire16539 ) ;
 assign n_n9356 = ( wire15941 ) | ( wire15942 ) ;
 assign n_n8734 = ( wire4948 ) | ( wire4949 ) | ( wire4950 ) | ( wire16494 ) ;
 assign n_n8733 = ( n_n9353  &  n_n8484 ) | ( n_n9353  &  wire16513 ) | ( n_n8484  &  wire16513 ) | ( n_n9353  &  wire16514 ) | ( n_n8484  &  wire16514 ) ;
 assign wire2460 = ( n_n8734 ) | ( n_n9353  &  n_n8484 ) | ( n_n9353  &  n_n8807 ) | ( n_n8484  &  n_n8807 ) ;
 assign n_n8784 = ( wire4962 ) | ( wire4963 ) | ( wire4964 ) | ( wire16519 ) ;
 assign n_n8373 = ( n_n9416  &  n_n8783 ) | ( n_n9416  &  wire16518 ) | ( n_n8783  &  wire16518 ) | ( n_n9416  &  wire16519 ) | ( n_n8783  &  wire16519 ) ;
 assign n_n7864 = ( wire15953 ) | ( wire15954 ) ;
 assign n_n8876 = ( (~ n_n8603)  &  n_n8923 ) | ( n_n8923  &  n_n8798 ) | ( n_n8603  &  (~ n_n8923)  &  (~ n_n8798) ) ;
 assign n_n9072 = ( wire15959 ) | ( wire15960 ) ;
 assign n_n7787 = ( wire15965 ) | ( wire15966 ) ;
 assign n_n8976 = ( n_n8911  &  n_n8978 ) | ( n_n8933  &  n_n8978 ) | ( n_n8978  &  n_n8932 ) | ( (~ n_n8911)  &  (~ n_n8933)  &  (~ n_n8978)  &  (~ n_n8932) ) ;
 assign n_n7637 = ( n_n9034  &  n_n9031 ) | ( n_n9034  &  n_n8993 ) | ( n_n9034  &  n_n8204 ) | ( (~ n_n9034)  &  (~ n_n9031)  &  (~ n_n8993)  &  (~ n_n8204) ) ;
 assign n_n9553 = ( wire15971 ) | ( wire15972 ) ;
 assign n_n9627 = ( (~ wire16245)  &  (~ wire16246)  &  wire16262 ) | ( (~ wire16245)  &  (~ wire16246)  &  wire16263 ) | ( wire16245  &  (~ wire16262)  &  (~ wire16263) ) | ( wire16246  &  (~ wire16262)  &  (~ wire16263) ) ;
 assign n_n8450 = ( wire4990 ) | ( wire4991 ) | ( wire4992 ) | ( wire16479 ) ;
 assign n_n8448 = ( n_n8419  &  n_n8418 ) | ( n_n8419  &  wire16543 ) | ( n_n8418  &  wire16543 ) | ( n_n8419  &  wire16544 ) | ( n_n8418  &  wire16544 ) ;
 assign n_n8324 = ( wire4983 ) | ( wire4984 ) | ( wire4985 ) | ( wire16534 ) ;
 assign n_n8820 = ( n_n9537  &  n_n8373 ) | ( n_n9537  &  wire16523 ) | ( n_n8373  &  wire16523 ) | ( n_n9537  &  wire16524 ) | ( n_n8373  &  wire16524 ) ;
 assign n_n8936 = ( wire4969 ) | ( wire4970 ) | ( wire4971 ) | ( wire16524 ) ;
 assign n_n8740 = ( wire4934 ) | ( wire4935 ) | ( wire4936 ) | ( wire16504 ) ;
 assign n_n8822 = ( wire4899 ) | ( wire4900 ) | ( wire4901 ) | ( wire16529 ) ;
 assign n_n8807 = ( wire4941 ) | ( wire4942 ) | ( wire4943 ) | ( wire16514 ) ;
 assign n_n9216 = ( wire15977 ) | ( wire15978 ) ;
 assign n_n8606 = ( n_n8913  &  n_n9011 ) | ( n_n8964  &  n_n9011 ) | ( n_n9011  &  n_n8493 ) | ( (~ n_n8913)  &  (~ n_n8964)  &  (~ n_n9011)  &  (~ n_n8493) ) ;
 assign n_n9010 = ( wire15983 ) | ( wire15984 ) ;
 assign n_n8823 = ( wire15989 ) | ( wire15990 ) ;
 assign n_n9029 = ( n_n9031  &  n_n8993 ) | ( n_n9031  &  n_n8204 ) | ( (~ n_n9031)  &  (~ n_n8993)  &  (~ n_n8204) ) ;
 assign n_n9288 = ( wire15995 ) | ( wire15996 ) ;
 assign n_n9114 = ( (~ n_n8603)  &  n_n8869 ) | ( n_n8923  &  n_n8869 ) | ( n_n8798  &  n_n8869 ) | ( n_n8603  &  (~ n_n8923)  &  (~ n_n8798)  &  (~ n_n8869) ) ;
 assign n_n9435 = ( wire16001 ) | ( wire16002 ) ;
 assign n_n9152 = ( n_n8631  &  n_n8847 ) | ( n_n8847  &  n_n8561 ) | ( n_n8847  &  n_n8342 ) | ( (~ n_n8631)  &  (~ n_n8847)  &  (~ n_n8561)  &  (~ n_n8342) ) ;
 assign n_n8846 = ( wire16007 ) | ( wire16008 ) ;
 assign nen3_2 = ( nsr1_2  &  n_n7476  &  nlc1_2 ) | ( (~ preset_0_0_)  &  nsr1_2  &  (~ nlc1_2) ) ;
 assign n_n8806 = ( wire16013 ) | ( wire16014 ) ;
 assign n_n8420 = ( wire4877 ) | ( wire4878 ) | ( wire4879 ) | ( wire16544 ) ;
 assign n_n7543 = ( (~ wire16639)  &  (~ wire16640)  &  wire16656 ) | ( (~ wire16639)  &  (~ wire16640)  &  wire16657 ) | ( wire16639  &  (~ wire16656)  &  (~ wire16657) ) | ( wire16640  &  (~ wire16656)  &  (~ wire16657) ) ;
 assign n_n8694 = ( (~ n_n7306)  &  n_n9248  &  n_n9247 ) ;
 assign n_n9385 = ( (~ wire16212)  &  (~ wire16213)  &  wire16229 ) | ( (~ wire16212)  &  (~ wire16213)  &  wire16230 ) | ( wire16212  &  (~ wire16229)  &  (~ wire16230) ) | ( wire16213  &  (~ wire16229)  &  (~ wire16230) ) ;
 assign n_n9384 = ( wire16245  &  wire16262 ) | ( wire16246  &  wire16262 ) | ( wire16245  &  wire16263 ) | ( wire16246  &  wire16263 ) ;
 assign nrq2_9 = ( preset_0_0_  &  nsr1_2  &  (~ nlc1_2)  &  (~ ndn2_2) ) ;
 assign wire2372 = ( nsr3_13  &  ndn3_12 ) | ( (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire2373 = ( nen3_36  &  (~ ndn3_36) ) | ( (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire2374 = ( (~ ndn3_29)  &  ndn3_28 ) | ( nen3_39  &  (~ ndn3_39) ) ;
 assign wire2375 = ( ndn3_42  &  (~ ndn3_44) ) | ( (~ ndn3_34)  &  nen3_34 ) ;
 assign wire2377 = ( (~ ndn3_19)  &  nen3_19 ) | ( (~ ndn3_28)  &  nen3_28 ) ;
 assign wire2380 = ( ndn3_39  &  (~ ndn3_40) ) | ( ndn3_25  &  (~ ndn3_26) ) ;
 assign wire2381 = ( (~ ndn3_42)  &  ndn3_40 ) | ( ndn3_29  &  (~ ndn3_32) ) ;
 assign wire2383 = ( (~ ndn3_17)  &  ndn3_16 ) | ( (~ ndn3_27)  &  ndn3_26 ) ;
 assign n_n9583 = ( (~ wire16081)  &  (~ wire16082)  &  wire16097 ) | ( (~ wire16081)  &  (~ wire16082)  &  wire16098 ) | ( wire16081  &  (~ wire16097)  &  (~ wire16098) ) | ( wire16082  &  (~ wire16097)  &  (~ wire16098) ) ;
 assign n_n7997 = ( (~ wire16377)  &  (~ wire16378)  &  wire16394 ) | ( (~ wire16377)  &  (~ wire16378)  &  wire16395 ) | ( wire16377  &  (~ wire16394)  &  (~ wire16395) ) | ( wire16378  &  (~ wire16394)  &  (~ wire16395) ) ;
 assign n_n9639 = ( n_n8930  &  n_n8929 ) | ( (~ n_n8930)  &  wire16027 ) | ( (~ n_n8930)  &  wire16028 ) ;
 assign n_n8493 = ( n_n8631 ) | ( n_n8847 ) | ( n_n8561 ) | ( n_n8342 ) ;
 assign n_n8019 = ( n_n7784  &  n_n7872 ) | ( (~ n_n7784)  &  n_n7872  &  wire5311 ) | ( n_n7784  &  (~ n_n7872)  &  wire5311 ) | ( (~ n_n7784)  &  n_n7872  &  wire5312 ) | ( n_n7784  &  (~ n_n7872)  &  wire5312 ) ;
 assign n_n7573 = ( (~ wire16278)  &  (~ wire16279)  &  wire16295 ) | ( (~ wire16278)  &  (~ wire16279)  &  wire16296 ) | ( wire16278  &  (~ wire16295)  &  (~ wire16296) ) | ( wire16279  &  (~ wire16295)  &  (~ wire16296) ) ;
 assign n_n7869 = ( (~ wire16114)  &  (~ wire16115)  &  wire16130 ) | ( (~ wire16114)  &  (~ wire16115)  &  wire16131 ) | ( wire16114  &  (~ wire16130)  &  (~ wire16131) ) | ( wire16115  &  (~ wire16130)  &  (~ wire16131) ) ;
 assign n_n8028 = ( n_n9124  &  n_n9389 ) | ( (~ n_n9124)  &  n_n9389  &  wire5338 ) | ( n_n9124  &  (~ n_n9389)  &  wire5338 ) | ( (~ n_n9124)  &  n_n9389  &  wire5339 ) | ( n_n9124  &  (~ n_n9389)  &  wire5339 ) ;
 assign n_n8953 = ( (~ wire16179)  &  (~ wire16180)  &  wire16196 ) | ( (~ wire16179)  &  (~ wire16180)  &  wire16197 ) | ( wire16179  &  (~ wire16196)  &  (~ wire16197) ) | ( wire16180  &  (~ wire16196)  &  (~ wire16197) ) ;
 assign n_n9197 = ( wire2372 ) | ( wire16464 ) | ( wire16465 ) | ( wire16466 ) ;
 assign n_n8667 = ( (~ n_n9198)  &  (~ n_n8668) ) | ( (~ n_n8668)  &  (~ n_n9639)  &  n_n9197 ) ;
 assign n_n7566 = ( n_n9332  &  n_n8321 ) | ( (~ n_n9332)  &  n_n8321  &  wire5184 ) | ( n_n9332  &  (~ n_n8321)  &  wire5184 ) | ( (~ n_n9332)  &  n_n8321  &  wire5185 ) | ( n_n9332  &  (~ n_n8321)  &  wire5185 ) ;
 assign n_n8154 = ( (~ wire16311)  &  (~ wire16312)  &  wire16328 ) | ( (~ wire16311)  &  (~ wire16312)  &  wire16329 ) | ( wire16311  &  (~ wire16328)  &  (~ wire16329) ) | ( wire16312  &  (~ wire16328)  &  (~ wire16329) ) ;
 assign n_n7818 = ( wire5495 ) | ( wire5496 ) | ( wire16110 ) | ( wire16115 ) ;
 assign n_n7597 = ( wire5477 ) | ( wire5478 ) | ( wire16126 ) | ( wire16131 ) ;
 assign n_n8314 = ( (~ wire16445)  &  (~ wire16446)  &  wire16461 ) | ( (~ wire16445)  &  (~ wire16446)  &  wire16462 ) | ( wire16445  &  (~ wire16461)  &  (~ wire16462) ) | ( wire16446  &  (~ wire16461)  &  (~ wire16462) ) ;
 assign n_n9040 = ( wire5402 ) | ( wire5403 ) | ( wire16208 ) | ( wire16213 ) ;
 assign n_n9307 = ( wire5420 ) | ( wire5421 ) | ( wire16225 ) | ( wire16230 ) ;
 assign n_n9332 = ( wire5227 ) | ( wire5228 ) | ( wire16340 ) | ( wire16345 ) ;
 assign n_n8321 = ( wire5165 ) | ( wire5166 ) | ( wire16357 ) | ( wire16362 ) ;
 assign n_n7311 = ( (~ wire16573)  &  (~ wire16574)  &  wire16590 ) | ( (~ wire16573)  &  (~ wire16574)  &  wire16591 ) | ( wire16573  &  (~ wire16590)  &  (~ wire16591) ) | ( wire16574  &  (~ wire16590)  &  (~ wire16591) ) ;
 assign n_n7544 = ( n_n8315  &  n_n8316 ) | ( (~ n_n8315)  &  n_n8316  &  wire5069 ) | ( n_n8315  &  (~ n_n8316)  &  wire5069 ) | ( (~ n_n8315)  &  n_n8316  &  wire5070 ) | ( n_n8315  &  (~ n_n8316)  &  wire5070 ) ;
 assign n_n8320 = ( (~ wire16344)  &  (~ wire16345)  &  wire16361 ) | ( (~ wire16344)  &  (~ wire16345)  &  wire16362 ) | ( wire16344  &  (~ wire16361)  &  (~ wire16362) ) | ( wire16345  &  (~ wire16361)  &  (~ wire16362) ) ;
 assign n_n8156 = ( wire5124 ) | ( wire5125 ) | ( wire16307 ) | ( wire16312 ) ;
 assign n_n8155 = ( wire5142 ) | ( wire5143 ) | ( wire16324 ) | ( wire16329 ) ;
 assign n_n9124 = ( wire5457 ) | ( wire5458 ) | ( wire16142 ) | ( wire16147 ) ;
 assign n_n9389 = ( wire5319 ) | ( wire5320 ) | ( wire16159 ) | ( wire16164 ) ;
 assign n_n7784 = ( wire5553 ) | ( wire5554 ) | ( wire16041 ) | ( wire16046 ) ;
 assign n_n7872 = ( wire5292 ) | ( wire5293 ) | ( wire16060 ) | ( wire16065 ) ;
 assign n_n8126 = ( wire4787 ) | ( wire4788 ) | ( wire16569 ) | ( wire16574 ) ;
 assign n_n8125 = ( wire4768 ) | ( wire4769 ) | ( wire16586 ) | ( wire16591 ) ;
 assign n_n9478 = ( (~ wire16146)  &  (~ wire16147)  &  wire16163 ) | ( (~ wire16146)  &  (~ wire16147)  &  wire16164 ) | ( wire16146  &  (~ wire16163)  &  (~ wire16164) ) | ( wire16147  &  (~ wire16163)  &  (~ wire16164) ) ;
 assign n_n8865 = ( (~ wire16607)  &  (~ wire16608)  &  wire16623 ) | ( (~ wire16607)  &  (~ wire16608)  &  wire16624 ) | ( wire16607  &  (~ wire16623)  &  (~ wire16624) ) | ( wire16608  &  (~ wire16623)  &  (~ wire16624) ) ;
 assign n_n8579 = ( wire4864 ) | ( wire4865 ) | ( wire4866 ) | ( wire16549 ) ;
 assign n_n8342 = ( n_n9034 ) | ( n_n9031 ) | ( n_n8993 ) | ( n_n8204 ) ;
 assign n_n8932 = ( (~ n_n8603) ) | ( n_n8923 ) | ( n_n8798 ) | ( n_n8869 ) ;
 assign n_n7274 = ( n_n9247  &  wire16463 ) | ( (~ n_n9247)  &  n_n9639  &  wire16469 ) ;
 assign n_n7218 = ( (~ wire16410)  &  (~ wire16411)  &  wire16427 ) | ( (~ wire16410)  &  (~ wire16411)  &  wire16428 ) | ( wire16410  &  (~ wire16427)  &  (~ wire16428) ) | ( wire16411  &  (~ wire16427)  &  (~ wire16428) ) ;
 assign n_n8315 = ( wire5032 ) | ( wire5033 ) | ( wire16441 ) | ( wire16446 ) ;
 assign n_n7939 = ( (~ wire16045)  &  (~ wire16046)  &  wire16064 ) | ( (~ wire16045)  &  (~ wire16046)  &  wire16065 ) | ( wire16045  &  (~ wire16064)  &  (~ wire16065) ) | ( wire16046  &  (~ wire16064)  &  (~ wire16065) ) ;
 assign n_n8204 = ( n_n8911 ) | ( n_n8933 ) | ( n_n8978 ) | ( n_n8932 ) ;
 assign n_n8316 = ( wire5051 ) | ( wire5052 ) | ( wire16457 ) | ( wire16462 ) ;
 assign n_n9258 = ( wire5270 ) | ( wire5271 ) | ( wire16274 ) | ( wire16279 ) ;
 assign n_n9587 = ( wire5251 ) | ( wire5252 ) | ( wire16291 ) | ( wire16296 ) ;
 assign wire2364 = ( (~ preset)  &  ndn3_34  &  n_n8580 ) | ( (~ preset)  &  (~ nen3_34)  &  n_n8580 ) ;
 assign wire2379 = ( (~ preset)  &  ndn3_46  &  n_n8428 ) | ( (~ preset)  &  (~ ndn3_44)  &  n_n8428 ) ;
 assign wire2382 = ( (~ preset)  &  n_n9333  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire2470 = ( (~ preset)  &  ngfdn_3  &  n_n9145 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n9145 ) ;
 assign wire2471 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46  &  n_n9629 ) ;
 assign wire2472 = ( (~ preset)  &  ndn3_17  &  n_n8811 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8811 ) ;
 assign wire2474 = ( (~ preset)  &  (~ nen3_36)  &  n_n7844 ) | ( (~ preset)  &  ndn3_36  &  n_n7844 ) ;
 assign wire2475 = ( (~ preset)  &  nrq3_36  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_36  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire2480 = ( (~ preset)  &  (~ ndn3_17)  &  n_n9131 ) | ( (~ preset)  &  ndn3_18  &  n_n9131 ) ;
 assign wire2482 = ( (~ preset)  &  ngfdn_3  &  n_n8948 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n8948 ) ;
 assign wire2484 = ( (~ preset)  &  psv26_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2485 = ( (~ preset)  &  ndn3_2  &  n_n9405 ) | ( (~ preset)  &  n_n9405  &  (~ nen3_2) ) ;
 assign wire2488 = ( (~ preset)  &  nsr3_35  &  n_n7928 ) | ( (~ preset)  &  ndn3_35  &  n_n7928 ) ;
 assign wire2490 = ( (~ preset)  &  (~ ndn3_25)  &  n_n7453 ) | ( (~ preset)  &  ndn3_26  &  n_n7453 ) ;
 assign wire2492 = ( (~ preset)  &  (~ ndn3_25)  &  n_n7485 ) | ( (~ preset)  &  ndn3_26  &  n_n7485 ) ;
 assign wire2493 = ( (~ preset)  &  ndn_latch3_26  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_26  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire2494 = ( (~ preset)  &  (~ ndn3_9)  &  n_n9345 ) | ( (~ preset)  &  ndn3_11  &  n_n9345 ) ;
 assign wire2498 = ( (~ preset)  &  ndn3_37  &  n_n7788 ) | ( (~ preset)  &  nsr3_37  &  n_n7788 ) ;
 assign wire2502 = ( (~ preset)  &  nsr3_35  &  n_n8078 ) | ( (~ preset)  &  ndn3_35  &  n_n8078 ) ;
 assign wire2504 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7288 ) | ( (~ preset)  &  ndn3_50  &  n_n7288 ) ;
 assign wire2505 = ( (~ preset)  &  ngfdn_3  &  n_n9282  &  (~ ndn3_50) ) ;
 assign wire2506 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7862 ) | ( (~ preset)  &  ndn3_40  &  n_n7862 ) ;
 assign wire2508 = ( (~ preset)  &  psv18_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2509 = ( (~ preset)  &  ndn3_2  &  n_n6976 ) | ( (~ preset)  &  n_n6976  &  (~ nen3_2) ) ;
 assign wire2512 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7344 ) | ( (~ preset)  &  ndn3_50  &  n_n7344 ) ;
 assign wire2513 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n9570 ) ;
 assign wire2514 = ( (~ preset)  &  nsr3_38  &  n_n9590 ) | ( (~ preset)  &  ndn3_38  &  n_n9590 ) ;
 assign wire2516 = ( (~ preset)  &  ndn3_46  &  n_n7203 ) | ( (~ preset)  &  (~ ndn3_44)  &  n_n7203 ) ;
 assign wire2517 = ( (~ preset)  &  n_n9125  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire2518 = ( (~ preset)  &  psv38_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2519 = ( (~ preset)  &  ndn3_2  &  n_n8139 ) | ( (~ preset)  &  n_n8139  &  (~ nen3_2) ) ;
 assign wire2522 = ( (~ preset)  &  (~ nen3_39)  &  n_n8991 ) | ( (~ preset)  &  ndn3_39  &  n_n8991 ) ;
 assign wire2524 = ( (~ preset)  &  ngfdn_3  &  n_n8895 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n8895 ) ;
 assign wire2525 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7570  &  ndn3_46 ) ;
 assign wire2526 = ( (~ preset)  &  nsr3_38  &  n_n7920 ) | ( (~ preset)  &  ndn3_38  &  n_n7920 ) ;
 assign wire2528 = ( (~ preset)  &  (~ ndn3_42)  &  n_n7156 ) | ( (~ preset)  &  ndn3_44  &  n_n7156 ) ;
 assign wire2529 = ( (~ preset)  &  n_n8609  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire2532 = ( (~ preset)  &  (~ ndn3_39)  &  n_n6974 ) | ( (~ preset)  &  ndn3_40  &  n_n6974 ) ;
 assign wire2534 = ( (~ preset)  &  (~ nen3_22)  &  n_n7500 ) | ( (~ preset)  &  ndn3_22  &  n_n7500 ) ;
 assign wire2535 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9460 ) ;
 assign wire2542 = ( (~ preset)  &  (~ ndn3_17)  &  n_n9048 ) | ( (~ preset)  &  ndn3_18  &  n_n9048 ) ;
 assign wire2543 = ( (~ preset)  &  nrq3_18  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_18  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire2544 = ( (~ preset)  &  psv38_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2545 = ( (~ preset)  &  ndn3_2  &  n_n9262 ) | ( (~ preset)  &  n_n9262  &  (~ nen3_2) ) ;
 assign wire2548 = ( (~ preset)  &  (~ nen3_22)  &  n_n7076 ) | ( (~ preset)  &  ndn3_22  &  n_n7076 ) ;
 assign wire2549 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n8462 ) ;
 assign wire2550 = ( (~ preset)  &  (~ ndn3_42)  &  n_n9632 ) | ( (~ preset)  &  ndn3_44  &  n_n9632 ) ;
 assign wire2554 = ( (~ preset)  &  ndn3_37  &  n_n9505 ) | ( (~ preset)  &  nsr3_37  &  n_n9505 ) ;
 assign wire2558 = ( (~ preset)  &  psv18_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2559 = ( (~ preset)  &  ndn3_2  &  n_n9594 ) | ( (~ preset)  &  n_n9594  &  (~ nen3_2) ) ;
 assign wire2564 = ( (~ preset)  &  psv18_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2565 = ( (~ preset)  &  ndn3_2  &  n_n7886 ) | ( (~ preset)  &  n_n7886  &  (~ nen3_2) ) ;
 assign wire2568 = ( (~ preset)  &  ndn3_4  &  n_n9269 ) | ( (~ preset)  &  (~ ndn3_2)  &  n_n9269 ) ;
 assign wire2569 = ( (~ preset)  &  nrq3_4  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_4  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire2570 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7111 ) | ( (~ preset)  &  ndn3_50  &  n_n7111 ) ;
 assign wire2571 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n9028 ) ;
 assign wire2572 = ( (~ preset)  &  psv2_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2573 = ( (~ preset)  &  ndn3_2  &  n_n9606 ) | ( (~ preset)  &  n_n9606  &  (~ nen3_2) ) ;
 assign wire2576 = ( (~ preset)  &  ndn3_42  &  n_n7927 ) | ( (~ preset)  &  (~ ndn3_40)  &  n_n7927 ) ;
 assign wire2578 = ( (~ preset)  &  (~ ndn3_39)  &  n_n8206 ) | ( (~ preset)  &  ndn3_40  &  n_n8206 ) ;
 assign wire2580 = ( (~ preset)  &  ndn3_27  &  n_n7601 ) | ( (~ preset)  &  n_n7601  &  (~ ndn3_26) ) ;
 assign wire2581 = ( (~ preset)  &  ndn_latch3_27  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_27  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire2584 = ( (~ preset)  &  nsr3_38  &  n_n9392 ) | ( (~ preset)  &  n_n9392  &  ndn3_38 ) ;
 assign wire2586 = ( (~ preset)  &  (~ ndn3_9)  &  n_n9133 ) | ( (~ preset)  &  ndn3_11  &  n_n9133 ) ;
 assign wire2588 = ( (~ preset)  &  nsr3_35  &  n_n7874 ) | ( (~ preset)  &  ndn3_35  &  n_n7874 ) ;
 assign wire2590 = ( n_n8354  &  n_n8353  &  wire16790 ) | ( n_n8354  &  n_n8355  &  wire16790 ) | ( n_n8353  &  n_n8355  &  wire16790 ) ;
 assign wire2591 = ( (~ n_n8419)  &  wire2395  &  (~ n_n8418)  &  n_n8420 ) | ( (~ n_n8419)  &  wire2395  &  n_n8418  &  (~ n_n8420) ) ;
 assign wire2592 = ( n_n8419  &  wire2363  &  (~ n_n8418)  &  (~ n_n8420) ) ;
 assign wire2593 = ( (~ preset)  &  n_n8419  &  (~ n_n7274) ) ;
 assign wire2594 = ( (~ preset)  &  (~ nen3_36)  &  n_n7664 ) | ( (~ preset)  &  ndn3_36  &  n_n7664 ) ;
 assign wire2595 = ( (~ preset)  &  nrq3_36  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_36  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire2596 = ( (~ preset)  &  ndn3_9  &  n_n9051 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n9051 ) ;
 assign wire2597 = ( (~ preset)  &  nrq3_9  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_9  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire2598 = ( (~ preset)  &  ndn3_27  &  n_n9077 ) | ( (~ preset)  &  n_n9077  &  (~ ndn3_26) ) ;
 assign wire2606 = ( (~ preset)  &  psv13_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2607 = ( (~ preset)  &  ndn3_2  &  n_n9604 ) | ( (~ preset)  &  n_n9604  &  (~ nen3_2) ) ;
 assign wire2612 = ( (~ preset)  &  ndn3_29  &  n_n8937 ) | ( (~ preset)  &  (~ ndn3_28)  &  n_n8937 ) ;
 assign wire2613 = ( (~ preset)  &  ndn_latch3_29  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_29  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire2614 = ( (~ preset)  &  psv39_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2615 = ( (~ preset)  &  ndn3_2  &  n_n8416 ) | ( (~ preset)  &  n_n8416  &  (~ nen3_2) ) ;
 assign wire2630 = ( (~ preset)  &  nsr3_20  &  n_n7653 ) | ( (~ preset)  &  n_n7653  &  ndn3_20 ) ;
 assign wire2634 = ( (~ preset)  &  psv33_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2635 = ( (~ preset)  &  ndn3_2  &  n_n9348 ) | ( (~ preset)  &  n_n9348  &  (~ nen3_2) ) ;
 assign wire2638 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7136 ) | ( (~ preset)  &  ndn3_40  &  n_n7136 ) ;
 assign wire2640 = ( (~ preset)  &  psv26_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2641 = ( (~ preset)  &  ndn3_2  &  n_n8051 ) | ( (~ preset)  &  n_n8051  &  (~ nen3_2) ) ;
 assign wire2648 = ( (~ preset)  &  ngfdn_3  &  n_n8850 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n8850 ) ;
 assign wire2649 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n9573  &  ndn3_46 ) ;
 assign wire2655 = ( n_n8806  &  wire4421 ) | ( n_n8806  &  n_n8667  &  wire16682 ) ;
 assign wire2656 = ( n_n8561  &  wire2363  &  n_n8342 ) | ( (~ n_n8561)  &  wire2363  &  (~ n_n8342) ) ;
 assign wire2657 = ( (~ preset)  &  (~ ndn3_17)  &  n_n8058 ) | ( (~ preset)  &  ndn3_18  &  n_n8058 ) ;
 assign wire2659 = ( (~ preset)  &  psv26_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2660 = ( (~ preset)  &  ndn3_2  &  n_n8192 ) | ( (~ preset)  &  n_n8192  &  (~ nen3_2) ) ;
 assign wire2665 = ( (~ preset)  &  nsr3_38  &  n_n7949 ) | ( (~ preset)  &  n_n7949  &  ndn3_38 ) ;
 assign wire2673 = ( (~ preset)  &  ndn3_9  &  n_n7792 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n7792 ) ;
 assign wire2675 = ( (~ preset)  &  psv18_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2676 = ( (~ preset)  &  ndn3_2  &  n_n9232 ) | ( (~ preset)  &  n_n9232  &  (~ nen3_2) ) ;
 assign wire2679 = ( (~ preset)  &  psv13_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2680 = ( (~ preset)  &  ndn3_2  &  n_n7815 ) | ( (~ preset)  &  n_n7815  &  (~ nen3_2) ) ;
 assign wire2683 = ( (~ preset)  &  psv2_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2684 = ( (~ preset)  &  ndn3_2  &  n_n7881 ) | ( (~ preset)  &  n_n7881  &  (~ nen3_2) ) ;
 assign wire2687 = ( (~ preset)  &  psv18_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2688 = ( (~ preset)  &  ndn3_2  &  n_n8033 ) | ( (~ preset)  &  n_n8033  &  (~ nen3_2) ) ;
 assign wire2691 = ( (~ preset)  &  nsr3_14  &  n_n9525 ) | ( (~ preset)  &  n_n9525  &  ndn3_14 ) ;
 assign wire2697 = ( (~ preset)  &  psv2_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2698 = ( (~ preset)  &  ndn3_2  &  n_n8770 ) | ( (~ preset)  &  n_n8770  &  (~ nen3_2) ) ;
 assign wire2701 = ( pinp_6_6_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2702 = ( (~ preset)  &  ndn3_2  &  n_n7644 ) | ( (~ preset)  &  n_n7644  &  (~ nen3_2) ) ;
 assign wire2703 = ( (~ preset)  &  ndn3_19  &  n_n8151 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n8151 ) ;
 assign wire2704 = ( (~ preset)  &  nrq3_19  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_19  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire2705 = ( (~ preset)  &  ndn3_17  &  n_n8226 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8226 ) ;
 assign wire2709 = ( (~ preset)  &  ndn3_23  &  n_n8841 ) | ( (~ preset)  &  nsr3_23  &  n_n8841 ) ;
 assign wire2711 = ( (~ preset)  &  ndn3_19  &  n_n8280 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n8280 ) ;
 assign wire2712 = ( (~ preset)  &  nrq3_19  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_19  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire2713 = ( (~ preset)  &  ndn3_23  &  n_n7846 ) | ( (~ preset)  &  nsr3_23  &  n_n7846 ) ;
 assign wire2715 = ( (~ preset)  &  ndn3_42  &  n_n7678 ) | ( (~ preset)  &  (~ ndn3_40)  &  n_n7678 ) ;
 assign wire2716 = ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40  &  n_n7862 ) ;
 assign wire2717 = ( (~ preset)  &  ndn3_27  &  n_n7666 ) | ( (~ preset)  &  n_n7666  &  (~ ndn3_26) ) ;
 assign wire2718 = ( (~ preset)  &  ndn_latch3_27  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_27  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire2719 = ( (~ preset)  &  (~ nen3_22)  &  n_n9520 ) | ( (~ preset)  &  ndn3_22  &  n_n9520 ) ;
 assign wire2721 = ( (~ preset)  &  psv39_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2722 = ( (~ preset)  &  ndn3_2  &  n_n7956 ) | ( (~ preset)  &  n_n7956  &  (~ nen3_2) ) ;
 assign wire2725 = ( (~ preset)  &  ndn3_30  &  n_n7732 ) | ( (~ preset)  &  nsr3_30  &  n_n7732 ) ;
 assign wire2727 = ( (~ preset)  &  ndn3_28  &  n_n7859 ) | ( (~ preset)  &  (~ nen3_28)  &  n_n7859 ) ;
 assign wire2731 = ( pinp_12_12_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2732 = ( (~ preset)  &  ndn3_2  &  n_n8108 ) | ( (~ preset)  &  n_n8108  &  (~ nen3_2) ) ;
 assign wire2735 = ( (~ preset)  &  (~ nen3_22)  &  n_n9026 ) | ( (~ preset)  &  ndn3_22  &  n_n9026 ) ;
 assign wire2736 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n7236 ) ;
 assign wire2737 = ( (~ preset)  &  psv38_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2738 = ( (~ preset)  &  ndn3_2  &  n_n8088 ) | ( (~ preset)  &  n_n8088  &  (~ nen3_2) ) ;
 assign wire2743 = ( (~ preset)  &  psv38_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2744 = ( (~ preset)  &  ndn3_2  &  n_n9225 ) | ( (~ preset)  &  n_n9225  &  (~ nen3_2) ) ;
 assign wire2747 = ( (~ preset)  &  ndn3_42  &  n_n8102 ) | ( (~ preset)  &  (~ ndn3_40)  &  n_n8102 ) ;
 assign wire2748 = ( (~ preset)  &  (~ ndn3_42)  &  n_n9542  &  ndn3_40 ) ;
 assign wire2749 = ( (~ preset)  &  ndn3_4  &  n_n9347 ) | ( (~ preset)  &  (~ ndn3_2)  &  n_n9347 ) ;
 assign wire2751 = ( (~ preset)  &  ngfdn_3  &  n_n7130 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n7130 ) ;
 assign wire2752 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7527  &  ndn3_46 ) ;
 assign wire2755 = ( (~ preset)  &  ndn3_46  &  n_n7444 ) | ( (~ preset)  &  (~ ndn3_44)  &  n_n7444 ) ;
 assign wire2757 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9542 ) | ( (~ preset)  &  n_n9542  &  ndn3_40 ) ;
 assign wire2758 = ( wire2371  &  (~ n_n8865)  &  wire4672 ) | ( wire2371  &  (~ n_n8865)  &  wire4673 ) | ( wire2371  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire2762 = ( (~ preset)  &  ndn3_42  &  n_n8371 ) | ( (~ preset)  &  n_n8371  &  (~ ndn3_40) ) ;
 assign wire2763 = ( (~ preset)  &  (~ ndn3_42)  &  n_n9452  &  ndn3_40 ) ;
 assign wire2764 = ( (~ preset)  &  (~ nen3_36)  &  n_n9455 ) | ( (~ preset)  &  ndn3_36  &  n_n9455 ) ;
 assign wire2768 = ( (~ preset)  &  (~ nen3_36)  &  n_n9261 ) | ( (~ preset)  &  ndn3_36  &  n_n9261 ) ;
 assign wire2769 = ( (~ preset)  &  nrq3_36  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_36  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire2772 = ( (~ preset)  &  ndn3_42  &  n_n7022 ) | ( (~ preset)  &  n_n7022  &  (~ ndn3_40) ) ;
 assign wire2773 = ( (~ preset)  &  n_n8959  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire2774 = ( (~ preset)  &  ndn3_42  &  n_n8303 ) | ( (~ preset)  &  n_n8303  &  (~ ndn3_40) ) ;
 assign wire2775 = ( (~ preset)  &  n_n8957  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire2776 = ( (~ preset)  &  ndn3_28  &  n_n9593 ) | ( (~ preset)  &  (~ nen3_28)  &  n_n9593 ) ;
 assign wire2777 = ( (~ preset)  &  ndn_latch3_28  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_28  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire2780 = ( (~ preset)  &  (~ ndn3_42)  &  n_n7435 ) | ( (~ preset)  &  ndn3_44  &  n_n7435 ) ;
 assign wire2781 = ( (~ preset)  &  ndn3_42  &  (~ ndn3_44)  &  n_n7927 ) ;
 assign wire2782 = ( (~ preset)  &  ndn3_28  &  n_n9313 ) | ( (~ preset)  &  (~ nen3_28)  &  n_n9313 ) ;
 assign wire2783 = ( (~ preset)  &  ndn_latch3_28  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_28  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire2784 = ( (~ preset)  &  ndn3_23  &  n_n9522 ) | ( (~ preset)  &  nsr3_23  &  n_n9522 ) ;
 assign wire2788 = ( (~ preset)  &  nsr3_35  &  n_n9488 ) | ( (~ preset)  &  ndn3_35  &  n_n9488 ) ;
 assign wire2790 = ( (~ preset)  &  (~ ndn3_42)  &  n_n9237 ) | ( (~ preset)  &  ndn3_44  &  n_n9237 ) ;
 assign wire2792 = ( (~ preset)  &  (~ ndn3_42)  &  n_n9239 ) | ( (~ preset)  &  ndn3_44  &  n_n9239 ) ;
 assign wire2794 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9452 ) | ( (~ preset)  &  n_n9452  &  ndn3_40 ) ;
 assign wire2796 = ( (~ preset)  &  ndn3_13  &  n_n9498 ) | ( (~ preset)  &  nsr3_13  &  n_n9498 ) ;
 assign wire2798 = ( (~ preset)  &  (~ ndn3_42)  &  n_n8439 ) | ( (~ preset)  &  ndn3_44  &  n_n8439 ) ;
 assign wire2799 = ( (~ preset)  &  n_n7757  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire2800 = ( (~ preset)  &  (~ ndn3_42)  &  n_n8146 ) | ( (~ preset)  &  ndn3_44  &  n_n8146 ) ;
 assign wire2801 = ( (~ preset)  &  n_n8024  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire2806 = ( (~ preset)  &  ngfdn_3  &  n_n9376 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n9376 ) ;
 assign wire2807 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8436  &  ndn3_46 ) ;
 assign wire2809 = ( n_n8846  &  wire4421 ) | ( n_n8846  &  n_n8667  &  wire16682 ) ;
 assign wire2810 = ( wire2363  &  n_n9152 ) ;
 assign wire2811 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7843 ) | ( (~ preset)  &  ndn3_50  &  n_n7843 ) ;
 assign wire2812 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n8256 ) ;
 assign wire2813 = ( (~ preset)  &  psv18_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2814 = ( (~ preset)  &  n_n8966  &  ndn3_2 ) | ( (~ preset)  &  n_n8966  &  (~ nen3_2) ) ;
 assign wire2819 = ( (~ preset)  &  ndn3_46  &  n_n7674 ) | ( (~ preset)  &  (~ ndn3_44)  &  n_n7674 ) ;
 assign wire2820 = ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44  &  n_n9237 ) ;
 assign wire2821 = ( (~ preset)  &  ndn3_17  &  n_n8727 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8727 ) ;
 assign wire2823 = ( (~ preset)  &  ndn3_46  &  n_n6910 ) | ( (~ preset)  &  (~ ndn3_44)  &  n_n6910 ) ;
 assign wire2824 = ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44  &  n_n9239 ) ;
 assign wire2825 = ( (~ preset)  &  nsr3_38  &  n_n9081 ) | ( (~ preset)  &  n_n9081  &  ndn3_38 ) ;
 assign wire2827 = ( (~ preset)  &  psv26_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2828 = ( (~ preset)  &  n_n7688  &  ndn3_2 ) | ( (~ preset)  &  n_n7688  &  (~ nen3_2) ) ;
 assign wire2831 = ( (~ preset)  &  ndn3_25  &  n_n9338 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n9338 ) ;
 assign wire2833 = ( (~ preset)  &  nsr3_38  &  n_n9061 ) | ( (~ preset)  &  n_n9061  &  ndn3_38 ) ;
 assign wire2835 = ( (~ preset)  &  (~ nen3_16)  &  n_n7686 ) | ( (~ preset)  &  ndn3_16  &  n_n7686 ) ;
 assign wire2836 = ( (~ preset)  &  nrq3_16  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_16  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire2837 = ( (~ preset)  &  psv33_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2838 = ( (~ preset)  &  n_n8267  &  ndn3_2 ) | ( (~ preset)  &  n_n8267  &  (~ nen3_2) ) ;
 assign wire2841 = ( (~ preset)  &  psv39_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2842 = ( (~ preset)  &  n_n8116  &  ndn3_2 ) | ( (~ preset)  &  n_n8116  &  (~ nen3_2) ) ;
 assign wire2845 = ( (~ preset)  &  (~ ndn3_9)  &  n_n8296 ) | ( (~ preset)  &  ndn3_11  &  n_n8296 ) ;
 assign wire2846 = ( (~ preset)  &  nrq3_11  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_11  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire2847 = ( (~ preset)  &  ndn3_13  &  n_n8344 ) | ( (~ preset)  &  nsr3_13  &  n_n8344 ) ;
 assign wire2851 = ( (~ preset)  &  ndn3_37  &  n_n8326 ) | ( (~ preset)  &  nsr3_37  &  n_n8326 ) ;
 assign wire2855 = ( pinp_0_0_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2856 = ( (~ preset)  &  n_n8011  &  ndn3_2 ) | ( (~ preset)  &  n_n8011  &  (~ nen3_2) ) ;
 assign wire2857 = ( (~ preset)  &  ndn3_17  &  n_n8583 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8583 ) ;
 assign wire2864 = ( n_n9435  &  wire4421 ) | ( n_n9435  &  n_n8667  &  wire16682 ) ;
 assign wire2865 = ( n_n8993  &  wire2363  &  n_n8204 ) | ( (~ n_n8993)  &  wire2363  &  (~ n_n8204) ) ;
 assign wire2869 = ( n_n9288  &  wire4421 ) | ( n_n9288  &  n_n8667  &  wire16682 ) ;
 assign wire2870 = ( wire2363  &  n_n9114 ) ;
 assign wire2871 = ( (~ preset)  &  (~ ndn3_29)  &  n_n8628 ) | ( (~ preset)  &  n_n8628  &  ndn3_32 ) ;
 assign wire2872 = ( (~ preset)  &  ndn_latch3_32  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_32  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire2875 = ( (~ preset)  &  psv18_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2876 = ( (~ preset)  &  n_n8586  &  ndn3_2 ) | ( (~ preset)  &  n_n8586  &  (~ nen3_2) ) ;
 assign wire2879 = ( (~ preset)  &  ndn3_23  &  n_n9340 ) | ( (~ preset)  &  nsr3_23  &  n_n9340 ) ;
 assign wire2885 = ( (~ preset)  &  psv18_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2886 = ( (~ preset)  &  n_n8408  &  ndn3_2 ) | ( (~ preset)  &  n_n8408  &  (~ nen3_2) ) ;
 assign wire2891 = ( (~ preset)  &  psv26_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2892 = ( (~ preset)  &  n_n9603  &  ndn3_2 ) | ( (~ preset)  &  n_n9603  &  (~ nen3_2) ) ;
 assign wire2895 = ( (~ preset)  &  nsr3_35  &  n_n7682 ) | ( (~ preset)  &  ndn3_35  &  n_n7682 ) ;
 assign wire2897 = ( (~ preset)  &  psv26_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2898 = ( (~ preset)  &  n_n9322  &  ndn3_2 ) | ( (~ preset)  &  n_n9322  &  (~ nen3_2) ) ;
 assign wire2903 = ( (~ preset)  &  psv33_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2904 = ( (~ preset)  &  n_n7511  &  ndn3_2 ) | ( (~ preset)  &  n_n7511  &  (~ nen3_2) ) ;
 assign wire2907 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7121 ) | ( (~ preset)  &  n_n7121  &  ndn3_40 ) ;
 assign wire2908 = ( (~ preset)  &  ndn3_39  &  n_n7626  &  (~ ndn3_40) ) ;
 assign wire2909 = ( (~ preset)  &  (~ ndn3_42)  &  n_n8468 ) | ( (~ preset)  &  n_n8468  &  ndn3_44 ) ;
 assign wire2910 = ( wire2369  &  (~ n_n8865)  &  wire4672 ) | ( wire2369  &  (~ n_n8865)  &  wire4673 ) | ( wire2369  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire2915 = ( n_n8823  &  wire4421 ) | ( n_n8823  &  n_n8667  &  wire16682 ) ;
 assign wire2916 = ( n_n9031  &  n_n8993  &  wire2363 ) | ( n_n9031  &  wire2363  &  n_n8204 ) | ( (~ n_n9031)  &  (~ n_n8993)  &  wire2363  &  (~ n_n8204) ) ;
 assign wire2917 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9424 ) | ( (~ preset)  &  n_n9424  &  ndn3_40 ) ;
 assign wire2918 = ( (~ preset)  &  ndn3_39  &  (~ ndn3_40)  &  n_n7346 ) ;
 assign wire2919 = ( (~ preset)  &  ndn3_7  &  n_n9404 ) | ( (~ preset)  &  (~ ndn3_4)  &  n_n9404 ) ;
 assign wire2925 = ( (~ preset)  &  nsr3_13  &  n_n9402 ) | ( (~ preset)  &  ndn3_15  &  n_n9402 ) ;
 assign wire2929 = ( (~ preset)  &  (~ ndn3_39)  &  n_n8361 ) | ( (~ preset)  &  n_n8361  &  ndn3_40 ) ;
 assign wire2930 = ( (~ preset)  &  n_n9611  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire2931 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7366 ) | ( (~ preset)  &  n_n7366  &  ndn3_40 ) ;
 assign wire2932 = ( (~ preset)  &  n_n9613  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire2933 = ( (~ preset)  &  nsr3_14  &  n_n9344 ) | ( (~ preset)  &  n_n9344  &  ndn3_14 ) ;
 assign wire2935 = ( (~ preset)  &  ndn3_46  &  n_n7083 ) | ( (~ preset)  &  n_n7083  &  (~ ndn3_44) ) ;
 assign wire2937 = ( (~ preset)  &  (~ ndn3_42)  &  n_n8188 ) | ( (~ preset)  &  n_n8188  &  ndn3_44 ) ;
 assign wire2938 = ( wire2369  &  (~ n_n7939)  &  wire5311 ) | ( wire2369  &  (~ n_n7939)  &  wire5312 ) | ( wire2369  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire2939 = ( (~ preset)  &  nsr3_14  &  n_n9178 ) | ( (~ preset)  &  n_n9178  &  ndn3_14 ) ;
 assign wire2941 = ( (~ preset)  &  (~ ndn3_39)  &  n_n8644 ) | ( (~ preset)  &  n_n8644  &  ndn3_40 ) ;
 assign wire2942 = ( (~ preset)  &  n_n8543  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire2943 = ( (~ preset)  &  (~ ndn3_42)  &  n_n8670 ) | ( (~ preset)  &  n_n8670  &  ndn3_44 ) ;
 assign wire2945 = ( (~ preset)  &  psv33_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2946 = ( (~ preset)  &  n_n9136  &  ndn3_2 ) | ( (~ preset)  &  n_n9136  &  (~ nen3_2) ) ;
 assign wire2949 = ( (~ preset)  &  ndn3_34  &  n_n9390 ) | ( (~ preset)  &  n_n9390  &  (~ nen3_34) ) ;
 assign wire2951 = ( (~ preset)  &  ndn3_4  &  n_n8789 ) | ( (~ preset)  &  n_n8789  &  (~ ndn3_2) ) ;
 assign wire2953 = ( (~ preset)  &  ndn3_27  &  n_n9046 ) | ( (~ preset)  &  n_n9046  &  (~ ndn3_26) ) ;
 assign wire2954 = ( (~ preset)  &  ndn_latch3_27  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_27  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire2955 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8938 ) | ( (~ preset)  &  n_n8938  &  ndn3_26 ) ;
 assign wire2956 = ( (~ preset)  &  ndn_latch3_26  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_26  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire2957 = ( (~ preset)  &  ndn3_46  &  n_n7402 ) | ( (~ preset)  &  n_n7402  &  (~ ndn3_44) ) ;
 assign wire2958 = ( (~ preset)  &  n_n9635  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire2961 = ( (~ preset)  &  psv26_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2962 = ( (~ preset)  &  n_n9067  &  ndn3_2 ) | ( (~ preset)  &  n_n9067  &  (~ nen3_2) ) ;
 assign wire2965 = ( (~ preset)  &  (~ ndn3_42)  &  n_n7715 ) | ( (~ preset)  &  n_n7715  &  ndn3_44 ) ;
 assign wire2966 = ( (~ preset)  &  n_n9486  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire2967 = ( (~ preset)  &  (~ nen3_22)  &  n_n6980 ) | ( (~ preset)  &  ndn3_22  &  n_n6980 ) ;
 assign wire2968 = ( (~ preset)  &  n_n9273  &  nen3_22  &  (~ ndn3_22) ) ;
 assign wire2969 = ( (~ preset)  &  psv38_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2970 = ( (~ preset)  &  n_n8779  &  ndn3_2 ) | ( (~ preset)  &  n_n8779  &  (~ nen3_2) ) ;
 assign wire2974 = ( n_n9010  &  wire4421 ) | ( n_n9010  &  n_n8667  &  wire16682 ) ;
 assign wire2975 = ( wire2363  &  n_n8606 ) ;
 assign wire2976 = ( (~ preset)  &  ndn3_17  &  n_n8729 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8729 ) ;
 assign wire2977 = ( (~ preset)  &  nrq3_17  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_17  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire2978 = ( (~ preset)  &  ndn3_46  &  n_n8916 ) | ( (~ preset)  &  n_n8916  &  (~ ndn3_44) ) ;
 assign wire2979 = ( (~ preset)  &  (~ ndn3_46)  &  n_n8670  &  ndn3_44 ) ;
 assign wire2980 = ( (~ preset)  &  psv2_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2981 = ( (~ preset)  &  n_n7827  &  ndn3_2 ) | ( (~ preset)  &  n_n7827  &  (~ nen3_2) ) ;
 assign wire2984 = ( (~ preset)  &  psv13_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2985 = ( (~ preset)  &  n_n9119  &  ndn3_2 ) | ( (~ preset)  &  n_n9119  &  (~ nen3_2) ) ;
 assign wire2988 = ( (~ preset)  &  psv2_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2989 = ( (~ preset)  &  n_n7744  &  ndn3_2 ) | ( (~ preset)  &  n_n7744  &  (~ nen3_2) ) ;
 assign wire2992 = ( (~ preset)  &  nsr3_14  &  n_n8909 ) | ( (~ preset)  &  n_n8909  &  ndn3_14 ) ;
 assign wire2994 = ( (~ preset)  &  psv13_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire2995 = ( (~ preset)  &  n_n8619  &  ndn3_2 ) | ( (~ preset)  &  n_n8619  &  (~ nen3_2) ) ;
 assign wire2998 = ( (~ preset)  &  nsr3_14  &  n_n8535 ) | ( (~ preset)  &  n_n8535  &  ndn3_14 ) ;
 assign wire3000 = ( (~ preset)  &  (~ ndn3_19)  &  n_n9255 ) | ( (~ preset)  &  ndn3_21  &  n_n9255 ) ;
 assign wire3001 = ( (~ preset)  &  nrq3_21  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_21  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3002 = ( (~ preset)  &  nsr3_14  &  n_n7969 ) | ( (~ preset)  &  n_n7969  &  ndn3_14 ) ;
 assign wire3004 = ( (~ preset)  &  (~ nen3_22)  &  n_n9493 ) | ( (~ preset)  &  ndn3_22  &  n_n9493 ) ;
 assign wire3006 = ( (~ preset)  &  n_n8657  &  nsr3_20 ) | ( (~ preset)  &  n_n8657  &  ndn3_20 ) ;
 assign wire3010 = ( (~ preset)  &  ndn3_37  &  n_n8636 ) | ( (~ preset)  &  n_n8636  &  nsr3_37 ) ;
 assign wire3014 = ( (~ preset)  &  ndn3_37  &  n_n8477 ) | ( (~ preset)  &  n_n8477  &  nsr3_37 ) ;
 assign wire3018 = ( (~ preset)  &  psv2_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3019 = ( (~ preset)  &  n_n7890  &  ndn3_2 ) | ( (~ preset)  &  n_n7890  &  (~ nen3_2) ) ;
 assign wire3025 = ( n_n9216  &  wire4421 ) | ( n_n9216  &  n_n8667  &  wire16682 ) ;
 assign wire3026 = ( (~ n_n8603)  &  n_n8798  &  wire2363 ) | ( n_n8603  &  (~ n_n8798)  &  wire2363 ) ;
 assign wire3027 = ( (~ preset)  &  psv38_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3028 = ( (~ preset)  &  n_n7665  &  ndn3_2 ) | ( (~ preset)  &  n_n7665  &  (~ nen3_2) ) ;
 assign wire3032 = ( wire2363  &  n_n7274  &  wire16775 ) ;
 assign wire3034 = ( (~ preset)  &  n_n9353  &  (~ n_n7274) ) ;
 assign wire3037 = ( (~ preset)  &  ndn3_19  &  n_n9139 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n9139 ) ;
 assign wire3038 = ( (~ preset)  &  nrq3_19  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_19  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3041 = ( (~ preset)  &  ndn3_28  &  n_n8839 ) | ( (~ preset)  &  (~ nen3_28)  &  n_n8839 ) ;
 assign wire3045 = ( (~ preset)  &  (~ nen3_22)  &  n_n8185 ) | ( (~ preset)  &  ndn3_22  &  n_n8185 ) ;
 assign wire3046 = ( (~ preset)  &  nen3_22  &  n_n9304  &  (~ ndn3_22) ) ;
 assign wire3049 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9155 ) | ( (~ preset)  &  n_n9155  &  ndn3_40 ) ;
 assign wire3051 = ( (~ preset)  &  ngfdn_3  &  n_n9508 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n9508 ) ;
 assign wire3052 = ( n_n7098  &  (~ n_n8314)  &  wire5069 ) | ( n_n7098  &  (~ n_n8314)  &  wire5070 ) | ( n_n7098  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire3053 = ( (~ preset)  &  (~ ndn3_29)  &  n_n9126 ) | ( (~ preset)  &  n_n9126  &  ndn3_32 ) ;
 assign wire3055 = ( (~ preset)  &  ndn3_46  &  n_n9629 ) | ( (~ preset)  &  n_n9629  &  (~ ndn3_44) ) ;
 assign wire3056 = ( wire2370  &  (~ n_n8865)  &  wire4672 ) | ( wire2370  &  (~ n_n8865)  &  wire4673 ) | ( wire2370  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire3059 = ( (~ preset)  &  (~ nen3_16)  &  n_n9317 ) | ( (~ preset)  &  ndn3_16  &  n_n9317 ) ;
 assign wire3060 = ( (~ preset)  &  nrq3_16  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_16  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3061 = ( (~ preset)  &  nsr3_13  &  n_n9600 ) | ( (~ preset)  &  ndn3_15  &  n_n9600 ) ;
 assign wire3062 = ( (~ preset)  &  nrq3_15  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_15  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3065 = ( n_n9537  &  n_n8373  &  wire16768 ) | ( n_n9537  &  n_n8936  &  wire16768 ) | ( n_n8373  &  n_n8936  &  wire16768 ) ;
 assign wire3066 = ( (~ n_n8821)  &  wire2395  &  (~ n_n8820)  &  n_n8822 ) | ( (~ n_n8821)  &  wire2395  &  n_n8820  &  (~ n_n8822) ) ;
 assign wire3067 = ( n_n8821  &  wire2363  &  (~ n_n8820)  &  (~ n_n8822) ) ;
 assign wire3068 = ( (~ preset)  &  n_n8821  &  (~ n_n7274) ) ;
 assign wire3073 = ( (~ preset)  &  n_n7074  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7074  &  ndn3_44 ) ;
 assign wire3074 = ( (~ preset)  &  n_n9355  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire3075 = ( (~ preset)  &  n_n8249  &  ndn3_42 ) | ( (~ preset)  &  n_n8249  &  (~ ndn3_40) ) ;
 assign wire3081 = ( (~ preset)  &  psv26_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3082 = ( (~ preset)  &  n_n8617  &  ndn3_2 ) | ( (~ preset)  &  n_n8617  &  (~ nen3_2) ) ;
 assign wire3085 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7069 ) | ( (~ preset)  &  ndn3_50  &  n_n7069 ) ;
 assign wire3086 = ( (~ preset)  &  ngfdn_3  &  n_n7324  &  (~ ndn3_50) ) ;
 assign wire3087 = ( (~ preset)  &  psv33_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3088 = ( (~ preset)  &  n_n9053  &  ndn3_2 ) | ( (~ preset)  &  n_n9053  &  (~ nen3_2) ) ;
 assign wire3091 = ( (~ preset)  &  ndn3_27  &  n_n9129 ) | ( (~ preset)  &  n_n9129  &  (~ ndn3_26) ) ;
 assign wire3095 = ( (~ preset)  &  ndn3_13  &  n_n9320 ) | ( (~ preset)  &  nsr3_13  &  n_n9320 ) ;
 assign wire3101 = ( (~ preset)  &  psv13_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3102 = ( (~ preset)  &  n_n8502  &  ndn3_2 ) | ( (~ preset)  &  n_n8502  &  (~ nen3_2) ) ;
 assign wire3107 = ( (~ preset)  &  psv18_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3108 = ( (~ preset)  &  n_n9230  &  ndn3_2 ) | ( (~ preset)  &  n_n9230  &  (~ nen3_2) ) ;
 assign wire3113 = ( (~ preset)  &  psv38_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3114 = ( (~ preset)  &  n_n7600  &  ndn3_2 ) | ( (~ preset)  &  n_n7600  &  (~ nen3_2) ) ;
 assign wire3117 = ( (~ preset)  &  nsr3_14  &  n_n8221 ) | ( (~ preset)  &  n_n8221  &  ndn3_14 ) ;
 assign wire3121 = ( (~ preset)  &  ndn3_25  &  n_n9595 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n9595 ) ;
 assign wire3122 = ( (~ preset)  &  ndn_latch3_25  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_25  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3123 = ( (~ preset)  &  (~ ndn3_9)  &  n_n7642 ) | ( (~ preset)  &  ndn3_11  &  n_n7642 ) ;
 assign wire3125 = ( pinp_8_8_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3126 = ( (~ preset)  &  n_n7697  &  ndn3_2 ) | ( (~ preset)  &  n_n7697  &  (~ nen3_2) ) ;
 assign wire3127 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7108 ) | ( (~ preset)  &  n_n7108  &  ndn3_40 ) ;
 assign wire3128 = ( (~ preset)  &  n_n8794  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire3129 = ( (~ preset)  &  (~ nen3_16)  &  n_n7810 ) | ( (~ preset)  &  ndn3_16  &  n_n7810 ) ;
 assign wire3131 = ( (~ preset)  &  ngfdn_3  &  n_n7781 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n7781 ) ;
 assign wire3132 = ( n_n7098  &  (~ n_n8320)  &  wire5184 ) | ( n_n7098  &  (~ n_n8320)  &  wire5185 ) | ( n_n7098  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire3135 = ( (~ preset)  &  ngfdn_3  &  n_n7606 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n7606 ) ;
 assign wire3139 = ( (~ preset)  &  (~ ndn3_19)  &  n_n9460 ) | ( (~ preset)  &  ndn3_21  &  n_n9460 ) ;
 assign wire3140 = ( (~ preset)  &  nrq3_21  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_21  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3143 = ( (~ preset)  &  ndn3_25  &  n_n8473 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n8473 ) ;
 assign wire3155 = ( (~ preset)  &  ndn3_29  &  n_n8224 ) | ( (~ preset)  &  (~ ndn3_28)  &  n_n8224 ) ;
 assign wire3157 = ( (~ preset)  &  psv39_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3158 = ( (~ preset)  &  n_n7837  &  ndn3_2 ) | ( (~ preset)  &  n_n7837  &  (~ nen3_2) ) ;
 assign wire3165 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8581 ) | ( (~ preset)  &  n_n8581  &  ndn3_26 ) ;
 assign wire3167 = ( (~ preset)  &  (~ ndn3_19)  &  n_n8213 ) | ( (~ preset)  &  ndn3_21  &  n_n8213 ) ;
 assign wire3168 = ( (~ preset)  &  nrq3_21  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_21  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3171 = ( (~ preset)  &  ndn3_30  &  n_n9092 ) | ( (~ preset)  &  nsr3_30  &  n_n9092 ) ;
 assign wire3177 = ( (~ preset)  &  (~ nen3_22)  &  n_n8781 ) | ( (~ preset)  &  ndn3_22  &  n_n8781 ) ;
 assign wire3178 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9255 ) ;
 assign wire3179 = ( (~ preset)  &  nsr3_35  &  n_n7990 ) | ( (~ preset)  &  ndn3_35  &  n_n7990 ) ;
 assign wire3183 = ( (~ preset)  &  n_n8470  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n8470  &  ndn3_44 ) ;
 assign wire3185 = ( (~ preset)  &  ndn3_30  &  n_n9394 ) | ( (~ preset)  &  nsr3_30  &  n_n9394 ) ;
 assign wire3187 = ( (~ preset)  &  n_n9355  &  ndn3_42 ) | ( (~ preset)  &  n_n9355  &  (~ ndn3_40) ) ;
 assign wire3188 = ( wire2368  &  (~ n_n8865)  &  wire4672 ) | ( wire2368  &  (~ n_n8865)  &  wire4673 ) | ( wire2368  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire3189 = ( (~ preset)  &  (~ nen3_22)  &  n_n7739 ) | ( (~ preset)  &  ndn3_22  &  n_n7739 ) ;
 assign wire3191 = ( n_n8930  &  wire16759 ) | ( (~ n_n9639)  &  wire16759 ) | ( (~ wire16469)  &  wire16759 ) ;
 assign wire3192 = ( (~ n_n8930)  &  n_n9639  &  wire16469  &  wire16760 ) ;
 assign wire3193 = ( (~ preset)  &  (~ nen3_22)  &  n_n7728 ) | ( (~ preset)  &  ndn3_22  &  n_n7728 ) ;
 assign wire3195 = ( (~ preset)  &  n_n8045  &  ndn3_42 ) | ( (~ preset)  &  n_n8045  &  (~ ndn3_40) ) ;
 assign wire3196 = ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40  &  n_n7136 ) ;
 assign wire3197 = ( (~ preset)  &  (~ nen3_36)  &  n_n9128 ) | ( (~ preset)  &  n_n9128  &  ndn3_36 ) ;
 assign wire3199 = ( (~ preset)  &  ndn3_28  &  n_n9159 ) | ( (~ preset)  &  n_n9159  &  (~ nen3_28) ) ;
 assign wire3205 = ( (~ preset)  &  nsr3_35  &  n_n9591 ) | ( (~ preset)  &  ndn3_35  &  n_n9591 ) ;
 assign wire3207 = ( (~ preset)  &  nsr3_35  &  n_n9393 ) | ( (~ preset)  &  ndn3_35  &  n_n9393 ) ;
 assign wire3211 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8263 ) | ( (~ preset)  &  ndn3_50  &  n_n8263 ) ;
 assign wire3212 = ( (~ preset)  &  ngfdn_3  &  n_n8081  &  (~ ndn3_50) ) ;
 assign wire3213 = ( (~ preset)  &  (~ ndn3_9)  &  n_n7848 ) | ( (~ preset)  &  ndn3_11  &  n_n7848 ) ;
 assign wire3214 = ( (~ preset)  &  nrq3_11  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_11  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3215 = ( (~ preset)  &  (~ nen3_39)  &  n_n7626 ) | ( (~ preset)  &  ndn3_39  &  n_n7626 ) ;
 assign wire3216 = ( (~ preset)  &  nrq3_39  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_39  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3217 = ( (~ preset)  &  ndn3_46  &  n_n9421 ) | ( (~ preset)  &  n_n9421  &  (~ ndn3_44) ) ;
 assign wire3218 = ( (~ preset)  &  n_n7691  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire3219 = ( (~ preset)  &  ndn3_9  &  n_n7849 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n7849 ) ;
 assign wire3220 = ( (~ preset)  &  nrq3_9  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_9  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3221 = ( (~ preset)  &  nsr3_38  &  n_n7873 ) | ( (~ preset)  &  n_n7873  &  ndn3_38 ) ;
 assign wire3223 = ( (~ preset)  &  psv33_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3224 = ( (~ preset)  &  n_n7914  &  ndn3_2 ) | ( (~ preset)  &  n_n7914  &  (~ nen3_2) ) ;
 assign wire3227 = ( (~ preset)  &  ndn3_9  &  n_n7668 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n7668 ) ;
 assign wire3228 = ( (~ preset)  &  nrq3_9  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_9  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3231 = ( (~ preset)  &  ndn3_30  &  n_n7925 ) | ( (~ preset)  &  nsr3_30  &  n_n7925 ) ;
 assign wire3233 = ( (~ preset)  &  ngfdn_3  &  n_n8256 ) | ( (~ preset)  &  (~ ndn3_46)  &  n_n8256 ) ;
 assign wire3235 = ( (~ preset)  &  ndn3_23  &  n_n7711 ) | ( (~ preset)  &  nsr3_23  &  n_n7711 ) ;
 assign wire3239 = ( (~ preset)  &  ndn3_4  &  n_n7971 ) | ( (~ preset)  &  n_n7971  &  (~ ndn3_2) ) ;
 assign wire3243 = ( (~ preset)  &  n_n8064  &  nsr3_20 ) | ( (~ preset)  &  n_n8064  &  ndn3_20 ) ;
 assign wire3245 = ( (~ preset)  &  (~ nen3_22)  &  n_n7932 ) | ( (~ preset)  &  ndn3_22  &  n_n7932 ) ;
 assign wire3247 = ( (~ preset)  &  nsr3_13  &  n_n8233 ) | ( (~ preset)  &  ndn3_15  &  n_n8233 ) ;
 assign wire3248 = ( (~ preset)  &  nrq3_15  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_15  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3251 = ( (~ preset)  &  ndn3_25  &  n_n8003 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n8003 ) ;
 assign wire3253 = ( n_n9416  &  n_n8783  &  wire16754 ) | ( n_n9416  &  n_n8784  &  wire16754 ) | ( n_n8783  &  n_n8784  &  wire16754 ) ;
 assign wire3254 = ( (~ n_n9537)  &  wire2395  &  (~ n_n8373)  &  n_n8936 ) | ( (~ n_n9537)  &  wire2395  &  n_n8373  &  (~ n_n8936) ) ;
 assign wire3255 = ( n_n9537  &  wire2363  &  (~ n_n8373)  &  (~ n_n8936) ) ;
 assign wire3256 = ( (~ preset)  &  n_n9537  &  (~ n_n7274) ) ;
 assign wire3257 = ( n_n9638  &  n_n8979  &  wire16748 ) | ( n_n9638  &  n_n7432  &  wire16748 ) | ( n_n8979  &  n_n7432  &  wire16748 ) ;
 assign wire3258 = ( (~ n_n9448)  &  wire2395  &  (~ n_n8323)  &  n_n8324 ) | ( (~ n_n9448)  &  wire2395  &  n_n8323  &  (~ n_n8324) ) ;
 assign wire3259 = ( n_n9448  &  wire2363  &  (~ n_n8323)  &  (~ n_n8324) ) ;
 assign wire3260 = ( (~ preset)  &  n_n9448  &  (~ n_n7274) ) ;
 assign wire3261 = ( (~ preset)  &  ndn3_46  &  n_n9221 ) | ( (~ preset)  &  n_n9221  &  (~ ndn3_44) ) ;
 assign wire3263 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9104 ) | ( (~ preset)  &  n_n9104  &  ndn3_40 ) ;
 assign wire3267 = ( (~ preset)  &  (~ ndn3_29)  &  n_n8277 ) | ( (~ preset)  &  n_n8277  &  ndn3_32 ) ;
 assign wire3268 = ( (~ preset)  &  ndn_latch3_32  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_32  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3269 = ( (~ preset)  &  ndn3_19  &  n_n8743 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n8743 ) ;
 assign wire3270 = ( (~ preset)  &  nrq3_19  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_19  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3271 = ( (~ preset)  &  psv33_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3272 = ( (~ preset)  &  n_n7554  &  ndn3_2 ) | ( (~ preset)  &  n_n7554  &  (~ nen3_2) ) ;
 assign wire3277 = ( n_n8419  &  n_n8418  &  wire16742 ) | ( n_n8419  &  n_n8420  &  wire16742 ) | ( n_n8418  &  n_n8420  &  wire16742 ) ;
 assign wire3278 = ( (~ n_n8449)  &  wire2395  &  (~ n_n8450)  &  n_n8448 ) | ( (~ n_n8449)  &  wire2395  &  n_n8450  &  (~ n_n8448) ) ;
 assign wire3279 = ( n_n8449  &  wire2363  &  (~ n_n8450)  &  (~ n_n8448) ) ;
 assign wire3280 = ( (~ preset)  &  n_n8449  &  (~ n_n7274) ) ;
 assign wire3281 = ( (~ preset)  &  (~ nen3_22)  &  n_n8384 ) | ( (~ preset)  &  ndn3_22  &  n_n8384 ) ;
 assign wire3282 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n8464 ) ;
 assign wire3283 = ( (~ preset)  &  psv38_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3284 = ( (~ preset)  &  n_n9212  &  ndn3_2 ) | ( (~ preset)  &  n_n9212  &  (~ nen3_2) ) ;
 assign wire3289 = ( (~ preset)  &  (~ ndn3_9)  &  n_n9050 ) | ( (~ preset)  &  ndn3_11  &  n_n9050 ) ;
 assign wire3290 = ( (~ preset)  &  nrq3_11  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_11  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3291 = ( (~ preset)  &  ngfdn_3  &  n_n9570 ) | ( (~ preset)  &  n_n9570  &  (~ ndn3_46) ) ;
 assign wire3292 = ( n_n7098  &  (~ n_n7939)  &  wire5311 ) | ( n_n7098  &  (~ n_n7939)  &  wire5312 ) | ( n_n7098  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire3293 = ( (~ preset)  &  ngfdn_3  &  n_n9028 ) | ( (~ preset)  &  n_n9028  &  (~ ndn3_46) ) ;
 assign wire3295 = ( (~ preset)  &  ngfdn_3  &  n_n9626 ) | ( (~ preset)  &  n_n9626  &  (~ ndn3_46) ) ;
 assign wire3299 = ( (~ preset)  &  psv39_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3300 = ( (~ preset)  &  n_n9605  &  ndn3_2 ) | ( (~ preset)  &  n_n9605  &  (~ nen3_2) ) ;
 assign wire3303 = ( (~ preset)  &  nsr3_35  &  n_n6968 ) | ( (~ preset)  &  n_n6968  &  ndn3_35 ) ;
 assign wire3307 = ( (~ preset)  &  (~ ndn3_39)  &  n_n7390 ) | ( (~ preset)  &  n_n7390  &  ndn3_40 ) ;
 assign wire3308 = ( (~ preset)  &  ndn3_39  &  (~ ndn3_40)  &  n_n7334 ) ;
 assign wire3309 = ( (~ preset)  &  psv33_7_7_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3310 = ( (~ preset)  &  n_n9270  &  ndn3_2 ) | ( (~ preset)  &  n_n9270  &  (~ nen3_2) ) ;
 assign wire3313 = ( (~ preset)  &  n_n7284  &  ndn3_46 ) | ( (~ preset)  &  n_n7284  &  (~ ndn3_44) ) ;
 assign wire3314 = ( (~ preset)  &  n_n7898  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire3315 = ( (~ preset)  &  ndn3_13  &  n_n9403 ) | ( (~ preset)  &  nsr3_13  &  n_n9403 ) ;
 assign wire3317 = ( (~ preset)  &  ndn3_34  &  n_n9308 ) | ( (~ preset)  &  n_n9308  &  (~ nen3_34) ) ;
 assign wire3318 = ( (~ preset)  &  nrq3_34  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_34  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3319 = ( (~ preset)  &  (~ ndn3_11)  &  n_n8584 ) | ( (~ preset)  &  ndn3_12  &  n_n8584 ) ;
 assign wire3321 = ( (~ preset)  &  psv26_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3322 = ( (~ preset)  &  n_n7946  &  ndn3_2 ) | ( (~ preset)  &  n_n7946  &  (~ nen3_2) ) ;
 assign wire3325 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7420 ) | ( (~ preset)  &  ndn3_50  &  n_n7420 ) ;
 assign wire3326 = ( (~ preset)  &  n_n7558  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign wire3327 = ( (~ preset)  &  psv18_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3328 = ( (~ preset)  &  n_n7737  &  ndn3_2 ) | ( (~ preset)  &  n_n7737  &  (~ nen3_2) ) ;
 assign wire3331 = ( (~ preset)  &  psv39_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3332 = ( (~ preset)  &  n_n8506  &  ndn3_2 ) | ( (~ preset)  &  n_n8506  &  (~ nen3_2) ) ;
 assign wire3335 = ( (~ preset)  &  (~ ndn3_29)  &  n_n7598 ) | ( (~ preset)  &  n_n7598  &  ndn3_32 ) ;
 assign wire3336 = ( (~ preset)  &  ndn_latch3_32  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_32  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3337 = ( (~ preset)  &  n_n8328  &  ndn3_37 ) | ( (~ preset)  &  n_n8328  &  nsr3_37 ) ;
 assign wire3342 = ( n_n9553  &  wire4421 ) | ( n_n9553  &  n_n8667  &  wire16682 ) ;
 assign wire3343 = ( wire2363  &  n_n7637 ) ;
 assign wire3346 = ( (~ preset)  &  (~ ndn3_25)  &  n_n9205 ) | ( (~ preset)  &  n_n9205  &  ndn3_26 ) ;
 assign wire3348 = ( (~ preset)  &  (~ nen3_22)  &  n_n8004 ) | ( (~ preset)  &  ndn3_22  &  n_n8004 ) ;
 assign wire3349 = ( wire2367  &  (~ n_n8865)  &  wire4672 ) | ( wire2367  &  (~ n_n8865)  &  wire4673 ) | ( wire2367  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire3350 = ( (~ preset)  &  n_n8061  &  ndn3_42 ) | ( (~ preset)  &  n_n8061  &  (~ ndn3_40) ) ;
 assign wire3351 = ( (~ preset)  &  n_n9104  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire3352 = ( (~ preset)  &  psv39_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3353 = ( (~ preset)  &  n_n9121  &  ndn3_2 ) | ( (~ preset)  &  n_n9121  &  (~ nen3_2) ) ;
 assign wire3356 = ( (~ preset)  &  n_n8436  &  ndn3_46 ) | ( (~ preset)  &  n_n8436  &  (~ ndn3_44) ) ;
 assign wire3357 = ( wire2370  &  (~ n_n8320)  &  wire5184 ) | ( wire2370  &  (~ n_n8320)  &  wire5185 ) | ( wire2370  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire3360 = ( (~ preset)  &  n_n9309  &  ndn3_42 ) | ( (~ preset)  &  n_n9309  &  (~ ndn3_40) ) ;
 assign wire3362 = ( (~ preset)  &  n_n9259  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9259  &  ndn3_44 ) ;
 assign wire3364 = ( (~ preset)  &  (~ nsr1_2)  &  n_n7476 ) | ( (~ preset)  &  n_n7476  &  nlc1_2 ) ;
 assign wire3365 = ( (~ preset_0_0_)  &  (~ preset)  &  nsr1_2  &  (~ nlc1_2) ) ;
 assign wire3366 = ( (~ preset)  &  psv26_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3367 = ( (~ preset)  &  n_n7424  &  ndn3_2 ) | ( (~ preset)  &  n_n7424  &  (~ nen3_2) ) ;
 assign wire3370 = ( (~ preset)  &  psv33_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3371 = ( (~ preset)  &  n_n7604  &  ndn3_2 ) | ( (~ preset)  &  n_n7604  &  (~ nen3_2) ) ;
 assign wire3374 = ( (~ preset)  &  ndn3_27  &  n_n7649 ) | ( (~ preset)  &  n_n7649  &  (~ ndn3_26) ) ;
 assign wire3376 = ( (~ preset)  &  ngfdn_3  &  n_n7976 ) | ( (~ preset)  &  n_n7976  &  (~ ndn3_46) ) ;
 assign wire3377 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8765  &  ndn3_46 ) ;
 assign wire3378 = ( (~ preset)  &  ndn3_34  &  n_n8898 ) | ( (~ preset)  &  n_n8898  &  (~ nen3_34) ) ;
 assign wire3379 = ( (~ preset)  &  nrq3_34  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_34  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3380 = ( (~ preset)  &  ndn3_34  &  n_n8222 ) | ( (~ preset)  &  n_n8222  &  (~ nen3_34) ) ;
 assign wire3382 = ( (~ preset)  &  n_n7964  &  ndn3_46 ) | ( (~ preset)  &  n_n7964  &  (~ ndn3_44) ) ;
 assign wire3383 = ( (~ preset)  &  n_n9041  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire3384 = ( (~ preset)  &  n_n7706  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7706  &  ndn3_44 ) ;
 assign wire3386 = ( (~ preset)  &  (~ ndn3_11)  &  n_n9318 ) | ( (~ preset)  &  ndn3_12  &  n_n9318 ) ;
 assign wire3387 = ( (~ preset)  &  ndn_latch3_12  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_12  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3388 = ( pinp_7_7_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3389 = ( (~ preset)  &  n_n9271  &  ndn3_2 ) | ( (~ preset)  &  n_n9271  &  (~ nen3_2) ) ;
 assign wire3390 = ( (~ preset)  &  (~ ndn3_29)  &  n_n9042 ) | ( (~ preset)  &  n_n9042  &  ndn3_32 ) ;
 assign wire3391 = ( (~ preset)  &  ndn_latch3_32  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_32  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3401 = ( n_n7787  &  wire4421 ) | ( n_n7787  &  n_n8667  &  wire16682 ) ;
 assign wire3402 = ( wire2363  &  n_n8976 ) ;
 assign wire3406 = ( n_n9072  &  wire4421 ) | ( n_n9072  &  n_n8667  &  wire16682 ) ;
 assign wire3407 = ( (~ n_n8603)  &  n_n8923  &  wire2363 ) | ( n_n8923  &  n_n8798  &  wire2363 ) | ( n_n8603  &  (~ n_n8923)  &  (~ n_n8798)  &  wire2363 ) ;
 assign wire3410 = ( n_n9248  &  (~ n_n9247)  &  wire16734 ) | ( n_n9248  &  (~ n_n9246)  &  wire16734 ) ;
 assign wire3411 = ( (~ preset)  &  n_n9248  &  n_n9247  &  (~ n_n9246) ) ;
 assign wire3414 = ( (~ preset)  &  (~ ndn3_19)  &  n_n9252 ) | ( (~ preset)  &  ndn3_21  &  n_n9252 ) ;
 assign wire3415 = ( (~ preset)  &  nrq3_21  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_21  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3416 = ( (~ preset)  &  (~ ndn3_39)  &  n_n9576 ) | ( (~ preset)  &  n_n9576  &  ndn3_40 ) ;
 assign wire3422 = ( (~ preset)  &  n_n6920  &  ndn3_46 ) | ( (~ preset)  &  n_n6920  &  (~ ndn3_44) ) ;
 assign wire3423 = ( (~ preset)  &  (~ ndn3_46)  &  n_n8470  &  ndn3_44 ) ;
 assign wire3424 = ( (~ preset)  &  psv38_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3425 = ( (~ preset)  &  n_n7692  &  ndn3_2 ) | ( (~ preset)  &  n_n7692  &  (~ nen3_2) ) ;
 assign wire3428 = ( (~ preset)  &  psv2_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3429 = ( (~ preset)  &  n_n9023  &  ndn3_2 ) | ( (~ preset)  &  n_n9023  &  (~ nen3_2) ) ;
 assign wire3432 = ( (~ preset)  &  nsr3_38  &  n_n9059 ) | ( (~ preset)  &  n_n9059  &  ndn3_38 ) ;
 assign wire3446 = ( (~ preset)  &  (~ nen3_22)  &  n_n7809 ) | ( (~ preset)  &  ndn3_22  &  n_n7809 ) ;
 assign wire3447 = ( wire2367  &  (~ n_n8314)  &  wire5069 ) | ( wire2367  &  (~ n_n8314)  &  wire5070 ) | ( wire2367  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire3448 = ( (~ preset)  &  ndn3_28  &  n_n8889 ) | ( (~ preset)  &  n_n8889  &  (~ nen3_28) ) ;
 assign wire3449 = ( (~ preset)  &  ndn_latch3_28  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_28  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3450 = ( (~ preset)  &  (~ nen3_36)  &  n_n8253 ) | ( (~ preset)  &  n_n8253  &  ndn3_36 ) ;
 assign wire3451 = ( (~ preset)  &  nrq3_36  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_36  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3452 = ( (~ preset)  &  ndn3_27  &  n_n7845 ) | ( (~ preset)  &  n_n7845  &  (~ ndn3_26) ) ;
 assign wire3453 = ( (~ preset)  &  ndn_latch3_27  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_27  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3456 = ( (~ preset)  &  n_n8989  &  ndn3_42 ) | ( (~ preset)  &  n_n8989  &  (~ ndn3_40) ) ;
 assign wire3457 = ( wire2368  &  (~ n_n8320)  &  wire5184 ) | ( wire2368  &  (~ n_n8320)  &  wire5185 ) | ( wire2368  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire3458 = ( (~ preset)  &  (~ ndn3_29)  &  n_n8223 ) | ( (~ preset)  &  n_n8223  &  ndn3_32 ) ;
 assign wire3462 = ( (~ preset)  &  n_n9171  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9171  &  ndn3_44 ) ;
 assign wire3466 = ( (~ preset)  &  ndn3_13  &  n_n7879 ) | ( (~ preset)  &  nsr3_13  &  n_n7879 ) ;
 assign wire3468 = ( (~ preset)  &  ndn3_13  &  n_n9186 ) | ( (~ preset)  &  nsr3_13  &  n_n9186 ) ;
 assign wire3474 = ( (~ preset)  &  nsr3_38  &  n_n7885 ) | ( (~ preset)  &  n_n7885  &  ndn3_38 ) ;
 assign wire3476 = ( (~ preset)  &  n_n7966  &  ndn3_37 ) | ( (~ preset)  &  n_n7966  &  nsr3_37 ) ;
 assign wire3480 = ( (~ preset)  &  ngfdn_3  &  n_n8081 ) | ( (~ preset)  &  n_n8081  &  (~ ndn3_46) ) ;
 assign wire3481 = ( n_n7098  &  (~ n_n8865)  &  wire4672 ) | ( n_n7098  &  (~ n_n8865)  &  wire4673 ) | ( n_n7098  &  n_n8865  &  (~ wire4672)  &  (~ wire4673) ) ;
 assign wire3482 = ( (~ preset)  &  ngfdn_3  &  n_n9219 ) | ( (~ preset)  &  n_n9219  &  (~ ndn3_46) ) ;
 assign wire3484 = ( (~ preset)  &  n_n9043  &  ndn3_37 ) | ( (~ preset)  &  n_n9043  &  nsr3_37 ) ;
 assign wire3489 = ( n_n7864  &  wire4421 ) | ( n_n7864  &  n_n8667  &  wire16682 ) ;
 assign wire3490 = ( n_n8933  &  wire2363  &  n_n8932 ) | ( (~ n_n8933)  &  wire2363  &  (~ n_n8932) ) ;
 assign wire3495 = ( (~ preset)  &  (~ ndn3_39)  &  n_n8100 ) | ( (~ preset)  &  n_n8100  &  ndn3_40 ) ;
 assign wire3496 = ( (~ preset)  &  n_n8871  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire3497 = ( (~ preset)  &  nsr3_14  &  n_n9266 ) | ( (~ preset)  &  n_n9266  &  ndn3_14 ) ;
 assign wire3501 = ( (~ preset)  &  ndn3_19  &  n_n7429 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n7429 ) ;
 assign wire3502 = ( (~ preset)  &  nrq3_19  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_19  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3505 = ( (~ preset)  &  n_n8791  &  ndn3_4 ) | ( (~ preset)  &  n_n8791  &  (~ ndn3_2) ) ;
 assign wire3506 = ( (~ preset)  &  nrq3_4  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_4  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3507 = ( (~ preset)  &  (~ nen3_39)  &  n_n7624 ) | ( (~ preset)  &  ndn3_39  &  n_n7624 ) ;
 assign wire3515 = ( (~ preset)  &  n_n9535  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9535  &  ndn3_44 ) ;
 assign wire3516 = ( (~ preset)  &  n_n9309  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire3517 = ( (~ preset)  &  ndn3_13  &  n_n8396 ) | ( (~ preset)  &  nsr3_13  &  n_n8396 ) ;
 assign wire3519 = ( (~ preset)  &  ndn3_7  &  n_n7813 ) | ( (~ preset)  &  n_n7813  &  (~ ndn3_4) ) ;
 assign wire3521 = ( (~ preset)  &  psv38_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3522 = ( (~ preset)  &  n_n7509  &  ndn3_2 ) | ( (~ preset)  &  n_n7509  &  (~ nen3_2) ) ;
 assign wire3525 = ( (~ preset)  &  ndn3_30  &  n_n7980 ) | ( (~ preset)  &  nsr3_30  &  n_n7980 ) ;
 assign wire3527 = ( (~ preset)  &  ndn3_23  &  n_n7667 ) | ( (~ preset)  &  nsr3_23  &  n_n7667 ) ;
 assign wire3529 = ( (~ preset)  &  n_n7761  &  nsr3_20 ) | ( (~ preset)  &  n_n7761  &  ndn3_20 ) ;
 assign wire3531 = ( (~ preset)  &  ndn3_25  &  n_n7683 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n7683 ) ;
 assign wire3532 = ( (~ preset)  &  ndn_latch3_25  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_25  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3535 = ( (~ preset)  &  ndn3_29  &  n_n8177 ) | ( (~ preset)  &  (~ ndn3_28)  &  n_n8177 ) ;
 assign wire3536 = ( (~ preset)  &  ndn_latch3_29  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_29  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3537 = ( (~ preset)  &  n_n7793  &  ndn3_4 ) | ( (~ preset)  &  n_n7793  &  (~ ndn3_2) ) ;
 assign wire3541 = ( (~ preset)  &  psv2_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3542 = ( (~ preset)  &  n_n7817  &  ndn3_2 ) | ( (~ preset)  &  n_n7817  &  (~ nen3_2) ) ;
 assign wire3545 = ( (~ preset)  &  n_n7225  &  nsr3_20 ) | ( (~ preset)  &  n_n7225  &  ndn3_20 ) ;
 assign wire3547 = ( (~ preset)  &  ndn3_30  &  n_n7808 ) | ( (~ preset)  &  nsr3_30  &  n_n7808 ) ;
 assign wire3549 = ( (~ preset)  &  n_n6963  &  ndn3_42 ) | ( (~ preset)  &  n_n6963  &  (~ ndn3_40) ) ;
 assign wire3550 = ( (~ preset)  &  n_n9155  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire3551 = ( (~ preset)  &  (~ nen3_22)  &  n_n7392 ) | ( (~ preset)  &  ndn3_22  &  n_n7392 ) ;
 assign wire3552 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9586 ) ;
 assign wire3553 = ( (~ preset)  &  psv33_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3554 = ( (~ preset)  &  n_n9302  &  ndn3_2 ) | ( (~ preset)  &  n_n9302  &  (~ nen3_2) ) ;
 assign wire3557 = ( (~ preset)  &  n_n9458  &  ndn3_34 ) | ( (~ preset)  &  n_n9458  &  (~ nen3_34) ) ;
 assign wire3565 = ( (~ preset)  &  n_n8801  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n8801  &  ndn3_44 ) ;
 assign wire3566 = ( (~ preset)  &  n_n8247  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire3567 = ( (~ preset)  &  psv18_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3568 = ( (~ preset)  &  n_n9396  &  ndn3_2 ) | ( (~ preset)  &  n_n9396  &  (~ nen3_2) ) ;
 assign wire3571 = ( (~ preset)  &  (~ nen3_22)  &  n_n7231 ) | ( (~ preset)  &  ndn3_22  &  n_n7231 ) ;
 assign wire3572 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n8093 ) ;
 assign wire3573 = ( (~ preset)  &  ndn3_30  &  n_n9312 ) | ( (~ preset)  &  nsr3_30  &  n_n9312 ) ;
 assign wire3575 = ( (~ preset)  &  (~ nen3_22)  &  n_n8856 ) | ( (~ preset)  &  ndn3_22  &  n_n8856 ) ;
 assign wire3576 = ( wire2367  &  (~ n_n7939)  &  wire5311 ) | ( wire2367  &  (~ n_n7939)  &  wire5312 ) | ( wire2367  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire3581 = ( (~ n_n8667)  &  (~ wire4421)  &  wire16729 ) | ( (~ wire4421)  &  (~ wire16682)  &  wire16729 ) ;
 assign wire3582 = ( n_n8603  &  (~ wire2363)  &  (~ wire15947)  &  (~ wire15948) ) ;
 assign wire3586 = ( n_n9434  &  n_n8880  &  wire16721 ) | ( n_n9434  &  n_n8431  &  wire16721 ) | ( n_n8880  &  n_n8431  &  wire16721 ) ;
 assign wire3587 = ( (~ n_n9416)  &  wire2395  &  (~ n_n8783)  &  n_n8784 ) | ( (~ n_n9416)  &  wire2395  &  n_n8783  &  (~ n_n8784) ) ;
 assign wire3588 = ( n_n9416  &  wire2363  &  (~ n_n8783)  &  (~ n_n8784) ) ;
 assign wire3589 = ( (~ preset)  &  n_n9416  &  (~ n_n7274) ) ;
 assign wire3590 = ( (~ preset)  &  psv39_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3591 = ( (~ preset)  &  n_n9324  &  ndn3_2 ) | ( (~ preset)  &  n_n9324  &  (~ nen3_2) ) ;
 assign wire3594 = ( (~ preset)  &  psv33_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3595 = ( (~ preset)  &  n_n9182  &  ndn3_2 ) | ( (~ preset)  &  n_n9182  &  (~ nen3_2) ) ;
 assign wire3600 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n9278 ) | ( (~ preset)  &  n_n9278  &  ndn3_50 ) ;
 assign wire3601 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n7781 ) ;
 assign wire3602 = ( (~ preset)  &  ndn3_9  &  n_n8014 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n8014 ) ;
 assign wire3604 = ( (~ preset)  &  ndn3_9  &  n_n8961 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n8961 ) ;
 assign wire3606 = ( (~ preset)  &  psv13_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3607 = ( (~ preset)  &  n_n7880  &  ndn3_2 ) | ( (~ preset)  &  n_n7880  &  (~ nen3_2) ) ;
 assign wire3610 = ( (~ preset)  &  psv13_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3611 = ( (~ preset)  &  n_n7766  &  ndn3_2 ) | ( (~ preset)  &  n_n7766  &  (~ nen3_2) ) ;
 assign wire3614 = ( (~ preset)  &  nsr3_13  &  n_n7687 ) | ( (~ preset)  &  ndn3_15  &  n_n7687 ) ;
 assign wire3615 = ( (~ preset)  &  nrq3_15  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_15  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3618 = ( (~ preset)  &  n_n7685  &  nsr3_20 ) | ( (~ preset)  &  n_n7685  &  ndn3_20 ) ;
 assign wire3620 = ( (~ preset)  &  ndn3_17  &  n_n8281 ) | ( (~ preset)  &  (~ ndn3_16)  &  n_n8281 ) ;
 assign wire3621 = ( (~ preset)  &  nrq3_17  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_17  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3622 = ( pinp_2_2_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3623 = ( (~ preset)  &  n_n8009  &  ndn3_2 ) | ( (~ preset)  &  n_n8009  &  (~ nen3_2) ) ;
 assign wire3624 = ( (~ preset)  &  ndn3_7  &  n_n7825 ) | ( (~ preset)  &  n_n7825  &  (~ ndn3_4) ) ;
 assign wire3625 = ( (~ preset)  &  ndn_latch3_7  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_7  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3630 = ( (~ preset)  &  nsr3_13  &  n_n7878 ) | ( (~ preset)  &  ndn3_15  &  n_n7878 ) ;
 assign wire3632 = ( (~ preset)  &  n_n7395  &  ndn3_42 ) | ( (~ preset)  &  n_n7395  &  (~ ndn3_40) ) ;
 assign wire3633 = ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40  &  n_n8206 ) ;
 assign wire3636 = ( (~ preset)  &  ndn3_28  &  n_n9327 ) | ( (~ preset)  &  n_n9327  &  (~ nen3_28) ) ;
 assign wire3638 = ( (~ preset)  &  ndn3_23  &  n_n9176 ) | ( (~ preset)  &  nsr3_23  &  n_n9176 ) ;
 assign wire3640 = ( (~ preset)  &  (~ ndn3_19)  &  n_n7756 ) | ( (~ preset)  &  ndn3_21  &  n_n7756 ) ;
 assign wire3644 = ( (~ preset)  &  (~ ndn3_19)  &  n_n8464 ) | ( (~ preset)  &  ndn3_21  &  n_n8464 ) ;
 assign wire3646 = ( (~ preset)  &  nsr3_35  &  n_n7734 ) | ( (~ preset)  &  n_n7734  &  ndn3_35 ) ;
 assign wire3648 = ( (~ preset)  &  psv26_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3649 = ( (~ preset)  &  n_n9500  &  ndn3_2 ) | ( (~ preset)  &  n_n9500  &  (~ nen3_2) ) ;
 assign wire3654 = ( (~ preset)  &  nsr3_35  &  n_n7650 ) | ( (~ preset)  &  n_n7650  &  ndn3_35 ) ;
 assign wire3656 = ( (~ preset)  &  nsr3_35  &  n_n7807 ) | ( (~ preset)  &  n_n7807  &  ndn3_35 ) ;
 assign wire3668 = ( (~ preset)  &  (~ nen3_39)  &  n_n8794 ) | ( (~ preset)  &  n_n8794  &  ndn3_39 ) ;
 assign wire3670 = ( (~ preset)  &  (~ nen3_22)  &  n_n7360 ) | ( (~ preset)  &  ndn3_22  &  n_n7360 ) ;
 assign wire3671 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n7756 ) ;
 assign wire3672 = ( (~ preset)  &  (~ ndn3_11)  &  n_n8984 ) | ( (~ preset)  &  n_n8984  &  ndn3_12 ) ;
 assign wire3676 = ( (~ preset)  &  (~ ndn3_11)  &  n_n9599 ) | ( (~ preset)  &  n_n9599  &  ndn3_12 ) ;
 assign wire3677 = ( (~ preset)  &  ndn_latch3_12  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_12  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3678 = ( (~ preset)  &  psv13_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3679 = ( (~ preset)  &  n_n7866  &  ndn3_2 ) | ( (~ preset)  &  n_n7866  &  (~ nen3_2) ) ;
 assign wire3684 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8486 ) | ( (~ preset)  &  n_n8486  &  ndn3_50 ) ;
 assign wire3685 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n9626 ) ;
 assign wire3686 = ( (~ preset)  &  psv18_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3687 = ( (~ preset)  &  n_n9314  &  ndn3_2 ) | ( (~ preset)  &  n_n9314  &  (~ nen3_2) ) ;
 assign wire3690 = ( (~ preset)  &  n_n8073  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8073  &  ndn3_40 ) ;
 assign wire3691 = ( (~ preset)  &  ndn3_39  &  n_n7624  &  (~ ndn3_40) ) ;
 assign wire3692 = ( (~ preset)  &  n_n7896  &  ndn3_46 ) | ( (~ preset)  &  n_n7896  &  (~ ndn3_44) ) ;
 assign wire3694 = ( pinp_9_9_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3695 = ( (~ preset)  &  n_n9349  &  ndn3_2 ) | ( (~ preset)  &  n_n9349  &  (~ nen3_2) ) ;
 assign wire3696 = ( (~ preset)  &  psv13_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3697 = ( (~ preset)  &  n_n9323  &  ndn3_2 ) | ( (~ preset)  &  n_n9323  &  (~ nen3_2) ) ;
 assign wire3700 = ( (~ preset)  &  pinp_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3701 = ( (~ preset)  &  n_n9183  &  ndn3_2 ) | ( (~ preset)  &  n_n9183  &  (~ nen3_2) ) ;
 assign wire3702 = ( (~ preset)  &  (~ nen3_22)  &  n_n8854 ) | ( (~ preset)  &  ndn3_22  &  n_n8854 ) ;
 assign wire3704 = ( pinp_3_3_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3705 = ( (~ preset)  &  n_n9137  &  ndn3_2 ) | ( (~ preset)  &  n_n9137  &  (~ nen3_2) ) ;
 assign wire3713 = ( (~ preset)  &  nsr3_13  &  n_n9319 ) | ( (~ preset)  &  ndn3_15  &  n_n9319 ) ;
 assign wire3714 = ( (~ preset)  &  nrq3_15  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_15  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3715 = ( n_n9353  &  n_n8484  &  wire16714 ) | ( n_n9353  &  n_n8807  &  wire16714 ) | ( n_n8484  &  n_n8807  &  wire16714 ) ;
 assign wire3719 = ( (~ preset)  &  ndn3_28  &  n_n9395 ) | ( (~ preset)  &  n_n9395  &  (~ nen3_28) ) ;
 assign wire3721 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7923 ) | ( (~ preset)  &  n_n7923  &  ndn3_50 ) ;
 assign wire3722 = ( (~ preset)  &  n_n7779  &  ngfdn_3  &  (~ ndn3_50) ) ;
 assign wire3723 = ( (~ preset)  &  ndn3_13  &  n_n8833 ) | ( (~ preset)  &  nsr3_13  &  n_n8833 ) ;
 assign wire3725 = ( (~ preset)  &  (~ ndn3_9)  &  n_n8276 ) | ( (~ preset)  &  ndn3_11  &  n_n8276 ) ;
 assign wire3726 = ( (~ preset)  &  nrq3_11  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_11  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3731 = ( (~ preset)  &  n_n7514  &  ndn3_46 ) | ( (~ preset)  &  n_n7514  &  (~ ndn3_44) ) ;
 assign wire3732 = ( (~ preset)  &  (~ ndn3_46)  &  n_n8188  &  ndn3_44 ) ;
 assign wire3733 = ( (~ preset)  &  psv33_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3734 = ( (~ preset)  &  n_n8456  &  ndn3_2 ) | ( (~ preset)  &  n_n8456  &  (~ nen3_2) ) ;
 assign wire3737 = ( (~ preset)  &  psv39_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3738 = ( (~ preset)  &  n_n8504  &  ndn3_2 ) | ( (~ preset)  &  n_n8504  &  (~ nen3_2) ) ;
 assign wire3741 = ( (~ preset)  &  ndn3_30  &  n_n7950 ) | ( (~ preset)  &  nsr3_30  &  n_n7950 ) ;
 assign wire3743 = ( (~ preset)  &  ndn3_25  &  n_n9315 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n9315 ) ;
 assign wire3744 = ( (~ preset)  &  ndn_latch3_25  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_25  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3745 = ( (~ preset)  &  (~ ndn3_17)  &  n_n8402 ) | ( (~ preset)  &  ndn3_18  &  n_n8402 ) ;
 assign wire3749 = ( (~ preset)  &  (~ nen3_22)  &  n_n7684 ) | ( (~ preset)  &  ndn3_22  &  n_n7684 ) ;
 assign wire3757 = ( (~ preset)  &  (~ nen3_36)  &  n_n8552 ) | ( (~ preset)  &  n_n8552  &  ndn3_36 ) ;
 assign wire3761 = ( (~ preset)  &  psv39_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3762 = ( (~ preset)  &  n_n7835  &  ndn3_2 ) | ( (~ preset)  &  n_n7835  &  (~ nen3_2) ) ;
 assign wire3765 = ( (~ preset)  &  psv2_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3766 = ( (~ preset)  &  n_n7689  &  ndn3_2 ) | ( (~ preset)  &  n_n7689  &  (~ nen3_2) ) ;
 assign wire3769 = ( (~ preset)  &  n_n9494  &  nsr3_20 ) | ( (~ preset)  &  n_n9494  &  ndn3_20 ) ;
 assign wire3773 = ( (~ preset)  &  ndn3_19  &  n_n8982 ) | ( (~ preset)  &  (~ nen3_19)  &  n_n8982 ) ;
 assign wire3775 = ( (~ preset)  &  n_n8095  &  nsr3_35 ) | ( (~ preset)  &  n_n8095  &  ndn3_35 ) ;
 assign wire3783 = ( (~ preset)  &  ndn3_30  &  n_n8900 ) | ( (~ preset)  &  nsr3_30  &  n_n8900 ) ;
 assign wire3787 = ( (~ preset)  &  n_n8210  &  nsr3_14 ) | ( (~ preset)  &  n_n8210  &  ndn3_14 ) ;
 assign wire3791 = ( (~ preset)  &  n_n8626  &  ndn3_34 ) | ( (~ preset)  &  n_n8626  &  (~ nen3_34) ) ;
 assign wire3792 = ( (~ preset)  &  nrq3_34  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_34  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3797 = ( (~ preset)  &  n_n7988  &  nsr3_35 ) | ( (~ preset)  &  n_n7988  &  ndn3_35 ) ;
 assign wire3799 = ( (~ preset)  &  (~ nen3_39)  &  n_n8906 ) | ( (~ preset)  &  n_n8906  &  ndn3_39 ) ;
 assign wire3800 = ( (~ preset)  &  nrq3_39  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_39  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3801 = ( (~ preset)  &  ndn3_9  &  n_n9268 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n9268 ) ;
 assign wire3802 = ( (~ preset)  &  nrq3_9  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_9  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3805 = ( (~ preset)  &  ndn3_17  &  n_n8983 ) | ( (~ preset)  &  n_n8983  &  (~ ndn3_16) ) ;
 assign wire3807 = ( (~ preset)  &  n_n7256  &  ndn3_46 ) | ( (~ preset)  &  n_n7256  &  (~ ndn3_44) ) ;
 assign wire3808 = ( (~ preset)  &  n_n9171  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire3809 = ( (~ preset)  &  ndn3_17  &  n_n8939 ) | ( (~ preset)  &  n_n8939  &  (~ ndn3_16) ) ;
 assign wire3810 = ( (~ preset)  &  nrq3_17  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_17  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3811 = ( (~ preset)  &  psv2_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3812 = ( (~ preset)  &  n_n8739  &  ndn3_2 ) | ( (~ preset)  &  n_n8739  &  (~ nen3_2) ) ;
 assign wire3817 = ( (~ preset)  &  n_n9366  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n9366  &  ndn3_40 ) ;
 assign wire3818 = ( (~ preset)  &  ndn3_39  &  n_n7464  &  (~ ndn3_40) ) ;
 assign wire3819 = ( (~ preset)  &  nsr3_38  &  n_n9310 ) | ( (~ preset)  &  n_n9310  &  ndn3_38 ) ;
 assign wire3821 = ( (~ preset)  &  n_n7570  &  ndn3_46 ) | ( (~ preset)  &  n_n7570  &  (~ ndn3_44) ) ;
 assign wire3822 = ( wire2370  &  (~ n_n8314)  &  wire5069 ) | ( wire2370  &  (~ n_n8314)  &  wire5070 ) | ( wire2370  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire3823 = ( (~ preset)  &  (~ ndn3_29)  &  n_n9470 ) | ( (~ preset)  &  n_n9470  &  ndn3_32 ) ;
 assign wire3824 = ( (~ preset)  &  ndn_latch3_32  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_32  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire3825 = ( (~ preset)  &  n_n9623  &  ndn3_42 ) | ( (~ preset)  &  n_n9623  &  (~ ndn3_40) ) ;
 assign wire3827 = ( (~ preset)  &  n_n9609  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n9609  &  ndn3_40 ) ;
 assign wire3829 = ( (~ preset)  &  psv2_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3830 = ( (~ preset)  &  n_n9325  &  ndn3_2 ) | ( (~ preset)  &  n_n9325  &  (~ nen3_2) ) ;
 assign wire3833 = ( (~ preset)  &  (~ nen3_16)  &  n_n9342 ) | ( (~ preset)  &  n_n9342  &  ndn3_16 ) ;
 assign wire3837 = ( pinp_1_1_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3838 = ( (~ preset)  &  n_n9054  &  ndn3_2 ) | ( (~ preset)  &  n_n9054  &  (~ nen3_2) ) ;
 assign wire3839 = ( (~ preset)  &  (~ nen3_22)  &  n_n7822 ) | ( (~ preset)  &  ndn3_22  &  n_n7822 ) ;
 assign wire3843 = ( (~ preset)  &  psv39_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3844 = ( (~ preset)  &  n_n9502  &  ndn3_2 ) | ( (~ preset)  &  n_n9502  &  (~ nen3_2) ) ;
 assign wire3847 = ( (~ preset)  &  ndn3_29  &  n_n8741 ) | ( (~ preset)  &  (~ ndn3_28)  &  n_n8741 ) ;
 assign wire3848 = ( (~ preset)  &  ndn_latch3_29  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_29  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3849 = ( (~ preset)  &  n_n9371  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n9371  &  ndn3_40 ) ;
 assign wire3850 = ( (~ preset)  &  n_n8611  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire3851 = ( (~ preset)  &  n_n8980  &  ndn3_34 ) | ( (~ preset)  &  n_n8980  &  (~ nen3_34) ) ;
 assign wire3853 = ( (~ preset)  &  psv26_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3854 = ( (~ preset)  &  n_n7743  &  ndn3_2 ) | ( (~ preset)  &  n_n7743  &  (~ nen3_2) ) ;
 assign wire3857 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n9429 ) | ( (~ preset)  &  n_n9429  &  ndn3_50 ) ;
 assign wire3858 = ( (~ preset)  &  ngfdn_3  &  n_n7217  &  (~ ndn3_50) ) ;
 assign wire3859 = ( (~ preset)  &  n_n6961  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n6961  &  ndn3_44 ) ;
 assign wire3860 = ( (~ preset)  &  n_n8989  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire3861 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8809 ) | ( (~ preset)  &  n_n8809  &  ndn3_26 ) ;
 assign wire3863 = ( (~ preset)  &  n_n8340  &  ndn3_46 ) | ( (~ preset)  &  n_n8340  &  (~ ndn3_44) ) ;
 assign wire3864 = ( (~ preset)  &  (~ ndn3_46)  &  n_n8468  &  ndn3_44 ) ;
 assign wire3865 = ( (~ preset)  &  psv39_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3866 = ( (~ preset)  &  n_n7936  &  ndn3_2 ) | ( (~ preset)  &  n_n7936  &  (~ nen3_2) ) ;
 assign wire3875 = ( (~ preset)  &  n_n8430  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8430  &  ndn3_40 ) ;
 assign wire3876 = ( (~ preset)  &  n_n9106  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire3877 = ( (~ preset)  &  (~ nen3_22)  &  n_n9596 ) | ( (~ preset)  &  ndn3_22  &  n_n9596 ) ;
 assign wire3879 = ( (~ preset)  &  (~ nen3_16)  &  n_n7876 ) | ( (~ preset)  &  n_n7876  &  ndn3_16 ) ;
 assign wire3886 = ( n_n9356  &  wire4421 ) | ( n_n9356  &  n_n8667  &  wire16682 ) ;
 assign wire3887 = ( n_n8911  &  n_n8933  &  wire2363 ) | ( n_n8911  &  wire2363  &  n_n8932 ) | ( (~ n_n8911)  &  (~ n_n8933)  &  wire2363  &  (~ n_n8932) ) ;
 assign wire3888 = ( (~ preset)  &  ndn3_25  &  n_n7887 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n7887 ) ;
 assign wire3889 = ( (~ preset)  &  ndn_latch3_25  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_25  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire3892 = ( (~ preset)  &  n_n8760  &  ndn3_4 ) | ( (~ preset)  &  n_n8760  &  (~ ndn3_2) ) ;
 assign wire3893 = ( (~ preset)  &  nrq3_4  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_4  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3894 = ( (~ preset)  &  ndn3_23  &  n_n9264 ) | ( (~ preset)  &  nsr3_23  &  n_n9264 ) ;
 assign wire3896 = ( (~ preset)  &  psv39_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3897 = ( (~ preset)  &  n_n7657  &  ndn3_2 ) | ( (~ preset)  &  n_n7657  &  (~ nen3_2) ) ;
 assign wire3902 = ( (~ preset)  &  n_n9102  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n9102  &  ndn3_40 ) ;
 assign wire3903 = ( wire2371  &  (~ n_n8320)  &  wire5184 ) | ( wire2371  &  (~ n_n8320)  &  wire5185 ) | ( wire2371  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire3904 = ( (~ preset)  &  n_n9316  &  nsr3_20 ) | ( (~ preset)  &  n_n9316  &  ndn3_20 ) ;
 assign wire3906 = ( (~ preset)  &  ndn3_30  &  n_n7929 ) | ( (~ preset)  &  nsr3_30  &  n_n7929 ) ;
 assign wire3908 = ( (~ preset)  &  n_n7962  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n7962  &  ndn3_40 ) ;
 assign wire3909 = ( wire2371  &  (~ n_n9478)  &  wire5338 ) | ( wire2371  &  (~ n_n9478)  &  wire5339 ) | ( wire2371  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire3910 = ( (~ preset)  &  psv18_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3911 = ( (~ preset)  &  n_n7930  &  ndn3_2 ) | ( (~ preset)  &  n_n7930  &  (~ nen3_2) ) ;
 assign wire3914 = ( (~ preset)  &  (~ ndn3_29)  &  n_n8864 ) | ( (~ preset)  &  n_n8864  &  ndn3_32 ) ;
 assign wire3918 = ( n_n9448  &  n_n8323  &  wire16707 ) | ( n_n9448  &  n_n8324  &  wire16707 ) | ( n_n8323  &  n_n8324  &  wire16707 ) ;
 assign wire3919 = ( (~ n_n8354)  &  wire2395  &  (~ n_n8353)  &  n_n8355 ) | ( (~ n_n8354)  &  wire2395  &  n_n8353  &  (~ n_n8355) ) ;
 assign wire3920 = ( n_n8354  &  wire2363  &  (~ n_n8353)  &  (~ n_n8355) ) ;
 assign wire3921 = ( (~ preset)  &  n_n8354  &  (~ n_n7274) ) ;
 assign wire3928 = ( (~ preset)  &  (~ nen3_36)  &  n_n7789 ) | ( (~ preset)  &  n_n7789  &  ndn3_36 ) ;
 assign wire3930 = ( (~ preset)  &  (~ nen3_39)  &  n_n8543 ) | ( (~ preset)  &  n_n8543  &  ndn3_39 ) ;
 assign wire3931 = ( (~ preset)  &  nrq3_39  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_39  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire3932 = ( (~ preset)  &  n_n8480  &  ndn3_37 ) | ( (~ preset)  &  n_n8480  &  nsr3_37 ) ;
 assign wire3936 = ( (~ preset)  &  nsr3_38  &  n_n9487 ) | ( (~ preset)  &  n_n9487  &  ndn3_38 ) ;
 assign wire3938 = ( (~ preset)  &  (~ nen3_36)  &  n_n7967 ) | ( (~ preset)  &  n_n7967  &  ndn3_36 ) ;
 assign wire3940 = ( (~ preset)  &  ndn3_17  &  n_n8744 ) | ( (~ preset)  &  n_n8744  &  (~ ndn3_16) ) ;
 assign wire3941 = ( (~ preset)  &  nrq3_17  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_17  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3942 = ( (~ preset)  &  n_n8022  &  ndn3_42 ) | ( (~ preset)  &  n_n8022  &  (~ ndn3_40) ) ;
 assign wire3943 = ( wire2368  &  (~ n_n8314)  &  wire5069 ) | ( wire2368  &  (~ n_n8314)  &  wire5070 ) | ( wire2368  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire3944 = ( (~ preset)  &  ndn3_30  &  n_n9592 ) | ( (~ preset)  &  nsr3_30  &  n_n9592 ) ;
 assign wire3949 = ( (~ preset)  &  ndn3_29  &  n_n8808 ) | ( (~ preset)  &  (~ ndn3_28)  &  n_n8808 ) ;
 assign wire3951 = ( (~ preset)  &  (~ nen3_36)  &  n_n9044 ) | ( (~ preset)  &  n_n9044  &  ndn3_36 ) ;
 assign wire3952 = ( (~ preset)  &  nrq3_36  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_36  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire3953 = ( (~ preset)  &  psv39_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3954 = ( (~ preset)  &  n_n9407  &  ndn3_2 ) | ( (~ preset)  &  n_n9407  &  (~ nen3_2) ) ;
 assign wire3964 = ( (~ preset)  &  n_n9132  &  nsr3_14 ) | ( (~ preset)  &  n_n9132  &  ndn3_14 ) ;
 assign wire3966 = ( (~ preset)  &  n_n9337  &  ndn3_27 ) | ( (~ preset)  &  n_n9337  &  (~ ndn3_26) ) ;
 assign wire3968 = ( (~ preset)  &  ngfdn_3  &  n_n8589 ) | ( (~ preset)  &  n_n8589  &  (~ ndn3_46) ) ;
 assign wire3969 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46  &  n_n9221 ) ;
 assign wire3972 = ( (~ preset)  &  (~ ndn3_17)  &  n_n7603 ) | ( (~ preset)  &  ndn3_18  &  n_n7603 ) ;
 assign wire3973 = ( (~ preset)  &  nrq3_18  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_18  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire3975 = ( n_n8963  &  wire4421 ) | ( n_n8963  &  n_n8667  &  wire16682 ) ;
 assign wire3976 = ( n_n8913  &  n_n8964  &  wire2363 ) | ( n_n8964  &  wire2363  &  n_n8493 ) | ( (~ n_n8913)  &  (~ n_n8964)  &  wire2363  &  (~ n_n8493) ) ;
 assign wire3977 = ( (~ preset)  &  psv38_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3978 = ( (~ preset)  &  n_n8638  &  ndn3_2 ) | ( (~ preset)  &  n_n8638  &  (~ nen3_2) ) ;
 assign wire3981 = ( (~ preset)  &  (~ nen3_22)  &  n_n7017 ) | ( (~ preset)  &  ndn3_22  &  n_n7017 ) ;
 assign wire3982 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9087 ) ;
 assign wire3983 = ( (~ preset)  &  ndn3_25  &  n_n9397 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n9397 ) ;
 assign wire3989 = ( (~ preset)  &  nsr3_13  &  n_n8519 ) | ( (~ preset)  &  n_n8519  &  ndn3_15 ) ;
 assign wire3991 = ( (~ preset)  &  (~ nen3_22)  &  n_n9368 ) | ( (~ preset)  &  ndn3_22  &  n_n9368 ) ;
 assign wire3993 = ( (~ preset)  &  n_n8750  &  ndn3_42 ) | ( (~ preset)  &  n_n8750  &  (~ ndn3_40) ) ;
 assign wire3994 = ( (~ preset)  &  n_n7962  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire3995 = ( (~ preset)  &  ndn3_23  &  n_n7968 ) | ( (~ preset)  &  nsr3_23  &  n_n7968 ) ;
 assign wire3997 = ( pinp_14_14_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire3998 = ( (~ preset)  &  n_n8000  &  ndn3_2 ) | ( (~ preset)  &  n_n8000  &  (~ nen3_2) ) ;
 assign wire4001 = ( pinp_11_11_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4002 = ( (~ preset)  &  n_n8986  &  ndn3_2 ) | ( (~ preset)  &  n_n8986  &  (~ nen3_2) ) ;
 assign wire4003 = ( (~ preset)  &  ndn3_28  &  n_n7820 ) | ( (~ preset)  &  n_n7820  &  (~ nen3_28) ) ;
 assign wire4004 = ( (~ preset)  &  ndn_latch3_28  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_28  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4007 = ( (~ preset)  &  n_n9333  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9333  &  ndn3_44 ) ;
 assign wire4008 = ( wire2369  &  (~ n_n8320)  &  wire5184 ) | ( wire2369  &  (~ n_n8320)  &  wire5185 ) | ( wire2369  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire4009 = ( (~ preset)  &  ndn3_23  &  n_n9047 ) | ( (~ preset)  &  nsr3_23  &  n_n9047 ) ;
 assign wire4013 = ( (~ preset)  &  ndn3_19  &  n_n8810 ) | ( (~ preset)  &  n_n8810  &  (~ nen3_19) ) ;
 assign wire4015 = ( (~ preset)  &  n_n8381  &  nsr3_14 ) | ( (~ preset)  &  n_n8381  &  ndn3_14 ) ;
 assign wire4017 = ( (~ preset)  &  n_n9041  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9041  &  ndn3_44 ) ;
 assign wire4019 = ( (~ preset)  &  (~ ndn3_19)  &  n_n8093 ) | ( (~ preset)  &  n_n8093  &  ndn3_21 ) ;
 assign wire4020 = ( (~ preset)  &  nrq3_21  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_21  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire4021 = ( (~ preset)  &  n_n7102  &  ndn3_42 ) | ( (~ preset)  &  n_n7102  &  (~ ndn3_40) ) ;
 assign wire4022 = ( (~ preset)  &  n_n9609  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4027 = ( n_n8449  &  n_n8450  &  wire16690 ) | ( n_n8449  &  n_n8448  &  wire16690 ) | ( n_n8450  &  n_n8448  &  wire16690 ) ;
 assign wire4028 = ( (~ n_n8549)  &  wire2395  &  (~ n_n8522)  &  n_n8521 ) | ( (~ n_n8549)  &  wire2395  &  n_n8522  &  (~ n_n8521) ) ;
 assign wire4029 = ( n_n8549  &  wire2363  &  (~ n_n8522)  &  (~ n_n8521) ) ;
 assign wire4030 = ( (~ preset)  &  n_n8549  &  (~ n_n7274) ) ;
 assign wire4033 = ( (~ preset)  &  nsr3_38  &  n_n7681 ) | ( (~ preset)  &  n_n7681  &  ndn3_38 ) ;
 assign wire4037 = ( (~ preset)  &  ndn3_9  &  n_n9346 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n9346 ) ;
 assign wire4041 = ( (~ preset)  &  psv38_9_9_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4042 = ( (~ preset)  &  n_n9336  &  ndn3_2 ) | ( (~ preset)  &  n_n9336  &  (~ nen3_2) ) ;
 assign wire4045 = ( (~ preset)  &  ndn3_9  &  n_n9134 ) | ( (~ preset)  &  (~ ndn3_7)  &  n_n9134 ) ;
 assign wire4047 = ( (~ preset)  &  psv18_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4048 = ( (~ preset)  &  n_n9491  &  ndn3_2 ) | ( (~ preset)  &  n_n9491  &  (~ nen3_2) ) ;
 assign wire4051 = ( (~ preset)  &  (~ ndn3_29)  &  n_n9334 ) | ( (~ preset)  &  n_n9334  &  ndn3_32 ) ;
 assign wire4053 = ( (~ preset)  &  psv38_1_1_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4054 = ( (~ preset)  &  n_n9045  &  ndn3_2 ) | ( (~ preset)  &  n_n9045  &  (~ nen3_2) ) ;
 assign wire4059 = ( (~ preset)  &  ngfdn_3  &  n_n9282 ) | ( (~ preset)  &  n_n9282  &  (~ ndn3_46) ) ;
 assign wire4071 = ( (~ preset)  &  ndn3_23  &  n_n8697 ) | ( (~ preset)  &  nsr3_23  &  n_n8697 ) ;
 assign wire4073 = ( (~ preset)  &  n_n7875  &  nsr3_20 ) | ( (~ preset)  &  n_n7875  &  ndn3_20 ) ;
 assign wire4075 = ( (~ preset)  &  n_n9036  &  ndn3_42 ) | ( (~ preset)  &  n_n9036  &  (~ ndn3_40) ) ;
 assign wire4077 = ( (~ preset)  &  n_n7527  &  ndn3_46 ) | ( (~ preset)  &  n_n7527  &  (~ ndn3_44) ) ;
 assign wire4081 = ( (~ preset)  &  n_n7454  &  ndn3_19 ) | ( (~ preset)  &  n_n7454  &  (~ nen3_19) ) ;
 assign wire4083 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8369 ) | ( (~ preset)  &  n_n8369  &  ndn3_50 ) ;
 assign wire4084 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n9508 ) ;
 assign wire4085 = ( (~ preset)  &  n_n9263  &  ndn3_27 ) | ( (~ preset)  &  n_n9263  &  (~ ndn3_26) ) ;
 assign wire4086 = ( (~ preset)  &  ndn_latch3_27  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_27  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire4087 = ( (~ preset)  &  n_n8153  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n8153  &  ndn3_12 ) ;
 assign wire4088 = ( (~ preset)  &  ndn_latch3_12  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_12  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4091 = ( (~ preset)  &  ngfdn_3  &  n_n9004 ) | ( (~ preset)  &  n_n9004  &  (~ ndn3_46) ) ;
 assign wire4092 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8951  &  ndn3_46 ) ;
 assign wire4093 = ( (~ preset)  &  n_n8049  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n8049  &  ndn3_44 ) ;
 assign wire4094 = ( (~ preset)  &  n_n9589  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4099 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n9148 ) | ( (~ preset)  &  n_n9148  &  ndn3_50 ) ;
 assign wire4100 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n7606 ) ;
 assign wire4101 = ( (~ preset)  &  n_n7498  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7498  &  ndn3_44 ) ;
 assign wire4102 = ( (~ preset)  &  n_n9391  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4103 = ( (~ preset)  &  n_n7824  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n7824  &  ndn3_12 ) ;
 assign wire4104 = ( (~ preset)  &  ndn_latch3_12  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_12  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4105 = ( (~ preset)  &  (~ nen3_22)  &  n_n7777 ) | ( (~ preset)  &  ndn3_22  &  n_n7777 ) ;
 assign wire4106 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9100 ) ;
 assign wire4107 = ( (~ preset)  &  psv13_4_4_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4108 = ( (~ preset)  &  n_n7826  &  ndn3_2 ) | ( (~ preset)  &  n_n7826  &  (~ nen3_2) ) ;
 assign wire4113 = ( (~ preset)  &  n_n8777  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8777  &  ndn3_40 ) ;
 assign wire4114 = ( (~ preset)  &  ndn3_39  &  (~ ndn3_40)  &  n_n8858 ) ;
 assign wire4117 = ( (~ preset)  &  psv33_10_10_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4118 = ( (~ preset)  &  n_n9300  &  ndn3_2 ) | ( (~ preset)  &  n_n9300  &  (~ nen3_2) ) ;
 assign wire4123 = ( (~ preset)  &  (~ ndn3_17)  &  n_n7847 ) | ( (~ preset)  &  ndn3_18  &  n_n7847 ) ;
 assign wire4124 = ( (~ preset)  &  nrq3_18  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_18  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4125 = ( (~ preset)  &  (~ nen3_22)  &  n_n7760 ) | ( (~ preset)  &  ndn3_22  &  n_n7760 ) ;
 assign wire4129 = ( (~ preset)  &  ngfdn_3  &  n_n8466 ) | ( (~ preset)  &  n_n8466  &  (~ ndn3_46) ) ;
 assign wire4133 = ( (~ preset)  &  ndn3_23  &  n_n7911 ) | ( (~ preset)  &  nsr3_23  &  n_n7911 ) ;
 assign wire4135 = ( (~ preset)  &  n_n8582  &  ndn3_19 ) | ( (~ preset)  &  n_n8582  &  (~ nen3_19) ) ;
 assign wire4139 = ( (~ preset)  &  n_n7790  &  ndn3_27 ) | ( (~ preset)  &  n_n7790  &  (~ ndn3_26) ) ;
 assign wire4141 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8279 ) | ( (~ preset)  &  n_n8279  &  ndn3_26 ) ;
 assign wire4142 = ( (~ preset)  &  ndn_latch3_26  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_26  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4143 = ( (~ preset)  &  psv2_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4144 = ( (~ preset)  &  n_n9387  &  ndn3_2 ) | ( (~ preset)  &  n_n9387  &  (~ nen3_2) ) ;
 assign wire4147 = ( (~ preset)  &  n_n9589  &  ndn3_42 ) | ( (~ preset)  &  n_n9589  &  (~ ndn3_40) ) ;
 assign wire4149 = ( (~ preset)  &  n_n8951  &  ndn3_46 ) | ( (~ preset)  &  n_n8951  &  (~ ndn3_44) ) ;
 assign wire4151 = ( (~ preset)  &  n_n9573  &  ndn3_46 ) | ( (~ preset)  &  n_n9573  &  (~ ndn3_44) ) ;
 assign wire4152 = ( wire2370  &  (~ n_n9478)  &  wire5338 ) | ( wire2370  &  (~ n_n9478)  &  wire5339 ) | ( wire2370  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire4155 = ( (~ preset)  &  n_n8659  &  nsr3_14 ) | ( (~ preset)  &  n_n8659  &  ndn3_14 ) ;
 assign wire4157 = ( (~ preset)  &  n_n8681  &  ndn3_42 ) | ( (~ preset)  &  n_n8681  &  (~ ndn3_40) ) ;
 assign wire4158 = ( (~ preset)  &  n_n8996  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4159 = ( (~ preset)  &  n_n8042  &  nsr3_14 ) | ( (~ preset)  &  n_n8042  &  ndn3_14 ) ;
 assign wire4161 = ( (~ preset)  &  ndn3_29  &  n_n8941 ) | ( (~ preset)  &  n_n8941  &  (~ ndn3_28) ) ;
 assign wire4163 = ( (~ preset)  &  psv33_6_6_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4164 = ( (~ preset)  &  n_n7643  &  ndn3_2 ) | ( (~ preset)  &  n_n7643  &  (~ nen3_2) ) ;
 assign wire4171 = ( (~ preset)  &  ngfdn_3  &  n_n7775 ) | ( (~ preset)  &  n_n7775  &  (~ ndn3_46) ) ;
 assign wire4172 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46  &  n_n7083 ) ;
 assign wire4173 = ( (~ preset)  &  ngfdn_3  &  n_n9096 ) | ( (~ preset)  &  n_n9096  &  (~ ndn3_46) ) ;
 assign wire4174 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n8258  &  ndn3_46 ) ;
 assign wire4175 = ( (~ preset)  &  ndn3_13  &  n_n9189 ) | ( (~ preset)  &  n_n9189  &  nsr3_13 ) ;
 assign wire4177 = ( (~ preset)  &  (~ ndn3_17)  &  n_n9341 ) | ( (~ preset)  &  ndn3_18  &  n_n9341 ) ;
 assign wire4179 = ( (~ preset)  &  ndn3_13  &  n_n8260 ) | ( (~ preset)  &  n_n8260  &  nsr3_13 ) ;
 assign wire4181 = ( (~ preset)  &  n_n7918  &  nsr3_38 ) | ( (~ preset)  &  n_n7918  &  ndn3_38 ) ;
 assign wire4183 = ( (~ preset)  &  n_n8996  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8996  &  ndn3_40 ) ;
 assign wire4185 = ( (~ preset)  &  n_n7806  &  nsr3_38 ) | ( (~ preset)  &  n_n7806  &  ndn3_38 ) ;
 assign wire4187 = ( (~ preset)  &  n_n8024  &  ndn3_42 ) | ( (~ preset)  &  n_n8024  &  (~ ndn3_40) ) ;
 assign wire4189 = ( (~ preset)  &  n_n8678  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n8678  &  ndn3_44 ) ;
 assign wire4190 = ( (~ preset)  &  n_n7948  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4191 = ( (~ preset)  &  n_n9432  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9432  &  ndn3_44 ) ;
 assign wire4192 = ( (~ preset)  &  n_n9036  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4193 = ( (~ preset)  &  psv38_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4194 = ( (~ preset)  &  n_n9174  &  ndn3_2 ) | ( (~ preset)  &  n_n9174  &  (~ nen3_2) ) ;
 assign wire4197 = ( (~ preset)  &  n_n7757  &  ndn3_42 ) | ( (~ preset)  &  n_n7757  &  (~ ndn3_40) ) ;
 assign wire4199 = ( (~ preset)  &  n_n7831  &  ndn3_30 ) | ( (~ preset)  &  n_n7831  &  nsr3_30 ) ;
 assign wire4201 = ( (~ preset)  &  psv13_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4202 = ( (~ preset)  &  n_n9501  &  ndn3_2 ) | ( (~ preset)  &  n_n9501  &  (~ nen3_2) ) ;
 assign wire4205 = ( (~ preset)  &  n_n8445  &  nsr3_38 ) | ( (~ preset)  &  n_n8445  &  ndn3_38 ) ;
 assign wire4207 = ( (~ preset)  &  psv2_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4208 = ( (~ preset)  &  n_n9408  &  ndn3_2 ) | ( (~ preset)  &  n_n9408  &  (~ nen3_2) ) ;
 assign wire4211 = ( (~ preset)  &  n_n9489  &  ndn3_30 ) | ( (~ preset)  &  n_n9489  &  nsr3_30 ) ;
 assign wire4213 = ( (~ preset)  &  ndn3_25  &  n_n7821 ) | ( (~ preset)  &  (~ ndn3_22)  &  n_n7821 ) ;
 assign wire4214 = ( (~ preset)  &  ndn_latch3_25  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_25  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4215 = ( (~ preset)  &  ngfdn_3  &  n_n7217 ) | ( (~ preset)  &  n_n7217  &  (~ ndn3_46) ) ;
 assign wire4220 = ( (~ preset)  &  n_n9321  &  ndn3_7 ) | ( (~ preset)  &  n_n9321  &  (~ ndn3_4) ) ;
 assign wire4221 = ( (~ preset)  &  ndn_latch3_7  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_7  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire4222 = ( (~ preset)  &  n_n8843  &  nsr3_20 ) | ( (~ preset)  &  n_n8843  &  ndn3_20 ) ;
 assign wire4224 = ( (~ preset)  &  ndn3_23  &  n_n7641 ) | ( (~ preset)  &  n_n7641  &  nsr3_23 ) ;
 assign wire4226 = ( (~ preset)  &  n_n8258  &  ndn3_46 ) | ( (~ preset)  &  n_n8258  &  (~ ndn3_44) ) ;
 assign wire4228 = ( (~ preset)  &  n_n8247  &  ndn3_42 ) | ( (~ preset)  &  n_n8247  &  (~ ndn3_40) ) ;
 assign wire4230 = ( (~ preset)  &  n_n8957  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8957  &  ndn3_40 ) ;
 assign wire4232 = ( (~ preset)  &  n_n8959  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8959  &  ndn3_40 ) ;
 assign wire4233 = ( wire2371  &  (~ n_n7939)  &  wire5311 ) | ( wire2371  &  (~ n_n7939)  &  wire5312 ) | ( wire2371  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire4234 = ( (~ preset)  &  psv26_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4235 = ( (~ preset)  &  n_n7954  &  ndn3_2 ) | ( (~ preset)  &  n_n7954  &  (~ nen3_2) ) ;
 assign wire4238 = ( (~ preset)  &  ndn3_13  &  n_n9601 ) | ( (~ preset)  &  n_n9601  &  nsr3_13 ) ;
 assign wire4240 = ( (~ preset)  &  n_n9465  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9465  &  ndn3_44 ) ;
 assign wire4241 = ( (~ preset)  &  n_n8022  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4242 = ( (~ preset)  &  psv26_0_0_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4243 = ( (~ preset)  &  n_n7656  &  ndn3_2 ) | ( (~ preset)  &  n_n7656  &  (~ nen3_2) ) ;
 assign wire4246 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8998 ) | ( (~ preset)  &  n_n8998  &  ndn3_26 ) ;
 assign wire4248 = ( (~ preset)  &  n_n8282  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n8282  &  ndn3_12 ) ;
 assign wire4249 = ( (~ preset)  &  ndn_latch3_12  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_12  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4250 = ( (~ preset)  &  ngfdn_3  &  n_n7546 ) | ( (~ preset)  &  n_n7546  &  (~ ndn3_46) ) ;
 assign wire4251 = ( (~ preset)  &  n_n9235  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign wire4254 = ( (~ preset)  &  n_n7174  &  ndn3_46 ) | ( (~ preset)  &  n_n7174  &  (~ ndn3_44) ) ;
 assign wire4255 = ( (~ preset)  &  (~ ndn3_46)  &  ndn3_44  &  n_n9632 ) ;
 assign wire4256 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8742 ) | ( (~ preset)  &  n_n8742  &  ndn3_26 ) ;
 assign wire4257 = ( (~ preset)  &  ndn_latch3_26  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  ndn_latch3_26  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire4258 = ( (~ preset)  &  n_n8006  &  ndn3_7 ) | ( (~ preset)  &  n_n8006  &  (~ ndn3_4) ) ;
 assign wire4260 = ( (~ preset)  &  psv13_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4261 = ( (~ preset)  &  n_n8414  &  ndn3_2 ) | ( (~ preset)  &  n_n8414  &  (~ nen3_2) ) ;
 assign wire4264 = ( (~ preset)  &  psv13_8_8_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4265 = ( (~ preset)  &  n_n7955  &  ndn3_2 ) | ( (~ preset)  &  n_n7955  &  (~ nen3_2) ) ;
 assign wire4272 = ( (~ preset)  &  n_n7160  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n7160  &  ndn3_40 ) ;
 assign wire4273 = ( (~ preset)  &  n_n8906  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire4274 = ( (~ preset)  &  psv33_13_13_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4275 = ( (~ preset)  &  n_n9098  &  ndn3_2 ) | ( (~ preset)  &  n_n9098  &  (~ nen3_2) ) ;
 assign wire4278 = ( (~ preset)  &  (~ ndn3_29)  &  n_n7640 ) | ( (~ preset)  &  n_n7640  &  ndn3_32 ) ;
 assign wire4280 = ( (~ preset)  &  n_n7803  &  ndn3_7 ) | ( (~ preset)  &  n_n7803  &  (~ ndn3_4) ) ;
 assign wire4281 = ( (~ preset)  &  ndn_latch3_7  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_7  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4282 = ( (~ preset)  &  psv33_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4283 = ( (~ preset)  &  n_n8086  &  ndn3_2 ) | ( (~ preset)  &  n_n8086  &  (~ nen3_2) ) ;
 assign wire4288 = ( (~ preset)  &  (~ nen3_22)  &  n_n9339 ) | ( (~ preset)  &  ndn3_22  &  n_n9339 ) ;
 assign wire4289 = ( wire2367  &  (~ n_n8320)  &  wire5184 ) | ( wire2367  &  (~ n_n8320)  &  wire5185 ) | ( wire2367  &  n_n8320  &  (~ wire5184)  &  (~ wire5185) ) ;
 assign wire4290 = ( pinp_4_4_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4291 = ( (~ preset)  &  n_n8736  &  ndn3_2 ) | ( (~ preset)  &  n_n8736  &  (~ nen3_2) ) ;
 assign wire4292 = ( (~ preset)  &  n_n8005  &  (~ nen3_16) ) | ( (~ preset)  &  n_n8005  &  ndn3_16 ) ;
 assign wire4294 = ( (~ preset)  &  n_n7823  &  (~ nen3_16) ) | ( (~ preset)  &  n_n7823  &  ndn3_16 ) ;
 assign wire4295 = ( (~ preset)  &  nrq3_16  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_16  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4296 = ( (~ preset)  &  (~ ndn3_25)  &  n_n8545 ) | ( (~ preset)  &  n_n8545  &  ndn3_26 ) ;
 assign wire4297 = ( (~ preset)  &  ndn_latch3_26  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  ndn_latch3_26  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4302 = ( (~ preset)  &  n_n8219  &  nsr3_20 ) | ( (~ preset)  &  n_n8219  &  ndn3_20 ) ;
 assign wire4304 = ( (~ preset)  &  n_n7236  &  (~ ndn3_19) ) | ( (~ preset)  &  n_n7236  &  ndn3_21 ) ;
 assign wire4310 = ( (~ preset)  &  ndn3_29  &  n_n7428 ) | ( (~ preset)  &  n_n7428  &  (~ ndn3_28) ) ;
 assign wire4311 = ( (~ preset)  &  ndn_latch3_29  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  ndn_latch3_29  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4314 = ( (~ preset)  &  n_n9597  &  nsr3_20 ) | ( (~ preset)  &  n_n9597  &  ndn3_20 ) ;
 assign wire4316 = ( pinp_10_10_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4317 = ( (~ preset)  &  n_n8110  &  ndn3_2 ) | ( (~ preset)  &  n_n8110  &  (~ nen3_2) ) ;
 assign wire4318 = ( (~ preset)  &  n_n9391  &  ndn3_42 ) | ( (~ preset)  &  n_n9391  &  (~ ndn3_40) ) ;
 assign wire4319 = ( wire2368  &  (~ n_n9478)  &  wire5338 ) | ( wire2368  &  (~ n_n9478)  &  wire5339 ) | ( wire2368  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire4320 = ( (~ preset)  &  n_n7758  &  ndn3_30 ) | ( (~ preset)  &  n_n7758  &  nsr3_30 ) ;
 assign wire4322 = ( (~ preset)  &  ndn3_29  &  n_n8278 ) | ( (~ preset)  &  n_n8278  &  (~ ndn3_28) ) ;
 assign wire4323 = ( (~ preset)  &  ndn_latch3_29  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_29  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4326 = ( (~ preset)  &  n_n9125  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9125  &  ndn3_44 ) ;
 assign wire4327 = ( wire2369  &  (~ n_n9478)  &  wire5338 ) | ( wire2369  &  (~ n_n9478)  &  wire5339 ) | ( wire2369  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire4328 = ( (~ preset)  &  n_n9169  &  ndn3_42 ) | ( (~ preset)  &  n_n9169  &  (~ ndn3_40) ) ;
 assign wire4329 = ( (~ preset)  &  (~ ndn3_42)  &  ndn3_40  &  n_n6974 ) ;
 assign wire4330 = ( (~ preset)  &  psv38_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4331 = ( (~ preset)  &  n_n9223  &  ndn3_2 ) | ( (~ preset)  &  n_n9223  &  (~ nen3_2) ) ;
 assign wire4344 = ( (~ preset)  &  n_n9135  &  ndn3_4 ) | ( (~ preset)  &  n_n9135  &  (~ ndn3_2) ) ;
 assign wire4346 = ( (~ preset)  &  n_n7898  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7898  &  ndn3_44 ) ;
 assign wire4350 = ( (~ preset)  &  n_n8765  &  ndn3_46 ) | ( (~ preset)  &  n_n8765  &  (~ ndn3_44) ) ;
 assign wire4352 = ( (~ preset)  &  n_n7908  &  ndn3_37 ) | ( (~ preset)  &  n_n7908  &  nsr3_37 ) ;
 assign wire4354 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7462 ) | ( (~ preset)  &  n_n7462  &  ndn3_50 ) ;
 assign wire4355 = ( (~ preset)  &  ngfdn_3  &  n_n9219  &  (~ ndn3_50) ) ;
 assign wire4358 = ( (~ preset)  &  n_n7384  &  ndn3_46 ) | ( (~ preset)  &  n_n7384  &  (~ ndn3_44) ) ;
 assign wire4360 = ( (~ preset)  &  n_n9613  &  (~ nen3_39) ) | ( (~ preset)  &  n_n9613  &  ndn3_39 ) ;
 assign wire4361 = ( (~ preset)  &  nrq3_39  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_39  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4364 = ( (~ preset)  &  psv13_3_3_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4365 = ( (~ preset)  &  n_n9406  &  ndn3_2 ) | ( (~ preset)  &  n_n9406  &  (~ nen3_2) ) ;
 assign wire4370 = ( (~ preset)  &  n_n9611  &  (~ nen3_39) ) | ( (~ preset)  &  n_n9611  &  ndn3_39 ) ;
 assign wire4372 = ( (~ preset)  &  ngfdn_3  &  n_n7324 ) | ( (~ preset)  &  n_n7324  &  (~ ndn3_46) ) ;
 assign wire4374 = ( (~ preset)  &  n_n9335  &  ndn3_37 ) | ( (~ preset)  &  n_n9335  &  nsr3_37 ) ;
 assign wire4376 = ( (~ preset)  &  n_n9127  &  ndn3_37 ) | ( (~ preset)  &  n_n9127  &  nsr3_37 ) ;
 assign wire4378 = ( (~ preset_0_0_)  &  (~ ngfdn_3)  &  nsr1_2 ) | ( (~ ngfdn_3)  &  nsr1_2  &  nlc1_2 ) ;
 assign wire4380 = ( (~ preset)  &  n_n9400  &  (~ nen3_16) ) | ( (~ preset)  &  n_n9400  &  ndn3_16 ) ;
 assign wire4382 = ( (~ preset)  &  n_n9343  &  nsr3_13 ) | ( (~ preset)  &  n_n9343  &  ndn3_15 ) ;
 assign wire4384 = ( (~ preset)  &  n_n7054  &  ndn3_42 ) | ( (~ preset)  &  n_n7054  &  (~ ndn3_40) ) ;
 assign wire4385 = ( (~ preset)  &  n_n9576  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4386 = ( (~ preset)  &  n_n7948  &  ndn3_42 ) | ( (~ preset)  &  n_n7948  &  (~ ndn3_40) ) ;
 assign wire4388 = ( (~ preset)  &  n_n7783  &  ndn3_46 ) | ( (~ preset)  &  n_n7783  &  (~ ndn3_44) ) ;
 assign wire4389 = ( wire2370  &  (~ n_n7939)  &  wire5311 ) | ( wire2370  &  (~ n_n7939)  &  wire5312 ) | ( wire2370  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire4390 = ( (~ preset)  &  ndn3_23  &  n_n7602 ) | ( (~ preset)  &  n_n7602  &  nsr3_23 ) ;
 assign wire4392 = ( (~ preset)  &  n_n7740  &  nsr3_20 ) | ( (~ preset)  &  n_n7740  &  ndn3_20 ) ;
 assign wire4394 = ( (~ preset)  &  n_n7691  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7691  &  ndn3_44 ) ;
 assign wire4396 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n9483 ) | ( (~ preset)  &  n_n9483  &  ndn3_50 ) ;
 assign wire4397 = ( (~ preset)  &  ngfdn_3  &  (~ ndn3_50)  &  n_n8948 ) ;
 assign wire4398 = ( (~ preset)  &  n_n9049  &  nsr3_14 ) | ( (~ preset)  &  n_n9049  &  ndn3_14 ) ;
 assign wire4400 = ( (~ preset)  &  n_n9588  &  ndn3_34 ) | ( (~ preset)  &  n_n9588  &  (~ nen3_34) ) ;
 assign wire4401 = ( (~ preset)  &  nrq3_34  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_34  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire4404 = ( (~ preset)  &  (~ ndn3_9)  &  n_n7791 ) | ( (~ preset)  &  n_n7791  &  ndn3_11 ) ;
 assign wire4406 = ( (~ preset)  &  n_n7857  &  ndn3_46 ) | ( (~ preset)  &  n_n7857  &  (~ ndn3_44) ) ;
 assign wire4407 = ( (~ preset)  &  n_n7706  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire4411 = ( n_n8630  &  wire4421 ) | ( n_n8630  &  n_n8667  &  wire16682 ) ;
 assign wire4412 = ( n_n8631  &  n_n8561  &  wire2363 ) | ( n_n8631  &  wire2363  &  n_n8342 ) | ( (~ n_n8631)  &  (~ n_n8561)  &  wire2363  &  (~ n_n8342) ) ;
 assign wire4416 = ( n_n9056  &  wire4421 ) | ( n_n9056  &  n_n8667  &  wire16682 ) ;
 assign wire4417 = ( n_n8913  &  wire2363  &  n_n8493 ) | ( (~ n_n8913)  &  wire2363  &  (~ n_n8493) ) ;
 assign wire4421 = ( (~ preset)  &  (~ n_n9247)  &  n_n9639  &  wire16469 ) ;
 assign wire4424 = ( (~ preset)  &  psv13_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4425 = ( (~ preset)  &  n_n8114  &  ndn3_2 ) | ( (~ preset)  &  n_n8114  &  (~ nen3_2) ) ;
 assign wire4428 = ( (~ preset)  &  psv39_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4429 = ( (~ preset)  &  n_n8491  &  ndn3_2 ) | ( (~ preset)  &  n_n8491  &  (~ nen3_2) ) ;
 assign wire4432 = ( (~ preset)  &  (~ nen3_22)  &  n_n8175 ) | ( (~ preset)  &  n_n8175  &  ndn3_22 ) ;
 assign wire4433 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9252 ) ;
 assign wire4434 = ( (~ preset)  &  ndn3_13  &  n_n9257 ) | ( (~ preset)  &  n_n9257  &  nsr3_13 ) ;
 assign wire4436 = ( (~ preset)  &  n_n8091  &  (~ ngfdn_3) ) | ( (~ preset)  &  n_n8091  &  ndn3_50 ) ;
 assign wire4437 = ( (~ preset)  &  ngfdn_3  &  n_n8466  &  (~ ndn3_50) ) ;
 assign wire4440 = ( (~ preset)  &  n_n8066  &  nsr3_14 ) | ( (~ preset)  &  n_n8066  &  ndn3_14 ) ;
 assign wire4444 = ( (~ preset)  &  psv13_2_2_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4445 = ( (~ preset)  &  n_n8053  &  ndn3_2 ) | ( (~ preset)  &  n_n8053  &  (~ nen3_2) ) ;
 assign wire4448 = ( (~ preset)  &  n_n7811  &  nsr3_13 ) | ( (~ preset)  &  n_n7811  &  ndn3_15 ) ;
 assign wire4450 = ( (~ preset)  &  ndn3_13  &  n_n7934 ) | ( (~ preset)  &  n_n7934  &  nsr3_13 ) ;
 assign wire4452 = ( (~ preset)  &  n_n7735  &  ndn3_30 ) | ( (~ preset)  &  n_n7735  &  nsr3_30 ) ;
 assign wire4456 = ( (~ preset)  &  n_n7651  &  ndn3_30 ) | ( (~ preset)  &  n_n7651  &  nsr3_30 ) ;
 assign wire4460 = ( (~ preset)  &  n_n9412  &  (~ ndn3_19) ) | ( (~ preset)  &  n_n9412  &  ndn3_21 ) ;
 assign wire4462 = ( (~ preset)  &  (~ nen3_22)  &  n_n9398 ) | ( (~ preset)  &  n_n9398  &  ndn3_22 ) ;
 assign wire4463 = ( wire2367  &  (~ n_n9478)  &  wire5338 ) | ( wire2367  &  (~ n_n9478)  &  wire5339 ) | ( wire2367  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire4464 = ( (~ preset)  &  n_n9064  &  nsr3_20 ) | ( (~ preset)  &  n_n9064  &  ndn3_20 ) ;
 assign wire4468 = ( (~ preset)  &  psv2_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4469 = ( (~ preset)  &  n_n8007  &  ndn3_2 ) | ( (~ preset)  &  n_n8007  &  (~ nen3_2) ) ;
 assign wire4472 = ( pinp_15_15_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4473 = ( (~ preset)  &  n_n8482  &  ndn3_2 ) | ( (~ preset)  &  n_n8482  &  (~ nen3_2) ) ;
 assign wire4474 = ( (~ preset)  &  psv2_14_14_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4475 = ( (~ preset)  &  n_n7937  &  ndn3_2 ) | ( (~ preset)  &  n_n7937  &  (~ nen3_2) ) ;
 assign wire4480 = ( pinp_13_13_  &  (~ preset)  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4481 = ( (~ preset)  &  n_n7850  &  ndn3_2 ) | ( (~ preset)  &  n_n7850  &  (~ nen3_2) ) ;
 assign wire4488 = ( n_n9512  &  n_n8734  &  wire16676 ) | ( n_n9512  &  n_n8733  &  wire16676 ) | ( n_n8734  &  n_n8733  &  wire16676 ) ;
 assign wire4489 = ( (~ n_n9434)  &  wire2395  &  (~ n_n8880)  &  n_n8431 ) | ( (~ n_n9434)  &  wire2395  &  n_n8880  &  (~ n_n8431) ) ;
 assign wire4490 = ( n_n9434  &  wire2363  &  (~ n_n8880)  &  (~ n_n8431) ) ;
 assign wire4491 = ( (~ preset)  &  n_n9434  &  (~ n_n7274) ) ;
 assign wire4494 = ( (~ preset)  &  n_n9399  &  nsr3_20 ) | ( (~ preset)  &  n_n9399  &  ndn3_20 ) ;
 assign wire4496 = ( (~ preset)  &  n_n8333  &  ndn3_28 ) | ( (~ preset)  &  n_n8333  &  (~ nen3_28) ) ;
 assign wire4497 = ( (~ preset)  &  ndn_latch3_28  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_28  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4498 = ( (~ preset)  &  psv18_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4499 = ( (~ preset)  &  n_n7759  &  ndn3_2 ) | ( (~ preset)  &  n_n7759  &  (~ nen3_2) ) ;
 assign wire4502 = ( (~ preset)  &  n_n8661  &  nsr3_14 ) | ( (~ preset)  &  n_n8661  &  ndn3_14 ) ;
 assign wire4504 = ( (~ preset)  &  n_n8132  &  ndn3_42 ) | ( (~ preset)  &  n_n8132  &  (~ ndn3_40) ) ;
 assign wire4505 = ( (~ preset)  &  n_n8150  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4508 = ( (~ preset)  &  n_n8488  &  (~ nen3_22) ) | ( (~ preset)  &  n_n8488  &  ndn3_22 ) ;
 assign wire4509 = ( (~ preset)  &  nen3_22  &  n_n9412  &  (~ ndn3_22) ) ;
 assign wire4510 = ( (~ preset)  &  ndn3_13  &  n_n7953 ) | ( (~ preset)  &  n_n7953  &  nsr3_13 ) ;
 assign wire4518 = ( (~ preset)  &  n_n7179  &  ngfdn_3 ) | ( (~ preset)  &  n_n7179  &  (~ ndn3_46) ) ;
 assign wire4519 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7783  &  ndn3_46 ) ;
 assign wire4520 = ( (~ preset)  &  n_n9265  &  (~ ndn3_17) ) | ( (~ preset)  &  n_n9265  &  ndn3_18 ) ;
 assign wire4521 = ( (~ preset)  &  nrq3_18  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_18  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire4522 = ( (~ preset)  &  n_n9052  &  ndn3_4 ) | ( (~ preset)  &  n_n9052  &  (~ ndn3_2) ) ;
 assign wire4523 = ( (~ preset)  &  nrq3_4  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_4  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire4526 = ( (~ preset)  &  n_n9106  &  (~ nen3_39) ) | ( (~ preset)  &  n_n9106  &  ndn3_39 ) ;
 assign wire4527 = ( (~ preset)  &  nrq3_39  &  (~ n_n9385)  &  n_n9384 ) | ( (~ preset)  &  nrq3_39  &  n_n9385  &  (~ n_n9384) ) ;
 assign wire4530 = ( (~ preset)  &  n_n8702  &  (~ nen3_22) ) | ( (~ preset)  &  n_n8702  &  ndn3_22 ) ;
 assign wire4531 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n8213 ) ;
 assign wire4532 = ( (~ preset)  &  n_n7190  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7190  &  ndn3_44 ) ;
 assign wire4533 = ( (~ preset)  &  n_n8249  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4534 = ( (~ preset)  &  n_n9635  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n9635  &  ndn3_44 ) ;
 assign wire4535 = ( wire2369  &  (~ n_n8314)  &  wire5069 ) | ( wire2369  &  (~ n_n8314)  &  wire5070 ) | ( wire2369  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire4536 = ( (~ preset)  &  n_n8001  &  nsr3_38 ) | ( (~ preset)  &  n_n8001  &  ndn3_38 ) ;
 assign wire4538 = ( (~ preset)  &  n_n9000  &  ndn3_25 ) | ( (~ preset)  &  n_n9000  &  (~ ndn3_22) ) ;
 assign wire4544 = ( (~ preset)  &  n_n9598  &  (~ nen3_16) ) | ( (~ preset)  &  n_n9598  &  ndn3_16 ) ;
 assign wire4545 = ( (~ preset)  &  nrq3_16  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_16  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire4546 = ( (~ preset)  &  n_n8786  &  ndn3_7 ) | ( (~ preset)  &  n_n8786  &  (~ ndn3_4) ) ;
 assign wire4548 = ( (~ preset)  &  n_n9602  &  ndn3_7 ) | ( (~ preset)  &  n_n9602  &  (~ ndn3_4) ) ;
 assign wire4549 = ( (~ preset)  &  ndn_latch3_7  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  ndn_latch3_7  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire4582 = ( (~ preset)  &  n_n8981  &  ndn3_29 ) | ( (~ preset)  &  n_n8981  &  (~ ndn3_28) ) ;
 assign wire4588 = ( (~ preset)  &  n_n8308  &  ndn3_46 ) | ( (~ preset)  &  n_n8308  &  (~ ndn3_44) ) ;
 assign wire4590 = ( (~ preset)  &  n_n8609  &  ndn3_42 ) | ( (~ preset)  &  n_n8609  &  (~ ndn3_40) ) ;
 assign wire4591 = ( wire2368  &  (~ n_n7939)  &  wire5311 ) | ( wire2368  &  (~ n_n7939)  &  wire5312 ) | ( wire2368  &  n_n7939  &  (~ wire5311)  &  (~ wire5312) ) ;
 assign wire4592 = ( (~ preset)  &  n_n8699  &  nsr3_20 ) | ( (~ preset)  &  n_n8699  &  ndn3_20 ) ;
 assign wire4594 = ( (~ preset)  &  ndn3_23  &  n_n8533 ) | ( (~ preset)  &  n_n8533  &  nsr3_23 ) ;
 assign wire4598 = ( (~ preset)  &  n_n9273  &  (~ ndn3_19) ) | ( (~ preset)  &  n_n9273  &  ndn3_21 ) ;
 assign wire4600 = ( (~ preset)  &  n_n9311  &  nsr3_35 ) | ( (~ preset)  &  n_n9311  &  ndn3_35 ) ;
 assign wire4602 = ( (~ preset)  &  n_n7148  &  (~ ndn3_42) ) | ( (~ preset)  &  n_n7148  &  ndn3_44 ) ;
 assign wire4603 = ( (~ preset)  &  n_n9623  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4606 = ( (~ preset)  &  n_n8227  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n8227  &  ndn3_12 ) ;
 assign wire4614 = ( (~ preset)  &  n_n7970  &  (~ ndn3_9) ) | ( (~ preset)  &  n_n7970  &  ndn3_11 ) ;
 assign wire4618 = ( (~ preset)  &  n_n7581  &  (~ nen3_22) ) | ( (~ preset)  &  n_n7581  &  ndn3_22 ) ;
 assign wire4619 = ( (~ preset)  &  nen3_22  &  (~ ndn3_22)  &  n_n9351 ) ;
 assign wire4620 = ( (~ preset)  &  n_n9008  &  ndn3_9 ) | ( (~ preset)  &  n_n9008  &  (~ ndn3_7) ) ;
 assign wire4621 = ( (~ preset)  &  nrq3_9  &  (~ n_n7869)  &  n_n8028 ) | ( (~ preset)  &  nrq3_9  &  n_n7869  &  (~ n_n8028) ) ;
 assign wire4624 = ( (~ preset)  &  psv26_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4625 = ( (~ preset)  &  n_n7814  &  ndn3_2 ) | ( (~ preset)  &  n_n7814  &  (~ nen3_2) ) ;
 assign wire4628 = ( (~ preset)  &  n_n7877  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n7877  &  ndn3_12 ) ;
 assign wire4630 = ( (~ preset)  &  psv26_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4631 = ( (~ preset)  &  n_n7765  &  ndn3_2 ) | ( (~ preset)  &  n_n7765  &  (~ nen3_2) ) ;
 assign wire4634 = ( (~ preset)  &  n_n8758  &  ndn3_7 ) | ( (~ preset)  &  n_n8758  &  (~ ndn3_4) ) ;
 assign wire4635 = ( (~ preset)  &  ndn_latch3_7  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  ndn_latch3_7  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4636 = ( (~ preset)  &  n_n7332  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n7332  &  ndn3_40 ) ;
 assign wire4637 = ( (~ preset)  &  ndn3_39  &  (~ ndn3_40)  &  n_n8991 ) ;
 assign wire4640 = ( (~ preset)  &  psv39_12_12_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4641 = ( (~ preset)  &  n_n7816  &  ndn3_2 ) | ( (~ preset)  &  n_n7816  &  (~ nen3_2) ) ;
 assign wire4644 = ( (~ preset)  &  n_n7812  &  ndn3_13 ) | ( (~ preset)  &  n_n7812  &  nsr3_13 ) ;
 assign wire4646 = ( (~ preset)  &  n_n8394  &  ndn3_13 ) | ( (~ preset)  &  n_n8394  &  nsr3_13 ) ;
 assign wire4648 = ( (~ preset)  &  n_n8152  &  ndn3_17 ) | ( (~ preset)  &  n_n8152  &  (~ ndn3_16) ) ;
 assign wire4649 = ( (~ preset)  &  nrq3_17  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_17  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4650 = ( (~ preset)  &  n_n8597  &  (~ ndn3_17) ) | ( (~ preset)  &  n_n8597  &  ndn3_18 ) ;
 assign wire4651 = ( (~ preset)  &  nrq3_18  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_18  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4652 = ( (~ preset)  &  n_n7889  &  nsr3_13 ) | ( (~ preset)  &  n_n7889  &  ndn3_15 ) ;
 assign wire4653 = ( (~ preset)  &  nrq3_15  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_15  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4654 = ( (~ preset)  &  n_n7888  &  (~ nen3_16) ) | ( (~ preset)  &  n_n7888  &  ndn3_16 ) ;
 assign wire4655 = ( (~ preset)  &  nrq3_16  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_16  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4660 = ( (~ preset)  &  n_n8225  &  ndn3_19 ) | ( (~ preset)  &  n_n8225  &  (~ nen3_19) ) ;
 assign wire4662 = ( (~ preset)  &  n_n7599  &  ndn3_37 ) | ( (~ preset)  &  n_n7599  &  nsr3_37 ) ;
 assign wire4664 = ( (~ preset)  &  n_n7558  &  ngfdn_3 ) | ( (~ preset)  &  n_n7558  &  (~ ndn3_46) ) ;
 assign wire4665 = ( n_n7098  &  (~ n_n9478)  &  wire5338 ) | ( n_n7098  &  (~ n_n9478)  &  wire5339 ) | ( n_n7098  &  n_n9478  &  (~ wire5338)  &  (~ wire5339) ) ;
 assign wire4666 = ( (~ preset)  &  n_n8377  &  ndn3_7 ) | ( (~ preset)  &  n_n8377  &  (~ ndn3_4) ) ;
 assign wire4668 = ( (~ preset)  &  n_n8208  &  (~ ndn3_17) ) | ( (~ preset)  &  n_n8208  &  ndn3_18 ) ;
 assign wire4672 = ( n_n7543  &  n_n8126  &  n_n8125 ) | ( n_n7543  &  n_n7544  &  (~ n_n8126)  &  n_n8125 ) | ( n_n7543  &  n_n7544  &  n_n8126  &  (~ n_n8125) ) ;
 assign wire4673 = ( wire16639  &  wire16656 ) | ( wire16640  &  wire16656 ) | ( wire16639  &  wire16657 ) | ( wire16640  &  wire16657 ) ;
 assign wire4678 = ( n_n9568  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n9568 ) ;
 assign wire4679 = ( n_n8772  &  wire16030 ) | ( (~ ndn3_17)  &  n_n8772  &  ndn3_16 ) ;
 assign wire4684 = ( (~ ndn3_7)  &  ndn3_4  &  n_n7914 ) ;
 assign wire4685 = ( ndn3_11  &  (~ ndn3_12)  &  n_n7913 ) ;
 assign wire4686 = ( n_n7908  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4687 = ( (~ ndn3_27)  &  n_n7932  &  ndn3_26 ) ;
 assign wire4688 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n9632 ) ;
 assign wire4689 = ( nen3_16  &  (~ ndn3_16)  &  n_n8535 ) ;
 assign wire4690 = ( ndn3_29  &  n_n7910  &  (~ ndn3_32) ) ;
 assign wire4691 = ( n_n7909  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire4692 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7912 ) ;
 assign wire4693 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7911 ) ;
 assign wire4694 = ( n_n8512  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire4695 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8106 ) ;
 assign wire4696 = ( n_n7935  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n7935 ) ;
 assign wire4697 = ( n_n7936  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n7936 ) ;
 assign wire4701 = ( n_n7937  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire4702 = ( nen3_39  &  (~ ndn3_39)  &  n_n7928 ) ;
 assign wire4703 = ( (~ ndn3_9)  &  n_n8114  &  ndn3_7 ) ;
 assign wire4704 = ( (~ ngfdn_3)  &  n_n9108  &  ndn3_46 ) ;
 assign wire4705 = ( ndn3_9  &  (~ ndn3_11)  &  n_n7946 ) ;
 assign wire4706 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7933 ) ;
 assign wire4707 = ( n_n7931  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire4708 = ( (~ ndn3_46)  &  ndn3_44  &  n_n7927 ) ;
 assign wire4709 = ( n_n8445  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4710 = ( (~ ndn3_34)  &  n_n8425  &  nen3_34 ) ;
 assign wire4711 = ( nen3_36  &  n_n7929  &  (~ ndn3_36) ) ;
 assign wire4712 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8516 ) ;
 assign wire4713 = ( nen3_22  &  (~ ndn3_22)  &  n_n8219 ) ;
 assign wire4714 = ( n_n7934  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire4717 = ( n_n7971  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n7971 ) ;
 assign wire4718 = ( n_n8014  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n8014 ) ;
 assign wire4723 = ( (~ ndn3_7)  &  n_n8456  &  ndn3_4 ) ;
 assign wire4724 = ( n_n7970  &  ndn3_11  &  (~ ndn3_12) ) ;
 assign wire4725 = ( n_n7966  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4726 = ( (~ ndn3_27)  &  n_n8004  &  ndn3_26 ) ;
 assign wire4727 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8468 ) ;
 assign wire4728 = ( nen3_16  &  (~ ndn3_16)  &  n_n7969 ) ;
 assign wire4729 = ( ndn3_29  &  n_n9077  &  (~ ndn3_32) ) ;
 assign wire4730 = ( n_n7967  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire4731 = ( n_n8208  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire4732 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7968 ) ;
 assign wire4733 = ( n_n8864  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire4734 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8519 ) ;
 assign wire4735 = ( n_n8006  &  wire16047 ) | ( n_n8006  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire4736 = ( n_n8491  &  wire16048 ) | ( (~ ndn3_25)  &  n_n8491  &  ndn3_22 ) ;
 assign wire4740 = ( n_n8007  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire4741 = ( nen3_39  &  (~ ndn3_39)  &  n_n8078 ) ;
 assign wire4742 = ( (~ ndn3_9)  &  ndn3_7  &  n_n8502 ) ;
 assign wire4743 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8580 ) ;
 assign wire4744 = ( ndn3_9  &  (~ ndn3_11)  &  n_n8192 ) ;
 assign wire4745 = ( n_n8005  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire4746 = ( (~ ndn3_28)  &  n_n8003  &  nen3_28 ) ;
 assign wire4747 = ( (~ ndn3_46)  &  n_n9355  &  ndn3_44 ) ;
 assign wire4748 = ( n_n8001  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4749 = ( (~ ndn3_34)  &  n_n8839  &  nen3_34 ) ;
 assign wire4750 = ( nen3_36  &  n_n8900  &  (~ ndn3_36) ) ;
 assign wire4751 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8584 ) ;
 assign wire4752 = ( nen3_22  &  (~ ndn3_22)  &  n_n8064 ) ;
 assign wire4753 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n8344 ) ;
 assign wire4760 = ( (~ preset)  &  n_n8775  &  ndn3_4 ) | ( (~ preset)  &  n_n8775  &  (~ ndn3_2) ) ;
 assign wire4761 = ( (~ preset)  &  nrq3_4  &  (~ n_n7311)  &  n_n7544 ) | ( (~ preset)  &  nrq3_4  &  n_n7311  &  (~ n_n7544) ) ;
 assign wire4768 = ( n_n8758  &  wire16047 ) | ( n_n8758  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire4769 = ( n_n8504  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n8504 ) ;
 assign wire4773 = ( (~ ndn3_4)  &  n_n7890  &  ndn3_2 ) ;
 assign wire4774 = ( nen3_39  &  n_n7988  &  (~ ndn3_39) ) ;
 assign wire4775 = ( (~ ndn3_9)  &  n_n8414  &  ndn3_7 ) ;
 assign wire4776 = ( (~ ngfdn_3)  &  n_n8626  &  ndn3_46 ) ;
 assign wire4777 = ( ndn3_9  &  (~ ndn3_11)  &  n_n9067 ) ;
 assign wire4778 = ( n_n7888  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire4779 = ( (~ ndn3_28)  &  n_n7887  &  nen3_28 ) ;
 assign wire4780 = ( n_n9623  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire4781 = ( n_n7885  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire4782 = ( n_n8333  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire4783 = ( nen3_36  &  (~ ndn3_36)  &  n_n9092 ) ;
 assign wire4784 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8282 ) ;
 assign wire4785 = ( nen3_22  &  n_n9064  &  (~ ndn3_22) ) ;
 assign wire4786 = ( n_n8394  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire4787 = ( n_n8775  &  wire16029 ) | ( n_n8775  &  nen3_22  &  (~ ndn3_22) ) ;
 assign wire4788 = ( n_n7849  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n7849 ) ;
 assign wire4793 = ( n_n9098  &  (~ ndn3_7)  &  ndn3_4 ) ;
 assign wire4794 = ( ndn3_11  &  (~ ndn3_12)  &  n_n7848 ) ;
 assign wire4795 = ( n_n8480  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4796 = ( (~ ndn3_27)  &  n_n9520  &  ndn3_26 ) ;
 assign wire4797 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8470 ) ;
 assign wire4798 = ( nen3_16  &  (~ ndn3_16)  &  n_n8909 ) ;
 assign wire4799 = ( ndn3_29  &  n_n7845  &  (~ ndn3_32) ) ;
 assign wire4800 = ( ndn3_39  &  (~ ndn3_40)  &  n_n7844 ) ;
 assign wire4801 = ( n_n7847  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire4802 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7846 ) ;
 assign wire4803 = ( (~ ndn3_46)  &  n_n8277  &  ndn3_44 ) ;
 assign wire4804 = ( n_n7889  &  ndn3_17  &  (~ ndn3_18) ) ;
 assign wire4805 = ( (~ preset)  &  n_n7452  &  ndn3_29 ) | ( (~ preset)  &  n_n7452  &  (~ ndn3_28) ) ;
 assign wire4809 = ( n_n8821  &  n_n8820  &  wire16554 ) | ( n_n8821  &  n_n8822  &  wire16554 ) | ( n_n8820  &  n_n8822  &  wire16554 ) ;
 assign wire4810 = ( (~ n_n9638)  &  wire2395  &  (~ n_n8979)  &  n_n7432 ) | ( (~ n_n9638)  &  wire2395  &  n_n8979  &  (~ n_n7432) ) ;
 assign wire4811 = ( n_n9638  &  wire2363  &  (~ n_n8979)  &  (~ n_n7432) ) ;
 assign wire4812 = ( (~ preset)  &  n_n9638  &  (~ n_n7274) ) ;
 assign wire4817 = ( (~ preset)  &  n_n7522  &  ndn3_42 ) | ( (~ preset)  &  n_n7522  &  (~ ndn3_40) ) ;
 assign wire4818 = ( (~ preset)  &  n_n9102  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire4819 = ( (~ preset)  &  n_n9235  &  ndn3_46 ) | ( (~ preset)  &  n_n9235  &  (~ ndn3_44) ) ;
 assign wire4821 = ( (~ preset)  &  n_n9486  &  ndn3_42 ) | ( (~ preset)  &  n_n9486  &  (~ ndn3_40) ) ;
 assign wire4823 = ( (~ preset)  &  ndn3_23  &  n_n9130 ) | ( (~ preset)  &  n_n9130  &  nsr3_23 ) ;
 assign wire4827 = ( (~ preset)  &  psv38_11_11_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4828 = ( (~ preset)  &  n_n7709  &  ndn3_2 ) | ( (~ preset)  &  n_n7709  &  (~ nen3_2) ) ;
 assign wire4833 = ( (~ preset)  &  n_n7819  &  nsr3_35 ) | ( (~ preset)  &  n_n7819  &  ndn3_35 ) ;
 assign wire4843 = ( (~ preset)  &  psv18_15_15_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire4844 = ( (~ preset)  &  n_n8002  &  ndn3_2 ) | ( (~ preset)  &  n_n8002  &  (~ nen3_2) ) ;
 assign wire4847 = ( (~ preset)  &  n_n9467  &  ndn3_34 ) | ( (~ preset)  &  n_n9467  &  (~ nen3_34) ) ;
 assign wire4848 = ( (~ preset)  &  nrq3_34  &  (~ n_n7566)  &  n_n8154 ) | ( (~ preset)  &  nrq3_34  &  n_n7566  &  (~ n_n8154) ) ;
 assign wire4851 = ( (~ preset)  &  n_n9548  &  ngfdn_3 ) | ( (~ preset)  &  n_n9548  &  (~ ndn3_46) ) ;
 assign wire4852 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7384  &  ndn3_46 ) ;
 assign wire4857 = ( (~ preset)  &  n_n7707  &  ndn3_37 ) | ( (~ preset)  &  n_n7707  &  nsr3_37 ) ;
 assign wire4861 = ( (~ preset)  &  n_n8557  &  (~ n_n7274) ) ;
 assign wire4864 = ( nsr3_13  &  ndn3_12  &  n_n8584 ) | ( (~ nsr3_13)  &  nsr3_14  &  n_n8584 ) ;
 assign wire4865 = ( ndn3_17  &  n_n8583  &  nsr3_20 ) ;
 assign wire4866 = ( ndn3_29  &  n_n8941  &  nsr3_35 ) ;
 assign wire4867 = ( n_n8864  &  nsr3_37  &  nen3_34 ) ;
 assign wire4868 = ( nsr3_30  &  n_n8581  &  ndn3_26 ) ;
 assign wire4869 = ( nsr3_38  &  nen3_36  &  n_n8580 ) ;
 assign wire4870 = ( nsr3_23  &  n_n8582  &  ndn3_19 ) ;
 assign wire4877 = ( n_n8227  &  nsr3_13  &  ndn3_12 ) | ( n_n8227  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4878 = ( ndn3_17  &  nsr3_20  &  n_n8226 ) ;
 assign wire4879 = ( ndn3_29  &  nsr3_35  &  n_n8224 ) ;
 assign wire4880 = ( n_n8223  &  nsr3_37  &  nen3_34 ) ;
 assign wire4881 = ( nsr3_30  &  n_n9205  &  ndn3_26 ) ;
 assign wire4882 = ( nsr3_38  &  nen3_36  &  n_n8222 ) ;
 assign wire4883 = ( n_n8225  &  nsr3_23  &  ndn3_19 ) ;
 assign wire4886 = ( n_n8203  &  nsr3_13  &  ndn3_12 ) | ( n_n8203  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4887 = ( ndn3_17  &  n_n9019  &  nsr3_20 ) ;
 assign wire4888 = ( ndn3_29  &  nsr3_35  &  n_n8201 ) ;
 assign wire4889 = ( n_n9110  &  nsr3_37  &  nen3_34 ) ;
 assign wire4890 = ( nsr3_30  &  n_n9615  &  ndn3_26 ) ;
 assign wire4891 = ( nsr3_38  &  nen3_36  &  n_n9516 ) ;
 assign wire4892 = ( n_n8202  &  nsr3_23  &  ndn3_19 ) ;
 assign wire4899 = ( n_n7951  &  nsr3_13  &  ndn3_12 ) | ( n_n7951  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4900 = ( ndn3_17  &  n_n8753  &  nsr3_20 ) ;
 assign wire4901 = ( ndn3_29  &  n_n7474  &  nsr3_35 ) ;
 assign wire4902 = ( n_n9518  &  nsr3_37  &  nen3_34 ) ;
 assign wire4903 = ( nsr3_30  &  n_n9286  &  ndn3_26 ) ;
 assign wire4904 = ( nsr3_38  &  nen3_36  &  n_n7947 ) ;
 assign wire4905 = ( nsr3_23  &  ndn3_19  &  n_n7588 ) ;
 assign wire4918 = ( n_n9141  &  nsr3_13  &  ndn3_12 ) | ( n_n9141  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4919 = ( ndn3_17  &  n_n7375  &  nsr3_20 ) ;
 assign wire4920 = ( n_n7373  &  ndn3_29  &  nsr3_35 ) ;
 assign wire4921 = ( n_n8499  &  nsr3_37  &  nen3_34 ) ;
 assign wire4922 = ( nsr3_30  &  n_n7487  &  ndn3_26 ) ;
 assign wire4923 = ( nsr3_38  &  nen3_36  &  n_n8135 ) ;
 assign wire4924 = ( nsr3_23  &  ndn3_19  &  n_n7374 ) ;
 assign wire4927 = ( n_n9015  &  nsr3_13  &  ndn3_12 ) | ( n_n9015  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4928 = ( ndn3_17  &  n_n8104  &  nsr3_20 ) ;
 assign wire4929 = ( ndn3_29  &  nsr3_35  &  n_n8828 ) ;
 assign wire4930 = ( n_n7670  &  nsr3_37  &  nen3_34 ) ;
 assign wire4931 = ( n_n7341  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4932 = ( n_n8862  &  nsr3_38  &  nen3_36 ) ;
 assign wire4933 = ( nsr3_23  &  ndn3_19  &  n_n7342 ) ;
 assign wire4934 = ( nsr3_13  &  ndn3_12  &  n_n9318 ) | ( (~ nsr3_13)  &  nsr3_14  &  n_n9318 ) ;
 assign wire4935 = ( ndn3_17  &  n_n8744  &  nsr3_20 ) ;
 assign wire4936 = ( ndn3_29  &  n_n8741  &  nsr3_35 ) ;
 assign wire4937 = ( n_n9042  &  nsr3_37  &  nen3_34 ) ;
 assign wire4938 = ( n_n8742  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4939 = ( nsr3_38  &  nen3_36  &  n_n9308 ) ;
 assign wire4940 = ( nsr3_23  &  ndn3_19  &  n_n8743 ) ;
 assign wire4941 = ( n_n9401  &  nsr3_13  &  ndn3_12 ) | ( n_n9401  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4942 = ( ndn3_17  &  nsr3_20  &  n_n8811 ) ;
 assign wire4943 = ( ndn3_29  &  n_n8808  &  nsr3_35 ) ;
 assign wire4944 = ( n_n9126  &  nsr3_37  &  nen3_34 ) ;
 assign wire4945 = ( nsr3_30  &  n_n8809  &  ndn3_26 ) ;
 assign wire4946 = ( nsr3_38  &  nen3_36  &  n_n9390 ) ;
 assign wire4947 = ( nsr3_23  &  ndn3_19  &  n_n8810 ) ;
 assign wire4948 = ( n_n7824  &  nsr3_13  &  ndn3_12 ) | ( n_n7824  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4949 = ( ndn3_17  &  n_n8729  &  nsr3_20 ) ;
 assign wire4950 = ( ndn3_29  &  n_n7428  &  nsr3_35 ) ;
 assign wire4951 = ( n_n7598  &  nsr3_37  &  nen3_34 ) ;
 assign wire4952 = ( nsr3_30  &  ndn3_26  &  n_n7485 ) ;
 assign wire4953 = ( nsr3_38  &  nen3_36  &  n_n8898 ) ;
 assign wire4954 = ( nsr3_23  &  ndn3_19  &  n_n7429 ) ;
 assign wire4955 = ( nsr3_13  &  ndn3_12  &  n_n9496 ) | ( (~ nsr3_13)  &  nsr3_14  &  n_n9496 ) ;
 assign wire4956 = ( ndn3_17  &  n_n8884  &  nsr3_20 ) ;
 assign wire4957 = ( ndn3_29  &  nsr3_35  &  n_n8881 ) ;
 assign wire4958 = ( n_n9473  &  nsr3_37  &  nen3_34 ) ;
 assign wire4959 = ( n_n8882  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4960 = ( n_n9485  &  nsr3_38  &  nen3_36 ) ;
 assign wire4961 = ( n_n8883  &  nsr3_23  &  ndn3_19 ) ;
 assign wire4962 = ( n_n7877  &  nsr3_13  &  ndn3_12 ) | ( n_n7877  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4963 = ( ndn3_17  &  n_n8727  &  nsr3_20 ) ;
 assign wire4964 = ( n_n7452  &  ndn3_29  &  nsr3_35 ) ;
 assign wire4965 = ( n_n7640  &  nsr3_37  &  nen3_34 ) ;
 assign wire4966 = ( nsr3_30  &  ndn3_26  &  n_n7453 ) ;
 assign wire4967 = ( nsr3_38  &  nen3_36  &  n_n9458 ) ;
 assign wire4968 = ( nsr3_23  &  n_n7454  &  ndn3_19 ) ;
 assign wire4969 = ( nsr3_13  &  n_n9599  &  ndn3_12 ) | ( (~ nsr3_13)  &  n_n9599  &  nsr3_14 ) ;
 assign wire4970 = ( ndn3_17  &  n_n8939  &  nsr3_20 ) ;
 assign wire4971 = ( ndn3_29  &  nsr3_35  &  n_n8937 ) ;
 assign wire4972 = ( n_n9470  &  nsr3_37  &  nen3_34 ) ;
 assign wire4973 = ( nsr3_30  &  n_n8938  &  ndn3_26 ) ;
 assign wire4974 = ( n_n9588  &  nsr3_38  &  nen3_36 ) ;
 assign wire4975 = ( nsr3_23  &  ndn3_19  &  n_n9139 ) ;
 assign wire4976 = ( nsr3_13  &  n_n8984  &  ndn3_12 ) | ( (~ nsr3_13)  &  n_n8984  &  nsr3_14 ) ;
 assign wire4977 = ( ndn3_17  &  n_n8983  &  nsr3_20 ) ;
 assign wire4978 = ( n_n8981  &  ndn3_29  &  nsr3_35 ) ;
 assign wire4979 = ( n_n9334  &  nsr3_37  &  nen3_34 ) ;
 assign wire4980 = ( n_n8998  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4981 = ( nsr3_38  &  nen3_36  &  n_n8980 ) ;
 assign wire4982 = ( nsr3_23  &  ndn3_19  &  n_n8982 ) ;
 assign wire4983 = ( n_n8153  &  nsr3_13  &  ndn3_12 ) | ( n_n8153  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4984 = ( n_n8152  &  ndn3_17  &  nsr3_20 ) ;
 assign wire4985 = ( ndn3_29  &  nsr3_35  &  n_n8177 ) ;
 assign wire4986 = ( nsr3_37  &  n_n8628  &  nen3_34 ) ;
 assign wire4987 = ( n_n8545  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4988 = ( n_n9467  &  nsr3_38  &  nen3_36 ) ;
 assign wire4989 = ( nsr3_23  &  ndn3_19  &  n_n8151 ) ;
 assign wire4990 = ( n_n8282  &  nsr3_13  &  ndn3_12 ) | ( n_n8282  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire4991 = ( ndn3_17  &  n_n8281  &  nsr3_20 ) ;
 assign wire4992 = ( ndn3_29  &  n_n8278  &  nsr3_35 ) ;
 assign wire4993 = ( n_n8277  &  nsr3_37  &  nen3_34 ) ;
 assign wire4994 = ( n_n8279  &  nsr3_30  &  ndn3_26 ) ;
 assign wire4995 = ( nsr3_38  &  nen3_36  &  n_n8626 ) ;
 assign wire4996 = ( nsr3_23  &  ndn3_19  &  n_n8280 ) ;
 assign wire4997 = ( nsr3_13  &  ndn3_12  &  n_n8516 ) | ( (~ nsr3_13)  &  nsr3_14  &  n_n8516 ) ;
 assign wire4998 = ( ndn3_17  &  n_n8515  &  nsr3_20 ) ;
 assign wire4999 = ( ndn3_29  &  nsr3_35  &  n_n8513 ) ;
 assign wire5000 = ( n_n8512  &  nsr3_37  &  nen3_34 ) ;
 assign wire5001 = ( nsr3_30  &  n_n9203  &  ndn3_26 ) ;
 assign wire5002 = ( nsr3_38  &  nen3_36  &  n_n9108 ) ;
 assign wire5003 = ( nsr3_23  &  ndn3_19  &  n_n8514 ) ;
 assign wire5004 = ( (~ preset)  &  n_n6991  &  ngfdn_3 ) | ( (~ preset)  &  n_n6991  &  (~ ndn3_46) ) ;
 assign wire5005 = ( (~ preset)  &  (~ ngfdn_3)  &  n_n7896  &  ndn3_46 ) ;
 assign wire5006 = ( (~ preset)  &  n_n7271  &  ngfdn_3 ) | ( (~ preset)  &  n_n7271  &  (~ ndn3_46) ) ;
 assign wire5007 = ( (~ preset)  &  n_n8308  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign wire5008 = ( (~ preset)  &  n_n7252  &  ngfdn_3 ) | ( (~ preset)  &  n_n7252  &  (~ ndn3_46) ) ;
 assign wire5009 = ( (~ preset)  &  (~ ngfdn_3)  &  ndn3_46  &  n_n7444 ) ;
 assign wire5010 = ( (~ preset)  &  n_n8871  &  (~ nen3_39) ) | ( (~ preset)  &  n_n8871  &  ndn3_39 ) ;
 assign wire5012 = ( (~ preset)  &  n_n8592  &  ndn3_46 ) | ( (~ preset)  &  n_n8592  &  (~ ndn3_44) ) ;
 assign wire5013 = ( (~ preset)  &  n_n9259  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5022 = ( (~ preset)  &  n_n9401  &  (~ ndn3_11) ) | ( (~ preset)  &  n_n9401  &  ndn3_12 ) ;
 assign wire5026 = ( (~ preset)  &  n_n8150  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n8150  &  ndn3_40 ) ;
 assign wire5027 = ( wire2371  &  (~ n_n8314)  &  wire5069 ) | ( wire2371  &  (~ n_n8314)  &  wire5070 ) | ( wire2371  &  n_n8314  &  (~ wire5069)  &  (~ wire5070) ) ;
 assign wire5032 = ( n_n7813  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n7813 ) ;
 assign wire5033 = ( n_n7816  &  wire16048 ) | ( n_n7816  &  (~ ndn3_25)  &  ndn3_22 ) ;
 assign wire5037 = ( n_n7817  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5038 = ( nen3_39  &  n_n7807  &  (~ ndn3_39) ) ;
 assign wire5039 = ( (~ ndn3_9)  &  ndn3_7  &  n_n7815 ) ;
 assign wire5040 = ( (~ ngfdn_3)  &  n_n8222  &  ndn3_46 ) ;
 assign wire5041 = ( n_n7814  &  ndn3_9  &  (~ ndn3_11) ) ;
 assign wire5042 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7810 ) ;
 assign wire5043 = ( (~ ndn3_28)  &  n_n8473  &  nen3_28 ) ;
 assign wire5044 = ( n_n8022  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5045 = ( n_n7806  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5046 = ( (~ ndn3_34)  &  n_n7859  &  nen3_34 ) ;
 assign wire5047 = ( nen3_36  &  n_n7808  &  (~ ndn3_36) ) ;
 assign wire5048 = ( n_n8227  &  ndn3_17  &  (~ ndn3_18) ) ;
 assign wire5049 = ( nen3_22  &  (~ ndn3_22)  &  n_n8657 ) ;
 assign wire5050 = ( n_n7812  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5051 = ( n_n7793  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n7793 ) ;
 assign wire5052 = ( n_n7792  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n7792 ) ;
 assign wire5057 = ( (~ ndn3_7)  &  ndn3_4  &  n_n8267 ) ;
 assign wire5058 = ( n_n7791  &  ndn3_11  &  (~ ndn3_12) ) ;
 assign wire5059 = ( (~ ndn3_42)  &  ndn3_40  &  n_n7788 ) ;
 assign wire5060 = ( (~ ndn3_27)  &  n_n7809  &  ndn3_26 ) ;
 assign wire5061 = ( n_n9635  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign wire5062 = ( nen3_16  &  (~ ndn3_16)  &  n_n9525 ) ;
 assign wire5063 = ( ndn3_29  &  n_n7790  &  (~ ndn3_32) ) ;
 assign wire5064 = ( n_n7789  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5065 = ( ndn3_19  &  (~ ndn3_21)  &  n_n8402 ) ;
 assign wire5066 = ( (~ ndn3_25)  &  ndn3_22  &  n_n8841 ) ;
 assign wire5067 = ( n_n8223  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5068 = ( ndn3_17  &  n_n7811  &  (~ ndn3_18) ) ;
 assign wire5069 = ( wire16410  &  wire16427 ) | ( wire16411  &  wire16427 ) | ( wire16410  &  wire16428 ) | ( wire16411  &  wire16428 ) ;
 assign wire5070 = ( n_n8156  &  n_n8155  &  n_n7218 ) | ( n_n7566  &  (~ n_n8156)  &  n_n8155  &  n_n7218 ) | ( n_n7566  &  n_n8156  &  (~ n_n8155)  &  n_n7218 ) ;
 assign wire5071 = ( (~ preset)  &  psv2_5_5_  &  (~ ndn3_2)  &  nen3_2 ) ;
 assign wire5072 = ( (~ preset)  &  n_n9503  &  ndn3_2 ) | ( (~ preset)  &  n_n9503  &  (~ nen3_2) ) ;
 assign wire5077 = ( (~ preset)  &  n_n7779  &  ngfdn_3 ) | ( (~ preset)  &  n_n7779  &  (~ ndn3_46) ) ;
 assign wire5083 = ( n_n7764  &  wire16047 ) | ( nen3_16  &  n_n7764  &  (~ ndn3_16) ) ;
 assign wire5084 = ( n_n8506  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n8506 ) ;
 assign wire5088 = ( n_n9387  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5089 = ( nen3_39  &  (~ ndn3_39)  &  n_n7990 ) ;
 assign wire5090 = ( (~ ndn3_9)  &  ndn3_7  &  n_n7766 ) ;
 assign wire5091 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n9516 ) ;
 assign wire5092 = ( n_n7765  &  ndn3_9  &  (~ ndn3_11) ) ;
 assign wire5093 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7762 ) ;
 assign wire5094 = ( (~ ndn3_28)  &  nen3_28  &  n_n8852 ) ;
 assign wire5095 = ( n_n7757  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5096 = ( n_n7918  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5097 = ( n_n9157  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5098 = ( n_n7758  &  nen3_36  &  (~ ndn3_36) ) ;
 assign wire5099 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8203 ) ;
 assign wire5100 = ( nen3_22  &  (~ ndn3_22)  &  n_n7761 ) ;
 assign wire5101 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n8396 ) ;
 assign wire5102 = ( n_n7901  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n7901 ) ;
 assign wire5103 = ( n_n7713  &  wire16030 ) | ( (~ ndn3_17)  &  n_n7713  &  ndn3_16 ) ;
 assign wire5108 = ( n_n8086  &  (~ ndn3_7)  &  ndn3_4 ) ;
 assign wire5109 = ( ndn3_11  &  (~ ndn3_12)  &  n_n9210 ) ;
 assign wire5110 = ( n_n7707  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5111 = ( n_n7760  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5112 = ( (~ ngfdn_3)  &  n_n7706  &  ndn3_46 ) ;
 assign wire5113 = ( n_n8066  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5114 = ( ndn3_29  &  n_n7710  &  (~ ndn3_32) ) ;
 assign wire5115 = ( n_n7708  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5116 = ( n_n7712  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5117 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7711 ) ;
 assign wire5118 = ( n_n9110  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5119 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7763 ) ;
 assign wire5124 = ( n_n8760  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n8760 ) ;
 assign wire5125 = ( n_n7668  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n7668 ) ;
 assign wire5130 = ( n_n9300  &  (~ ndn3_7)  &  ndn3_4 ) ;
 assign wire5131 = ( ndn3_11  &  n_n8276  &  (~ ndn3_12) ) ;
 assign wire5132 = ( (~ ndn3_42)  &  ndn3_40  &  n_n9505 ) ;
 assign wire5133 = ( (~ ndn3_27)  &  n_n7684  &  ndn3_26 ) ;
 assign wire5134 = ( (~ ngfdn_3)  &  n_n7898  &  ndn3_46 ) ;
 assign wire5135 = ( nen3_16  &  (~ ndn3_16)  &  n_n8221 ) ;
 assign wire5136 = ( ndn3_29  &  n_n7666  &  (~ ndn3_32) ) ;
 assign wire5137 = ( ndn3_39  &  (~ ndn3_40)  &  n_n7664 ) ;
 assign wire5138 = ( n_n8597  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5139 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7667 ) ;
 assign wire5140 = ( (~ ndn3_46)  &  ndn3_44  &  n_n8628 ) ;
 assign wire5141 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7687 ) ;
 assign wire5142 = ( n_n7803  &  wire16047 ) | ( n_n7803  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5143 = ( n_n8116  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n8116 ) ;
 assign wire5147 = ( n_n7689  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5148 = ( nen3_39  &  (~ ndn3_39)  &  n_n7682 ) ;
 assign wire5149 = ( (~ ndn3_9)  &  ndn3_7  &  n_n9119 ) ;
 assign wire5150 = ( n_n9467  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign wire5151 = ( ndn3_9  &  (~ ndn3_11)  &  n_n7688 ) ;
 assign wire5152 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7686 ) ;
 assign wire5153 = ( (~ ndn3_28)  &  n_n7683  &  nen3_28 ) ;
 assign wire5154 = ( n_n8024  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5155 = ( n_n7681  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5156 = ( (~ ndn3_34)  &  n_n8889  &  nen3_34 ) ;
 assign wire5157 = ( nen3_36  &  (~ ndn3_36)  &  n_n7732 ) ;
 assign wire5158 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8153 ) ;
 assign wire5159 = ( nen3_22  &  (~ ndn3_22)  &  n_n7685 ) ;
 assign wire5160 = ( n_n9257  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5165 = ( n_n8786  &  wire16047 ) | ( n_n8786  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5166 = ( n_n8416  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n8416 ) ;
 assign wire5170 = ( n_n8739  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5171 = ( nen3_39  &  (~ ndn3_39)  &  n_n6968 ) ;
 assign wire5172 = ( (~ ndn3_9)  &  ndn3_7  &  n_n7866 ) ;
 assign wire5173 = ( (~ ngfdn_3)  &  n_n8980  &  ndn3_46 ) ;
 assign wire5174 = ( ndn3_9  &  (~ ndn3_11)  &  n_n7424 ) ;
 assign wire5175 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9342 ) ;
 assign wire5176 = ( (~ ndn3_28)  &  nen3_28  &  n_n9338 ) ;
 assign wire5177 = ( n_n8989  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5178 = ( ndn3_42  &  (~ ndn3_44)  &  n_n7920 ) ;
 assign wire5179 = ( (~ ndn3_34)  &  n_n9159  &  nen3_34 ) ;
 assign wire5180 = ( n_n7831  &  nen3_36  &  (~ ndn3_36) ) ;
 assign wire5181 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8984 ) ;
 assign wire5182 = ( nen3_22  &  (~ ndn3_22)  &  n_n7225 ) ;
 assign wire5183 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n8833 ) ;
 assign wire5184 = ( wire16377  &  wire16394 ) | ( wire16378  &  wire16394 ) | ( wire16377  &  wire16395 ) | ( wire16378  &  wire16395 ) ;
 assign wire5185 = ( n_n7997  &  n_n9258  &  n_n9587 ) | ( n_n7997  &  n_n8019  &  (~ n_n9258)  &  n_n9587 ) | ( n_n7997  &  n_n8019  &  n_n9258  &  (~ n_n9587) ) ;
 assign wire5188 = ( n_n8375  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n8375 ) ;
 assign wire5189 = ( n_n7956  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n7956 ) ;
 assign wire5193 = ( n_n9023  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5194 = ( nen3_39  &  n_n8095  &  (~ ndn3_39) ) ;
 assign wire5195 = ( (~ ndn3_9)  &  n_n7955  &  ndn3_7 ) ;
 assign wire5196 = ( (~ ngfdn_3)  &  n_n7947  &  ndn3_46 ) ;
 assign wire5197 = ( ndn3_9  &  n_n7954  &  (~ ndn3_11) ) ;
 assign wire5198 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9021 ) ;
 assign wire5199 = ( n_n9618  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire5200 = ( n_n7948  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5201 = ( ndn3_42  &  (~ ndn3_44)  &  n_n7949 ) ;
 assign wire5202 = ( n_n8891  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5203 = ( nen3_36  &  n_n7950  &  (~ ndn3_36) ) ;
 assign wire5204 = ( ndn3_17  &  n_n7951  &  (~ ndn3_18) ) ;
 assign wire5205 = ( nen3_22  &  (~ ndn3_22)  &  n_n8843 ) ;
 assign wire5206 = ( n_n7953  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5209 = ( n_n7696  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n7696 ) ;
 assign wire5210 = ( n_n7695  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n7695 ) ;
 assign wire5215 = ( (~ ndn3_7)  &  n_n9302  &  ndn3_4 ) ;
 assign wire5216 = ( ndn3_11  &  (~ ndn3_12)  &  n_n7694 ) ;
 assign wire5217 = ( (~ ndn3_42)  &  n_n8326  &  ndn3_40 ) ;
 assign wire5218 = ( (~ ndn3_27)  &  n_n8854  &  ndn3_26 ) ;
 assign wire5219 = ( (~ ngfdn_3)  &  n_n7691  &  ndn3_46 ) ;
 assign wire5220 = ( nen3_16  &  n_n8659  &  (~ ndn3_16) ) ;
 assign wire5221 = ( ndn3_29  &  n_n7693  &  (~ ndn3_32) ) ;
 assign wire5222 = ( n_n8410  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5223 = ( n_n8599  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5224 = ( (~ ndn3_25)  &  ndn3_22  &  n_n8697 ) ;
 assign wire5225 = ( n_n9518  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5226 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7952 ) ;
 assign wire5227 = ( n_n9347  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n9347 ) ;
 assign wire5228 = ( n_n9346  &  wire16030 ) | ( (~ ndn3_17)  &  n_n9346  &  ndn3_16 ) ;
 assign wire5233 = ( (~ ndn3_7)  &  ndn3_4  &  n_n9348 ) ;
 assign wire5234 = ( ndn3_11  &  (~ ndn3_12)  &  n_n9345 ) ;
 assign wire5235 = ( n_n9335  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5236 = ( n_n9339  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5237 = ( (~ ngfdn_3)  &  n_n9333  &  ndn3_46 ) ;
 assign wire5238 = ( nen3_16  &  (~ ndn3_16)  &  n_n9344 ) ;
 assign wire5239 = ( ndn3_29  &  n_n9337  &  (~ ndn3_32) ) ;
 assign wire5240 = ( ndn3_39  &  n_n9455  &  (~ ndn3_40) ) ;
 assign wire5241 = ( n_n9341  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5242 = ( (~ ndn3_25)  &  ndn3_22  &  n_n9340 ) ;
 assign wire5243 = ( n_n9334  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5244 = ( ndn3_17  &  n_n9343  &  (~ ndn3_18) ) ;
 assign wire5245 = ( (~ preset)  &  n_n9267  &  (~ ndn3_9) ) | ( (~ preset)  &  n_n9267  &  ndn3_11 ) ;
 assign wire5246 = ( (~ preset)  &  nrq3_11  &  (~ n_n8019)  &  n_n7573 ) | ( (~ preset)  &  nrq3_11  &  n_n8019  &  (~ n_n7573) ) ;
 assign wire5251 = ( n_n9602  &  wire16047 ) | ( n_n9602  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5252 = ( n_n9605  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n9605 ) ;
 assign wire5256 = ( (~ ndn3_4)  &  ndn3_2  &  n_n9606 ) ;
 assign wire5257 = ( nen3_39  &  (~ ndn3_39)  &  n_n9591 ) ;
 assign wire5258 = ( (~ ndn3_9)  &  ndn3_7  &  n_n9604 ) ;
 assign wire5259 = ( (~ ngfdn_3)  &  n_n9588  &  ndn3_46 ) ;
 assign wire5260 = ( ndn3_9  &  (~ ndn3_11)  &  n_n9603 ) ;
 assign wire5261 = ( n_n9598  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5262 = ( (~ ndn3_28)  &  n_n9595  &  nen3_28 ) ;
 assign wire5263 = ( n_n9589  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5264 = ( ndn3_42  &  (~ ndn3_44)  &  n_n9590 ) ;
 assign wire5265 = ( (~ ndn3_34)  &  n_n9593  &  nen3_34 ) ;
 assign wire5266 = ( nen3_36  &  n_n9592  &  (~ ndn3_36) ) ;
 assign wire5267 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9599 ) ;
 assign wire5268 = ( nen3_22  &  (~ ndn3_22)  &  n_n9597 ) ;
 assign wire5269 = ( n_n9601  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5270 = ( n_n9269  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n9269 ) ;
 assign wire5271 = ( n_n9268  &  wire16030 ) | ( (~ ndn3_17)  &  n_n9268  &  ndn3_16 ) ;
 assign wire5276 = ( (~ ndn3_7)  &  ndn3_4  &  n_n9270 ) ;
 assign wire5277 = ( n_n9267  &  ndn3_11  &  (~ ndn3_12) ) ;
 assign wire5278 = ( n_n9260  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5279 = ( n_n9596  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5280 = ( (~ ngfdn_3)  &  n_n9259  &  ndn3_46 ) ;
 assign wire5281 = ( nen3_16  &  (~ ndn3_16)  &  n_n9266 ) ;
 assign wire5282 = ( ndn3_29  &  n_n9263  &  (~ ndn3_32) ) ;
 assign wire5283 = ( ndn3_39  &  n_n9261  &  (~ ndn3_40) ) ;
 assign wire5284 = ( n_n9265  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5285 = ( (~ ndn3_25)  &  ndn3_22  &  n_n9264 ) ;
 assign wire5286 = ( n_n9470  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5287 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9600 ) ;
 assign wire5292 = ( n_n8377  &  wire16047 ) | ( n_n8377  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5293 = ( n_n9121  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n9121 ) ;
 assign wire5297 = ( (~ ndn3_4)  &  ndn3_2  &  n_n7881 ) ;
 assign wire5298 = ( nen3_39  &  (~ ndn3_39)  &  n_n7874 ) ;
 assign wire5299 = ( (~ ndn3_9)  &  ndn3_7  &  n_n7880 ) ;
 assign wire5300 = ( (~ ngfdn_3)  &  n_n9458  &  ndn3_46 ) ;
 assign wire5301 = ( ndn3_9  &  (~ ndn3_11)  &  n_n8051 ) ;
 assign wire5302 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7876 ) ;
 assign wire5303 = ( n_n9000  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire5304 = ( n_n8609  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5305 = ( n_n7873  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5306 = ( n_n9327  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5307 = ( nen3_36  &  n_n7980  &  (~ ndn3_36) ) ;
 assign wire5308 = ( n_n7877  &  ndn3_17  &  (~ ndn3_18) ) ;
 assign wire5309 = ( nen3_22  &  (~ ndn3_22)  &  n_n7875 ) ;
 assign wire5310 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n7879 ) ;
 assign wire5311 = ( n_n9583  &  n_n7818  &  n_n7597 ) | ( n_n9583  &  n_n8028  &  (~ n_n7818)  &  n_n7597 ) | ( n_n9583  &  n_n8028  &  n_n7818  &  (~ n_n7597) ) ;
 assign wire5312 = ( wire16081  &  wire16097 ) | ( wire16082  &  wire16097 ) | ( wire16081  &  wire16098 ) | ( wire16082  &  wire16098 ) ;
 assign wire5319 = ( n_n9404  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n9404 ) ;
 assign wire5320 = ( n_n9407  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n9407 ) ;
 assign wire5324 = ( n_n9408  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5325 = ( nen3_39  &  (~ ndn3_39)  &  n_n9393 ) ;
 assign wire5326 = ( (~ ndn3_9)  &  n_n9406  &  ndn3_7 ) ;
 assign wire5327 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n9390 ) ;
 assign wire5328 = ( ndn3_9  &  (~ ndn3_11)  &  n_n9405 ) ;
 assign wire5329 = ( n_n9400  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5330 = ( (~ ndn3_28)  &  n_n9397  &  nen3_28 ) ;
 assign wire5331 = ( n_n9391  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5332 = ( ndn3_42  &  (~ ndn3_44)  &  n_n9392 ) ;
 assign wire5333 = ( n_n9395  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5334 = ( nen3_36  &  n_n9394  &  (~ ndn3_36) ) ;
 assign wire5335 = ( n_n9401  &  ndn3_17  &  (~ ndn3_18) ) ;
 assign wire5336 = ( nen3_22  &  n_n9399  &  (~ ndn3_22) ) ;
 assign wire5337 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n9403 ) ;
 assign wire5338 = ( wire16179  &  wire16196 ) | ( wire16180  &  wire16196 ) | ( wire16179  &  wire16197 ) | ( wire16180  &  wire16197 ) ;
 assign wire5339 = ( n_n8953  &  n_n9040  &  n_n9307 ) | ( n_n9384  &  n_n8953  &  (~ n_n9040)  &  n_n9307 ) | ( n_n9384  &  n_n8953  &  n_n9040  &  (~ n_n9307) ) ;
 assign wire5342 = ( n_n7742  &  wire16047 ) | ( n_n7742  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5343 = ( n_n7837  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n7837 ) ;
 assign wire5347 = ( (~ ndn3_4)  &  n_n7744  &  ndn3_2 ) ;
 assign wire5348 = ( nen3_39  &  n_n7734  &  (~ ndn3_39) ) ;
 assign wire5349 = ( (~ ndn3_9)  &  n_n8053  &  ndn3_7 ) ;
 assign wire5350 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8135 ) ;
 assign wire5351 = ( ndn3_9  &  (~ ndn3_11)  &  n_n7743 ) ;
 assign wire5352 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7741 ) ;
 assign wire5353 = ( n_n7738  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire5354 = ( n_n8247  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5355 = ( n_n9059  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5356 = ( n_n7736  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5357 = ( n_n7735  &  nen3_36  &  (~ ndn3_36) ) ;
 assign wire5358 = ( n_n9141  &  ndn3_17  &  (~ ndn3_18) ) ;
 assign wire5359 = ( nen3_22  &  n_n7740  &  (~ ndn3_22) ) ;
 assign wire5360 = ( n_n9189  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5363 = ( n_n7655  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n7655 ) ;
 assign wire5364 = ( n_n7657  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n7657 ) ;
 assign wire5368 = ( (~ ndn3_4)  &  ndn3_2  &  n_n8770 ) ;
 assign wire5369 = ( nen3_39  &  n_n7650  &  (~ ndn3_39) ) ;
 assign wire5370 = ( (~ ndn3_9)  &  ndn3_7  &  n_n8619 ) ;
 assign wire5371 = ( (~ ngfdn_3)  &  n_n8862  &  ndn3_46 ) ;
 assign wire5372 = ( ndn3_9  &  n_n7656  &  (~ ndn3_11) ) ;
 assign wire5373 = ( n_n7654  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5374 = ( (~ ndn3_28)  &  n_n7652  &  nen3_28 ) ;
 assign wire5375 = ( (~ ndn3_46)  &  n_n8249  &  ndn3_44 ) ;
 assign wire5376 = ( ndn3_42  &  (~ ndn3_44)  &  n_n9061 ) ;
 assign wire5377 = ( (~ ndn3_34)  &  n_n9075  &  nen3_34 ) ;
 assign wire5378 = ( n_n7651  &  nen3_36  &  (~ ndn3_36) ) ;
 assign wire5379 = ( ndn3_17  &  n_n9015  &  (~ ndn3_18) ) ;
 assign wire5380 = ( nen3_22  &  (~ ndn3_22)  &  n_n7653 ) ;
 assign wire5381 = ( n_n8260  &  (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire5382 = ( n_n8641  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n8641 ) ;
 assign wire5383 = ( n_n9566  &  wire16030 ) | ( (~ ndn3_17)  &  n_n9566  &  ndn3_16 ) ;
 assign wire5388 = ( (~ ndn3_7)  &  ndn3_4  &  n_n7511 ) ;
 assign wire5389 = ( ndn3_11  &  (~ ndn3_12)  &  n_n8075 ) ;
 assign wire5390 = ( (~ ndn3_42)  &  n_n8477  &  ndn3_40 ) ;
 assign wire5391 = ( (~ ndn3_27)  &  n_n7728  &  ndn3_26 ) ;
 assign wire5392 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8670 ) ;
 assign wire5393 = ( nen3_16  &  n_n8210  &  (~ ndn3_16) ) ;
 assign wire5394 = ( ndn3_29  &  (~ ndn3_32)  &  n_n8526 ) ;
 assign wire5395 = ( n_n7995  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5396 = ( ndn3_19  &  (~ ndn3_21)  &  n_n7510 ) ;
 assign wire5397 = ( (~ ndn3_25)  &  ndn3_22  &  n_n9522 ) ;
 assign wire5398 = ( n_n7670  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5399 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7661 ) ;
 assign wire5402 = ( n_n9052  &  wire16029 ) | ( n_n9052  &  nen3_22  &  (~ ndn3_22) ) ;
 assign wire5403 = ( n_n9051  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n9051 ) ;
 assign wire5408 = ( (~ ndn3_7)  &  ndn3_4  &  n_n9053 ) ;
 assign wire5409 = ( ndn3_11  &  (~ ndn3_12)  &  n_n9050 ) ;
 assign wire5410 = ( n_n9043  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5411 = ( n_n9368  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5412 = ( (~ ngfdn_3)  &  n_n9041  &  ndn3_46 ) ;
 assign wire5413 = ( n_n9049  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5414 = ( ndn3_29  &  n_n9046  &  (~ ndn3_32) ) ;
 assign wire5415 = ( n_n9044  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5416 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9048 ) ;
 assign wire5417 = ( (~ ndn3_25)  &  ndn3_22  &  n_n9047 ) ;
 assign wire5418 = ( n_n9042  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5419 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9319 ) ;
 assign wire5420 = ( n_n9321  &  wire16047 ) | ( n_n9321  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5421 = ( n_n9324  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n9324 ) ;
 assign wire5425 = ( n_n9325  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5426 = ( n_n9311  &  nen3_39  &  (~ ndn3_39) ) ;
 assign wire5427 = ( (~ ndn3_9)  &  ndn3_7  &  n_n9323 ) ;
 assign wire5428 = ( (~ ngfdn_3)  &  n_n9308  &  ndn3_46 ) ;
 assign wire5429 = ( ndn3_9  &  (~ ndn3_11)  &  n_n9322 ) ;
 assign wire5430 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9317 ) ;
 assign wire5431 = ( (~ ndn3_28)  &  n_n9315  &  nen3_28 ) ;
 assign wire5432 = ( n_n9309  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5433 = ( n_n9310  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5434 = ( (~ ndn3_34)  &  n_n9313  &  nen3_34 ) ;
 assign wire5435 = ( nen3_36  &  n_n9312  &  (~ ndn3_36) ) ;
 assign wire5436 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9318 ) ;
 assign wire5437 = ( nen3_22  &  (~ ndn3_22)  &  n_n9316 ) ;
 assign wire5438 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n9320 ) ;
 assign wire5439 = ( n_n7553  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n7553 ) ;
 assign wire5440 = ( n_n9563  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n9563 ) ;
 assign wire5445 = ( (~ ndn3_7)  &  ndn3_4  &  n_n7554 ) ;
 assign wire5446 = ( n_n8298  &  ndn3_11  &  (~ ndn3_12) ) ;
 assign wire5447 = ( (~ ndn3_42)  &  n_n8636  &  ndn3_40 ) ;
 assign wire5448 = ( (~ ndn3_27)  &  n_n7739  &  ndn3_26 ) ;
 assign wire5449 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n9239 ) ;
 assign wire5450 = ( nen3_16  &  n_n8381  &  (~ ndn3_16) ) ;
 assign wire5451 = ( n_n7552  &  ndn3_29  &  (~ ndn3_32) ) ;
 assign wire5452 = ( ndn3_39  &  n_n7993  &  (~ ndn3_40) ) ;
 assign wire5453 = ( n_n8035  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5454 = ( n_n8533  &  (~ ndn3_25)  &  ndn3_22 ) ;
 assign wire5455 = ( n_n8499  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5456 = ( ndn3_17  &  n_n9528  &  (~ ndn3_18) ) ;
 assign wire5457 = ( n_n9135  &  wire16029 ) | ( nen3_22  &  n_n9135  &  (~ ndn3_22) ) ;
 assign wire5458 = ( n_n9134  &  wire16030 ) | ( (~ ndn3_17)  &  n_n9134  &  ndn3_16 ) ;
 assign wire5463 = ( (~ ndn3_7)  &  ndn3_4  &  n_n9136 ) ;
 assign wire5464 = ( ndn3_11  &  (~ ndn3_12)  &  n_n9133 ) ;
 assign wire5465 = ( n_n9127  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5466 = ( n_n9398  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5467 = ( (~ ngfdn_3)  &  n_n9125  &  ndn3_46 ) ;
 assign wire5468 = ( nen3_16  &  n_n9132  &  (~ ndn3_16) ) ;
 assign wire5469 = ( ndn3_29  &  n_n9129  &  (~ ndn3_32) ) ;
 assign wire5470 = ( ndn3_39  &  n_n9128  &  (~ ndn3_40) ) ;
 assign wire5471 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9131 ) ;
 assign wire5472 = ( n_n9130  &  (~ ndn3_25)  &  ndn3_22 ) ;
 assign wire5473 = ( (~ ndn3_46)  &  n_n9126  &  ndn3_44 ) ;
 assign wire5474 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9402 ) ;
 assign wire5477 = ( n_n8791  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n8791 ) ;
 assign wire5478 = ( n_n9008  &  wire16030 ) | ( n_n9008  &  (~ ndn3_17)  &  ndn3_16 ) ;
 assign wire5483 = ( (~ ndn3_7)  &  ndn3_4  &  n_n7604 ) ;
 assign wire5484 = ( ndn3_11  &  (~ ndn3_12)  &  n_n8296 ) ;
 assign wire5485 = ( n_n7599  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5486 = ( n_n7822  &  (~ ndn3_27)  &  ndn3_26 ) ;
 assign wire5487 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n9237 ) ;
 assign wire5488 = ( nen3_16  &  n_n8042  &  (~ ndn3_16) ) ;
 assign wire5489 = ( ndn3_29  &  (~ ndn3_32)  &  n_n7601 ) ;
 assign wire5490 = ( ndn3_39  &  n_n8253  &  (~ ndn3_40) ) ;
 assign wire5491 = ( ndn3_19  &  n_n7603  &  (~ ndn3_21) ) ;
 assign wire5492 = ( (~ ndn3_25)  &  n_n7602  &  ndn3_22 ) ;
 assign wire5493 = ( n_n7598  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5494 = ( ndn3_17  &  (~ ndn3_18)  &  n_n8233 ) ;
 assign wire5495 = ( n_n7825  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n7825 ) ;
 assign wire5496 = ( n_n7835  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n7835 ) ;
 assign wire5500 = ( (~ ndn3_4)  &  n_n7827  &  ndn3_2 ) ;
 assign wire5501 = ( n_n7819  &  nen3_39  &  (~ ndn3_39) ) ;
 assign wire5502 = ( (~ ndn3_9)  &  n_n7826  &  ndn3_7 ) ;
 assign wire5503 = ( (~ ngfdn_3)  &  n_n8898  &  ndn3_46 ) ;
 assign wire5504 = ( ndn3_9  &  (~ ndn3_11)  &  n_n8617 ) ;
 assign wire5505 = ( n_n7823  &  ndn3_19  &  (~ ndn3_21) ) ;
 assign wire5506 = ( n_n7821  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire5507 = ( n_n9036  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5508 = ( ndn3_42  &  (~ ndn3_44)  &  n_n9081 ) ;
 assign wire5509 = ( n_n7820  &  (~ ndn3_34)  &  nen3_34 ) ;
 assign wire5510 = ( nen3_36  &  n_n7925  &  (~ ndn3_36) ) ;
 assign wire5511 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7824 ) ;
 assign wire5512 = ( n_n8699  &  nen3_22  &  (~ ndn3_22) ) ;
 assign wire5513 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n9186 ) ;
 assign wire5516 = ( n_n9499  &  wire16047 ) | ( nen3_16  &  (~ ndn3_16)  &  n_n9499 ) ;
 assign wire5517 = ( n_n9502  &  wire16048 ) | ( (~ ndn3_25)  &  ndn3_22  &  n_n9502 ) ;
 assign wire5521 = ( n_n9503  &  (~ ndn3_4)  &  ndn3_2 ) ;
 assign wire5522 = ( nen3_39  &  (~ ndn3_39)  &  n_n9488 ) ;
 assign wire5523 = ( (~ ndn3_9)  &  n_n9501  &  ndn3_7 ) ;
 assign wire5524 = ( n_n9485  &  (~ ngfdn_3)  &  ndn3_46 ) ;
 assign wire5525 = ( ndn3_9  &  (~ ndn3_11)  &  n_n9500 ) ;
 assign wire5526 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9495 ) ;
 assign wire5527 = ( n_n9492  &  (~ ndn3_28)  &  nen3_28 ) ;
 assign wire5528 = ( n_n9486  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5529 = ( n_n9487  &  ndn3_42  &  (~ ndn3_44) ) ;
 assign wire5530 = ( (~ ndn3_34)  &  n_n9490  &  nen3_34 ) ;
 assign wire5531 = ( n_n9489  &  nen3_36  &  (~ ndn3_36) ) ;
 assign wire5532 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9496 ) ;
 assign wire5533 = ( nen3_22  &  (~ ndn3_22)  &  n_n9494 ) ;
 assign wire5534 = ( (~ nsr3_13)  &  (~ ndn3_15)  &  n_n9498 ) ;
 assign wire5535 = ( n_n9181  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n9181 ) ;
 assign wire5536 = ( n_n9180  &  wire16030 ) | ( n_n9180  &  (~ ndn3_17)  &  ndn3_16 ) ;
 assign wire5541 = ( (~ ndn3_7)  &  n_n9182  &  ndn3_4 ) ;
 assign wire5542 = ( ndn3_11  &  (~ ndn3_12)  &  n_n9179 ) ;
 assign wire5543 = ( n_n9172  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5544 = ( (~ ndn3_27)  &  n_n9493  &  ndn3_26 ) ;
 assign wire5545 = ( (~ ngfdn_3)  &  n_n9171  &  ndn3_46 ) ;
 assign wire5546 = ( nen3_16  &  (~ ndn3_16)  &  n_n9178 ) ;
 assign wire5547 = ( ndn3_29  &  n_n9175  &  (~ ndn3_32) ) ;
 assign wire5548 = ( ndn3_39  &  n_n9173  &  (~ ndn3_40) ) ;
 assign wire5549 = ( ndn3_19  &  (~ ndn3_21)  &  n_n9177 ) ;
 assign wire5550 = ( (~ ndn3_25)  &  ndn3_22  &  n_n9176 ) ;
 assign wire5551 = ( n_n9473  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5552 = ( ndn3_17  &  (~ ndn3_18)  &  n_n9497 ) ;
 assign wire5553 = ( n_n8789  &  wire16029 ) | ( nen3_22  &  (~ ndn3_22)  &  n_n8789 ) ;
 assign wire5554 = ( n_n8961  &  wire16030 ) | ( (~ ndn3_17)  &  ndn3_16  &  n_n8961 ) ;
 assign wire5559 = ( n_n7643  &  (~ ndn3_7)  &  ndn3_4 ) ;
 assign wire5560 = ( ndn3_11  &  (~ ndn3_12)  &  n_n7642 ) ;
 assign wire5561 = ( n_n8328  &  (~ ndn3_42)  &  ndn3_40 ) ;
 assign wire5562 = ( (~ ndn3_27)  &  n_n8856  &  ndn3_26 ) ;
 assign wire5563 = ( (~ ngfdn_3)  &  ndn3_46  &  n_n8188 ) ;
 assign wire5564 = ( n_n8661  &  nen3_16  &  (~ ndn3_16) ) ;
 assign wire5565 = ( ndn3_29  &  n_n7649  &  (~ ndn3_32) ) ;
 assign wire5566 = ( n_n8552  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5567 = ( ndn3_19  &  (~ ndn3_21)  &  n_n8058 ) ;
 assign wire5568 = ( (~ ndn3_25)  &  ndn3_22  &  n_n7641 ) ;
 assign wire5569 = ( n_n7640  &  (~ ndn3_46)  &  ndn3_44 ) ;
 assign wire5570 = ( ndn3_17  &  (~ ndn3_18)  &  n_n7878 ) ;
 assign wire5571 = ( (~ preset)  &  n_n7726  &  (~ ndn3_39) ) | ( (~ preset)  &  n_n7726  &  ndn3_40 ) ;
 assign wire5572 = ( (~ preset)  &  n_n7376  &  ndn3_39  &  (~ ndn3_40) ) ;
 assign wire5573 = ( (~ preset)  &  n_n9260  &  ndn3_37 ) | ( (~ preset)  &  n_n9260  &  nsr3_37 ) ;
 assign wire5575 = ( (~ preset)  &  n_n9172  &  ndn3_37 ) | ( (~ preset)  &  n_n9172  &  nsr3_37 ) ;
 assign wire5579 = ( (~ nsr3_13)  &  n_n8649  &  nsr3_14 ) ;
 assign wire5580 = ( ndn3_17  &  n_n8648  &  nsr3_20 ) ;
 assign wire5581 = ( nsr3_13  &  ndn3_12  &  n_n8650 ) ;
 assign wire5582 = ( ndn3_29  &  nsr3_35  &  n_n8796 ) ;
 assign wire5583 = ( n_n8647  &  nsr3_37  &  nen3_34 ) ;
 assign wire5584 = ( n_n9242  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5585 = ( nsr3_38  &  nen3_36  &  n_n8646 ) ;
 assign wire5586 = ( nsr3_23  &  ndn3_19  &  n_n9013 ) ;
 assign wire5587 = ( (~ nsr3_13)  &  nsr3_14  &  n_n7629 ) ;
 assign wire5588 = ( ndn3_17  &  nsr3_20  &  n_n7628 ) ;
 assign wire5589 = ( nsr3_13  &  ndn3_12  &  n_n7630 ) ;
 assign wire5590 = ( n_n8613  &  ndn3_29  &  nsr3_35 ) ;
 assign wire5591 = ( n_n8875  &  nsr3_37  &  nen3_34 ) ;
 assign wire5592 = ( nsr3_30  &  n_n8141  &  ndn3_26 ) ;
 assign wire5593 = ( nsr3_38  &  nen3_36  &  n_n7627 ) ;
 assign wire5594 = ( nsr3_23  &  n_n7983  &  ndn3_19 ) ;
 assign wire5595 = ( (~ nsr3_13)  &  nsr3_14  &  n_n9165 ) ;
 assign wire5596 = ( ndn3_17  &  n_n9164  &  nsr3_20 ) ;
 assign wire5597 = ( nsr3_13  &  ndn3_12  &  n_n9166 ) ;
 assign wire5598 = ( ndn3_29  &  nsr3_35  &  n_n9161 ) ;
 assign wire5599 = ( n_n9160  &  nsr3_37  &  nen3_34 ) ;
 assign wire5600 = ( nsr3_30  &  n_n9162  &  ndn3_26 ) ;
 assign wire5601 = ( nsr3_38  &  nen3_36  &  n_n9578 ) ;
 assign wire5602 = ( nsr3_23  &  ndn3_19  &  n_n9163 ) ;
 assign wire5603 = ( (~ nsr3_13)  &  n_n8240  &  nsr3_14 ) ;
 assign wire5604 = ( ndn3_17  &  n_n8239  &  nsr3_20 ) ;
 assign wire5605 = ( nsr3_13  &  ndn3_12  &  n_n8241 ) ;
 assign wire5606 = ( ndn3_29  &  nsr3_35  &  n_n8312 ) ;
 assign wire5607 = ( n_n8236  &  nsr3_37  &  nen3_34 ) ;
 assign wire5608 = ( n_n8237  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5609 = ( nsr3_38  &  n_n8235  &  nen3_36 ) ;
 assign wire5610 = ( nsr3_23  &  ndn3_19  &  n_n8238 ) ;
 assign wire5611 = ( (~ nsr3_13)  &  nsr3_14  &  n_n8574 ) ;
 assign wire5612 = ( n_n8573  &  ndn3_17  &  nsr3_20 ) ;
 assign wire5613 = ( nsr3_13  &  ndn3_12  &  n_n8575 ) ;
 assign wire5614 = ( ndn3_29  &  n_n8572  &  nsr3_35 ) ;
 assign wire5615 = ( n_n8571  &  nsr3_37  &  nen3_34 ) ;
 assign wire5616 = ( nsr3_30  &  n_n8970  &  ndn3_26 ) ;
 assign wire5617 = ( nsr3_38  &  nen3_36  &  n_n8570 ) ;
 assign wire5618 = ( n_n9150  &  nsr3_23  &  ndn3_19 ) ;
 assign wire5619 = ( n_n9362  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire5620 = ( ndn3_17  &  n_n9552  &  nsr3_20 ) ;
 assign wire5621 = ( nsr3_13  &  ndn3_12  &  n_n9363 ) ;
 assign wire5622 = ( ndn3_29  &  nsr3_35  &  n_n9359 ) ;
 assign wire5623 = ( n_n9358  &  nsr3_37  &  nen3_34 ) ;
 assign wire5624 = ( nsr3_30  &  n_n9360  &  ndn3_26 ) ;
 assign wire5625 = ( nsr3_38  &  nen3_36  &  n_n9357 ) ;
 assign wire5626 = ( n_n9361  &  nsr3_23  &  ndn3_19 ) ;
 assign wire5627 = ( (~ nsr3_13)  &  nsr3_14  &  n_n9292 ) ;
 assign wire5628 = ( ndn3_17  &  n_n9291  &  nsr3_20 ) ;
 assign wire5629 = ( n_n9410  &  nsr3_13  &  ndn3_12 ) ;
 assign wire5630 = ( ndn3_29  &  nsr3_35  &  n_n9289 ) ;
 assign wire5631 = ( n_n9539  &  nsr3_37  &  nen3_34 ) ;
 assign wire5632 = ( n_n9290  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5633 = ( nsr3_38  &  nen3_36  &  n_n9296 ) ;
 assign wire5634 = ( nsr3_23  &  ndn3_19  &  n_n9298 ) ;
 assign wire5635 = ( (~ nsr3_13)  &  n_n8273  &  nsr3_14 ) ;
 assign wire5636 = ( ndn3_17  &  n_n8272  &  nsr3_20 ) ;
 assign wire5637 = ( nsr3_13  &  n_n8274  &  ndn3_12 ) ;
 assign wire5638 = ( ndn3_29  &  n_n8348  &  nsr3_35 ) ;
 assign wire5639 = ( n_n8269  &  nsr3_37  &  nen3_34 ) ;
 assign wire5640 = ( n_n8270  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5641 = ( n_n8508  &  nsr3_38  &  nen3_36 ) ;
 assign wire5642 = ( nsr3_23  &  ndn3_19  &  n_n8271 ) ;
 assign wire5643 = ( n_n9560  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire5644 = ( ndn3_17  &  n_n9559  &  nsr3_20 ) ;
 assign wire5645 = ( n_n9561  &  nsr3_13  &  ndn3_12 ) ;
 assign wire5646 = ( ndn3_29  &  nsr3_35  &  n_n9556 ) ;
 assign wire5647 = ( n_n9555  &  nsr3_37  &  nen3_34 ) ;
 assign wire5648 = ( n_n9557  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5649 = ( n_n9554  &  nsr3_38  &  nen3_36 ) ;
 assign wire5650 = ( nsr3_23  &  ndn3_19  &  n_n9558 ) ;
 assign wire5651 = ( (~ nsr3_13)  &  n_n9510  &  nsr3_14 ) ;
 assign wire5652 = ( ndn3_17  &  n_n7854  &  nsr3_20 ) ;
 assign wire5653 = ( n_n8037  &  nsr3_13  &  ndn3_12 ) ;
 assign wire5654 = ( ndn3_29  &  nsr3_35  &  n_n7852 ) ;
 assign wire5655 = ( nsr3_37  &  n_n8756  &  nen3_34 ) ;
 assign wire5656 = ( nsr3_30  &  n_n8972  &  ndn3_26 ) ;
 assign wire5657 = ( nsr3_38  &  nen3_36  &  n_n8171 ) ;
 assign wire5658 = ( nsr3_23  &  ndn3_19  &  n_n7853 ) ;
 assign wire5659 = ( (~ nsr3_13)  &  n_n7771  &  nsr3_14 ) ;
 assign wire5660 = ( ndn3_17  &  nsr3_20  &  n_n7770 ) ;
 assign wire5661 = ( nsr3_13  &  ndn3_12  &  n_n7961 ) ;
 assign wire5662 = ( ndn3_29  &  n_n9331  &  nsr3_35 ) ;
 assign wire5663 = ( n_n7768  &  nsr3_37  &  nen3_34 ) ;
 assign wire5664 = ( nsr3_30  &  n_n7769  &  ndn3_26 ) ;
 assign wire5665 = ( n_n8173  &  nsr3_38  &  nen3_36 ) ;
 assign wire5666 = ( nsr3_23  &  ndn3_19  &  n_n8803 ) ;
 assign wire5667 = ( n_n8199  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire5668 = ( n_n9280  &  ndn3_17  &  nsr3_20 ) ;
 assign wire5669 = ( nsr3_13  &  ndn3_12  &  n_n8200 ) ;
 assign wire5670 = ( ndn3_29  &  nsr3_35  &  n_n8197 ) ;
 assign wire5671 = ( n_n8710  &  nsr3_37  &  nen3_34 ) ;
 assign wire5672 = ( nsr3_30  &  n_n8366  &  ndn3_26 ) ;
 assign wire5673 = ( n_n8196  &  nsr3_38  &  nen3_36 ) ;
 assign wire5674 = ( nsr3_23  &  ndn3_19  &  n_n8198 ) ;
 assign wire5675 = ( (~ nsr3_13)  &  nsr3_14  &  n_n9441 ) ;
 assign wire5676 = ( ndn3_17  &  n_n9550  &  nsr3_20 ) ;
 assign wire5677 = ( n_n9442  &  nsr3_13  &  ndn3_12 ) ;
 assign wire5678 = ( ndn3_29  &  n_n9438  &  nsr3_35 ) ;
 assign wire5679 = ( n_n9437  &  nsr3_37  &  nen3_34 ) ;
 assign wire5680 = ( nsr3_30  &  n_n9439  &  ndn3_26 ) ;
 assign wire5681 = ( nsr3_38  &  nen3_36  &  n_n9436 ) ;
 assign wire5682 = ( nsr3_23  &  ndn3_19  &  n_n9440 ) ;
 assign wire5683 = ( (~ nsr3_13)  &  n_n7584  &  nsr3_14 ) ;
 assign wire5684 = ( ndn3_17  &  nsr3_20  &  n_n8447 ) ;
 assign wire5685 = ( nsr3_13  &  ndn3_12  &  n_n8691 ) ;
 assign wire5686 = ( ndn3_29  &  n_n8968  &  nsr3_35 ) ;
 assign wire5687 = ( n_n7582  &  nsr3_37  &  nen3_34 ) ;
 assign wire5688 = ( n_n7583  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5689 = ( nsr3_38  &  nen3_36  &  n_n8016 ) ;
 assign wire5690 = ( nsr3_23  &  ndn3_19  &  n_n7985 ) ;
 assign wire5691 = ( (~ nsr3_13)  &  nsr3_14  &  n_n7704 ) ;
 assign wire5692 = ( ndn3_17  &  n_n8685  &  nsr3_20 ) ;
 assign wire5693 = ( nsr3_13  &  ndn3_12  &  n_n8577 ) ;
 assign wire5694 = ( ndn3_29  &  nsr3_35  &  n_n9294 ) ;
 assign wire5695 = ( nsr3_37  &  n_n8118  &  nen3_34 ) ;
 assign wire5696 = ( n_n7702  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5697 = ( nsr3_38  &  nen3_36  &  n_n7701 ) ;
 assign wire5698 = ( nsr3_23  &  n_n7703  &  ndn3_19 ) ;
 assign wire5699 = ( n_n8531  &  (~ nsr3_13)  &  nsr3_14 ) ;
 assign wire5700 = ( ndn3_17  &  n_n8530  &  nsr3_20 ) ;
 assign wire5701 = ( nsr3_13  &  n_n8615  &  ndn3_12 ) ;
 assign wire5702 = ( ndn3_29  &  nsr3_35  &  n_n9275 ) ;
 assign wire5703 = ( n_n8529  &  nsr3_37  &  nen3_34 ) ;
 assign wire5704 = ( n_n9244  &  nsr3_30  &  ndn3_26 ) ;
 assign wire5705 = ( nsr3_38  &  nen3_36  &  n_n8528 ) ;
 assign wire5706 = ( nsr3_23  &  n_n8935  &  ndn3_19 ) ;
 assign wire15923 = ( wire5699 ) | ( wire5700 ) | ( wire5701 ) | ( wire5702 ) ;
 assign wire15924 = ( wire5703 ) | ( wire5704 ) | ( wire5705 ) | ( wire5706 ) ;
 assign wire15929 = ( wire5603 ) | ( wire5604 ) | ( wire5605 ) | ( wire5606 ) ;
 assign wire15930 = ( wire5607 ) | ( wire5608 ) | ( wire5609 ) | ( wire5610 ) ;
 assign wire15935 = ( wire5611 ) | ( wire5612 ) | ( wire5613 ) | ( wire5614 ) ;
 assign wire15936 = ( wire5615 ) | ( wire5616 ) | ( wire5617 ) | ( wire5618 ) ;
 assign wire15941 = ( wire5619 ) | ( wire5620 ) | ( wire5621 ) | ( wire5622 ) ;
 assign wire15942 = ( wire5623 ) | ( wire5624 ) | ( wire5625 ) | ( wire5626 ) ;
 assign wire15947 = ( wire5683 ) | ( wire5684 ) | ( wire5685 ) | ( wire5686 ) ;
 assign wire15948 = ( wire5687 ) | ( wire5688 ) | ( wire5689 ) | ( wire5690 ) ;
 assign wire15953 = ( wire5691 ) | ( wire5692 ) | ( wire5693 ) | ( wire5694 ) ;
 assign wire15954 = ( wire5695 ) | ( wire5696 ) | ( wire5697 ) | ( wire5698 ) ;
 assign wire15959 = ( wire5587 ) | ( wire5588 ) | ( wire5589 ) | ( wire5590 ) ;
 assign wire15960 = ( wire5591 ) | ( wire5592 ) | ( wire5593 ) | ( wire5594 ) ;
 assign wire15965 = ( wire5659 ) | ( wire5660 ) | ( wire5661 ) | ( wire5662 ) ;
 assign wire15966 = ( wire5663 ) | ( wire5664 ) | ( wire5665 ) | ( wire5666 ) ;
 assign wire15971 = ( wire5643 ) | ( wire5644 ) | ( wire5645 ) | ( wire5646 ) ;
 assign wire15972 = ( wire5647 ) | ( wire5648 ) | ( wire5649 ) | ( wire5650 ) ;
 assign wire15977 = ( wire5595 ) | ( wire5596 ) | ( wire5597 ) | ( wire5598 ) ;
 assign wire15978 = ( wire5599 ) | ( wire5600 ) | ( wire5601 ) | ( wire5602 ) ;
 assign wire15983 = ( wire5579 ) | ( wire5580 ) | ( wire5581 ) | ( wire5582 ) ;
 assign wire15984 = ( wire5583 ) | ( wire5584 ) | ( wire5585 ) | ( wire5586 ) ;
 assign wire15989 = ( wire5651 ) | ( wire5652 ) | ( wire5653 ) | ( wire5654 ) ;
 assign wire15990 = ( wire5655 ) | ( wire5656 ) | ( wire5657 ) | ( wire5658 ) ;
 assign wire15995 = ( wire5627 ) | ( wire5628 ) | ( wire5629 ) | ( wire5630 ) ;
 assign wire15996 = ( wire5631 ) | ( wire5632 ) | ( wire5633 ) | ( wire5634 ) ;
 assign wire16001 = ( wire5675 ) | ( wire5676 ) | ( wire5677 ) | ( wire5678 ) ;
 assign wire16002 = ( wire5679 ) | ( wire5680 ) | ( wire5681 ) | ( wire5682 ) ;
 assign wire16007 = ( wire5635 ) | ( wire5636 ) | ( wire5637 ) | ( wire5638 ) ;
 assign wire16008 = ( wire5639 ) | ( wire5640 ) | ( wire5641 ) | ( wire5642 ) ;
 assign wire16013 = ( wire5667 ) | ( wire5668 ) | ( wire5669 ) | ( wire5670 ) ;
 assign wire16014 = ( wire5671 ) | ( wire5672 ) | ( wire5673 ) | ( wire5674 ) ;
 assign wire16015 = ( wire15923 ) | ( wire15924 ) | ( wire15929 ) | ( wire15930 ) ;
 assign wire16016 = ( wire15935 ) | ( wire15936 ) | ( wire15941 ) | ( wire15942 ) ;
 assign wire16017 = ( wire15947 ) | ( wire15948 ) | ( wire15953 ) | ( wire15954 ) ;
 assign wire16018 = ( wire15959 ) | ( wire15960 ) | ( wire15965 ) | ( wire15966 ) ;
 assign wire16019 = ( wire15971 ) | ( wire15972 ) | ( wire15977 ) | ( wire15978 ) ;
 assign wire16020 = ( wire15983 ) | ( wire15984 ) | ( wire15989 ) | ( wire15990 ) ;
 assign wire16021 = ( wire15995 ) | ( wire15996 ) | ( wire16001 ) | ( wire16002 ) ;
 assign wire16022 = ( wire16007 ) | ( wire16008 ) | ( wire16013 ) | ( wire16014 ) ;
 assign wire16027 = ( wire16015 ) | ( wire16016 ) | ( wire16017 ) | ( wire16018 ) ;
 assign wire16028 = ( wire16019 ) | ( wire16020 ) | ( wire16021 ) | ( wire16022 ) ;
 assign wire16029 = ( (~ ndn3_9)  &  ndn3_7 ) | ( ndn3_25  &  (~ ndn3_26) ) ;
 assign wire16030 = ( ndn3_9  &  (~ ndn3_11) ) | ( (~ nsr3_13)  &  (~ ndn3_15) ) ;
 assign wire16037 = ( n_n8779  &  wire2375 ) | ( n_n7876  &  wire2377 ) ;
 assign wire16038 = ( n_n7644  &  wire2373 ) | ( n_n9000  &  wire2374 ) ;
 assign wire16039 = ( wire5559 ) | ( wire5560 ) | ( wire5561 ) | ( wire5562 ) ;
 assign wire16040 = ( wire5563 ) | ( wire5564 ) | ( wire5565 ) | ( wire5566 ) ;
 assign wire16041 = ( wire5567 ) | ( wire5568 ) | ( wire5569 ) | ( wire5570 ) ;
 assign wire16045 = ( wire5553 ) | ( wire5554 ) | ( wire16041 ) ;
 assign wire16046 = ( wire16037 ) | ( wire16038 ) | ( wire16039 ) | ( wire16040 ) ;
 assign wire16047 = ( (~ ndn3_19)  &  nen3_19 ) | ( ndn3_11  &  (~ ndn3_12) ) ;
 assign wire16048 = ( (~ ndn3_29)  &  ndn3_28 ) | ( (~ ndn3_7)  &  ndn3_4 ) ;
 assign wire16056 = ( n_n9230  &  wire2381 ) | ( n_n7878  &  wire2383 ) ;
 assign wire16057 = ( wire5297 ) | ( wire5298 ) | ( n_n8856  &  wire2380 ) ;
 assign wire16058 = ( wire5299 ) | ( wire5300 ) | ( wire5301 ) | ( wire5302 ) ;
 assign wire16059 = ( wire5303 ) | ( wire5304 ) | ( wire5305 ) | ( wire5306 ) ;
 assign wire16060 = ( wire5307 ) | ( wire5308 ) | ( wire5309 ) | ( wire5310 ) ;
 assign wire16064 = ( wire5292 ) | ( wire5293 ) | ( wire16060 ) ;
 assign wire16065 = ( wire16056 ) | ( wire16057 ) | ( wire16058 ) | ( wire16059 ) ;
 assign wire16073 = ( n_n9491  &  wire2381 ) | ( n_n9497  &  wire2383 ) ;
 assign wire16074 = ( wire5521 ) | ( wire5522 ) | ( n_n9493  &  wire2380 ) ;
 assign wire16075 = ( wire5523 ) | ( wire5524 ) | ( wire5525 ) | ( wire5526 ) ;
 assign wire16076 = ( wire5527 ) | ( wire5528 ) | ( wire5529 ) | ( wire5530 ) ;
 assign wire16077 = ( wire5531 ) | ( wire5532 ) | ( wire5533 ) | ( wire5534 ) ;
 assign wire16081 = ( wire5516 ) | ( wire5517 ) | ( wire16077 ) ;
 assign wire16082 = ( wire16073 ) | ( wire16074 ) | ( wire16075 ) | ( wire16076 ) ;
 assign wire16089 = ( n_n9174  &  wire2375 ) | ( n_n9495  &  wire2377 ) ;
 assign wire16090 = ( n_n9183  &  wire2373 ) | ( n_n9492  &  wire2374 ) ;
 assign wire16091 = ( wire5541 ) | ( wire5542 ) | ( wire5543 ) | ( wire5544 ) ;
 assign wire16092 = ( wire5545 ) | ( wire5546 ) | ( wire5547 ) | ( wire5548 ) ;
 assign wire16093 = ( wire5549 ) | ( wire5550 ) | ( wire5551 ) | ( wire5552 ) ;
 assign wire16097 = ( wire5535 ) | ( wire5536 ) | ( wire16093 ) ;
 assign wire16098 = ( wire16089 ) | ( wire16090 ) | ( wire16091 ) | ( wire16092 ) ;
 assign wire16106 = ( n_n9232  &  wire2381 ) | ( n_n8233  &  wire2383 ) ;
 assign wire16107 = ( wire5500 ) | ( wire5501 ) | ( n_n7822  &  wire2380 ) ;
 assign wire16108 = ( wire5502 ) | ( wire5503 ) | ( wire5504 ) | ( wire5505 ) ;
 assign wire16109 = ( wire5506 ) | ( wire5507 ) | ( wire5508 ) | ( wire5509 ) ;
 assign wire16110 = ( wire5510 ) | ( wire5511 ) | ( wire5512 ) | ( wire5513 ) ;
 assign wire16114 = ( wire5495 ) | ( wire5496 ) | ( wire16110 ) ;
 assign wire16115 = ( wire16106 ) | ( wire16107 ) | ( wire16108 ) | ( wire16109 ) ;
 assign wire16122 = ( n_n7600  &  wire2375 ) | ( n_n7823  &  wire2377 ) ;
 assign wire16123 = ( n_n8736  &  wire2373 ) | ( n_n7821  &  wire2374 ) ;
 assign wire16124 = ( wire5483 ) | ( wire5484 ) | ( wire5485 ) | ( wire5486 ) ;
 assign wire16125 = ( wire5487 ) | ( wire5488 ) | ( wire5489 ) | ( wire5490 ) ;
 assign wire16126 = ( wire5491 ) | ( wire5492 ) | ( wire5493 ) | ( wire5494 ) ;
 assign wire16130 = ( wire5477 ) | ( wire5478 ) | ( wire16126 ) ;
 assign wire16131 = ( wire16122 ) | ( wire16123 ) | ( wire16124 ) | ( wire16125 ) ;
 assign wire16138 = ( n_n9212  &  wire2375 ) | ( n_n9400  &  wire2377 ) ;
 assign wire16139 = ( n_n9137  &  wire2373 ) | ( n_n9397  &  wire2374 ) ;
 assign wire16140 = ( wire5463 ) | ( wire5464 ) | ( wire5465 ) | ( wire5466 ) ;
 assign wire16141 = ( wire5467 ) | ( wire5468 ) | ( wire5469 ) | ( wire5470 ) ;
 assign wire16142 = ( wire5471 ) | ( wire5472 ) | ( wire5473 ) | ( wire5474 ) ;
 assign wire16146 = ( wire5457 ) | ( wire5458 ) | ( wire16142 ) ;
 assign wire16147 = ( wire16138 ) | ( wire16139 ) | ( wire16140 ) | ( wire16141 ) ;
 assign wire16155 = ( n_n9396  &  wire2381 ) | ( n_n9402  &  wire2383 ) ;
 assign wire16156 = ( wire5324 ) | ( wire5325 ) | ( n_n9398  &  wire2380 ) ;
 assign wire16157 = ( wire5326 ) | ( wire5327 ) | ( wire5328 ) | ( wire5329 ) ;
 assign wire16158 = ( wire5330 ) | ( wire5331 ) | ( wire5332 ) | ( wire5333 ) ;
 assign wire16159 = ( wire5334 ) | ( wire5335 ) | ( wire5336 ) | ( wire5337 ) ;
 assign wire16163 = ( wire5319 ) | ( wire5320 ) | ( wire16159 ) ;
 assign wire16164 = ( wire16155 ) | ( wire16156 ) | ( wire16157 ) | ( wire16158 ) ;
 assign wire16171 = ( n_n8638  &  wire2375 ) | ( n_n7741  &  wire2377 ) ;
 assign wire16172 = ( n_n8009  &  wire2373 ) | ( n_n7738  &  wire2374 ) ;
 assign wire16173 = ( wire5445 ) | ( wire5446 ) | ( wire5447 ) | ( wire5448 ) ;
 assign wire16174 = ( wire5449 ) | ( wire5450 ) | ( wire5451 ) | ( wire5452 ) ;
 assign wire16175 = ( wire5453 ) | ( wire5454 ) | ( wire5455 ) | ( wire5456 ) ;
 assign wire16179 = ( wire5439 ) | ( wire5440 ) | ( wire16175 ) ;
 assign wire16180 = ( wire16171 ) | ( wire16172 ) | ( wire16173 ) | ( wire16174 ) ;
 assign wire16188 = ( n_n7737  &  wire2381 ) | ( n_n9528  &  wire2383 ) ;
 assign wire16189 = ( wire5347 ) | ( wire5348 ) | ( n_n7739  &  wire2380 ) ;
 assign wire16190 = ( wire5349 ) | ( wire5350 ) | ( wire5351 ) | ( wire5352 ) ;
 assign wire16191 = ( wire5353 ) | ( wire5354 ) | ( wire5355 ) | ( wire5356 ) ;
 assign wire16192 = ( wire5357 ) | ( wire5358 ) | ( wire5359 ) | ( wire5360 ) ;
 assign wire16196 = ( wire5342 ) | ( wire5343 ) | ( wire16192 ) ;
 assign wire16197 = ( wire16188 ) | ( wire16189 ) | ( wire16190 ) | ( wire16191 ) ;
 assign wire16204 = ( n_n9045  &  wire2375 ) | ( n_n9317  &  wire2377 ) ;
 assign wire16205 = ( n_n9054  &  wire2373 ) | ( n_n9315  &  wire2374 ) ;
 assign wire16206 = ( wire5408 ) | ( wire5409 ) | ( wire5410 ) | ( wire5411 ) ;
 assign wire16207 = ( wire5412 ) | ( wire5413 ) | ( wire5414 ) | ( wire5415 ) ;
 assign wire16208 = ( wire5416 ) | ( wire5417 ) | ( wire5418 ) | ( wire5419 ) ;
 assign wire16212 = ( wire5402 ) | ( wire5403 ) | ( wire16208 ) ;
 assign wire16213 = ( wire16204 ) | ( wire16205 ) | ( wire16206 ) | ( wire16207 ) ;
 assign wire16221 = ( n_n9314  &  wire2381 ) | ( n_n9319  &  wire2383 ) ;
 assign wire16222 = ( wire5425 ) | ( wire5426 ) | ( n_n9368  &  wire2380 ) ;
 assign wire16223 = ( wire5427 ) | ( wire5428 ) | ( wire5429 ) | ( wire5430 ) ;
 assign wire16224 = ( wire5431 ) | ( wire5432 ) | ( wire5433 ) | ( wire5434 ) ;
 assign wire16225 = ( wire5435 ) | ( wire5436 ) | ( wire5437 ) | ( wire5438 ) ;
 assign wire16229 = ( wire5420 ) | ( wire5421 ) | ( wire16225 ) ;
 assign wire16230 = ( wire16221 ) | ( wire16222 ) | ( wire16223 ) | ( wire16224 ) ;
 assign wire16237 = ( n_n7509  &  wire2375 ) | ( n_n7654  &  wire2377 ) ;
 assign wire16238 = ( n_n8011  &  wire2373 ) | ( n_n7652  &  wire2374 ) ;
 assign wire16239 = ( wire5388 ) | ( wire5389 ) | ( wire5390 ) | ( wire5391 ) ;
 assign wire16240 = ( wire5392 ) | ( wire5393 ) | ( wire5394 ) | ( wire5395 ) ;
 assign wire16241 = ( wire5396 ) | ( wire5397 ) | ( wire5398 ) | ( wire5399 ) ;
 assign wire16245 = ( wire5382 ) | ( wire5383 ) | ( wire16241 ) ;
 assign wire16246 = ( wire16237 ) | ( wire16238 ) | ( wire16239 ) | ( wire16240 ) ;
 assign wire16254 = ( n_n8033  &  wire2381 ) | ( n_n7661  &  wire2383 ) ;
 assign wire16255 = ( wire5368 ) | ( wire5369 ) | ( n_n7728  &  wire2380 ) ;
 assign wire16256 = ( wire5370 ) | ( wire5371 ) | ( wire5372 ) | ( wire5373 ) ;
 assign wire16257 = ( wire5374 ) | ( wire5375 ) | ( wire5376 ) | ( wire5377 ) ;
 assign wire16258 = ( wire5378 ) | ( wire5379 ) | ( wire5380 ) | ( wire5381 ) ;
 assign wire16262 = ( wire5363 ) | ( wire5364 ) | ( wire16258 ) ;
 assign wire16263 = ( wire16254 ) | ( wire16255 ) | ( wire16256 ) | ( wire16257 ) ;
 assign wire16270 = ( n_n9262  &  wire2375 ) | ( n_n9598  &  wire2377 ) ;
 assign wire16271 = ( n_n9271  &  wire2373 ) | ( n_n9595  &  wire2374 ) ;
 assign wire16272 = ( wire5276 ) | ( wire5277 ) | ( wire5278 ) | ( wire5279 ) ;
 assign wire16273 = ( wire5280 ) | ( wire5281 ) | ( wire5282 ) | ( wire5283 ) ;
 assign wire16274 = ( wire5284 ) | ( wire5285 ) | ( wire5286 ) | ( wire5287 ) ;
 assign wire16278 = ( wire5270 ) | ( wire5271 ) | ( wire16274 ) ;
 assign wire16279 = ( wire16270 ) | ( wire16271 ) | ( wire16272 ) | ( wire16273 ) ;
 assign wire16287 = ( n_n9594  &  wire2381 ) | ( n_n9600  &  wire2383 ) ;
 assign wire16288 = ( wire5256 ) | ( wire5257 ) | ( n_n9596  &  wire2380 ) ;
 assign wire16289 = ( wire5258 ) | ( wire5259 ) | ( wire5260 ) | ( wire5261 ) ;
 assign wire16290 = ( wire5262 ) | ( wire5263 ) | ( wire5264 ) | ( wire5265 ) ;
 assign wire16291 = ( wire5266 ) | ( wire5267 ) | ( wire5268 ) | ( wire5269 ) ;
 assign wire16295 = ( wire5251 ) | ( wire5252 ) | ( wire16291 ) ;
 assign wire16296 = ( wire16287 ) | ( wire16288 ) | ( wire16289 ) | ( wire16290 ) ;
 assign wire16303 = ( n_n7665  &  wire2375 ) | ( n_n7686  &  wire2377 ) ;
 assign wire16304 = ( n_n8110  &  wire2373 ) | ( n_n7683  &  wire2374 ) ;
 assign wire16305 = ( wire5130 ) | ( wire5131 ) | ( wire5132 ) | ( wire5133 ) ;
 assign wire16306 = ( wire5134 ) | ( wire5135 ) | ( wire5136 ) | ( wire5137 ) ;
 assign wire16307 = ( wire5138 ) | ( wire5139 ) | ( wire5140 ) | ( wire5141 ) ;
 assign wire16311 = ( wire5124 ) | ( wire5125 ) | ( wire16307 ) ;
 assign wire16312 = ( wire16303 ) | ( wire16304 ) | ( wire16305 ) | ( wire16306 ) ;
 assign wire16320 = ( n_n8586  &  wire2381 ) | ( n_n7687  &  wire2383 ) ;
 assign wire16321 = ( wire5147 ) | ( wire5148 ) | ( n_n7684  &  wire2380 ) ;
 assign wire16322 = ( wire5149 ) | ( wire5150 ) | ( wire5151 ) | ( wire5152 ) ;
 assign wire16323 = ( wire5153 ) | ( wire5154 ) | ( wire5155 ) | ( wire5156 ) ;
 assign wire16324 = ( wire5157 ) | ( wire5158 ) | ( wire5159 ) | ( wire5160 ) ;
 assign wire16328 = ( wire5142 ) | ( wire5143 ) | ( wire16324 ) ;
 assign wire16329 = ( wire16320 ) | ( wire16321 ) | ( wire16322 ) | ( wire16323 ) ;
 assign wire16336 = ( n_n9336  &  wire2375 ) | ( n_n9342  &  wire2377 ) ;
 assign wire16337 = ( n_n9349  &  wire2373 ) | ( n_n9338  &  wire2374 ) ;
 assign wire16338 = ( wire5233 ) | ( wire5234 ) | ( wire5235 ) | ( wire5236 ) ;
 assign wire16339 = ( wire5237 ) | ( wire5238 ) | ( wire5239 ) | ( wire5240 ) ;
 assign wire16340 = ( wire5241 ) | ( wire5242 ) | ( wire5243 ) | ( wire5244 ) ;
 assign wire16344 = ( wire5227 ) | ( wire5228 ) | ( wire16340 ) ;
 assign wire16345 = ( wire16336 ) | ( wire16337 ) | ( wire16338 ) | ( wire16339 ) ;
 assign wire16353 = ( n_n6976  &  wire2381 ) | ( n_n9343  &  wire2383 ) ;
 assign wire16354 = ( wire5170 ) | ( wire5171 ) | ( n_n9339  &  wire2380 ) ;
 assign wire16355 = ( wire5172 ) | ( wire5173 ) | ( wire5174 ) | ( wire5175 ) ;
 assign wire16356 = ( wire5176 ) | ( wire5177 ) | ( wire5178 ) | ( wire5179 ) ;
 assign wire16357 = ( wire5180 ) | ( wire5181 ) | ( wire5182 ) | ( wire5183 ) ;
 assign wire16361 = ( wire5165 ) | ( wire5166 ) | ( wire16357 ) ;
 assign wire16362 = ( wire16353 ) | ( wire16354 ) | ( wire16355 ) | ( wire16356 ) ;
 assign wire16369 = ( n_n7692  &  wire2375 ) | ( n_n9021  &  wire2377 ) ;
 assign wire16370 = ( n_n7697  &  wire2373 ) | ( n_n9618  &  wire2374 ) ;
 assign wire16371 = ( wire5215 ) | ( wire5216 ) | ( wire5217 ) | ( wire5218 ) ;
 assign wire16372 = ( wire5219 ) | ( wire5220 ) | ( wire5221 ) | ( wire5222 ) ;
 assign wire16373 = ( wire5223 ) | ( wire5224 ) | ( wire5225 ) | ( wire5226 ) ;
 assign wire16377 = ( wire5209 ) | ( wire5210 ) | ( wire16373 ) ;
 assign wire16378 = ( wire16369 ) | ( wire16370 ) | ( wire16371 ) | ( wire16372 ) ;
 assign wire16386 = ( n_n8966  &  wire2381 ) | ( n_n7952  &  wire2383 ) ;
 assign wire16387 = ( wire5193 ) | ( wire5194 ) | ( n_n8854  &  wire2380 ) ;
 assign wire16388 = ( wire5195 ) | ( wire5196 ) | ( wire5197 ) | ( wire5198 ) ;
 assign wire16389 = ( wire5199 ) | ( wire5200 ) | ( wire5201 ) | ( wire5202 ) ;
 assign wire16390 = ( wire5203 ) | ( wire5204 ) | ( wire5205 ) | ( wire5206 ) ;
 assign wire16394 = ( wire5188 ) | ( wire5189 ) | ( wire16390 ) ;
 assign wire16395 = ( wire16386 ) | ( wire16387 ) | ( wire16388 ) | ( wire16389 ) ;
 assign wire16402 = ( n_n7709  &  wire2375 ) | ( n_n7762  &  wire2377 ) ;
 assign wire16403 = ( n_n8986  &  wire2373 ) | ( n_n8852  &  wire2374 ) ;
 assign wire16404 = ( wire5108 ) | ( wire5109 ) | ( wire5110 ) | ( wire5111 ) ;
 assign wire16405 = ( wire5112 ) | ( wire5113 ) | ( wire5114 ) | ( wire5115 ) ;
 assign wire16406 = ( wire5116 ) | ( wire5117 ) | ( wire5118 ) | ( wire5119 ) ;
 assign wire16410 = ( wire5102 ) | ( wire5103 ) | ( wire16406 ) ;
 assign wire16411 = ( wire16402 ) | ( wire16403 ) | ( wire16404 ) | ( wire16405 ) ;
 assign wire16419 = ( n_n7759  &  wire2381 ) | ( n_n7763  &  wire2383 ) ;
 assign wire16420 = ( wire5088 ) | ( wire5089 ) | ( n_n7760  &  wire2380 ) ;
 assign wire16421 = ( wire5090 ) | ( wire5091 ) | ( wire5092 ) | ( wire5093 ) ;
 assign wire16422 = ( wire5094 ) | ( wire5095 ) | ( wire5096 ) | ( wire5097 ) ;
 assign wire16423 = ( wire5098 ) | ( wire5099 ) | ( wire5100 ) | ( wire5101 ) ;
 assign wire16427 = ( wire5083 ) | ( wire5084 ) | ( wire16423 ) ;
 assign wire16428 = ( wire16419 ) | ( wire16420 ) | ( wire16421 ) | ( wire16422 ) ;
 assign wire16437 = ( n_n8408  &  wire2381 ) | ( n_n7811  &  wire2383 ) ;
 assign wire16438 = ( wire5037 ) | ( wire5038 ) | ( n_n7809  &  wire2380 ) ;
 assign wire16439 = ( wire5039 ) | ( wire5040 ) | ( wire5041 ) | ( wire5042 ) ;
 assign wire16440 = ( wire5043 ) | ( wire5044 ) | ( wire5045 ) | ( wire5046 ) ;
 assign wire16441 = ( wire5047 ) | ( wire5048 ) | ( wire5049 ) | ( wire5050 ) ;
 assign wire16445 = ( wire5032 ) | ( wire5033 ) | ( wire16441 ) ;
 assign wire16446 = ( wire16437 ) | ( wire16438 ) | ( wire16439 ) | ( wire16440 ) ;
 assign wire16453 = ( n_n8088  &  wire2375 ) | ( n_n7810  &  wire2377 ) ;
 assign wire16454 = ( n_n8108  &  wire2373 ) | ( n_n8473  &  wire2374 ) ;
 assign wire16455 = ( wire5057 ) | ( wire5058 ) | ( wire5059 ) | ( wire5060 ) ;
 assign wire16456 = ( wire5061 ) | ( wire5062 ) | ( wire5063 ) | ( wire5064 ) ;
 assign wire16457 = ( wire5065 ) | ( wire5066 ) | ( wire5067 ) | ( wire5068 ) ;
 assign wire16461 = ( wire5051 ) | ( wire5052 ) | ( wire16457 ) ;
 assign wire16462 = ( wire16453 ) | ( wire16454 ) | ( wire16455 ) | ( wire16456 ) ;
 assign wire16463 = ( n_n9248  &  (~ n_n7306) ) ;
 assign wire16464 = ( nsr3_23  &  ndn3_19 ) | ( nsr3_38  &  nen3_36 ) ;
 assign wire16465 = ( nsr3_37  &  nen3_34 ) | ( nsr3_30  &  ndn3_26 ) ;
 assign wire16466 = ( ndn3_29  &  nsr3_35 ) | ( ndn3_17  &  nsr3_20 ) ;
 assign wire16469 = ( n_n9197  &  n_n9198 ) ;
 assign wire16473 = ( wire4997 ) | ( wire4998 ) | ( wire4999 ) ;
 assign wire16474 = ( wire5000 ) | ( wire5001 ) | ( wire5002 ) | ( wire5003 ) ;
 assign wire16478 = ( wire4990 ) | ( wire4991 ) | ( wire4992 ) ;
 assign wire16479 = ( wire4993 ) | ( wire4994 ) | ( wire4995 ) | ( wire4996 ) ;
 assign wire16483 = ( wire4976 ) | ( wire4977 ) | ( wire4978 ) ;
 assign wire16484 = ( wire4979 ) | ( wire4980 ) | ( wire4981 ) | ( wire4982 ) ;
 assign wire16488 = ( wire4955 ) | ( wire4956 ) | ( wire4957 ) ;
 assign wire16489 = ( wire4958 ) | ( wire4959 ) | ( wire4960 ) | ( wire4961 ) ;
 assign wire16493 = ( wire4948 ) | ( wire4949 ) | ( wire4950 ) ;
 assign wire16494 = ( wire4951 ) | ( wire4952 ) | ( wire4953 ) | ( wire4954 ) ;
 assign wire16498 = ( wire4927 ) | ( wire4928 ) | ( wire4929 ) ;
 assign wire16499 = ( wire4930 ) | ( wire4931 ) | ( wire4932 ) | ( wire4933 ) ;
 assign wire16503 = ( wire4934 ) | ( wire4935 ) | ( wire4936 ) ;
 assign wire16504 = ( wire4937 ) | ( wire4938 ) | ( wire4939 ) | ( wire4940 ) ;
 assign wire16508 = ( wire4918 ) | ( wire4919 ) | ( wire4920 ) ;
 assign wire16509 = ( wire4921 ) | ( wire4922 ) | ( wire4923 ) | ( wire4924 ) ;
 assign wire16513 = ( wire4941 ) | ( wire4942 ) | ( wire4943 ) ;
 assign wire16514 = ( wire4944 ) | ( wire4945 ) | ( wire4946 ) | ( wire4947 ) ;
 assign wire16518 = ( wire4962 ) | ( wire4963 ) | ( wire4964 ) ;
 assign wire16519 = ( wire4965 ) | ( wire4966 ) | ( wire4967 ) | ( wire4968 ) ;
 assign wire16523 = ( wire4969 ) | ( wire4970 ) | ( wire4971 ) ;
 assign wire16524 = ( wire4972 ) | ( wire4973 ) | ( wire4974 ) | ( wire4975 ) ;
 assign wire16528 = ( wire4899 ) | ( wire4900 ) | ( wire4901 ) ;
 assign wire16529 = ( wire4902 ) | ( wire4903 ) | ( wire4904 ) | ( wire4905 ) ;
 assign wire16533 = ( wire4983 ) | ( wire4984 ) | ( wire4985 ) ;
 assign wire16534 = ( wire4986 ) | ( wire4987 ) | ( wire4988 ) | ( wire4989 ) ;
 assign wire16538 = ( wire4886 ) | ( wire4887 ) | ( wire4888 ) ;
 assign wire16539 = ( wire4889 ) | ( wire4890 ) | ( wire4891 ) | ( wire4892 ) ;
 assign wire16543 = ( wire4877 ) | ( wire4878 ) | ( wire4879 ) ;
 assign wire16544 = ( wire4880 ) | ( wire4881 ) | ( wire4882 ) | ( wire4883 ) ;
 assign wire16549 = ( wire4867 ) | ( wire4868 ) | ( wire4869 ) | ( wire4870 ) ;
 assign wire16550 = ( (~ n_n8557)  &  wire2363  &  n_n7274 ) ;
 assign wire16551 = ( wire2363  &  n_n8557 ) ;
 assign wire16554 = ( n_n9638  &  wire2363  &  wire16483 ) | ( n_n9638  &  wire2363  &  wire16484 ) ;
 assign wire16565 = ( n_n9225  &  wire2375 ) | ( n_n7888  &  wire2377 ) ;
 assign wire16566 = ( n_n7850  &  wire2373 ) | ( n_n7887  &  wire2374 ) ;
 assign wire16567 = ( wire4793 ) | ( wire4794 ) | ( wire4795 ) | ( wire4796 ) ;
 assign wire16568 = ( wire4797 ) | ( wire4798 ) | ( wire4799 ) | ( wire4800 ) ;
 assign wire16569 = ( wire4801 ) | ( wire4802 ) | ( wire4803 ) | ( wire4804 ) ;
 assign wire16573 = ( wire4787 ) | ( wire4788 ) | ( wire16569 ) ;
 assign wire16574 = ( wire16565 ) | ( wire16566 ) | ( wire16567 ) | ( wire16568 ) ;
 assign wire16582 = ( n_n7886  &  wire2381 ) | ( n_n7889  &  wire2383 ) ;
 assign wire16583 = ( wire4773 ) | ( wire4774 ) | ( n_n9520  &  wire2380 ) ;
 assign wire16584 = ( wire4775 ) | ( wire4776 ) | ( wire4777 ) | ( wire4778 ) ;
 assign wire16585 = ( wire4779 ) | ( wire4780 ) | ( wire4781 ) | ( wire4782 ) ;
 assign wire16586 = ( wire4783 ) | ( wire4784 ) | ( wire4785 ) | ( wire4786 ) ;
 assign wire16590 = ( wire4768 ) | ( wire4769 ) | ( wire16586 ) ;
 assign wire16591 = ( wire16582 ) | ( wire16583 ) | ( wire16584 ) | ( wire16585 ) ;
 assign wire16599 = ( n_n8002  &  wire2381 ) | ( n_n8519  &  wire2383 ) ;
 assign wire16600 = ( wire4740 ) | ( wire4741 ) | ( n_n8004  &  wire2380 ) ;
 assign wire16601 = ( wire4742 ) | ( wire4743 ) | ( wire4744 ) | ( wire4745 ) ;
 assign wire16602 = ( wire4746 ) | ( wire4747 ) | ( wire4748 ) | ( wire4749 ) ;
 assign wire16603 = ( wire4750 ) | ( wire4751 ) | ( wire4752 ) | ( wire4753 ) ;
 assign wire16607 = ( wire4735 ) | ( wire4736 ) | ( wire16603 ) ;
 assign wire16608 = ( wire16599 ) | ( wire16600 ) | ( wire16601 ) | ( wire16602 ) ;
 assign wire16615 = ( n_n9223  &  wire2375 ) | ( n_n8005  &  wire2377 ) ;
 assign wire16616 = ( n_n8482  &  wire2373 ) | ( n_n8003  &  wire2374 ) ;
 assign wire16617 = ( wire4723 ) | ( wire4724 ) | ( wire4725 ) | ( wire4726 ) ;
 assign wire16618 = ( wire4727 ) | ( wire4728 ) | ( wire4729 ) | ( wire4730 ) ;
 assign wire16619 = ( wire4731 ) | ( wire4732 ) | ( wire4733 ) | ( wire4734 ) ;
 assign wire16623 = ( wire4717 ) | ( wire4718 ) | ( wire16619 ) ;
 assign wire16624 = ( wire16615 ) | ( wire16616 ) | ( wire16617 ) | ( wire16618 ) ;
 assign wire16631 = ( n_n8139  &  wire2375 ) | ( n_n7933  &  wire2377 ) ;
 assign wire16632 = ( n_n8000  &  wire2373 ) | ( n_n7931  &  wire2374 ) ;
 assign wire16633 = ( wire4684 ) | ( wire4685 ) | ( wire4686 ) | ( wire4687 ) ;
 assign wire16634 = ( wire4688 ) | ( wire4689 ) | ( wire4690 ) | ( wire4691 ) ;
 assign wire16635 = ( wire4692 ) | ( wire4693 ) | ( wire4694 ) | ( wire4695 ) ;
 assign wire16639 = ( wire4678 ) | ( wire4679 ) | ( wire16635 ) ;
 assign wire16640 = ( wire16631 ) | ( wire16632 ) | ( wire16633 ) | ( wire16634 ) ;
 assign wire16648 = ( n_n7930  &  wire2381 ) | ( n_n8106  &  wire2383 ) ;
 assign wire16649 = ( wire4701 ) | ( wire4702 ) | ( n_n7932  &  wire2380 ) ;
 assign wire16650 = ( wire4703 ) | ( wire4704 ) | ( wire4705 ) | ( wire4706 ) ;
 assign wire16651 = ( wire4707 ) | ( wire4708 ) | ( wire4709 ) | ( wire4710 ) ;
 assign wire16652 = ( wire4711 ) | ( wire4712 ) | ( wire4713 ) | ( wire4714 ) ;
 assign wire16656 = ( wire4696 ) | ( wire4697 ) | ( wire16652 ) ;
 assign wire16657 = ( wire16648 ) | ( wire16649 ) | ( wire16650 ) | ( wire16651 ) ;
 assign wire16661 = ( (~ n_n8603)  &  (~ n_n8798)  &  (~ n_n8869) ) ;
 assign wire16662 = ( (~ n_n8933)  &  (~ n_n8876)  &  n_n8694  &  n_n8932 ) | ( n_n8933  &  (~ n_n8876)  &  n_n8694  &  (~ n_n8932) ) ;
 assign wire16663 = ( (~ n_n8911)  &  n_n8933  &  wire16661 ) | ( (~ n_n8911)  &  n_n8932  &  wire16661 ) | ( n_n8911  &  (~ n_n8933)  &  (~ n_n8932)  &  wire16661 ) ;
 assign wire16664 = ( (~ n_n8976)  &  wire16662 ) ;
 assign wire16667 = ( (~ n_n8993)  &  (~ n_n7637)  &  n_n8204  &  wire16663 ) | ( n_n8993  &  (~ n_n7637)  &  (~ n_n8204)  &  wire16663 ) ;
 assign wire16668 = ( (~ n_n8561)  &  (~ n_n9029)  &  n_n8342  &  wire16664 ) | ( n_n8561  &  (~ n_n9029)  &  (~ n_n8342)  &  wire16664 ) ;
 assign wire16670 = ( (~ n_n9152)  &  wire16668 ) ;
 assign wire16671 = ( (~ n_n8913)  &  (~ n_n8403)  &  n_n8493  &  wire16667 ) | ( n_n8913  &  (~ n_n8403)  &  (~ n_n8493)  &  wire16667 ) ;
 assign wire16674 = ( preset ) | ( (~ n_n9198) ) | ( (~ n_n9639) ) | ( (~ n_n9197) ) ;
 assign wire16676 = ( n_n9434  &  wire2363  &  wire16488 ) | ( n_n9434  &  wire2363  &  wire16489 ) ;
 assign wire16682 = ( (~ n_n9639)  &  (~ preset) ) ;
 assign wire16686 = ( preset ) | ( pdn ) | ( nsr3_23  &  (~ nak3_13) ) ;
 assign wire16687 = ( preset ) | ( pdn ) | ( nsr3_13  &  (~ nak3_13) ) ;
 assign wire16688 = ( preset ) | ( pdn ) | ( nsr3_38  &  (~ nak3_13) ) ;
 assign wire16690 = ( n_n8549  &  wire2363  &  wire16473 ) | ( n_n8549  &  wire2363  &  wire16474 ) ;
 assign wire16698 = ( n_n8652  &  wire2363  &  (~ n_n8653) ) | ( (~ n_n8652)  &  wire2363  &  n_n8653  &  n_n7274 ) ;
 assign wire16701 = ( (~ n_n8707)  &  (~ n_n8706)  &  wire16508 ) | ( (~ n_n8707)  &  (~ n_n8706)  &  wire16509 ) | ( (~ n_n8707)  &  n_n8706  &  (~ wire16508)  &  (~ wire16509) ) ;
 assign wire16703 = ( n_n8707  &  wire2363  &  n_n8706  &  n_n8708 ) | ( n_n8707  &  wire2363  &  (~ n_n8706)  &  (~ n_n8708) ) ;
 assign wire16704 = ( wire16703 ) | ( wire2363  &  n_n7274  &  wire16701 ) ;
 assign wire16705 = ( preset ) | ( pdn ) | ( nsr3_30  &  (~ ndn3_26) ) ;
 assign wire16707 = ( n_n8354  &  wire2363  &  wire16538 ) | ( n_n8354  &  wire2363  &  wire16539 ) ;
 assign wire16714 = ( n_n9512  &  wire2363  &  wire16493 ) | ( n_n9512  &  wire2363  &  wire16494 ) ;
 assign wire16715 = ( wire2363  &  wire2460  &  n_n7274 ) ;
 assign wire16716 = ( wire2363  &  n_n9512 ) ;
 assign wire16717 = ( wire3715 ) | ( (~ preset)  &  n_n9512  &  (~ n_n7274) ) ;
 assign wire16719 = ( preset ) | ( pdn ) | ( nsr3_35  &  (~ nak3_13) ) ;
 assign wire16721 = ( n_n9416  &  wire2363  &  wire16518 ) | ( n_n9416  &  wire2363  &  wire16519 ) ;
 assign wire16726 = ( pdn ) | ( preset  &  (~ nak3_13) ) | ( (~ nak3_13)  &  nsr3_14 ) ;
 assign wire16727 = ( (~ n_n8603)  &  (~ n_n8667)  &  (~ wire4421) ) | ( (~ n_n8603)  &  (~ wire4421)  &  (~ wire16682) ) ;
 assign wire16728 = ( (~ n_n8603)  &  (~ wire15947)  &  (~ wire15948) ) ;
 assign wire16729 = ( (~ wire2363)  &  n_n8603 ) ;
 assign wire16732 = ( (~ wire2451)  &  wire16727 ) | ( (~ wire2451)  &  wire16728 ) ;
 assign wire16734 = ( (~ preset)  &  n_n9198  &  n_n9639  &  n_n9197 ) ;
 assign wire16742 = ( n_n8449  &  wire2363  &  wire16478 ) | ( n_n8449  &  wire2363  &  wire16479 ) ;
 assign wire16748 = ( n_n9448  &  wire2363  &  wire16533 ) | ( n_n9448  &  wire2363  &  wire16534 ) ;
 assign wire16754 = ( n_n9537  &  wire2363  &  wire16523 ) | ( n_n9537  &  wire2363  &  wire16524 ) ;
 assign wire16759 = ( n_n8929  &  (~ preset) ) ;
 assign wire16760 = ( (~ preset)  &  wire16027 ) | ( (~ preset)  &  wire16028 ) ;
 assign wire16763 = ( (~ n_n9284)  &  (~ n_n8537)  &  wire16503 ) | ( (~ n_n9284)  &  (~ n_n8537)  &  wire16504 ) | ( (~ n_n9284)  &  n_n8537  &  (~ wire16503)  &  (~ wire16504) ) ;
 assign wire16765 = ( n_n9284  &  wire2363  &  n_n8537  &  n_n8740 ) | ( n_n9284  &  wire2363  &  (~ n_n8537)  &  (~ n_n8740) ) ;
 assign wire16766 = ( wire16765 ) | ( wire2363  &  n_n7274  &  wire16763 ) ;
 assign wire16768 = ( n_n8821  &  wire2363  &  wire16528 ) | ( n_n8821  &  wire2363  &  wire16529 ) ;
 assign wire16775 = ( (~ n_n9353)  &  (~ n_n8484)  &  wire16513 ) | ( (~ n_n9353)  &  (~ n_n8484)  &  wire16514 ) | ( (~ n_n9353)  &  n_n8484  &  (~ wire16513)  &  (~ wire16514) ) ;
 assign wire16777 = ( n_n9353  &  wire2363  &  n_n8484  &  n_n8807 ) | ( n_n9353  &  wire2363  &  (~ n_n8484)  &  (~ n_n8807) ) ;
 assign wire16782 = ( preset ) | ( pdn ) | ( nsr3_37  &  (~ nen3_34) ) ;
 assign wire16786 = ( preset ) | ( pdn ) | ( (~ nak3_13)  &  nsr3_20 ) ;
 assign wire16790 = ( n_n8419  &  wire2363  &  wire16543 ) | ( n_n8419  &  wire2363  &  wire16544 ) ;


endmodule

