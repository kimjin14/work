module tseng (
	i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, 
	i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, 
	o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, 
	o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, 
	o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_43_, 
	o_30_, o_44_, o_41_, o_42_, o_20_, o_45_, o_10_, o_9_, o_7_, o_8_, 
	o_5_, o_6_, o_3_, o_4_);

input i_9_;
input i_10_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_14_;
input i_3_;
input i_13_;
input i_4_;
input i_12_;
input i_1_;
input i_11_;
input i_2_;
input i_0_;
input i_15_;
output o_1_;
output o_19_;
output o_2_;
output o_0_;
output o_29_;
output o_39_;
output o_38_;
output o_25_;
output o_12_;
output o_37_;
output o_26_;
output o_11_;
output o_36_;
output o_27_;
output o_14_;
output o_35_;
output o_28_;
output o_13_;
output o_34_;
output o_21_;
output o_16_;
output o_40_;
output o_33_;
output o_22_;
output o_15_;
output o_32_;
output o_23_;
output o_18_;
output o_31_;
output o_24_;
output o_17_;
output o_43_;
output o_30_;
output o_44_;
output o_41_;
output o_42_;
output o_20_;
output o_45_;
output o_10_;
output o_9_;
output o_7_;
output o_8_;
output o_5_;
output o_6_;
output o_3_;
output o_4_;
wire wire428;
wire n_n5144;
wire wire736;
wire n_n162;
wire n_n65;
wire n_n71;
wire n_n9;
wire wire343;
wire n_n38;
wire n_n373;
wire n_n374;
wire n_n969;
wire n_n4721;
wire n_n519;
wire n_n4597;
wire wire140;
wire wire390;
wire wire393;
wire wire712;
wire n_n31;
wire n_n30;
wire n_n4161;
wire wire132;
wire wire137;
wire wire599;
wire wire695;
wire n_n17;
wire n_n2229;
wire n_n2220;
wire n_n2232;
wire n_n2227;
wire n_n2226;
wire n_n2228;
wire n_n2234;
wire n_n4106;
wire n_n7241;
wire n_n7240;
wire n_n51;
wire n_n13;
wire n_n4;
wire wire77;
wire wire431;
wire wire529;
wire wire568;
wire wire569;
wire n_n53;
wire n_n3795;
wire n_n3787;
wire n_n3789;
wire wire157;
wire wire213;
wire n_n36;
wire n_n34;
wire n_n2622;
wire n_n3454;
wire n_n3456;
wire n_n7263;
wire n_n14;
wire n_n7265;
wire n_n7267;
wire n_n2998;
wire wire253;
wire n_n4308;
wire n_n6271;
wire n_n6267;
wire n_n3085;
wire n_n6266;
wire n_n6270;
wire n_n6269;
wire n_n6268;
wire n_n5052;
wire n_n5055;
wire wire608;
wire n_n10;
wire wire525;
wire n_n33;
wire n_n2732;
wire n_n2728;
wire n_n2721;
wire wire587;
wire wire767;
wire n_n6;
wire n_n135;
wire wire267;
wire n_n3389;
wire n_n5;
wire wire145;
wire wire388;
wire wire770;
wire n_n3166;
wire n_n144;
wire n_n7346;
wire n_n3;
wire n_n2;
wire wire708;
wire n_n18;
wire n_n5319;
wire wire430;
wire wire684;
wire wire748;
wire n_n16;
wire n_n197;
wire n_n212;
wire n_n2748;
wire n_n2747;
wire n_n101;
wire n_n42;
wire n_n4755;
wire wire172;
wire wire381;
wire wire662;
wire n_n3028;
wire n_n4845;
wire n_n184;
wire n_n163;
wire n_n161;
wire n_n6005;
wire wire419;
wire wire445;
wire wire446;
wire n_n3179;
wire wire95;
wire n_n743;
wire wire777;
wire wire776;
wire wire775;
wire wire185;
wire n_n7252;
wire n_n7253;
wire wire389;
wire wire454;
wire wire706;
wire wire742;
wire wire779;
wire wire783;
wire wire781;
wire wire707;
wire n_n46;
wire wire168;
wire n_n47;
wire n_n138;
wire wire214;
wire n_n5107;
wire n_n41;
wire wire245;
wire n_n108;
wire n_n148;
wire wire90;
wire n_n5000;
wire n_n1434;
wire n_n1408;
wire wire789;
wire n_n1426;
wire wire791;
wire n_n1416;
wire wire793;
wire wire422;
wire wire797;
wire wire796;
wire wire55;
wire wire207;
wire n_n1520;
wire wire800;
wire wire799;
wire n_n4581;
wire wire458;
wire wire541;
wire n_n125;
wire n_n3912;
wire n_n123;
wire wire570;
wire n_n1700;
wire wire803;
wire n_n4139;
wire n_n4206;
wire n_n1624;
wire wire85;
wire n_n4112;
wire n_n1594;
wire wire543;
wire wire808;
wire n_n4904;
wire n_n5037;
wire n_n4903;
wire wire544;
wire n_n4103;
wire wire52;
wire wire176;
wire n_n4007;
wire wire129;
wire wire142;
wire n_n4622;
wire wire182;
wire n_n5060;
wire n_n40;
wire n_n130;
wire wire134;
wire wire123;
wire n_n3276;
wire wire53;
wire n_n83;
wire n_n6445;
wire n_n7242;
wire n_n68;
wire wire344;
wire n_n19;
wire wire462;
wire wire817;
wire wire149;
wire wire130;
wire wire188;
wire n_n59;
wire wire226;
wire wire820;
wire wire819;
wire n_n2284;
wire n_n2241;
wire wire824;
wire n_n2253;
wire n_n61;
wire wire228;
wire wire827;
wire wire826;
wire n_n43;
wire wire139;
wire n_n117;
wire wire257;
wire wire313;
wire n_n129;
wire n_n166;
wire n_n127;
wire n_n39;
wire n_n82;
wire wire190;
wire wire334;
wire wire836;
wire n_n139;
wire wire838;
wire n_n1819;
wire n_n1870;
wire wire840;
wire n_n1800;
wire wire68;
wire n_n4591;
wire wire147;
wire wire98;
wire n_n2715;
wire n_n112;
wire n_n113;
wire wire844;
wire wire845;
wire wire542;
wire wire614;
wire wire850;
wire wire849;
wire n_n5109;
wire wire677;
wire wire852;
wire n_n140;
wire n_n142;
wire wire856;
wire n_n116;
wire wire255;
wire wire601;
wire wire859;
wire n_n157;
wire wire733;
wire wire743;
wire n_n213;
wire n_n199;
wire wire723;
wire wire729;
wire n_n95;
wire n_n200;
wire wire726;
wire n_n216;
wire wire724;
wire n_n103;
wire n_n191;
wire n_n89;
wire n_n207;
wire n_n177;
wire wire716;
wire n_n173;
wire n_n170;
wire wire720;
wire n_n169;
wire n_n204;
wire wire717;
wire wire730;
wire wire718;
wire n_n156;
wire wire722;
wire n_n154;
wire n_n205;
wire n_n150;
wire n_n149;
wire n_n151;
wire wire719;
wire wire721;
wire n_n141;
wire n_n115;
wire n_n209;
wire n_n134;
wire wire725;
wire n_n55;
wire wire728;
wire n_n54;
wire n_n126;
wire n_n124;
wire n_n92;
wire wire727;
wire n_n178;
wire n_n57;
wire wire715;
wire n_n48;
wire wire714;
wire n_n183;
wire n_n90;
wire n_n70;
wire n_n62;
wire n_n189;
wire n_n122;
wire n_n185;
wire n_n84;
wire n_n147;
wire n_n136;
wire n_n220;
wire n_n52;
wire n_n35;
wire n_n210;
wire n_n172;
wire n_n58;
wire n_n118;
wire n_n32;
wire n_n186;
wire n_n107;
wire n_n198;
wire n_n168;
wire n_n176;
wire n_n60;
wire n_n219;
wire n_n12;
wire n_n159;
wire wire151;
wire wire860;
wire n_n1442;
wire wire863;
wire wire865;
wire n_n4686;
wire wire247;
wire wire704;
wire n_n4231;
wire wire158;
wire wire155;
wire wire218;
wire wire180;
wire wire248;
wire n_n4460;
wire n_n4900;
wire wire867;
wire n_n4388;
wire n_n4441;
wire wire532;
wire wire575;
wire wire594;
wire wire660;
wire n_n4116;
wire wire156;
wire n_n77;
wire wire104;
wire n_n5111;
wire n_n5113;
wire wire868;
wire n_n7254;
wire n_n7248;
wire n_n3562;
wire wire63;
wire n_n3398;
wire wire143;
wire wire481;
wire n_n3050;
wire wire875;
wire n_n3033;
wire wire711;
wire wire878;
wire wire877;
wire wire879;
wire n_n2948;
wire n_n231;
wire wire308;
wire wire887;
wire wire189;
wire wire888;
wire wire896;
wire wire894;
wire wire561;
wire n_n2239;
wire wire899;
wire wire902;
wire wire133;
wire wire376;
wire wire904;
wire n_n1862;
wire wire583;
wire wire911;
wire n_n1799;
wire wire126;
wire wire913;
wire n_n2881;
wire n_n1708;
wire wire916;
wire n_n1717;
wire wire639;
wire wire564;
wire wire924;
wire n_n1170;
wire wire925;
wire wire928;
wire n_n4674;
wire n_n78;
wire n_n974;
wire wire933;
wire n_n7260;
wire n_n275;
wire wire551;
wire wire751;
wire n_n202;
wire n_n215;
wire n_n72;
wire n_n63;
wire n_n131;
wire n_n201;
wire n_n182;
wire n_n132;
wire n_n143;
wire n_n137;
wire n_n128;
wire n_n190;
wire n_n214;
wire n_n196;
wire n_n64;
wire n_n175;
wire n_n171;
wire n_n218;
wire n_n7264;
wire n_n74;
wire wire118;
wire wire566;
wire wire670;
wire n_n4808;
wire wire683;
wire wire524;
wire wire672;
wire n_n4564;
wire wire709;
wire n_n4169;
wire wire942;
wire n_n155;
wire wire60;
wire wire359;
wire n_n1514;
wire wire597;
wire n_n4996;
wire n_n4994;
wire wire511;
wire wire946;
wire n_n4120;
wire wire122;
wire wire443;
wire n_n4240;
wire n_n4154;
wire wire144;
wire wire654;
wire wire739;
wire wire279;
wire n_n4600;
wire n_n4602;
wire wire605;
wire wire146;
wire wire59;
wire n_n5075;
wire wire498;
wire wire951;
wire n_n6492;
wire wire152;
wire n_n3413;
wire wire546;
wire wire674;
wire n_n3889;
wire wire671;
wire wire463;
wire wire958;
wire wire960;
wire wire959;
wire n_n2813;
wire wire181;
wire n_n2265;
wire wire93;
wire wire968;
wire wire971;
wire n_n5739;
wire n_n2340;
wire n_n5743;
wire wire440;
wire wire447;
wire wire973;
wire n_n2259;
wire wire975;
wire wire979;
wire wire978;
wire wire980;
wire n_n2249;
wire wire397;
wire wire984;
wire wire989;
wire wire988;
wire wire993;
wire n_n1809;
wire wire685;
wire n_n5011;
wire wire81;
wire n_n1517;
wire wire457;
wire wire572;
wire wire1003;
wire wire1006;
wire n_n832;
wire wire1012;
wire wire1017;
wire n_n102;
wire n_n56;
wire n_n133;
wire n_n4915;
wire wire1021;
wire wire1023;
wire wire1022;
wire wire224;
wire n_n4981;
wire wire1030;
wire wire127;
wire wire70;
wire n_n4620;
wire n_n4131;
wire n_n4109;
wire wire249;
wire wire571;
wire wire620;
wire wire549;
wire wire621;
wire n_n4102;
wire n_n3417;
wire n_n6384;
wire n_n3419;
wire wire1036;
wire n_n3421;
wire wire391;
wire wire1042;
wire wire1041;
wire wire745;
wire wire231;
wire wire1044;
wire wire1049;
wire n_n2266;
wire wire526;
wire n_n2310;
wire wire1052;
wire wire1056;
wire n_n2257;
wire wire1060;
wire wire1064;
wire wire250;
wire wire227;
wire wire1069;
wire n_n5019;
wire wire1070;
wire n_n5033;
wire wire65;
wire wire111;
wire wire760;
wire wire1072;
wire wire1075;
wire wire1077;
wire wire1079;
wire n_n972;
wire wire48;
wire wire1084;
wire wire1089;
wire wire1087;
wire wire1090;
wire n_n259;
wire n_n164;
wire n_n111;
wire wire186;
wire n_n5103;
wire wire212;
wire n_n5067;
wire wire1096;
wire wire208;
wire wire591;
wire wire515;
wire wire657;
wire n_n4424;
wire wire518;
wire wire653;
wire wire694;
wire n_n4404;
wire wire503;
wire wire666;
wire n_n4397;
wire n_n4312;
wire wire141;
wire wire135;
wire n_n4476;
wire n_n4449;
wire n_n4566;
wire wire46;
wire wire51;
wire n_n1553;
wire wire209;
wire n_n5059;
wire n_n5058;
wire wire577;
wire wire1115;
wire wire1114;
wire wire1116;
wire wire1117;
wire wire1120;
wire wire1124;
wire wire1126;
wire wire1129;
wire wire1132;
wire wire1135;
wire wire74;
wire wire1136;
wire wire83;
wire wire384;
wire wire1143;
wire wire1145;
wire wire1147;
wire wire1150;
wire wire1152;
wire wire500;
wire wire1154;
wire wire1153;
wire n_n3415;
wire wire1160;
wire wire1159;
wire n_n7262;
wire n_n73;
wire n_n211;
wire wire150;
wire n_n1606;
wire wire1170;
wire n_n4623;
wire n_n3979;
wire wire361;
wire wire363;
wire wire426;
wire wire442;
wire wire1173;
wire wire1174;
wire wire1177;
wire wire1176;
wire wire1179;
wire wire1178;
wire wire377;
wire n_n4247;
wire wire655;
wire wire1190;
wire wire1189;
wire wire1188;
wire wire1194;
wire wire136;
wire wire364;
wire wire1197;
wire wire1196;
wire wire1195;
wire n_n1843;
wire n_n1826;
wire wire1200;
wire wire1199;
wire n_n1803;
wire n_n1824;
wire wire1201;
wire wire1205;
wire wire62;
wire wire1207;
wire wire1211;
wire n_n1542;
wire n_n4641;
wire wire693;
wire wire1214;
wire wire1216;
wire wire154;
wire wire1218;
wire n_n369;
wire wire335;
wire wire747;
wire wire100;
wire wire153;
wire wire234;
wire wire652;
wire n_n4518;
wire wire1224;
wire wire125;
wire n_n7266;
wire wire1229;
wire n_n3054;
wire wire131;
wire n_n2770;
wire wire1234;
wire wire412;
wire wire1239;
wire n_n1913;
wire n_n3638;
wire wire1242;
wire wire1244;
wire wire1243;
wire wire1246;
wire n_n1811;
wire wire1247;
wire wire1251;
wire wire1255;
wire wire1257;
wire n_n817;
wire wire167;
wire n_n799;
wire wire1259;
wire wire1261;
wire wire1260;
wire wire1263;
wire wire449;
wire wire656;
wire wire686;
wire wire1271;
wire n_n4692;
wire wire1277;
wire wire175;
wire wire383;
wire wire1279;
wire wire1281;
wire wire1285;
wire wire69;
wire wire276;
wire wire1287;
wire wire1286;
wire wire473;
wire wire1290;
wire wire1289;
wire wire1292;
wire wire557;
wire wire1294;
wire wire1293;
wire n_n1566;
wire wire88;
wire wire1295;
wire n_n1575;
wire wire1297;
wire wire124;
wire wire1302;
wire wire1305;
wire wire1311;
wire wire80;
wire n_n2859;
wire n_n4657;
wire wire160;
wire wire78;
wire wire651;
wire n_n3570;
wire n_n3573;
wire wire1319;
wire n_n3823;
wire wire1321;
wire wire537;
wire wire1326;
wire n_n5070;
wire wire217;
wire n_n3037;
wire wire469;
wire wire1331;
wire wire115;
wire wire673;
wire n_n3029;
wire wire1336;
wire wire173;
wire n_n2733;
wire wire1341;
wire wire378;
wire wire1345;
wire wire1343;
wire wire1342;
wire wire1347;
wire wire1346;
wire n_n784;
wire wire629;
wire n_n752;
wire wire1354;
wire wire1357;
wire wire244;
wire wire1363;
wire wire1366;
wire wire1367;
wire wire479;
wire wire222;
wire n_n3525;
wire wire1375;
wire n_n3561;
wire n_n3825;
wire wire1378;
wire n_n3180;
wire wire1381;
wire wire1383;
wire n_n3170;
wire wire1386;
wire wire1390;
wire wire1389;
wire wire170;
wire wire1395;
wire wire1401;
wire wire1404;
wire wire1405;
wire wire219;
wire n_n371;
wire wire1416;
wire wire1415;
wire wire1414;
wire wire759;
wire wire1417;
wire wire645;
wire wire664;
wire wire171;
wire wire394;
wire wire1420;
wire n_n3592;
wire n_n3834;
wire n_n3833;
wire wire1425;
wire wire1424;
wire wire1427;
wire wire1432;
wire wire1436;
wire wire1437;
wire n_n772;
wire wire1440;
wire wire1444;
wire n_n326;
wire wire1446;
wire wire86;
wire wire240;
wire wire497;
wire wire1450;
wire wire636;
wire n_n3578;
wire wire47;
wire wire1459;
wire wire1463;
wire n_n2956;
wire wire1465;
wire n_n3601;
wire wire197;
wire wire1470;
wire wire1469;
wire wire401;
wire wire1477;
wire wire1476;
wire wire1480;
wire wire1479;
wire wire1478;
wire wire1483;
wire wire1482;
wire n_n225;
wire n_n5021;
wire wire128;
wire wire565;
wire wire1488;
wire wire579;
wire wire648;
wire wire681;
wire wire1489;
wire wire504;
wire n_n3800;
wire n_n3514;
wire wire1491;
wire n_n3802;
wire n_n3511;
wire wire690;
wire wire1493;
wire wire1496;
wire wire1495;
wire wire1498;
wire wire1497;
wire wire1500;
wire wire1499;
wire wire1503;
wire wire1504;
wire wire1507;
wire wire1510;
wire wire1513;
wire wire1512;
wire wire689;
wire wire1519;
wire wire1520;
wire wire1523;
wire n_n3176;
wire wire1524;
wire wire1527;
wire wire315;
wire wire1537;
wire wire1539;
wire n_n1163;
wire wire348;
wire wire385;
wire wire675;
wire wire1544;
wire wire270;
wire wire1553;
wire wire1556;
wire wire1558;
wire wire1560;
wire wire1562;
wire wire1568;
wire wire1570;
wire wire560;
wire wire688;
wire wire432;
wire wire1576;
wire n_n3555;
wire wire1580;
wire wire1579;
wire wire1578;
wire wire1581;
wire wire1582;
wire wire1587;
wire wire1590;
wire wire1592;
wire wire1595;
wire wire57;
wire wire434;
wire wire538;
wire wire539;
wire wire1601;
wire n_n2777;
wire wire1602;
wire wire607;
wire wire640;
wire wire584;
wire wire1605;
wire wire1613;
wire wire1617;
wire n_n3485;
wire wire698;
wire n_n3467;
wire n_n3510;
wire wire1625;
wire wire578;
wire n_n2754;
wire wire1627;
wire n_n2630;
wire wire642;
wire wire1628;
wire wire407;
wire wire1630;
wire wire1632;
wire n_n765;
wire wire635;
wire wire1633;
wire n_n745;
wire wire346;
wire wire1636;
wire wire1640;
wire wire1639;
wire n_n302;
wire wire1641;
wire n_n301;
wire n_n3473;
wire wire1648;
wire n_n3470;
wire n_n2642;
wire wire1649;
wire wire1655;
wire wire1658;
wire n_n768;
wire wire1659;
wire n_n746;
wire wire697;
wire wire1668;
wire wire1666;
wire n_n304;
wire n_n3501;
wire n_n3500;
wire wire1674;
wire n_n834;
wire wire107;
wire wire1675;
wire n_n769;
wire wire1679;
wire n_n747;
wire wire1684;
wire wire296;
wire wire1689;
wire wire696;
wire n_n3542;
wire n_n3482;
wire n_n3487;
wire n_n3460;
wire wire1695;
wire wire1704;
wire wire1706;
wire wire1709;
wire wire1708;
wire wire1707;
wire n_n748;
wire wire1717;
wire wire1716;
wire wire1720;
wire wire1723;
wire wire606;
wire wire1730;
wire wire1729;
wire n_n2626;
wire wire263;
wire wire1735;
wire wire165;
wire wire1739;
wire wire1738;
wire wire1741;
wire wire1740;
wire wire1743;
wire wire1742;
wire n_n333;
wire wire256;
wire wire1748;
wire wire1747;
wire n_n3492;
wire n_n3491;
wire wire1751;
wire n_n3462;
wire n_n3489;
wire n_n3451;
wire wire1754;
wire wire1753;
wire wire1756;
wire wire1758;
wire wire1761;
wire wire1766;
wire wire1775;
wire wire1779;
wire wire1778;
wire wire1777;
wire wire1780;
wire n_n2684;
wire wire1782;
wire wire1786;
wire n_n1801;
wire wire1789;
wire n_n4419;
wire wire1791;
wire wire1794;
wire n_n4399;
wire wire1807;
wire wire1809;
wire wire225;
wire wire1811;
wire wire1812;
wire wire1814;
wire wire49;
wire wire50;
wire wire54;
wire wire56;
wire wire72;
wire wire75;
wire wire79;
wire wire82;
wire wire84;
wire wire87;
wire wire92;
wire wire94;
wire wire99;
wire wire108;
wire wire110;
wire wire116;
wire wire117;
wire wire120;
wire wire121;
wire wire148;
wire wire161;
wire wire415;
wire wire162;
wire wire438;
wire wire163;
wire wire399;
wire wire164;
wire wire340;
wire wire284;
wire wire166;
wire wire339;
wire wire169;
wire wire174;
wire wire177;
wire wire179;
wire wire183;
wire wire184;
wire wire187;
wire wire425;
wire wire192;
wire wire193;
wire wire424;
wire wire194;
wire wire195;
wire wire358;
wire wire196;
wire wire198;
wire wire199;
wire wire362;
wire wire200;
wire wire366;
wire wire201;
wire wire202;
wire wire203;
wire wire204;
wire wire205;
wire wire206;
wire wire210;
wire wire211;
wire wire215;
wire wire216;
wire wire220;
wire wire221;
wire wire223;
wire wire229;
wire wire230;
wire wire232;
wire wire233;
wire wire235;
wire wire236;
wire wire237;
wire wire238;
wire wire239;
wire wire241;
wire wire242;
wire wire243;
wire wire246;
wire wire251;
wire wire252;
wire wire254;
wire wire258;
wire wire259;
wire wire260;
wire wire261;
wire wire262;
wire wire264;
wire wire265;
wire wire268;
wire wire269;
wire wire271;
wire wire272;
wire wire273;
wire wire274;
wire wire275;
wire wire277;
wire wire278;
wire wire280;
wire wire281;
wire wire282;
wire wire283;
wire wire289;
wire wire290;
wire wire291;
wire wire292;
wire wire293;
wire wire294;
wire wire295;
wire wire297;
wire wire298;
wire wire299;
wire wire300;
wire wire301;
wire wire302;
wire wire303;
wire wire304;
wire wire305;
wire wire306;
wire wire307;
wire wire309;
wire wire310;
wire wire311;
wire wire312;
wire wire314;
wire wire316;
wire wire317;
wire wire318;
wire wire319;
wire wire320;
wire wire321;
wire wire322;
wire wire323;
wire wire324;
wire wire325;
wire wire326;
wire wire327;
wire wire328;
wire wire329;
wire wire330;
wire wire331;
wire wire332;
wire wire333;
wire wire336;
wire wire337;
wire wire338;
wire wire341;
wire wire342;
wire wire345;
wire wire347;
wire wire349;
wire wire351;
wire wire352;
wire wire354;
wire wire357;
wire wire368;
wire wire369;
wire wire370;
wire wire371;
wire wire372;
wire wire373;
wire wire374;
wire wire375;
wire wire380;
wire wire398;
wire wire400;
wire wire402;
wire wire403;
wire wire405;
wire wire406;
wire wire408;
wire wire409;
wire wire410;
wire wire413;
wire wire414;
wire wire416;
wire wire417;
wire wire418;
wire wire1840;
wire wire1844;
wire wire1853;
wire wire1862;
wire wire1864;
wire wire1902;
wire wire795;
wire wire805;
wire wire815;
wire wire890;
wire wire994;
wire wire1128;
wire wire1131;
wire wire1203;
wire wire1209;
wire wire1253;
wire wire1328;
wire wire1356;
wire wire1409;
wire wire1447;
wire wire1522;
wire wire1550;
wire wire1557;
wire wire1619;
wire wire1638;
wire wire1643;
wire wire1661;
wire wire1768;
wire wire1842;
wire wire138;
wire wire439;
wire wire441;
wire wire467;
wire wire499;
wire wire501;
wire wire507;
wire wire508;
wire wire510;
wire wire513;
wire wire516;
wire wire520;
wire wire552;
wire wire556;
wire wire1906;
wire wire1907;
wire wire1908;
wire wire1910;
wire wire1912;
wire wire1914;
wire wire1916;
wire wire1936;
wire wire1937;
wire wire1938;
wire wire1939;
wire wire1940;
wire wire1945;
wire wire1946;
wire wire1949;
wire wire1950;
wire wire1951;
wire wire1960;
wire wire1961;
wire wire1962;
wire wire1968;
wire wire1971;
wire wire1972;
wire wire1976;
wire wire1979;
wire wire1982;
wire wire1983;
wire wire1987;
wire wire1988;
wire wire1990;
wire wire1991;
wire wire1992;
wire wire1993;
wire wire1995;
wire wire1996;
wire wire1997;
wire wire1998;
wire wire1999;
wire wire2000;
wire wire2004;
wire wire2017;
wire wire2026;
wire wire2027;
wire wire2032;
wire wire2035;
wire wire2040;
wire wire2041;
wire wire2045;
wire wire2051;
wire wire2062;
wire wire2068;
wire wire2070;
wire wire2078;
wire wire2079;
wire wire2080;
wire wire2083;
wire wire2099;
wire wire2108;
wire wire2119;
wire wire2124;
wire wire2125;
wire wire2130;
wire wire2134;
wire wire2136;
wire wire2139;
wire wire2141;
wire wire2146;
wire wire2149;
wire wire2153;
wire wire2155;
wire wire2156;
wire wire2157;
wire wire2163;
wire wire2169;
wire wire2172;
wire wire2174;
wire wire2176;
wire wire2177;
wire wire2179;
wire wire2180;
wire wire2181;
wire wire2182;
wire wire2190;
wire wire2191;
wire wire2195;
wire wire2197;
wire wire2204;
wire wire2205;
wire wire2218;
wire wire2229;
wire wire2232;
wire wire2233;
wire wire2239;
wire wire2240;
wire wire2242;
wire wire2243;
wire wire2245;
wire wire2257;
wire wire2269;
wire wire2277;
wire wire2278;
wire wire2281;
wire wire2282;
wire wire2283;
wire wire2287;
wire wire2290;
wire wire2293;
wire wire2294;
wire wire2295;
wire wire2296;
wire wire2302;
wire wire2303;
wire wire2308;
wire wire2310;
wire wire2311;
wire wire2323;
wire wire2324;
wire wire2329;
wire wire2331;
wire wire2335;
wire wire2336;
wire wire2340;
wire wire2341;
wire wire2343;
wire wire2344;
wire wire2345;
wire wire2346;
wire wire2349;
wire wire2350;
wire wire2351;
wire wire2352;
wire wire2353;
wire wire2356;
wire wire2359;
wire wire2362;
wire wire2364;
wire wire2365;
wire wire2370;
wire wire2371;
wire wire2372;
wire wire2373;
wire wire2374;
wire wire2375;
wire wire2379;
wire wire2380;
wire wire2382;
wire wire2384;
wire wire2393;
wire wire2398;
wire wire2404;
wire wire2405;
wire wire2407;
wire wire2410;
wire wire2415;
wire wire2417;
wire wire2418;
wire wire2424;
wire wire2427;
wire wire2428;
wire wire2435;
wire wire2442;
wire wire2448;
wire wire2449;
wire wire2451;
wire wire2452;
wire wire2462;
wire wire2463;
wire wire2464;
wire wire2468;
wire wire2475;
wire wire2480;
wire wire2481;
wire wire2487;
wire wire2488;
wire wire2489;
wire wire2490;
wire wire2493;
wire wire2498;
wire wire2513;
wire wire2516;
wire wire2518;
wire wire2522;
wire wire2523;
wire wire2524;
wire wire2525;
wire wire2526;
wire wire2532;
wire wire2537;
wire wire2540;
wire wire2543;
wire wire2545;
wire wire2548;
wire wire2549;
wire wire2556;
wire wire2557;
wire wire2558;
wire wire2559;
wire wire2560;
wire wire2565;
wire wire2567;
wire wire2568;
wire wire2576;
wire wire2578;
wire wire2579;
wire wire2584;
wire wire2585;
wire wire2588;
wire wire2594;
wire wire2595;
wire wire2598;
wire wire2599;
wire wire2606;
wire wire2610;
wire wire2614;
wire wire2615;
wire wire2618;
wire wire2630;
wire wire2631;
wire wire2634;
wire wire2635;
wire wire2636;
wire wire2638;
wire wire2643;
wire wire2645;
wire wire2646;
wire wire2657;
wire wire2666;
wire wire2669;
wire wire2676;
wire wire2679;
wire wire2686;
wire wire2691;
wire wire2692;
wire wire2693;
wire wire2700;
wire wire2702;
wire wire2703;
wire wire2704;
wire wire2705;
wire wire2712;
wire wire2713;
wire wire2717;
wire wire2718;
wire wire2720;
wire wire2721;
wire wire2724;
wire wire2726;
wire wire2728;
wire wire2729;
wire wire2730;
wire wire2731;
wire wire2733;
wire wire2738;
wire wire2739;
wire wire2740;
wire wire2741;
wire wire2743;
wire wire2744;
wire wire2746;
wire wire2748;
wire wire2750;
wire wire2751;
wire wire2775;
wire wire2776;
wire wire2784;
wire wire2785;
wire wire2791;
wire wire2797;
wire wire2801;
wire wire2802;
wire wire2808;
wire wire2809;
wire wire2814;
wire wire2815;
wire wire2817;
wire wire2825;
wire wire2828;
wire wire2831;
wire wire2842;
wire wire2843;
wire wire2848;
wire wire2849;
wire wire2850;
wire wire2851;
wire wire2853;
wire wire2861;
wire wire2865;
wire wire2866;
wire wire2870;
wire wire2875;
wire wire2896;
wire wire2897;
wire wire2900;
wire wire2901;
wire wire2909;
wire wire2910;
wire wire2911;
wire wire2914;
wire wire2915;
wire wire2923;
wire wire2937;
wire wire2939;
wire wire2940;
wire wire2943;
wire wire2944;
wire wire2952;
wire wire2953;
wire wire2958;
wire wire2959;
wire wire2962;
wire wire2964;
wire wire2965;
wire wire2970;
wire wire2974;
wire wire2975;
wire wire2977;
wire wire2979;
wire wire2981;
wire wire2985;
wire wire2995;
wire wire3001;
wire wire3006;
wire wire3008;
wire wire3013;
wire wire3014;
wire wire3015;
wire wire3020;
wire wire3027;
wire wire3032;
wire wire3044;
wire wire3059;
wire wire3060;
wire wire3066;
wire wire3067;
wire wire3068;
wire wire3069;
wire wire3078;
wire wire3079;
wire wire3080;
wire wire3081;
wire wire3093;
wire wire3098;
wire wire3102;
wire wire3111;
wire wire3113;
wire wire3118;
wire wire3123;
wire wire3124;
wire wire3128;
wire wire3135;
wire wire3136;
wire wire3142;
wire wire3143;
wire wire3154;
wire wire3155;
wire wire3177;
wire wire3194;
wire wire3195;
wire wire3201;
wire wire3202;
wire wire3209;
wire wire3210;
wire wire3217;
wire wire3219;
wire wire3220;
wire wire3222;
wire wire3223;
wire wire3224;
wire wire3225;
wire wire3229;
wire wire3230;
wire wire3232;
wire wire3233;
wire wire3234;
wire wire3244;
wire wire3245;
wire wire3248;
wire wire3256;
wire wire3257;
wire wire3258;
wire wire3264;
wire wire3271;
wire wire3275;
wire wire3279;
wire wire3280;
wire wire3291;
wire wire3292;
wire wire3296;
wire wire3298;
wire wire3299;
wire wire3300;
wire wire3301;
wire wire3308;
wire wire3312;
wire wire3313;
wire wire3325;
wire wire3328;
wire wire3333;
wire wire3337;
wire wire3338;
wire wire3342;
wire wire3343;
wire wire3349;
wire wire3353;
wire wire3374;
wire wire3375;
wire wire3376;
wire wire3385;
wire wire3392;
wire wire3396;
wire wire3397;
wire wire3403;
wire wire3404;
wire wire3409;
wire wire3410;
wire wire3415;
wire wire3425;
wire wire3433;
wire wire3434;
wire wire3435;
wire wire3437;
wire wire3438;
wire wire3439;
wire wire3442;
wire wire3451;
wire wire3461;
wire wire3469;
wire wire3470;
wire wire3471;
wire wire3472;
wire wire3479;
wire wire3480;
wire wire3484;
wire wire3496;
wire wire3497;
wire wire3498;
wire wire3515;
wire wire3516;
wire wire3520;
wire wire3524;
wire wire3526;
wire wire3527;
wire wire3531;
wire wire3533;
wire wire3545;
wire wire3550;
wire wire3551;
wire wire3563;
wire wire3570;
wire wire3575;
wire wire3580;
wire wire3581;
wire wire3588;
wire wire3594;
wire wire3601;
wire wire3607;
wire wire3621;
wire wire3622;
wire wire3624;
wire wire3628;
wire wire3629;
wire wire3643;
wire wire3653;
wire wire3658;
wire wire3662;
wire wire3665;
wire wire3671;
wire wire3676;
wire wire3685;
wire wire3690;
wire wire3696;
wire wire3700;
wire wire3701;
wire wire3702;
wire wire3710;
wire wire3723;
wire wire3747;
wire wire3755;
wire wire3759;
wire wire3767;
wire wire3773;
wire wire3774;
wire wire3810;
wire wire3811;
wire wire3820;
wire wire3828;
wire wire3829;
wire wire3835;
wire wire3836;
wire wire3850;
wire wire3851;
wire wire3866;
wire wire3885;
wire wire3886;
wire wire3887;
wire wire3895;
wire wire3896;
wire wire3897;
wire wire3899;
wire wire3900;
wire wire3901;
wire wire3957;
wire wire3958;
wire wire3964;
wire wire3973;
wire wire3985;
wire wire3990;
wire wire3991;
wire wire3996;
wire wire3997;
wire wire3998;
wire wire4013;
wire wire4020;
wire wire4021;
wire wire4026;
wire wire4027;
wire wire4043;
wire wire4048;
wire wire4060;
wire wire4064;
wire wire4065;
wire wire4067;
wire wire4080;
wire wire4088;
wire wire4102;
wire wire4103;
wire wire4104;
wire wire4113;
wire wire4126;
wire wire4130;
wire wire4143;
wire wire4151;
wire wire4158;
wire wire4159;
wire wire4172;
wire wire4182;
wire wire4185;
wire wire4186;
wire wire4217;
wire wire4220;
wire wire4221;
wire wire4223;
wire wire4228;
wire wire4229;
wire wire4230;
wire wire4233;
wire wire4234;
wire wire4252;
wire wire4253;
wire wire4260;
wire wire4263;
wire wire4285;
wire wire4286;
wire wire4291;
wire wire4320;
wire wire4323;
wire wire4324;
wire wire4334;
wire wire4341;
wire wire4343;
wire wire4344;
wire wire4354;
wire wire4355;
wire wire4365;
wire wire4372;
wire wire4376;
wire wire4382;
wire wire4393;
wire wire4395;
wire wire4396;
wire wire4419;
wire wire4420;
wire wire4427;
wire wire4428;
wire wire4429;
wire wire4430;
wire wire4434;
wire wire4453;
wire wire4454;
wire wire4458;
wire wire4459;
wire wire4460;
wire wire4470;
wire wire4474;
wire wire4475;
wire wire4481;
wire wire4485;
wire wire4486;
wire wire4491;
wire wire4496;
wire wire4500;
wire wire4503;
wire wire4504;
wire wire4505;
wire wire4506;
wire wire4508;
wire wire4509;
wire wire4510;
wire wire4520;
wire wire4523;
wire wire4526;
wire wire4531;
wire wire4539;
wire wire4544;
wire wire4545;
wire wire4548;
wire wire4549;
wire wire4550;
wire wire4551;
wire wire4554;
wire wire4558;
wire wire4561;
wire wire4562;
wire wire4568;
wire wire4569;
wire wire4572;
wire wire4573;
wire wire4576;
wire wire4581;
wire wire4591;
wire wire4602;
wire wire4619;
wire wire4620;
wire wire4628;
wire wire4638;
wire wire4639;
wire wire4643;
wire wire4644;
wire wire4649;
wire wire4651;
wire wire4655;
wire wire4658;
wire wire4659;
wire wire4662;
wire wire4663;
wire wire4669;
wire wire4671;
wire wire4676;
wire wire4680;
wire wire4684;
wire wire4685;
wire wire4701;
wire wire4735;
wire wire4739;
wire wire4740;
wire wire4743;
wire wire4750;
wire wire4751;
wire wire4752;
wire wire4753;
wire wire4765;
wire wire4768;
wire wire4771;
wire wire4780;
wire wire4786;
wire wire4805;
wire wire4818;
wire wire4819;
wire wire4820;
wire wire4821;
wire wire4822;
wire wire4827;
wire wire4828;
wire wire4829;
wire wire4830;
wire wire4831;
wire wire4832;
wire wire4838;
wire wire4839;
wire wire4842;
wire wire4857;
wire wire4858;
wire wire4859;
wire wire4860;
wire wire4863;
wire wire4864;
wire wire4869;
wire wire4870;
wire wire4888;
wire wire4890;
wire wire4891;
wire wire4900;
wire wire4904;
wire wire4905;
wire wire4908;
wire wire4919;
wire wire4924;
wire wire4933;
wire wire4934;
wire wire4935;
wire wire4937;
wire wire4941;
wire wire4942;
wire wire4948;
wire wire4950;
wire wire4953;
wire wire4960;
wire wire4961;
wire wire4965;
wire wire4966;
wire wire4974;
wire wire4981;
wire wire4982;
wire wire4986;
wire wire4993;
wire wire4998;
wire wire5022;
wire wire5023;
wire wire5024;
wire wire5025;
wire wire5026;
wire wire5027;
wire wire5032;
wire wire5057;
wire wire5067;
wire wire5068;
wire wire16857;
wire wire16861;
wire wire16863;
wire wire16865;
wire wire16866;
wire wire16867;
wire wire16870;
wire wire16871;
wire wire16872;
wire wire16876;
wire wire16877;
wire wire16880;
wire wire16884;
wire wire16885;
wire wire16886;
wire wire16888;
wire wire16889;
wire wire16890;
wire wire16892;
wire wire16896;
wire wire16897;
wire wire16898;
wire wire16908;
wire wire16909;
wire wire16910;
wire wire16911;
wire wire16924;
wire wire16929;
wire wire16930;
wire wire16933;
wire wire16936;
wire wire16940;
wire wire16941;
wire wire16943;
wire wire16946;
wire wire16950;
wire wire16952;
wire wire16953;
wire wire16954;
wire wire16957;
wire wire16960;
wire wire16961;
wire wire16962;
wire wire16964;
wire wire16966;
wire wire16968;
wire wire16972;
wire wire16974;
wire wire16975;
wire wire16976;
wire wire16980;
wire wire16987;
wire wire16988;
wire wire16990;
wire wire16991;
wire wire16993;
wire wire16994;
wire wire16995;
wire wire16996;
wire wire16997;
wire wire17000;
wire wire17001;
wire wire17003;
wire wire17007;
wire wire17013;
wire wire17014;
wire wire17016;
wire wire17018;
wire wire17019;
wire wire17023;
wire wire17025;
wire wire17028;
wire wire17033;
wire wire17034;
wire wire17035;
wire wire17038;
wire wire17039;
wire wire17041;
wire wire17042;
wire wire17044;
wire wire17045;
wire wire17047;
wire wire17049;
wire wire17050;
wire wire17052;
wire wire17053;
wire wire17055;
wire wire17056;
wire wire17058;
wire wire17060;
wire wire17061;
wire wire17063;
wire wire17064;
wire wire17067;
wire wire17070;
wire wire17071;
wire wire17072;
wire wire17074;
wire wire17076;
wire wire17079;
wire wire17081;
wire wire17082;
wire wire17083;
wire wire17089;
wire wire17093;
wire wire17094;
wire wire17096;
wire wire17100;
wire wire17102;
wire wire17106;
wire wire17108;
wire wire17109;
wire wire17114;
wire wire17115;
wire wire17116;
wire wire17117;
wire wire17119;
wire wire17120;
wire wire17121;
wire wire17122;
wire wire17123;
wire wire17125;
wire wire17127;
wire wire17128;
wire wire17129;
wire wire17132;
wire wire17134;
wire wire17136;
wire wire17137;
wire wire17139;
wire wire17140;
wire wire17141;
wire wire17145;
wire wire17146;
wire wire17149;
wire wire17150;
wire wire17152;
wire wire17153;
wire wire17154;
wire wire17156;
wire wire17158;
wire wire17159;
wire wire17164;
wire wire17166;
wire wire17169;
wire wire17170;
wire wire17172;
wire wire17174;
wire wire17175;
wire wire17176;
wire wire17178;
wire wire17181;
wire wire17184;
wire wire17185;
wire wire17186;
wire wire17187;
wire wire17190;
wire wire17191;
wire wire17193;
wire wire17196;
wire wire17198;
wire wire17201;
wire wire17202;
wire wire17203;
wire wire17206;
wire wire17209;
wire wire17212;
wire wire17213;
wire wire17215;
wire wire17217;
wire wire17220;
wire wire17224;
wire wire17226;
wire wire17228;
wire wire17229;
wire wire17231;
wire wire17234;
wire wire17238;
wire wire17239;
wire wire17241;
wire wire17243;
wire wire17245;
wire wire17246;
wire wire17247;
wire wire17249;
wire wire17251;
wire wire17253;
wire wire17256;
wire wire17257;
wire wire17258;
wire wire17259;
wire wire17260;
wire wire17265;
wire wire17266;
wire wire17268;
wire wire17271;
wire wire17272;
wire wire17275;
wire wire17276;
wire wire17277;
wire wire17280;
wire wire17281;
wire wire17284;
wire wire17285;
wire wire17287;
wire wire17288;
wire wire17289;
wire wire17290;
wire wire17291;
wire wire17292;
wire wire17294;
wire wire17295;
wire wire17297;
wire wire17298;
wire wire17299;
wire wire17301;
wire wire17303;
wire wire17305;
wire wire17307;
wire wire17309;
wire wire17310;
wire wire17313;
wire wire17314;
wire wire17317;
wire wire17319;
wire wire17321;
wire wire17322;
wire wire17324;
wire wire17325;
wire wire17327;
wire wire17329;
wire wire17333;
wire wire17335;
wire wire17336;
wire wire17337;
wire wire17338;
wire wire17339;
wire wire17341;
wire wire17342;
wire wire17343;
wire wire17345;
wire wire17347;
wire wire17349;
wire wire17350;
wire wire17352;
wire wire17353;
wire wire17357;
wire wire17358;
wire wire17359;
wire wire17360;
wire wire17361;
wire wire17363;
wire wire17364;
wire wire17365;
wire wire17367;
wire wire17368;
wire wire17374;
wire wire17377;
wire wire17379;
wire wire17382;
wire wire17383;
wire wire17384;
wire wire17385;
wire wire17388;
wire wire17389;
wire wire17390;
wire wire17391;
wire wire17392;
wire wire17393;
wire wire17394;
wire wire17395;
wire wire17397;
wire wire17398;
wire wire17400;
wire wire17401;
wire wire17405;
wire wire17407;
wire wire17408;
wire wire17410;
wire wire17416;
wire wire17417;
wire wire17418;
wire wire17420;
wire wire17426;
wire wire17428;
wire wire17431;
wire wire17433;
wire wire17434;
wire wire17435;
wire wire17436;
wire wire17438;
wire wire17439;
wire wire17440;
wire wire17441;
wire wire17443;
wire wire17445;
wire wire17446;
wire wire17447;
wire wire17448;
wire wire17450;
wire wire17452;
wire wire17453;
wire wire17454;
wire wire17456;
wire wire17457;
wire wire17458;
wire wire17459;
wire wire17462;
wire wire17465;
wire wire17466;
wire wire17467;
wire wire17468;
wire wire17469;
wire wire17470;
wire wire17471;
wire wire17472;
wire wire17478;
wire wire17479;
wire wire17480;
wire wire17483;
wire wire17484;
wire wire17486;
wire wire17490;
wire wire17493;
wire wire17498;
wire wire17499;
wire wire17501;
wire wire17504;
wire wire17505;
wire wire17507;
wire wire17509;
wire wire17510;
wire wire17513;
wire wire17514;
wire wire17516;
wire wire17518;
wire wire17521;
wire wire17522;
wire wire17528;
wire wire17529;
wire wire17533;
wire wire17534;
wire wire17535;
wire wire17537;
wire wire17539;
wire wire17541;
wire wire17542;
wire wire17543;
wire wire17545;
wire wire17548;
wire wire17549;
wire wire17550;
wire wire17552;
wire wire17553;
wire wire17554;
wire wire17555;
wire wire17557;
wire wire17558;
wire wire17559;
wire wire17560;
wire wire17562;
wire wire17563;
wire wire17565;
wire wire17566;
wire wire17568;
wire wire17569;
wire wire17570;
wire wire17573;
wire wire17574;
wire wire17575;
wire wire17576;
wire wire17578;
wire wire17579;
wire wire17581;
wire wire17582;
wire wire17585;
wire wire17586;
wire wire17587;
wire wire17588;
wire wire17591;
wire wire17592;
wire wire17593;
wire wire17594;
wire wire17596;
wire wire17599;
wire wire17600;
wire wire17601;
wire wire17602;
wire wire17604;
wire wire17605;
wire wire17606;
wire wire17608;
wire wire17610;
wire wire17612;
wire wire17615;
wire wire17622;
wire wire17626;
wire wire17627;
wire wire17629;
wire wire17631;
wire wire17632;
wire wire17635;
wire wire17638;
wire wire17639;
wire wire17640;
wire wire17646;
wire wire17647;
wire wire17650;
wire wire17651;
wire wire17654;
wire wire17656;
wire wire17657;
wire wire17659;
wire wire17660;
wire wire17662;
wire wire17663;
wire wire17667;
wire wire17668;
wire wire17671;
wire wire17672;
wire wire17674;
wire wire17676;
wire wire17677;
wire wire17679;
wire wire17681;
wire wire17682;
wire wire17684;
wire wire17685;
wire wire17686;
wire wire17688;
wire wire17690;
wire wire17691;
wire wire17692;
wire wire17693;
wire wire17695;
wire wire17696;
wire wire17697;
wire wire17698;
wire wire17700;
wire wire17701;
wire wire17704;
wire wire17705;
wire wire17706;
wire wire17708;
wire wire17709;
wire wire17710;
wire wire17712;
wire wire17716;
wire wire17717;
wire wire17721;
wire wire17724;
wire wire17725;
wire wire17726;
wire wire17729;
wire wire17732;
wire wire17735;
wire wire17739;
wire wire17740;
wire wire17741;
wire wire17744;
wire wire17746;
wire wire17747;
wire wire17748;
wire wire17750;
wire wire17752;
wire wire17753;
wire wire17756;
wire wire17757;
wire wire17760;
wire wire17761;
wire wire17764;
wire wire17765;
wire wire17766;
wire wire17767;
wire wire17772;
wire wire17773;
wire wire17776;
wire wire17778;
wire wire17779;
wire wire17781;
wire wire17783;
wire wire17786;
wire wire17787;
wire wire17793;
wire wire17796;
wire wire17798;
wire wire17800;
wire wire17801;
wire wire17805;
wire wire17806;
wire wire17808;
wire wire17810;
wire wire17812;
wire wire17813;
wire wire17816;
wire wire17817;
wire wire17818;
wire wire17819;
wire wire17821;
wire wire17822;
wire wire17824;
wire wire17825;
wire wire17826;
wire wire17827;
wire wire17830;
wire wire17831;
wire wire17832;
wire wire17836;
wire wire17837;
wire wire17839;
wire wire17840;
wire wire17841;
wire wire17842;
wire wire17843;
wire wire17844;
wire wire17845;
wire wire17848;
wire wire17849;
wire wire17850;
wire wire17852;
wire wire17853;
wire wire17854;
wire wire17858;
wire wire17860;
wire wire17861;
wire wire17862;
wire wire17864;
wire wire17865;
wire wire17867;
wire wire17868;
wire wire17869;
wire wire17870;
wire wire17872;
wire wire17873;
wire wire17876;
wire wire17877;
wire wire17880;
wire wire17881;
wire wire17884;
wire wire17887;
wire wire17889;
wire wire17891;
wire wire17893;
wire wire17894;
wire wire17896;
wire wire17897;
wire wire17898;
wire wire17901;
wire wire17903;
wire wire17906;
wire wire17908;
wire wire17909;
wire wire17911;
wire wire17913;
wire wire17915;
wire wire17916;
wire wire17918;
wire wire17919;
wire wire17920;
wire wire17921;
wire wire17924;
wire wire17926;
wire wire17931;
wire wire17934;
wire wire17935;
wire wire17940;
wire wire17941;
wire wire17942;
wire wire17944;
wire wire17947;
wire wire17948;
wire wire17951;
wire wire17952;
wire wire17954;
wire wire17955;
wire wire17958;
wire wire17959;
wire wire17960;
wire wire17963;
wire wire17964;
wire wire17965;
wire wire17968;
wire wire17970;
wire wire17971;
wire wire17972;
wire wire17976;
wire wire17977;
wire wire17979;
wire wire17980;
wire wire17985;
wire wire17987;
wire wire17988;
wire wire17989;
wire wire17993;
wire wire17995;
wire wire17996;
wire wire17999;
wire wire18000;
wire wire18001;
wire wire18002;
wire wire18003;
wire wire18004;
wire wire18007;
wire wire18010;
wire wire18012;
wire wire18013;
wire wire18014;
wire wire18017;
wire wire18018;
wire wire18019;
wire wire18021;
wire wire18023;
wire wire18024;
wire wire18026;
wire wire18027;
wire wire18028;
wire wire18032;
wire wire18035;
wire wire18036;
wire wire18039;
wire wire18044;
wire wire18049;
wire wire18050;
wire wire18051;
wire wire18053;
wire wire18057;
wire wire18058;
wire wire18063;
wire wire18064;
wire wire18067;
wire wire18068;
wire wire18069;
wire wire18071;
wire wire18074;
wire wire18075;
wire wire18076;
wire wire18078;
wire wire18081;
wire wire18082;
wire wire18083;
wire wire18085;
wire wire18087;
wire wire18088;
wire wire18089;
wire wire18091;
wire wire18092;
wire wire18096;
wire wire18097;
wire wire18098;
wire wire18102;
wire wire18103;
wire wire18104;
wire wire18106;
wire wire18107;
wire wire18111;
wire wire18113;
wire wire18117;
wire wire18119;
wire wire18120;
wire wire18122;
wire wire18125;
wire wire18128;
wire wire18129;
wire wire18132;
wire wire18134;
wire wire18135;
wire wire18136;
wire wire18137;
wire wire18140;
wire wire18141;
wire wire18142;
wire wire18144;
wire wire18145;
wire wire18146;
wire wire18148;
wire wire18150;
wire wire18154;
wire wire18155;
wire wire18157;
wire wire18158;
wire wire18159;
wire wire18160;
wire wire18161;
wire wire18163;
wire wire18164;
wire wire18167;
wire wire18168;
wire wire18169;
wire wire18172;
wire wire18173;
wire wire18174;
wire wire18178;
wire wire18180;
wire wire18182;
wire wire18184;
wire wire18185;
wire wire18186;
wire wire18187;
wire wire18188;
wire wire18190;
wire wire18191;
wire wire18192;
wire wire18193;
wire wire18194;
wire wire18196;
wire wire18198;
wire wire18199;
wire wire18200;
wire wire18201;
wire wire18202;
wire wire18205;
wire wire18206;
wire wire18209;
wire wire18210;
wire wire18212;
wire wire18213;
wire wire18214;
wire wire18215;
wire wire18220;
wire wire18221;
wire wire18222;
wire wire18225;
wire wire18230;
wire wire18232;
wire wire18234;
wire wire18237;
wire wire18238;
wire wire18242;
wire wire18243;
wire wire18244;
wire wire18245;
wire wire18251;
wire wire18252;
wire wire18253;
wire wire18260;
wire wire18264;
wire wire18266;
wire wire18267;
wire wire18268;
wire wire18269;
wire wire18270;
wire wire18272;
wire wire18273;
wire wire18278;
wire wire18281;
wire wire18283;
wire wire18287;
wire wire18288;
wire wire18290;
wire wire18292;
wire wire18294;
wire wire18295;
wire wire18297;
wire wire18298;
wire wire18299;
wire wire18300;
wire wire18301;
wire wire18302;
wire wire18307;
wire wire18310;
wire wire18311;
wire wire18316;
wire wire18318;
wire wire18321;
wire wire18323;
wire wire18324;
wire wire18325;
wire wire18328;
wire wire18329;
wire wire18330;
wire wire18332;
wire wire18334;
wire wire18337;
wire wire18342;
wire wire18345;
wire wire18348;
wire wire18352;
wire wire18353;
wire wire18354;
wire wire18355;
wire wire18358;
wire wire18360;
wire wire18361;
wire wire18367;
wire wire18370;
wire wire18371;
wire wire18372;
wire wire18374;
wire wire18375;
wire wire18377;
wire wire18384;
wire wire18385;
wire wire18386;
wire wire18388;
wire wire18391;
wire wire18393;
wire wire18394;
wire wire18397;
wire wire18398;
wire wire18401;
wire wire18402;
wire wire18403;
wire wire18408;
wire wire18409;
wire wire18411;
wire wire18413;
wire wire18414;
wire wire18416;
wire wire18418;
wire wire18420;
wire wire18421;
wire wire18422;
wire wire18424;
wire wire18425;
wire wire18426;
wire wire18429;
wire wire18432;
wire wire18433;
wire wire18434;
wire wire18436;
wire wire18437;
wire wire18444;
wire wire18445;
wire wire18450;
wire wire18452;
wire wire18454;
wire wire18455;
wire wire18457;
wire wire18461;
wire wire18462;
wire wire18467;
wire wire18469;
wire wire18471;
wire wire18474;
wire wire18475;
wire wire18476;
wire wire18481;
wire wire18482;
wire wire18486;
wire wire18487;
wire wire18488;
wire wire18490;
wire wire18492;
wire wire18493;
wire wire18495;
wire wire18496;
wire wire18498;
wire wire18499;
wire wire18504;
wire wire18505;
wire wire18507;
wire wire18508;
wire wire18509;
wire wire18510;
wire wire18512;
wire wire18517;
wire wire18521;
wire wire18522;
wire wire18526;
wire wire18527;
wire wire18528;
wire wire18529;
wire wire18533;
wire wire18534;
wire wire18537;
wire wire18540;
wire wire18541;
wire wire18546;
wire wire18547;
wire wire18548;
wire wire18553;
wire wire18555;
wire wire18559;
wire wire18560;
wire wire18562;
wire wire18564;
wire wire18565;
wire wire18567;
wire wire18568;
wire wire18572;
wire wire18575;
wire wire18576;
wire wire18577;
wire wire18578;
wire wire18581;
wire wire18582;
wire wire18583;
wire wire18586;
wire wire18587;
wire wire18588;
wire wire18593;
wire wire18594;
wire wire18596;
wire wire18598;
wire wire18600;
wire wire18602;
wire wire18603;
wire wire18605;
wire wire18607;
wire wire18608;
wire wire18609;
wire wire18611;
wire wire18614;
wire wire18616;
wire wire18617;
wire wire18619;
wire wire18621;
wire wire18623;
wire wire18624;
wire wire18625;
wire wire18626;
wire wire18631;
wire wire18632;
wire wire18635;
wire wire18637;
wire wire18638;
wire wire18641;
wire wire18642;
wire wire18644;
wire wire18645;
wire wire18646;
wire wire18649;
wire wire18650;
wire wire18652;
wire wire18653;
wire wire18655;
wire wire18656;
wire wire18657;
wire wire18662;
wire wire18663;
wire wire18665;
wire wire18668;
wire wire18669;
wire wire18670;
wire wire18671;
wire wire18676;
wire wire18677;
wire wire18679;
wire wire18680;
wire wire18682;
wire wire18683;
wire wire18685;
wire wire18686;
wire wire18687;
wire wire18688;
wire wire18691;
wire wire18692;
wire wire18694;
wire wire18695;
wire wire18696;
wire wire18701;
wire wire18702;
wire wire18703;
wire wire18704;
wire wire18705;
wire wire18706;
wire wire18707;
wire wire18709;
wire wire18711;
wire wire18712;
wire wire18714;
wire wire18715;
wire wire18718;
wire wire18719;
wire wire18720;
wire wire18725;
wire wire18726;
wire wire18731;
wire wire18732;
wire wire18735;
wire wire18736;
wire wire18737;
wire wire18738;
wire wire18744;
wire wire18749;
wire wire18750;
wire wire18752;
wire wire18755;
wire wire18756;
wire wire18757;
wire wire18760;
wire wire18761;
wire wire18763;
wire wire18767;
wire wire18768;
wire wire18769;
wire wire18770;
wire wire18771;
wire wire18773;
wire wire18776;
wire wire18777;
wire wire18780;
wire wire18783;
wire wire18784;
wire wire18786;
wire wire18788;
wire wire18789;
wire wire18790;
wire wire18792;
wire wire18793;
wire wire18795;
wire wire18801;
wire wire18802;
wire wire18803;
wire wire18804;
wire wire18807;
wire wire18809;
wire wire18810;
wire wire18811;
wire wire18812;
wire wire18814;
wire wire18815;
wire wire18816;
wire wire18818;
wire wire18821;
wire wire18824;
wire wire18826;
wire wire18828;
wire wire18830;
wire wire18831;
wire wire18832;
wire wire18833;
wire wire18834;
wire wire18835;
wire wire18837;
wire wire18838;
wire wire18839;
wire wire18841;
wire wire18845;
wire wire18846;
wire wire18847;
wire wire18850;
wire wire18852;
wire wire18854;
wire wire18855;
wire wire18857;
wire wire18858;
wire wire18859;
wire wire18863;
wire wire18865;
wire wire18866;
wire wire18871;
wire wire18872;
wire wire18874;
wire wire18877;
wire wire18878;
wire wire18879;
wire wire18882;
wire wire18883;
wire wire18884;
wire wire18885;
wire wire18889;
wire wire18890;
wire wire18891;
wire wire18892;
wire wire18894;
wire wire18895;
wire wire18897;
wire wire18898;
wire wire18901;
wire wire18908;
wire wire18911;
wire wire18912;
wire wire18913;
wire wire18914;
wire wire18916;
wire wire18917;
wire wire18918;
wire wire18919;
wire wire18921;
wire wire18922;
wire wire18923;
wire wire18924;
wire wire18925;
wire wire18926;
wire wire18928;
wire wire18929;
wire wire18930;
wire wire18931;
wire wire18932;
wire wire18934;
wire wire18935;
wire wire18936;
wire wire18938;
wire wire18939;
wire wire18941;
wire wire18943;
wire wire18944;
wire wire18945;
wire wire18947;
wire wire18949;
wire wire18950;
wire wire18951;
wire wire18955;
wire wire18956;
wire wire18958;
wire wire18959;
wire wire18961;
wire wire18962;
wire wire18965;
wire wire18966;
wire wire18968;
wire wire18969;
wire wire18970;
wire wire18971;
wire wire18972;
wire wire18973;
wire wire18975;
wire wire18976;
wire wire18978;
wire wire18980;
wire wire18981;
wire wire18985;
wire wire18986;
wire wire18991;
wire wire18992;
wire wire18993;
wire wire18997;
wire wire18998;
wire wire19001;
wire wire19003;
wire wire19004;
wire wire19005;
wire wire19006;
wire wire19008;
wire wire19009;
wire wire19010;
wire wire19011;
wire wire19013;
wire wire19015;
wire wire19016;
wire wire19020;
wire wire19021;
wire wire19023;
wire wire19025;
wire wire19027;
wire wire19029;
wire wire19030;
wire wire19031;
wire wire19033;
wire wire19034;
wire wire19036;
wire wire19038;
wire wire19043;
wire wire19044;
wire wire19047;
wire wire19048;
wire wire19050;
wire wire19053;
wire wire19054;
wire wire19055;
wire wire19057;
wire wire19062;
wire wire19063;
wire wire19069;
wire wire19071;
wire wire19072;
wire wire19074;
wire wire19075;
wire wire19076;
wire wire19077;
wire wire19078;
wire wire19079;
wire wire19083;
wire wire19084;
wire wire19087;
wire wire19089;
wire wire19090;
wire wire19094;
wire wire19097;
wire wire19098;
wire wire19099;
wire wire19103;
wire wire19104;
wire wire19106;
wire wire19108;
wire wire19109;
wire wire19110;
wire wire19113;
wire wire19116;
wire wire19118;
wire wire19119;
wire wire19123;
wire wire19125;
wire wire19126;
wire wire19127;
wire wire19128;
wire wire19129;
wire wire19130;
wire wire19134;
wire wire19138;
wire wire19144;
wire wire19146;
wire wire19147;
wire wire19148;
wire wire19150;
wire wire19152;
wire wire19153;
wire wire19158;
wire wire19163;
wire wire19164;
wire wire19168;
wire wire19169;
wire wire19170;
wire wire19174;
wire wire19177;
wire wire19178;
wire wire19179;
wire wire19182;
wire wire19185;
wire wire19186;
wire wire19189;
wire wire19190;
wire wire19192;
wire wire19193;
wire wire19194;
wire wire19196;
wire wire19197;
wire wire19200;
wire wire19201;
wire wire19202;
wire wire19204;
wire wire19208;
wire wire19210;
wire wire19211;
wire wire19212;
wire wire19213;
wire wire19216;
wire wire19219;
wire wire19220;
wire wire19221;
wire wire19226;
wire wire19227;
wire wire19232;
wire wire19233;
wire wire19234;
wire wire19238;
wire wire19239;
wire wire19240;
wire wire19241;
wire wire19243;
wire wire19245;
wire wire19246;
wire wire19248;
wire wire19249;
wire wire19250;
wire wire19253;
wire wire19256;
wire wire19258;
wire wire19259;
wire wire19260;
wire wire19263;
wire wire19268;
wire wire19269;
wire wire19270;
wire wire19272;
wire wire19273;
wire wire19274;
wire wire19276;
wire wire19277;
wire wire19278;
wire wire19279;
wire wire19281;
wire wire19283;
wire wire19284;
wire wire19285;
wire wire19286;
wire wire19289;
wire wire19290;
wire wire19291;
wire wire19294;
wire wire19295;
wire wire19297;
wire wire19299;
wire wire19301;
wire wire19302;
wire wire19304;
wire wire19306;
wire wire19307;
wire wire19308;
wire wire19309;
wire wire19310;
wire wire19312;
wire wire19315;
wire wire19316;
wire wire19317;
wire wire19318;
wire wire19320;
wire wire19324;
wire wire19325;
wire wire19326;
wire wire19328;
wire wire19332;
wire wire19337;
wire wire19338;
wire wire19339;
wire wire19343;
wire wire19344;
wire wire19346;
wire wire19347;
wire wire19348;
wire wire19349;
wire wire19351;
wire wire19354;
wire wire19355;
wire wire19359;
wire wire19362;
wire wire19363;
wire wire19364;
wire wire19366;
wire wire19368;
wire wire19369;
wire wire19370;
wire wire19375;
wire wire19376;
wire wire19380;
wire wire19381;
wire wire19387;
wire wire19388;
wire wire19389;
wire wire19393;
wire wire19395;
wire wire19396;
wire wire19400;
wire wire19401;
wire wire19402;
wire wire19403;
wire wire19405;
wire wire19406;
wire wire19408;
wire wire19409;
wire wire19411;
wire wire19412;
wire wire19413;
wire wire19414;
wire wire19417;
wire wire19420;
wire wire19423;
wire wire19424;
wire wire19426;
wire wire19427;
wire wire19429;
wire wire19430;
wire wire19431;
wire wire19436;
wire wire19437;
wire wire19438;
wire wire19440;
wire wire19441;
wire wire19442;
wire wire19443;
wire wire19446;
wire wire19447;
wire wire19448;
wire wire19449;
wire wire19450;
wire wire19452;
wire wire19453;
wire wire19454;
wire wire19455;
wire wire19456;
wire wire19458;
wire wire19459;
wire wire19461;
wire wire19464;
wire wire19466;
wire wire19469;
wire wire19471;
wire wire19472;
wire wire19476;
wire wire19477;
wire wire19479;
wire wire19480;
wire wire19481;
wire wire19485;
wire wire19486;
wire wire19490;
wire wire19491;
wire wire19494;
wire wire19496;
wire wire19497;
wire wire19498;
wire wire19499;
wire wire19500;
wire wire19504;
wire wire19506;
wire wire19510;
wire wire19513;
wire wire19516;
wire wire19519;
wire wire19520;
wire wire19521;
wire wire19523;
wire wire19526;
wire wire19527;
wire wire19528;
wire wire19529;
wire wire19530;
wire wire19531;
wire wire19532;
wire wire19533;
wire wire19535;
wire wire19536;
wire wire19538;
wire wire19539;
wire wire19541;
wire wire19542;
wire wire19543;
wire wire19544;
wire wire19545;
wire wire19548;
wire wire19549;
wire wire19552;
wire wire19556;
wire wire19557;
wire wire19560;
wire wire19565;
wire wire19567;
wire wire19569;
wire wire19574;
wire wire19576;
wire wire19577;
wire wire19580;
wire wire19581;
wire wire19582;
wire wire19583;
wire wire19584;
wire wire19587;
wire wire19588;
wire wire19589;
wire wire19591;
wire wire19596;
wire wire19599;
wire wire19600;
wire wire19602;
wire wire19603;
wire wire19605;
wire wire19607;
wire wire19608;
wire wire19610;
wire wire19612;
wire wire19613;
wire wire19614;
wire wire19617;
wire wire19619;
wire wire19620;
wire wire19621;
wire wire19623;
wire wire19624;
wire wire19629;
wire wire19630;
wire wire19633;
wire wire19636;
wire wire19637;
wire wire19638;
wire wire19640;
wire wire19641;
wire wire19644;
wire wire19645;
wire wire19646;
wire wire19647;
wire wire19648;
wire wire19650;
wire wire19652;
wire wire19653;
wire wire19654;
wire wire19656;
wire wire19657;
wire wire19658;
wire wire19659;
wire wire19660;
wire wire19663;
wire wire19666;
wire wire19667;
wire wire19668;
wire wire19670;
wire wire19671;
wire wire19672;
wire wire19674;
wire wire19675;
wire wire19676;
wire wire19677;
wire wire19680;
wire wire19682;
wire wire19683;
wire wire19687;
wire wire19688;
wire wire19689;
wire wire19691;
wire wire19693;
wire wire19694;
wire wire19695;
wire wire19698;
wire wire19700;
wire wire19701;
wire wire19702;
wire wire19704;
wire wire19706;
wire wire19707;
wire wire19708;
wire wire19709;
wire wire19710;
wire wire19714;
wire wire19716;
wire wire19717;
wire wire19718;
wire wire19721;
wire wire19722;
wire wire19724;
wire wire19725;
wire wire19726;
wire wire19727;
wire wire19728;
wire wire19730;
wire wire19731;
wire wire19732;
wire wire19733;
wire wire19734;
wire wire19735;
wire wire19738;
wire wire19739;
wire wire19744;
wire wire19745;
wire wire19746;
wire wire19747;
wire wire19750;
wire wire19751;
wire wire19752;
wire wire19756;
wire wire19757;
wire wire19758;
wire wire19759;
wire wire19760;
wire wire19764;
wire wire19765;
wire wire19766;
wire wire19767;
wire wire19769;
wire wire19770;
wire wire19774;
wire wire19775;
wire wire19777;
wire wire19778;
wire wire19779;
wire wire19780;
wire wire19782;
wire wire19783;
wire wire19786;
wire wire19787;
wire wire19792;
wire wire19793;
wire wire19796;
wire wire19798;
wire wire19799;
wire wire19800;
wire wire19801;
wire wire19802;
wire wire19803;
wire wire19804;
wire wire19807;
wire wire19808;
wire wire19812;
wire wire19813;
wire wire19820;
wire wire19823;
wire wire19824;
wire wire19825;
wire wire19827;
wire wire19828;
wire wire19829;
wire wire19830;
wire wire19831;
wire wire19834;
wire wire19835;
wire wire19837;
wire wire19838;
wire wire19839;
wire wire19841;
wire wire19842;
wire wire19843;
wire wire19845;
wire wire19846;
wire wire19847;
wire wire19848;
wire wire19850;
wire wire19853;
wire wire19854;
wire wire19856;
wire wire19858;
wire wire19859;
wire wire19861;
wire wire19862;
wire wire19864;
wire wire19865;
wire wire19867;
wire wire19868;
wire wire19869;
wire wire19871;
wire wire19874;
wire wire19875;
wire wire19876;
wire wire19878;
wire wire19879;
wire wire19880;
wire wire19882;
wire wire19884;
wire wire19886;
wire wire19887;
wire wire19888;
wire wire19890;
wire wire19891;
wire wire19893;
wire wire19895;
wire wire19898;
wire wire19899;
wire wire19901;
wire wire19904;
wire wire19905;
wire wire19907;
wire wire19909;
wire wire19910;
wire wire19911;
wire wire19912;
wire wire19913;
wire wire19914;
wire wire19916;
wire wire19917;
wire wire19920;
wire wire19922;
wire wire19923;
wire wire19925;
wire wire19926;
wire wire19928;
wire wire19929;
wire wire19930;
wire wire19933;
wire wire19935;
wire wire19938;
wire wire19939;
wire wire19941;
wire wire19943;
wire wire19944;
wire wire19946;
assign o_1_ = ( wire5057 ) | ( wire16866 ) | ( wire16870 ) | ( wire16872 ) ;
 assign o_19_ = ( n_n5144 ) | ( wire736  &  wire16876 ) ;
 assign o_2_ = ( wire16877 ) | ( wire736  &  n_n162 ) ;
 assign o_0_ = ( n_n225 ) | ( wire16897 ) | ( wire16898 ) ;
 assign o_29_ = ( wire5026 ) | ( wire5027 ) | ( wire16911 ) ;
 assign o_39_ = ( n_n4721 ) | ( wire16933 ) ;
 assign o_38_ = ( n_n4397 ) | ( n_n4399 ) | ( wire17159 ) | ( wire17175 ) ;
 assign o_25_ = ( n_n5144 ) | ( n_n17  &  n_n159  &  wire17176 ) ;
 assign o_12_ = ( n_n2220 ) | ( wire17401 ) | ( wire17407 ) | ( wire17408 ) ;
 assign o_37_ = ( n_n4103 ) | ( n_n4102 ) | ( wire17582 ) | ( wire17586 ) ;
 assign o_26_ = ( n_n5144 ) | ( wire17600 ) | ( wire17601 ) | ( wire17602 ) ;
 assign o_11_ = ( wire17604 ) | ( wire17612 ) | ( n_n4  &  wire1495 ) ;
 assign o_36_ = ( wire17848 ) | ( wire17849 ) ;
 assign o_27_ = ( n_n5144 ) | ( wire17860 ) | ( wire17861 ) | ( wire17862 ) ;
 assign o_14_ = ( wire17876 ) | ( wire17877 ) | ( wire17913 ) | ( wire17915 ) ;
 assign o_35_ = ( wire18141 ) | ( wire18142 ) | ( wire18144 ) | ( wire18148 ) ;
 assign o_28_ = ( n_n2998 ) | ( wire18154 ) | ( wire18155 ) | ( wire18167 ) ;
 assign o_13_ = ( wire18212 ) | ( wire18213 ) | ( wire18215 ) | ( wire18225 ) ;
 assign o_34_ = ( wire18214 ) | ( wire18215 ) | ( wire18292 ) | ( wire18297 ) ;
 assign o_21_ = ( wire18299 ) | ( n_n10  &  wire185 ) | ( n_n10  &  wire270 ) ;
 assign o_16_ = ( n_n2721 ) | ( wire3442 ) | ( wire18310 ) | ( wire18311 ) ;
 assign o_40_ = ( n_n5144 ) | ( wire3439 ) | ( n_n135  &  wire267 ) ;
 assign o_33_ = ( n_n259 ) | ( wire18323 ) | ( wire18329 ) | ( wire18330 ) ;
 assign o_22_ = ( wire18332 ) | ( n_n14  &  wire185 ) | ( n_n14  &  wire270 ) ;
 assign o_15_ = ( n_n5144 ) | ( n_n2684 ) | ( wire18354 ) | ( wire18355 ) ;
 assign o_32_ = ( n_n3166 ) | ( wire18436 ) | ( wire18437 ) | ( wire18490 ) ;
 assign o_23_ = ( wire18498 ) | ( wire18499 ) | ( wire18508 ) | ( wire18512 ) ;
 assign o_18_ = ( wire18526 ) | ( wire18527 ) | ( wire18565 ) | ( wire18567 ) ;
 assign o_31_ = ( wire3194 ) | ( wire18568 ) | ( wire18572 ) ;
 assign o_24_ = ( n_n5144 ) | ( n_n16  &  n_n159  &  wire17176 ) ;
 assign o_17_ = ( n_n2748 ) | ( wire18621 ) | ( wire18623 ) ;
 assign o_43_ = ( wire18682 ) | ( wire18683 ) | ( wire18685 ) | ( wire18695 ) ;
 assign o_30_ = ( n_n3028 ) | ( wire18214 ) | ( wire18215 ) | ( wire18292 ) ;
 assign o_44_ = ( n_n4845 ) | ( wire18792 ) | ( wire18795 ) ;
 assign o_41_ = ( n_n5144 ) | ( wire2962 ) ;
 assign o_42_ = ( wire18802 ) | ( wire18803 ) | ( wire18807 ) ;
 assign o_20_ = ( n_n5144 ) | ( wire736  &  wire18809 ) ;
 assign o_45_ = ( wire18436 ) | ( wire18437 ) | ( wire18490 ) | ( wire18818 ) ;
 assign o_10_ = ( n_n5144 ) | ( wire19029 ) | ( wire19030 ) | ( wire19036 ) ;
 assign o_9_ = ( wire19348 ) | ( wire19349 ) | ( wire19458 ) | ( wire19459 ) ;
 assign o_7_ = ( n_n743 ) | ( wire19682 ) | ( wire19683 ) | ( wire19689 ) ;
 assign o_8_ = ( i_3_  &  (~ i_1_)  &  i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign o_5_ = ( wire19868 ) | ( wire19869 ) | ( wire19871 ) | ( wire19914 ) ;
 assign o_6_ = ( wire19922 ) | ( n_n5  &  wire238 ) | ( n_n5  &  wire19916 ) ;
 assign o_3_ = ( n_n259 ) | ( wire18323 ) | ( wire19928 ) ;
 assign o_4_ = ( n_n275 ) | ( wire441 ) | ( wire19941 ) | ( wire19946 ) ;
 assign wire428 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign n_n5144 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire736 = ( n_n184  &  n_n163  &  wire725  &  n_n35 ) ;
 assign n_n162 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n65 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign n_n71 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign n_n9 = ( n_n162  &  n_n124  &  n_n159 ) ;
 assign wire343 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign n_n38 = ( n_n124  &  n_n48  &  n_n220 ) ;
 assign n_n373 = ( wire5024 ) | ( n_n38  &  wire244 ) ;
 assign n_n374 = ( wire5022 ) | ( wire140  &  n_n39 ) ;
 assign n_n969 = ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) | ( n_n39  &  n_n132 ) ;
 assign n_n4721 = ( n_n39  &  wire244 ) | ( n_n38  &  wire1595 ) | ( n_n39  &  wire1595 ) ;
 assign n_n519 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign n_n4597 = ( n_n38  &  n_n134 ) | ( n_n38  &  n_n132 ) | ( n_n39  &  n_n132 ) ;
 assign wire140 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire390 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) ;
 assign wire393 = ( n_n38  &  n_n177  &  wire719 ) ;
 assign wire712 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n52 ) ;
 assign n_n31 = ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign n_n30 = ( n_n162  &  n_n220  &  n_n35 ) ;
 assign n_n4161 = ( n_n30  &  wire143 ) | ( n_n30  &  wire154 ) | ( n_n30  &  wire47 ) ;
 assign wire132 = ( n_n170  &  wire720 ) | ( n_n170  &  wire722 ) | ( n_n170  &  wire715 ) ;
 assign wire137 = ( wire723  &  n_n177 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire727 ) ;
 assign wire599 = ( n_n4449 ) | ( wire17164 ) | ( n_n30  &  wire1864 ) ;
 assign wire695 = ( n_n31  &  wire146 ) | ( n_n31  &  wire131 ) ;
 assign n_n17 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n2229 = ( wire4680 ) | ( wire17198 ) | ( wire17213 ) ;
 assign n_n2220 = ( n_n2239 ) | ( wire4643 ) | ( wire17234 ) | ( wire17249 ) ;
 assign n_n2232 = ( n_n2259 ) | ( wire17256 ) | ( wire17257 ) | ( wire17277 ) ;
 assign n_n2227 = ( wire4561 ) | ( wire4562 ) | ( wire17303 ) | ( wire17305 ) ;
 assign n_n2226 = ( n_n2241 ) | ( wire17321 ) | ( wire17322 ) | ( wire17327 ) ;
 assign n_n2228 = ( n_n2249 ) | ( wire17341 ) | ( wire17342 ) | ( wire17347 ) ;
 assign n_n2234 = ( n_n2265 ) | ( n_n2266 ) | ( wire17379 ) ;
 assign n_n4106 = ( wire599 ) | ( n_n4120 ) | ( wire4434 ) | ( wire17420 ) ;
 assign n_n7241 = ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign n_n7240 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) ;
 assign n_n51 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign n_n13 = ( n_n159  &  n_n111  &  wire747 ) ;
 assign n_n4 = ( n_n35  &  n_n159  &  n_n111 ) ;
 assign wire77 = ( wire717  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire431 = ( i_7_  &  i_6_  &  n_n19  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire529 = ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n111 ) ;
 assign wire568 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign wire569 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign n_n53 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign n_n3795 = ( n_n3825 ) | ( wire4060 ) | ( wire17726 ) | ( wire17729 ) ;
 assign n_n3787 = ( n_n3800 ) | ( n_n3802 ) | ( wire17798 ) ;
 assign n_n3789 = ( wire17831 ) | ( wire17832 ) | ( wire17836 ) | ( wire17839 ) ;
 assign wire157 = ( n_n156  &  wire719 ) | ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign wire213 = ( i_8_  &  n_n162  &  n_n157  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n157  &  n_n220 ) ;
 assign n_n36 = ( (~ i_7_)  &  (~ i_6_)  &  wire714  &  n_n218 ) ;
 assign n_n34 = ( n_n220  &  n_n35  &  n_n218 ) ;
 assign n_n2622 = ( wire597 ) | ( wire620 ) | ( n_n2630 ) | ( wire17884 ) ;
 assign n_n3454 = ( n_n3467 ) | ( wire17934 ) | ( wire17935 ) ;
 assign n_n3456 = ( n_n3473 ) | ( wire17958 ) | ( wire17959 ) | ( wire17968 ) ;
 assign n_n7263 = ( (~ i_7_)  &  (~ i_6_)  &  n_n48  &  n_n219 ) ;
 assign n_n14 = ( n_n161  &  n_n48  &  n_n159 ) ;
 assign n_n7265 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign n_n7267 = ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign n_n2998 = ( wire3628 ) | ( wire3629 ) | ( wire18150 ) ;
 assign wire253 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire717 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire717 ) ;
 assign n_n4308 = ( wire157  &  n_n161  &  n_n48  &  n_n220 ) ;
 assign n_n6271 = ( n_n177  &  n_n124  &  n_n220  &  n_n111 ) ;
 assign n_n6267 = ( n_n156  &  n_n126  &  n_n220  &  n_n111 ) ;
 assign n_n3085 = ( wire4260 ) | ( wire17554 ) | ( n_n47  &  wire152 ) ;
 assign n_n6266 = ( n_n177  &  n_n126  &  n_n220  &  n_n111 ) ;
 assign n_n6270 = ( n_n170  &  n_n126  &  n_n220  &  n_n111 ) ;
 assign n_n6269 = ( n_n149  &  n_n124  &  n_n220  &  n_n111 ) ;
 assign n_n6268 = ( n_n170  &  n_n124  &  n_n220  &  n_n111 ) ;
 assign n_n5052 = ( n_n17  &  wire245  &  n_n48  &  wire714 ) ;
 assign n_n5055 = ( n_n40  &  n_n57 ) | ( n_n41  &  wire144 ) ;
 assign wire608 = ( wire3469 ) | ( n_n41  &  wire122 ) ;
 assign n_n10 = ( n_n162  &  n_n161  &  n_n159 ) ;
 assign wire525 = ( n_n149  &  wire725  &  wire751 ) | ( n_n149  &  wire725  &  wire18298 ) ;
 assign n_n33 = ( n_n162  &  n_n200  &  n_n220 ) ;
 assign n_n2732 = ( n_n162  &  n_n17  &  wire714  &  wire1417 ) ;
 assign n_n2728 = ( n_n33  &  wire55 ) | ( n_n33  &  wire149 ) | ( n_n33  &  wire127 ) ;
 assign n_n2721 = ( wire675 ) | ( wire3451 ) | ( wire18301 ) | ( wire18302 ) ;
 assign wire587 = ( wire132  &  n_n33 ) | ( n_n33  &  wire126 ) ;
 assign wire767 = ( wire172 ) | ( wire147 ) | ( wire158 ) | ( wire133 ) ;
 assign n_n6 = ( n_n48  &  n_n35  &  n_n159 ) ;
 assign n_n135 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire267 = ( n_n126  &  n_n159  &  n_n111 ) | ( n_n159  &  n_n111  &  wire747 ) ;
 assign n_n3389 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign n_n5 = ( n_n124  &  n_n159  &  n_n111 ) ;
 assign wire145 = ( wire729  &  n_n191 ) | ( n_n191  &  wire730 ) ;
 assign wire388 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n219 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n219 ) ;
 assign wire770 = ( wire729  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign n_n3166 = ( n_n3179 ) | ( wire18374 ) | ( wire18375 ) | ( wire18377 ) ;
 assign n_n144 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire717 ) ;
 assign n_n7346 = ( i_7_  &  i_6_  &  n_n159  &  n_n218 ) ;
 assign n_n3 = ( n_n124  &  n_n159  &  n_n218 ) ;
 assign n_n2 = ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire708 = ( wire430 ) | ( wire77  &  n_n2 ) ;
 assign n_n18 = ( i_7_  &  i_6_ ) ;
 assign n_n5319 = ( i_5_  &  n_n157  &  n_n159  &  wire17176 ) ;
 assign wire430 = ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n218 ) ;
 assign wire684 = ( i_3_  &  i_4_  &  n_n159  &  wire17587 ) ;
 assign wire748 = ( i_5_  &  i_3_  &  i_4_  &  n_n159 ) ;
 assign n_n16 = ( (~ i_7_)  &  i_6_ ) ;
 assign n_n197 = ( n_n200  &  n_n220  &  n_n218 ) ;
 assign n_n212 = ( i_7_  &  (~ i_6_)  &  wire714  &  n_n218 ) ;
 assign n_n2748 = ( n_n4441 ) | ( wire575 ) | ( wire18577 ) | ( wire18578 ) ;
 assign n_n2747 = ( n_n2754 ) | ( wire18593 ) | ( wire18594 ) ;
 assign n_n101 = ( n_n162  &  n_n124  &  n_n220 ) ;
 assign n_n42 = ( n_n162  &  n_n161  &  n_n220 ) ;
 assign n_n4755 = ( wire3128 ) | ( wire18624 ) | ( wire18625 ) | ( wire18626 ) ;
 assign wire172 = ( n_n191  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n191  &  wire728 ) ;
 assign wire381 = ( n_n156  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n156  &  wire728 ) ;
 assign wire662 = ( n_n43  &  wire63 ) | ( n_n43  &  wire48 ) ;
 assign n_n3028 = ( wire608 ) | ( wire18711 ) | ( wire18712 ) | ( wire18719 ) ;
 assign n_n4845 = ( wire2977 ) | ( wire18783 ) | ( wire18789 ) | ( wire18790 ) ;
 assign n_n184 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n163 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n161 = ( i_7_  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n6005 = ( n_n200  &  n_n149  &  n_n220  &  n_n111 ) ;
 assign wire419 = ( n_n156  &  n_n220  &  n_n111  &  wire17072 ) ;
 assign wire445 = ( n_n177  &  n_n220  &  n_n111  &  wire17072 ) ;
 assign wire446 = ( n_n200  &  n_n170  &  n_n220  &  n_n111 ) ;
 assign n_n3179 = ( wire3469 ) | ( wire3470 ) | ( wire18360 ) | ( wire18361 ) ;
 assign wire95 = ( wire717  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign n_n743 = ( n_n799 ) | ( wire2310 ) | ( wire2311 ) | ( wire19504 ) ;
 assign wire777 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire776 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire775 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire185 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign n_n7252 = ( i_7_  &  i_6_  &  n_n162  &  n_n219 ) ;
 assign n_n7253 = ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n219 ) ;
 assign wire389 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n19 ) ;
 assign wire454 = ( wire3248 ) | ( wire77  &  n_n5 ) ;
 assign wire706 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n162  &  n_n219 ) ;
 assign wire742 = ( n_n126  &  n_n159  &  n_n111 ) ;
 assign wire779 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire783 = ( n_n126  &  n_n159  &  n_n111 ) | ( n_n159  &  n_n111  &  wire747 ) ;
 assign wire781 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire707 = ( wire430 ) | ( n_n2  &  wire185 ) ;
 assign n_n46 = ( n_n161  &  n_n48  &  n_n220 ) ;
 assign wire168 = ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire724 ) ;
 assign n_n47 = ( i_7_  &  i_6_  &  n_n48  &  wire714 ) ;
 assign n_n138 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire214 = ( n_n216  &  wire721 ) | ( n_n216  &  wire725 ) ;
 assign n_n5107 = ( n_n47  &  n_n138 ) | ( n_n46  &  wire214 ) ;
 assign n_n41 = ( i_7_  &  (~ i_6_)  &  n_n48  &  wire714 ) ;
 assign wire245 = ( n_n149  &  wire719 ) | ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign n_n108 = ( n_n162  &  n_n126  &  n_n220 ) ;
 assign n_n148 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign wire90 = ( wire729  &  n_n156 ) | ( wire726  &  n_n156 ) ;
 assign n_n5000 = ( n_n101  &  n_n148 ) | ( n_n108  &  wire90 ) ;
 assign n_n1434 = ( n_n31  &  wire98 ) | ( n_n30  &  n_n102 ) ;
 assign n_n1408 = ( n_n71  &  n_n31 ) | ( n_n30  &  wire118 ) ;
 assign wire789 = ( wire120 ) | ( wire179 ) | ( wire324 ) | ( wire18720 ) ;
 assign n_n1426 = ( n_n31  &  n_n117 ) | ( n_n30  &  wire98 ) ;
 assign wire791 = ( n_n89 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign n_n1416 = ( n_n31  &  wire53 ) | ( n_n30  &  n_n77 ) ;
 assign wire793 = ( wire53 ) | ( wire117 ) | ( wire281 ) | ( wire294 ) ;
 assign wire422 = ( n_n125  &  wire85 ) | ( n_n125  &  wire142 ) ;
 assign wire797 = ( n_n132 ) | ( wire150 ) | ( wire80 ) | ( wire78 ) ;
 assign wire796 = ( n_n55 ) | ( wire80 ) | ( wire78 ) | ( wire252 ) ;
 assign wire55 = ( wire720  &  n_n149 ) | ( wire722  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire207 = ( wire720  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign n_n1520 = ( n_n38  &  wire207 ) | ( n_n39  &  n_n150 ) ;
 assign wire800 = ( wire155 ) | ( wire205 ) | ( wire215 ) | ( wire17490 ) ;
 assign wire799 = ( n_n148 ) | ( wire234 ) | ( wire86 ) | ( wire84 ) ;
 assign n_n4581 = ( n_n220  &  n_n35  &  n_n218  &  wire181 ) ;
 assign wire458 = ( n_n36  &  wire134 ) | ( n_n36  &  wire156 ) ;
 assign wire541 = ( n_n36  &  wire176 ) | ( n_n36  &  wire123 ) ;
 assign n_n125 = ( n_n126  &  n_n220  &  n_n218 ) ;
 assign n_n3912 = ( wire4393 ) | ( n_n125  &  n_n216  &  wire719 ) ;
 assign n_n123 = ( n_n124  &  n_n220  &  n_n218 ) ;
 assign wire570 = ( wire90  &  n_n125 ) | ( n_n125  &  wire205 ) ;
 assign n_n1700 = ( n_n148  &  n_n125 ) | ( n_n123  &  wire60 ) ;
 assign wire803 = ( wire60 ) | ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign n_n4139 = ( wire4365 ) | ( wire17470 ) | ( wire17471 ) | ( wire17472 ) ;
 assign n_n4206 = ( wire4829 ) | ( n_n46  &  n_n199  &  wire720 ) ;
 assign n_n1624 = ( wire4354 ) | ( wire4355 ) | ( n_n47  &  n_n214 ) ;
 assign wire85 = ( n_n216  &  wire722 ) | ( n_n216  &  wire727 ) | ( n_n216  &  wire715 ) ;
 assign n_n4112 = ( n_n4139 ) | ( wire17478 ) | ( wire17479 ) | ( wire17486 ) ;
 assign n_n1594 = ( n_n46  &  n_n155 ) | ( n_n47  &  wire60 ) ;
 assign wire543 = ( wire17082 ) | ( n_n46  &  wire1842 ) | ( n_n46  &  wire17081 ) ;
 assign wire808 = ( n_n148 ) | ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign n_n4904 = ( n_n108  &  wire85 ) | ( n_n108  &  wire142 ) | ( n_n108  &  wire180 ) ;
 assign n_n5037 = ( wire447 ) | ( wire4320 ) | ( n_n108  &  n_n214 ) ;
 assign n_n4903 = ( n_n5033 ) | ( n_n101  &  wire219 ) | ( n_n101  &  wire108 ) ;
 assign wire544 = ( wire4935 ) | ( n_n108  &  wire1844 ) ;
 assign n_n4103 = ( n_n4112 ) | ( wire543 ) | ( wire17501 ) | ( wire17514 ) ;
 assign wire52 = ( n_n191  &  wire716 ) | ( n_n191  &  wire717 ) | ( n_n191  &  wire718 ) ;
 assign wire176 = ( wire729  &  n_n156 ) | ( wire726  &  n_n156 ) | ( wire724  &  n_n156 ) ;
 assign n_n4007 = ( n_n161  &  wire176  &  n_n48  &  n_n220 ) ;
 assign wire129 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( wire724  &  n_n191 ) ;
 assign wire142 = ( wire723  &  n_n216 ) | ( n_n216  &  wire716 ) | ( n_n216  &  wire730 ) ;
 assign n_n4622 = ( n_n17  &  wire142  &  n_n48  &  wire714 ) ;
 assign wire182 = ( n_n177  &  wire719 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign n_n5060 = ( n_n17  &  wire182  &  n_n48  &  wire714 ) ;
 assign n_n40 = ( n_n200  &  n_n48  &  n_n220 ) ;
 assign n_n130 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire134 = ( wire720  &  n_n156 ) | ( n_n156  &  wire722 ) | ( n_n156  &  wire715 ) ;
 assign wire123 = ( wire716  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign n_n3276 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n48 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n48 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n48 ) ;
 assign wire53 = ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) ;
 assign n_n83 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign n_n6445 = ( n_n41  &  wire729  &  n_n177 ) ;
 assign n_n7242 = ( i_7_  &  i_6_  &  n_n19  &  n_n48 ) ;
 assign n_n68 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire344 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire730 ) ;
 assign n_n19 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire462 = ( i_7_  &  i_6_  &  n_n19  &  n_n218 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n218 ) ;
 assign wire817 = ( i_5_  &  (~ i_3_)  &  i_4_ ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire149 = ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) | ( wire724  &  n_n170 ) ;
 assign wire130 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire724 ) ;
 assign wire188 = ( i_8_  &  n_n17  &  n_n220  &  n_n218 ) | ( (~ i_8_)  &  n_n17  &  n_n220  &  n_n218 ) ;
 assign n_n59 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire226 = ( i_8_  &  n_n157  &  n_n220  &  n_n218 ) | ( (~ i_8_)  &  n_n157  &  n_n220  &  n_n218 ) ;
 assign wire820 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire819 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign n_n2284 = ( wire4558 ) | ( wire17307 ) | ( wire226  &  wire819 ) ;
 assign n_n2241 = ( n_n2284 ) | ( wire4554 ) | ( wire17314 ) ;
 assign wire824 = ( wire129 ) | ( wire130 ) | ( wire304 ) | ( wire306 ) ;
 assign n_n2253 = ( wire4701 ) | ( wire17178 ) | ( n_n46  &  wire824 ) ;
 assign n_n61 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) ;
 assign wire228 = ( i_8_  &  n_n162  &  n_n16  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n16  &  n_n220 ) ;
 assign wire827 = ( n_n147 ) | ( n_n63 ) | ( wire60 ) | ( wire351 ) ;
 assign wire826 = ( n_n154 ) | ( n_n63 ) | ( wire60 ) | ( wire377 ) ;
 assign n_n43 = ( i_7_  &  i_6_  &  n_n162  &  wire714 ) ;
 assign wire139 = ( n_n184  &  wire716 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire718 ) ;
 assign n_n117 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire257 = ( i_15_  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n213  &  n_n191 ) ;
 assign wire313 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) ;
 assign n_n129 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign n_n166 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire716 ) ;
 assign n_n127 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign n_n39 = ( n_n126  &  n_n48  &  n_n220 ) ;
 assign n_n82 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) ;
 assign wire190 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire334 = ( i_8_  &  n_n16  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n16  &  n_n48  &  n_n220 ) ;
 assign wire836 = ( n_n177  &  wire716 ) | ( n_n177  &  wire715 ) | ( n_n170  &  wire715 ) ;
 assign n_n139 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) ;
 assign wire838 = ( wire260 ) | ( wire373 ) | ( n_n216  &  wire721 ) ;
 assign n_n1819 = ( wire2896 ) | ( wire2900 ) | ( wire2901 ) | ( wire18863 ) ;
 assign n_n1870 = ( wire18865 ) | ( wire18866 ) | ( n_n36  &  wire143 ) ;
 assign wire840 = ( wire257 ) | ( n_n95 ) | ( wire74 ) | ( wire136 ) ;
 assign n_n1800 = ( n_n1819 ) | ( wire18857 ) | ( wire18858 ) | ( wire18874 ) ;
 assign wire68 = ( n_n199  &  wire723 ) | ( n_n199  &  wire730 ) | ( n_n199  &  wire727 ) ;
 assign n_n4591 = ( wire68  &  n_n220  &  n_n35  &  n_n218 ) ;
 assign wire147 = ( wire716  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire718 ) ;
 assign wire98 = ( n_n191  &  wire720 ) | ( n_n191  &  wire715 ) ;
 assign n_n2715 = ( n_n161  &  n_n220  &  wire63  &  n_n218 ) ;
 assign n_n112 = ( n_n161  &  n_n220  &  n_n218 ) ;
 assign n_n113 = ( i_7_  &  i_6_  &  wire714  &  n_n218 ) ;
 assign wire844 = ( wire155 ) | ( wire127 ) | ( wire227 ) | ( wire232 ) ;
 assign wire845 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire542 = ( n_n36  &  n_n148 ) | ( n_n34  &  wire127 ) ;
 assign wire614 = ( n_n36  &  wire729  &  n_n156 ) ;
 assign wire850 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire849 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign n_n5109 = ( n_n65  &  n_n46 ) | ( n_n47  &  wire118 ) ;
 assign wire677 = ( n_n47  &  wire133 ) | ( n_n47  &  wire127 ) ;
 assign wire852 = ( wire118 ) | ( wire234 ) | ( wire75 ) | ( wire19119 ) ;
 assign n_n140 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) ;
 assign n_n142 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) ;
 assign wire856 = ( wire290 ) | ( wire720  &  n_n156 ) | ( n_n156  &  wire715 ) ;
 assign n_n116 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire255 = ( i_8_  &  n_n16  &  n_n220  &  n_n218 ) | ( (~ i_8_)  &  n_n16  &  n_n220  &  n_n218 ) ;
 assign wire601 = ( n_n125  &  n_n216  &  wire719 ) ;
 assign wire859 = ( wire199 ) | ( wire402 ) | ( wire19640 ) | ( wire19641 ) ;
 assign n_n157 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign wire733 = ( (~ i_1_)  &  i_2_  &  i_0_  &  n_n111 ) ;
 assign wire743 = ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n219 ) ;
 assign n_n213 = ( i_14_  &  i_13_  &  (~ i_12_) ) ;
 assign n_n199 = ( (~ i_9_)  &  i_10_  &  i_11_ ) ;
 assign wire723 = ( i_14_  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign wire729 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign n_n95 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire729 ) ;
 assign n_n200 = ( i_7_  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire726 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign n_n216 = ( i_9_  &  i_10_  &  i_11_ ) ;
 assign wire724 = ( (~ i_14_)  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign n_n103 = ( i_9_  &  i_10_  &  i_11_  &  wire724 ) ;
 assign n_n191 = ( i_9_  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n89 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign n_n207 = ( (~ i_14_)  &  i_13_  &  i_12_ ) ;
 assign n_n177 = ( i_9_  &  (~ i_10_)  &  i_11_ ) ;
 assign wire716 = ( (~ i_14_)  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign n_n173 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire716 ) ;
 assign n_n170 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) ;
 assign wire720 = ( i_14_  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign n_n169 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign n_n204 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire717 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign wire730 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign wire718 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_  &  i_15_ ) ;
 assign n_n156 = ( i_9_  &  i_10_  &  (~ i_11_) ) ;
 assign wire722 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  i_15_ ) ;
 assign n_n154 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign n_n205 = ( (~ i_14_)  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n150 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign n_n149 = ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign n_n151 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire717 ) ;
 assign wire719 = ( i_14_  &  i_13_  &  i_12_  &  i_15_ ) ;
 assign wire721 = ( (~ i_14_)  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign n_n141 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) ;
 assign n_n115 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign n_n209 = ( i_14_  &  i_13_  &  i_12_ ) ;
 assign n_n134 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign wire725 = ( (~ i_14_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_15_) ) ;
 assign n_n55 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) ;
 assign wire728 = ( i_14_  &  (~ i_13_)  &  i_12_  &  (~ i_15_) ) ;
 assign n_n54 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign n_n126 = ( (~ i_7_)  &  i_8_  &  i_6_ ) ;
 assign n_n124 = ( (~ i_7_)  &  (~ i_8_)  &  i_6_ ) ;
 assign n_n92 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire730 ) ;
 assign wire727 = ( i_14_  &  i_13_  &  i_12_  &  (~ i_15_) ) ;
 assign n_n178 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign n_n57 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) ;
 assign wire715 = ( i_14_  &  i_13_  &  (~ i_12_)  &  i_15_ ) ;
 assign n_n48 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign wire714 = ( i_8_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n183 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign n_n90 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign n_n70 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire715 ) ;
 assign n_n62 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) ;
 assign n_n189 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign n_n122 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign n_n185 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign n_n84 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign n_n147 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign n_n136 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign n_n220 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n52 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign n_n35 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n210 = ( i_9_  &  i_10_  &  i_11_  &  wire722 ) ;
 assign n_n172 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire717 ) ;
 assign n_n58 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) ;
 assign n_n118 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign n_n32 = ( i_7_  &  (~ i_6_)  &  n_n162  &  wire714 ) ;
 assign n_n186 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire717 ) ;
 assign n_n107 = ( i_9_  &  i_10_  &  i_11_  &  wire715 ) ;
 assign n_n198 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire720 ) ;
 assign n_n168 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) ;
 assign n_n176 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) ;
 assign n_n60 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign n_n219 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n12 = ( n_n124  &  n_n48  &  n_n159 ) ;
 assign n_n159 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire151 = ( n_n199  &  wire720 ) | ( n_n199  &  wire722 ) | ( n_n199  &  wire715 ) ;
 assign wire860 = ( wire94 ) | ( wire184 ) | ( wire268 ) | ( wire18738 ) ;
 assign n_n1442 = ( n_n30  &  wire81 ) | ( n_n31  &  n_n102 ) ;
 assign wire863 = ( wire111 ) | ( wire162 ) | ( wire164 ) | ( wire341 ) ;
 assign wire865 = ( wire206 ) | ( wire243 ) | ( wire368 ) | ( wire18752 ) ;
 assign n_n4686 = ( n_n212  &  n_n140 ) | ( n_n197  &  wire153 ) ;
 assign wire247 = ( n_n199  &  wire721 ) | ( n_n199  &  wire725 ) | ( n_n199  &  wire728 ) ;
 assign wire704 = ( n_n212  &  n_n63 ) | ( n_n197  &  wire135 ) ;
 assign n_n4231 = ( n_n4686 ) | ( wire704 ) | ( n_n212  &  wire247 ) ;
 assign wire158 = ( wire729  &  n_n149 ) | ( wire726  &  n_n149 ) | ( wire724  &  n_n149 ) ;
 assign wire155 = ( wire723  &  n_n156 ) | ( wire716  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign wire218 = ( n_n199  &  wire719 ) | ( n_n199  &  wire721 ) | ( n_n199  &  wire728 ) ;
 assign wire180 = ( n_n216  &  wire724 ) | ( n_n216  &  wire717 ) | ( n_n216  &  wire718 ) ;
 assign wire248 = ( wire723  &  n_n156 ) | ( wire730  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign n_n4460 = ( n_n36  &  wire168 ) | ( n_n36  &  wire68 ) | ( n_n36  &  wire74 ) ;
 assign n_n4900 = ( n_n101  &  wire85 ) | ( n_n101  &  wire142 ) | ( n_n101  &  wire180 ) ;
 assign wire867 = ( wire155 ) | ( n_n155 ) | ( wire205 ) | ( wire215 ) ;
 assign n_n4388 = ( n_n200  &  n_n220  &  wire133  &  n_n218 ) ;
 assign n_n4441 = ( n_n4518 ) | ( wire17100 ) | ( n_n197  &  wire1224 ) ;
 assign wire532 = ( n_n212  &  wire133 ) | ( n_n212  &  wire127 ) ;
 assign wire575 = ( wire4739 ) | ( wire4740 ) | ( wire17102 ) ;
 assign wire594 = ( n_n197  &  wire55 ) | ( n_n212  &  wire176 ) ;
 assign wire660 = ( n_n212  &  wire134 ) | ( n_n212  &  wire156 ) ;
 assign n_n4116 = ( n_n4441 ) | ( wire575 ) | ( wire17521 ) | ( wire17522 ) ;
 assign wire156 = ( wire723  &  n_n156 ) | ( wire730  &  n_n156 ) | ( n_n156  &  wire727 ) ;
 assign n_n77 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire104 = ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign n_n5111 = ( n_n47  &  n_n77 ) | ( n_n46  &  wire104 ) ;
 assign n_n5113 = ( n_n46  &  n_n89 ) | ( n_n47  &  wire104 ) ;
 assign wire868 = ( wire98 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign n_n7254 = ( (~ i_7_)  &  i_6_  &  n_n162  &  n_n219 ) ;
 assign n_n7248 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n218 ) ;
 assign n_n3562 = ( wire168  &  n_n47 ) | ( n_n47  &  wire68 ) | ( n_n47  &  wire74 ) ;
 assign wire63 = ( wire723  &  n_n191 ) | ( n_n191  &  wire730 ) | ( n_n191  &  wire727 ) ;
 assign n_n3398 = ( n_n3562 ) | ( wire3601 ) | ( wire18168 ) | ( wire18169 ) ;
 assign wire143 = ( n_n216  &  wire716 ) | ( n_n216  &  wire717 ) | ( n_n216  &  wire718 ) ;
 assign wire481 = ( n_n47  &  wire154 ) | ( n_n47  &  wire47 ) ;
 assign n_n3050 = ( wire3594 ) | ( wire18172 ) | ( wire18173 ) | ( wire18174 ) ;
 assign wire875 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign n_n3033 = ( n_n3398 ) | ( n_n3050 ) | ( wire18180 ) ;
 assign wire711 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign wire878 = ( n_n65 ) | ( wire77 ) | ( n_n89 ) | ( wire87 ) ;
 assign wire877 = ( n_n161  &  n_n48  &  n_n159 ) | ( n_n124  &  n_n48  &  n_n159 ) ;
 assign wire879 = ( wire87 ) | ( wire729  &  n_n191 ) | ( wire729  &  n_n149 ) ;
 assign n_n2948 = ( i_7_  &  i_6_  &  n_n48  &  n_n219 ) | ( (~ i_7_)  &  i_6_  &  n_n48  &  n_n219 ) | ( i_7_  &  (~ i_6_)  &  n_n48  &  n_n219 ) ;
 assign n_n231 = ( wire431 ) | ( wire389 ) | ( n_n7242 ) | ( wire16880 ) ;
 assign wire308 = ( i_15_  &  n_n204  &  n_n156 ) | ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire887 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire189 = ( i_8_  &  n_n18  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n18  &  n_n48  &  n_n220 ) ;
 assign wire888 = ( n_n59 ) | ( wire158 ) | ( wire299 ) | ( wire417 ) ;
 assign wire896 = ( i_8_  &  n_n162  &  n_n18  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n18  &  n_n220 ) ;
 assign wire894 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire561 = ( n_n161  &  n_n48  &  n_n220  &  wire131 ) ;
 assign n_n2239 = ( wire4658 ) | ( wire4659 ) | ( wire17217 ) ;
 assign wire899 = ( wire129 ) | ( wire130 ) | ( wire304 ) | ( wire306 ) ;
 assign wire902 = ( wire308 ) | ( wire131 ) | ( wire200 ) | ( wire201 ) ;
 assign wire133 = ( wire716  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire376 = ( i_15_  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n213  &  n_n149 ) ;
 assign wire904 = ( i_15_  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n201 ) ;
 assign n_n1862 = ( wire2861 ) | ( wire18892 ) | ( n_n36  &  wire123 ) ;
 assign wire583 = ( n_n34  &  wire729  &  n_n170 ) ;
 assign wire911 = ( i_15_  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n213  &  n_n177 ) | ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) ;
 assign n_n1799 = ( n_n1862 ) | ( wire18897 ) | ( wire18898 ) | ( wire18901 ) ;
 assign wire126 = ( wire723  &  n_n170 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire727 ) ;
 assign wire913 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign n_n2881 = ( wire147  &  n_n126  &  n_n220  &  n_n218 ) ;
 assign n_n1708 = ( n_n123  &  n_n176 ) | ( n_n125  &  wire69 ) ;
 assign wire916 = ( wire118 ) | ( wire179 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n1717 = ( n_n125  &  n_n176 ) | ( n_n123  &  wire51 ) ;
 assign wire639 = ( n_n123  &  wire729  &  n_n170 ) ;
 assign wire564 = ( n_n33  &  wire133 ) | ( n_n33  &  wire127 ) ;
 assign wire924 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign n_n1170 = ( wire2610 ) | ( wire19138 ) | ( n_n32  &  wire924 ) ;
 assign wire925 = ( wire142 ) | ( wire70 ) | ( wire233 ) | ( wire251 ) ;
 assign wire928 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign n_n4674 = ( n_n125  &  n_n198 ) | ( n_n123  &  wire70 ) ;
 assign n_n78 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire724 ) ;
 assign n_n974 = ( wire53  &  n_n39 ) | ( n_n38  &  n_n78 ) ;
 assign wire933 = ( i_15_  &  n_n170  &  n_n205 ) | ( (~ i_15_)  &  n_n170  &  n_n205 ) | ( i_15_  &  n_n170  &  n_n215 ) ;
 assign n_n7260 = ( i_7_  &  i_6_  &  n_n48  &  n_n219 ) ;
 assign n_n275 = ( wire525 ) | ( n_n7266 ) | ( wire19929 ) | ( wire19933 ) ;
 assign wire551 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n218 ) ;
 assign wire751 = ( n_n126  &  n_n159  &  n_n218 ) ;
 assign n_n202 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) ;
 assign n_n215 = ( i_14_  &  (~ i_13_)  &  i_12_ ) ;
 assign n_n72 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire724 ) ;
 assign n_n63 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) ;
 assign n_n131 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) ;
 assign n_n201 = ( (~ i_14_)  &  i_13_  &  (~ i_12_) ) ;
 assign n_n182 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign n_n132 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) ;
 assign n_n143 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire726 ) ;
 assign n_n137 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign n_n128 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n190 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign n_n214 = ( i_9_  &  i_10_  &  i_11_  &  wire720 ) ;
 assign n_n196 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire722 ) ;
 assign n_n64 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) ;
 assign n_n175 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire722 ) ;
 assign n_n171 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign n_n218 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n7264 = ( i_7_  &  i_6_  &  n_n219  &  n_n218 ) ;
 assign n_n74 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire118 = ( wire720  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire566 = ( n_n33  &  wire55 ) | ( n_n33  &  wire149 ) ;
 assign wire670 = ( wire139  &  n_n32 ) | ( n_n32  &  wire128 ) ;
 assign n_n4808 = ( n_n162  &  n_n161  &  n_n220  &  wire128 ) ;
 assign wire683 = ( n_n43  &  wire124 ) | ( n_n43  &  wire128 ) ;
 assign wire524 = ( n_n43  &  n_n191  &  wire725 ) ;
 assign wire672 = ( n_n42  &  wire63 ) | ( n_n42  &  wire48 ) ;
 assign n_n4564 = ( n_n36  &  n_n140 ) | ( n_n34  &  wire153 ) ;
 assign wire709 = ( n_n36  &  n_n63 ) | ( n_n34  &  wire135 ) ;
 assign n_n4169 = ( n_n4564 ) | ( wire709 ) | ( n_n36  &  wire247 ) ;
 assign wire942 = ( n_n55 ) | ( wire80 ) | ( wire78 ) | ( wire252 ) ;
 assign n_n155 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire720 ) ;
 assign wire60 = ( wire729  &  n_n149 ) | ( wire726  &  n_n149 ) ;
 assign wire359 = ( n_n41  &  wire729  &  n_n216 ) | ( n_n41  &  wire726  &  n_n216 ) ;
 assign n_n1514 = ( n_n38  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign wire597 = ( wire432 ) | ( wire17034 ) | ( wire17035 ) ;
 assign n_n4996 = ( n_n108  &  n_n148 ) | ( n_n101  &  wire60 ) ;
 assign n_n4994 = ( n_n162  &  n_n126  &  n_n220  &  wire234 ) ;
 assign wire511 = ( n_n101  &  n_n155 ) | ( n_n108  &  wire60 ) ;
 assign wire946 = ( wire155 ) | ( wire234 ) | ( wire215 ) | ( wire220 ) ;
 assign n_n4120 = ( n_n4161 ) | ( wire449 ) | ( wire656 ) | ( wire17410 ) ;
 assign wire122 = ( n_n156  &  wire721 ) | ( n_n156  &  wire725 ) ;
 assign wire443 = ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) ;
 assign n_n4240 = ( n_n30  &  n_n128 ) | ( n_n31  &  wire122 ) ;
 assign n_n4154 = ( wire4965 ) | ( wire4966 ) | ( n_n31  &  n_n63 ) ;
 assign wire144 = ( n_n156  &  wire719 ) | ( n_n156  &  wire728 ) ;
 assign wire654 = ( n_n30  &  wire176 ) | ( n_n30  &  wire123 ) ;
 assign wire739 = ( n_n156  &  n_n220  &  n_n111 ) ;
 assign wire279 = ( n_n177  &  wire716 ) | ( n_n177  &  wire722 ) | ( n_n177  &  wire727 ) ;
 assign n_n4600 = ( n_n124  &  n_n48  &  n_n220  &  wire279 ) ;
 assign n_n4602 = ( n_n126  &  n_n48  &  n_n220  &  wire279 ) ;
 assign wire605 = ( n_n39  &  wire279 ) | ( n_n39  &  wire724  &  n_n177 ) ;
 assign wire146 = ( n_n177  &  wire716 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign wire59 = ( wire720  &  n_n156 ) | ( n_n156  &  wire715 ) ;
 assign n_n5075 = ( n_n65  &  n_n41 ) | ( n_n40  &  wire59 ) ;
 assign wire498 = ( n_n47  &  n_n89 ) | ( n_n46  &  wire54 ) ;
 assign wire951 = ( n_n117 ) | ( wire94 ) | ( wire184 ) | ( wire268 ) ;
 assign n_n6492 = ( n_n41  &  wire726  &  n_n156 ) ;
 assign wire152 = ( n_n149  &  wire721 ) | ( n_n149  &  wire725 ) | ( n_n149  &  wire728 ) ;
 assign n_n3413 = ( n_n71  &  n_n41 ) | ( n_n40  &  wire118 ) ;
 assign wire546 = ( wire137  &  n_n46 ) | ( n_n46  &  wire146 ) ;
 assign wire674 = ( n_n47  &  wire134 ) | ( n_n47  &  wire156 ) ;
 assign n_n3889 = ( wire137  &  n_n47 ) | ( n_n47  &  wire146 ) | ( n_n47  &  wire131 ) ;
 assign wire671 = ( n_n46  &  wire63 ) | ( n_n46  &  wire48 ) ;
 assign wire463 = ( i_7_  &  i_6_  &  n_n48  &  n_n219 ) | ( i_7_  &  (~ i_6_)  &  n_n48  &  n_n219 ) ;
 assign wire958 = ( wire132 ) | ( wire149 ) | ( wire126 ) ;
 assign wire960 = ( wire55 ) | ( wire158 ) | ( wire133 ) | ( wire127 ) ;
 assign wire959 = ( wire134 ) | ( wire123 ) | ( wire158 ) | ( wire156 ) ;
 assign n_n2813 = ( wire18555 ) | ( n_n125  &  wire1730 ) ;
 assign wire181 = ( wire729  &  n_n216 ) | ( wire726  &  n_n216 ) | ( n_n216  &  wire724 ) ;
 assign n_n2265 = ( wire4485 ) | ( wire4486 ) | ( wire17367 ) | ( wire17368 ) ;
 assign wire93 = ( wire726  &  n_n191 ) | ( wire724  &  n_n191 ) | ( n_n191  &  wire717 ) ;
 assign wire968 = ( i_8_  &  n_n162  &  n_n157  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n157  &  n_n220 ) ;
 assign wire971 = ( wire115 ) | ( wire116 ) | ( wire371 ) | ( wire17253 ) ;
 assign n_n5739 = ( n_n161  &  n_n216  &  n_n220  &  n_n111 ) ;
 assign n_n2340 = ( wire17258 ) | ( wire17259 ) | ( wire17260 ) ;
 assign n_n5743 = ( n_n161  &  n_n177  &  n_n220  &  n_n111 ) ;
 assign wire440 = ( n_n161  &  n_n191  &  n_n220  &  n_n111 ) ;
 assign wire447 = ( n_n161  &  n_n156  &  n_n220  &  n_n111 ) ;
 assign wire973 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( n_n191  &  wire725 ) ;
 assign n_n2259 = ( n_n2340 ) | ( wire4619 ) | ( wire4620 ) | ( wire17268 ) ;
 assign wire975 = ( wire117 ) | ( wire120 ) | ( wire366 ) | ( wire17272 ) ;
 assign wire979 = ( i_8_  &  n_n157  &  n_n220  &  n_n218 ) | ( (~ i_8_)  &  n_n157  &  n_n220  &  n_n218 ) ;
 assign wire978 = ( i_15_  &  n_n199  &  n_n211 ) | ( (~ i_15_)  &  n_n199  &  n_n211 ) | ( i_15_  &  n_n191  &  n_n211 ) | ( (~ i_15_)  &  n_n191  &  n_n211 ) ;
 assign wire980 = ( wire117 ) | ( wire120 ) | ( wire362 ) | ( wire366 ) ;
 assign n_n2249 = ( n_n2310 ) | ( wire17333 ) | ( wire17335 ) ;
 assign wire397 = ( n_n41  &  wire729  &  n_n177 ) | ( n_n41  &  wire726  &  n_n177 ) ;
 assign wire984 = ( n_n168 ) | ( n_n175 ) | ( wire229 ) | ( wire265 ) ;
 assign wire989 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire988 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire993 = ( wire302 ) | ( wire303 ) | ( wire316 ) | ( wire18831 ) ;
 assign n_n1809 = ( wire18832 ) | ( n_n31  &  wire993 ) ;
 assign wire685 = ( n_n108  &  wire123 ) | ( n_n108  &  wire156 ) ;
 assign n_n5011 = ( n_n108  &  n_n169 ) | ( n_n101  &  wire69 ) ;
 assign wire81 = ( n_n199  &  wire720 ) | ( n_n199  &  wire715 ) ;
 assign n_n1517 = ( n_n39  &  n_n143 ) | ( n_n38  &  wire110 ) ;
 assign wire457 = ( wire207  &  n_n39 ) | ( n_n38  &  n_n143 ) ;
 assign wire572 = ( n_n126  &  n_n48  &  n_n220  &  wire110 ) ;
 assign wire1003 = ( wire716  &  n_n170 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire715 ) ;
 assign wire1006 = ( n_n176 ) | ( wire179 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n832 = ( wire2239 ) | ( wire2240 ) | ( n_n42  &  n_n190 ) ;
 assign wire1012 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1017 = ( wire111 ) | ( wire291 ) | ( wire297 ) | ( wire19621 ) ;
 assign n_n102 = ( i_9_  &  i_10_  &  i_11_  &  wire729 ) ;
 assign n_n56 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) ;
 assign n_n133 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) ;
 assign n_n4915 = ( n_n162  &  wire172  &  n_n157  &  wire714 ) ;
 assign wire1021 = ( wire247 ) | ( wire116 ) | ( wire198 ) | ( wire18773 ) ;
 assign wire1023 = ( wire182 ) | ( wire186 ) | ( wire217 ) | ( wire18780 ) ;
 assign wire1022 = ( n_n132 ) | ( wire150 ) | ( wire256 ) | ( wire216 ) ;
 assign wire224 = ( wire724  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign n_n4981 = ( n_n101  &  n_n59 ) | ( n_n108  &  wire80 ) ;
 assign wire1030 = ( wire208 ) | ( wire225 ) | ( wire148 ) | ( wire17083 ) ;
 assign wire127 = ( wire723  &  n_n149 ) | ( wire730  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire70 = ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) ;
 assign n_n4620 = ( n_n41  &  n_n198 ) | ( n_n40  &  wire70 ) ;
 assign n_n4131 = ( wire17528 ) | ( wire17529 ) | ( n_n40  &  wire1173 ) ;
 assign n_n4109 = ( n_n4131 ) | ( wire17533 ) | ( wire17534 ) | ( wire17539 ) ;
 assign wire249 = ( wire723  &  n_n149 ) | ( wire730  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire571 = ( wire157  &  n_n40 ) | ( n_n40  &  n_n156  &  wire725 ) ;
 assign wire620 = ( n_n4460 ) | ( wire17033 ) ;
 assign wire549 = ( n_n41  &  wire85 ) | ( n_n41  &  wire142 ) | ( n_n41  &  n_n214 ) ;
 assign wire621 = ( n_n4476 ) | ( wire537 ) | ( wire4842 ) | ( wire17007 ) ;
 assign n_n4102 = ( n_n4109 ) | ( wire17552 ) | ( wire17553 ) | ( wire17566 ) ;
 assign n_n3417 = ( n_n41  &  n_n117 ) | ( n_n40  &  wire98 ) ;
 assign n_n6384 = ( n_n40  &  wire726  &  n_n216 ) ;
 assign n_n3419 = ( n_n41  &  wire98 ) | ( n_n40  &  n_n102 ) ;
 assign wire1036 = ( n_n89 ) | ( wire93 ) | ( wire241 ) | ( wire273 ) ;
 assign n_n3421 = ( n_n40  &  wire81 ) | ( n_n41  &  n_n102 ) ;
 assign wire391 = ( n_n41  &  n_n216  &  wire720 ) | ( n_n41  &  n_n216  &  wire715 ) ;
 assign wire1042 = ( n_n9 ) | ( n_n14 ) | ( n_n10 ) | ( n_n12 ) ;
 assign wire1041 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire745 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_  &  n_n111 ) ;
 assign wire231 = ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) ;
 assign wire1044 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire1049 = ( wire129 ) | ( wire131 ) | ( wire200 ) | ( wire304 ) ;
 assign n_n2266 = ( wire4481 ) | ( wire17374 ) | ( n_n212  &  wire1049 ) ;
 assign wire526 = ( n_n42  &  n_n59 ) | ( n_n135  &  n_n43 ) ;
 assign n_n2310 = ( wire524 ) | ( wire526 ) | ( wire4531 ) | ( wire17329 ) ;
 assign wire1052 = ( n_n210 ) | ( n_n196 ) | ( wire70 ) | ( wire374 ) ;
 assign wire1056 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign n_n2257 = ( wire4505 ) | ( wire4506 ) | ( wire4508 ) | ( wire4509 ) ;
 assign wire1060 = ( n_n175 ) | ( wire69 ) | ( wire229 ) | ( wire265 ) ;
 assign wire1064 = ( wire86 ) | ( wire263 ) | ( wire374 ) | ( wire17361 ) ;
 assign wire250 = ( wire723  &  n_n177 ) | ( n_n177  &  wire716 ) | ( n_n177  &  wire730 ) ;
 assign wire227 = ( wire720  &  n_n156 ) | ( n_n156  &  wire727 ) | ( n_n156  &  wire715 ) ;
 assign wire1069 = ( n_n176 ) | ( wire179 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n5019 = ( n_n101  &  n_n190 ) | ( n_n108  &  wire62 ) ;
 assign wire1070 = ( wire139 ) | ( wire128 ) | ( wire54 ) | ( wire19179 ) ;
 assign n_n5033 = ( n_n101  &  n_n198 ) | ( n_n108  &  wire86 ) ;
 assign wire65 = ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) ;
 assign wire111 = ( n_n216  &  wire720 ) | ( n_n216  &  wire715 ) ;
 assign wire760 = ( n_n220  &  n_n111  &  wire1902  &  wire16987 ) ;
 assign wire1072 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire1075 = ( wire385 ) | ( wire108 ) | ( wire19196 ) | ( wire19197 ) ;
 assign wire1077 = ( wire98 ) | ( wire51 ) | ( wire148 ) | ( wire277 ) ;
 assign wire1079 = ( wire51 ) | ( wire276 ) | ( wire211 ) | ( wire271 ) ;
 assign n_n972 = ( n_n38  &  n_n84 ) | ( n_n39  &  wire110 ) ;
 assign wire48 = ( n_n191  &  wire720 ) | ( n_n191  &  wire722 ) | ( n_n191  &  wire715 ) ;
 assign wire1084 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) | ( i_15_  &  n_n191  &  n_n209 ) ;
 assign wire1089 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1087 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1090 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign n_n259 = ( wire3433 ) | ( wire3434 ) | ( wire18316 ) ;
 assign n_n164 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign n_n111 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign wire186 = ( n_n170  &  wire721 ) | ( n_n170  &  wire725 ) ;
 assign n_n5103 = ( n_n47  &  n_n132 ) | ( n_n46  &  wire186 ) ;
 assign wire212 = ( n_n216  &  wire719 ) | ( n_n216  &  wire728 ) ;
 assign n_n5067 = ( n_n41  &  n_n61 ) | ( n_n40  &  wire212 ) ;
 assign wire1096 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign wire208 = ( n_n170  &  wire722 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire715 ) ;
 assign wire591 = ( n_n108  &  wire208 ) | ( n_n108  &  wire148 ) ;
 assign wire515 = ( n_n125  &  n_n177  &  wire725 ) ;
 assign wire657 = ( n_n5743 ) | ( wire4948 ) ;
 assign n_n4424 = ( wire17013 ) | ( wire17014 ) | ( n_n40  &  wire1789 ) ;
 assign wire518 = ( n_n40  &  n_n176 ) | ( n_n41  &  wire69 ) ;
 assign wire653 = ( n_n40  &  wire224 ) | ( n_n40  &  wire57 ) ;
 assign wire694 = ( n_n41  &  wire208 ) | ( n_n41  &  wire148 ) ;
 assign n_n4404 = ( n_n4424 ) | ( wire17018 ) | ( wire17019 ) | ( wire17025 ) ;
 assign wire503 = ( n_n126  &  n_n48  &  n_n220  &  wire104 ) ;
 assign wire666 = ( n_n46  &  wire182 ) | ( n_n47  &  wire150 ) ;
 assign n_n4397 = ( n_n4404 ) | ( wire17049 ) | ( wire17050 ) | ( wire17064 ) ;
 assign n_n4312 = ( wire157  &  n_n18  &  n_n48  &  wire714 ) ;
 assign wire141 = ( n_n216  &  wire721 ) | ( n_n216  &  wire725 ) | ( n_n216  &  wire728 ) ;
 assign wire135 = ( n_n199  &  wire719 ) | ( n_n199  &  wire728 ) ;
 assign n_n4476 = ( n_n41  &  wire219 ) | ( n_n41  &  wire108 ) | ( n_n41  &  wire258 ) ;
 assign n_n4449 = ( n_n31  &  wire168 ) | ( n_n31  &  wire68 ) | ( n_n31  &  wire74 ) ;
 assign n_n4566 = ( n_n157  &  wire714  &  n_n218  &  wire125 ) ;
 assign wire46 = ( n_n177  &  wire720 ) | ( n_n177  &  wire722 ) | ( n_n177  &  wire715 ) ;
 assign wire51 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) ;
 assign n_n1553 = ( n_n41  &  n_n176 ) | ( n_n40  &  wire51 ) ;
 assign wire209 = ( n_n170  &  wire719 ) | ( n_n170  &  wire728 ) ;
 assign n_n5059 = ( n_n41  &  n_n57 ) | ( n_n40  &  wire209 ) ;
 assign n_n5058 = ( n_n41  &  n_n132 ) | ( n_n40  &  wire186 ) ;
 assign wire577 = ( n_n47  &  wire143 ) | ( n_n47  &  wire181 ) ;
 assign wire1115 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire1114 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire1116 = ( wire724  &  n_n177 ) | ( n_n177  &  wire722 ) | ( n_n170  &  wire722 ) ;
 assign wire1117 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1120 = ( wire730  &  n_n156 ) | ( wire726  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire1124 = ( wire164 ) | ( wire358 ) | ( wire243 ) | ( wire17395 ) ;
 assign wire1126 = ( wire723  &  n_n156 ) | ( wire718  &  n_n156 ) | ( wire723  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire1129 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign wire1132 = ( wire303 ) | ( wire321 ) | ( wire326 ) | ( wire327 ) ;
 assign wire1135 = ( wire197 ) | ( wire203 ) | ( wire309 ) | ( wire323 ) ;
 assign wire74 = ( n_n199  &  wire716 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire718 ) ;
 assign wire1136 = ( i_15_  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n199  &  n_n201 ) ;
 assign wire83 = ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign wire384 = ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n177  &  wire715 ) ;
 assign wire1143 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire1145 = ( wire52 ) | ( wire98 ) | ( wire51 ) | ( wire330 ) ;
 assign wire1147 = ( wire276 ) | ( wire211 ) | ( wire271 ) | ( wire19221 ) ;
 assign wire1150 = ( wire142 ) | ( n_n102 ) | ( wire233 ) | ( wire251 ) ;
 assign wire1152 = ( n_n172 ) | ( wire179 ) | ( wire223 ) | ( wire271 ) ;
 assign wire500 = ( n_n17  &  n_n48  &  wire714  &  wire51 ) ;
 assign wire1154 = ( wire52 ) | ( wire63 ) | ( wire276 ) | ( wire211 ) ;
 assign wire1153 = ( n_n183 ) | ( wire184 ) | ( wire246 ) | ( wire254 ) ;
 assign n_n3415 = ( n_n41  &  wire53 ) | ( n_n40  &  n_n77 ) ;
 assign wire1160 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1159 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n7262 = ( (~ i_7_)  &  i_6_  &  n_n48  &  n_n219 ) ;
 assign n_n73 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire718 ) ;
 assign n_n211 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire150 = ( n_n170  &  wire721 ) | ( n_n170  &  wire725 ) | ( n_n170  &  wire728 ) ;
 assign n_n1606 = ( n_n46  &  n_n169 ) | ( n_n47  &  wire57 ) ;
 assign wire1170 = ( n_n176 ) | ( wire224 ) | ( wire250 ) | ( wire100 ) ;
 assign n_n4623 = ( n_n17  &  wire85  &  n_n48  &  wire714 ) ;
 assign n_n3979 = ( wire90  &  n_n40 ) | ( n_n41  &  n_n142 ) ;
 assign wire361 = ( n_n40  &  wire729  &  n_n216 ) | ( n_n40  &  wire726  &  n_n216 ) ;
 assign wire363 = ( n_n41  &  wire729  &  n_n156 ) | ( n_n41  &  wire726  &  n_n156 ) ;
 assign wire426 = ( n_n41  &  wire215 ) | ( n_n41  &  wire720  &  n_n156 ) ;
 assign wire442 = ( n_n41  &  wire155 ) | ( n_n41  &  wire205 ) ;
 assign wire1173 = ( n_n148 ) | ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign wire1174 = ( wire54 ) | ( wire94 ) | ( wire184 ) | ( wire268 ) ;
 assign wire1177 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1176 = ( wire1177 ) | ( wire729  &  n_n156 ) ;
 assign wire1179 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1178 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire377 = ( wire724  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign n_n4247 = ( n_n162  &  n_n157  &  wire714  &  wire158 ) ;
 assign wire655 = ( n_n31  &  n_n216  &  wire725 ) ;
 assign wire1190 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1189 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1188 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) ;
 assign wire1194 = ( wire380 ) | ( wire18986 ) ;
 assign wire136 = ( i_15_  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n213  &  n_n199 ) ;
 assign wire364 = ( i_15_  &  n_n213  &  n_n216 ) | ( (~ i_15_)  &  n_n213  &  n_n216 ) ;
 assign wire1197 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1196 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1195 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign n_n1843 = ( wire18834 ) | ( n_n31  &  wire1197 ) ;
 assign n_n1826 = ( n_n46  &  wire1401 ) | ( n_n47  &  wire1401 ) | ( n_n47  &  wire331 ) ;
 assign wire1200 = ( wire197 ) | ( wire203 ) | ( wire309 ) | ( wire323 ) ;
 assign wire1199 = ( i_8_  &  n_n18  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n18  &  n_n48  &  n_n220 ) ;
 assign n_n1803 = ( n_n1826 ) | ( wire18961 ) | ( wire18962 ) | ( wire18966 ) ;
 assign n_n1824 = ( wire18981 ) | ( n_n46  &  wire1768 ) | ( n_n46  &  wire18980 ) ;
 assign wire1201 = ( wire312 ) | ( wire326 ) | ( wire327 ) | ( wire331 ) ;
 assign wire1205 = ( wire261 ) | ( wire264 ) | ( wire375 ) | ( wire19001 ) ;
 assign wire62 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) ;
 assign wire1207 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1211 = ( wire92 ) | ( wire232 ) | ( wire19413 ) | ( wire19414 ) ;
 assign n_n1542 = ( n_n41  &  n_n148 ) | ( n_n40  &  wire60 ) ;
 assign n_n4641 = ( n_n46  &  n_n214 ) | ( n_n47  &  wire70 ) ;
 assign wire693 = ( n_n47  &  wire68 ) | ( n_n47  &  wire74 ) ;
 assign wire1214 = ( wire86 ) | ( wire162 ) | ( wire169 ) | ( wire19320 ) ;
 assign wire1216 = ( n_n155 ) | ( wire148 ) | ( wire274 ) | ( wire277 ) ;
 assign wire154 = ( wire723  &  n_n216 ) | ( n_n216  &  wire730 ) | ( n_n216  &  wire727 ) ;
 assign wire1218 = ( i_15_  &  n_n216  &  n_n205 ) | ( (~ i_15_)  &  n_n216  &  n_n205 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign n_n369 = ( wire2083 ) | ( n_n34  &  wire154 ) | ( n_n34  &  wire1218 ) ;
 assign wire335 = ( n_n216  &  wire720 ) | ( n_n216  &  wire727 ) ;
 assign wire747 = ( (~ i_7_)  &  i_8_  &  (~ i_6_) ) ;
 assign wire100 = ( n_n177  &  wire722 ) | ( n_n177  &  wire727 ) | ( n_n177  &  wire715 ) ;
 assign wire153 = ( n_n199  &  wire721 ) | ( n_n199  &  wire725 ) ;
 assign wire234 = ( wire723  &  n_n149 ) | ( wire716  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire652 = ( n_n46  &  wire218 ) | ( n_n47  &  wire141 ) ;
 assign n_n4518 = ( n_n212  &  wire143 ) | ( n_n212  &  wire154 ) | ( n_n212  &  wire47 ) ;
 assign wire1224 = ( wire168 ) | ( wire68 ) | ( wire151 ) | ( wire74 ) ;
 assign wire125 = ( n_n216  &  wire719 ) | ( n_n216  &  wire721 ) | ( n_n216  &  wire728 ) ;
 assign n_n7266 = ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n218 ) ;
 assign wire1229 = ( n_n161  &  n_n48  &  n_n159 ) | ( n_n124  &  n_n48  &  n_n159 ) ;
 assign n_n3054 = ( wire18706 ) | ( wire18707 ) | ( n_n92  &  wire1229 ) ;
 assign wire131 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) | ( wire724  &  n_n177 ) ;
 assign n_n2770 = ( wire137  &  n_n197 ) | ( n_n197  &  wire146 ) | ( n_n197  &  wire131 ) ;
 assign wire1234 = ( wire116 ) | ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire412 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) ;
 assign wire1239 = ( i_15_  &  n_n191  &  n_n204 ) | ( i_15_  &  n_n191  &  n_n201 ) | ( (~ i_15_)  &  n_n191  &  n_n201 ) ;
 assign n_n1913 = ( wire18938 ) | ( wire18939 ) ;
 assign n_n3638 = ( wire139  &  n_n157  &  wire714  &  n_n218 ) ;
 assign wire1242 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1244 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1243 = ( i_8_  &  n_n16  &  n_n220  &  n_n218 ) | ( (~ i_8_)  &  n_n16  &  n_n220  &  n_n218 ) ;
 assign wire1246 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign n_n1811 = ( n_n31  &  wire1246 ) | ( n_n30  &  wire1246 ) | ( n_n30  &  wire309 ) ;
 assign wire1247 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1251 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1255 = ( wire98 ) | ( wire63 ) | ( wire206 ) | ( wire330 ) ;
 assign wire1257 = ( n_n177  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign n_n817 = ( n_n974 ) | ( wire4869 ) | ( n_n38  &  wire104 ) ;
 assign wire167 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n209 ) ;
 assign n_n799 = ( wire2329 ) | ( wire2331 ) | ( wire19480 ) | ( wire19481 ) ;
 assign wire1259 = ( wire320 ) | ( wire19660 ) ;
 assign wire1261 = ( wire98 ) | ( wire195 ) | ( wire320 ) | ( wire19663 ) ;
 assign wire1260 = ( n_n118 ) | ( wire104 ) | ( wire54 ) | ( wire195 ) ;
 assign wire1263 = ( wire182 ) | ( n_n177  &  wire725 ) ;
 assign wire449 = ( n_n31  &  wire134 ) | ( n_n31  &  wire156 ) ;
 assign wire656 = ( n_n31  &  wire176 ) | ( n_n31  &  wire123 ) ;
 assign wire686 = ( wire132  &  n_n47 ) | ( n_n47  &  wire126 ) ;
 assign wire1271 = ( wire132 ) | ( wire149 ) | ( wire147 ) | ( wire126 ) ;
 assign n_n4692 = ( n_n200  &  n_n220  &  n_n218  &  wire46 ) ;
 assign wire1277 = ( i_8_  &  n_n162  &  n_n18  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n18  &  n_n220 ) ;
 assign wire175 = ( i_15_  &  n_n213  &  n_n156 ) | ( (~ i_15_)  &  n_n213  &  n_n156 ) ;
 assign wire383 = ( i_15_  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n213  &  n_n177 ) ;
 assign wire1279 = ( i_15_  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n191  &  n_n201 ) ;
 assign wire1281 = ( n_n137 ) | ( wire302 ) | ( wire316 ) | ( wire403 ) ;
 assign wire1285 = ( wire312 ) | ( wire326 ) | ( wire327 ) | ( wire331 ) ;
 assign wire69 = ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) ;
 assign wire276 = ( n_n184  &  wire720 ) | ( n_n184  &  wire727 ) | ( n_n184  &  wire715 ) ;
 assign wire1287 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire1286 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire473 = ( n_n115  &  n_n32 ) | ( n_n33  &  n_n137 ) ;
 assign wire1290 = ( wire179 ) | ( wire223 ) | ( wire239 ) | ( wire19253 ) ;
 assign wire1289 = ( wire155 ) | ( wire227 ) | ( wire232 ) | ( wire19250 ) ;
 assign wire1292 = ( wire155 ) | ( wire227 ) | ( wire232 ) | ( wire19260 ) ;
 assign wire557 = ( n_n212  &  wire147 ) | ( n_n212  &  wire126 ) ;
 assign wire1294 = ( n_n77 ) | ( wire148 ) | ( wire274 ) | ( wire277 ) ;
 assign wire1293 = ( wire53 ) | ( wire179 ) | ( wire223 ) | ( wire239 ) ;
 assign n_n1566 = ( n_n43  &  n_n115 ) | ( n_n42  &  wire65 ) ;
 assign wire88 = ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) ;
 assign wire1295 = ( n_n216  &  wire717 ) | ( n_n216  &  wire718 ) | ( n_n216  &  wire727 ) ;
 assign n_n1575 = ( n_n43  &  n_n183 ) | ( n_n42  &  wire62 ) ;
 assign wire1297 = ( wire184 ) | ( wire246 ) | ( wire254 ) | ( wire349 ) ;
 assign wire124 = ( n_n184  &  wire720 ) | ( n_n184  &  wire722 ) | ( n_n184  &  wire715 ) ;
 assign wire1302 = ( n_n72 ) | ( wire199 ) | ( wire290 ) | ( wire19464 ) ;
 assign wire1305 = ( wire98 ) | ( wire195 ) | ( wire320 ) | ( wire19469 ) ;
 assign wire1311 = ( wire329 ) | ( wire726  &  n_n170 ) ;
 assign wire80 = ( n_n177  &  wire719 ) | ( n_n177  &  wire728 ) ;
 assign n_n2859 = ( n_n123  &  n_n63 ) | ( n_n125  &  wire171 ) ;
 assign n_n4657 = ( wire182  &  n_n126  &  n_n220  &  n_n218 ) ;
 assign wire160 = ( n_n191  &  wire721 ) | ( n_n191  &  wire725 ) ;
 assign wire78 = ( n_n177  &  wire721 ) | ( n_n177  &  wire725 ) ;
 assign wire651 = ( wire157  &  n_n47 ) | ( n_n46  &  wire174 ) ;
 assign n_n3570 = ( n_n108  &  wire176 ) | ( n_n108  &  wire123 ) | ( n_n108  &  wire156 ) ;
 assign n_n3573 = ( wire137  &  n_n108 ) | ( n_n108  &  wire146 ) | ( n_n108  &  wire46 ) ;
 assign wire1319 = ( wire137 ) | ( wire146 ) | ( wire46 ) | ( wire131 ) ;
 assign n_n3823 = ( n_n3573 ) | ( wire4182 ) | ( n_n101  &  wire1319 ) ;
 assign wire1321 = ( wire214 ) | ( n_n134 ) | ( wire222 ) | ( wire174 ) ;
 assign wire537 = ( wire85  &  n_n40 ) | ( wire142  &  n_n40 ) ;
 assign wire1326 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign n_n5070 = ( wire214  &  n_n41 ) | ( n_n40  &  n_n140 ) ;
 assign wire217 = ( n_n184  &  wire719 ) | ( n_n184  &  wire721 ) | ( n_n184  &  wire728 ) ;
 assign n_n3037 = ( wire3496 ) | ( wire3497 ) | ( wire18272 ) | ( wire18273 ) ;
 assign wire469 = ( wire724  &  n_n177 ) | ( n_n177  &  wire717 ) ;
 assign wire1331 = ( wire53 ) | ( wire117 ) | ( wire281 ) | ( wire294 ) ;
 assign wire115 = ( wire726  &  n_n149 ) | ( wire724  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire673 = ( n_n40  &  wire247 ) | ( n_n41  &  wire218 ) ;
 assign n_n3029 = ( n_n3037 ) | ( wire3484 ) | ( wire18283 ) | ( wire18288 ) ;
 assign wire1336 = ( wire157 ) | ( wire186 ) | ( wire209 ) | ( wire174 ) ;
 assign wire173 = ( n_n149  &  wire721 ) | ( n_n149  &  wire725 ) ;
 assign n_n2733 = ( n_n33  &  wire173 ) | ( n_n33  &  n_n149  &  wire719 ) ;
 assign wire1341 = ( i_15_  &  n_n213  &  n_n216 ) | ( (~ i_15_)  &  n_n213  &  n_n216 ) | ( (~ i_15_)  &  n_n216  &  n_n209 ) ;
 assign wire378 = ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire1345 = ( i_8_  &  n_n162  &  n_n16  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n16  &  n_n220 ) ;
 assign wire1343 = ( n_n199  &  wire720 ) | ( n_n199  &  wire727 ) | ( n_n199  &  wire715 ) ;
 assign wire1342 = ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1347 = ( wire48 ) | ( wire167 ) | ( wire124 ) | ( wire165 ) ;
 assign wire1346 = ( wire167 ) | ( wire124 ) | ( wire165 ) | ( wire280 ) ;
 assign n_n784 = ( wire2302 ) | ( wire2303 ) | ( wire19510 ) ;
 assign wire629 = ( n_n200  &  n_n220  &  n_n218  &  wire47 ) ;
 assign n_n752 = ( n_n784 ) | ( wire2308 ) | ( wire19506 ) | ( wire19516 ) ;
 assign wire1354 = ( wire166 ) | ( wire269 ) | ( wire275 ) | ( wire278 ) ;
 assign wire1357 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire244 = ( wire723  &  n_n156 ) | ( wire720  &  n_n156 ) | ( n_n156  &  wire727 ) ;
 assign wire1363 = ( wire140 ) | ( wire244 ) | ( wire282 ) | ( wire283 ) ;
 assign wire1366 = ( wire296 ) | ( wire262 ) | ( wire332 ) | ( wire342 ) ;
 assign wire1367 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire479 = ( n_n125  &  wire155 ) | ( n_n125  &  n_n155 ) | ( n_n125  &  wire215 ) ;
 assign wire222 = ( n_n191  &  wire719 ) | ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) ;
 assign n_n3525 = ( wire137  &  n_n36 ) | ( n_n36  &  wire146 ) | ( n_n36  &  wire131 ) ;
 assign wire1375 = ( n_n177  &  n_n220  &  n_n111 ) | ( n_n156  &  n_n220  &  n_n111 ) ;
 assign n_n3561 = ( n_n47  &  wire52 ) | ( n_n47  &  wire63 ) | ( n_n47  &  wire48 ) ;
 assign n_n3825 = ( n_n3578 ) | ( wire4067 ) | ( wire17716 ) | ( wire17717 ) ;
 assign wire1378 = ( wire52 ) | ( wire129 ) | ( wire63 ) | ( wire48 ) ;
 assign n_n3180 = ( wire3496 ) | ( wire3497 ) | ( wire18454 ) | ( wire18455 ) ;
 assign wire1381 = ( wire132 ) | ( wire149 ) | ( wire147 ) | ( wire126 ) ;
 assign wire1383 = ( wire55 ) | ( wire158 ) | ( wire133 ) | ( wire127 ) ;
 assign n_n3170 = ( n_n3180 ) | ( wire18461 ) | ( wire18462 ) | ( wire18469 ) ;
 assign wire1386 = ( wire168 ) | ( wire68 ) | ( wire151 ) | ( wire74 ) ;
 assign wire1390 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) ;
 assign wire1389 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire730 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire730 ) ;
 assign wire170 = ( wire729  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire1395 = ( wire247 ) | ( wire125 ) | ( wire160 ) | ( wire18534 ) ;
 assign wire1401 = ( wire292 ) | ( wire311 ) | ( wire317 ) | ( wire319 ) ;
 assign wire1404 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1405 = ( n_n191  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n191  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire219 = ( n_n199  &  wire722 ) | ( n_n199  &  wire727 ) | ( n_n199  &  wire715 ) ;
 assign n_n371 = ( wire712 ) | ( wire2080 ) | ( n_n34  &  n_n198 ) ;
 assign wire1416 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1415 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1414 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire759 = ( n_n149  &  n_n220  &  n_n111 ) ;
 assign wire1417 = ( n_n184  &  wire719 ) | ( n_n184  &  wire725 ) | ( n_n184  &  wire728 ) ;
 assign wire645 = ( n_n40  &  wire155 ) | ( n_n40  &  wire205 ) ;
 assign wire664 = ( n_n41  &  wire234 ) | ( n_n41  &  wire84 ) ;
 assign wire171 = ( n_n191  &  wire719 ) | ( n_n191  &  wire728 ) ;
 assign wire394 = ( n_n125  &  wire224 ) | ( n_n125  &  wire250 ) | ( n_n125  &  wire57 ) ;
 assign wire1420 = ( wire240 ) | ( wire187 ) | ( wire210 ) | ( wire17741 ) ;
 assign n_n3592 = ( n_n125  &  wire240 ) | ( n_n125  &  wire187 ) | ( n_n125  &  wire210 ) ;
 assign n_n3834 = ( wire648 ) | ( wire681 ) | ( wire17766 ) | ( wire17767 ) ;
 assign n_n3833 = ( n_n2770 ) | ( n_n4692 ) | ( n_n3601 ) | ( wire504 ) ;
 assign wire1425 = ( n_n51 ) | ( wire245 ) | ( wire122 ) | ( wire144 ) ;
 assign wire1424 = ( n_n128 ) | ( wire122 ) | ( wire144 ) | ( wire152 ) ;
 assign wire1427 = ( n_n124  &  n_n48  &  n_n159 ) | ( n_n48  &  n_n35  &  n_n159 ) ;
 assign wire1432 = ( n_n65 ) | ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign wire1436 = ( wire90 ) | ( wire175 ) | ( wire198 ) | ( wire19099 ) ;
 assign wire1437 = ( wire48 ) | ( wire167 ) | ( wire124 ) | ( wire165 ) ;
 assign n_n772 = ( wire19599 ) | ( wire19600 ) | ( n_n46  &  wire1437 ) ;
 assign wire1440 = ( n_n60 ) | ( wire235 ) | ( wire236 ) | ( wire413 ) ;
 assign wire1444 = ( wire166 ) | ( wire269 ) | ( wire275 ) | ( wire278 ) ;
 assign n_n326 = ( n_n46  &  wire1444 ) | ( n_n47  &  wire1444 ) | ( n_n47  &  wire325 ) ;
 assign wire1446 = ( wire244 ) | ( wire235 ) | ( wire236 ) | ( wire19701 ) ;
 assign wire86 = ( wire729  &  n_n216 ) | ( wire726  &  n_n216 ) ;
 assign wire240 = ( wire724  &  n_n191 ) | ( n_n191  &  wire717 ) | ( n_n191  &  wire718 ) ;
 assign wire497 = ( n_n41  &  n_n190 ) | ( n_n41  &  wire187 ) | ( n_n41  &  wire210 ) ;
 assign wire1450 = ( n_n190 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire636 = ( wire157  &  n_n36 ) | ( n_n34  &  wire174 ) ;
 assign n_n3578 = ( n_n108  &  wire143 ) | ( n_n108  &  wire181 ) | ( n_n108  &  wire154 ) ;
 assign wire47 = ( n_n216  &  wire720 ) | ( n_n216  &  wire722 ) | ( n_n216  &  wire715 ) ;
 assign wire1459 = ( wire120 ) | ( wire179 ) | ( wire324 ) | ( wire18253 ) ;
 assign wire1463 = ( (~ i_7_)  &  i_6_ ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n2956 = ( n_n7254 ) | ( wire551 ) | ( wire4223 ) | ( wire17588 ) ;
 assign wire1465 = ( wire176 ) | ( wire134 ) | ( wire123 ) | ( wire156 ) ;
 assign n_n3601 = ( n_n212  &  wire134 ) | ( n_n212  &  wire123 ) | ( n_n212  &  wire156 ) ;
 assign wire197 = ( i_15_  &  n_n213  &  n_n216 ) | ( (~ i_15_)  &  n_n213  &  n_n216 ) | ( i_15_  &  n_n216  &  n_n207 ) ;
 assign wire1470 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1469 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire401 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1477 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1476 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1480 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire1479 = ( n_n177  &  wire720 ) | ( n_n170  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n170  &  wire727 ) ;
 assign wire1478 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1483 = ( n_n164 ) | ( wire110 ) | ( wire336 ) | ( wire19895 ) ;
 assign wire1482 = ( n_n185 ) | ( wire161 ) | ( wire336 ) | ( wire19895 ) ;
 assign n_n225 = ( n_n231 ) | ( wire16886 ) | ( wire736  &  n_n162 ) ;
 assign n_n5021 = ( n_n108  &  n_n190 ) | ( n_n101  &  wire86 ) ;
 assign wire128 = ( n_n184  &  wire723 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire727 ) ;
 assign wire565 = ( n_n197  &  wire134 ) | ( n_n197  &  wire156 ) ;
 assign wire1488 = ( wire144 ) | ( n_n156  &  wire721 ) | ( n_n156  &  wire725 ) ;
 assign wire579 = ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) ;
 assign wire648 = ( wire137  &  n_n212 ) | ( n_n212  &  wire46 ) ;
 assign wire681 = ( n_n197  &  wire63 ) | ( n_n197  &  wire48 ) ;
 assign wire1489 = ( wire137 ) | ( wire146 ) | ( wire46 ) ;
 assign wire504 = ( n_n212  &  wire146 ) | ( n_n212  &  wire131 ) ;
 assign n_n3800 = ( wire449 ) | ( wire656 ) | ( wire3985 ) | ( wire17787 ) ;
 assign n_n3514 = ( n_n31  &  wire52 ) | ( n_n31  &  wire63 ) | ( n_n31  &  wire48 ) ;
 assign wire1491 = ( wire63 ) | ( wire143 ) | ( wire48 ) | ( wire154 ) ;
 assign n_n3802 = ( n_n3514 ) | ( wire17793 ) | ( n_n30  &  wire1491 ) ;
 assign n_n3511 = ( n_n31  &  wire137 ) | ( n_n31  &  wire146 ) | ( n_n31  &  wire131 ) ;
 assign wire690 = ( n_n30  &  wire137 ) | ( n_n30  &  wire46 ) ;
 assign wire1493 = ( wire52 ) | ( wire129 ) | ( wire63 ) | ( wire48 ) ;
 assign wire1496 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1495 = ( n_n65 ) | ( wire95 ) | ( n_n89 ) | ( wire87 ) ;
 assign wire1498 = ( n_n82 ) | ( wire230 ) | ( wire260 ) | ( wire373 ) ;
 assign wire1497 = ( n_n70 ) | ( wire230 ) | ( wire347 ) | ( wire352 ) ;
 assign wire1500 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1499 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire1503 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1504 = ( wire133 ) | ( wire60 ) | ( wire127 ) | ( wire227 ) ;
 assign wire1507 = ( wire210 ) | ( wire349 ) | ( wire357 ) | ( wire19328 ) ;
 assign wire1510 = ( wire314 ) | ( n_n184  &  wire726 ) ;
 assign wire1513 = ( n_n178 ) | ( wire259 ) | ( wire337 ) | ( wire19831 ) ;
 assign wire1512 = ( n_n202 ) | ( wire337 ) | ( wire338 ) | ( wire19831 ) ;
 assign wire689 = ( wire157  &  n_n212 ) | ( n_n197  &  wire174 ) ;
 assign wire1519 = ( wire172 ) | ( wire51 ) | ( wire240 ) | ( wire210 ) ;
 assign wire1520 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire1523 = ( wire145 ) | ( n_n151 ) | ( n_n186 ) | ( wire370 ) ;
 assign n_n3176 = ( wire707 ) | ( wire18367 ) | ( n_n2  &  wire1523 ) ;
 assign wire1524 = ( i_5_  &  (~ i_3_)  &  i_4_  &  n_n19 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n19 ) | ( i_5_  &  (~ i_3_)  &  (~ i_4_)  &  n_n19 ) | ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_)  &  n_n19 ) ;
 assign wire1527 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire315 = ( wire729  &  n_n149 ) | ( wire726  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire1537 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire1539 = ( wire155 ) | ( wire232 ) | ( wire19442 ) | ( wire19443 ) ;
 assign n_n1163 = ( wire19446 ) | ( n_n30  &  wire1539 ) ;
 assign wire348 = ( i_15_  &  n_n191  &  n_n205 ) | ( (~ i_15_)  &  n_n191  &  n_n205 ) ;
 assign wire385 = ( i_15_  &  n_n199  &  n_n205 ) | ( (~ i_15_)  &  n_n199  &  n_n205 ) ;
 assign wire675 = ( n_n33  &  wire129 ) | ( n_n33  &  wire150 ) ;
 assign wire1544 = ( wire137 ) | ( n_n84 ) | ( wire146 ) | ( wire46 ) ;
 assign wire270 = ( wire729  &  n_n191 ) | ( n_n191  &  wire717 ) | ( n_n191  &  wire730 ) ;
 assign wire1553 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire1556 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1558 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire1560 = ( n_n199  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire1562 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire1568 = ( n_n202 ) | ( wire295 ) | ( wire333 ) | ( wire19882 ) ;
 assign wire1570 = ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) | ( i_15_  &  n_n156  &  n_n215 ) ;
 assign wire560 = ( n_n47  &  wire176 ) | ( n_n47  &  wire123 ) ;
 assign wire688 = ( n_n46  &  wire123 ) | ( n_n46  &  wire156 ) ;
 assign wire432 = ( n_n36  &  wire154 ) | ( n_n36  &  wire47 ) ;
 assign wire1576 = ( wire116 ) | ( wire198 ) | ( wire289 ) | ( wire18426 ) ;
 assign n_n3555 = ( n_n47  &  wire158 ) | ( n_n47  &  wire133 ) | ( n_n47  &  wire127 ) ;
 assign wire1580 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1579 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1578 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire1581 = ( wire385 ) | ( wire108 ) | ( wire19318 ) ;
 assign wire1582 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire1587 = ( wire335 ) | ( wire295 ) | ( wire333 ) | ( wire19835 ) ;
 assign wire1590 = ( wire314 ) | ( wire333 ) | ( wire338 ) | ( wire19901 ) ;
 assign wire1592 = ( n_n150 ) | ( wire248 ) | ( wire249 ) | ( wire19905 ) ;
 assign wire1595 = ( wire132 ) | ( wire46 ) | ( wire121 ) | ( wire280 ) ;
 assign wire57 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) ;
 assign wire434 = ( n_n39  &  n_n156  &  wire728 ) | ( n_n39  &  n_n149  &  wire728 ) ;
 assign wire538 = ( n_n125  &  wire108 ) | ( n_n125  &  wire258 ) ;
 assign wire539 = ( n_n125  &  wire180 ) | ( n_n125  &  wire86 ) ;
 assign wire1601 = ( wire17918 ) | ( wire17919 ) | ( wire17920 ) | ( wire17921 ) ;
 assign n_n2777 = ( n_n212  &  wire139 ) | ( n_n212  &  wire124 ) | ( n_n212  &  wire128 ) ;
 assign wire1602 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire607 = ( n_n34  &  wire146 ) | ( n_n34  &  wire131 ) ;
 assign wire640 = ( n_n34  &  wire63 ) | ( n_n34  &  wire48 ) ;
 assign wire584 = ( wire132  &  n_n36 ) | ( n_n36  &  wire126 ) ;
 assign wire1605 = ( wire107 ) | ( wire339 ) | ( wire187 ) | ( wire19523 ) ;
 assign wire1613 = ( wire335 ) | ( wire295 ) | ( wire333 ) | ( wire19767 ) ;
 assign wire1617 = ( wire99 ) | ( wire282 ) | ( wire283 ) | ( wire325 ) ;
 assign n_n3485 = ( wire674 ) | ( n_n3889 ) | ( wire686 ) | ( wire18028 ) ;
 assign wire698 = ( n_n125  &  wire208 ) | ( n_n125  &  wire148 ) ;
 assign n_n3467 = ( wire449 ) | ( wire656 ) | ( wire3820 ) | ( wire17926 ) ;
 assign n_n3510 = ( n_n31  &  wire132 ) | ( n_n31  &  wire147 ) | ( n_n31  &  wire126 ) ;
 assign wire1625 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire578 = ( n_n197  &  wire147 ) | ( n_n197  &  wire126 ) ;
 assign n_n2754 = ( wire3177 ) | ( wire18581 ) | ( wire18582 ) | ( wire18583 ) ;
 assign wire1627 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign n_n2630 = ( wire17880 ) | ( wire17881 ) | ( n_n34  &  wire1627 ) ;
 assign wire642 = ( n_n36  &  wire63 ) | ( n_n36  &  wire48 ) ;
 assign wire1628 = ( wire124 ) | ( wire47 ) | ( wire165 ) | ( wire322 ) ;
 assign wire407 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1630 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1632 = ( wire55 ) | ( wire134 ) | ( wire163 ) | ( wire194 ) ;
 assign n_n765 = ( n_n41  &  wire1632 ) | ( n_n40  &  wire1632 ) | ( n_n40  &  wire280 ) ;
 assign wire635 = ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) ;
 assign wire1633 = ( wire720  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign n_n745 = ( n_n817 ) | ( wire19556 ) | ( wire19557 ) | ( wire19560 ) ;
 assign wire346 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) ;
 assign wire1636 = ( n_n60 ) | ( wire235 ) | ( wire236 ) | ( wire19796 ) ;
 assign wire1640 = ( wire296 ) | ( wire262 ) | ( wire332 ) | ( wire342 ) ;
 assign wire1639 = ( i_8_  &  n_n18  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n18  &  n_n48  &  n_n220 ) ;
 assign n_n302 = ( n_n326 ) | ( wire19786 ) | ( wire19787 ) | ( wire19793 ) ;
 assign wire1641 = ( wire282 ) | ( wire283 ) | ( wire325 ) | ( wire354 ) ;
 assign n_n301 = ( wire2017 ) | ( wire19799 ) | ( wire19812 ) ;
 assign n_n3473 = ( wire458 ) | ( n_n3525 ) | ( wire584 ) | ( wire17960 ) ;
 assign wire1648 = ( wire211 ) | ( wire242 ) | ( wire272 ) | ( wire17944 ) ;
 assign n_n3470 = ( wire17947 ) | ( wire17948 ) | ( n_n32  &  wire1648 ) ;
 assign n_n2642 = ( n_n36  &  wire158 ) | ( n_n36  &  wire133 ) | ( n_n36  &  wire127 ) ;
 assign wire1649 = ( n_n138 ) | ( n_n63 ) | ( wire135 ) | ( wire153 ) ;
 assign wire1655 = ( wire209 ) | ( wire217 ) | ( wire174 ) | ( wire18611 ) ;
 assign wire1658 = ( i_8_  &  n_n162  &  n_n18  &  n_n220 ) | ( (~ i_8_)  &  n_n162  &  n_n18  &  n_n220 ) ;
 assign n_n768 = ( n_n832 ) | ( wire2232 ) | ( wire2233 ) | ( wire19569 ) ;
 assign wire1659 = ( wire132 ) | ( wire46 ) | ( wire121 ) | ( wire280 ) ;
 assign n_n746 = ( n_n768 ) | ( wire2242 ) | ( wire2243 ) | ( wire19574 ) ;
 assign wire697 = ( n_n43  &  n_n191  &  wire720 ) ;
 assign wire1668 = ( i_8_  &  n_n18  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n18  &  n_n48  &  n_n220 ) ;
 assign wire1666 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign n_n304 = ( n_n333 ) | ( wire19846 ) | ( wire19847 ) | ( wire19859 ) ;
 assign n_n3501 = ( wire579 ) | ( wire648 ) | ( n_n2777 ) | ( wire18122 ) ;
 assign n_n3500 = ( wire557 ) | ( n_n3601 ) | ( wire504 ) | ( wire18125 ) ;
 assign wire1674 = ( wire55 ) | ( wire163 ) | ( wire194 ) | ( wire19577 ) ;
 assign n_n834 = ( wire2218 ) | ( wire19584 ) | ( n_n43  &  n_n190 ) ;
 assign wire107 = ( n_n184  &  wire722 ) | ( n_n184  &  wire727 ) | ( n_n184  &  wire715 ) ;
 assign wire1675 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign n_n769 = ( n_n834 ) | ( wire19587 ) | ( wire19588 ) | ( wire19591 ) ;
 assign wire1679 = ( wire132 ) | ( wire121 ) | ( wire280 ) ;
 assign n_n747 = ( n_n769 ) | ( wire19582 ) | ( wire19583 ) | ( wire19596 ) ;
 assign wire1684 = ( wire415 ) | ( wire269 ) | ( wire275 ) | ( wire342 ) ;
 assign wire296 = ( n_n199  &  wire723 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire727 ) ;
 assign wire1689 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire696 = ( n_n41  &  wire224 ) | ( n_n41  &  wire250 ) ;
 assign n_n3542 = ( n_n41  &  wire224 ) | ( n_n41  &  wire250 ) | ( n_n41  &  wire100 ) ;
 assign n_n3482 = ( wire683 ) | ( wire3767 ) | ( wire17979 ) | ( wire17980 ) ;
 assign n_n3487 = ( n_n3562 ) | ( wire481 ) | ( wire577 ) | ( wire18032 ) ;
 assign n_n3460 = ( n_n3485 ) | ( n_n3487 ) | ( wire18039 ) ;
 assign wire1695 = ( wire143 ) | ( wire181 ) | ( wire154 ) | ( wire47 ) ;
 assign wire1704 = ( i_8_  &  n_n17  &  n_n48  &  n_n220 ) | ( (~ i_8_)  &  n_n17  &  n_n48  &  n_n220 ) ;
 assign wire1706 = ( wire320 ) | ( wire19624 ) ;
 assign wire1709 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1708 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire1707 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign n_n748 = ( wire2182 ) | ( wire19614 ) | ( wire19617 ) | ( wire19619 ) ;
 assign wire1717 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1716 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire1720 = ( i_15_  &  n_n191  &  n_n205 ) | ( (~ i_15_)  &  n_n191  &  n_n205 ) | ( i_15_  &  n_n191  &  n_n215 ) | ( (~ i_15_)  &  n_n191  &  n_n215 ) ;
 assign wire1723 = ( wire107 ) | ( wire211 ) | ( wire272 ) | ( wire18657 ) ;
 assign wire606 = ( wire137  &  n_n34 ) | ( n_n34  &  wire46 ) ;
 assign wire1730 = ( wire129 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign wire1729 = ( wire130 ) | ( wire139 ) | ( wire124 ) | ( wire128 ) ;
 assign n_n2626 = ( n_n2642 ) | ( wire17896 ) | ( wire17897 ) | ( wire17898 ) ;
 assign wire263 = ( n_n216  &  wire724 ) | ( n_n216  &  wire717 ) | ( n_n216  &  wire730 ) ;
 assign wire1735 = ( wire261 ) | ( wire264 ) | ( wire375 ) | ( wire19013 ) ;
 assign wire165 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n209 ) ;
 assign wire1739 = ( wire132 ) | ( wire55 ) | ( wire121 ) | ( wire163 ) ;
 assign wire1738 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire1741 = ( n_n84 ) | ( wire279 ) | ( wire54 ) | ( wire195 ) ;
 assign wire1740 = ( wire53 ) | ( n_n118 ) | ( wire195 ) | ( wire237 ) ;
 assign wire1743 = ( wire118 ) | ( wire279 ) | ( wire199 ) | ( wire19633 ) ;
 assign wire1742 = ( n_n72 ) | ( wire118 ) | ( wire59 ) | ( wire290 ) ;
 assign n_n333 = ( wire1946 ) | ( wire1949 ) | ( wire1950 ) | ( wire19854 ) ;
 assign wire256 = ( n_n184  &  wire721 ) | ( n_n184  &  wire725 ) ;
 assign wire1748 = ( wire68 ) | ( wire151 ) | ( wire74 ) | ( wire47 ) ;
 assign wire1747 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_ ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_) ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n_n3492 = ( n_n3578 ) | ( wire18044 ) | ( n_n108  &  wire1748 ) ;
 assign n_n3491 = ( n_n108  &  wire18049 ) | ( n_n108  &  wire18050 ) | ( n_n108  &  wire18051 ) ;
 assign wire1751 = ( wire381 ) | ( n_n130 ) | ( wire186 ) | ( wire209 ) ;
 assign n_n3462 = ( n_n3492 ) | ( n_n3491 ) | ( wire18057 ) | ( wire18058 ) ;
 assign n_n3489 = ( n_n3570 ) | ( n_n108  &  wire18063 ) | ( n_n108  &  wire18064 ) ;
 assign n_n3451 = ( n_n3460 ) | ( n_n3462 ) | ( wire18078 ) ;
 assign wire1754 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1753 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire1756 = ( wire237 ) | ( wire19630 ) ;
 assign wire1758 = ( n_n84 ) | ( wire279 ) | ( wire237 ) | ( wire19654 ) ;
 assign wire1761 = ( n_n171 ) | ( wire329 ) | ( wire336 ) | ( wire19856 ) ;
 assign wire1766 = ( n_n137 ) | ( wire302 ) | ( wire316 ) | ( wire18978 ) ;
 assign wire1775 = ( wire111 ) | ( wire291 ) | ( wire297 ) | ( wire19672 ) ;
 assign wire1779 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1778 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1777 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire1780 = ( i_15_  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n205  &  n_n149 ) ;
 assign n_n2684 = ( wire697 ) | ( wire3403 ) | ( wire18342 ) | ( wire18345 ) ;
 assign wire1782 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign wire1786 = ( wire51 ) | ( wire240 ) | ( wire187 ) | ( wire210 ) ;
 assign n_n1801 = ( wire2713 ) | ( wire19021 ) | ( wire19023 ) ;
 assign wire1789 = ( n_n169 ) | ( wire208 ) | ( wire225 ) | ( wire148 ) ;
 assign n_n4419 = ( wire4974 ) | ( wire16952 ) | ( wire16953 ) | ( wire16954 ) ;
 assign wire1791 = ( n_n138 ) | ( n_n63 ) | ( wire135 ) | ( wire153 ) ;
 assign wire1794 = ( n_n189 ) | ( wire202 ) | ( wire307 ) | ( wire17339 ) ;
 assign n_n4399 = ( wire17149 ) | ( wire17150 ) ;
 assign wire1807 = ( wire160 ) | ( wire171 ) | ( wire242 ) | ( wire18004 ) ;
 assign wire1809 = ( n_n103 ) | ( wire291 ) | ( wire297 ) | ( wire19500 ) ;
 assign wire225 = ( wire724  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire718 ) ;
 assign wire1811 = ( wire381 ) | ( wire186 ) | ( wire209 ) | ( wire18007 ) ;
 assign wire1812 = ( wire218 ) | ( wire60 ) | ( wire220 ) | ( wire18014 ) ;
 assign wire1814 = ( wire209 ) | ( wire217 ) | ( wire174 ) | ( wire17903 ) ;
 assign wire49 = ( n_n216  &  wire721 ) | ( n_n216  &  wire728 ) ;
 assign wire50 = ( wire717  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire54 = ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) ;
 assign wire56 = ( n_n216  &  wire717 ) | ( n_n216  &  wire718 ) ;
 assign wire72 = ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire75 = ( wire717  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire79 = ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign wire82 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire84 = ( wire722  &  n_n149 ) | ( n_n149  &  wire727 ) | ( n_n149  &  wire715 ) ;
 assign wire87 = ( n_n191  &  wire717 ) | ( n_n191  &  wire730 ) ;
 assign wire92 = ( n_n199  &  wire721 ) | ( n_n199  &  wire728 ) ;
 assign wire94 = ( n_n184  &  wire726 ) | ( n_n184  &  wire724 ) | ( n_n184  &  wire717 ) ;
 assign wire99 = ( n_n177  &  wire730 ) | ( n_n177  &  wire718 ) ;
 assign wire108 = ( n_n199  &  wire723 ) | ( n_n199  &  wire716 ) | ( n_n199  &  wire730 ) ;
 assign wire110 = ( wire720  &  n_n156 ) | ( n_n156  &  wire727 ) ;
 assign wire116 = ( wire726  &  n_n156 ) | ( wire724  &  n_n156 ) | ( wire717  &  n_n156 ) ;
 assign wire117 = ( wire726  &  n_n170 ) | ( wire724  &  n_n170 ) | ( n_n170  &  wire717 ) ;
 assign wire120 = ( wire726  &  n_n177 ) | ( wire724  &  n_n177 ) | ( n_n177  &  wire717 ) ;
 assign wire121 = ( i_15_  &  n_n207  &  n_n170 ) | ( (~ i_15_)  &  n_n207  &  n_n170 ) | ( (~ i_15_)  &  n_n170  &  n_n209 ) ;
 assign wire148 = ( wire723  &  n_n170 ) | ( wire716  &  n_n170 ) | ( n_n170  &  wire730 ) ;
 assign wire161 = ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) ;
 assign wire415 = ( n_n216  &  wire730 ) | ( n_n216  &  wire718 ) ;
 assign wire162 = ( n_n216  &  wire716 ) | ( n_n216  &  wire730 ) | ( n_n216  &  wire718 ) ;
 assign wire438 = ( i_15_  &  n_n207  &  n_n149 ) | ( (~ i_15_)  &  n_n207  &  n_n149 ) ;
 assign wire163 = ( i_15_  &  n_n207  &  n_n149 ) | ( (~ i_15_)  &  n_n207  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n209 ) ;
 assign wire399 = ( n_n216  &  wire724 ) | ( n_n216  &  wire717 ) ;
 assign wire164 = ( wire726  &  n_n216 ) | ( n_n216  &  wire724 ) | ( n_n216  &  wire717 ) ;
 assign wire340 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) ;
 assign wire284 = ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) ;
 assign wire166 = ( wire723  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) ;
 assign wire339 = ( i_15_  &  n_n191  &  n_n207 ) | ( (~ i_15_)  &  n_n191  &  n_n207 ) ;
 assign wire169 = ( wire723  &  n_n216 ) | ( n_n216  &  wire727 ) ;
 assign wire174 = ( n_n177  &  wire721 ) | ( n_n177  &  wire725 ) | ( n_n177  &  wire728 ) ;
 assign wire177 = ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) ;
 assign wire179 = ( n_n177  &  wire716 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire718 ) ;
 assign wire183 = ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) ;
 assign wire184 = ( n_n184  &  wire716 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire718 ) ;
 assign wire187 = ( n_n191  &  wire722 ) | ( n_n191  &  wire727 ) | ( n_n191  &  wire715 ) ;
 assign wire425 = ( i_15_  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n207 ) ;
 assign wire192 = ( i_15_  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n207 ) | ( (~ i_15_)  &  n_n199  &  n_n209 ) ;
 assign wire193 = ( i_15_  &  n_n199  &  n_n204 ) | ( i_15_  &  n_n199  &  n_n211 ) | ( (~ i_15_)  &  n_n199  &  n_n211 ) ;
 assign wire424 = ( i_15_  &  n_n207  &  n_n156 ) | ( (~ i_15_)  &  n_n207  &  n_n156 ) ;
 assign wire194 = ( i_15_  &  n_n207  &  n_n156 ) | ( (~ i_15_)  &  n_n207  &  n_n156 ) | ( (~ i_15_)  &  n_n156  &  n_n209 ) ;
 assign wire195 = ( n_n184  &  wire716 ) | ( n_n184  &  wire722 ) | ( n_n184  &  wire727 ) ;
 assign wire358 = ( i_15_  &  n_n216  &  n_n211 ) | ( (~ i_15_)  &  n_n216  &  n_n211 ) ;
 assign wire196 = ( i_15_  &  n_n216  &  n_n204 ) | ( i_15_  &  n_n216  &  n_n211 ) | ( (~ i_15_)  &  n_n216  &  n_n211 ) ;
 assign wire198 = ( wire716  &  n_n156 ) | ( wire730  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire199 = ( wire716  &  n_n149 ) | ( wire722  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire362 = ( i_15_  &  n_n177  &  n_n211 ) | ( (~ i_15_)  &  n_n177  &  n_n211 ) ;
 assign wire200 = ( i_15_  &  n_n177  &  n_n204 ) | ( i_15_  &  n_n177  &  n_n211 ) | ( (~ i_15_)  &  n_n177  &  n_n211 ) ;
 assign wire366 = ( i_15_  &  n_n170  &  n_n211 ) | ( (~ i_15_)  &  n_n170  &  n_n211 ) ;
 assign wire201 = ( i_15_  &  n_n170  &  n_n204 ) | ( i_15_  &  n_n170  &  n_n211 ) | ( (~ i_15_)  &  n_n170  &  n_n211 ) ;
 assign wire202 = ( n_n184  &  wire724 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire730 ) ;
 assign wire203 = ( n_n199  &  wire729 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire718 ) ;
 assign wire204 = ( n_n149  &  wire719 ) | ( n_n149  &  wire728 ) ;
 assign wire205 = ( wire724  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire206 = ( n_n199  &  wire716 ) | ( n_n199  &  wire730 ) | ( n_n199  &  wire718 ) ;
 assign wire210 = ( wire723  &  n_n191 ) | ( n_n191  &  wire716 ) | ( n_n191  &  wire730 ) ;
 assign wire211 = ( n_n184  &  wire723 ) | ( n_n184  &  wire716 ) | ( n_n184  &  wire730 ) ;
 assign wire215 = ( n_n156  &  wire722 ) | ( n_n156  &  wire727 ) | ( n_n156  &  wire715 ) ;
 assign wire216 = ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire220 = ( wire724  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire221 = ( wire716  &  n_n149 ) | ( wire730  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire223 = ( i_15_  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n177  &  n_n209 ) ;
 assign wire229 = ( wire724  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire730 ) ;
 assign wire230 = ( wire723  &  n_n170 ) | ( wire716  &  n_n170 ) | ( n_n170  &  wire718 ) ;
 assign wire232 = ( i_15_  &  n_n204  &  n_n156 ) | ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) ;
 assign wire233 = ( n_n216  &  wire720 ) | ( n_n216  &  wire727 ) | ( n_n216  &  wire715 ) ;
 assign wire235 = ( i_15_  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n205  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n211 ) ;
 assign wire236 = ( wire723  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire237 = ( wire716  &  n_n170 ) | ( n_n170  &  wire722 ) | ( n_n170  &  wire727 ) ;
 assign wire238 = ( wire87 ) | ( wire729  &  n_n149 ) ;
 assign wire239 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) | ( n_n177  &  wire717 ) ;
 assign wire241 = ( n_n191  &  wire716 ) | ( n_n191  &  wire730 ) | ( n_n191  &  wire718 ) ;
 assign wire242 = ( n_n184  &  wire721 ) | ( n_n184  &  wire725 ) | ( n_n184  &  wire728 ) ;
 assign wire243 = ( n_n199  &  wire726 ) | ( n_n199  &  wire724 ) | ( n_n199  &  wire717 ) ;
 assign wire246 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n209 ) ;
 assign wire251 = ( i_15_  &  n_n216  &  n_n204 ) | ( i_15_  &  n_n216  &  n_n205 ) | ( (~ i_15_)  &  n_n216  &  n_n205 ) ;
 assign wire252 = ( n_n170  &  wire719 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire254 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire717 ) ;
 assign wire258 = ( n_n199  &  wire724 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire718 ) ;
 assign wire259 = ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) ;
 assign wire260 = ( wire723  &  n_n156 ) | ( wire716  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire261 = ( wire723  &  n_n216 ) | ( n_n216  &  wire716 ) | ( n_n216  &  wire718 ) ;
 assign wire262 = ( i_15_  &  n_n216  &  n_n205 ) | ( (~ i_15_)  &  n_n216  &  n_n205 ) | ( (~ i_15_)  &  n_n216  &  n_n211 ) ;
 assign wire264 = ( n_n199  &  wire723 ) | ( n_n199  &  wire716 ) | ( n_n199  &  wire718 ) ;
 assign wire265 = ( wire724  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire730 ) ;
 assign wire268 = ( n_n184  &  wire723 ) | ( n_n184  &  wire722 ) | ( n_n184  &  wire727 ) ;
 assign wire269 = ( n_n184  &  wire723 ) | ( n_n184  &  wire720 ) | ( n_n184  &  wire727 ) ;
 assign wire271 = ( i_15_  &  n_n184  &  n_n204 ) | ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) ;
 assign wire272 = ( n_n184  &  wire724 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire718 ) ;
 assign wire273 = ( wire723  &  n_n191 ) | ( n_n191  &  wire722 ) | ( n_n191  &  wire727 ) ;
 assign wire274 = ( i_15_  &  n_n170  &  n_n204 ) | ( i_15_  &  n_n170  &  n_n205 ) | ( (~ i_15_)  &  n_n170  &  n_n205 ) ;
 assign wire275 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) ;
 assign wire277 = ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) | ( n_n170  &  wire715 ) ;
 assign wire278 = ( i_15_  &  n_n191  &  n_n205 ) | ( (~ i_15_)  &  n_n191  &  n_n205 ) | ( (~ i_15_)  &  n_n191  &  n_n211 ) ;
 assign wire280 = ( i_15_  &  n_n207  &  n_n177 ) | ( (~ i_15_)  &  n_n207  &  n_n177 ) | ( (~ i_15_)  &  n_n177  &  n_n209 ) ;
 assign wire281 = ( wire716  &  n_n170 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire718 ) ;
 assign wire282 = ( i_15_  &  n_n170  &  n_n205 ) | ( (~ i_15_)  &  n_n170  &  n_n205 ) | ( (~ i_15_)  &  n_n170  &  n_n211 ) ;
 assign wire283 = ( wire723  &  n_n170 ) | ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) ;
 assign wire289 = ( wire723  &  n_n156 ) | ( n_n156  &  wire722 ) | ( n_n156  &  wire727 ) ;
 assign wire290 = ( wire716  &  n_n156 ) | ( n_n156  &  wire722 ) | ( n_n156  &  wire727 ) ;
 assign wire291 = ( n_n216  &  wire716 ) | ( n_n216  &  wire722 ) | ( n_n216  &  wire727 ) ;
 assign wire292 = ( wire729  &  n_n191 ) | ( n_n191  &  wire717 ) | ( n_n191  &  wire718 ) ;
 assign wire293 = ( wire729  &  n_n191 ) | ( n_n191  &  wire717 ) ;
 assign wire294 = ( wire723  &  n_n170 ) | ( n_n170  &  wire722 ) | ( n_n170  &  wire727 ) ;
 assign wire295 = ( n_n199  &  wire723 ) | ( n_n199  &  wire730 ) | ( n_n199  &  wire718 ) ;
 assign wire297 = ( n_n199  &  wire716 ) | ( n_n199  &  wire722 ) | ( n_n199  &  wire727 ) ;
 assign wire298 = ( wire723  &  n_n149 ) | ( wire722  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire299 = ( i_15_  &  n_n204  &  n_n149 ) | ( i_15_  &  n_n149  &  n_n211 ) | ( (~ i_15_)  &  n_n149  &  n_n211 ) ;
 assign wire300 = ( i_15_  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n149  &  n_n209 ) ;
 assign wire301 = ( i_15_  &  n_n191  &  n_n211 ) | ( (~ i_15_)  &  n_n191  &  n_n211 ) ;
 assign wire302 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire303 = ( wire729  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire304 = ( i_15_  &  n_n184  &  n_n204 ) | ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) ;
 assign wire305 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) ;
 assign wire306 = ( i_15_  &  n_n191  &  n_n204 ) | ( i_15_  &  n_n191  &  n_n211 ) | ( (~ i_15_)  &  n_n191  &  n_n211 ) ;
 assign wire307 = ( wire724  &  n_n191 ) | ( n_n191  &  wire717 ) | ( n_n191  &  wire730 ) ;
 assign wire309 = ( wire729  &  n_n216 ) | ( n_n216  &  wire717 ) | ( n_n216  &  wire718 ) ;
 assign wire310 = ( n_n184  &  wire723 ) | ( n_n184  &  wire716 ) | ( n_n184  &  wire718 ) ;
 assign wire311 = ( i_15_  &  n_n184  &  n_n213 ) | ( (~ i_15_)  &  n_n184  &  n_n213 ) | ( i_15_  &  n_n184  &  n_n207 ) ;
 assign wire312 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire718 ) ;
 assign wire314 = ( n_n184  &  wire723 ) | ( n_n184  &  wire730 ) | ( n_n184  &  wire718 ) ;
 assign wire316 = ( i_15_  &  n_n213  &  n_n149 ) | ( (~ i_15_)  &  n_n213  &  n_n149 ) | ( i_15_  &  n_n207  &  n_n149 ) ;
 assign wire317 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire718 ) ;
 assign wire318 = ( wire723  &  n_n191 ) | ( n_n191  &  wire716 ) | ( n_n191  &  wire718 ) ;
 assign wire319 = ( i_15_  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n213  &  n_n191 ) | ( i_15_  &  n_n191  &  n_n207 ) ;
 assign wire320 = ( n_n191  &  wire716 ) | ( n_n191  &  wire722 ) | ( n_n191  &  wire727 ) ;
 assign wire321 = ( i_15_  &  n_n213  &  n_n156 ) | ( (~ i_15_)  &  n_n213  &  n_n156 ) | ( i_15_  &  n_n207  &  n_n156 ) ;
 assign wire322 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n209 ) ;
 assign wire323 = ( i_15_  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n213  &  n_n199 ) | ( i_15_  &  n_n199  &  n_n207 ) ;
 assign wire324 = ( wire723  &  n_n177 ) | ( n_n177  &  wire722 ) | ( n_n177  &  wire727 ) ;
 assign wire325 = ( wire723  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) ;
 assign wire326 = ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) | ( i_15_  &  n_n207  &  n_n170 ) ;
 assign wire327 = ( wire729  &  n_n170 ) | ( n_n170  &  wire717 ) | ( n_n170  &  wire718 ) ;
 assign wire328 = ( i_15_  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n213  &  n_n199 ) | ( (~ i_15_)  &  n_n199  &  n_n209 ) ;
 assign wire329 = ( wire723  &  n_n170 ) | ( n_n170  &  wire730 ) | ( n_n170  &  wire718 ) ;
 assign wire330 = ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire717 ) ;
 assign wire331 = ( i_15_  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n213  &  n_n177 ) | ( i_15_  &  n_n207  &  n_n177 ) ;
 assign wire332 = ( i_15_  &  n_n199  &  n_n205 ) | ( (~ i_15_)  &  n_n199  &  n_n205 ) | ( (~ i_15_)  &  n_n199  &  n_n211 ) ;
 assign wire333 = ( wire723  &  n_n216 ) | ( n_n216  &  wire730 ) | ( n_n216  &  wire718 ) ;
 assign wire336 = ( wire723  &  n_n177 ) | ( n_n177  &  wire730 ) | ( n_n177  &  wire718 ) ;
 assign wire337 = ( wire723  &  n_n191 ) | ( n_n191  &  wire730 ) | ( n_n191  &  wire718 ) ;
 assign wire338 = ( n_n184  &  wire720 ) | ( n_n184  &  wire727 ) ;
 assign wire341 = ( wire723  &  n_n216 ) | ( n_n216  &  wire722 ) | ( n_n216  &  wire727 ) ;
 assign wire342 = ( wire723  &  n_n216 ) | ( n_n216  &  wire720 ) | ( n_n216  &  wire727 ) ;
 assign wire345 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire347 = ( wire723  &  n_n149 ) | ( wire716  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire349 = ( i_15_  &  n_n191  &  n_n204 ) | ( i_15_  &  n_n191  &  n_n205 ) | ( (~ i_15_)  &  n_n191  &  n_n205 ) ;
 assign wire351 = ( wire724  &  n_n149 ) | ( wire717  &  n_n149 ) | ( wire730  &  n_n149 ) ;
 assign wire352 = ( wire729  &  n_n170 ) | ( n_n170  &  wire717 ) ;
 assign wire354 = ( i_15_  &  n_n177  &  n_n205 ) | ( (~ i_15_)  &  n_n177  &  n_n205 ) | ( (~ i_15_)  &  n_n177  &  n_n211 ) ;
 assign wire357 = ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) | ( n_n191  &  wire715 ) ;
 assign wire368 = ( n_n199  &  wire723 ) | ( n_n199  &  wire722 ) | ( n_n199  &  wire727 ) ;
 assign wire369 = ( i_15_  &  n_n149  &  n_n211 ) | ( (~ i_15_)  &  n_n149  &  n_n211 ) ;
 assign wire370 = ( wire729  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign wire371 = ( i_15_  &  n_n156  &  n_n211 ) | ( (~ i_15_)  &  n_n156  &  n_n211 ) ;
 assign wire372 = ( wire729  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire730  &  n_n156 ) ;
 assign wire373 = ( wire729  &  n_n156 ) | ( wire717  &  n_n156 ) ;
 assign wire374 = ( n_n199  &  wire724 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire730 ) ;
 assign wire375 = ( wire729  &  n_n216 ) | ( n_n216  &  wire717 ) ;
 assign wire380 = ( wire723  &  n_n177 ) | ( n_n177  &  wire716 ) | ( n_n177  &  wire718 ) ;
 assign wire398 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire400 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) ;
 assign wire402 = ( wire724  &  n_n156 ) | ( n_n199  &  wire719 ) ;
 assign wire403 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire405 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire406 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire408 = ( wire726  &  n_n156 ) | ( n_n199  &  wire728 ) ;
 assign wire409 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire410 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire413 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire414 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire416 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire417 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire418 = ( i_9_  &  i_10_  &  i_11_  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire1840 = ( n_n198 ) | ( wire219 ) | ( wire108 ) | ( wire258 ) ;
 assign wire1844 = ( wire219 ) | ( wire108 ) | ( wire258 ) | ( wire16980 ) ;
 assign wire1853 = ( n_n198 ) | ( wire219 ) | ( wire108 ) | ( wire258 ) ;
 assign wire1862 = ( n_n216  &  wire719 ) | ( n_n199  &  wire725 ) ;
 assign wire1864 = ( wire168 ) | ( wire68 ) | ( wire151 ) | ( wire74 ) ;
 assign wire1902 = ( (~ i_9_)  &  i_10_  &  i_11_ ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign wire795 = ( wire117 ) | ( wire281 ) | ( wire294 ) ;
 assign wire805 = ( wire234 ) | ( wire84 ) | ( wire220 ) ;
 assign wire815 = ( n_n124  &  n_n159  &  n_n111 ) | ( n_n35  &  n_n159  &  n_n111 ) ;
 assign wire890 = ( wire158 ) | ( wire299 ) | ( n_n191  &  wire725 ) ;
 assign wire994 = ( wire302 ) | ( wire303 ) | ( wire316 ) ;
 assign wire1128 = ( wire723  &  n_n156 ) | ( wire723  &  n_n149 ) | ( wire718  &  n_n149 ) ;
 assign wire1131 = ( wire292 ) | ( wire311 ) | ( wire317 ) ;
 assign wire1203 = ( wire312 ) | ( wire326 ) | ( wire327 ) ;
 assign wire1209 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire1253 = ( n_n177  &  wire721 ) | ( n_n170  &  wire721 ) | ( n_n170  &  wire728 ) ;
 assign wire1328 = ( wire115 ) | ( wire221 ) | ( wire298 ) ;
 assign wire1356 = ( wire269 ) | ( wire275 ) | ( wire278 ) ;
 assign wire1409 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire1447 = ( wire244 ) | ( wire235 ) | ( wire236 ) ;
 assign wire1522 = ( wire130 ) | ( wire139 ) | ( wire128 ) ;
 assign wire1550 = ( n_n124  &  n_n159  &  n_n111 ) | ( n_n35  &  n_n159  &  n_n111 ) ;
 assign wire1557 = ( n_n170  &  wire721 ) | ( n_n177  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire1619 = ( wire282 ) | ( wire283 ) | ( wire325 ) ;
 assign wire1638 = ( wire235 ) | ( wire236 ) | ( n_n191  &  wire728 ) ;
 assign wire1643 = ( wire282 ) | ( wire283 ) | ( wire354 ) ;
 assign wire1661 = ( wire132 ) | ( wire46 ) | ( wire121 ) ;
 assign wire1768 = ( wire302 ) | ( wire316 ) | ( n_n191  &  wire721 ) ;
 assign wire1842 = ( wire219 ) | ( wire108 ) | ( wire258 ) ;
 assign wire138 = ( n_n2  &  wire270 ) | ( n_n2  &  wire372 ) ;
 assign wire439 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n48 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n48 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n48 ) ;
 assign wire441 = ( n_n65  &  n_n3 ) | ( n_n3  &  wire87 ) | ( n_n3  &  wire19935 ) ;
 assign wire467 = ( n_n5  &  wire145 ) | ( n_n5  &  n_n151 ) | ( n_n5  &  wire370 ) ;
 assign wire499 = ( n_n30  &  wire249 ) | ( n_n30  &  wire110 ) | ( n_n30  &  wire19905 ) ;
 assign wire501 = ( n_n162  &  n_n157  &  wire714  &  wire1592 ) ;
 assign wire507 = ( n_n31  &  wire337 ) | ( n_n31  &  wire338 ) | ( n_n31  &  wire19899 ) ;
 assign wire508 = ( n_n162  &  n_n220  &  n_n35  &  wire1590 ) ;
 assign wire510 = ( n_n30  &  wire284 ) | ( n_n30  &  wire337 ) ;
 assign wire513 = ( n_n31  &  wire314 ) | ( n_n31  &  n_n184  &  wire726 ) ;
 assign wire516 = ( n_n162  &  n_n157  &  wire714  &  wire1483 ) ;
 assign wire520 = ( n_n31  &  wire161 ) | ( n_n31  &  wire329 ) ;
 assign wire552 = ( n_n30  &  wire248 ) | ( n_n30  &  n_n64 ) | ( n_n30  &  wire408 ) ;
 assign wire556 = ( n_n36  &  wire19888 ) | ( n_n36  &  wire718  &  n_n149 ) ;
 assign wire1906 = ( n_n220  &  n_n35  &  n_n218  &  wire1779 ) ;
 assign wire1907 = ( n_n30  &  wire335 ) | ( n_n30  &  wire295 ) | ( n_n30  &  wire19882 ) ;
 assign wire1908 = ( n_n162  &  n_n157  &  wire714  &  wire1568 ) ;
 assign wire1910 = ( n_n33  &  wire278 ) | ( n_n33  &  wire19879 ) ;
 assign wire1912 = ( n_n184  &  wire728  &  n_n32 ) ;
 assign wire1914 = ( n_n32  &  wire269 ) | ( n_n32  &  wire275 ) ;
 assign wire1916 = ( n_n33  &  wire236 ) | ( n_n33  &  wire282 ) | ( n_n33  &  wire19874 ) ;
 assign wire1936 = ( n_n17  &  wire714  &  n_n218  &  wire1363 ) ;
 assign wire1937 = ( n_n197  &  wire283 ) | ( n_n197  &  wire325 ) | ( n_n197  &  wire19820 ) ;
 assign wire1938 = ( n_n200  &  n_n220  &  n_n218  &  wire1354 ) ;
 assign wire1939 = ( n_n212  &  wire325 ) | ( n_n212  &  wire354 ) | ( n_n212  &  wire1356 ) ;
 assign wire1940 = ( n_n123  &  wire259 ) | ( n_n123  &  wire329 ) | ( n_n123  &  wire19856 ) ;
 assign wire1945 = ( wire207  &  n_n125 ) | ( n_n125  &  wire416 ) | ( n_n125  &  wire19848 ) ;
 assign wire1946 = ( n_n123  &  wire408 ) | ( n_n123  &  wire19850 ) | ( n_n123  &  wire19853 ) ;
 assign wire1949 = ( n_n123  &  wire248 ) | ( n_n123  &  wire110 ) ;
 assign wire1950 = ( n_n125  &  wire249 ) | ( n_n125  &  wire726  &  n_n149 ) ;
 assign wire1951 = ( n_n108  &  wire335 ) | ( n_n108  &  wire333 ) ;
 assign wire1960 = ( n_n123  &  wire336 ) | ( n_n123  &  wire726  &  n_n177 ) ;
 assign wire1961 = ( n_n125  &  wire248 ) | ( n_n125  &  wire110 ) ;
 assign wire1962 = ( n_n125  &  n_n202 ) | ( n_n125  &  wire295 ) | ( n_n125  &  wire19835 ) ;
 assign wire1968 = ( n_n126  &  n_n220  &  n_n218  &  wire1513 ) ;
 assign wire1971 = ( n_n125  &  wire314 ) | ( n_n125  &  wire338 ) ;
 assign wire1972 = ( n_n125  &  wire335 ) | ( n_n125  &  wire333 ) ;
 assign wire1976 = ( n_n197  &  n_n60 ) | ( n_n197  &  wire235 ) | ( n_n197  &  wire19827 ) ;
 assign wire1979 = ( wire140  &  n_n197 ) | ( n_n197  &  wire244 ) ;
 assign wire1982 = ( n_n101  &  wire259 ) | ( n_n101  &  wire336 ) | ( n_n101  &  wire19770 ) ;
 assign wire1983 = ( n_n108  &  wire248 ) | ( n_n108  &  wire161 ) | ( n_n108  &  wire19774 ) ;
 assign wire1987 = ( n_n108  &  n_n202 ) | ( n_n108  &  wire295 ) | ( n_n108  &  wire19767 ) ;
 assign wire1988 = ( n_n162  &  n_n124  &  n_n220  &  wire1613 ) ;
 assign wire1990 = ( n_n101  &  wire338 ) | ( n_n101  &  wire726  &  n_n216 ) ;
 assign wire1991 = ( n_n108  &  wire337 ) | ( n_n108  &  wire19766 ) ;
 assign wire1992 = ( n_n108  &  wire259 ) | ( n_n108  &  wire336 ) | ( n_n108  &  wire19760 ) ;
 assign wire1993 = ( n_n101  &  wire284 ) | ( n_n101  &  wire329 ) | ( n_n101  &  wire19764 ) ;
 assign wire1995 = ( n_n101  &  wire314 ) | ( n_n101  &  n_n184  &  wire726 ) ;
 assign wire1996 = ( n_n108  &  wire314 ) | ( n_n108  &  wire338 ) ;
 assign wire1997 = ( n_n108  &  wire207 ) | ( n_n108  &  wire726  &  n_n156 ) ;
 assign wire1998 = ( n_n101  &  wire249 ) | ( n_n101  &  wire19759 ) ;
 assign wire1999 = ( n_n161  &  n_n48  &  n_n220  &  wire1641 ) ;
 assign wire2000 = ( wire140  &  n_n47 ) | ( n_n47  &  wire244 ) | ( n_n47  &  wire1643 ) ;
 assign wire2004 = ( n_n43  &  wire63 ) | ( n_n43  &  wire348 ) ;
 assign wire2017 = ( n_n46  &  wire1638 ) | ( n_n46  &  wire19798 ) ;
 assign wire2026 = ( n_n101  &  wire248 ) | ( n_n101  &  wire409 ) | ( n_n101  &  wire19780 ) ;
 assign wire2027 = ( n_n108  &  wire249 ) | ( n_n108  &  wire19782 ) | ( n_n108  &  wire19783 ) ;
 assign wire2032 = ( n_n101  &  wire408 ) | ( n_n101  &  wire19778 ) ;
 assign wire2035 = ( n_n40  &  wire166 ) | ( n_n40  &  wire278 ) | ( n_n40  &  wire1619 ) ;
 assign wire2040 = ( n_n42  &  wire63 ) | ( n_n42  &  wire348 ) ;
 assign wire2041 = ( n_n43  &  wire346 ) | ( n_n43  &  n_n191  &  wire728 ) ;
 assign wire2045 = ( n_n41  &  wire415 ) | ( n_n41  &  wire169 ) ;
 assign wire2051 = ( n_n41  &  wire275 ) | ( n_n41  &  wire278 ) | ( n_n41  &  wire19744 ) ;
 assign wire2062 = ( n_n36  &  wire156 ) | ( n_n36  &  wire19727 ) | ( n_n36  &  wire19728 ) ;
 assign wire2068 = ( n_n36  &  wire19724 ) | ( n_n36  &  wire726  &  n_n177 ) ;
 assign wire2070 = ( n_n34  &  wire128 ) | ( n_n34  &  wire348 ) ;
 assign wire2078 = ( n_n34  &  wire346 ) | ( n_n34  &  n_n191  &  wire720 ) ;
 assign wire2079 = ( n_n36  &  wire128 ) | ( n_n36  &  wire19716 ) ;
 assign wire2080 = ( n_n36  &  wire154 ) | ( n_n36  &  wire19714 ) ;
 assign wire2083 = ( n_n36  &  wire385 ) | ( n_n36  &  n_n191  &  wire720 ) ;
 assign wire2099 = ( n_n3  &  wire270 ) | ( n_n3  &  wire372 ) ;
 assign wire2108 = ( n_n162  &  n_n220  &  n_n35  &  wire1415 ) ;
 assign wire2119 = ( n_n125  &  n_n103 ) | ( n_n125  &  wire297 ) | ( n_n125  &  wire19672 ) ;
 assign wire2124 = ( n_n212  &  n_n138 ) | ( n_n212  &  wire163 ) | ( n_n212  &  wire405 ) ;
 assign wire2125 = ( n_n197  &  n_n138 ) | ( n_n197  &  wire407 ) | ( n_n197  &  wire163 ) ;
 assign wire2130 = ( n_n197  &  wire134 ) | ( n_n197  &  wire194 ) ;
 assign wire2134 = ( n_n124  &  n_n220  &  n_n218  &  wire1261 ) ;
 assign wire2136 = ( n_n123  &  wire54 ) | ( n_n123  &  n_n216  &  wire724 ) ;
 assign wire2139 = ( n_n125  &  wire111 ) | ( n_n125  &  wire291 ) ;
 assign wire2141 = ( n_n123  &  wire104 ) | ( n_n123  &  wire237 ) | ( n_n123  &  wire19654 ) ;
 assign wire2146 = ( n_n112  &  wire187 ) | ( n_n112  &  n_n191  &  wire720 ) ;
 assign wire2149 = ( n_n126  &  n_n220  &  n_n218  &  wire1089 ) ;
 assign wire2153 = ( n_n108  &  wire111 ) | ( n_n108  &  wire291 ) ;
 assign wire2155 = ( n_n123  &  wire279 ) | ( n_n123  &  wire724  &  n_n177 ) ;
 assign wire2156 = ( n_n125  &  wire59 ) | ( n_n125  &  wire290 ) ;
 assign wire2157 = ( n_n125  &  n_n72 ) | ( n_n125  &  wire118 ) | ( n_n125  &  wire401 ) ;
 assign wire2163 = ( n_n125  &  wire199 ) | ( n_n125  &  wire724  &  n_n149 ) ;
 assign wire2169 = ( n_n101  &  wire104 ) | ( n_n101  &  wire724  &  n_n170 ) ;
 assign wire2172 = ( n_n162  &  n_n126  &  n_n220  &  wire1741 ) ;
 assign wire2174 = ( n_n108  &  wire104 ) | ( n_n184  &  n_n108  &  wire724 ) ;
 assign wire2176 = ( n_n108  &  n_n103 ) | ( n_n108  &  wire297 ) | ( n_n108  &  wire19621 ) ;
 assign wire2177 = ( n_n162  &  n_n124  &  n_n220  &  wire1017 ) ;
 assign wire2179 = ( n_n101  &  wire54 ) | ( n_n101  &  n_n216  &  wire724 ) ;
 assign wire2180 = ( n_n108  &  wire320 ) | ( n_n108  &  wire19620 ) ;
 assign wire2181 = ( n_n47  &  wire47 ) | ( n_n47  &  wire192 ) | ( n_n47  &  wire322 ) ;
 assign wire2182 = ( n_n46  &  wire192 ) | ( n_n46  &  wire322 ) ;
 assign wire2190 = ( n_n101  &  wire290 ) | ( n_n101  &  wire406 ) | ( n_n101  &  wire19605 ) ;
 assign wire2191 = ( n_n108  &  wire199 ) | ( n_n108  &  wire19607 ) | ( n_n108  &  wire19608 ) ;
 assign wire2195 = ( n_n101  &  wire402 ) | ( n_n101  &  wire19602 ) ;
 assign wire2197 = ( n_n184  &  wire228  &  wire719 ) ;
 assign wire2204 = ( n_n47  &  wire134 ) | ( n_n47  &  wire1679 ) | ( n_n47  &  wire194 ) ;
 assign wire2205 = ( wire132  &  n_n46 ) | ( n_n46  &  wire121 ) | ( n_n46  &  wire280 ) ;
 assign wire2218 = ( n_n43  &  wire339 ) | ( n_n43  &  wire187 ) ;
 assign wire2229 = ( n_n40  &  wire48 ) | ( n_n40  &  wire167 ) | ( n_n40  &  wire1661 ) ;
 assign wire2232 = ( n_n40  &  wire151 ) | ( n_n40  &  wire192 ) ;
 assign wire2233 = ( n_n41  &  wire151 ) | ( n_n41  &  wire322 ) ;
 assign wire2239 = ( n_n42  &  wire339 ) | ( n_n42  &  wire187 ) ;
 assign wire2240 = ( n_n43  &  wire340 ) | ( n_n43  &  n_n191  &  wire719 ) ;
 assign wire2242 = ( n_n200  &  n_n48  &  n_n220  &  wire1628 ) ;
 assign wire2243 = ( n_n41  &  wire124 ) | ( n_n41  &  wire165 ) | ( n_n41  &  wire19565 ) ;
 assign wire2245 = ( wire207  &  n_n124  &  n_n48  &  n_n220 ) ;
 assign wire2257 = ( n_n17  &  n_n48  &  wire714  &  wire1630 ) ;
 assign wire2269 = ( n_n36  &  wire85 ) | ( n_n36  &  wire19535 ) ;
 assign wire2277 = ( n_n34  &  wire208 ) | ( n_n34  &  wire100 ) | ( n_n34  &  wire19530 ) ;
 assign wire2278 = ( n_n36  &  wire208 ) | ( n_n36  &  wire19530 ) | ( n_n36  &  wire19531 ) ;
 assign wire2281 = ( n_n34  &  wire19528 ) | ( n_n34  &  wire724  &  n_n177 ) ;
 assign wire2282 = ( n_n36  &  wire215 ) | ( n_n36  &  wire19529 ) ;
 assign wire2283 = ( n_n34  &  n_n190 ) | ( n_n34  &  wire107 ) | ( n_n34  &  wire340 ) ;
 assign wire2287 = ( n_n34  &  wire339 ) | ( n_n34  &  wire187 ) ;
 assign wire2290 = ( n_n34  &  wire219 ) | ( n_n34  &  wire425 ) ;
 assign wire2293 = ( n_n36  &  wire425 ) | ( n_n36  &  n_n191  &  wire720 ) ;
 assign wire2294 = ( n_n34  &  wire85 ) | ( n_n34  &  wire19519 ) ;
 assign wire2295 = ( n_n212  &  wire47 ) | ( n_n212  &  wire192 ) | ( n_n212  &  wire322 ) ;
 assign wire2296 = ( n_n197  &  wire151 ) | ( n_n197  &  wire192 ) | ( n_n197  &  wire322 ) ;
 assign wire2302 = ( n_n212  &  wire134 ) | ( n_n212  &  wire121 ) | ( n_n212  &  wire194 ) ;
 assign wire2303 = ( n_n197  &  wire55 ) | ( n_n197  &  wire121 ) | ( n_n197  &  wire280 ) ;
 assign wire2308 = ( n_n200  &  n_n220  &  n_n218  &  wire1347 ) ;
 assign wire2310 = ( n_n30  &  wire111 ) | ( n_n30  &  wire297 ) | ( n_n30  &  wire19500 ) ;
 assign wire2311 = ( n_n162  &  n_n157  &  wire714  &  wire1809 ) ;
 assign wire2323 = ( n_n36  &  wire84 ) | ( n_n36  &  wire438 ) | ( n_n36  &  wire19486 ) ;
 assign wire2324 = ( n_n34  &  wire84 ) | ( n_n34  &  wire424 ) | ( n_n34  &  wire19490 ) ;
 assign wire2329 = ( n_n162  &  n_n200  &  n_n220  &  wire167 ) ;
 assign wire2331 = ( n_n184  &  wire719  &  n_n32 ) ;
 assign wire2335 = ( n_n30  &  wire53 ) | ( n_n30  &  wire237 ) | ( n_n30  &  wire19472 ) ;
 assign wire2336 = ( n_n31  &  wire104 ) | ( n_n31  &  wire279 ) | ( n_n31  &  wire19476 ) ;
 assign wire2340 = ( n_n31  &  n_n90 ) | ( n_n31  &  wire195 ) | ( n_n31  &  wire19469 ) ;
 assign wire2341 = ( n_n162  &  n_n220  &  n_n35  &  wire1305 ) ;
 assign wire2343 = ( n_n30  &  wire291 ) | ( n_n30  &  n_n216  &  wire724 ) ;
 assign wire2344 = ( n_n31  &  wire98 ) | ( n_n31  &  wire320 ) ;
 assign wire2345 = ( n_n30  &  wire59 ) | ( n_n30  &  wire199 ) | ( n_n30  &  wire19464 ) ;
 assign wire2346 = ( n_n162  &  n_n157  &  wire714  &  wire1302 ) ;
 assign wire2349 = ( n_n30  &  n_n142 ) | ( n_n30  &  wire290 ) | ( n_n30  &  wire402 ) ;
 assign wire2350 = ( n_n31  &  wire59 ) | ( n_n31  &  wire724  &  n_n170 ) ;
 assign wire2351 = ( n_n30  &  wire279 ) | ( n_n30  &  wire19461 ) ;
 assign wire2352 = ( n_n30  &  wire19447 ) | ( n_n30  &  wire19448 ) ;
 assign wire2353 = ( n_n31  &  wire19449 ) | ( n_n31  &  wire19450 ) ;
 assign wire2356 = ( n_n31  &  wire19440 ) | ( n_n31  &  wire19441 ) ;
 assign wire2359 = ( n_n30  &  wire72 ) | ( n_n30  &  wire19438 ) ;
 assign wire2362 = ( n_n31  &  wire221 ) | ( n_n31  &  wire232 ) | ( n_n31  &  wire19436 ) ;
 assign wire2364 = ( n_n38  &  wire53 ) | ( n_n38  &  wire19426 ) ;
 assign wire2365 = ( n_n39  &  wire384 ) | ( n_n39  &  wire19427 ) ;
 assign wire2370 = ( n_n40  &  wire65 ) | ( n_n40  &  wire1557 ) ;
 assign wire2371 = ( n_n17  &  n_n48  &  wire714  &  wire1556 ) ;
 assign wire2372 = ( n_n40  &  wire82 ) | ( n_n40  &  wire19424 ) ;
 assign wire2373 = ( n_n17  &  n_n48  &  wire714  &  wire1404 ) ;
 assign wire2374 = ( n_n40  &  wire133 ) | ( n_n40  &  wire127 ) ;
 assign wire2375 = ( n_n41  &  wire227 ) | ( n_n41  &  wire221 ) | ( n_n41  &  wire19420 ) ;
 assign wire2379 = ( n_n41  &  wire19411 ) | ( n_n41  &  wire19412 ) ;
 assign wire2380 = ( n_n200  &  n_n48  &  n_n220  &  wire1211 ) ;
 assign wire2382 = ( n_n40  &  wire155 ) | ( n_n40  &  wire227 ) ;
 assign wire2384 = ( n_n34  &  wire223 ) | ( n_n34  &  wire274 ) ;
 assign wire2393 = ( n_n34  &  wire184 ) | ( n_n34  &  wire246 ) | ( n_n34  &  wire254 ) ;
 assign wire2398 = ( n_n36  &  wire179 ) | ( n_n36  &  wire223 ) | ( n_n36  &  wire239 ) ;
 assign wire2404 = ( n_n34  &  wire179 ) | ( n_n34  &  wire239 ) ;
 assign wire2405 = ( n_n157  &  wire714  &  n_n218  &  wire227 ) ;
 assign wire2407 = ( n_n30  &  wire274 ) | ( n_n30  &  wire277 ) | ( n_n30  &  wire19387 ) ;
 assign wire2410 = ( n_n31  &  wire155 ) | ( n_n31  &  wire227 ) | ( n_n31  &  wire69 ) ;
 assign wire2415 = ( n_n31  &  wire276 ) | ( n_n31  &  wire211 ) | ( n_n31  &  wire19375 ) ;
 assign wire2417 = ( n_n34  &  wire70 ) | ( n_n34  &  wire233 ) ;
 assign wire2418 = ( n_n36  &  wire206 ) | ( n_n36  &  wire328 ) | ( n_n36  &  wire330 ) ;
 assign wire2424 = ( n_n34  &  wire142 ) | ( n_n34  &  wire251 ) ;
 assign wire2427 = ( n_n38  &  n_n173 ) | ( n_n38  &  wire249 ) | ( n_n38  &  wire384 ) ;
 assign wire2428 = ( n_n126  &  n_n48  &  n_n220  &  wire1003 ) ;
 assign wire2435 = ( n_n36  &  wire142 ) | ( n_n36  &  wire233 ) | ( n_n36  &  wire251 ) ;
 assign wire2442 = ( n_n46  &  wire57 ) | ( n_n46  &  wire281 ) | ( n_n46  &  wire19339 ) ;
 assign wire2448 = ( n_n46  &  wire139 ) | ( n_n46  &  wire62 ) | ( n_n46  &  wire128 ) ;
 assign wire2449 = ( n_n47  &  wire349 ) | ( n_n47  &  wire357 ) | ( n_n47  &  wire19337 ) ;
 assign wire2451 = ( wire137  &  n_n47 ) | ( n_n47  &  wire146 ) | ( n_n47  &  wire254 ) ;
 assign wire2452 = ( n_n161  &  n_n48  &  n_n220  &  wire1507 ) ;
 assign wire2462 = ( n_n18  &  n_n48  &  wire714  &  wire81 ) ;
 assign wire2463 = ( n_n101  &  wire123 ) | ( n_n101  &  wire88 ) | ( n_n101  &  wire1409 ) ;
 assign wire2464 = ( n_n108  &  wire1409 ) | ( n_n108  &  wire19315 ) ;
 assign wire2468 = ( n_n108  &  wire72 ) | ( n_n108  &  wire19312 ) ;
 assign wire2475 = ( n_n18  &  n_n48  &  wire714  &  wire1341 ) ;
 assign wire2480 = ( n_n101  &  wire53 ) | ( n_n101  &  wire147 ) | ( n_n101  &  wire126 ) ;
 assign wire2481 = ( n_n108  &  wire79 ) | ( n_n108  &  wire19297 ) ;
 assign wire2487 = ( n_n101  &  wire241 ) | ( n_n101  &  wire19295 ) ;
 assign wire2488 = ( n_n162  &  n_n126  &  n_n220  &  wire384 ) ;
 assign wire2489 = ( n_n101  &  wire315 ) | ( n_n101  &  wire221 ) | ( n_n101  &  wire19289 ) ;
 assign wire2490 = ( n_n108  &  wire75 ) | ( n_n108  &  wire19290 ) | ( n_n108  &  wire19291 ) ;
 assign wire2493 = ( n_n101  &  wire384 ) | ( n_n101  &  wire79 ) | ( n_n101  &  wire19279 ) ;
 assign wire2498 = ( n_n125  &  wire251 ) | ( n_n125  &  wire328 ) ;
 assign wire2513 = ( n_n200  &  n_n220  &  n_n218  &  wire1292 ) ;
 assign wire2516 = ( n_n200  &  n_n220  &  n_n218  &  wire1290 ) ;
 assign wire2518 = ( n_n212  &  wire72 ) | ( n_n212  &  wire19246 ) ;
 assign wire2522 = ( n_n17  &  wire714  &  n_n218  &  wire1560 ) ;
 assign wire2523 = ( n_n197  &  wire92 ) | ( n_n197  &  wire19245 ) ;
 assign wire2524 = ( n_n17  &  wire714  &  n_n218  &  wire1558 ) ;
 assign wire2525 = ( n_n197  &  wire72 ) | ( n_n197  &  wire19243 ) ;
 assign wire2526 = ( n_n123  &  n_n183 ) | ( n_n123  &  wire233 ) | ( n_n123  &  wire251 ) ;
 assign wire2532 = ( n_n197  &  wire68 ) | ( n_n197  &  wire81 ) | ( n_n197  &  wire74 ) ;
 assign wire2537 = ( n_n212  &  n_n198 ) | ( n_n212  &  wire206 ) | ( n_n212  &  wire328 ) ;
 assign wire2540 = ( n_n197  &  wire63 ) | ( n_n197  &  wire184 ) | ( n_n197  &  wire19226 ) ;
 assign wire2543 = ( n_n197  &  wire233 ) | ( n_n197  &  wire246 ) | ( n_n197  &  wire19219 ) ;
 assign wire2545 = ( n_n125  &  wire142 ) | ( n_n125  &  wire233 ) ;
 assign wire2548 = ( n_n71  &  n_n123 ) | ( n_n123  &  wire49 ) | ( n_n123  &  wire92 ) ;
 assign wire2549 = ( n_n126  &  n_n220  &  wire928  &  n_n218 ) ;
 assign wire2556 = ( n_n124  &  n_n220  &  n_n218  &  wire1562 ) ;
 assign wire2557 = ( n_n125  &  wire88 ) | ( n_n125  &  wire19204 ) ;
 assign wire2558 = ( n_n124  &  n_n220  &  n_n218  &  wire1251 ) ;
 assign wire2559 = ( n_n125  &  wire83 ) | ( n_n125  &  wire1253 ) ;
 assign wire2560 = ( n_n101  &  wire143 ) | ( n_n101  &  wire111 ) | ( n_n101  &  wire154 ) ;
 assign wire2565 = ( n_n108  &  wire241 ) | ( n_n108  &  wire19194 ) ;
 assign wire2567 = ( n_n220  &  wire1072  &  n_n111  &  wire16987 ) ;
 assign wire2568 = ( n_n101  &  wire206 ) | ( n_n101  &  wire328 ) | ( n_n101  &  wire330 ) ;
 assign wire2576 = ( n_n101  &  wire276 ) | ( n_n101  &  wire211 ) | ( n_n101  &  wire19185 ) ;
 assign wire2578 = ( n_n123  &  wire148 ) | ( n_n123  &  wire274 ) | ( n_n123  &  wire277 ) ;
 assign wire2579 = ( n_n125  &  wire179 ) | ( n_n125  &  wire223 ) | ( n_n125  &  wire19174 ) ;
 assign wire2584 = ( n_n125  &  wire276 ) | ( n_n125  &  wire211 ) | ( n_n125  &  wire271 ) ;
 assign wire2585 = ( n_n123  &  wire184 ) | ( n_n123  &  wire246 ) | ( n_n123  &  wire19168 ) ;
 assign wire2588 = ( n_n125  &  wire227 ) | ( n_n125  &  wire232 ) ;
 assign wire2594 = ( n_n125  &  wire315 ) | ( n_n125  &  wire221 ) | ( n_n125  &  wire300 ) ;
 assign wire2595 = ( wire844  &  n_n124  &  n_n220  &  n_n218 ) ;
 assign wire2598 = ( wire52  &  n_n112 ) | ( wire98  &  n_n112 ) | ( n_n112  &  wire51 ) ;
 assign wire2599 = ( n_n113  &  wire211 ) | ( n_n113  &  wire271 ) | ( n_n113  &  wire19150 ) ;
 assign wire2606 = ( n_n31  &  wire206 ) | ( n_n31  &  wire328 ) | ( n_n31  &  wire19144 ) ;
 assign wire2610 = ( n_n33  &  wire210 ) | ( n_n33  &  wire349 ) | ( n_n33  &  wire357 ) ;
 assign wire2614 = ( n_n30  &  wire68 ) | ( n_n30  &  wire74 ) ;
 assign wire2615 = ( n_n31  &  wire142 ) | ( n_n31  &  wire233 ) | ( n_n31  &  wire251 ) ;
 assign wire2618 = ( n_n33  &  wire19128 ) | ( n_n33  &  wire19129 ) ;
 assign wire2630 = ( n_n18  &  n_n48  &  wire714  &  wire1582 ) ;
 assign wire2631 = ( n_n46  &  wire49 ) | ( n_n46  &  wire19113 ) | ( n_n46  &  wire19116 ) ;
 assign wire2634 = ( n_n18  &  n_n48  &  wire714  &  wire1553 ) ;
 assign wire2635 = ( n_n46  &  wire90 ) | ( n_n46  &  n_n62 ) | ( n_n46  &  wire19110 ) ;
 assign wire2636 = ( n_n43  &  wire210 ) | ( n_n43  &  wire357 ) ;
 assign wire2638 = ( n_n18  &  n_n48  &  wire714  &  wire1503 ) ;
 assign wire2643 = ( n_n161  &  n_n48  &  n_n220  &  wire1500 ) ;
 assign wire2645 = ( n_n41  &  wire206 ) | ( n_n41  &  wire328 ) | ( n_n41  &  wire330 ) ;
 assign wire2646 = ( n_n40  &  wire68 ) | ( n_n40  &  wire74 ) | ( n_n40  &  wire19094 ) ;
 assign wire2657 = ( n_n17  &  n_n48  &  wire714  &  wire1295 ) ;
 assign wire2666 = ( n_n42  &  wire210 ) | ( n_n42  &  wire349 ) ;
 assign wire2669 = ( n_n41  &  wire147 ) | ( n_n41  &  wire126 ) ;
 assign wire2676 = ( n_n17  &  n_n48  &  wire714  &  wire1154 ) ;
 assign wire2679 = ( wire52  &  n_n40 ) | ( n_n40  &  wire63 ) | ( n_n40  &  wire277 ) ;
 assign wire2686 = ( n_n33  &  wire148 ) | ( n_n33  &  wire274 ) | ( n_n33  &  wire19053 ) ;
 assign wire2691 = ( n_n36  &  wire83 ) | ( n_n36  &  wire1209 ) ;
 assign wire2692 = ( n_n34  &  wire118 ) | ( n_n34  &  wire60 ) ;
 assign wire2693 = ( n_n36  &  wire221 ) | ( n_n36  &  wire232 ) | ( n_n36  &  wire19047 ) ;
 assign wire2700 = ( n_n34  &  wire227 ) | ( n_n34  &  wire232 ) | ( n_n34  &  wire19043 ) ;
 assign wire2702 = ( n_n220  &  n_n35  &  n_n218  &  wire1143 ) ;
 assign wire2703 = ( n_n36  &  wire88 ) | ( n_n36  &  wire19038 ) ;
 assign wire2704 = ( n_n30  &  wire197 ) | ( n_n30  &  wire203 ) | ( n_n30  &  wire323 ) ;
 assign wire2705 = ( n_n31  &  wire203 ) | ( n_n31  &  wire309 ) | ( n_n31  &  wire323 ) ;
 assign wire2712 = ( n_n41  &  wire230 ) | ( n_n41  &  wire352 ) | ( n_n41  &  wire19016 ) ;
 assign wire2713 = ( n_n40  &  wire230 ) | ( n_n40  &  wire400 ) | ( n_n40  &  wire19020 ) ;
 assign wire2717 = ( n_n40  &  n_n107 ) | ( n_n40  &  wire264 ) | ( n_n40  &  wire19013 ) ;
 assign wire2718 = ( n_n17  &  n_n48  &  wire714  &  wire1735 ) ;
 assign wire2720 = ( n_n184  &  wire721  &  wire1277 ) | ( n_n191  &  wire721  &  wire1277 ) ;
 assign wire2721 = ( n_n162  &  n_n161  &  wire52  &  n_n220 ) ;
 assign wire2724 = ( wire1704  &  wire318 ) | ( n_n191  &  wire715  &  wire1704 ) ;
 assign wire2726 = ( n_n41  &  wire305 ) | ( n_n41  &  wire310 ) ;
 assign wire2728 = ( n_n41  &  wire293 ) | ( n_n184  &  n_n41  &  wire715 ) ;
 assign wire2729 = ( n_n40  &  wire310 ) | ( n_n40  &  wire19008 ) ;
 assign wire2730 = ( n_n40  &  wire293 ) | ( n_n40  &  n_n170  &  wire715 ) ;
 assign wire2731 = ( n_n41  &  wire380 ) | ( n_n41  &  wire19006 ) ;
 assign wire2733 = ( n_n101  &  n_n107 ) | ( n_n101  &  wire264 ) | ( n_n101  &  wire19001 ) ;
 assign wire2738 = ( n_n101  &  wire261 ) | ( n_n101  &  wire375 ) ;
 assign wire2739 = ( n_n108  &  wire318 ) | ( n_n108  &  n_n191  &  wire715 ) ;
 assign wire2740 = ( n_n101  &  wire293 ) | ( n_n101  &  wire318 ) | ( n_n101  &  wire18993 ) ;
 assign wire2741 = ( n_n108  &  wire310 ) | ( n_n108  &  wire400 ) | ( n_n108  &  wire18997 ) ;
 assign wire2743 = ( n_n108  &  wire293 ) | ( n_n184  &  n_n108  &  wire715 ) ;
 assign wire2744 = ( n_n101  &  wire310 ) | ( n_n101  &  wire18992 ) ;
 assign wire2746 = ( n_n162  &  n_n126  &  n_n220  &  wire1498 ) ;
 assign wire2748 = ( n_n108  &  wire352 ) | ( n_n108  &  n_n156  &  wire715 ) ;
 assign wire2750 = ( n_n161  &  n_n48  &  n_n220  &  wire1201 ) ;
 assign wire2751 = ( n_n47  &  wire303 ) | ( n_n47  &  wire321 ) | ( n_n47  &  wire1203 ) ;
 assign wire2775 = ( n_n108  &  wire345 ) | ( n_n108  &  wire347 ) | ( n_n108  &  wire18956 ) ;
 assign wire2776 = ( n_n101  &  wire260 ) | ( n_n101  &  wire18958 ) | ( n_n101  &  wire18959 ) ;
 assign wire2784 = ( n_n123  &  wire147 ) | ( n_n123  &  wire18944 ) ;
 assign wire2785 = ( n_n125  &  wire146 ) | ( n_n125  &  wire183 ) | ( n_n125  &  wire18945 ) ;
 assign wire2791 = ( wire1244  &  wire1243 ) ;
 assign wire2797 = ( n_n220  &  n_n111  &  wire412  &  wire16987 ) ;
 assign wire2801 = ( n_n113  &  wire305 ) | ( n_n113  &  wire310 ) ;
 assign wire2802 = ( n_n112  &  wire318 ) | ( n_n112  &  n_n191  &  wire715 ) ;
 assign wire2808 = ( n_n123  &  wire123 ) | ( n_n123  &  wire175 ) ;
 assign wire2809 = ( n_n125  &  wire133 ) | ( n_n125  &  wire729  &  n_n149 ) ;
 assign wire2814 = ( n_n123  &  wire146 ) | ( n_n123  &  wire729  &  n_n177 ) ;
 assign wire2815 = ( n_n125  &  wire123 ) | ( n_n125  &  wire175 ) ;
 assign wire2817 = ( n_n123  &  wire143 ) | ( n_n123  &  wire364 ) ;
 assign wire2825 = ( n_n125  &  wire143 ) | ( n_n125  &  wire364 ) ;
 assign wire2828 = ( n_n197  &  n_n137 ) | ( n_n197  &  wire302 ) | ( n_n197  &  wire18921 ) ;
 assign wire2831 = ( n_n197  &  wire303 ) | ( n_n197  &  wire321 ) ;
 assign wire2842 = ( n_n123  &  wire139 ) | ( n_n184  &  n_n123  &  wire729 ) ;
 assign wire2843 = ( n_n125  &  wire139 ) | ( n_n125  &  wire313 ) ;
 assign wire2848 = ( n_n17  &  wire714  &  n_n218  &  wire1132 ) ;
 assign wire2849 = ( n_n197  &  wire326 ) | ( n_n197  &  wire327 ) | ( n_n197  &  wire18908 ) ;
 assign wire2850 = ( n_n200  &  n_n220  &  n_n218  &  wire1129 ) ;
 assign wire2851 = ( n_n212  &  wire312 ) | ( n_n212  &  wire331 ) | ( n_n212  &  wire1131 ) ;
 assign wire2853 = ( n_n36  &  wire183 ) | ( n_n36  &  wire18894 ) ;
 assign wire2861 = ( n_n34  &  wire376 ) | ( n_n34  &  wire729  &  n_n177 ) ;
 assign wire2865 = ( n_n34  &  wire139 ) | ( n_n34  &  wire313 ) | ( n_n34  &  n_n89 ) ;
 assign wire2866 = ( n_n36  &  n_n89 ) | ( n_n36  &  wire146 ) | ( n_n36  &  wire383 ) ;
 assign wire2870 = ( n_n34  &  wire257 ) | ( n_n34  &  n_n184  &  wire729 ) ;
 assign wire2875 = ( n_n34  &  n_n139 ) | ( n_n34  &  wire175 ) | ( n_n34  &  wire18879 ) ;
 assign wire2896 = ( n_n40  &  wire838 ) | ( n_n40  &  n_n70 ) | ( n_n40  &  wire347 ) ;
 assign wire2897 = ( n_n41  &  n_n141 ) | ( n_n41  &  wire260 ) | ( n_n41  &  wire373 ) ;
 assign wire2900 = ( n_n40  &  wire345 ) | ( n_n40  &  n_n156  &  wire715 ) ;
 assign wire2901 = ( n_n41  &  wire347 ) | ( n_n41  &  wire18859 ) ;
 assign wire2909 = ( n_n126  &  n_n48  &  n_n220  &  wire1126 ) ;
 assign wire2910 = ( n_n38  &  wire1128 ) | ( n_n38  &  wire18852 ) ;
 assign wire2911 = ( n_n17  &  n_n48  &  wire714  &  wire988 ) ;
 assign wire2914 = ( n_n33  &  wire293 ) | ( n_n33  &  wire18847 ) ;
 assign wire2915 = ( n_n162  &  n_n157  &  wire714  &  wire197 ) ;
 assign wire2923 = ( n_n65  &  n_n2 ) | ( n_n2  &  wire87 ) | ( n_n2  &  wire18835 ) ;
 assign wire2937 = ( wire213  &  n_n199  &  wire721 ) ;
 assign wire2939 = ( n_n32  &  wire305 ) | ( n_n32  &  wire310 ) ;
 assign wire2940 = ( n_n33  &  wire230 ) | ( n_n33  &  wire318 ) | ( n_n33  &  wire18824 ) ;
 assign wire2943 = ( n_n33  &  wire347 ) | ( n_n33  &  wire352 ) | ( n_n33  &  wire18821 ) ;
 assign wire2944 = ( n_n184  &  wire715  &  n_n32 ) ;
 assign wire2952 = ( n_n3  &  wire95 ) | ( wire95  &  wire18810 ) ;
 assign wire2953 = ( wire729  &  n_n156  &  n_n12 ) | ( wire729  &  n_n156  &  wire18811 ) ;
 assign wire2958 = ( n_n9  &  wire95 ) | ( n_n6  &  wire95 ) | ( wire95  &  n_n12 ) ;
 assign wire2959 = ( n_n71  &  n_n9 ) | ( n_n71  &  n_n6 ) | ( n_n71  &  n_n5 ) ;
 assign wire2962 = ( n_n162  &  n_n184  &  n_n163  &  n_n161 ) ;
 assign wire2964 = ( n_n31  &  wire118 ) | ( n_n31  &  wire221 ) | ( n_n31  &  wire298 ) ;
 assign wire2965 = ( n_n162  &  n_n220  &  n_n35  &  wire1096 ) ;
 assign wire2970 = ( n_n30  &  wire152 ) | ( n_n30  &  wire18784 ) ;
 assign wire2974 = ( n_n30  &  wire59 ) | ( n_n30  &  wire289 ) ;
 assign wire2975 = ( n_n31  &  wire115 ) | ( n_n31  &  wire729  &  n_n149 ) ;
 assign wire2977 = ( n_n162  &  n_n220  &  n_n35  &  wire1023 ) ;
 assign wire2979 = ( n_n30  &  wire172 ) | ( n_n30  &  wire209 ) ;
 assign wire2981 = ( n_n31  &  wire218 ) | ( n_n31  &  wire212 ) | ( n_n31  &  wire18771 ) ;
 assign wire2985 = ( n_n33  &  wire147 ) | ( n_n33  &  wire158 ) ;
 assign wire2995 = ( n_n33  &  wire52 ) | ( n_n33  &  wire63 ) | ( n_n33  &  wire222 ) ;
 assign wire3001 = ( n_n30  &  n_n95 ) | ( n_n30  &  wire111 ) | ( n_n30  &  wire341 ) ;
 assign wire3006 = ( n_n30  &  wire206 ) | ( n_n30  &  wire243 ) | ( n_n30  &  wire368 ) ;
 assign wire3008 = ( n_n33  &  n_n191  &  wire725 ) ;
 assign wire3013 = ( n_n162  &  n_n220  &  n_n35  &  wire860 ) ;
 assign wire3014 = ( n_n31  &  wire268 ) | ( n_n31  &  wire273 ) | ( n_n31  &  wire18744 ) ;
 assign wire3015 = ( n_n30  &  wire162 ) | ( n_n30  &  wire164 ) ;
 assign wire3020 = ( n_n31  &  n_n83 ) | ( n_n31  &  wire120 ) | ( n_n31  &  wire795 ) ;
 assign wire3027 = ( n_n31  &  wire179 ) | ( n_n31  &  wire184 ) | ( n_n31  &  wire18731 ) ;
 assign wire3032 = ( n_n31  &  wire116 ) | ( n_n31  &  wire198 ) | ( n_n31  &  wire18725 ) ;
 assign wire3044 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) ;
 assign wire3059 = ( n_n162  &  n_n16  &  n_n19 ) | ( n_n16  &  n_n19  &  n_n48 ) ;
 assign wire3060 = ( n_n18  &  n_n19  &  n_n218 ) | ( n_n18  &  n_n19  &  n_n111 ) ;
 assign wire3066 = ( wire344  &  wire815 ) | ( wire344  &  wire18696 ) ;
 assign wire3067 = ( n_n6  &  n_n68 ) | ( n_n68  &  wire398 ) | ( n_n68  &  wire815 ) ;
 assign wire3068 = ( n_n162  &  wire381  &  n_n124  &  n_n220 ) ;
 assign wire3069 = ( n_n162  &  wire172  &  n_n161  &  n_n220 ) ;
 assign wire3078 = ( n_n101  &  wire80 ) | ( n_n101  &  wire78 ) ;
 assign wire3079 = ( wire381  &  n_n108 ) | ( n_n108  &  wire18687 ) ;
 assign wire3080 = ( n_n108  &  wire173 ) | ( n_n108  &  wire204 ) ;
 assign wire3081 = ( n_n101  &  wire245 ) | ( n_n101  &  wire18686 ) ;
 assign wire3093 = ( n_n108  &  wire107 ) | ( n_n108  &  wire211 ) | ( n_n108  &  wire18676 ) ;
 assign wire3098 = ( n_n108  &  wire240 ) | ( n_n108  &  wire187 ) | ( n_n108  &  wire18662 ) ;
 assign wire3102 = ( n_n101  &  wire234 ) | ( n_n101  &  wire220 ) ;
 assign wire3111 = ( n_n108  &  wire222 ) | ( n_n108  &  wire242 ) | ( n_n108  &  wire18649 ) ;
 assign wire3113 = ( n_n101  &  wire155 ) | ( n_n101  &  wire205 ) | ( n_n101  &  wire215 ) ;
 assign wire3118 = ( n_n108  &  wire225 ) | ( n_n108  &  wire205 ) | ( n_n108  &  wire18635 ) ;
 assign wire3123 = ( n_n42  &  wire256 ) | ( n_n42  &  wire216 ) ;
 assign wire3124 = ( wire130  &  n_n43 ) | ( n_n43  &  n_n116 ) | ( n_n43  &  wire242 ) ;
 assign wire3128 = ( n_n42  &  wire130 ) | ( n_n42  &  wire124 ) ;
 assign wire3135 = ( n_n212  &  wire152 ) | ( n_n212  &  n_n149  &  wire719 ) ;
 assign wire3136 = ( wire157  &  n_n197 ) | ( n_n197  &  wire204 ) | ( n_n197  &  wire18617 ) ;
 assign wire3142 = ( n_n197  &  wire171 ) | ( n_n197  &  wire252 ) | ( n_n197  &  wire18609 ) ;
 assign wire3143 = ( n_n17  &  wire714  &  n_n218  &  wire1655 ) ;
 assign wire3154 = ( n_n197  &  wire242 ) | ( n_n197  &  n_n184  &  wire719 ) ;
 assign wire3155 = ( n_n212  &  wire247 ) | ( n_n212  &  wire160 ) | ( n_n212  &  wire171 ) ;
 assign wire3177 = ( n_n212  &  wire147 ) | ( n_n212  &  wire126 ) ;
 assign wire3194 = ( i_5_  &  n_n18  &  n_n159  &  wire17176 ) ;
 assign wire3195 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n159  &  n_n111 ) ;
 assign wire3201 = ( wire168  &  n_n123 ) | ( n_n123  &  wire68 ) | ( n_n123  &  wire151 ) ;
 assign wire3202 = ( n_n125  &  wire181 ) | ( n_n125  &  wire154 ) | ( n_n125  &  wire18559 ) ;
 assign wire3209 = ( n_n124  &  n_n220  &  n_n218  &  wire1695 ) ;
 assign wire3210 = ( n_n125  &  wire63 ) | ( n_n125  &  wire48 ) | ( n_n125  &  wire18553 ) ;
 assign wire3217 = ( n_n123  &  wire125 ) | ( n_n123  &  wire242 ) | ( n_n123  &  wire18540 ) ;
 assign wire3219 = ( n_n123  &  wire174 ) | ( n_n123  &  wire252 ) | ( n_n123  &  wire18529 ) ;
 assign wire3220 = ( n_n126  &  n_n220  &  n_n218  &  wire1336 ) ;
 assign wire3222 = ( n_n123  &  wire160 ) | ( n_n123  &  wire171 ) ;
 assign wire3223 = ( n_n125  &  wire217 ) | ( n_n125  &  wire18528 ) ;
 assign wire3224 = ( n_n123  &  wire147 ) | ( n_n123  &  wire958 ) | ( n_n123  &  wire46 ) ;
 assign wire3225 = ( wire132  &  n_n125 ) | ( n_n125  &  wire149 ) | ( n_n125  &  wire126 ) ;
 assign wire3229 = ( n_n123  &  wire129 ) | ( n_n123  &  wire63 ) | ( n_n123  &  wire48 ) ;
 assign wire3230 = ( n_n125  &  wire146 ) | ( n_n125  &  wire46 ) | ( n_n125  &  wire18521 ) ;
 assign wire3232 = ( n_n126  &  n_n220  &  n_n218  &  wire1465 ) ;
 assign wire3233 = ( n_n123  &  wire146 ) | ( n_n123  &  wire127 ) | ( n_n123  &  wire18517 ) ;
 assign wire3234 = ( n_n65  &  n_n2 ) | ( n_n2  &  n_n89 ) | ( n_n2  &  wire87 ) ;
 assign wire3244 = ( wire145  &  n_n3 ) | ( n_n3  &  n_n186 ) | ( n_n3  &  wire170 ) ;
 assign wire3245 = ( n_n4  &  wire185 ) | ( n_n4  &  wire270 ) ;
 assign wire3248 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) ;
 assign wire3256 = ( n_n65  &  n_n9 ) | ( n_n9  &  n_n89 ) | ( n_n9  &  wire87 ) ;
 assign wire3257 = ( n_n65  &  n_n10 ) | ( wire77  &  n_n10 ) | ( n_n10  &  wire87 ) ;
 assign wire3258 = ( n_n41  &  wire1386 ) | ( n_n41  &  n_n216  &  wire724 ) ;
 assign wire3264 = ( n_n40  &  wire154 ) | ( n_n40  &  wire124 ) | ( n_n40  &  wire18481 ) ;
 assign wire3271 = ( n_n41  &  wire143 ) | ( n_n41  &  wire154 ) ;
 assign wire3275 = ( n_n41  &  wire134 ) | ( n_n41  &  wire123 ) | ( n_n41  &  wire18467 ) ;
 assign wire3279 = ( n_n40  &  wire198 ) | ( n_n40  &  wire289 ) ;
 assign wire3280 = ( n_n41  &  wire133 ) | ( n_n41  &  wire127 ) | ( n_n41  &  wire18457 ) ;
 assign wire3291 = ( n_n17  &  n_n48  &  wire714  &  wire1381 ) ;
 assign wire3292 = ( n_n40  &  wire146 ) | ( n_n40  &  wire46 ) | ( n_n40  &  wire18450 ) ;
 assign wire3296 = ( wire129  &  n_n40 ) | ( n_n40  &  wire147 ) | ( n_n40  &  wire18444 ) ;
 assign wire3298 = ( n_n17  &  n_n48  &  wire714  &  wire1520 ) ;
 assign wire3299 = ( n_n40  &  wire63 ) | ( n_n40  &  wire48 ) | ( n_n40  &  wire1522 ) ;
 assign wire3300 = ( n_n46  &  wire53 ) | ( n_n46  &  wire294 ) ;
 assign wire3301 = ( n_n47  &  wire120 ) | ( n_n47  &  wire281 ) | ( n_n47  &  wire18432 ) ;
 assign wire3308 = ( n_n18  &  n_n48  &  wire714  &  wire1576 ) ;
 assign wire3312 = ( n_n46  &  wire111 ) | ( n_n46  &  wire341 ) ;
 assign wire3313 = ( n_n47  &  wire206 ) | ( n_n47  &  wire243 ) | ( n_n47  &  wire18416 ) ;
 assign wire3325 = ( n_n46  &  n_n102 ) | ( n_n46  &  wire162 ) | ( n_n46  &  wire164 ) ;
 assign wire3328 = ( n_n47  &  wire241 ) | ( n_n47  &  wire268 ) | ( n_n47  &  wire18408 ) ;
 assign wire3333 = ( n_n46  &  wire59 ) | ( n_n46  &  wire289 ) | ( n_n46  &  wire1328 ) ;
 assign wire3337 = ( n_n47  &  wire256 ) | ( n_n47  &  wire216 ) ;
 assign wire3338 = ( wire172  &  n_n46 ) | ( n_n46  &  wire217 ) | ( n_n46  &  wire18394 ) ;
 assign wire3342 = ( n_n47  &  wire218 ) | ( n_n47  &  wire212 ) | ( n_n47  &  wire18386 ) ;
 assign wire3343 = ( n_n46  &  wire247 ) | ( n_n46  &  wire116 ) | ( n_n46  &  wire18391 ) ;
 assign wire3349 = ( n_n47  &  wire179 ) | ( n_n47  &  wire184 ) | ( n_n47  &  wire18384 ) ;
 assign wire3353 = ( n_n46  &  n_n77 ) | ( n_n46  &  wire117 ) | ( n_n46  &  wire281 ) ;
 assign wire3374 = ( wire185  &  wire1427 ) | ( wire1427  &  wire270 ) | ( wire1427  &  wire372 ) ;
 assign wire3375 = ( n_n3  &  wire270 ) | ( n_n3  &  wire372 ) ;
 assign wire3376 = ( n_n161  &  wire185  &  n_n48  &  n_n159 ) ;
 assign wire3385 = ( n_n138  &  n_n43 ) | ( n_n43  &  wire62 ) | ( n_n43  &  wire272 ) ;
 assign wire3392 = ( n_n43  &  wire107 ) | ( n_n43  &  wire211 ) ;
 assign wire3396 = ( n_n42  &  wire217 ) | ( n_n42  &  n_n184  &  wire725 ) ;
 assign wire3397 = ( wire172  &  n_n43 ) | ( n_n43  &  wire216 ) ;
 assign wire3403 = ( n_n112  &  wire222 ) | ( n_n112  &  n_n191  &  wire725 ) ;
 assign wire3404 = ( n_n42  &  wire107 ) | ( n_n42  &  wire211 ) | ( n_n42  &  wire272 ) ;
 assign wire3409 = ( wire52  &  n_n112 ) | ( wire129  &  n_n112 ) | ( n_n112  &  wire48 ) ;
 assign wire3410 = ( n_n113  &  wire124 ) | ( n_n113  &  wire128 ) | ( n_n113  &  wire18337 ) ;
 assign wire3415 = ( n_n5  &  wire145 ) | ( n_n5  &  n_n151 ) | ( n_n5  &  wire370 ) ;
 assign wire3425 = ( n_n4  &  wire185 ) | ( n_n4  &  wire87 ) ;
 assign wire3433 = ( n_n5  &  n_n144 ) | ( n_n5  &  n_n186 ) | ( n_n5  &  wire170 ) ;
 assign wire3434 = ( n_n4  &  wire95 ) | ( n_n4  &  wire729  &  n_n191 ) ;
 assign wire3435 = ( i_7_  &  i_6_  &  n_n159  &  n_n111 ) ;
 assign wire3437 = ( n_n9  &  wire145 ) | ( n_n9  &  n_n186 ) | ( n_n9  &  wire170 ) ;
 assign wire3438 = ( n_n10  &  n_n144 ) | ( n_n10  &  n_n186 ) | ( n_n10  &  wire170 ) ;
 assign wire3439 = ( n_n6  &  wire185 ) | ( n_n6  &  wire270 ) | ( n_n6  &  wire372 ) ;
 assign wire3442 = ( n_n162  &  wire767  &  n_n200  &  n_n220 ) ;
 assign wire3451 = ( n_n33  &  wire52 ) | ( n_n33  &  wire63 ) ;
 assign wire3461 = ( n_n184  &  wire721  &  n_n32 ) ;
 assign wire3469 = ( n_n40  &  wire152 ) | ( n_n40  &  n_n149  &  wire719 ) ;
 assign wire3470 = ( n_n17  &  n_n48  &  wire714  &  wire122 ) ;
 assign wire3471 = ( n_n40  &  wire198 ) | ( n_n40  &  wire289 ) ;
 assign wire3472 = ( n_n17  &  n_n48  &  wire714  &  wire115 ) ;
 assign wire3479 = ( n_n40  &  wire116 ) | ( n_n40  &  wire729  &  n_n156 ) ;
 assign wire3480 = ( n_n17  &  n_n48  &  wire714  &  wire212 ) ;
 assign wire3484 = ( n_n41  &  wire198 ) | ( n_n41  &  wire221 ) | ( n_n41  &  wire18281 ) ;
 assign wire3496 = ( wire172  &  n_n41 ) | ( n_n41  &  n_n191  &  wire719 ) ;
 assign wire3497 = ( n_n40  &  n_n216  &  wire721 ) | ( n_n40  &  n_n216  &  wire725 ) ;
 assign wire3498 = ( n_n41  &  wire256 ) | ( n_n41  &  wire216 ) ;
 assign wire3515 = ( n_n200  &  n_n48  &  n_n220  &  wire1459 ) ;
 assign wire3516 = ( n_n41  &  wire289 ) | ( n_n41  &  wire294 ) | ( n_n41  &  wire18260 ) ;
 assign wire3520 = ( n_n40  &  wire94 ) | ( n_n40  &  wire241 ) | ( n_n40  &  wire18251 ) ;
 assign wire3524 = ( n_n41  &  wire104 ) | ( n_n41  &  wire179 ) | ( n_n41  &  wire324 ) ;
 assign wire3526 = ( n_n41  &  wire243 ) | ( n_n41  &  n_n199  &  wire729 ) ;
 assign wire3527 = ( n_n40  &  wire243 ) | ( n_n40  &  wire341 ) | ( n_n40  &  wire18242 ) ;
 assign wire3531 = ( n_n41  &  wire81 ) | ( n_n41  &  wire206 ) | ( n_n41  &  wire368 ) ;
 assign wire3533 = ( n_n41  &  wire162 ) | ( n_n41  &  wire399 ) | ( n_n41  &  wire341 ) ;
 assign wire3545 = ( n_n40  &  wire162 ) | ( n_n40  &  wire184 ) | ( n_n40  &  wire18230 ) ;
 assign wire3550 = ( n_n40  &  wire122 ) | ( n_n40  &  wire144 ) ;
 assign wire3551 = ( n_n41  &  n_n149  &  wire725 ) ;
 assign wire3563 = ( n_n46  &  wire158 ) | ( n_n46  &  wire133 ) ;
 assign wire3570 = ( n_n46  &  wire171 ) | ( n_n46  &  wire252 ) | ( n_n46  &  wire18194 ) ;
 assign wire3575 = ( n_n46  &  wire135 ) | ( n_n46  &  wire153 ) | ( n_n46  &  wire125 ) ;
 assign wire3580 = ( n_n47  &  wire160 ) | ( n_n47  &  wire171 ) ;
 assign wire3581 = ( n_n46  &  wire242 ) | ( n_n46  &  wire18188 ) ;
 assign wire3588 = ( n_n47  &  wire52 ) | ( n_n47  &  wire139 ) | ( n_n47  &  wire128 ) ;
 assign wire3594 = ( n_n46  &  wire68 ) | ( n_n46  &  wire74 ) ;
 assign wire3601 = ( n_n46  &  wire143 ) | ( n_n46  &  wire154 ) ;
 assign wire3607 = ( n_n18  &  n_n48  &  wire714  &  wire152 ) ;
 assign wire3621 = ( wire253  &  n_n6 ) | ( wire253  &  wire398 ) | ( wire253  &  wire1550 ) ;
 assign wire3622 = ( wire717  &  n_n156  &  wire1550 ) | ( wire717  &  n_n156  &  wire18157 ) ;
 assign wire3624 = ( n_n162  &  n_n19  &  n_n157 ) | ( n_n19  &  n_n157  &  n_n48 ) ;
 assign wire3628 = ( wire253  &  n_n10 ) | ( wire253  &  n_n12 ) ;
 assign wire3629 = ( n_n9  &  n_n151 ) | ( n_n6  &  n_n151 ) | ( n_n151  &  n_n12 ) ;
 assign wire3643 = ( n_n212  &  wire68 ) | ( n_n212  &  wire74 ) ;
 assign wire3653 = ( n_n125  &  wire84 ) | ( n_n125  &  wire205 ) | ( n_n125  &  wire18117 ) ;
 assign wire3658 = ( n_n125  &  wire211 ) | ( n_n125  &  wire272 ) | ( n_n125  &  wire18111 ) ;
 assign wire3662 = ( n_n125  &  wire18102 ) | ( n_n125  &  wire18103 ) | ( n_n125  &  wire18104 ) ;
 assign wire3665 = ( n_n125  &  wire70 ) | ( n_n125  &  wire219 ) | ( n_n125  &  wire18092 ) ;
 assign wire3671 = ( n_n212  &  wire18087 ) | ( n_n212  &  wire18088 ) ;
 assign wire3676 = ( n_n212  &  wire18081 ) | ( n_n212  &  wire18082 ) | ( n_n212  &  wire18083 ) ;
 assign wire3685 = ( n_n108  &  wire18067 ) | ( n_n108  &  wire18068 ) | ( n_n108  &  wire18069 ) ;
 assign wire3690 = ( n_n113  &  wire94 ) | ( n_n113  &  wire184 ) | ( n_n113  &  wire18053 ) ;
 assign wire3696 = ( n_n220  &  n_n111  &  wire1747  &  wire16987 ) ;
 assign wire3700 = ( n_n113  &  wire54 ) | ( n_n113  &  wire268 ) ;
 assign wire3701 = ( wire245  &  n_n125 ) | ( n_n125  &  n_n149  &  wire725 ) ;
 assign wire3702 = ( n_n47  &  wire139 ) | ( n_n47  &  wire128 ) ;
 assign wire3710 = ( n_n220  &  n_n111  &  wire412  &  wire17072 ) ;
 assign wire3723 = ( wire53  &  n_n39 ) | ( n_n39  &  n_n143 ) | ( n_n39  &  wire237 ) ;
 assign wire3747 = ( n_n41  &  wire225 ) | ( n_n41  &  n_n170  &  wire720 ) ;
 assign wire3755 = ( n_n41  &  wire211 ) | ( n_n41  &  wire272 ) | ( n_n41  &  wire17993 ) ;
 assign wire3759 = ( n_n43  &  wire256 ) | ( n_n43  &  wire216 ) ;
 assign wire3767 = ( wire130  &  n_n43 ) | ( n_n43  &  wire222 ) ;
 assign wire3773 = ( n_n47  &  wire17970 ) | ( n_n47  &  wire17971 ) | ( n_n47  &  wire17972 ) ;
 assign wire3774 = ( n_n149  &  n_n126  &  n_n220  &  n_n111 ) ;
 assign wire3810 = ( n_n32  &  wire107 ) | ( n_n184  &  wire720  &  n_n32 ) ;
 assign wire3811 = ( n_n36  &  wire17940 ) | ( n_n36  &  wire17941 ) | ( n_n36  &  wire17942 ) ;
 assign wire3820 = ( n_n31  &  wire55 ) | ( n_n31  &  wire133 ) | ( n_n31  &  wire127 ) ;
 assign wire3828 = ( n_n36  &  wire152 ) | ( n_n36  &  n_n149  &  wire719 ) ;
 assign wire3829 = ( wire157  &  n_n34 ) | ( n_n34  &  wire204 ) | ( n_n34  &  wire17909 ) ;
 assign wire3835 = ( n_n34  &  wire171 ) | ( n_n34  &  wire252 ) | ( n_n34  &  wire17901 ) ;
 assign wire3836 = ( n_n157  &  wire714  &  n_n218  &  wire1814 ) ;
 assign wire3850 = ( n_n34  &  wire242 ) | ( n_n34  &  n_n184  &  wire719 ) ;
 assign wire3851 = ( n_n36  &  wire247 ) | ( n_n36  &  wire160 ) | ( n_n36  &  wire171 ) ;
 assign wire3866 = ( wire132  &  n_n34 ) | ( n_n34  &  wire149 ) | ( n_n34  &  wire46 ) ;
 assign wire3885 = ( i_7_  &  (~ i_6_)  &  n_n19  &  wire817 ) ;
 assign wire3886 = ( i_7_  &  i_6_  &  wire748 ) | ( i_7_  &  i_6_  &  wire733 ) ;
 assign wire3887 = ( i_7_  &  i_6_  &  n_n162  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n162  &  n_n19 ) ;
 assign wire3895 = ( n_n4  &  wire145 ) | ( n_n6  &  wire145 ) | ( n_n5  &  wire145 ) ;
 assign wire3896 = ( n_n9  &  n_n186 ) | ( n_n6  &  n_n186 ) | ( n_n5  &  n_n186 ) ;
 assign wire3897 = ( n_n4  &  n_n191  &  wire717 ) | ( n_n191  &  wire717  &  wire1044 ) ;
 assign wire3899 = ( i_5_  &  n_n159  &  wire231  &  wire17176 ) ;
 assign wire3900 = ( n_n9  &  wire145 ) | ( n_n10  &  wire145 ) | ( wire145  &  n_n12 ) ;
 assign wire3901 = ( n_n14  &  n_n186 ) | ( n_n10  &  n_n186 ) | ( n_n186  &  n_n12 ) ;
 assign wire3957 = ( n_n36  &  wire172 ) | ( n_n36  &  wire80 ) | ( n_n36  &  wire78 ) ;
 assign wire3958 = ( n_n34  &  wire144 ) | ( n_n34  &  wire222 ) | ( n_n34  &  wire17808 ) ;
 assign wire3964 = ( n_n34  &  wire214 ) | ( n_n34  &  wire212 ) ;
 assign wire3973 = ( n_n30  &  wire52 ) | ( n_n30  &  wire129 ) | ( n_n30  &  wire146 ) ;
 assign wire3985 = ( n_n30  &  wire134 ) | ( n_n30  &  wire156 ) ;
 assign wire3990 = ( n_n31  &  wire157 ) | ( n_n31  &  wire80 ) | ( n_n31  &  wire78 ) ;
 assign wire3991 = ( n_n30  &  wire222 ) | ( n_n30  &  wire174 ) | ( n_n30  &  wire17781 ) ;
 assign wire3996 = ( n_n30  &  wire214 ) | ( n_n30  &  wire212 ) ;
 assign wire3997 = ( n_n31  &  n_n191  &  wire719 ) ;
 assign wire3998 = ( n_n197  &  wire143 ) | ( n_n197  &  wire154 ) ;
 assign wire4013 = ( n_n125  &  wire180 ) | ( n_n125  &  n_n190 ) | ( n_n125  &  wire86 ) ;
 assign wire4020 = ( n_n212  &  wire172 ) | ( n_n212  &  n_n191  &  wire719 ) ;
 assign wire4021 = ( n_n197  &  wire214 ) | ( n_n197  &  wire212 ) ;
 assign wire4026 = ( n_n212  &  wire80 ) | ( n_n212  &  wire78 ) ;
 assign wire4027 = ( n_n197  &  n_n59 ) | ( n_n197  &  wire144 ) | ( n_n197  &  wire222 ) ;
 assign wire4043 = ( n_n123  &  wire100 ) | ( n_n123  &  wire215 ) | ( n_n123  &  wire17739 ) ;
 assign wire4048 = ( wire172  &  n_n123 ) | ( n_n138  &  n_n123 ) | ( n_n123  &  wire125 ) ;
 assign wire4060 = ( n_n112  &  wire241 ) | ( n_n112  &  wire273 ) | ( n_n112  &  wire17724 ) ;
 assign wire4064 = ( n_n123  &  wire80 ) | ( n_n123  &  wire78 ) ;
 assign wire4065 = ( wire381  &  n_n125 ) | ( n_n125  &  n_n156  &  wire719 ) ;
 assign wire4067 = ( n_n101  &  wire143 ) | ( n_n101  &  wire154 ) | ( n_n101  &  wire47 ) ;
 assign wire4080 = ( n_n46  &  wire143 ) | ( n_n46  &  wire154 ) ;
 assign wire4088 = ( n_n46  &  wire52 ) | ( n_n46  &  wire129 ) ;
 assign wire4102 = ( n_n42  &  wire52 ) | ( n_n42  &  wire129 ) ;
 assign wire4103 = ( n_n162  &  n_n18  &  wire714  &  wire222 ) ;
 assign wire4104 = ( wire381  &  n_n41 ) | ( n_n41  &  wire160 ) | ( n_n41  &  wire171 ) ;
 assign wire4113 = ( n_n40  &  n_n155 ) | ( n_n40  &  wire125 ) | ( n_n40  &  wire215 ) ;
 assign wire4126 = ( n_n40  &  wire80 ) | ( n_n40  &  wire78 ) ;
 assign wire4130 = ( n_n42  &  wire160 ) | ( n_n42  &  wire171 ) ;
 assign wire4143 = ( n_n40  &  n_n176 ) | ( n_n40  &  wire250 ) | ( n_n40  &  wire100 ) ;
 assign wire4151 = ( n_n17  &  n_n48  &  wire714  &  wire240 ) ;
 assign wire4158 = ( n_n46  &  wire144 ) | ( n_n46  &  wire222 ) | ( n_n46  &  wire17632 ) ;
 assign wire4159 = ( n_n156  &  n_n124  &  n_n220  &  n_n111 ) ;
 assign wire4172 = ( wire172  &  n_n108 ) | ( n_n138  &  n_n108 ) | ( n_n108  &  wire78 ) ;
 assign wire4182 = ( n_n108  &  wire134 ) | ( n_n108  &  wire131 ) ;
 assign wire4185 = ( n_n108  &  wire125 ) | ( n_n108  &  n_n216  &  wire725 ) ;
 assign wire4186 = ( n_n101  &  wire134 ) | ( n_n101  &  wire123 ) | ( n_n101  &  wire17615 ) ;
 assign wire4217 = ( n_n4  &  wire170 ) | ( n_n6  &  wire170 ) | ( n_n5  &  wire170 ) ;
 assign wire4220 = ( i_3_  &  i_4_  &  n_n159  &  wire17591 ) ;
 assign wire4221 = ( n_n4  &  wire717  &  n_n149 ) | ( wire717  &  n_n149  &  wire1527 ) ;
 assign wire4223 = ( n_n162  &  n_n19  &  wire1463 ) | ( n_n19  &  n_n48  &  wire1463 ) ;
 assign wire4228 = ( n_n9  &  wire170 ) | ( n_n10  &  wire170 ) | ( n_n12  &  wire170 ) ;
 assign wire4229 = ( n_n14  &  n_n144 ) | ( n_n10  &  n_n144 ) | ( n_n144  &  n_n12 ) ;
 assign wire4230 = ( wire123  &  n_n200  &  n_n220  &  n_n218 ) ;
 assign wire4233 = ( n_n197  &  wire152 ) | ( n_n197  &  wire17569 ) ;
 assign wire4234 = ( n_n212  &  wire245 ) | ( n_n212  &  wire144 ) | ( n_n212  &  wire17570 ) ;
 assign wire4252 = ( n_n149  &  n_n126  &  n_n220  &  n_n111 ) ;
 assign wire4253 = ( n_n156  &  n_n124  &  n_n220  &  n_n111 ) ;
 assign wire4260 = ( n_n46  &  wire173 ) | ( n_n46  &  wire204 ) ;
 assign wire4263 = ( n_n124  &  n_n48  &  n_n220  &  wire249 ) ;
 assign wire4285 = ( n_n40  &  wire173 ) | ( n_n40  &  wire204 ) ;
 assign wire4286 = ( wire157  &  n_n41 ) | ( n_n41  &  wire152 ) | ( n_n41  &  wire17535 ) ;
 assign wire4291 = ( n_n40  &  wire215 ) | ( n_n40  &  wire720  &  n_n156 ) ;
 assign wire4320 = ( n_n149  &  n_n220  &  n_n111  &  wire16987 ) ;
 assign wire4323 = ( n_n123  &  wire173 ) | ( n_n123  &  wire204 ) ;
 assign wire4324 = ( n_n125  &  wire152 ) | ( n_n125  &  wire17468 ) ;
 assign wire4334 = ( n_n46  &  wire205 ) | ( n_n46  &  wire215 ) | ( n_n46  &  wire17498 ) ;
 assign wire4341 = ( n_n18  &  wire800  &  n_n48  &  wire714 ) ;
 assign wire4343 = ( n_n108  &  wire152 ) | ( n_n108  &  n_n149  &  wire719 ) ;
 assign wire4344 = ( wire157  &  n_n101 ) | ( n_n101  &  wire17480 ) ;
 assign wire4354 = ( n_n200  &  n_n156  &  n_n220  &  n_n111 ) ;
 assign wire4355 = ( n_n149  &  n_n220  &  n_n111  &  wire17072 ) ;
 assign wire4365 = ( n_n101  &  wire204 ) | ( n_n101  &  wire205 ) ;
 assign wire4372 = ( n_n162  &  n_n126  &  n_n220  &  wire141 ) ;
 assign wire4376 = ( n_n123  &  n_n155 ) | ( n_n123  &  wire215 ) | ( n_n123  &  wire805 ) ;
 assign wire4382 = ( n_n125  &  wire215 ) | ( n_n125  &  wire720  &  n_n156 ) ;
 assign wire4393 = ( wire90  &  n_n123 ) | ( n_n123  &  wire155 ) | ( n_n123  &  wire205 ) ;
 assign wire4395 = ( n_n34  &  wire152 ) | ( n_n34  &  wire17447 ) ;
 assign wire4396 = ( n_n36  &  wire245 ) | ( n_n36  &  wire144 ) | ( n_n36  &  wire17448 ) ;
 assign wire4419 = ( n_n30  &  wire152 ) | ( n_n30  &  wire125 ) | ( n_n30  &  wire17428 ) ;
 assign wire4420 = ( n_n162  &  n_n157  &  wire714  &  wire144 ) ;
 assign wire4427 = ( n_n31  &  wire245 ) | ( n_n31  &  n_n149  &  wire725 ) ;
 assign wire4428 = ( n_n162  &  n_n220  &  n_n35  &  wire144 ) ;
 assign wire4429 = ( n_n31  &  wire55 ) | ( n_n31  &  wire133 ) | ( n_n31  &  wire127 ) ;
 assign wire4430 = ( n_n30  &  wire156 ) | ( n_n30  &  wire133 ) | ( n_n30  &  wire17426 ) ;
 assign wire4434 = ( n_n33  &  wire234 ) | ( n_n33  &  wire84 ) | ( n_n33  &  wire17416 ) ;
 assign wire4453 = ( n_n123  &  wire93 ) | ( n_n123  &  wire177 ) | ( n_n123  &  wire17391 ) ;
 assign wire4454 = ( n_n125  &  wire93 ) | ( n_n125  &  wire362 ) | ( n_n125  &  wire17391 ) ;
 assign wire4458 = ( n_n123  &  wire94 ) | ( n_n184  &  n_n123  &  wire729 ) ;
 assign wire4459 = ( n_n125  &  wire94 ) | ( n_n125  &  wire177 ) ;
 assign wire4460 = ( n_n212  &  wire299 ) | ( n_n212  &  wire17385 ) ;
 assign wire4470 = ( n_n125  &  wire164 ) | ( n_n125  &  wire358 ) ;
 assign wire4474 = ( n_n212  &  wire193 ) | ( n_n212  &  wire196 ) | ( n_n212  &  wire306 ) ;
 assign wire4475 = ( n_n197  &  wire168 ) | ( n_n197  &  wire193 ) | ( n_n197  &  wire196 ) ;
 assign wire4481 = ( n_n197  &  wire130 ) | ( n_n197  &  wire304 ) | ( n_n197  &  wire306 ) ;
 assign wire4485 = ( n_n212  &  wire308 ) | ( n_n212  &  wire201 ) ;
 assign wire4486 = ( n_n197  &  wire200 ) | ( n_n197  &  wire201 ) | ( n_n197  &  wire299 ) ;
 assign wire4491 = ( n_n101  &  n_n210 ) | ( n_n101  &  wire374 ) | ( n_n101  &  wire17361 ) ;
 assign wire4496 = ( n_n108  &  wire307 ) | ( n_n108  &  n_n191  &  wire722 ) ;
 assign wire4500 = ( n_n108  &  wire69 ) | ( n_n108  &  wire229 ) | ( n_n108  &  wire17357 ) ;
 assign wire4503 = ( n_n101  &  wire351 ) | ( n_n101  &  wire722  &  n_n149 ) ;
 assign wire4504 = ( n_n108  &  wire90 ) | ( n_n108  &  wire377 ) ;
 assign wire4505 = ( n_n101  &  wire202 ) | ( n_n101  &  wire17349 ) | ( n_n101  &  wire17350 ) ;
 assign wire4506 = ( n_n108  &  wire265 ) | ( n_n108  &  wire17352 ) | ( n_n108  &  wire17353 ) ;
 assign wire4508 = ( n_n101  &  wire307 ) | ( n_n101  &  n_n191  &  wire722 ) ;
 assign wire4509 = ( n_n108  &  wire62 ) | ( n_n108  &  wire202 ) ;
 assign wire4510 = ( n_n40  &  n_n168 ) | ( n_n40  &  wire229 ) | ( n_n40  &  wire17343 ) ;
 assign wire4520 = ( n_n41  &  wire307 ) | ( n_n41  &  n_n191  &  wire722 ) ;
 assign wire4523 = ( n_n40  &  wire265 ) | ( n_n40  &  wire17336 ) ;
 assign wire4526 = ( n_n41  &  n_n196 ) | ( n_n41  &  wire263 ) | ( n_n41  &  wire374 ) ;
 assign wire4531 = ( n_n42  &  wire93 ) | ( n_n42  &  n_n184  &  wire725 ) ;
 assign wire4539 = ( n_n36  &  wire117 ) | ( n_n36  &  wire366 ) | ( n_n36  &  wire17324 ) ;
 assign wire4544 = ( n_n34  &  wire93 ) | ( n_n34  &  wire301 ) | ( n_n34  &  wire17317 ) ;
 assign wire4545 = ( n_n36  &  wire94 ) | ( n_n36  &  wire120 ) | ( n_n36  &  wire17319 ) ;
 assign wire4548 = ( n_n34  &  wire94 ) | ( n_n34  &  wire177 ) ;
 assign wire4549 = ( n_n36  &  wire93 ) | ( n_n36  &  wire729  &  n_n191 ) ;
 assign wire4550 = ( n_n34  &  wire369 ) | ( n_n34  &  wire729  &  n_n177 ) ;
 assign wire4551 = ( n_n36  &  wire116 ) | ( n_n36  &  wire371 ) ;
 assign wire4554 = ( n_n34  &  wire115 ) | ( n_n34  &  wire17310 ) | ( n_n34  &  wire17313 ) ;
 assign wire4558 = ( wire820  &  n_n157  &  wire714  &  n_n218 ) ;
 assign wire4561 = ( wire979  &  wire243 ) | ( n_n199  &  wire729  &  wire979 ) ;
 assign wire4562 = ( n_n34  &  wire164 ) | ( n_n34  &  wire358 ) ;
 assign wire4568 = ( n_n36  &  wire164 ) | ( n_n36  &  wire358 ) ;
 assign wire4569 = ( i_15_  &  n_n34  &  n_n199  &  n_n211 ) | ( (~ i_15_)  &  n_n34  &  n_n199  &  n_n211 ) ;
 assign wire4572 = ( n_n41  &  wire60 ) | ( n_n41  &  wire351 ) | ( n_n41  &  wire17292 ) ;
 assign wire4573 = ( n_n40  &  wire377 ) | ( n_n40  &  wire17294 ) | ( n_n40  &  wire17295 ) ;
 assign wire4576 = ( n_n40  &  wire351 ) | ( n_n40  &  wire722  &  n_n149 ) ;
 assign wire4581 = ( n_n38  &  wire1120 ) | ( n_n38  &  wire17287 ) ;
 assign wire4591 = ( n_n126  &  n_n48  &  n_n220  &  wire1116 ) ;
 assign wire4602 = ( n_n123  &  wire120 ) | ( n_n123  &  wire729  &  n_n177 ) ;
 assign wire4619 = ( n_n113  &  wire62 ) | ( n_n113  &  wire202 ) ;
 assign wire4620 = ( n_n112  &  wire307 ) | ( n_n112  &  n_n191  &  wire722 ) ;
 assign wire4628 = ( n_n30  &  wire149 ) | ( n_n30  &  wire200 ) | ( n_n30  &  wire201 ) ;
 assign wire4638 = ( n_n31  &  wire176 ) | ( n_n31  &  n_n59 ) | ( n_n31  &  wire299 ) ;
 assign wire4639 = ( n_n30  &  wire158 ) | ( n_n30  &  wire308 ) | ( n_n30  &  wire17238 ) ;
 assign wire4643 = ( n_n162  &  n_n220  &  n_n35  &  wire899 ) ;
 assign wire4644 = ( n_n31  &  wire130 ) | ( n_n31  &  wire304 ) | ( n_n31  &  wire306 ) ;
 assign wire4649 = ( n_n32  &  wire62 ) | ( n_n32  &  wire202 ) ;
 assign wire4651 = ( n_n33  &  wire229 ) | ( n_n33  &  wire307 ) | ( n_n33  &  wire17224 ) ;
 assign wire4655 = ( n_n33  &  n_n147 ) | ( n_n33  &  wire69 ) | ( n_n33  &  wire351 ) ;
 assign wire4658 = ( wire168  &  wire968 ) | ( wire968  &  wire193 ) | ( wire968  &  wire196 ) ;
 assign wire4659 = ( n_n33  &  n_n55 ) | ( n_n33  &  wire51 ) | ( n_n33  &  wire17215 ) ;
 assign wire4662 = ( n_n46  &  wire149 ) | ( n_n46  &  wire200 ) | ( n_n46  &  wire201 ) ;
 assign wire4663 = ( n_n47  &  wire308 ) | ( n_n47  &  wire131 ) | ( n_n47  &  wire201 ) ;
 assign wire4669 = ( wire896  &  wire301 ) | ( n_n184  &  wire729  &  wire896 ) ;
 assign wire4671 = ( n_n43  &  wire94 ) | ( n_n43  &  wire177 ) ;
 assign wire4676 = ( n_n42  &  wire94 ) | ( n_n42  &  wire177 ) ;
 assign wire4680 = ( n_n46  &  wire308 ) | ( n_n46  &  wire418 ) | ( n_n46  &  wire890 ) ;
 assign wire4684 = ( wire168  &  n_n47 ) | ( n_n47  &  wire193 ) | ( n_n47  &  wire196 ) ;
 assign wire4685 = ( n_n46  &  wire193 ) | ( n_n46  &  wire196 ) ;
 assign wire4701 = ( n_n47  &  wire200 ) | ( n_n47  &  wire304 ) | ( n_n47  &  wire306 ) ;
 assign wire4735 = ( n_n101  &  wire100 ) | ( n_n101  &  n_n177  &  wire720 ) ;
 assign wire4739 = ( n_n212  &  wire68 ) | ( n_n212  &  wire74 ) ;
 assign wire4740 = ( n_n197  &  wire143 ) | ( n_n197  &  wire154 ) ;
 assign wire4743 = ( n_n123  &  wire224 ) | ( n_n123  &  wire250 ) | ( n_n123  &  wire57 ) ;
 assign wire4750 = ( n_n123  &  wire141 ) | ( n_n123  &  n_n216  &  wire719 ) ;
 assign wire4751 = ( n_n126  &  n_n220  &  n_n218  &  wire153 ) ;
 assign wire4752 = ( n_n125  &  wire225 ) | ( n_n125  &  n_n170  &  wire720 ) ;
 assign wire4753 = ( n_n123  &  wire100 ) | ( n_n123  &  wire225 ) | ( n_n123  &  wire17132 ) ;
 assign wire4765 = ( n_n123  &  wire85 ) | ( n_n123  &  n_n216  &  wire720 ) ;
 assign wire4768 = ( n_n123  &  wire218 ) | ( n_n123  &  n_n199  &  wire725 ) ;
 assign wire4771 = ( wire137  &  n_n197 ) | ( n_n197  &  wire146 ) ;
 assign wire4780 = ( n_n126  &  n_n220  &  n_n218  &  wire219 ) ;
 assign wire4786 = ( n_n17  &  wire714  &  wire247  &  n_n218 ) ;
 assign wire4805 = ( n_n46  &  wire208 ) | ( n_n46  &  wire86 ) | ( n_n46  &  wire148 ) ;
 assign wire4818 = ( n_n18  &  n_n48  &  wire714  &  wire1030 ) ;
 assign wire4819 = ( n_n46  &  wire100 ) | ( n_n46  &  wire225 ) | ( n_n46  &  wire17089 ) ;
 assign wire4820 = ( n_n47  &  wire85 ) | ( n_n47  &  n_n216  &  wire720 ) ;
 assign wire4821 = ( n_n108  &  wire150 ) | ( n_n108  &  n_n170  &  wire719 ) ;
 assign wire4822 = ( n_n101  &  wire182 ) | ( n_n101  &  wire17074 ) ;
 assign wire4827 = ( n_n200  &  n_n177  &  n_n220  &  n_n111 ) ;
 assign wire4828 = ( n_n170  &  n_n220  &  n_n111  &  wire17072 ) ;
 assign wire4829 = ( n_n47  &  wire142 ) | ( n_n47  &  wire180 ) | ( n_n47  &  wire86 ) ;
 assign wire4830 = ( n_n46  &  n_n199  &  wire720 ) ;
 assign wire4831 = ( n_n101  &  wire224 ) | ( n_n101  &  wire209 ) ;
 assign wire4832 = ( n_n108  &  wire182 ) | ( n_n108  &  n_n57 ) | ( n_n108  &  wire141 ) ;
 assign wire4838 = ( n_n162  &  n_n124  &  n_n220  &  wire1862 ) ;
 assign wire4839 = ( n_n108  &  wire135 ) | ( n_n108  &  wire153 ) ;
 assign wire4842 = ( n_n40  &  n_n214 ) | ( n_n40  &  wire108 ) | ( n_n40  &  wire258 ) ;
 assign wire4857 = ( n_n47  &  wire182 ) | ( n_n47  &  n_n177  &  wire725 ) ;
 assign wire4858 = ( n_n161  &  n_n48  &  n_n220  &  wire209 ) ;
 assign wire4859 = ( n_n47  &  wire135 ) | ( n_n47  &  wire153 ) ;
 assign wire4860 = ( n_n46  &  wire141 ) | ( n_n46  &  wire17052 ) ;
 assign wire4863 = ( n_n38  &  wire53 ) | ( n_n38  &  wire237 ) ;
 assign wire4864 = ( n_n39  &  wire724  &  n_n177 ) ;
 assign wire4869 = ( n_n39  &  wire237 ) | ( n_n39  &  wire724  &  n_n170 ) ;
 assign wire4870 = ( n_n124  &  n_n48  &  n_n220  &  wire104 ) ;
 assign wire4888 = ( n_n157  &  wire714  &  wire151  &  n_n218 ) ;
 assign wire4890 = ( n_n41  &  wire225 ) | ( n_n41  &  n_n170  &  wire720 ) ;
 assign wire4891 = ( n_n40  &  wire250 ) | ( n_n40  &  wire100 ) | ( n_n40  &  wire69 ) ;
 assign wire4900 = ( n_n17  &  n_n48  &  wire714  &  wire150 ) ;
 assign wire4904 = ( n_n40  &  wire141 ) | ( n_n40  &  n_n216  &  wire719 ) ;
 assign wire4905 = ( n_n17  &  n_n48  &  wire714  &  wire153 ) ;
 assign wire4908 = ( n_n40  &  wire218 ) | ( n_n40  &  n_n199  &  wire725 ) ;
 assign wire4919 = ( n_n40  &  wire219 ) | ( n_n40  &  n_n199  &  wire720 ) ;
 assign wire4924 = ( n_n108  &  wire100 ) | ( n_n108  &  n_n177  &  wire720 ) ;
 assign wire4933 = ( n_n108  &  wire224 ) | ( n_n108  &  wire57 ) ;
 assign wire4934 = ( n_n101  &  n_n170  &  wire720 ) ;
 assign wire4935 = ( n_n101  &  n_n214 ) | ( n_n101  &  wire70 ) | ( n_n101  &  wire258 ) ;
 assign wire4937 = ( n_n101  &  wire219 ) | ( n_n101  &  wire108 ) ;
 assign wire4941 = ( n_n125  &  wire150 ) | ( n_n125  &  n_n170  &  wire719 ) ;
 assign wire4942 = ( n_n123  &  wire182 ) | ( n_n123  &  wire209 ) | ( n_n123  &  wire16988 ) ;
 assign wire4948 = ( n_n170  &  n_n220  &  n_n111  &  wire16987 ) ;
 assign wire4950 = ( n_n199  &  n_n220  &  n_n111  &  wire16987 ) ;
 assign wire4953 = ( n_n30  &  wire126 ) | ( n_n30  &  wire150 ) | ( n_n30  &  wire16972 ) ;
 assign wire4960 = ( n_n31  &  wire80 ) | ( n_n31  &  wire78 ) ;
 assign wire4961 = ( n_n30  &  wire146 ) | ( n_n30  &  wire125 ) | ( n_n30  &  wire16964 ) ;
 assign wire4965 = ( n_n30  &  wire135 ) | ( n_n30  &  wire153 ) ;
 assign wire4966 = ( n_n31  &  wire247 ) | ( n_n31  &  n_n199  &  wire719 ) ;
 assign wire4974 = ( wire132  &  n_n34 ) | ( n_n34  &  wire149 ) ;
 assign wire4981 = ( n_n34  &  wire150 ) | ( n_n34  &  wire16946 ) ;
 assign wire4982 = ( n_n157  &  wire714  &  n_n218  &  wire942 ) ;
 assign wire4986 = ( n_n157  &  wire714  &  wire247  &  n_n218 ) ;
 assign wire4993 = ( n_n33  &  wire225 ) | ( n_n33  &  wire148 ) | ( n_n33  &  wire16940 ) ;
 assign wire4998 = ( wire140  &  n_n124  &  n_n48  &  n_n220 ) ;
 assign wire5022 = ( n_n38  &  wire235 ) | ( n_n38  &  wire236 ) ;
 assign wire5023 = ( wire140  &  n_n126  &  n_n48  &  n_n220 ) ;
 assign wire5024 = ( n_n39  &  wire235 ) | ( n_n39  &  wire236 ) ;
 assign wire5025 = ( n_n124  &  n_n48  &  n_n220  &  wire244 ) ;
 assign wire5026 = ( n_n65  &  n_n5 ) | ( n_n65  &  wire398 ) | ( n_n65  &  wire16908 ) ;
 assign wire5027 = ( wire343  &  n_n5 ) | ( wire343  &  wire16908 ) | ( wire343  &  wire16909 ) ;
 assign wire5032 = ( wire729  &  n_n156  &  n_n12 ) ;
 assign wire5057 = ( n_n35  &  wire5067  &  wire16861 ) | ( n_n35  &  wire5068  &  wire16861 ) ;
 assign wire5067 = ( n_n184  &  wire725  &  n_n111 ) ;
 assign wire5068 = ( n_n184  &  wire717  &  n_n48 ) ;
 assign wire16857 = ( n_n162  &  n_n163  &  n_n200 ) ;
 assign wire16861 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign wire16863 = ( i_3_  &  n_n219 ) | ( n_n157  &  n_n219  &  n_n111 ) ;
 assign wire16865 = ( n_n7263 ) | ( n_n7264 ) | ( n_n135  &  wire16857 ) ;
 assign wire16866 = ( wire16863 ) | ( wire463 ) ;
 assign wire16867 = ( n_n3389 ) | ( n_n7252 ) | ( n_n7262 ) ;
 assign wire16870 = ( wire388 ) | ( wire16865 ) | ( wire16867 ) ;
 assign wire16871 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16872 = ( wire428 ) | ( wire16871 ) ;
 assign wire16876 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign wire16877 = ( n_n5144 ) | ( n_n184  &  wire725  &  wire16857 ) ;
 assign wire16880 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire16884 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n218 ) ;
 assign wire16885 = ( i_3_  &  (~ i_1_)  &  i_2_  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16886 = ( n_n3276 ) | ( wire462 ) | ( wire16884 ) | ( wire16885 ) ;
 assign wire16888 = ( i_3_  &  (~ i_1_)  &  i_2_  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire16889 = ( n_n17  &  n_n219  &  n_n218 ) | ( n_n17  &  n_n219  &  n_n111 ) ;
 assign wire16890 = ( n_n162  &  n_n18  &  n_n219 ) | ( n_n18  &  n_n219  &  n_n111 ) ;
 assign wire16892 = ( n_n7263 ) | ( wire711 ) | ( n_n7264 ) ;
 assign wire16896 = ( wire388 ) | ( n_n2948 ) | ( wire16889 ) | ( wire16890 ) ;
 assign wire16897 = ( wire569 ) | ( wire16888 ) | ( wire16892 ) | ( wire16896 ) ;
 assign wire16898 = ( i_2_  &  (~ i_0_) ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  i_0_ ) | ( i_3_  &  (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign wire16908 = ( n_n48  &  n_n35  &  n_n159 ) | ( n_n35  &  n_n159  &  n_n111 ) ;
 assign wire16909 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire16910 = ( n_n5144 ) | ( n_n9  &  wire729  &  n_n156 ) ;
 assign wire16911 = ( wire5032 ) | ( wire16910 ) | ( wire1042  &  wire1041 ) ;
 assign wire16924 = ( n_n5144 ) | ( n_n39  &  n_n177  &  wire719 ) ;
 assign wire16929 = ( wire390 ) | ( wire393 ) | ( wire712 ) | ( wire16924 ) ;
 assign wire16930 = ( n_n969 ) | ( n_n519 ) | ( n_n4597 ) | ( wire4998 ) ;
 assign wire16933 = ( n_n373 ) | ( n_n374 ) | ( wire16929 ) | ( wire16930 ) ;
 assign wire16936 = ( i_15_  &  n_n170  &  n_n215 ) | ( (~ i_15_)  &  n_n170  &  n_n215 ) ;
 assign wire16940 = ( wire186 ) | ( wire208 ) | ( wire69 ) | ( wire16936 ) ;
 assign wire16941 = ( n_n33  &  n_n132 ) | ( n_n34  &  wire78 ) ;
 assign wire16943 = ( wire443 ) | ( wire16941 ) | ( n_n31  &  wire143 ) ;
 assign wire16946 = ( n_n177  &  wire719 ) | ( n_n170  &  wire719 ) | ( n_n177  &  wire728 ) ;
 assign wire16950 = ( wire4981 ) | ( n_n34  &  n_n63 ) | ( n_n34  &  wire125 ) ;
 assign wire16952 = ( n_n34  &  wire147 ) | ( n_n34  &  wire181 ) ;
 assign wire16953 = ( wire137  &  n_n36 ) | ( n_n34  &  wire126 ) ;
 assign wire16954 = ( n_n36  &  wire146 ) | ( n_n36  &  wire46 ) | ( n_n36  &  wire131 ) ;
 assign wire16957 = ( n_n36  &  wire147 ) | ( n_n36  &  wire125 ) ;
 assign wire16960 = ( wire607 ) | ( wire16957 ) | ( n_n36  &  wire149 ) ;
 assign wire16961 = ( wire584 ) | ( wire606 ) | ( wire16960 ) ;
 assign wire16962 = ( n_n4169 ) | ( n_n4419 ) | ( wire4982 ) | ( wire16950 ) ;
 assign wire16964 = ( n_n170  &  wire719 ) | ( n_n216  &  wire725 ) ;
 assign wire16966 = ( n_n31  &  wire125 ) | ( n_n30  &  wire131 ) ;
 assign wire16968 = ( wire655 ) | ( wire4961 ) | ( wire4965 ) | ( wire4966 ) ;
 assign wire16972 = ( wire149 ) | ( wire147 ) | ( wire80 ) | ( wire78 ) ;
 assign wire16974 = ( n_n3510 ) | ( n_n31  &  n_n55 ) | ( n_n31  &  wire252 ) ;
 assign wire16975 = ( wire690 ) | ( wire4953 ) | ( n_n31  &  wire149 ) ;
 assign wire16976 = ( wire4960 ) | ( wire16966 ) | ( wire16968 ) | ( wire16974 ) ;
 assign wire16980 = ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire720 ) ;
 assign wire16987 = ( i_7_  &  i_8_  &  i_6_ ) ;
 assign wire16988 = ( n_n170  &  wire721 ) | ( n_n177  &  wire725 ) | ( n_n170  &  wire725 ) ;
 assign wire16990 = ( n_n125  &  n_n57 ) | ( n_n108  &  n_n214 ) ;
 assign wire16991 = ( n_n5739 ) | ( n_n5743 ) | ( wire4948 ) | ( wire4950 ) ;
 assign wire16993 = ( wire4941 ) | ( wire16990 ) | ( wire16991 ) ;
 assign wire16994 = ( wire4942 ) | ( n_n4904 ) ;
 assign wire16995 = ( n_n108  &  wire250 ) | ( n_n101  &  wire86 ) ;
 assign wire16996 = ( wire4924 ) | ( n_n101  &  wire208 ) ;
 assign wire16997 = ( n_n5033 ) | ( wire4937 ) | ( wire16995 ) ;
 assign wire17000 = ( n_n4900 ) | ( wire4933 ) | ( wire4934 ) | ( wire16997 ) ;
 assign wire17001 = ( wire544 ) | ( wire16993 ) | ( wire16994 ) | ( wire16996 ) ;
 assign wire17003 = ( n_n41  &  wire180 ) | ( n_n41  &  n_n202 ) | ( n_n41  &  n_n102 ) ;
 assign wire17007 = ( n_n41  &  n_n198 ) | ( n_n41  &  wire70 ) | ( n_n40  &  wire70 ) ;
 assign wire17013 = ( wire397 ) | ( wire361 ) | ( n_n40  &  wire180 ) ;
 assign wire17014 = ( wire696 ) | ( n_n41  &  n_n176 ) | ( n_n41  &  wire100 ) ;
 assign wire17016 = ( n_n41  &  wire141 ) | ( n_n41  &  wire135 ) ;
 assign wire17018 = ( n_n5060 ) | ( n_n5059 ) | ( n_n5058 ) | ( wire4900 ) ;
 assign wire17019 = ( wire4904 ) | ( wire4905 ) | ( wire4908 ) | ( wire17016 ) ;
 assign wire17023 = ( wire518 ) | ( wire4890 ) | ( n_n41  &  n_n142 ) ;
 assign wire17025 = ( wire653 ) | ( wire694 ) | ( wire4891 ) | ( wire17023 ) ;
 assign wire17028 = ( n_n34  &  wire168 ) | ( n_n34  &  wire74 ) ;
 assign wire17033 = ( n_n34  &  wire143 ) | ( n_n34  &  wire154 ) | ( n_n34  &  wire47 ) ;
 assign wire17034 = ( n_n34  &  wire68 ) | ( n_n36  &  wire143 ) ;
 assign wire17035 = ( n_n34  &  wire151 ) | ( n_n36  &  wire181 ) ;
 assign wire17038 = ( n_n38  &  n_n84 ) | ( n_n39  &  n_n132 ) ;
 assign wire17039 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n134 ) | ( n_n38  &  n_n132 ) ;
 assign wire17041 = ( n_n4597 ) | ( wire17038 ) | ( wire17039 ) ;
 assign wire17042 = ( n_n40  &  n_n57 ) | ( n_n39  &  wire104 ) ;
 assign wire17044 = ( n_n38  &  wire279 ) | ( n_n39  &  wire279 ) ;
 assign wire17045 = ( n_n974 ) | ( wire17042 ) | ( wire182  &  n_n40 ) ;
 assign wire17047 = ( wire4863 ) | ( wire4864 ) | ( wire4869 ) | ( wire4870 ) ;
 assign wire17049 = ( wire4888 ) | ( wire17028 ) | ( wire17044 ) | ( wire17047 ) ;
 assign wire17050 = ( wire597 ) | ( wire620 ) | ( wire17041 ) | ( wire17045 ) ;
 assign wire17052 = ( n_n216  &  wire719 ) | ( n_n199  &  wire725 ) ;
 assign wire17053 = ( n_n47  &  n_n142 ) | ( n_n46  &  wire57 ) ;
 assign wire17055 = ( n_n5103 ) | ( wire652 ) | ( wire17053 ) ;
 assign wire17056 = ( wire4857 ) | ( wire4858 ) | ( wire4859 ) | ( wire4860 ) ;
 assign wire17058 = ( n_n6271 ) | ( n_n6270 ) | ( n_n46  &  n_n57 ) ;
 assign wire17060 = ( n_n6266 ) | ( n_n6268 ) | ( wire666 ) | ( wire17058 ) ;
 assign wire17061 = ( wire549 ) | ( wire4919 ) | ( wire17003 ) ;
 assign wire17063 = ( wire621 ) | ( wire17055 ) | ( wire17056 ) ;
 assign wire17064 = ( wire17060 ) | ( wire17061 ) | ( wire17063 ) ;
 assign wire17067 = ( n_n108  &  n_n142 ) | ( n_n101  &  wire57 ) ;
 assign wire17070 = ( wire4831 ) | ( n_n101  &  wire218 ) | ( n_n101  &  wire141 ) ;
 assign wire17071 = ( wire4832 ) | ( wire4838 ) | ( wire4839 ) | ( wire17067 ) ;
 assign wire17072 = ( i_7_  &  i_8_  &  (~ i_6_) ) ;
 assign wire17074 = ( n_n170  &  wire721 ) | ( n_n177  &  wire725 ) | ( n_n170  &  wire725 ) ;
 assign wire17076 = ( wire445 ) | ( wire446 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire17079 = ( wire4820 ) | ( wire4821 ) | ( wire4822 ) | ( wire17076 ) ;
 assign wire17081 = ( wire85 ) | ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) ;
 assign wire17082 = ( n_n4641 ) | ( n_n47  &  wire1840 ) ;
 assign wire17083 = ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) | ( n_n170  &  wire720 ) ;
 assign wire17089 = ( n_n176 ) | ( wire224 ) | ( wire250 ) | ( wire69 ) ;
 assign wire17093 = ( n_n1606 ) | ( n_n46  &  wire142 ) | ( n_n46  &  wire180 ) ;
 assign wire17094 = ( wire4805 ) | ( n_n47  &  wire1170 ) ;
 assign wire17096 = ( wire4818 ) | ( wire4819 ) | ( wire17093 ) | ( wire17094 ) ;
 assign wire17100 = ( n_n212  &  wire151 ) | ( n_n212  &  wire181 ) ;
 assign wire17102 = ( n_n212  &  wire168 ) | ( n_n197  &  wire47 ) ;
 assign wire17106 = ( n_n197  &  n_n63 ) | ( n_n125  &  n_n214 ) ;
 assign wire17108 = ( wire422 ) | ( wire17106 ) | ( n_n197  &  wire125 ) ;
 assign wire17109 = ( n_n197  &  wire797 ) | ( n_n212  &  wire796 ) ;
 assign wire17114 = ( wire538 ) | ( n_n125  &  wire180 ) | ( n_n125  &  wire86 ) ;
 assign wire17115 = ( n_n4674 ) | ( wire4780 ) | ( n_n123  &  wire1853 ) ;
 assign wire17116 = ( n_n212  &  wire149 ) | ( n_n197  &  wire131 ) ;
 assign wire17117 = ( n_n197  &  wire46 ) | ( n_n212  &  wire125 ) ;
 assign wire17119 = ( n_n4686 ) | ( wire704 ) | ( wire4786 ) | ( wire17117 ) ;
 assign wire17120 = ( wire4771 ) | ( wire17116 ) | ( wire17119 ) ;
 assign wire17121 = ( wire17108 ) | ( wire17109 ) | ( wire17114 ) | ( wire17115 ) ;
 assign wire17122 = ( n_n125  &  wire141 ) | ( n_n125  &  wire135 ) ;
 assign wire17123 = ( n_n123  &  wire142 ) | ( n_n125  &  wire70 ) ;
 assign wire17125 = ( n_n123  &  n_n169 ) | ( n_n125  &  n_n176 ) ;
 assign wire17127 = ( n_n123  &  wire180 ) | ( n_n125  &  wire100 ) ;
 assign wire17128 = ( wire17125 ) | ( wire17127 ) | ( n_n123  &  wire86 ) ;
 assign wire17129 = ( wire394 ) | ( wire4765 ) | ( wire17123 ) ;
 assign wire17132 = ( wire208 ) | ( wire69 ) | ( wire148 ) ;
 assign wire17134 = ( n_n1708 ) | ( wire698 ) | ( wire4752 ) ;
 assign wire17136 = ( n_n125  &  wire182 ) | ( n_n125  &  n_n216  &  wire719 ) ;
 assign wire17137 = ( wire4768 ) | ( wire17122 ) | ( wire17136 ) ;
 assign wire17139 = ( wire4743 ) | ( wire4750 ) | ( wire4751 ) | ( wire17137 ) ;
 assign wire17140 = ( wire4753 ) | ( wire17128 ) | ( wire17129 ) | ( wire17134 ) ;
 assign wire17141 = ( wire132  &  n_n212 ) | ( n_n197  &  wire149 ) ;
 assign wire17145 = ( wire17141 ) | ( wire132  &  n_n197 ) | ( n_n197  &  wire181 ) ;
 assign wire17146 = ( wire557 ) | ( wire648 ) | ( wire504 ) | ( wire578 ) ;
 assign wire17149 = ( n_n4441 ) | ( wire575 ) | ( wire17145 ) | ( wire17146 ) ;
 assign wire17150 = ( wire17120 ) | ( wire17121 ) | ( wire17139 ) | ( wire17140 ) ;
 assign wire17152 = ( n_n101  &  wire225 ) | ( n_n108  &  wire225 ) | ( n_n101  &  wire148 ) ;
 assign wire17153 = ( n_n5011 ) | ( wire591 ) | ( n_n101  &  wire250 ) ;
 assign wire17154 = ( wire4735 ) | ( wire17152 ) | ( n_n108  &  wire69 ) ;
 assign wire17156 = ( n_n4206 ) | ( wire17070 ) | ( wire17071 ) | ( wire17079 ) ;
 assign wire17158 = ( wire543 ) | ( wire17000 ) | ( wire17001 ) | ( wire17096 ) ;
 assign wire17159 = ( wire17153 ) | ( wire17154 ) | ( wire17156 ) | ( wire17158 ) ;
 assign wire17164 = ( n_n31  &  wire151 ) | ( n_n31  &  wire181 ) ;
 assign wire17166 = ( n_n5144 ) | ( n_n30  &  wire181 ) ;
 assign wire17169 = ( wire17166 ) | ( n_n31  &  wire137 ) | ( n_n31  &  wire46 ) ;
 assign wire17170 = ( n_n4161 ) | ( wire695 ) | ( n_n30  &  wire132 ) ;
 assign wire17172 = ( wire599 ) | ( wire4993 ) | ( wire16943 ) ;
 assign wire17174 = ( wire16961 ) | ( wire16962 ) | ( wire16975 ) | ( wire16976 ) ;
 assign wire17175 = ( wire17169 ) | ( wire17170 ) | ( wire17172 ) | ( wire17174 ) ;
 assign wire17176 = ( i_4_  &  i_3_ ) ;
 assign wire17178 = ( n_n47  &  wire129 ) | ( n_n47  &  wire130 ) ;
 assign wire17181 = ( n_n135  &  n_n101 ) | ( n_n135  &  n_n108 ) | ( n_n101  &  wire1179 ) ;
 assign wire17184 = ( n_n101  &  wire90 ) | ( n_n101  &  n_n61 ) | ( n_n108  &  n_n61 ) ;
 assign wire17185 = ( wire17181 ) | ( wire17184 ) | ( n_n108  &  wire1178 ) ;
 assign wire17186 = ( n_n108  &  wire827 ) | ( n_n101  &  wire826 ) ;
 assign wire17187 = ( n_n51  &  n_n101 ) | ( n_n53  &  n_n101 ) | ( n_n51  &  n_n108 ) ;
 assign wire17190 = ( wire4685 ) | ( n_n46  &  wire168 ) | ( n_n46  &  wire181 ) ;
 assign wire17191 = ( wire4684 ) | ( wire17187 ) | ( n_n47  &  wire181 ) ;
 assign wire17193 = ( n_n2253 ) | ( wire17185 ) | ( wire17186 ) ;
 assign wire17196 = ( n_n46  &  n_n61 ) | ( n_n47  &  n_n61 ) | ( n_n47  &  n_n63 ) ;
 assign wire17198 = ( n_n4007 ) | ( wire17196 ) | ( n_n47  &  wire888 ) ;
 assign wire17201 = ( n_n43  &  wire93 ) | ( n_n43  &  wire729  &  n_n191 ) ;
 assign wire17202 = ( n_n46  &  n_n156  &  wire725 ) | ( n_n47  &  n_n156  &  wire725 ) ;
 assign wire17203 = ( n_n46  &  n_n57 ) | ( n_n46  &  wire894 ) | ( n_n47  &  wire894 ) ;
 assign wire17206 = ( wire4669 ) | ( wire4676 ) | ( wire17201 ) | ( wire17202 ) ;
 assign wire17209 = ( n_n47  &  wire176 ) | ( n_n47  &  wire149 ) ;
 assign wire17212 = ( wire561 ) | ( wire4662 ) | ( wire4663 ) | ( wire17209 ) ;
 assign wire17213 = ( wire4671 ) | ( wire17203 ) | ( wire17206 ) | ( wire17212 ) ;
 assign wire17215 = ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire17217 = ( n_n135  &  n_n32 ) | ( n_n31  &  wire181 ) ;
 assign wire17220 = ( n_n32  &  n_n182 ) | ( n_n33  &  wire60 ) ;
 assign wire17224 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire17226 = ( n_n36  &  n_n156  &  wire725 ) | ( n_n36  &  n_n149  &  wire725 ) ;
 assign wire17228 = ( wire4649 ) | ( wire17226 ) | ( n_n34  &  wire1056 ) ;
 assign wire17229 = ( wire4651 ) | ( wire4655 ) | ( wire17220 ) ;
 assign wire17231 = ( n_n31  &  wire129 ) | ( n_n30  &  wire181 ) ;
 assign wire17234 = ( wire4644 ) | ( wire17228 ) | ( wire17229 ) | ( wire17231 ) ;
 assign wire17238 = ( wire176 ) | ( wire299 ) | ( wire418 ) ;
 assign wire17239 = ( n_n31  &  wire158 ) | ( n_n31  &  n_n216  &  wire725 ) ;
 assign wire17241 = ( wire4638 ) | ( wire17239 ) | ( wire213  &  n_n61 ) ;
 assign wire17243 = ( n_n31  &  wire1189 ) | ( n_n31  &  wire1188 ) | ( n_n30  &  wire1188 ) ;
 assign wire17245 = ( n_n31  &  wire149 ) | ( n_n30  &  wire131 ) ;
 assign wire17246 = ( wire17243 ) | ( wire17245 ) | ( n_n30  &  wire1190 ) ;
 assign wire17247 = ( wire4628 ) | ( n_n31  &  wire902 ) ;
 assign wire17249 = ( wire4639 ) | ( wire17241 ) | ( wire17246 ) | ( wire17247 ) ;
 assign wire17251 = ( n_n135  &  n_n125 ) | ( n_n135  &  n_n123 ) | ( n_n125  &  wire1177 ) ;
 assign wire17253 = ( (~ i_15_)  &  n_n149  &  n_n201 ) | ( i_15_  &  n_n149  &  n_n211 ) | ( (~ i_15_)  &  n_n149  &  n_n211 ) ;
 assign wire17256 = ( n_n71  &  n_n125 ) | ( n_n125  &  wire115 ) | ( n_n125  &  wire17253 ) ;
 assign wire17257 = ( wire17251 ) | ( n_n123  &  wire971 ) | ( n_n123  &  wire1176 ) ;
 assign wire17258 = ( n_n53  &  n_n123 ) | ( n_n125  &  n_n57 ) ;
 assign wire17259 = ( n_n125  &  wire1115 ) | ( n_n123  &  wire1114 ) ;
 assign wire17260 = ( wire255  &  n_n55 ) | ( n_n113  &  n_n182 ) ;
 assign wire17265 = ( n_n5739 ) | ( wire440 ) | ( n_n108  &  n_n210 ) ;
 assign wire17266 = ( n_n5743 ) | ( wire447 ) | ( n_n135  &  n_n113 ) ;
 assign wire17268 = ( wire17265 ) | ( wire17266 ) | ( n_n112  &  wire973 ) ;
 assign wire17271 = ( i_15_  &  n_n177  &  n_n211 ) | ( (~ i_15_)  &  n_n177  &  n_n211 ) | ( i_15_  &  n_n170  &  n_n211 ) | ( (~ i_15_)  &  n_n170  &  n_n211 ) ;
 assign wire17272 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire17275 = ( n_n123  &  n_n77 ) | ( n_n123  &  wire117 ) | ( n_n123  &  wire17271 ) ;
 assign wire17276 = ( wire4602 ) | ( n_n125  &  wire975 ) | ( n_n125  &  wire1234 ) ;
 assign wire17277 = ( wire17276 ) | ( wire17275 ) ;
 assign wire17280 = ( n_n53  &  n_n40 ) | ( n_n38  &  n_n168 ) ;
 assign wire17281 = ( n_n51  &  wire190 ) | ( wire334  &  n_n78 ) ;
 assign wire17284 = ( n_n53  &  n_n41 ) | ( n_n41  &  wire1117 ) | ( n_n40  &  wire1117 ) ;
 assign wire17285 = ( n_n135  &  n_n41 ) | ( n_n135  &  n_n40 ) | ( n_n41  &  n_n57 ) | ( n_n40  &  n_n57 ) ;
 assign wire17287 = ( wire724  &  n_n177 ) | ( n_n177  &  wire722 ) ;
 assign wire17288 = ( n_n39  &  wire1120 ) | ( n_n39  &  wire726  &  n_n156 ) ;
 assign wire17289 = ( wire4581 ) | ( wire17284 ) | ( wire17285 ) ;
 assign wire17290 = ( wire4591 ) | ( wire17280 ) | ( wire17281 ) | ( wire17288 ) ;
 assign wire17291 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire377 ) ;
 assign wire17292 = ( wire722  &  n_n149 ) | ( n_n216  &  wire725 ) ;
 assign wire17294 = ( n_n156  &  wire722 ) | ( n_n216  &  wire725 ) ;
 assign wire17295 = ( wire729  &  n_n156 ) | ( wire726  &  n_n156 ) | ( wire729  &  n_n149 ) | ( wire726  &  n_n149 ) ;
 assign wire17297 = ( wire4572 ) | ( wire190  &  n_n199  &  wire725 ) ;
 assign wire17298 = ( wire4573 ) | ( wire4576 ) | ( wire17291 ) ;
 assign wire17299 = ( n_n38  &  n_n150 ) | ( n_n36  &  n_n102 ) ;
 assign wire17301 = ( n_n36  &  wire978 ) | ( n_n34  &  n_n102 ) ;
 assign wire17303 = ( wire4568 ) | ( wire4569 ) | ( wire17299 ) | ( wire17301 ) ;
 assign wire17305 = ( wire17289 ) | ( wire17290 ) | ( wire17297 ) | ( wire17298 ) ;
 assign wire17307 = ( n_n34  &  n_n216  &  wire725 ) | ( n_n34  &  n_n191  &  wire725 ) ;
 assign wire17309 = ( (~ i_15_)  &  n_n149  &  n_n201 ) | ( i_15_  &  n_n149  &  n_n211 ) | ( (~ i_15_)  &  n_n149  &  n_n211 ) ;
 assign wire17310 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign wire17313 = ( wire116 ) | ( wire371 ) | ( n_n199  &  wire725 ) ;
 assign wire17314 = ( n_n36  &  n_n63 ) | ( n_n36  &  wire115 ) | ( n_n36  &  wire17309 ) ;
 assign wire17317 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire729 ) ;
 assign wire17319 = ( i_15_  &  n_n184  &  n_n211 ) | ( (~ i_15_)  &  n_n184  &  n_n211 ) | ( i_15_  &  n_n177  &  n_n211 ) | ( (~ i_15_)  &  n_n177  &  n_n211 ) ;
 assign wire17321 = ( wire4544 ) | ( n_n36  &  n_n184  &  wire729 ) ;
 assign wire17322 = ( wire4545 ) | ( wire4548 ) | ( wire4549 ) ;
 assign wire17324 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire17325 = ( wire614 ) | ( wire583 ) | ( wire4550 ) | ( wire4551 ) ;
 assign wire17327 = ( wire4539 ) | ( wire17325 ) | ( n_n34  &  wire980 ) ;
 assign wire17329 = ( n_n42  &  n_n89 ) | ( n_n41  &  n_n210 ) ;
 assign wire17333 = ( n_n41  &  n_n202 ) | ( n_n41  &  n_n102 ) | ( n_n41  &  wire70 ) ;
 assign wire17335 = ( wire4526 ) | ( n_n40  &  wire1052 ) ;
 assign wire17336 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) | ( n_n177  &  wire722 ) ;
 assign wire17337 = ( n_n41  &  wire69 ) | ( n_n41  &  n_n156  &  wire722 ) ;
 assign wire17338 = ( n_n40  &  n_n202 ) | ( n_n40  &  n_n102 ) | ( n_n40  &  wire263 ) ;
 assign wire17339 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire722 ) ;
 assign wire17341 = ( n_n41  &  wire51 ) | ( n_n41  &  wire202 ) | ( n_n41  &  wire17339 ) ;
 assign wire17342 = ( wire4520 ) | ( wire17338 ) | ( n_n40  &  wire1794 ) ;
 assign wire17343 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) ;
 assign wire17345 = ( wire397 ) | ( wire4523 ) | ( wire17337 ) ;
 assign wire17347 = ( wire4510 ) | ( wire17345 ) | ( n_n41  &  wire984 ) ;
 assign wire17349 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire17350 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) ;
 assign wire17352 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire722 ) ;
 assign wire17353 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) ;
 assign wire17357 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire722 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire722 ) ;
 assign wire17358 = ( wire4503 ) | ( wire4504 ) | ( n_n101  &  wire57 ) ;
 assign wire17359 = ( wire4500 ) | ( n_n101  &  wire1060 ) ;
 assign wire17360 = ( n_n101  &  wire86 ) | ( n_n101  &  wire263 ) ;
 assign wire17361 = ( n_n199  &  wire729 ) | ( n_n199  &  wire726 ) | ( n_n199  &  wire722 ) ;
 assign wire17363 = ( wire4491 ) | ( wire4496 ) | ( wire17360 ) ;
 assign wire17364 = ( wire17363 ) | ( n_n108  &  wire1064 ) ;
 assign wire17365 = ( n_n2257 ) | ( wire17358 ) | ( wire17359 ) ;
 assign wire17367 = ( n_n212  &  wire176 ) | ( n_n197  &  wire149 ) ;
 assign wire17368 = ( n_n212  &  wire149 ) | ( n_n197  &  wire131 ) ;
 assign wire17374 = ( n_n197  &  wire129 ) | ( n_n212  &  wire130 ) ;
 assign wire17377 = ( n_n212  &  wire168 ) | ( n_n197  &  wire181 ) | ( n_n212  &  wire181 ) ;
 assign wire17379 = ( wire4474 ) | ( wire4475 ) | ( wire17377 ) ;
 assign wire17382 = ( n_n51  &  n_n197 ) | ( n_n53  &  n_n197 ) | ( n_n51  &  n_n212 ) | ( n_n53  &  n_n212 ) ;
 assign wire17383 = ( n_n197  &  wire176 ) | ( n_n212  &  n_n63 ) ;
 assign wire17384 = ( n_n197  &  n_n61 ) | ( n_n212  &  n_n61 ) | ( n_n197  &  wire308 ) ;
 assign wire17385 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire725 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire725 ) ;
 assign wire17388 = ( n_n197  &  n_n55 ) | ( n_n212  &  n_n55 ) | ( n_n197  &  wire887 ) ;
 assign wire17389 = ( wire4460 ) | ( n_n197  &  wire158 ) | ( n_n212  &  wire158 ) ;
 assign wire17390 = ( wire17383 ) | ( wire17384 ) | ( wire17388 ) ;
 assign wire17391 = ( (~ i_15_)  &  n_n191  &  n_n201 ) | ( i_15_  &  n_n191  &  n_n211 ) | ( (~ i_15_)  &  n_n191  &  n_n211 ) ;
 assign wire17392 = ( n_n125  &  n_n117 ) | ( n_n123  &  n_n102 ) ;
 assign wire17393 = ( wire4458 ) | ( wire4459 ) | ( wire17392 ) ;
 assign wire17394 = ( wire4454 ) | ( wire4453 ) ;
 assign wire17395 = ( (~ i_15_)  &  n_n199  &  n_n201 ) | ( i_15_  &  n_n199  &  n_n211 ) | ( (~ i_15_)  &  n_n199  &  n_n211 ) ;
 assign wire17397 = ( n_n125  &  n_n102 ) | ( n_n125  &  wire243 ) | ( n_n125  &  wire17395 ) ;
 assign wire17398 = ( wire4470 ) | ( wire17382 ) | ( n_n123  &  wire1124 ) ;
 assign wire17400 = ( wire17389 ) | ( wire17390 ) | ( wire17393 ) | ( wire17394 ) ;
 assign wire17401 = ( n_n5144 ) | ( wire17190 ) | ( wire17191 ) | ( wire17193 ) ;
 assign wire17405 = ( n_n2234 ) | ( wire17397 ) | ( wire17398 ) | ( wire17400 ) ;
 assign wire17407 = ( n_n2229 ) | ( n_n2232 ) | ( n_n2227 ) | ( n_n2226 ) ;
 assign wire17408 = ( n_n2228 ) | ( wire17364 ) | ( wire17365 ) | ( wire17405 ) ;
 assign wire17410 = ( n_n30  &  wire55 ) | ( n_n30  &  wire181 ) ;
 assign wire17416 = ( wire152 ) | ( wire220 ) | ( wire720  &  n_n149 ) ;
 assign wire17417 = ( n_n33  &  wire60 ) | ( n_n33  &  n_n149  &  wire719 ) ;
 assign wire17418 = ( n_n31  &  wire143 ) | ( n_n34  &  wire122 ) ;
 assign wire17420 = ( wire443 ) | ( wire17417 ) | ( wire17418 ) ;
 assign wire17426 = ( wire134 ) | ( wire158 ) | ( wire127 ) ;
 assign wire17428 = ( n_n156  &  wire721 ) | ( n_n216  &  wire725 ) | ( n_n156  &  wire725 ) ;
 assign wire17431 = ( wire654 ) | ( n_n31  &  wire125 ) ;
 assign wire17433 = ( wire4419 ) | ( wire4427 ) | ( n_n30  &  wire144 ) ;
 assign wire17434 = ( n_n4240 ) | ( n_n4154 ) | ( wire4420 ) | ( wire17431 ) ;
 assign wire17435 = ( n_n4247 ) | ( wire4429 ) | ( wire4430 ) | ( wire17433 ) ;
 assign wire17436 = ( n_n34  &  wire133 ) | ( n_n34  &  wire181 ) ;
 assign wire17438 = ( wire541 ) | ( n_n34  &  wire55 ) | ( n_n34  &  wire158 ) ;
 assign wire17439 = ( wire458 ) | ( wire17436 ) | ( n_n34  &  wire127 ) ;
 assign wire17440 = ( n_n34  &  wire134 ) | ( n_n34  &  wire123 ) ;
 assign wire17441 = ( n_n34  &  wire176 ) | ( n_n34  &  wire156 ) ;
 assign wire17443 = ( n_n36  &  wire55 ) | ( n_n36  &  wire127 ) ;
 assign wire17445 = ( wire17441 ) | ( n_n36  &  wire133 ) | ( n_n36  &  wire125 ) ;
 assign wire17446 = ( wire17440 ) | ( wire17443 ) | ( n_n36  &  wire158 ) ;
 assign wire17447 = ( n_n156  &  wire719 ) | ( n_n149  &  wire719 ) | ( n_n156  &  wire728 ) ;
 assign wire17448 = ( n_n156  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n149  &  wire725 ) ;
 assign wire17450 = ( n_n34  &  wire125 ) | ( n_n34  &  n_n216  &  wire725 ) ;
 assign wire17452 = ( n_n4564 ) | ( wire709 ) | ( wire4396 ) | ( wire4986 ) ;
 assign wire17453 = ( wire4395 ) | ( wire17450 ) | ( wire17452 ) ;
 assign wire17454 = ( wire17438 ) | ( wire17439 ) | ( wire17445 ) | ( wire17446 ) ;
 assign wire17456 = ( wire4768 ) | ( wire17122 ) | ( wire157  &  n_n125 ) ;
 assign wire17457 = ( wire601 ) | ( wire4393 ) | ( wire4750 ) | ( wire4751 ) ;
 assign wire17458 = ( n_n123  &  wire86 ) | ( n_n123  &  wire720  &  n_n149 ) ;
 assign wire17459 = ( n_n125  &  wire155 ) | ( n_n123  &  wire180 ) ;
 assign wire17462 = ( wire570 ) | ( wire4765 ) | ( wire17123 ) | ( wire17458 ) ;
 assign wire17465 = ( n_n1700 ) | ( n_n125  &  wire803 ) ;
 assign wire17466 = ( wire4376 ) | ( wire4382 ) | ( wire17459 ) | ( wire17462 ) ;
 assign wire17467 = ( wire17456 ) | ( wire17457 ) | ( wire17465 ) ;
 assign wire17468 = ( n_n149  &  wire719 ) | ( n_n156  &  wire725 ) ;
 assign wire17469 = ( n_n101  &  wire90 ) | ( n_n108  &  n_n142 ) ;
 assign wire17470 = ( n_n53  &  n_n108 ) | ( n_n101  &  wire218 ) ;
 assign wire17471 = ( wire157  &  n_n108 ) | ( n_n101  &  wire141 ) ;
 assign wire17472 = ( wire4372 ) | ( wire4838 ) | ( wire4839 ) | ( wire17469 ) ;
 assign wire17478 = ( wire511 ) | ( n_n108  &  wire84 ) | ( n_n108  &  wire220 ) ;
 assign wire17479 = ( n_n4996 ) | ( n_n4994 ) | ( n_n101  &  wire946 ) ;
 assign wire17480 = ( n_n149  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n149  &  wire725 ) ;
 assign wire17483 = ( wire4343 ) | ( n_n47  &  wire85 ) ;
 assign wire17484 = ( n_n6005 ) | ( wire419 ) | ( n_n1624 ) | ( wire4344 ) ;
 assign wire17486 = ( wire4829 ) | ( wire4830 ) | ( wire17483 ) | ( wire17484 ) ;
 assign wire17490 = ( wire729  &  n_n156 ) | ( wire726  &  n_n156 ) | ( wire720  &  n_n156 ) ;
 assign wire17493 = ( n_n46  &  wire799 ) | ( n_n46  &  wire142 ) | ( n_n46  &  wire180 ) ;
 assign wire17498 = ( wire155 ) | ( wire60 ) | ( wire220 ) ;
 assign wire17499 = ( n_n1594 ) | ( n_n47  &  wire808 ) ;
 assign wire17501 = ( wire4334 ) | ( wire4341 ) | ( wire17493 ) | ( wire17499 ) ;
 assign wire17504 = ( n_n5000 ) | ( n_n101  &  wire86 ) | ( n_n101  &  wire84 ) ;
 assign wire17505 = ( n_n4900 ) | ( n_n108  &  wire867 ) ;
 assign wire17507 = ( n_n5739 ) | ( wire4950 ) | ( n_n53  &  n_n123 ) ;
 assign wire17509 = ( n_n5037 ) | ( wire17507 ) | ( wire157  &  n_n123 ) ;
 assign wire17510 = ( n_n4904 ) | ( wire4323 ) | ( wire4324 ) ;
 assign wire17513 = ( n_n4903 ) | ( wire17504 ) | ( wire17505 ) | ( wire17509 ) ;
 assign wire17514 = ( wire544 ) | ( wire17510 ) | ( wire17513 ) ;
 assign wire17516 = ( n_n212  &  wire55 ) | ( n_n197  &  wire181 ) ;
 assign wire17518 = ( n_n212  &  wire123 ) | ( n_n197  &  wire127 ) ;
 assign wire17521 = ( wire17518 ) | ( n_n197  &  wire158 ) | ( n_n197  &  wire133 ) ;
 assign wire17522 = ( wire532 ) | ( wire594 ) | ( wire660 ) | ( wire17516 ) ;
 assign wire17528 = ( wire361 ) | ( wire363 ) | ( n_n40  &  wire180 ) ;
 assign wire17529 = ( wire426 ) | ( n_n41  &  wire155 ) | ( n_n41  &  wire205 ) ;
 assign wire17533 = ( wire4291 ) | ( n_n41  &  wire60 ) | ( n_n41  &  wire220 ) ;
 assign wire17534 = ( n_n3979 ) | ( n_n1542 ) | ( wire645 ) | ( wire664 ) ;
 assign wire17535 = ( n_n149  &  wire719 ) | ( n_n156  &  wire725 ) ;
 assign wire17537 = ( wire4285 ) | ( wire4908 ) | ( wire17016 ) ;
 assign wire17539 = ( wire4286 ) | ( wire4904 ) | ( wire4905 ) | ( wire17537 ) ;
 assign wire17541 = ( n_n38  &  wire726  &  n_n156 ) | ( n_n38  &  n_n156  &  wire728 ) ;
 assign wire17542 = ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) | ( n_n39  &  n_n52 ) ;
 assign wire17543 = ( n_n1514 ) | ( wire17541 ) | ( wire17542 ) ;
 assign wire17545 = ( n_n38  &  wire248 ) | ( n_n39  &  wire248 ) ;
 assign wire17548 = ( n_n1520 ) | ( wire571 ) | ( n_n39  &  wire110 ) ;
 assign wire17549 = ( n_n1517 ) | ( wire17545 ) | ( n_n39  &  wire249 ) ;
 assign wire17550 = ( wire457 ) | ( wire4263 ) | ( wire4888 ) | ( wire17028 ) ;
 assign wire17552 = ( n_n4460 ) | ( wire17033 ) | ( wire17550 ) ;
 assign wire17553 = ( wire597 ) | ( wire17543 ) | ( wire17548 ) | ( wire17549 ) ;
 assign wire17554 = ( n_n47  &  n_n128 ) | ( n_n47  &  n_n156  &  wire725 ) ;
 assign wire17555 = ( n_n46  &  wire90 ) | ( n_n47  &  n_n142 ) ;
 assign wire17557 = ( wire652 ) | ( wire4260 ) | ( wire17554 ) ;
 assign wire17558 = ( n_n4312 ) | ( wire4859 ) | ( wire4860 ) | ( wire17555 ) ;
 assign wire17559 = ( wire4252 ) | ( wire4253 ) | ( n_n53  &  n_n46 ) ;
 assign wire17560 = ( n_n6267 ) | ( n_n6269 ) | ( wire157  &  n_n46 ) ;
 assign wire17562 = ( wire17559 ) | ( wire17560 ) | ( n_n47  &  wire152 ) ;
 assign wire17563 = ( wire549 ) | ( wire4919 ) | ( wire17003 ) ;
 assign wire17565 = ( wire621 ) | ( wire17557 ) | ( wire17558 ) ;
 assign wire17566 = ( wire17562 ) | ( wire17563 ) | ( wire17565 ) ;
 assign wire17568 = ( n_n125  &  n_n214 ) | ( n_n197  &  wire122 ) ;
 assign wire17569 = ( n_n156  &  wire719 ) | ( n_n149  &  wire719 ) | ( n_n156  &  wire728 ) ;
 assign wire17570 = ( n_n156  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n149  &  wire725 ) ;
 assign wire17573 = ( wire4233 ) | ( n_n197  &  n_n63 ) | ( n_n197  &  wire125 ) ;
 assign wire17574 = ( wire422 ) | ( wire4234 ) | ( wire17568 ) ;
 assign wire17575 = ( n_n197  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign wire17576 = ( wire565 ) | ( n_n212  &  wire158 ) ;
 assign wire17578 = ( n_n4231 ) | ( wire4230 ) | ( wire17575 ) | ( wire17576 ) ;
 assign wire17579 = ( wire17114 ) | ( wire17115 ) | ( wire17573 ) | ( wire17574 ) ;
 assign wire17581 = ( n_n4116 ) | ( wire17578 ) | ( wire17579 ) ;
 assign wire17582 = ( wire17466 ) | ( wire17467 ) | ( wire17581 ) ;
 assign wire17585 = ( wire17434 ) | ( wire17435 ) | ( wire17453 ) | ( wire17454 ) ;
 assign wire17586 = ( n_n5144 ) | ( n_n4106 ) | ( wire17585 ) ;
 assign wire17587 = ( i_7_  &  (~ i_5_)  &  i_6_ ) ;
 assign wire17588 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire17591 = ( (~ i_7_)  &  (~ i_5_)  &  i_6_ ) | ( i_7_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire17592 = ( wire4220 ) | ( wire170  &  wire1527 ) ;
 assign wire17593 = ( n_n9  &  n_n144 ) | ( n_n6  &  n_n144 ) | ( n_n5  &  n_n144 ) ;
 assign wire17594 = ( n_n162  &  n_n157  &  n_n219 ) | ( n_n157  &  n_n48  &  n_n219 ) ;
 assign wire17596 = ( n_n16  &  n_n48  &  n_n219 ) | ( n_n16  &  n_n219  &  n_n218 ) ;
 assign wire17599 = ( wire569 ) | ( wire17594 ) | ( n_n14  &  wire170 ) ;
 assign wire17600 = ( n_n7267 ) | ( wire684 ) | ( n_n2956 ) | ( wire17596 ) ;
 assign wire17601 = ( wire4228 ) | ( wire4229 ) | ( wire17599 ) ;
 assign wire17602 = ( wire4217 ) | ( wire4221 ) | ( wire17592 ) | ( wire17593 ) ;
 assign wire17604 = ( n_n71  &  n_n4 ) | ( n_n13  &  wire1496 ) ;
 assign wire17605 = ( n_n5144 ) | ( n_n19  &  n_n157  &  n_n111 ) ;
 assign wire17606 = ( i_7_  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire17608 = ( wire569 ) | ( n_n13  &  n_n149  &  wire725 ) ;
 assign wire17610 = ( wire529 ) | ( wire568 ) | ( n_n4  &  wire77 ) ;
 assign wire17612 = ( wire17605 ) | ( wire17606 ) | ( wire17608 ) | ( wire17610 ) ;
 assign wire17615 = ( wire176 ) | ( wire156 ) | ( wire212 ) ;
 assign wire17622 = ( wire445 ) | ( n_n53  &  n_n108 ) | ( wire157  &  n_n108 ) ;
 assign wire17626 = ( wire4172 ) | ( n_n4981 ) ;
 assign wire17627 = ( wire17622 ) | ( n_n101  &  wire1321 ) | ( n_n101  &  wire1488 ) ;
 assign wire17629 = ( n_n3570 ) | ( n_n3823 ) | ( wire4185 ) | ( wire4186 ) ;
 assign wire17631 = ( n_n46  &  n_n134 ) | ( n_n47  &  wire78 ) ;
 assign wire17632 = ( n_n156  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n156  &  wire725 ) ;
 assign wire17635 = ( n_n6266 ) | ( n_n47  &  n_n156  &  wire725 ) ;
 assign wire17638 = ( wire4159 ) | ( wire172  &  n_n47 ) | ( n_n47  &  wire80 ) ;
 assign wire17639 = ( n_n6271 ) | ( n_n6267 ) | ( wire17635 ) | ( wire17638 ) ;
 assign wire17640 = ( wire651 ) | ( wire4158 ) | ( wire17631 ) ;
 assign wire17646 = ( n_n1553 ) | ( wire500 ) | ( wire361 ) | ( wire4151 ) ;
 assign wire17647 = ( wire497 ) | ( n_n40  &  wire1450 ) ;
 assign wire17650 = ( n_n3542 ) | ( n_n41  &  n_n155 ) | ( n_n41  &  wire215 ) ;
 assign wire17651 = ( wire397 ) | ( wire653 ) | ( wire4143 ) ;
 assign wire17654 = ( n_n40  &  wire180 ) | ( n_n41  &  n_n214 ) | ( n_n40  &  n_n214 ) ;
 assign wire17656 = ( wire359 ) | ( wire537 ) | ( n_n59  &  n_n43 ) ;
 assign wire17657 = ( wire17654 ) | ( n_n41  &  wire142 ) | ( n_n41  &  wire180 ) ;
 assign wire17659 = ( n_n4623 ) | ( wire4130 ) | ( wire17656 ) | ( wire17657 ) ;
 assign wire17660 = ( wire17646 ) | ( wire17647 ) | ( wire17650 ) | ( wire17651 ) ;
 assign wire17662 = ( n_n41  &  wire182 ) | ( n_n41  &  n_n130 ) | ( n_n41  &  n_n57 ) ;
 assign wire17663 = ( n_n38  &  wire104 ) | ( n_n38  &  wire279 ) ;
 assign wire17667 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n134 ) | ( n_n38  &  wire110 ) ;
 assign wire17668 = ( n_n38  &  n_n150 ) | ( n_n39  &  n_n150 ) | ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) ;
 assign wire17671 = ( wire17668 ) | ( n_n38  &  wire248 ) | ( n_n39  &  wire248 ) ;
 assign wire17672 = ( wire605 ) | ( n_n972 ) | ( wire17663 ) | ( wire17667 ) ;
 assign wire17674 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire141 ) ;
 assign wire17676 = ( wire17674 ) | ( n_n40  &  wire155 ) | ( n_n40  &  wire205 ) ;
 assign wire17677 = ( n_n3979 ) | ( wire442 ) | ( wire4113 ) ;
 assign wire17679 = ( n_n40  &  n_n63 ) | ( n_n40  &  n_n191  &  wire719 ) ;
 assign wire17681 = ( wire503 ) | ( wire17679 ) | ( wire172  &  n_n40 ) ;
 assign wire17682 = ( wire4104 ) | ( n_n53  &  n_n40 ) | ( wire157  &  n_n40 ) ;
 assign wire17684 = ( wire4126 ) | ( wire17662 ) | ( wire17681 ) | ( wire17682 ) ;
 assign wire17685 = ( wire17671 ) | ( wire17672 ) | ( wire17676 ) | ( wire17677 ) ;
 assign wire17686 = ( n_n47  &  n_n63 ) | ( n_n46  &  wire212 ) ;
 assign wire17688 = ( n_n46  &  wire134 ) | ( n_n47  &  wire125 ) ;
 assign wire17690 = ( n_n5107 ) | ( wire688 ) | ( n_n46  &  wire176 ) ;
 assign wire17691 = ( wire560 ) | ( wire17686 ) | ( wire17688 ) ;
 assign wire17692 = ( wire52  &  n_n43 ) | ( wire129  &  n_n43 ) ;
 assign wire17693 = ( n_n42  &  wire63 ) | ( n_n43  &  wire63 ) | ( n_n42  &  wire48 ) | ( n_n43  &  wire48 ) ;
 assign wire17695 = ( wire4102 ) | ( wire4103 ) | ( wire17692 ) | ( wire17693 ) ;
 assign wire17696 = ( wire17639 ) | ( wire17640 ) | ( wire17690 ) | ( wire17691 ) ;
 assign wire17697 = ( wire17696 ) | ( wire17695 ) ;
 assign wire17698 = ( wire17659 ) | ( wire17660 ) | ( wire17684 ) | ( wire17685 ) ;
 assign wire17700 = ( wire419 ) | ( n_n200  &  wire1375 ) ;
 assign wire17701 = ( n_n46  &  wire181 ) | ( n_n46  &  wire47 ) ;
 assign wire17704 = ( wire481 ) | ( wire17700 ) | ( wire17701 ) ;
 assign wire17705 = ( n_n47  &  wire129 ) | ( n_n46  &  wire131 ) ;
 assign wire17706 = ( wire137  &  n_n46 ) | ( n_n46  &  wire146 ) | ( n_n46  &  wire46 ) ;
 assign wire17708 = ( wire4088 ) | ( wire17705 ) | ( n_n47  &  wire46 ) ;
 assign wire17709 = ( n_n3561 ) | ( n_n3889 ) ;
 assign wire17710 = ( wire674 ) | ( wire671 ) | ( wire17706 ) ;
 assign wire17712 = ( wire577 ) | ( wire4080 ) | ( wire17704 ) | ( wire17710 ) ;
 assign wire17716 = ( n_n5739 ) | ( wire440 ) | ( n_n112  &  wire160 ) ;
 assign wire17717 = ( n_n5743 ) | ( wire447 ) | ( n_n108  &  wire47 ) ;
 assign wire17721 = ( wire729  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire715 ) ;
 assign wire17724 = ( wire93 ) | ( wire171 ) | ( wire17721 ) ;
 assign wire17725 = ( wire157  &  n_n123 ) | ( n_n123  &  n_n156  &  wire725 ) ;
 assign wire17726 = ( wire515 ) | ( wire4064 ) | ( wire4065 ) | ( wire17725 ) ;
 assign wire17729 = ( n_n101  &  wire181 ) | ( n_n101  &  wire1378 ) | ( n_n108  &  wire1378 ) ;
 assign wire17732 = ( n_n125  &  wire141 ) | ( n_n125  &  wire160 ) ;
 assign wire17735 = ( n_n2859 ) | ( n_n4657 ) | ( wire4048 ) | ( wire17732 ) ;
 assign wire17739 = ( n_n155 ) | ( wire224 ) | ( wire250 ) | ( wire57 ) ;
 assign wire17740 = ( wire479 ) | ( wire90  &  n_n125 ) | ( n_n125  &  wire205 ) ;
 assign wire17741 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire17744 = ( n_n125  &  n_n176 ) | ( n_n125  &  wire51 ) | ( n_n123  &  wire51 ) ;
 assign wire17746 = ( wire394 ) | ( n_n123  &  wire1420 ) ;
 assign wire17747 = ( wire17744 ) | ( wire17746 ) | ( n_n125  &  wire100 ) ;
 assign wire17748 = ( n_n3912 ) | ( wire4043 ) | ( wire17735 ) | ( wire17740 ) ;
 assign wire17750 = ( n_n53  &  n_n212 ) | ( n_n197  &  n_n134 ) ;
 assign wire17752 = ( wire4027 ) | ( wire689 ) ;
 assign wire17753 = ( wire422 ) | ( wire4026 ) | ( wire17568 ) | ( wire17750 ) ;
 assign wire17756 = ( wire4020 ) | ( n_n212  &  wire176 ) | ( n_n212  &  n_n63 ) ;
 assign wire17757 = ( wire565 ) | ( wire4021 ) | ( wire4230 ) | ( wire17575 ) ;
 assign wire17760 = ( n_n123  &  wire180 ) | ( n_n123  &  wire86 ) ;
 assign wire17761 = ( n_n123  &  wire85 ) | ( n_n123  &  wire142 ) | ( n_n123  &  n_n214 ) ;
 assign wire17764 = ( n_n3592 ) | ( wire4013 ) | ( wire17760 ) | ( wire17761 ) ;
 assign wire17765 = ( wire17752 ) | ( wire17753 ) | ( wire17756 ) | ( wire17757 ) ;
 assign wire17766 = ( n_n197  &  wire52 ) | ( n_n197  &  wire129 ) ;
 assign wire17767 = ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) | ( n_n212  &  wire63 ) ;
 assign wire17772 = ( n_n197  &  wire181 ) | ( n_n212  &  wire48 ) ;
 assign wire17773 = ( n_n212  &  wire181 ) | ( n_n197  &  wire47 ) ;
 assign wire17776 = ( n_n4518 ) | ( wire3998 ) | ( wire17772 ) | ( wire17773 ) ;
 assign wire17778 = ( n_n3834 ) | ( n_n3833 ) | ( wire17776 ) ;
 assign wire17779 = ( wire17747 ) | ( wire17748 ) | ( wire17764 ) | ( wire17765 ) ;
 assign wire17781 = ( n_n177  &  wire719 ) | ( n_n191  &  wire725 ) ;
 assign wire17783 = ( n_n31  &  wire125 ) | ( n_n31  &  n_n216  &  wire725 ) ;
 assign wire17786 = ( n_n4915 ) | ( wire3991 ) | ( wire3996 ) | ( wire3997 ) ;
 assign wire17787 = ( n_n30  &  wire176 ) | ( n_n30  &  wire123 ) | ( n_n30  &  wire131 ) ;
 assign wire17793 = ( n_n31  &  wire129 ) | ( n_n30  &  wire181 ) ;
 assign wire17796 = ( n_n30  &  wire137 ) | ( n_n31  &  wire46 ) | ( n_n30  &  wire46 ) ;
 assign wire17798 = ( n_n3511 ) | ( wire3973 ) | ( wire17796 ) ;
 assign wire17800 = ( n_n36  &  n_n63 ) | ( n_n36  &  n_n191  &  wire719 ) ;
 assign wire17801 = ( n_n34  &  wire134 ) | ( n_n34  &  wire123 ) ;
 assign wire17805 = ( wire17801 ) | ( n_n34  &  wire176 ) | ( n_n34  &  wire156 ) ;
 assign wire17806 = ( wire541 ) | ( n_n4566 ) | ( wire3964 ) | ( wire17800 ) ;
 assign wire17808 = ( n_n156  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n156  &  wire725 ) ;
 assign wire17810 = ( n_n53  &  n_n36 ) | ( n_n34  &  n_n134 ) ;
 assign wire17812 = ( wire3957 ) | ( n_n33  &  n_n190 ) | ( n_n33  &  wire187 ) ;
 assign wire17813 = ( wire636 ) | ( wire3958 ) | ( wire17810 ) ;
 assign wire17816 = ( n_n33  &  n_n138 ) | ( n_n31  &  wire143 ) ;
 assign wire17817 = ( n_n31  &  wire181 ) | ( n_n30  &  wire47 ) ;
 assign wire17818 = ( wire17816 ) | ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) ;
 assign wire17819 = ( wire17817 ) | ( n_n33  &  wire1519 ) ;
 assign wire17821 = ( wire17805 ) | ( wire17806 ) | ( wire17812 ) | ( wire17813 ) ;
 assign wire17822 = ( n_n34  &  wire52 ) | ( n_n36  &  wire46 ) ;
 assign wire17824 = ( n_n38  &  n_n134 ) | ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) ;
 assign wire17825 = ( n_n34  &  wire143 ) | ( n_n34  &  wire181 ) ;
 assign wire17826 = ( n_n36  &  wire143 ) | ( n_n34  &  wire154 ) ;
 assign wire17827 = ( n_n36  &  wire181 ) | ( n_n34  &  wire47 ) ;
 assign wire17830 = ( wire432 ) | ( wire17824 ) | ( wire17827 ) ;
 assign wire17831 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17832 = ( n_n34  &  wire146 ) | ( n_n34  &  wire131 ) ;
 assign wire17836 = ( n_n3525 ) | ( wire17822 ) | ( n_n34  &  wire129 ) ;
 assign wire17837 = ( wire458 ) | ( wire640 ) | ( wire642 ) | ( wire606 ) ;
 assign wire17839 = ( wire17825 ) | ( wire17826 ) | ( wire17830 ) | ( wire17837 ) ;
 assign wire17840 = ( n_n5144 ) | ( wire213  &  n_n156  &  wire725 ) ;
 assign wire17841 = ( wire17840 ) | ( n_n30  &  wire157 ) ;
 assign wire17842 = ( wire3990 ) | ( wire17783 ) | ( wire17786 ) | ( wire17841 ) ;
 assign wire17843 = ( wire17626 ) | ( wire17627 ) | ( wire17629 ) | ( wire17842 ) ;
 assign wire17844 = ( n_n3795 ) | ( wire17708 ) | ( wire17709 ) | ( wire17712 ) ;
 assign wire17845 = ( n_n3787 ) | ( wire17818 ) | ( wire17819 ) | ( wire17821 ) ;
 assign wire17848 = ( wire17697 ) | ( wire17698 ) | ( wire17778 ) | ( wire17779 ) ;
 assign wire17849 = ( n_n3789 ) | ( wire17843 ) | ( wire17844 ) | ( wire17845 ) ;
 assign wire17850 = ( n_n162  &  n_n17  &  n_n219 ) | ( n_n17  &  n_n219  &  n_n218 ) ;
 assign wire17852 = ( wire17850 ) | ( wire463 ) ;
 assign wire17853 = ( wire568 ) | ( n_n7264 ) | ( n_n14  &  wire145 ) ;
 assign wire17854 = ( wire3899 ) | ( wire145  &  wire1044 ) ;
 assign wire17858 = ( n_n7252 ) | ( n_n7242 ) | ( wire3887 ) ;
 assign wire17860 = ( wire462 ) | ( wire3885 ) | ( wire3886 ) | ( wire17858 ) ;
 assign wire17861 = ( wire3900 ) | ( wire3901 ) | ( wire17852 ) | ( wire17853 ) ;
 assign wire17862 = ( wire3895 ) | ( wire3896 ) | ( wire3897 ) | ( wire17854 ) ;
 assign wire17864 = ( n_n36  &  wire123 ) | ( n_n34  &  wire127 ) ;
 assign wire17865 = ( wire137  &  n_n34 ) | ( n_n36  &  wire176 ) ;
 assign wire17867 = ( wire17864 ) | ( n_n34  &  wire146 ) | ( n_n34  &  wire131 ) ;
 assign wire17868 = ( wire458 ) | ( wire17865 ) | ( n_n34  &  wire55 ) ;
 assign wire17869 = ( wire640 ) | ( n_n36  &  wire130 ) ;
 assign wire17870 = ( n_n3525 ) | ( wire17822 ) | ( n_n34  &  wire129 ) ;
 assign wire17872 = ( n_n36  &  wire147 ) | ( n_n34  &  wire147 ) ;
 assign wire17873 = ( n_n36  &  wire149 ) | ( n_n34  &  wire126 ) ;
 assign wire17876 = ( wire584 ) | ( wire3866 ) | ( wire17872 ) | ( wire17873 ) ;
 assign wire17877 = ( wire17867 ) | ( wire17868 ) | ( wire17869 ) | ( wire17870 ) ;
 assign wire17880 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17881 = ( n_n36  &  wire139 ) | ( n_n36  &  wire124 ) | ( n_n36  &  wire128 ) ;
 assign wire17884 = ( n_n4581 ) | ( wire642 ) | ( wire4888 ) | ( wire17028 ) ;
 assign wire17887 = ( n_n34  &  n_n134 ) | ( n_n36  &  wire186 ) ;
 assign wire17889 = ( n_n34  &  wire176 ) | ( n_n34  &  n_n216  &  wire725 ) ;
 assign wire17891 = ( n_n36  &  wire125 ) | ( n_n34  &  wire125 ) ;
 assign wire17893 = ( n_n4564 ) | ( wire709 ) | ( wire17889 ) ;
 assign wire17894 = ( wire3850 ) | ( wire3851 ) | ( wire17891 ) ;
 assign wire17896 = ( n_n34  &  wire134 ) | ( n_n34  &  wire133 ) ;
 assign wire17897 = ( n_n34  &  wire123 ) | ( n_n34  &  wire156 ) ;
 assign wire17898 = ( n_n36  &  wire55 ) | ( n_n34  &  wire158 ) ;
 assign wire17901 = ( n_n191  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n170  &  wire725 ) ;
 assign wire17903 = ( n_n177  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire17906 = ( wire636 ) | ( wire3835 ) | ( wire17887 ) ;
 assign wire17908 = ( n_n2626 ) | ( wire17893 ) | ( wire17894 ) ;
 assign wire17909 = ( n_n149  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n149  &  wire725 ) ;
 assign wire17911 = ( n_n5144 ) | ( n_n36  &  n_n156  &  wire725 ) ;
 assign wire17913 = ( wire3828 ) | ( wire3829 ) | ( wire17911 ) ;
 assign wire17915 = ( n_n2622 ) | ( wire3836 ) | ( wire17906 ) | ( wire17908 ) ;
 assign wire17916 = ( n_n149  &  wire719 ) | ( n_n156  &  wire725 ) ;
 assign wire17918 = ( wire150 ) | ( wire152 ) ;
 assign wire17919 = ( wire153 ) | ( wire217 ) | ( n_n191  &  wire719 ) ;
 assign wire17920 = ( n_n135 ) | ( n_n132 ) | ( wire80 ) | ( wire78 ) ;
 assign wire17921 = ( wire157 ) | ( n_n63 ) | ( wire135 ) | ( wire17916 ) ;
 assign wire17924 = ( n_n31  &  wire172 ) | ( n_n31  &  wire125 ) ;
 assign wire17926 = ( n_n31  &  wire149 ) | ( n_n31  &  wire158 ) ;
 assign wire17931 = ( n_n31  &  wire129 ) | ( n_n31  &  wire46 ) ;
 assign wire17934 = ( n_n3510 ) | ( n_n31  &  wire1625 ) ;
 assign wire17935 = ( n_n4449 ) | ( n_n3514 ) | ( n_n3511 ) | ( wire17931 ) ;
 assign wire17940 = ( wire78 ) | ( wire217 ) | ( n_n170  &  wire719 ) ;
 assign wire17941 = ( n_n53 ) | ( n_n135 ) | ( wire80 ) | ( wire204 ) ;
 assign wire17942 = ( wire157 ) | ( wire172 ) | ( wire150 ) | ( wire173 ) ;
 assign wire17944 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire719 ) ;
 assign wire17947 = ( n_n31  &  wire143 ) | ( n_n31  &  wire181 ) ;
 assign wire17948 = ( n_n31  &  wire151 ) | ( n_n31  &  wire154 ) | ( n_n31  &  wire47 ) ;
 assign wire17951 = ( n_n36  &  wire176 ) | ( n_n36  &  wire123 ) | ( n_n36  &  wire1649 ) ;
 assign wire17952 = ( n_n2642 ) | ( n_n36  &  wire55 ) | ( n_n36  &  wire125 ) ;
 assign wire17954 = ( n_n3470 ) | ( wire3810 ) | ( wire3811 ) ;
 assign wire17955 = ( n_n39  &  n_n54 ) | ( n_n39  &  n_n52 ) | ( n_n39  &  n_n132 ) ;
 assign wire17958 = ( wire432 ) | ( n_n36  &  wire143 ) | ( n_n36  &  wire181 ) ;
 assign wire17959 = ( n_n4460 ) | ( wire17955 ) | ( n_n36  &  wire151 ) ;
 assign wire17960 = ( n_n36  &  wire149 ) | ( n_n36  &  wire147 ) ;
 assign wire17963 = ( n_n36  &  wire52 ) | ( n_n36  &  wire129 ) ;
 assign wire17964 = ( n_n36  &  wire139 ) | ( n_n36  &  wire46 ) ;
 assign wire17965 = ( n_n36  &  wire130 ) | ( n_n36  &  wire124 ) | ( n_n36  &  wire128 ) ;
 assign wire17968 = ( wire642 ) | ( wire17963 ) | ( wire17964 ) | ( wire17965 ) ;
 assign wire17970 = ( wire150 ) | ( n_n149  &  wire721 ) | ( n_n149  &  wire725 ) ;
 assign wire17971 = ( wire78 ) | ( wire217 ) | ( n_n170  &  wire719 ) ;
 assign wire17972 = ( n_n53 ) | ( n_n135 ) | ( wire80 ) | ( wire204 ) ;
 assign wire17976 = ( n_n6267 ) | ( n_n6266 ) | ( n_n6270 ) | ( wire3774 ) ;
 assign wire17977 = ( wire157  &  n_n47 ) | ( wire172  &  n_n47 ) ;
 assign wire17979 = ( wire52  &  n_n43 ) | ( n_n43  &  wire139 ) ;
 assign wire17980 = ( wire129  &  n_n43 ) | ( n_n43  &  wire63 ) | ( n_n43  &  wire48 ) ;
 assign wire17985 = ( n_n41  &  wire85 ) | ( n_n41  &  n_n198 ) | ( n_n41  &  n_n214 ) ;
 assign wire17987 = ( wire17985 ) | ( n_n41  &  wire142 ) | ( n_n41  &  wire180 ) ;
 assign wire17988 = ( wire524 ) | ( wire359 ) | ( n_n4476 ) | ( wire3759 ) ;
 assign wire17989 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire17993 = ( wire62 ) | ( wire240 ) | ( wire107 ) | ( wire17989 ) ;
 assign wire17995 = ( wire497 ) | ( n_n41  &  wire70 ) | ( n_n41  &  wire51 ) ;
 assign wire17996 = ( n_n41  &  n_n83 ) | ( n_n41  &  n_n171 ) | ( n_n41  &  wire69 ) ;
 assign wire17999 = ( wire694 ) | ( n_n3542 ) | ( wire17996 ) ;
 assign wire18000 = ( wire426 ) | ( wire3747 ) | ( wire17999 ) ;
 assign wire18001 = ( wire3755 ) | ( wire17987 ) | ( wire17988 ) | ( wire17995 ) ;
 assign wire18002 = ( n_n39  &  wire110 ) | ( n_n39  &  wire726  &  n_n156 ) ;
 assign wire18003 = ( wire207  &  n_n39 ) | ( n_n39  &  wire248 ) | ( n_n39  &  n_n78 ) ;
 assign wire18004 = ( n_n184  &  wire719 ) | ( n_n199  &  wire725 ) ;
 assign wire18007 = ( n_n156  &  wire719 ) | ( n_n149  &  wire725 ) ;
 assign wire18010 = ( n_n41  &  n_n57 ) | ( n_n39  &  wire104 ) ;
 assign wire18012 = ( wire18010 ) | ( n_n41  &  wire245 ) | ( n_n41  &  wire182 ) ;
 assign wire18013 = ( n_n41  &  wire1807 ) | ( n_n41  &  wire1811 ) ;
 assign wire18014 = ( wire720  &  n_n149 ) | ( n_n216  &  wire719 ) ;
 assign wire18017 = ( n_n71  &  n_n41 ) | ( n_n41  &  n_n150 ) | ( n_n41  &  wire141 ) ;
 assign wire18018 = ( wire442 ) | ( n_n41  &  wire234 ) | ( n_n41  &  wire84 ) ;
 assign wire18019 = ( wire18017 ) | ( n_n41  &  wire1812 ) ;
 assign wire18021 = ( n_n39  &  n_n177  &  wire719 ) | ( n_n39  &  n_n170  &  wire719 ) ;
 assign wire18023 = ( wire434 ) | ( wire18021 ) | ( n_n39  &  wire249 ) ;
 assign wire18024 = ( wire3723 ) | ( n_n39  &  n_n84 ) | ( n_n39  &  wire279 ) ;
 assign wire18026 = ( wire18002 ) | ( wire18003 ) | ( wire18023 ) | ( wire18024 ) ;
 assign wire18027 = ( wire18012 ) | ( wire18013 ) | ( wire18018 ) | ( wire18019 ) ;
 assign wire18028 = ( n_n47  &  wire149 ) | ( n_n47  &  wire147 ) ;
 assign wire18032 = ( wire419 ) | ( wire3710 ) | ( n_n47  &  wire151 ) ;
 assign wire18035 = ( n_n47  &  wire129 ) | ( n_n47  &  wire130 ) ;
 assign wire18036 = ( n_n47  &  wire46 ) | ( n_n47  &  wire124 ) ;
 assign wire18039 = ( n_n3561 ) | ( wire3702 ) | ( wire18035 ) | ( wire18036 ) ;
 assign wire18044 = ( wire3696 ) | ( n_n113  &  wire256 ) ;
 assign wire18049 = ( wire124 ) | ( wire48 ) ;
 assign wire18050 = ( wire168 ) | ( wire52 ) | ( wire128 ) ;
 assign wire18051 = ( wire129 ) | ( wire130 ) | ( wire139 ) | ( wire63 ) ;
 assign wire18053 = ( n_n184  &  wire729 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire18057 = ( wire3700 ) | ( wire3701 ) | ( n_n125  &  n_n57 ) ;
 assign wire18058 = ( wire3690 ) | ( n_n125  &  wire1751 ) ;
 assign wire18063 = ( wire135 ) | ( wire125 ) | ( n_n216  &  wire725 ) ;
 assign wire18064 = ( wire55 ) | ( wire158 ) | ( wire133 ) | ( wire127 ) ;
 assign wire18067 = ( n_n138 ) | ( n_n132 ) | ( wire153 ) | ( wire78 ) ;
 assign wire18068 = ( n_n53 ) | ( n_n135 ) | ( wire80 ) | ( wire204 ) ;
 assign wire18069 = ( wire172 ) | ( wire150 ) | ( wire217 ) | ( wire173 ) ;
 assign wire18071 = ( wire445 ) | ( wire157  &  n_n108 ) ;
 assign wire18074 = ( wire131 ) | ( wire126 ) ;
 assign wire18075 = ( wire132 ) | ( wire134 ) | ( wire149 ) | ( wire147 ) ;
 assign wire18076 = ( n_n108  &  wire1489 ) | ( n_n108  &  wire18074 ) | ( n_n108  &  wire18075 ) ;
 assign wire18078 = ( n_n3489 ) | ( wire3685 ) | ( wire18071 ) | ( wire18076 ) ;
 assign wire18081 = ( wire217 ) | ( wire150 ) ;
 assign wire18082 = ( n_n135 ) | ( n_n132 ) | ( wire80 ) | ( wire78 ) ;
 assign wire18083 = ( n_n53 ) | ( wire157 ) | ( wire173 ) | ( wire204 ) ;
 assign wire18085 = ( n_n125  &  wire85 ) | ( n_n125  &  wire142 ) | ( n_n125  &  n_n214 ) ;
 assign wire18087 = ( wire127 ) | ( wire153 ) | ( n_n191  &  wire719 ) ;
 assign wire18088 = ( wire172 ) | ( wire133 ) | ( n_n63 ) | ( wire135 ) ;
 assign wire18089 = ( n_n212  &  wire55 ) | ( n_n212  &  wire158 ) ;
 assign wire18091 = ( wire18089 ) | ( n_n212  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign wire18092 = ( (~ i_9_)  &  i_10_  &  i_11_  &  wire720 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire18096 = ( n_n3592 ) | ( wire538 ) | ( wire539 ) | ( wire3665 ) ;
 assign wire18097 = ( wire3671 ) | ( wire3676 ) | ( wire18085 ) | ( wire18091 ) ;
 assign wire18098 = ( n_n216  &  wire719 ) | ( n_n199  &  wire725 ) ;
 assign wire18102 = ( wire220 ) | ( wire234 ) ;
 assign wire18103 = ( wire60 ) | ( wire242 ) | ( n_n184  &  wire719 ) ;
 assign wire18104 = ( wire218 ) | ( wire160 ) | ( wire171 ) | ( wire18098 ) ;
 assign wire18106 = ( n_n125  &  wire182 ) | ( n_n125  &  wire141 ) ;
 assign wire18107 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire720 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire720 ) ;
 assign wire18111 = ( n_n176 ) | ( wire62 ) | ( wire107 ) | ( wire18107 ) ;
 assign wire18113 = ( wire394 ) | ( n_n125  &  wire51 ) | ( n_n125  &  wire100 ) ;
 assign wire18117 = ( n_n148 ) | ( wire90 ) | ( wire69 ) | ( wire225 ) ;
 assign wire18119 = ( wire479 ) | ( wire698 ) | ( wire3653 ) ;
 assign wire18120 = ( wire3658 ) | ( wire3662 ) | ( wire18106 ) | ( wire18113 ) ;
 assign wire18122 = ( n_n212  &  wire130 ) | ( n_n212  &  wire63 ) ;
 assign wire18125 = ( wire132  &  n_n212 ) | ( n_n212  &  wire149 ) ;
 assign wire18128 = ( n_n212  &  wire168 ) | ( n_n212  &  wire151 ) ;
 assign wire18129 = ( n_n212  &  wire181 ) | ( n_n212  &  wire48 ) ;
 assign wire18132 = ( n_n4518 ) | ( wire3643 ) | ( wire18128 ) | ( wire18129 ) ;
 assign wire18134 = ( n_n3501 ) | ( n_n3500 ) | ( wire18132 ) ;
 assign wire18135 = ( wire18096 ) | ( wire18097 ) | ( wire18119 ) | ( wire18120 ) ;
 assign wire18136 = ( n_n47  &  wire55 ) | ( n_n47  &  wire125 ) ;
 assign wire18137 = ( n_n47  &  wire176 ) | ( n_n47  &  wire123 ) | ( n_n47  &  wire1791 ) ;
 assign wire18140 = ( n_n3482 ) | ( wire3773 ) | ( wire17976 ) | ( wire17977 ) ;
 assign wire18141 = ( n_n3555 ) | ( wire18136 ) | ( wire18137 ) | ( wire18140 ) ;
 assign wire18142 = ( wire18000 ) | ( wire18001 ) | ( wire18026 ) | ( wire18027 ) ;
 assign wire18144 = ( n_n3451 ) | ( wire18134 ) | ( wire18135 ) ;
 assign wire18145 = ( n_n5144 ) | ( wire17924 ) | ( n_n31  &  wire1601 ) ;
 assign wire18146 = ( n_n3454 ) | ( wire17951 ) | ( wire17952 ) | ( wire17954 ) ;
 assign wire18148 = ( n_n3456 ) | ( wire18145 ) | ( wire18146 ) ;
 assign wire18150 = ( n_n9  &  n_n191  &  wire717 ) | ( n_n9  &  wire717  &  n_n149 ) ;
 assign wire18154 = ( wire3624 ) | ( n_n19  &  n_n157  &  n_n218 ) ;
 assign wire18155 = ( n_n7241 ) | ( n_n17  &  wire743 ) | ( n_n17  &  wire1524 ) ;
 assign wire18157 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire18158 = ( n_n5144 ) | ( n_n157  &  n_n48  &  n_n219 ) ;
 assign wire18159 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n111 ) ;
 assign wire18160 = ( n_n17  &  n_n48  &  n_n219 ) | ( n_n17  &  n_n219  &  n_n218 ) ;
 assign wire18161 = ( n_n162  &  n_n157  &  n_n219 ) | ( n_n157  &  n_n219  &  n_n218 ) ;
 assign wire18163 = ( wire18161 ) | ( wire18160 ) ;
 assign wire18164 = ( wire18158 ) | ( wire18159 ) | ( n_n14  &  wire253 ) ;
 assign wire18167 = ( wire3621 ) | ( wire3622 ) | ( wire18163 ) | ( wire18164 ) ;
 assign wire18168 = ( n_n46  &  wire181 ) | ( n_n47  &  wire48 ) ;
 assign wire18169 = ( n_n47  &  wire63 ) | ( n_n46  &  wire47 ) ;
 assign wire18172 = ( n_n46  &  wire168 ) | ( n_n47  &  wire181 ) ;
 assign wire18173 = ( n_n46  &  wire151 ) | ( n_n47  &  wire151 ) ;
 assign wire18174 = ( n_n47  &  wire143 ) | ( n_n47  &  wire154 ) | ( n_n47  &  wire47 ) ;
 assign wire18178 = ( n_n47  &  wire129 ) | ( n_n47  &  wire124 ) ;
 assign wire18180 = ( wire3588 ) | ( wire18178 ) | ( n_n46  &  wire875 ) ;
 assign wire18182 = ( n_n47  &  wire176 ) | ( n_n46  &  wire131 ) ;
 assign wire18184 = ( wire674 ) | ( n_n46  &  wire55 ) | ( n_n46  &  wire127 ) ;
 assign wire18185 = ( wire546 ) | ( wire18182 ) | ( n_n47  &  wire123 ) ;
 assign wire18186 = ( wire671 ) | ( n_n47  &  wire130 ) ;
 assign wire18187 = ( n_n3889 ) | ( wire4088 ) | ( n_n47  &  wire46 ) ;
 assign wire18188 = ( n_n184  &  wire719 ) | ( n_n216  &  wire725 ) ;
 assign wire18190 = ( n_n46  &  wire176 ) | ( n_n47  &  n_n63 ) ;
 assign wire18191 = ( n_n47  &  n_n140 ) | ( n_n47  &  wire247 ) | ( n_n47  &  wire125 ) ;
 assign wire18192 = ( wire18190 ) | ( wire3575 ) ;
 assign wire18193 = ( wire3580 ) | ( wire3581 ) | ( wire18191 ) ;
 assign wire18194 = ( n_n191  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n170  &  wire725 ) ;
 assign wire18196 = ( n_n177  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire18198 = ( wire217 ) | ( wire18196 ) ;
 assign wire18199 = ( wire186 ) | ( wire209 ) | ( wire174 ) ;
 assign wire18200 = ( wire651 ) | ( n_n46  &  n_n177  &  wire719 ) ;
 assign wire18201 = ( wire3570 ) | ( n_n47  &  wire18198 ) | ( n_n47  &  wire18199 ) ;
 assign wire18202 = ( n_n47  &  wire55 ) | ( n_n46  &  wire134 ) ;
 assign wire18205 = ( wire688 ) | ( n_n3555 ) | ( wire3563 ) | ( wire18202 ) ;
 assign wire18206 = ( wire18192 ) | ( wire18193 ) | ( wire18200 ) | ( wire18201 ) ;
 assign wire18209 = ( n_n47  &  wire149 ) | ( n_n46  &  wire46 ) ;
 assign wire18210 = ( wire132  &  n_n47 ) | ( n_n47  &  wire147 ) | ( n_n47  &  wire126 ) ;
 assign wire18212 = ( wire18209 ) | ( wire18210 ) | ( n_n46  &  wire1271 ) ;
 assign wire18213 = ( wire18184 ) | ( wire18185 ) | ( wire18186 ) | ( wire18187 ) ;
 assign wire18214 = ( wire18213 ) | ( wire18212 ) ;
 assign wire18215 = ( n_n3033 ) | ( wire18205 ) | ( wire18206 ) ;
 assign wire18220 = ( n_n5144 ) | ( n_n6271 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire18221 = ( n_n6267 ) | ( n_n6266 ) | ( n_n6270 ) | ( n_n6269 ) ;
 assign wire18222 = ( n_n6268 ) | ( n_n53  &  n_n46 ) | ( wire157  &  n_n46 ) ;
 assign wire18225 = ( n_n3085 ) | ( wire18220 ) | ( wire18221 ) | ( wire18222 ) ;
 assign wire18230 = ( wire54 ) | ( wire399 ) | ( wire268 ) ;
 assign wire18232 = ( n_n6384 ) | ( n_n3419 ) | ( n_n41  &  wire1036 ) ;
 assign wire18234 = ( n_n53  &  n_n46 ) | ( n_n41  &  n_n202 ) ;
 assign wire18237 = ( n_n4308 ) | ( n_n3421 ) | ( wire391 ) | ( wire18234 ) ;
 assign wire18238 = ( wire3533 ) | ( wire3607 ) | ( wire4260 ) | ( wire17554 ) ;
 assign wire18242 = ( wire111 ) | ( wire206 ) | ( wire368 ) ;
 assign wire18243 = ( wire3526 ) | ( wire3531 ) | ( n_n40  &  n_n95 ) ;
 assign wire18244 = ( wire3527 ) | ( wire3545 ) | ( wire18232 ) ;
 assign wire18245 = ( wire18237 ) | ( wire18238 ) | ( wire18243 ) ;
 assign wire18251 = ( wire93 ) | ( wire273 ) | ( n_n184  &  wire729 ) ;
 assign wire18252 = ( n_n3417 ) | ( n_n41  &  wire1174 ) ;
 assign wire18253 = ( wire729  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign wire18260 = ( n_n77 ) | ( wire59 ) | ( wire117 ) | ( wire281 ) ;
 assign wire18264 = ( n_n41  &  n_n83 ) | ( n_n41  &  n_n171 ) | ( n_n41  &  wire469 ) ;
 assign wire18266 = ( n_n3415 ) | ( wire18264 ) | ( n_n40  &  wire1331 ) ;
 assign wire18267 = ( wire3524 ) | ( wire18266 ) | ( n_n40  &  n_n89 ) ;
 assign wire18268 = ( wire3515 ) | ( wire3516 ) | ( wire3520 ) | ( wire18252 ) ;
 assign wire18269 = ( n_n138  &  n_n40 ) | ( n_n184  &  n_n40  &  wire725 ) ;
 assign wire18270 = ( n_n41  &  wire182 ) | ( wire172  &  n_n40 ) ;
 assign wire18272 = ( wire3498 ) | ( wire18269 ) | ( n_n40  &  wire217 ) ;
 assign wire18273 = ( n_n5067 ) | ( n_n5059 ) | ( wire18270 ) ;
 assign wire18278 = ( wire724  &  n_n156 ) | ( wire717  &  n_n156 ) ;
 assign wire18281 = ( wire118 ) | ( wire298 ) | ( wire18278 ) ;
 assign wire18283 = ( n_n6492 ) | ( n_n3413 ) | ( n_n40  &  wire1432 ) ;
 assign wire18287 = ( wire673 ) | ( wire3472 ) | ( wire3479 ) | ( wire3480 ) ;
 assign wire18288 = ( n_n5075 ) | ( n_n5070 ) | ( wire3471 ) | ( wire18287 ) ;
 assign wire18290 = ( n_n5144 ) | ( wire18244 ) | ( wire18245 ) ;
 assign wire18292 = ( n_n3029 ) | ( wire18267 ) | ( wire18268 ) | ( wire18290 ) ;
 assign wire18294 = ( wire3550 ) | ( wire3551 ) | ( wire182  &  n_n40 ) ;
 assign wire18295 = ( n_n5052 ) | ( n_n5055 ) | ( n_n5058 ) | ( wire4900 ) ;
 assign wire18297 = ( wire3469 ) | ( wire3470 ) | ( wire18294 ) | ( wire18295 ) ;
 assign wire18298 = ( n_n159  &  n_n218  &  wire747 ) ;
 assign wire18299 = ( n_n5144 ) | ( n_n51  &  wire751 ) | ( n_n51  &  wire18298 ) ;
 assign wire18300 = ( n_n33  &  n_n132 ) | ( n_n33  &  n_n149  &  wire728 ) ;
 assign wire18301 = ( n_n33  &  n_n128 ) | ( n_n33  &  wire48 ) | ( n_n33  &  wire173 ) ;
 assign wire18302 = ( wire130  &  n_n32 ) | ( wire139  &  n_n32 ) | ( n_n32  &  wire128 ) ;
 assign wire18307 = ( n_n5144 ) | ( n_n33  &  n_n191  &  wire719 ) ;
 assign wire18310 = ( wire587 ) | ( wire18307 ) | ( n_n32  &  wire124 ) ;
 assign wire18311 = ( n_n2732 ) | ( n_n2728 ) | ( wire3461 ) | ( wire18300 ) ;
 assign wire18316 = ( wire3435 ) | ( n_n4  &  wire729  &  n_n156 ) ;
 assign wire18318 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n111 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n111 ) ;
 assign wire18321 = ( wire431 ) | ( wire529 ) | ( wire18318 ) ;
 assign wire18323 = ( n_n7252 ) | ( wire389 ) | ( wire3425 ) | ( wire18321 ) ;
 assign wire18324 = ( n_n5144 ) | ( n_n157  &  n_n219  &  n_n111 ) ;
 assign wire18325 = ( wire18324 ) | ( n_n9  &  wire717  &  n_n149 ) ;
 assign wire18328 = ( n_n3389 ) | ( wire388 ) | ( n_n9  &  wire770 ) ;
 assign wire18329 = ( wire3415 ) | ( wire18325 ) | ( n_n10  &  wire145 ) ;
 assign wire18330 = ( wire3437 ) | ( wire3438 ) | ( wire18328 ) ;
 assign wire18332 = ( n_n5144 ) | ( wire267  &  n_n149  &  wire725 ) ;
 assign wire18334 = ( n_n184  &  wire719 ) | ( n_n184  &  wire725 ) | ( n_n184  &  wire728 ) ;
 assign wire18337 = ( wire130 ) | ( wire139 ) | ( wire18334 ) ;
 assign wire18342 = ( n_n113  &  n_n115 ) | ( n_n42  &  n_n183 ) ;
 assign wire18345 = ( wire3404 ) | ( n_n43  &  wire1786 ) ;
 assign wire18348 = ( wire526 ) | ( wire3397 ) | ( n_n42  &  n_n138 ) ;
 assign wire18352 = ( wire3385 ) | ( n_n42  &  n_n191  &  wire720 ) ;
 assign wire18353 = ( n_n1575 ) | ( wire3392 ) | ( n_n42  &  wire1782 ) ;
 assign wire18354 = ( n_n1566 ) | ( wire3396 ) | ( wire18348 ) | ( wire18352 ) ;
 assign wire18355 = ( n_n2715 ) | ( wire3409 ) | ( wire3410 ) | ( wire18353 ) ;
 assign wire18358 = ( n_n41  &  wire182 ) | ( wire182  &  n_n40 ) ;
 assign wire18360 = ( n_n5055 ) | ( n_n41  &  wire245 ) | ( n_n41  &  wire150 ) ;
 assign wire18361 = ( n_n5059 ) | ( n_n5058 ) | ( wire18358 ) ;
 assign wire18367 = ( n_n7346 ) | ( n_n5319 ) | ( n_n3  &  wire185 ) ;
 assign wire18370 = ( n_n7263 ) | ( n_n5319 ) | ( n_n7264 ) ;
 assign wire18371 = ( n_n7242 ) | ( wire463 ) | ( n_n7262 ) ;
 assign wire18372 = ( wire428 ) | ( n_n3276 ) | ( wire462 ) | ( wire16884 ) ;
 assign wire18374 = ( wire18372 ) | ( n_n14  &  wire270 ) ;
 assign wire18375 = ( wire3550 ) | ( wire3551 ) | ( wire18370 ) | ( wire18371 ) ;
 assign wire18377 = ( n_n3176 ) | ( wire3374 ) | ( wire3375 ) | ( wire3376 ) ;
 assign wire18384 = ( wire94 ) | ( wire324 ) | ( n_n184  &  wire729 ) ;
 assign wire18385 = ( n_n5113 ) | ( n_n46  &  wire868 ) ;
 assign wire18386 = ( n_n216  &  wire721 ) | ( n_n199  &  wire725 ) | ( n_n216  &  wire725 ) ;
 assign wire18388 = ( wire729  &  n_n156 ) | ( n_n199  &  wire719 ) ;
 assign wire18391 = ( wire212 ) | ( wire198 ) | ( wire18388 ) ;
 assign wire18393 = ( n_n5107 ) | ( wire3342 ) | ( wire172  &  n_n47 ) ;
 assign wire18394 = ( n_n191  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire18397 = ( n_n5103 ) | ( wire666 ) | ( wire3337 ) ;
 assign wire18398 = ( wire3338 ) | ( wire4857 ) | ( n_n46  &  wire209 ) ;
 assign wire18401 = ( n_n5109 ) | ( n_n47  &  wire1326 ) ;
 assign wire18402 = ( wire3333 ) | ( wire3343 ) | ( wire18393 ) ;
 assign wire18403 = ( wire18397 ) | ( wire18398 ) | ( wire18401 ) ;
 assign wire18408 = ( wire93 ) | ( wire54 ) | ( wire273 ) ;
 assign wire18409 = ( wire498 ) | ( n_n46  &  wire951 ) ;
 assign wire18411 = ( n_n5319 ) | ( n_n46  &  wire168 ) ;
 assign wire18413 = ( wire577 ) | ( n_n46  &  wire68 ) | ( n_n46  &  wire74 ) ;
 assign wire18414 = ( wire481 ) | ( wire18411 ) | ( n_n46  &  wire151 ) ;
 assign wire18416 = ( n_n199  &  wire723 ) | ( n_n199  &  wire729 ) | ( n_n199  &  wire727 ) ;
 assign wire18418 = ( n_n5319 ) | ( n_n47  &  wire151 ) ;
 assign wire18420 = ( wire3312 ) | ( wire3313 ) | ( wire18418 ) ;
 assign wire18421 = ( wire3325 ) | ( wire18420 ) | ( n_n47  &  wire98 ) ;
 assign wire18422 = ( wire3328 ) | ( wire18409 ) | ( wire18413 ) | ( wire18414 ) ;
 assign wire18424 = ( wire179 ) | ( wire120 ) ;
 assign wire18425 = ( wire118 ) | ( wire324 ) | ( wire729  &  n_n177 ) ;
 assign wire18426 = ( wire729  &  n_n156 ) | ( wire720  &  n_n156 ) | ( n_n156  &  wire715 ) ;
 assign wire18429 = ( n_n5111 ) | ( n_n46  &  wire18424 ) | ( n_n46  &  wire18425 ) ;
 assign wire18432 = ( wire117 ) | ( wire294 ) | ( wire729  &  n_n177 ) ;
 assign wire18433 = ( wire3300 ) | ( wire3353 ) | ( n_n47  &  wire53 ) ;
 assign wire18434 = ( wire3301 ) | ( wire3349 ) | ( wire18385 ) ;
 assign wire18436 = ( wire3308 ) | ( wire18429 ) | ( wire18433 ) | ( wire18434 ) ;
 assign wire18437 = ( wire18402 ) | ( wire18403 ) | ( wire18421 ) | ( wire18422 ) ;
 assign wire18444 = ( wire132 ) | ( wire52 ) | ( wire126 ) ;
 assign wire18445 = ( n_n41  &  n_n83 ) | ( n_n41  &  n_n171 ) | ( n_n41  &  wire1544 ) ;
 assign wire18450 = ( wire137 ) | ( wire149 ) | ( wire131 ) ;
 assign wire18452 = ( wire3296 ) | ( wire3298 ) | ( wire3299 ) | ( wire18445 ) ;
 assign wire18454 = ( wire3498 ) | ( wire18269 ) | ( n_n40  &  wire217 ) ;
 assign wire18455 = ( n_n5067 ) | ( wire673 ) | ( wire172  &  n_n40 ) ;
 assign wire18457 = ( wire726  &  n_n149 ) | ( wire724  &  n_n149 ) ;
 assign wire18461 = ( n_n5319 ) | ( n_n5075 ) | ( wire3479 ) | ( wire3480 ) ;
 assign wire18462 = ( n_n5070 ) | ( wire3279 ) | ( wire3280 ) ;
 assign wire18467 = ( wire55 ) | ( wire156 ) | ( wire724  &  n_n156 ) ;
 assign wire18469 = ( wire363 ) | ( wire3275 ) | ( n_n40  &  wire1383 ) ;
 assign wire18471 = ( n_n41  &  n_n210 ) | ( n_n41  &  n_n107 ) | ( n_n41  &  n_n214 ) ;
 assign wire18474 = ( n_n5319 ) | ( n_n46  &  n_n177  &  wire725 ) ;
 assign wire18475 = ( wire3271 ) | ( wire18471 ) | ( wire18474 ) ;
 assign wire18476 = ( n_n47  &  wire1425 ) | ( n_n46  &  wire1424 ) ;
 assign wire18481 = ( wire143 ) | ( wire47 ) | ( n_n216  &  wire724 ) ;
 assign wire18482 = ( wire361 ) | ( n_n41  &  wire1493 ) ;
 assign wire18486 = ( wire359 ) | ( wire3258 ) | ( n_n40  &  wire1386 ) ;
 assign wire18487 = ( wire3264 ) | ( wire18475 ) | ( wire18476 ) | ( wire18482 ) ;
 assign wire18488 = ( n_n5144 ) | ( wire3291 ) | ( wire3292 ) | ( wire18452 ) ;
 assign wire18490 = ( n_n3170 ) | ( wire18486 ) | ( wire18487 ) | ( wire18488 ) ;
 assign wire18492 = ( n_n7263 ) | ( n_n7265 ) | ( n_n7264 ) ;
 assign wire18493 = ( wire711 ) | ( n_n10  &  wire729  &  n_n191 ) ;
 assign wire18495 = ( wire18492 ) | ( wire18493 ) | ( wire878  &  wire877 ) ;
 assign wire18496 = ( wire529 ) | ( n_n9  &  wire77 ) | ( wire77  &  n_n6 ) ;
 assign wire18498 = ( wire3244 ) | ( n_n6  &  wire879 ) | ( n_n5  &  wire879 ) ;
 assign wire18499 = ( wire454 ) | ( wire3245 ) | ( wire18496 ) ;
 assign wire18504 = ( n_n3276 ) | ( wire462 ) | ( n_n2948 ) | ( wire16884 ) ;
 assign wire18505 = ( i_7_  &  i_6_  &  wire743 ) | ( (~ i_7_)  &  i_6_  &  wire743 ) | ( i_7_  &  (~ i_6_)  &  wire743 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire743 ) | ( i_7_  &  i_6_  &  wire745 ) | ( (~ i_7_)  &  i_6_  &  wire745 ) | ( i_7_  &  (~ i_6_)  &  wire745 ) | ( (~ i_7_)  &  (~ i_6_)  &  wire745 ) ;
 assign wire18507 = ( n_n231 ) | ( wire18504 ) | ( wire18505 ) ;
 assign wire18508 = ( wire3256 ) | ( wire3257 ) | ( wire18495 ) | ( wire18507 ) ;
 assign wire18509 = ( n_n5144 ) | ( n_n18  &  n_n159  &  n_n218 ) ;
 assign wire18510 = ( wire18509 ) | ( n_n3  &  wire717  &  n_n149 ) ;
 assign wire18512 = ( wire708 ) | ( wire3234 ) | ( wire18510 ) ;
 assign wire18517 = ( wire137 ) | ( wire55 ) | ( wire131 ) ;
 assign wire18521 = ( wire137 ) | ( wire130 ) | ( wire131 ) ;
 assign wire18522 = ( wire3229 ) | ( n_n123  &  wire52 ) ;
 assign wire18526 = ( wire3224 ) | ( wire3225 ) | ( n_n125  &  wire147 ) ;
 assign wire18527 = ( wire3230 ) | ( wire3232 ) | ( wire3233 ) | ( wire18522 ) ;
 assign wire18528 = ( n_n177  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire18529 = ( n_n177  &  wire719 ) | ( n_n170  &  wire725 ) ;
 assign wire18533 = ( wire3219 ) | ( wire3222 ) | ( wire3223 ) ;
 assign wire18534 = ( n_n199  &  wire719 ) | ( n_n216  &  wire725 ) ;
 assign wire18537 = ( n_n184  &  wire719 ) | ( n_n199  &  wire719 ) | ( n_n199  &  wire728 ) ;
 assign wire18540 = ( wire176 ) | ( wire153 ) | ( wire18537 ) ;
 assign wire18541 = ( n_n2859 ) | ( n_n125  &  wire1395 ) ;
 assign wire18546 = ( n_n123  &  wire133 ) | ( n_n123  &  wire959 ) ;
 assign wire18547 = ( wire18546 ) | ( n_n125  &  wire960 ) ;
 assign wire18548 = ( wire3217 ) | ( wire3220 ) | ( wire18533 ) | ( wire18541 ) ;
 assign wire18553 = ( wire168 ) | ( wire68 ) | ( wire74 ) ;
 assign wire18555 = ( n_n125  &  wire52 ) | ( n_n123  &  wire1729 ) ;
 assign wire18559 = ( wire151 ) | ( wire143 ) | ( wire47 ) ;
 assign wire18560 = ( wire3201 ) | ( n_n123  &  wire74 ) ;
 assign wire18562 = ( wire3202 ) | ( wire3209 ) | ( wire3210 ) | ( wire18560 ) ;
 assign wire18564 = ( n_n5144 ) | ( n_n53  &  n_n123 ) | ( wire157  &  n_n123 ) ;
 assign wire18565 = ( wire4323 ) | ( wire4324 ) | ( wire18564 ) ;
 assign wire18567 = ( n_n2813 ) | ( wire18547 ) | ( wire18548 ) | ( wire18562 ) ;
 assign wire18568 = ( n_n5144 ) | ( n_n18  &  n_n159  &  n_n218 ) ;
 assign wire18572 = ( n_n5319 ) | ( wire430 ) | ( wire684 ) | ( wire3195 ) ;
 assign wire18575 = ( n_n197  &  wire181 ) | ( n_n212  &  wire48 ) ;
 assign wire18576 = ( n_n212  &  wire52 ) | ( n_n212  &  wire129 ) | ( n_n212  &  wire63 ) ;
 assign wire18577 = ( n_n2777 ) | ( wire18575 ) ;
 assign wire18578 = ( wire18576 ) | ( n_n197  &  wire1602 ) ;
 assign wire18581 = ( wire132  &  n_n212 ) | ( n_n197  &  wire149 ) ;
 assign wire18582 = ( wire132  &  n_n197 ) | ( n_n212  &  wire149 ) ;
 assign wire18583 = ( n_n197  &  wire147 ) | ( n_n197  &  wire126 ) | ( n_n197  &  wire46 ) ;
 assign wire18586 = ( n_n197  &  wire52 ) | ( n_n212  &  wire130 ) ;
 assign wire18587 = ( n_n197  &  wire129 ) | ( n_n197  &  wire127 ) ;
 assign wire18588 = ( wire137  &  n_n212 ) | ( n_n212  &  wire46 ) ;
 assign wire18593 = ( wire594 ) | ( wire681 ) | ( wire504 ) | ( wire18586 ) ;
 assign wire18594 = ( n_n2770 ) | ( n_n3601 ) | ( wire18587 ) | ( wire18588 ) ;
 assign wire18596 = ( n_n197  &  n_n134 ) | ( n_n212  &  wire186 ) ;
 assign wire18598 = ( n_n197  &  wire125 ) | ( n_n197  &  n_n216  &  wire725 ) ;
 assign wire18600 = ( n_n197  &  wire176 ) | ( n_n212  &  wire125 ) ;
 assign wire18602 = ( n_n4686 ) | ( wire704 ) | ( wire18598 ) ;
 assign wire18603 = ( wire3154 ) | ( wire3155 ) | ( wire18600 ) ;
 assign wire18605 = ( n_n197  &  wire158 ) | ( n_n197  &  wire133 ) ;
 assign wire18607 = ( wire565 ) | ( n_n212  &  wire55 ) | ( n_n212  &  wire158 ) ;
 assign wire18608 = ( wire532 ) | ( wire18605 ) | ( n_n197  &  wire123 ) ;
 assign wire18609 = ( n_n191  &  wire721 ) | ( n_n191  &  wire725 ) | ( n_n170  &  wire725 ) ;
 assign wire18611 = ( n_n177  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire18614 = ( wire689 ) | ( wire3142 ) | ( wire18596 ) ;
 assign wire18616 = ( wire18602 ) | ( wire18603 ) | ( wire18607 ) | ( wire18608 ) ;
 assign wire18617 = ( n_n149  &  wire721 ) | ( n_n156  &  wire725 ) | ( n_n149  &  wire725 ) ;
 assign wire18619 = ( n_n5144 ) | ( n_n212  &  n_n156  &  wire725 ) ;
 assign wire18621 = ( wire3135 ) | ( wire3136 ) | ( wire18619 ) ;
 assign wire18623 = ( n_n2747 ) | ( wire3143 ) | ( wire18614 ) | ( wire18616 ) ;
 assign wire18624 = ( n_n42  &  wire139 ) | ( n_n43  &  wire139 ) ;
 assign wire18625 = ( wire52  &  n_n43 ) | ( wire129  &  n_n43 ) ;
 assign wire18626 = ( n_n43  &  wire124 ) | ( n_n42  &  wire128 ) | ( n_n43  &  wire128 ) ;
 assign wire18631 = ( wire672 ) | ( wire3123 ) | ( n_n59  &  n_n43 ) ;
 assign wire18632 = ( wire3124 ) | ( wire4102 ) | ( n_n43  &  wire222 ) ;
 assign wire18635 = ( wire155 ) | ( wire215 ) | ( wire720  &  n_n156 ) ;
 assign wire18637 = ( n_n101  &  wire224 ) | ( n_n101  &  wire250 ) | ( n_n101  &  wire57 ) ;
 assign wire18638 = ( wire4735 ) | ( wire18637 ) | ( n_n108  &  wire69 ) ;
 assign wire18641 = ( wire4372 ) | ( wire4838 ) | ( wire4839 ) | ( wire17469 ) ;
 assign wire18642 = ( wire3113 ) | ( n_n101  &  wire218 ) | ( n_n101  &  wire141 ) ;
 assign wire18644 = ( wire150 ) | ( n_n184  &  wire719 ) | ( n_n184  &  wire728 ) ;
 assign wire18645 = ( wire222 ) | ( wire256 ) | ( n_n170  &  wire719 ) ;
 assign wire18646 = ( n_n184  &  wire719 ) | ( n_n191  &  wire725 ) ;
 assign wire18649 = ( wire78 ) | ( wire252 ) | ( wire18646 ) ;
 assign wire18650 = ( n_n4981 ) | ( n_n101  &  wire18644 ) | ( n_n101  &  wire18645 ) ;
 assign wire18652 = ( n_n5000 ) | ( wire511 ) | ( n_n101  &  wire84 ) ;
 assign wire18653 = ( wire3102 ) | ( n_n108  &  wire84 ) | ( n_n108  &  wire220 ) ;
 assign wire18655 = ( n_n4996 ) | ( n_n4994 ) | ( wire18652 ) | ( wire18653 ) ;
 assign wire18656 = ( wire3111 ) | ( wire18641 ) | ( wire18642 ) | ( wire18650 ) ;
 assign wire18657 = ( n_n184  &  wire729 ) | ( n_n184  &  wire726 ) | ( n_n184  &  wire720 ) ;
 assign wire18662 = ( wire51 ) | ( wire210 ) | ( n_n184  &  wire720 ) ;
 assign wire18663 = ( n_n5021 ) | ( n_n101  &  wire1723 ) ;
 assign wire18665 = ( n_n5739 ) | ( wire440 ) | ( wire760 ) ;
 assign wire18668 = ( n_n4904 ) | ( n_n5037 ) | ( wire657 ) | ( wire18665 ) ;
 assign wire18669 = ( n_n4900 ) | ( n_n5033 ) | ( wire4937 ) ;
 assign wire18670 = ( wire4935 ) | ( wire18668 ) | ( n_n108  &  wire1844 ) ;
 assign wire18671 = ( wire3098 ) | ( wire18663 ) | ( wire18669 ) ;
 assign wire18676 = ( wire100 ) | ( wire272 ) | ( n_n177  &  wire720 ) ;
 assign wire18677 = ( n_n5019 ) | ( n_n101  &  wire1689 ) ;
 assign wire18679 = ( n_n101  &  wire208 ) | ( n_n101  &  wire225 ) | ( n_n101  &  wire148 ) ;
 assign wire18680 = ( n_n5011 ) | ( wire591 ) | ( n_n108  &  wire250 ) ;
 assign wire18682 = ( wire4933 ) | ( wire4934 ) | ( wire18679 ) | ( wire18680 ) ;
 assign wire18683 = ( wire3093 ) | ( wire3118 ) | ( wire18638 ) | ( wire18677 ) ;
 assign wire18685 = ( wire18655 ) | ( wire18656 ) | ( wire18670 ) | ( wire18671 ) ;
 assign wire18686 = ( n_n156  &  wire719 ) | ( n_n149  &  wire725 ) ;
 assign wire18687 = ( n_n156  &  wire719 ) | ( n_n170  &  wire725 ) ;
 assign wire18688 = ( n_n5144 ) | ( n_n42  &  n_n191  &  wire719 ) ;
 assign wire18691 = ( wire3068 ) | ( wire3080 ) | ( wire3081 ) | ( wire18688 ) ;
 assign wire18692 = ( wire662 ) | ( wire3069 ) | ( wire3078 ) | ( wire3079 ) ;
 assign wire18694 = ( n_n4755 ) | ( wire18631 ) | ( wire18632 ) ;
 assign wire18695 = ( wire18691 ) | ( wire18692 ) | ( wire18694 ) ;
 assign wire18696 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire18701 = ( n_n7240 ) | ( n_n7252 ) | ( wire3060 ) ;
 assign wire18702 = ( n_n7242 ) | ( n_n7254 ) | ( n_n7248 ) | ( wire3059 ) ;
 assign wire18703 = ( i_7_  &  i_6_  &  n_n219  &  n_n111 ) | ( (~ i_7_)  &  i_6_  &  n_n219  &  n_n111 ) ;
 assign wire18704 = ( n_n18  &  n_n48  &  n_n219 ) | ( n_n18  &  n_n219  &  n_n218 ) ;
 assign wire18705 = ( n_n16  &  n_n48  &  n_n219 ) | ( n_n16  &  n_n219  &  n_n218 ) ;
 assign wire18706 = ( wire18703 ) | ( n_n14  &  wire730  &  n_n149 ) ;
 assign wire18707 = ( wire18705 ) | ( wire18704 ) ;
 assign wire18709 = ( wire3044 ) | ( n_n41  &  wire245 ) ;
 assign wire18711 = ( n_n5058 ) | ( wire3550 ) | ( wire3551 ) | ( wire4900 ) ;
 assign wire18712 = ( n_n5055 ) | ( wire18709 ) | ( wire182  &  n_n40 ) ;
 assign wire18714 = ( n_n9  &  n_n74 ) | ( n_n9  &  wire1389 ) | ( n_n10  &  wire1389 ) ;
 assign wire18715 = ( n_n6  &  wire344 ) | ( n_n12  &  wire1390 ) ;
 assign wire18718 = ( wire3066 ) | ( wire3067 ) | ( wire18714 ) | ( wire18715 ) ;
 assign wire18719 = ( n_n3054 ) | ( wire18701 ) | ( wire18702 ) | ( wire18718 ) ;
 assign wire18720 = ( wire729  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign wire18725 = ( wire59 ) | ( wire289 ) | ( wire729  &  n_n170 ) ;
 assign wire18726 = ( n_n1408 ) | ( n_n30  &  wire789 ) ;
 assign wire18731 = ( wire104 ) | ( wire94 ) | ( wire324 ) ;
 assign wire18732 = ( n_n1426 ) | ( n_n30  &  wire791 ) ;
 assign wire18735 = ( n_n1416 ) | ( n_n30  &  wire793 ) ;
 assign wire18736 = ( wire3020 ) | ( wire3032 ) | ( wire18726 ) ;
 assign wire18737 = ( wire3027 ) | ( wire18732 ) | ( wire18735 ) ;
 assign wire18738 = ( n_n184  &  wire729 ) | ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) ;
 assign wire18744 = ( n_n89 ) | ( wire93 ) | ( wire54 ) | ( wire241 ) ;
 assign wire18749 = ( n_n1442 ) | ( wire3008 ) | ( wire3461 ) | ( wire18300 ) ;
 assign wire18750 = ( wire3006 ) | ( n_n31  &  wire863 ) ;
 assign wire18752 = ( n_n199  &  wire729 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire715 ) ;
 assign wire18755 = ( n_n1434 ) | ( wire3001 ) | ( wire3015 ) ;
 assign wire18756 = ( wire18755 ) | ( n_n31  &  wire865 ) ;
 assign wire18757 = ( wire3013 ) | ( wire3014 ) | ( wire18749 ) | ( wire18750 ) ;
 assign wire18760 = ( wire130  &  n_n32 ) | ( n_n33  &  wire48 ) ;
 assign wire18761 = ( n_n2733 ) | ( wire675 ) | ( n_n32  &  wire1417 ) ;
 assign wire18763 = ( n_n101  &  wire381 ) | ( n_n32  &  wire124 ) ;
 assign wire18767 = ( wire3078 ) | ( wire3079 ) | ( wire3080 ) | ( wire3081 ) ;
 assign wire18768 = ( wire587 ) | ( wire564 ) | ( wire566 ) | ( wire670 ) ;
 assign wire18769 = ( wire2985 ) | ( wire18763 ) | ( wire18767 ) ;
 assign wire18770 = ( wire2995 ) | ( wire18760 ) | ( wire18761 ) | ( wire18768 ) ;
 assign wire18771 = ( n_n216  &  wire721 ) | ( n_n199  &  wire725 ) | ( n_n216  &  wire725 ) ;
 assign wire18773 = ( wire729  &  n_n156 ) | ( n_n199  &  wire719 ) ;
 assign wire18776 = ( wire3996 ) | ( n_n31  &  wire172 ) | ( n_n31  &  n_n138 ) ;
 assign wire18777 = ( wire2981 ) | ( n_n30  &  wire1021 ) ;
 assign wire18780 = ( n_n191  &  wire719 ) | ( n_n184  &  wire725 ) ;
 assign wire18783 = ( wire2979 ) | ( n_n31  &  wire1022 ) | ( n_n31  &  wire1263 ) ;
 assign wire18784 = ( n_n156  &  wire721 ) | ( n_n177  &  wire725 ) | ( n_n156  &  wire725 ) ;
 assign wire18786 = ( n_n4240 ) | ( wire2970 ) | ( n_n31  &  wire144 ) ;
 assign wire18788 = ( wire2964 ) | ( wire2974 ) | ( wire2975 ) ;
 assign wire18789 = ( wire2965 ) | ( wire4427 ) | ( wire4428 ) | ( wire18786 ) ;
 assign wire18790 = ( wire18776 ) | ( wire18777 ) | ( wire18788 ) ;
 assign wire18792 = ( n_n5144 ) | ( wire18736 ) | ( wire18737 ) ;
 assign wire18793 = ( wire18756 ) | ( wire18757 ) | ( wire18769 ) | ( wire18770 ) ;
 assign wire18795 = ( wire18682 ) | ( wire18683 ) | ( wire18685 ) | ( wire18793 ) ;
 assign wire18801 = ( wire446 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire18802 = ( wire4354 ) | ( wire4355 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire18803 = ( n_n6271 ) | ( n_n6267 ) | ( n_n6270 ) | ( n_n6269 ) ;
 assign wire18804 = ( n_n5144 ) | ( n_n6266 ) | ( n_n6268 ) | ( n_n6005 ) ;
 assign wire18807 = ( wire419 ) | ( wire445 ) | ( wire18801 ) | ( wire18804 ) ;
 assign wire18809 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire18810 = ( n_n124  &  n_n159  &  n_n111 ) | ( n_n35  &  n_n159  &  n_n111 ) ;
 assign wire18811 = ( n_n124  &  n_n159  &  n_n218 ) | ( n_n35  &  n_n159  &  n_n218 ) ;
 assign wire18812 = ( n_n5319 ) | ( n_n4  &  wire729  &  n_n156 ) ;
 assign wire18814 = ( wire2953 ) | ( wire3550 ) | ( n_n51  &  n_n41 ) ;
 assign wire18815 = ( wire2952 ) | ( wire2958 ) | ( wire2959 ) | ( wire18812 ) ;
 assign wire18816 = ( n_n5319 ) | ( n_n2  &  wire95 ) ;
 assign wire18818 = ( n_n3179 ) | ( wire18814 ) | ( wire18815 ) | ( wire18816 ) ;
 assign wire18821 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire18824 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign wire18826 = ( n_n34  &  n_n133 ) | ( n_n36  &  wire1247 ) | ( n_n34  &  wire1247 ) ;
 assign wire18828 = ( wire2939 ) | ( wire2940 ) | ( wire18826 ) ;
 assign wire18830 = ( wire321 ) | ( n_n184  &  wire721 ) | ( n_n216  &  wire721 ) ;
 assign wire18831 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire18832 = ( wire2937 ) | ( n_n30  &  wire994 ) | ( n_n30  &  wire18830 ) ;
 assign wire18833 = ( n_n159  &  n_n218  &  wire747 ) ;
 assign wire18834 = ( n_n30  &  wire1196 ) | ( n_n31  &  wire1195 ) | ( n_n30  &  wire1195 ) ;
 assign wire18835 = ( wire95 ) | ( wire729  &  n_n191 ) | ( wire729  &  n_n156 ) ;
 assign wire18837 = ( wire551 ) | ( n_n191  &  wire725  &  wire18833 ) ;
 assign wire18838 = ( n_n30  &  n_n129 ) | ( n_n51  &  wire18298 ) ;
 assign wire18839 = ( wire428 ) | ( wire462 ) | ( n_n7264 ) ;
 assign wire18841 = ( wire18837 ) | ( wire18838 ) | ( wire18839 ) ;
 assign wire18845 = ( n_n31  &  wire1285 ) | ( n_n30  &  wire1285 ) | ( n_n31  &  wire321 ) ;
 assign wire18846 = ( n_n1843 ) | ( wire2923 ) | ( wire18841 ) | ( wire18845 ) ;
 assign wire18847 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire721 ) ;
 assign wire18850 = ( n_n41  &  n_n115 ) | ( n_n40  &  n_n115 ) | ( n_n40  &  wire989 ) ;
 assign wire18852 = ( n_n177  &  wire716 ) | ( n_n177  &  wire715 ) ;
 assign wire18854 = ( n_n40  &  n_n129 ) | ( n_n38  &  n_n82 ) ;
 assign wire18855 = ( n_n127  &  wire190 ) | ( n_n166  &  wire334 ) ;
 assign wire18857 = ( wire18854 ) | ( wire18855 ) | ( n_n39  &  wire836 ) ;
 assign wire18858 = ( wire2909 ) | ( wire2910 ) | ( wire2911 ) | ( wire18850 ) ;
 assign wire18859 = ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire18863 = ( wire2897 ) | ( wire190  &  n_n199  &  wire721 ) ;
 assign wire18865 = ( n_n36  &  n_n102 ) | ( n_n38  &  n_n73 ) ;
 assign wire18866 = ( n_n34  &  wire136 ) | ( n_n36  &  wire364 ) ;
 assign wire18871 = ( n_n34  &  n_n95 ) | ( n_n34  &  wire74 ) | ( n_n34  &  wire364 ) ;
 assign wire18872 = ( wire18871 ) | ( n_n34  &  wire143 ) | ( n_n34  &  n_n102 ) ;
 assign wire18874 = ( n_n1870 ) | ( wire18872 ) | ( n_n36  &  wire840 ) ;
 assign wire18877 = ( n_n34  &  wire1579 ) | ( n_n36  &  wire1578 ) | ( n_n34  &  wire1578 ) ;
 assign wire18878 = ( i_15_  &  n_n216  &  n_n201 ) | ( (~ i_15_)  &  n_n149  &  n_n201 ) ;
 assign wire18879 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire729 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire729 ) ;
 assign wire18882 = ( n_n36  &  wire133 ) | ( n_n36  &  wire376 ) | ( n_n36  &  wire18878 ) ;
 assign wire18883 = ( wire2875 ) | ( n_n34  &  wire123 ) | ( n_n34  &  wire133 ) ;
 assign wire18884 = ( wire18877 ) | ( wire18882 ) | ( n_n36  &  wire1580 ) ;
 assign wire18885 = ( n_n36  &  wire313 ) | ( n_n36  &  n_n184  &  wire729 ) ;
 assign wire18889 = ( n_n36  &  wire52 ) | ( n_n34  &  wire52 ) ;
 assign wire18890 = ( wire2866 ) | ( wire2865 ) ;
 assign wire18891 = ( n_n3638 ) | ( wire2870 ) | ( wire18885 ) | ( wire18889 ) ;
 assign wire18892 = ( n_n36  &  wire175 ) | ( n_n36  &  wire729  &  n_n156 ) ;
 assign wire18894 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire18895 = ( n_n36  &  wire147 ) | ( n_n34  &  n_n77 ) ;
 assign wire18897 = ( wire2853 ) | ( n_n34  &  wire911 ) ;
 assign wire18898 = ( wire18895 ) | ( n_n34  &  wire147 ) | ( n_n34  &  wire146 ) ;
 assign wire18901 = ( wire18883 ) | ( wire18884 ) | ( wire18890 ) | ( wire18891 ) ;
 assign wire18908 = ( wire312 ) | ( wire316 ) | ( wire331 ) ;
 assign wire18911 = ( n_n197  &  wire1135 ) | ( n_n212  &  wire1135 ) | ( n_n212  &  wire319 ) ;
 assign wire18912 = ( wire2848 ) | ( wire2849 ) | ( wire2850 ) | ( wire2851 ) ;
 assign wire18913 = ( n_n125  &  n_n117 ) | ( n_n123  &  n_n102 ) ;
 assign wire18914 = ( n_n123  &  wire313 ) | ( n_n125  &  wire383 ) ;
 assign wire18916 = ( n_n125  &  wire52 ) | ( n_n125  &  wire1279 ) | ( n_n123  &  wire1279 ) ;
 assign wire18917 = ( wire18913 ) | ( wire18914 ) | ( n_n123  &  wire52 ) ;
 assign wire18918 = ( wire2842 ) | ( wire2843 ) | ( wire18916 ) ;
 assign wire18919 = ( n_n197  &  n_n139 ) | ( n_n212  &  n_n139 ) | ( n_n212  &  n_n141 ) ;
 assign wire18921 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire18922 = ( wire2831 ) | ( wire18919 ) | ( wire188  &  n_n131 ) ;
 assign wire18923 = ( wire2828 ) | ( n_n212  &  wire1281 ) ;
 assign wire18924 = ( n_n197  &  n_n129 ) | ( n_n212  &  n_n129 ) | ( n_n197  &  n_n127 ) | ( n_n212  &  n_n127 ) ;
 assign wire18925 = ( n_n125  &  n_n102 ) | ( n_n123  &  wire74 ) ;
 assign wire18926 = ( n_n125  &  wire74 ) | ( n_n125  &  wire1136 ) | ( n_n123  &  wire1136 ) ;
 assign wire18928 = ( wire2825 ) | ( wire18924 ) | ( wire18926 ) ;
 assign wire18929 = ( wire2817 ) | ( wire18925 ) | ( wire18928 ) ;
 assign wire18930 = ( wire18917 ) | ( wire18918 ) | ( wire18922 ) | ( wire18923 ) ;
 assign wire18931 = ( n_n125  &  wire376 ) | ( n_n125  &  wire729  &  n_n156 ) ;
 assign wire18932 = ( n_n123  &  wire133 ) | ( n_n123  &  wire904 ) ;
 assign wire18934 = ( n_n125  &  n_n115 ) | ( n_n123  &  n_n115 ) | ( n_n125  &  wire1242 ) ;
 assign wire18935 = ( wire18934 ) | ( n_n71  &  n_n123 ) | ( n_n123  &  wire1242 ) ;
 assign wire18936 = ( wire2808 ) | ( wire2809 ) | ( wire18931 ) | ( wire18932 ) ;
 assign wire18938 = ( n_n113  &  n_n115 ) | ( n_n108  &  n_n107 ) ;
 assign wire18939 = ( wire760 ) | ( wire2797 ) | ( n_n112  &  wire1239 ) ;
 assign wire18941 = ( n_n113  &  n_n122 ) | ( wire255  &  n_n131 ) ;
 assign wire18943 = ( wire2791 ) | ( wire2801 ) | ( wire2802 ) | ( wire18941 ) ;
 assign wire18944 = ( i_15_  &  n_n213  &  n_n177 ) | ( (~ i_15_)  &  n_n213  &  n_n177 ) | ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) ;
 assign wire18945 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire729 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire729 ) ;
 assign wire18947 = ( n_n125  &  wire147 ) | ( n_n123  &  n_n77 ) ;
 assign wire18949 = ( wire2814 ) | ( wire2815 ) | ( wire18947 ) ;
 assign wire18950 = ( wire2784 ) | ( wire2785 ) | ( wire18949 ) ;
 assign wire18951 = ( n_n1913 ) | ( wire18935 ) | ( wire18936 ) | ( wire18943 ) ;
 assign wire18955 = ( n_n101  &  n_n115 ) | ( n_n108  &  n_n115 ) | ( n_n101  &  wire1470 ) ;
 assign wire18956 = ( n_n216  &  wire721 ) | ( n_n149  &  wire715 ) ;
 assign wire18958 = ( n_n216  &  wire721 ) | ( n_n156  &  wire715 ) ;
 assign wire18959 = ( wire729  &  n_n156 ) | ( wire717  &  n_n156 ) | ( wire729  &  n_n149 ) | ( wire717  &  n_n149 ) ;
 assign wire18961 = ( wire2775 ) | ( wire228  &  n_n199  &  wire721 ) ;
 assign wire18962 = ( wire2776 ) | ( wire18955 ) | ( n_n108  &  wire1469 ) ;
 assign wire18965 = ( n_n101  &  n_n129 ) | ( n_n101  &  n_n127 ) | ( n_n108  &  n_n127 ) ;
 assign wire18966 = ( wire18965 ) | ( wire1200  &  wire1199 ) ;
 assign wire18968 = ( n_n42  &  wire257 ) | ( n_n43  &  wire313 ) ;
 assign wire18969 = ( n_n43  &  wire139 ) | ( n_n42  &  n_n117 ) | ( n_n43  &  n_n117 ) ;
 assign wire18970 = ( n_n47  &  n_n129 ) | ( n_n43  &  n_n89 ) ;
 assign wire18971 = ( n_n46  &  wire1754 ) | ( n_n46  &  wire1753 ) | ( n_n47  &  wire1753 ) ;
 assign wire18972 = ( n_n43  &  wire257 ) | ( n_n42  &  wire313 ) ;
 assign wire18973 = ( wire52  &  n_n43 ) | ( n_n42  &  wire139 ) ;
 assign wire18975 = ( wire18973 ) | ( wire18972 ) ;
 assign wire18976 = ( wire18968 ) | ( wire18969 ) | ( wire18970 ) | ( wire18971 ) ;
 assign wire18978 = ( i_9_  &  i_10_  &  i_11_  &  wire721 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire721 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire721 ) ;
 assign wire18980 = ( wire303 ) | ( wire321 ) | ( wire410 ) ;
 assign wire18981 = ( n_n139  &  wire189 ) | ( n_n47  &  wire1766 ) ;
 assign wire18985 = ( wire2750 ) | ( wire2751 ) | ( wire18975 ) | ( wire18976 ) ;
 assign wire18986 = ( wire729  &  n_n177 ) | ( n_n177  &  wire717 ) | ( n_n177  &  wire715 ) ;
 assign wire18991 = ( wire2748 ) | ( n_n101  &  wire1194 ) | ( n_n101  &  wire1497 ) ;
 assign wire18992 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire715 ) ;
 assign wire18993 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire715 ) ;
 assign wire18997 = ( wire305 ) | ( wire380 ) | ( n_n177  &  wire715 ) ;
 assign wire18998 = ( wire2740 ) | ( wire2743 ) | ( wire2744 ) ;
 assign wire19001 = ( n_n199  &  wire729 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire715 ) ;
 assign wire19003 = ( wire2733 ) | ( wire2738 ) | ( wire2739 ) ;
 assign wire19004 = ( wire19003 ) | ( n_n108  &  wire1205 ) ;
 assign wire19005 = ( wire2741 ) | ( wire2746 ) | ( wire18991 ) | ( wire18998 ) ;
 assign wire19006 = ( n_n177  &  wire717 ) | ( n_n177  &  wire715 ) ;
 assign wire19008 = ( n_n184  &  wire729 ) | ( n_n184  &  wire717 ) | ( n_n184  &  wire715 ) ;
 assign wire19009 = ( wire2724 ) | ( n_n40  &  wire261 ) | ( n_n40  &  wire375 ) ;
 assign wire19010 = ( wire2726 ) | ( wire2728 ) | ( wire2729 ) ;
 assign wire19011 = ( n_n42  &  n_n89 ) | ( n_n41  &  n_n107 ) ;
 assign wire19013 = ( n_n199  &  wire729 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire715 ) ;
 assign wire19015 = ( wire2717 ) | ( wire2720 ) | ( wire2721 ) | ( wire19011 ) ;
 assign wire19016 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire715 ) | ( i_9_  &  i_10_  &  (~ i_11_)  &  wire715 ) ;
 assign wire19020 = ( wire352 ) | ( wire380 ) | ( n_n177  &  wire715 ) ;
 assign wire19021 = ( n_n6445 ) | ( wire2712 ) | ( wire2730 ) | ( wire2731 ) ;
 assign wire19023 = ( wire2718 ) | ( wire19009 ) | ( wire19010 ) | ( wire19015 ) ;
 assign wire19025 = ( wire18911 ) | ( wire18912 ) | ( wire18929 ) | ( wire18930 ) ;
 assign wire19027 = ( n_n1824 ) | ( wire18985 ) | ( wire19004 ) | ( wire19005 ) ;
 assign wire19029 = ( n_n1803 ) | ( wire18950 ) | ( wire18951 ) | ( wire19025 ) ;
 assign wire19030 = ( n_n1800 ) | ( n_n1799 ) | ( n_n1801 ) | ( wire19027 ) ;
 assign wire19031 = ( wire708 ) | ( wire473 ) | ( wire2914 ) | ( wire2915 ) ;
 assign wire19033 = ( wire2704 ) | ( wire2705 ) | ( wire19031 ) ;
 assign wire19034 = ( n_n1811 ) | ( wire2943 ) | ( wire2944 ) | ( wire18828 ) ;
 assign wire19036 = ( n_n1809 ) | ( wire18846 ) | ( wire19033 ) | ( wire19034 ) ;
 assign wire19038 = ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire19043 = ( n_n71 ) | ( wire155 ) | ( wire49 ) | ( wire92 ) ;
 assign wire19044 = ( wire2702 ) | ( wire2703 ) | ( n_n36  &  wire845 ) ;
 assign wire19047 = ( wire155 ) | ( wire315 ) | ( wire300 ) ;
 assign wire19048 = ( n_n71  &  n_n36 ) | ( n_n34  &  wire133 ) ;
 assign wire19050 = ( wire542 ) | ( wire2692 ) | ( wire19048 ) ;
 assign wire19053 = ( wire118 ) | ( wire277 ) | ( wire729  &  n_n170 ) ;
 assign wire19054 = ( n_n36  &  wire850 ) | ( n_n34  &  wire849 ) ;
 assign wire19055 = ( wire2691 ) | ( wire19054 ) | ( n_n34  &  wire1207 ) ;
 assign wire19057 = ( wire2693 ) | ( wire2700 ) | ( wire19044 ) | ( wire19050 ) ;
 assign wire19062 = ( wire397 ) | ( n_n3417 ) | ( n_n1553 ) ;
 assign wire19063 = ( wire2679 ) | ( n_n41  &  wire1152 ) ;
 assign wire19069 = ( n_n3419 ) | ( wire500 ) | ( n_n40  &  wire1153 ) ;
 assign wire19071 = ( wire239 ) | ( wire223 ) ;
 assign wire19072 = ( wire148 ) | ( wire179 ) | ( wire274 ) ;
 assign wire19074 = ( wire518 ) | ( n_n3415 ) | ( wire2669 ) ;
 assign wire19075 = ( wire19074 ) | ( n_n40  &  wire19071 ) | ( n_n40  &  wire19072 ) ;
 assign wire19076 = ( wire2676 ) | ( wire19062 ) | ( wire19063 ) | ( wire19069 ) ;
 assign wire19077 = ( n_n42  &  n_n89 ) | ( n_n43  &  wire65 ) ;
 assign wire19078 = ( n_n41  &  n_n107 ) | ( n_n41  &  n_n202 ) | ( n_n41  &  n_n214 ) ;
 assign wire19079 = ( n_n42  &  n_n115 ) | ( n_n42  &  n_n136 ) | ( n_n43  &  n_n136 ) ;
 assign wire19083 = ( n_n4622 ) | ( n_n3421 ) | ( n_n1566 ) | ( wire2657 ) ;
 assign wire19084 = ( wire2666 ) | ( wire19077 ) | ( wire19078 ) | ( wire19079 ) ;
 assign wire19087 = ( n_n42  &  wire139 ) | ( n_n43  &  n_n89 ) ;
 assign wire19089 = ( wire19087 ) | ( n_n42  &  wire54 ) | ( n_n42  &  wire357 ) ;
 assign wire19090 = ( n_n4808 ) | ( n_n1575 ) | ( n_n43  &  wire1297 ) ;
 assign wire19094 = ( wire142 ) | ( wire56 ) | ( wire233 ) ;
 assign wire19097 = ( n_n4620 ) | ( n_n6384 ) | ( wire2645 ) | ( wire2646 ) ;
 assign wire19098 = ( wire19083 ) | ( wire19084 ) | ( wire19089 ) | ( wire19090 ) ;
 assign wire19099 = ( wire717  &  n_n156 ) | ( n_n156  &  wire727 ) ;
 assign wire19103 = ( n_n6267 ) | ( n_n47  &  wire1499 ) ;
 assign wire19104 = ( n_n191  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire19106 = ( n_n6269 ) | ( wire4252 ) | ( wire4253 ) ;
 assign wire19108 = ( wire2636 ) | ( n_n46  &  wire72 ) | ( n_n46  &  wire19104 ) ;
 assign wire19109 = ( wire2638 ) | ( wire2643 ) | ( wire19103 ) | ( wire19106 ) ;
 assign wire19110 = ( wire717  &  n_n156 ) | ( n_n199  &  wire721 ) ;
 assign wire19113 = ( n_n191  &  wire728 ) | ( n_n156  &  wire727 ) ;
 assign wire19116 = ( wire175 ) | ( wire88 ) | ( wire198 ) ;
 assign wire19118 = ( n_n1594 ) | ( wire2630 ) | ( wire2634 ) | ( wire2635 ) ;
 assign wire19119 = ( wire726  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire19123 = ( n_n46  &  wire852 ) | ( n_n47  &  wire1436 ) ;
 assign wire19125 = ( wire2631 ) | ( wire19108 ) | ( wire19109 ) | ( wire19118 ) ;
 assign wire19126 = ( n_n5109 ) | ( wire677 ) | ( wire19123 ) | ( wire19125 ) ;
 assign wire19127 = ( wire19075 ) | ( wire19076 ) | ( wire19097 ) | ( wire19098 ) ;
 assign wire19128 = ( (~ i_15_)  &  n_n191  &  n_n201 ) | ( i_15_  &  n_n149  &  n_n201 ) ;
 assign wire19129 = ( n_n170  &  wire721 ) | ( n_n191  &  wire728 ) | ( n_n170  &  wire728 ) ;
 assign wire19130 = ( n_n33  &  n_n52 ) | ( n_n136  &  n_n32 ) ;
 assign wire19134 = ( wire473 ) | ( wire2615 ) | ( wire2618 ) | ( wire19130 ) ;
 assign wire19138 = ( n_n33  &  wire133 ) | ( n_n33  &  wire60 ) | ( n_n33  &  wire127 ) ;
 assign wire19144 = ( wire63 ) | ( wire330 ) | ( n_n199  &  wire720 ) ;
 assign wire19146 = ( n_n1434 ) | ( wire2606 ) | ( n_n30  &  wire925 ) ;
 assign wire19147 = ( n_n1442 ) | ( n_n1170 ) | ( wire2614 ) | ( wire19134 ) ;
 assign wire19148 = ( n_n125  &  wire1287 ) | ( n_n123  &  wire1286 ) ;
 assign wire19150 = ( n_n184  &  wire729 ) | ( n_n184  &  wire728 ) ;
 assign wire19152 = ( wire2598 ) | ( n_n112  &  wire63 ) ;
 assign wire19153 = ( wire2599 ) | ( wire19148 ) | ( n_n113  &  wire276 ) ;
 assign wire19158 = ( n_n1700 ) | ( wire2594 ) | ( n_n123  &  wire133 ) ;
 assign wire19163 = ( wire2588 ) | ( n_n71  &  n_n125 ) | ( n_n125  &  wire155 ) ;
 assign wire19164 = ( n_n2881 ) | ( n_n1708 ) | ( n_n123  &  wire916 ) ;
 assign wire19168 = ( wire98 ) | ( wire63 ) | ( wire254 ) ;
 assign wire19169 = ( n_n123  &  wire52 ) | ( n_n125  &  n_n117 ) ;
 assign wire19170 = ( wire2584 ) | ( wire19169 ) ;
 assign wire19174 = ( wire53 ) | ( wire126 ) | ( wire239 ) ;
 assign wire19177 = ( n_n1717 ) | ( wire639 ) | ( wire2578 ) | ( wire2579 ) ;
 assign wire19178 = ( wire2585 ) | ( wire19163 ) | ( wire19164 ) | ( wire19170 ) ;
 assign wire19179 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( n_n191  &  wire717 ) ;
 assign wire19182 = ( n_n184  &  wire729 ) | ( n_n191  &  wire727 ) ;
 assign wire19185 = ( wire257 ) | ( wire271 ) | ( wire19182 ) ;
 assign wire19186 = ( n_n5019 ) | ( n_n108  &  wire1070 ) ;
 assign wire19189 = ( n_n113  &  n_n115 ) | ( n_n108  &  wire111 ) ;
 assign wire19190 = ( wire760 ) | ( wire2567 ) | ( n_n112  &  wire65 ) ;
 assign wire19192 = ( wire19190 ) | ( n_n108  &  wire143 ) | ( n_n108  &  wire154 ) ;
 assign wire19193 = ( n_n5033 ) | ( wire2568 ) | ( wire19189 ) ;
 assign wire19194 = ( i_15_  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n213  &  n_n191 ) | ( (~ i_15_)  &  n_n191  &  n_n209 ) ;
 assign wire19196 = ( n_n199  &  wire729 ) | ( n_n199  &  wire727 ) ;
 assign wire19197 = ( n_n199  &  wire720 ) | ( n_n199  &  wire717 ) | ( n_n199  &  wire715 ) ;
 assign wire19200 = ( n_n5021 ) | ( wire2560 ) | ( wire2565 ) ;
 assign wire19201 = ( wire19200 ) | ( n_n108  &  wire1075 ) ;
 assign wire19202 = ( wire2576 ) | ( wire19186 ) | ( wire19192 ) | ( wire19193 ) ;
 assign wire19204 = ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) | ( n_n177  &  wire728 ) ;
 assign wire19208 = ( wire2556 ) | ( wire2557 ) | ( wire2558 ) | ( wire2559 ) ;
 assign wire19210 = ( wire2595 ) | ( wire19152 ) | ( wire19153 ) | ( wire19158 ) ;
 assign wire19211 = ( wire2548 ) | ( wire2549 ) | ( wire19208 ) | ( wire19210 ) ;
 assign wire19212 = ( wire19177 ) | ( wire19178 ) | ( wire19201 ) | ( wire19202 ) ;
 assign wire19213 = ( n_n212  &  n_n127 ) | ( n_n197  &  wire83 ) ;
 assign wire19216 = ( wire729  &  n_n216 ) | ( n_n184  &  wire720 ) ;
 assign wire19219 = ( wire142 ) | ( wire251 ) | ( wire19216 ) ;
 assign wire19220 = ( n_n212  &  wire63 ) | ( n_n212  &  wire1145 ) ;
 assign wire19221 = ( n_n184  &  wire729 ) | ( n_n177  &  wire720 ) ;
 assign wire19226 = ( wire98 ) | ( wire51 ) | ( wire254 ) ;
 assign wire19227 = ( n_n197  &  wire52 ) | ( n_n212  &  wire1147 ) ;
 assign wire19232 = ( wire2532 ) | ( n_n212  &  wire1150 ) ;
 assign wire19233 = ( wire2537 ) | ( wire19232 ) | ( n_n197  &  wire70 ) ;
 assign wire19234 = ( wire2540 ) | ( wire2543 ) | ( wire19220 ) | ( wire19227 ) ;
 assign wire19238 = ( n_n123  &  n_n102 ) | ( n_n125  &  wire51 ) ;
 assign wire19239 = ( n_n125  &  wire52 ) | ( n_n123  &  wire142 ) ;
 assign wire19240 = ( wire19239 ) | ( wire19238 ) ;
 assign wire19241 = ( wire2526 ) | ( n_n125  &  wire1255 ) ;
 assign wire19243 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) ;
 assign wire19245 = ( n_n216  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire19246 = ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire19248 = ( wire2518 ) | ( n_n197  &  wire1257 ) ;
 assign wire19249 = ( wire2522 ) | ( wire2523 ) | ( wire2524 ) | ( wire2525 ) ;
 assign wire19250 = ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) | ( wire729  &  n_n156 ) ;
 assign wire19253 = ( n_n177  &  wire720 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire19256 = ( n_n197  &  wire127 ) | ( n_n212  &  wire1289 ) ;
 assign wire19258 = ( wire221 ) | ( wire315 ) ;
 assign wire19259 = ( wire49 ) | ( wire300 ) | ( wire720  &  n_n149 ) ;
 assign wire19260 = ( wire729  &  n_n156 ) | ( wire729  &  n_n149 ) | ( wire726  &  n_n149 ) ;
 assign wire19263 = ( n_n4388 ) | ( n_n212  &  wire19258 ) | ( n_n212  &  wire19259 ) ;
 assign wire19268 = ( n_n212  &  wire147 ) | ( n_n212  &  wire126 ) | ( n_n212  &  wire1293 ) ;
 assign wire19269 = ( wire19268 ) | ( n_n197  &  wire1294 ) ;
 assign wire19270 = ( wire2513 ) | ( wire2516 ) | ( wire19256 ) | ( wire19263 ) ;
 assign wire19272 = ( n_n123  &  wire68 ) | ( n_n123  &  wire81 ) | ( n_n123  &  wire74 ) ;
 assign wire19273 = ( n_n4674 ) | ( wire2498 ) | ( n_n125  &  n_n102 ) ;
 assign wire19274 = ( wire2545 ) | ( wire19213 ) | ( wire19272 ) ;
 assign wire19276 = ( wire19240 ) | ( wire19241 ) | ( wire19248 ) | ( wire19249 ) ;
 assign wire19277 = ( wire19273 ) | ( wire19274 ) | ( wire19276 ) ;
 assign wire19278 = ( wire19233 ) | ( wire19234 ) | ( wire19269 ) | ( wire19270 ) ;
 assign wire19279 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) ;
 assign wire19281 = ( n_n170  &  wire717 ) | ( n_n170  &  wire727 ) ;
 assign wire19283 = ( wire19281 ) | ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) ;
 assign wire19284 = ( wire59 ) | ( wire69 ) | ( wire281 ) ;
 assign wire19285 = ( wire685 ) | ( n_n101  &  wire250 ) ;
 assign wire19286 = ( wire2493 ) | ( n_n108  &  wire19283 ) | ( n_n108  &  wire19284 ) ;
 assign wire19289 = ( wire156 ) | ( wire59 ) | ( wire300 ) ;
 assign wire19290 = ( wire729  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire19291 = ( wire726  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire19294 = ( n_n5000 ) | ( wire2490 ) | ( n_n108  &  wire234 ) ;
 assign wire19295 = ( wire729  &  n_n191 ) | ( wire726  &  n_n191 ) | ( n_n191  &  wire717 ) ;
 assign wire19297 = ( wire729  &  n_n177 ) | ( wire726  &  n_n177 ) ;
 assign wire19299 = ( n_n5011 ) | ( wire2481 ) | ( n_n108  &  wire250 ) ;
 assign wire19301 = ( wire2480 ) | ( wire2487 ) | ( wire2488 ) | ( wire19299 ) ;
 assign wire19302 = ( wire2489 ) | ( wire19285 ) | ( wire19286 ) | ( wire19294 ) ;
 assign wire19304 = ( n_n6005 ) | ( wire419 ) | ( n_n101  &  n_n129 ) ;
 assign wire19306 = ( wire729  &  n_n216 ) | ( wire726  &  n_n216 ) | ( n_n216  &  wire717 ) ;
 assign wire19307 = ( n_n108  &  n_n129 ) | ( n_n101  &  wire378 ) ;
 assign wire19308 = ( n_n46  &  wire1343 ) | ( wire1345  &  wire1342 ) ;
 assign wire19309 = ( wire19307 ) | ( n_n47  &  wire162 ) | ( n_n47  &  wire19306 ) ;
 assign wire19310 = ( n_n1624 ) | ( wire2475 ) | ( wire19304 ) | ( wire19308 ) ;
 assign wire19312 = ( n_n184  &  wire721 ) | ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire19315 = ( n_n191  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire19316 = ( wire2464 ) | ( n_n101  &  wire90 ) ;
 assign wire19317 = ( wire2463 ) | ( wire2468 ) | ( n_n101  &  wire1405 ) ;
 assign wire19318 = ( n_n199  &  wire729 ) | ( n_n199  &  wire717 ) ;
 assign wire19320 = ( n_n216  &  wire717 ) | ( n_n216  &  wire715 ) ;
 assign wire19324 = ( wire2462 ) | ( n_n46  &  wire1214 ) | ( n_n46  &  wire1581 ) ;
 assign wire19325 = ( n_n4641 ) | ( wire693 ) | ( wire19324 ) ;
 assign wire19326 = ( wire19309 ) | ( wire19310 ) | ( wire19316 ) | ( wire19317 ) ;
 assign wire19328 = ( i_15_  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n213  &  n_n170 ) | ( (~ i_15_)  &  n_n170  &  n_n209 ) ;
 assign wire19332 = ( n_n5113 ) | ( n_n1606 ) | ( wire2451 ) ;
 assign wire19337 = ( n_n183 ) | ( wire184 ) | ( wire210 ) | ( wire246 ) ;
 assign wire19338 = ( wire2448 ) | ( wire498 ) ;
 assign wire19339 = ( wire729  &  n_n170 ) | ( wire726  &  n_n170 ) | ( n_n170  &  wire717 ) ;
 assign wire19343 = ( n_n5111 ) | ( wire137  &  n_n46 ) | ( n_n46  &  wire146 ) ;
 assign wire19344 = ( wire2442 ) | ( n_n47  &  wire1216 ) ;
 assign wire19346 = ( wire2449 ) | ( wire2452 ) | ( wire19332 ) | ( wire19338 ) ;
 assign wire19347 = ( wire19301 ) | ( wire19302 ) | ( wire19325 ) | ( wire19326 ) ;
 assign wire19348 = ( wire19343 ) | ( wire19344 ) | ( wire19346 ) | ( wire19347 ) ;
 assign wire19349 = ( wire19211 ) | ( wire19212 ) | ( wire19277 ) | ( wire19278 ) ;
 assign wire19351 = ( n_n34  &  wire81 ) | ( n_n36  &  n_n102 ) ;
 assign wire19354 = ( n_n4591 ) | ( n_n1514 ) | ( wire17541 ) | ( wire17542 ) ;
 assign wire19355 = ( wire2435 ) | ( wire19351 ) | ( n_n38  &  wire248 ) ;
 assign wire19359 = ( n_n39  &  wire248 ) | ( n_n39  &  wire249 ) ;
 assign wire19362 = ( n_n1517 ) | ( wire457 ) | ( wire19359 ) ;
 assign wire19363 = ( n_n1520 ) | ( wire572 ) | ( wire2427 ) | ( wire2428 ) ;
 assign wire19364 = ( n_n36  &  wire98 ) | ( n_n34  &  n_n102 ) ;
 assign wire19366 = ( n_n36  &  n_n198 ) | ( n_n34  &  wire74 ) ;
 assign wire19368 = ( wire2418 ) | ( wire2424 ) | ( wire19364 ) ;
 assign wire19369 = ( wire2417 ) | ( wire19366 ) | ( wire19368 ) ;
 assign wire19370 = ( wire19354 ) | ( wire19355 ) | ( wire19362 ) | ( wire19363 ) ;
 assign wire19375 = ( wire52 ) | ( wire51 ) | ( wire271 ) ;
 assign wire19376 = ( n_n1426 ) | ( n_n30  &  wire913 ) ;
 assign wire19380 = ( n_n1416 ) | ( n_n31  &  wire147 ) | ( n_n31  &  wire126 ) ;
 assign wire19381 = ( wire2410 ) | ( n_n30  &  wire1069 ) ;
 assign wire19387 = ( wire52 ) | ( wire63 ) | ( wire51 ) | ( wire148 ) ;
 assign wire19388 = ( wire2407 ) | ( n_n31  &  wire1006 ) ;
 assign wire19389 = ( wire2415 ) | ( wire19376 ) | ( wire19380 ) | ( wire19381 ) ;
 assign wire19393 = ( n_n36  &  n_n176 ) | ( n_n36  &  n_n184  &  wire729 ) ;
 assign wire19395 = ( wire19393 ) | ( n_n34  &  wire52 ) | ( n_n34  &  wire63 ) ;
 assign wire19396 = ( wire2398 ) | ( n_n34  &  wire1077 ) ;
 assign wire19400 = ( n_n36  &  wire52 ) | ( n_n34  &  n_n183 ) ;
 assign wire19401 = ( wire19400 ) | ( n_n36  &  wire63 ) ;
 assign wire19402 = ( wire2393 ) | ( n_n36  &  wire1079 ) ;
 assign wire19403 = ( n_n34  &  n_n77 ) | ( n_n34  &  n_n177  &  wire720 ) ;
 assign wire19405 = ( n_n36  &  wire53 ) | ( n_n36  &  wire126 ) | ( n_n36  &  wire69 ) ;
 assign wire19406 = ( wire2384 ) | ( wire19403 ) | ( n_n36  &  wire147 ) ;
 assign wire19408 = ( wire2404 ) | ( wire2405 ) | ( wire19405 ) | ( wire19406 ) ;
 assign wire19409 = ( wire19395 ) | ( wire19396 ) | ( wire19401 ) | ( wire19402 ) ;
 assign wire19411 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire19412 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire19413 = ( i_15_  &  n_n184  &  n_n201 ) | ( (~ i_15_)  &  n_n156  &  n_n201 ) ;
 assign wire19414 = ( n_n216  &  wire721 ) | ( n_n184  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire19417 = ( wire2379 ) | ( wire2382 ) | ( n_n41  &  wire315 ) ;
 assign wire19420 = ( wire155 ) | ( wire50 ) | ( wire300 ) ;
 assign wire19423 = ( n_n6492 ) | ( n_n3413 ) | ( n_n1542 ) | ( wire2374 ) ;
 assign wire19424 = ( n_n177  &  wire721 ) | ( n_n156  &  wire721 ) | ( n_n156  &  wire728 ) ;
 assign wire19426 = ( wire716  &  n_n170 ) | ( n_n170  &  wire727 ) ;
 assign wire19427 = ( n_n177  &  wire716 ) | ( n_n170  &  wire720 ) ;
 assign wire19429 = ( wire2370 ) | ( wire2371 ) | ( wire2372 ) | ( wire2373 ) ;
 assign wire19430 = ( wire2364 ) | ( wire2365 ) | ( wire19429 ) ;
 assign wire19431 = ( wire2375 ) | ( wire2380 ) | ( wire19417 ) | ( wire19423 ) ;
 assign wire19436 = ( wire315 ) | ( wire300 ) | ( wire720  &  n_n149 ) ;
 assign wire19437 = ( n_n1408 ) | ( n_n30  &  wire1504 ) ;
 assign wire19438 = ( n_n184  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n191  &  wire728 ) ;
 assign wire19440 = ( n_n199  &  wire721 ) | ( n_n199  &  wire728 ) ;
 assign wire19441 = ( n_n216  &  wire721 ) | ( n_n191  &  wire721 ) | ( n_n216  &  wire728 ) | ( n_n191  &  wire728 ) ;
 assign wire19442 = ( wire729  &  n_n156 ) | ( n_n184  &  wire728 ) ;
 assign wire19443 = ( n_n199  &  wire721 ) | ( n_n216  &  wire721 ) | ( n_n199  &  wire728 ) | ( n_n216  &  wire728 ) ;
 assign wire19446 = ( wire2356 ) | ( wire2359 ) | ( n_n31  &  wire1537 ) ;
 assign wire19447 = ( n_n177  &  wire721 ) | ( n_n177  &  wire728 ) ;
 assign wire19448 = ( n_n156  &  wire721 ) | ( n_n149  &  wire721 ) | ( n_n156  &  wire728 ) | ( n_n149  &  wire728 ) ;
 assign wire19449 = ( n_n149  &  wire721 ) | ( n_n149  &  wire728 ) ;
 assign wire19450 = ( n_n170  &  wire721 ) | ( n_n156  &  wire721 ) | ( n_n170  &  wire728 ) | ( n_n156  &  wire728 ) ;
 assign wire19452 = ( wire2352 ) | ( wire2353 ) | ( wire2362 ) | ( wire19437 ) ;
 assign wire19453 = ( n_n5144 ) | ( wire2686 ) | ( wire19055 ) | ( wire19057 ) ;
 assign wire19454 = ( wire19146 ) | ( wire19147 ) | ( wire19369 ) | ( wire19370 ) ;
 assign wire19455 = ( wire19388 ) | ( wire19389 ) | ( wire19408 ) | ( wire19409 ) ;
 assign wire19456 = ( n_n1163 ) | ( wire19430 ) | ( wire19431 ) | ( wire19452 ) ;
 assign wire19458 = ( wire19456 ) | ( wire19455 ) ;
 assign wire19459 = ( wire19126 ) | ( wire19127 ) | ( wire19453 ) | ( wire19454 ) ;
 assign wire19461 = ( wire724  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire715 ) ;
 assign wire19464 = ( wire724  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire19466 = ( wire2345 ) | ( wire2349 ) | ( n_n31  &  wire1012 ) ;
 assign wire19469 = ( n_n184  &  wire724 ) | ( n_n184  &  wire720 ) | ( n_n184  &  wire715 ) ;
 assign wire19471 = ( wire2340 ) | ( wire2343 ) | ( wire2344 ) ;
 assign wire19472 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire724 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign wire19476 = ( wire53 ) | ( wire237 ) | ( wire724  &  n_n177 ) ;
 assign wire19477 = ( wire2335 ) | ( wire2350 ) | ( wire2351 ) ;
 assign wire19479 = ( wire2341 ) | ( wire2346 ) | ( wire19466 ) | ( wire19471 ) ;
 assign wire19480 = ( n_n33  &  n_n191  &  wire719 ) | ( n_n33  &  n_n149  &  wire719 ) ;
 assign wire19481 = ( n_n33  &  n_n132 ) | ( n_n31  &  wire111 ) ;
 assign wire19485 = ( n_n36  &  wire1708 ) | ( n_n36  &  wire1707 ) | ( n_n34  &  wire1707 ) ;
 assign wire19486 = ( wire720  &  n_n149 ) | ( n_n216  &  wire719 ) ;
 assign wire19490 = ( wire438 ) | ( wire215 ) | ( wire720  &  n_n156 ) ;
 assign wire19491 = ( wire2323 ) | ( wire19485 ) | ( n_n34  &  wire1709 ) ;
 assign wire19494 = ( n_n34  &  n_n177  &  wire719 ) | ( n_n34  &  n_n156  &  wire719 ) ;
 assign wire19496 = ( n_n33  &  wire48 ) | ( n_n32  &  wire124 ) ;
 assign wire19497 = ( wire226  &  n_n128 ) | ( n_n32  &  wire165 ) ;
 assign wire19498 = ( wire19494 ) | ( wire19496 ) | ( n_n36  &  wire1738 ) ;
 assign wire19499 = ( wire19497 ) | ( n_n33  &  wire1739 ) ;
 assign wire19500 = ( n_n199  &  wire724 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire715 ) ;
 assign wire19504 = ( wire2324 ) | ( wire19491 ) | ( wire19498 ) | ( wire19499 ) ;
 assign wire19506 = ( n_n212  &  wire46 ) | ( n_n212  &  wire1346 ) ;
 assign wire19510 = ( wire132  &  n_n197 ) | ( wire132  &  n_n212 ) | ( n_n197  &  wire46 ) ;
 assign wire19513 = ( n_n212  &  wire151 ) | ( n_n212  &  wire48 ) ;
 assign wire19516 = ( wire629 ) | ( wire2295 ) | ( wire2296 ) | ( wire19513 ) ;
 assign wire19519 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire19520 = ( n_n36  &  wire219 ) | ( n_n36  &  n_n199  &  wire720 ) ;
 assign wire19521 = ( n_n36  &  wire100 ) | ( n_n36  &  n_n177  &  wire720 ) ;
 assign wire19523 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire19526 = ( wire2283 ) | ( n_n34  &  n_n184  &  wire720 ) ;
 assign wire19527 = ( wire2287 ) | ( wire19521 ) | ( n_n36  &  wire1605 ) ;
 assign wire19528 = ( n_n177  &  wire716 ) | ( wire720  &  n_n149 ) ;
 assign wire19529 = ( i_15_  &  n_n207  &  n_n156 ) | ( (~ i_15_)  &  n_n207  &  n_n156 ) | ( i_15_  &  n_n156  &  n_n215 ) ;
 assign wire19530 = ( i_15_  &  n_n207  &  n_n170 ) | ( (~ i_15_)  &  n_n207  &  n_n170 ) | ( i_15_  &  n_n170  &  n_n215 ) ;
 assign wire19531 = ( i_15_  &  n_n207  &  n_n177 ) | ( (~ i_15_)  &  n_n207  &  n_n177 ) ;
 assign wire19532 = ( wire2281 ) | ( wire2282 ) | ( n_n34  &  n_n176 ) ;
 assign wire19533 = ( wire2278 ) | ( wire2277 ) ;
 assign wire19535 = ( i_15_  &  n_n216  &  n_n207 ) | ( (~ i_15_)  &  n_n216  &  n_n207 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire19536 = ( n_n38  &  n_n134 ) | ( n_n39  &  n_n132 ) ;
 assign wire19538 = ( wire2269 ) | ( wire19536 ) | ( n_n34  &  n_n198 ) ;
 assign wire19539 = ( wire2290 ) | ( wire2293 ) | ( wire2294 ) | ( wire19520 ) ;
 assign wire19541 = ( wire19526 ) | ( wire19527 ) | ( wire19532 ) | ( wire19533 ) ;
 assign wire19542 = ( n_n41  &  n_n130 ) | ( n_n39  &  wire104 ) ;
 assign wire19543 = ( n_n40  &  wire1160 ) | ( n_n41  &  wire1159 ) | ( n_n40  &  wire1159 ) ;
 assign wire19544 = ( n_n138  &  n_n40 ) | ( n_n41  &  n_n142 ) ;
 assign wire19545 = ( n_n41  &  n_n140 ) | ( n_n40  &  n_n140 ) | ( n_n40  &  wire407 ) ;
 assign wire19548 = ( n_n4602 ) | ( wire19542 ) | ( wire19543 ) | ( wire19544 ) ;
 assign wire19549 = ( wire2257 ) | ( wire4863 ) | ( wire4864 ) | ( wire19545 ) ;
 assign wire19552 = ( n_n38  &  wire110 ) | ( n_n38  &  n_n177  &  wire719 ) ;
 assign wire19556 = ( wire635 ) | ( wire19552 ) | ( n_n39  &  wire1633 ) ;
 assign wire19557 = ( n_n969 ) | ( n_n4600 ) | ( n_n972 ) | ( wire2245 ) ;
 assign wire19560 = ( n_n765 ) | ( wire19548 ) | ( wire19549 ) ;
 assign wire19565 = ( wire48 ) | ( wire167 ) | ( wire192 ) ;
 assign wire19567 = ( n_n42  &  n_n138 ) | ( n_n41  &  n_n210 ) ;
 assign wire19569 = ( wire391 ) | ( wire19567 ) | ( n_n116  &  wire1658 ) ;
 assign wire19574 = ( wire2229 ) | ( n_n41  &  wire1659 ) ;
 assign wire19576 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19577 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19580 = ( n_n46  &  n_n140 ) | ( n_n47  &  n_n140 ) | ( n_n47  &  n_n142 ) ;
 assign wire19581 = ( n_n47  &  wire55 ) | ( n_n46  &  wire134 ) ;
 assign wire19582 = ( wire19580 ) | ( n_n47  &  wire163 ) | ( n_n47  &  wire19576 ) ;
 assign wire19583 = ( wire19581 ) | ( n_n46  &  wire1674 ) ;
 assign wire19584 = ( n_n6271 ) | ( n_n6270 ) | ( n_n42  &  n_n183 ) ;
 assign wire19587 = ( n_n46  &  n_n134 ) | ( n_n43  &  n_n183 ) ;
 assign wire19588 = ( n_n46  &  n_n130 ) | ( n_n47  &  n_n130 ) | ( n_n46  &  wire1675 ) | ( n_n47  &  wire1675 ) ;
 assign wire19589 = ( n_n6266 ) | ( n_n6268 ) | ( n_n43  &  wire107 ) ;
 assign wire19591 = ( wire19589 ) | ( n_n42  &  wire107 ) | ( n_n42  &  wire340 ) ;
 assign wire19596 = ( wire2204 ) | ( wire2205 ) | ( n_n46  &  wire46 ) ;
 assign wire19599 = ( n_n47  &  wire48 ) | ( n_n47  &  wire124 ) ;
 assign wire19600 = ( n_n47  &  wire46 ) | ( n_n47  &  wire167 ) | ( n_n47  &  wire165 ) ;
 assign wire19602 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19603 = ( n_n108  &  wire401 ) | ( n_n108  &  n_n216  &  wire719 ) ;
 assign wire19605 = ( wire720  &  n_n156 ) | ( n_n156  &  wire719 ) | ( n_n156  &  wire715 ) ;
 assign wire19607 = ( wire724  &  n_n149 ) | ( n_n156  &  wire719 ) ;
 assign wire19608 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire719 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire719 ) ;
 assign wire19610 = ( wire445 ) | ( wire228  &  n_n170  &  wire719 ) ;
 assign wire19612 = ( wire2190 ) | ( wire2195 ) | ( wire2197 ) | ( wire19603 ) ;
 assign wire19613 = ( wire446 ) | ( wire4827 ) | ( wire4828 ) ;
 assign wire19614 = ( n_n47  &  wire151 ) | ( n_n46  &  wire47 ) ;
 assign wire19617 = ( wire2181 ) | ( wire19613 ) | ( n_n46  &  wire151 ) ;
 assign wire19619 = ( n_n772 ) | ( wire2191 ) | ( wire19610 ) | ( wire19612 ) ;
 assign wire19620 = ( wire724  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire715 ) ;
 assign wire19621 = ( n_n199  &  wire724 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire715 ) ;
 assign wire19623 = ( wire2176 ) | ( wire2179 ) | ( wire2180 ) ;
 assign wire19624 = ( wire724  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire715 ) ;
 assign wire19629 = ( wire2174 ) | ( n_n101  &  wire1706 ) | ( n_n101  &  wire1740 ) ;
 assign wire19630 = ( wire724  &  n_n170 ) | ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) ;
 assign wire19633 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire724 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire724 ) ;
 assign wire19636 = ( wire2169 ) | ( n_n108  &  wire1742 ) | ( n_n108  &  wire1756 ) ;
 assign wire19637 = ( wire19636 ) | ( n_n101  &  wire1743 ) ;
 assign wire19638 = ( wire2172 ) | ( wire2177 ) | ( wire19623 ) | ( wire19629 ) ;
 assign wire19640 = ( i_9_  &  i_10_  &  i_11_  &  wire719 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire719 ) ;
 assign wire19641 = ( wire724  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire715 ) ;
 assign wire19644 = ( n_n125  &  n_n142 ) | ( n_n125  &  n_n116 ) | ( n_n123  &  n_n116 ) ;
 assign wire19645 = ( wire2157 ) | ( wire19644 ) ;
 assign wire19646 = ( wire2163 ) | ( n_n123  &  wire856 ) | ( n_n123  &  wire859 ) ;
 assign wire19647 = ( n_n113  &  n_n116 ) | ( n_n112  &  wire1084 ) ;
 assign wire19648 = ( i_15_  &  n_n184  &  n_n207 ) | ( (~ i_15_)  &  n_n184  &  n_n207 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire19650 = ( n_n125  &  n_n132 ) | ( n_n123  &  n_n132 ) | ( n_n123  &  wire1087 ) ;
 assign wire19652 = ( wire19650 ) | ( n_n113  &  wire107 ) | ( n_n113  &  wire19648 ) ;
 assign wire19653 = ( wire2146 ) | ( wire2149 ) | ( wire2153 ) | ( wire19647 ) ;
 assign wire19654 = ( wire724  &  n_n170 ) | ( n_n170  &  wire720 ) | ( n_n170  &  wire715 ) ;
 assign wire19656 = ( wire2141 ) | ( wire2155 ) | ( wire2156 ) ;
 assign wire19657 = ( wire19656 ) | ( n_n125  &  wire1758 ) ;
 assign wire19658 = ( wire19645 ) | ( wire19646 ) | ( wire19652 ) | ( wire19653 ) ;
 assign wire19659 = ( n_n197  &  n_n130 ) | ( n_n212  &  n_n130 ) | ( n_n197  &  n_n128 ) | ( n_n212  &  n_n128 ) ;
 assign wire19660 = ( wire724  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire715 ) ;
 assign wire19663 = ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire724 ) ;
 assign wire19666 = ( wire2136 ) | ( n_n125  &  wire1259 ) | ( n_n125  &  wire1260 ) ;
 assign wire19667 = ( n_n197  &  n_n140 ) | ( n_n212  &  n_n140 ) | ( n_n212  &  n_n142 ) ;
 assign wire19668 = ( n_n212  &  wire55 ) | ( n_n197  &  n_n134 ) ;
 assign wire19670 = ( wire2124 ) | ( wire2130 ) | ( wire19667 ) ;
 assign wire19671 = ( wire2125 ) | ( wire19668 ) | ( wire188  &  n_n132 ) ;
 assign wire19672 = ( n_n199  &  wire724 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire715 ) ;
 assign wire19674 = ( wire2119 ) | ( wire2139 ) | ( wire19659 ) ;
 assign wire19675 = ( wire19674 ) | ( n_n123  &  wire1775 ) ;
 assign wire19676 = ( wire2134 ) | ( wire19666 ) | ( wire19670 ) | ( wire19671 ) ;
 assign wire19677 = ( n_n752 ) | ( wire19538 ) | ( wire19539 ) | ( wire19541 ) ;
 assign wire19680 = ( wire19637 ) | ( wire19638 ) | ( wire19657 ) | ( wire19658 ) ;
 assign wire19682 = ( n_n745 ) | ( n_n746 ) | ( n_n747 ) | ( n_n748 ) ;
 assign wire19683 = ( wire19675 ) | ( wire19676 ) | ( wire19677 ) | ( wire19680 ) ;
 assign wire19687 = ( n_n31  &  wire777 ) | ( n_n30  &  wire776 ) ;
 assign wire19688 = ( n_n5144 ) | ( wire19687 ) | ( wire213  &  wire775 ) ;
 assign wire19689 = ( wire2336 ) | ( wire19477 ) | ( wire19479 ) | ( wire19688 ) ;
 assign wire19691 = ( n_n31  &  wire1416 ) | ( n_n31  &  wire1414 ) | ( n_n30  &  wire1414 ) ;
 assign wire19693 = ( n_n7242 ) | ( n_n30  &  n_n156  &  wire728 ) ;
 assign wire19694 = ( n_n7263 ) | ( n_n3276 ) | ( n_n2948 ) ;
 assign wire19695 = ( n_n31  &  n_n52 ) | ( wire751  &  wire1367 ) ;
 assign wire19698 = ( wire2108 ) | ( wire19691 ) | ( wire19693 ) | ( wire19694 ) ;
 assign wire19700 = ( wire354 ) | ( wire140 ) ;
 assign wire19701 = ( wire730  &  n_n156 ) | ( wire718  &  n_n156 ) ;
 assign wire19702 = ( n_n6492 ) | ( n_n40  &  wire1447 ) | ( n_n40  &  wire19700 ) ;
 assign wire19704 = ( n_n41  &  n_n62 ) | ( n_n40  &  n_n62 ) | ( n_n40  &  wire1476 ) ;
 assign wire19706 = ( n_n177  &  wire720 ) | ( n_n170  &  wire720 ) | ( n_n177  &  wire727 ) | ( n_n170  &  wire727 ) ;
 assign wire19707 = ( n_n40  &  n_n58 ) | ( n_n41  &  wire1478 ) | ( n_n40  &  wire1478 ) ;
 assign wire19708 = ( n_n54  &  wire1480 ) | ( n_n38  &  wire1479 ) ;
 assign wire19709 = ( wire19707 ) | ( n_n39  &  wire244 ) | ( n_n39  &  wire19706 ) ;
 assign wire19710 = ( wire19704 ) | ( wire19708 ) | ( n_n41  &  wire1477 ) ;
 assign wire19714 = ( i_15_  &  n_n216  &  n_n205 ) | ( (~ i_15_)  &  n_n216  &  n_n205 ) | ( i_15_  &  n_n216  &  n_n215 ) ;
 assign wire19716 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( i_15_  &  n_n184  &  n_n215 ) ;
 assign wire19717 = ( n_n34  &  n_n183 ) | ( n_n36  &  n_n176 ) ;
 assign wire19718 = ( n_n34  &  wire63 ) | ( n_n36  &  wire348 ) ;
 assign wire19721 = ( wire19718 ) | ( wire137  &  n_n36 ) | ( n_n36  &  wire63 ) ;
 assign wire19722 = ( wire2070 ) | ( wire2078 ) | ( wire2079 ) | ( wire19717 ) ;
 assign wire19724 = ( n_n170  &  wire720 ) | ( n_n177  &  wire718 ) ;
 assign wire19725 = ( n_n34  &  wire126 ) | ( n_n34  &  wire933 ) ;
 assign wire19726 = ( n_n177  &  wire718 ) | ( wire720  &  n_n149 ) ;
 assign wire19727 = ( n_n170  &  wire718 ) | ( wire720  &  n_n156 ) ;
 assign wire19728 = ( (~ i_15_)  &  n_n170  &  n_n205 ) | ( i_15_  &  n_n156  &  n_n205 ) | ( (~ i_15_)  &  n_n156  &  n_n205 ) ;
 assign wire19730 = ( n_n34  &  n_n176 ) | ( n_n36  &  wire126 ) ;
 assign wire19731 = ( wire137  &  n_n34 ) | ( n_n34  &  n_n171 ) | ( n_n34  &  wire19726 ) ;
 assign wire19732 = ( wire19731 ) | ( wire19730 ) ;
 assign wire19733 = ( wire2062 ) | ( wire2068 ) | ( wire19725 ) ;
 assign wire19734 = ( n_n36  &  n_n198 ) | ( n_n34  &  wire385 ) ;
 assign wire19735 = ( n_n36  &  wire68 ) | ( n_n34  &  wire68 ) ;
 assign wire19738 = ( n_n369 ) | ( n_n371 ) | ( wire19734 ) | ( wire19735 ) ;
 assign wire19739 = ( wire19721 ) | ( wire19722 ) | ( wire19732 ) | ( wire19733 ) ;
 assign wire19744 = ( wire166 ) | ( wire269 ) | ( wire332 ) ;
 assign wire19745 = ( n_n40  &  wire1684 ) | ( n_n40  &  wire726  &  n_n216 ) ;
 assign wire19746 = ( n_n41  &  wire726  &  n_n216 ) | ( n_n41  &  n_n216  &  wire720 ) ;
 assign wire19747 = ( n_n42  &  n_n136 ) | ( n_n43  &  n_n136 ) | ( n_n42  &  n_n60 ) ;
 assign wire19750 = ( n_n41  &  wire296 ) | ( n_n40  &  wire296 ) | ( n_n40  &  wire332 ) ;
 assign wire19751 = ( wire2040 ) | ( wire2041 ) | ( n_n42  &  n_n190 ) ;
 assign wire19752 = ( wire2045 ) | ( wire19746 ) | ( wire19747 ) | ( wire19750 ) ;
 assign wire19756 = ( n_n41  &  wire1617 ) | ( n_n41  &  wire726  &  n_n177 ) ;
 assign wire19757 = ( wire2035 ) | ( wire2051 ) | ( wire19745 ) ;
 assign wire19758 = ( wire19751 ) | ( wire19752 ) | ( wire19756 ) ;
 assign wire19759 = ( wire726  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire19760 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign wire19764 = ( wire161 ) | ( wire337 ) | ( wire726  &  n_n191 ) ;
 assign wire19765 = ( wire1992 ) | ( wire1995 ) | ( wire1996 ) ;
 assign wire19766 = ( wire726  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) ;
 assign wire19767 = ( n_n199  &  wire726 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire727 ) ;
 assign wire19769 = ( wire1987 ) | ( wire1990 ) | ( wire1991 ) ;
 assign wire19770 = ( i_9_  &  (~ i_10_)  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire726 ) ;
 assign wire19774 = ( wire110 ) | ( wire329 ) | ( wire726  &  n_n170 ) ;
 assign wire19775 = ( wire1982 ) | ( wire1997 ) | ( wire1998 ) ;
 assign wire19777 = ( wire1988 ) | ( wire1993 ) | ( wire19765 ) | ( wire19769 ) ;
 assign wire19778 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire19779 = ( n_n101  &  n_n136 ) | ( n_n108  &  n_n136 ) | ( n_n108  &  wire1357 ) ;
 assign wire19780 = ( (~ i_15_)  &  n_n156  &  n_n209 ) | ( i_15_  &  n_n156  &  n_n215 ) | ( (~ i_15_)  &  n_n156  &  n_n215 ) ;
 assign wire19782 = ( i_9_  &  i_10_  &  (~ i_11_)  &  wire728 ) | ( (~ i_9_)  &  i_10_  &  (~ i_11_)  &  wire728 ) ;
 assign wire19783 = ( wire726  &  n_n149 ) | ( n_n177  &  wire728 ) ;
 assign wire19786 = ( wire419 ) | ( wire2027 ) | ( wire228  &  n_n56 ) ;
 assign wire19787 = ( wire2026 ) | ( wire2032 ) | ( wire19779 ) ;
 assign wire19792 = ( n_n6005 ) | ( wire4354 ) | ( wire4355 ) ;
 assign wire19793 = ( wire19792 ) | ( wire1640  &  wire1639 ) ;
 assign wire19796 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire19798 = ( wire140 ) | ( wire244 ) | ( wire414 ) ;
 assign wire19799 = ( n_n62  &  wire189 ) | ( n_n47  &  wire1636 ) ;
 assign wire19800 = ( n_n43  &  n_n183 ) | ( n_n42  &  wire346 ) ;
 assign wire19801 = ( n_n42  &  wire128 ) | ( n_n43  &  wire128 ) ;
 assign wire19802 = ( n_n42  &  n_n183 ) | ( n_n46  &  n_n58 ) ;
 assign wire19803 = ( i_8_  &  n_n16  &  wire739 ) | ( (~ i_8_)  &  n_n16  &  wire739 ) | ( i_8_  &  n_n16  &  wire759 ) | ( (~ i_8_)  &  n_n16  &  wire759 ) ;
 assign wire19804 = ( n_n43  &  n_n190 ) | ( wire189  &  wire1666 ) ;
 assign wire19807 = ( wire2004 ) | ( wire19802 ) | ( n_n54  &  wire1668 ) ;
 assign wire19808 = ( wire19800 ) | ( wire19801 ) | ( wire19803 ) | ( wire19804 ) ;
 assign wire19812 = ( wire1999 ) | ( wire2000 ) | ( wire19807 ) | ( wire19808 ) ;
 assign wire19813 = ( n_n302 ) | ( wire1983 ) | ( wire19775 ) | ( wire19777 ) ;
 assign wire19820 = ( wire236 ) | ( wire282 ) | ( wire354 ) ;
 assign wire19823 = ( n_n197  &  wire1366 ) | ( n_n212  &  wire1366 ) | ( n_n212  &  wire166 ) ;
 assign wire19824 = ( wire1936 ) | ( wire1937 ) | ( wire1938 ) | ( wire1939 ) ;
 assign wire19825 = ( n_n197  &  n_n62 ) | ( n_n212  &  n_n62 ) | ( n_n212  &  n_n64 ) ;
 assign wire19827 = ( i_9_  &  i_10_  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire19828 = ( wire1979 ) | ( wire19825 ) | ( wire188  &  n_n56 ) ;
 assign wire19829 = ( wire1976 ) | ( n_n212  &  wire1440 ) ;
 assign wire19830 = ( n_n197  &  n_n54 ) | ( n_n212  &  n_n54 ) | ( n_n197  &  n_n52 ) | ( n_n212  &  n_n52 ) ;
 assign wire19831 = ( wire726  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) ;
 assign wire19834 = ( wire1971 ) | ( n_n123  &  wire1510 ) | ( n_n123  &  wire1512 ) ;
 assign wire19835 = ( n_n199  &  wire726 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire727 ) ;
 assign wire19837 = ( wire1962 ) | ( wire1972 ) | ( wire19830 ) ;
 assign wire19838 = ( wire19837 ) | ( n_n123  &  wire1587 ) ;
 assign wire19839 = ( wire1968 ) | ( wire19828 ) | ( wire19829 ) | ( wire19834 ) ;
 assign wire19841 = ( n_n113  &  n_n183 ) | ( wire255  &  n_n56 ) ;
 assign wire19842 = ( n_n125  &  wire1717 ) | ( n_n123  &  wire1716 ) ;
 assign wire19843 = ( i_15_  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n205 ) | ( (~ i_15_)  &  n_n184  &  n_n215 ) ;
 assign wire19845 = ( n_n112  &  wire63 ) | ( n_n112  &  wire1720 ) ;
 assign wire19846 = ( wire1951 ) | ( n_n113  &  wire128 ) | ( n_n113  &  wire19843 ) ;
 assign wire19847 = ( wire19841 ) | ( wire19842 ) | ( wire19845 ) ;
 assign wire19848 = ( wire726  &  n_n156 ) | ( n_n216  &  wire728 ) ;
 assign wire19850 = ( wire726  &  n_n149 ) | ( n_n191  &  wire728 ) ;
 assign wire19853 = ( wire207 ) | ( wire249 ) | ( n_n216  &  wire728 ) ;
 assign wire19854 = ( wire1945 ) | ( n_n184  &  wire255  &  wire728 ) ;
 assign wire19856 = ( wire726  &  n_n170 ) | ( n_n170  &  wire720 ) | ( n_n170  &  wire727 ) ;
 assign wire19858 = ( wire1940 ) | ( wire1960 ) | ( wire1961 ) ;
 assign wire19859 = ( wire19858 ) | ( n_n125  &  wire1761 ) ;
 assign wire19861 = ( wire19823 ) | ( wire19824 ) | ( wire19838 ) | ( wire19839 ) ;
 assign wire19862 = ( n_n38  &  n_n54 ) | ( n_n39  &  n_n54 ) | ( n_n38  &  n_n52 ) ;
 assign wire19864 = ( n_n519 ) | ( wire19862 ) | ( n_n38  &  wire140 ) ;
 assign wire19865 = ( wire5022 ) | ( wire5023 ) | ( wire5024 ) | ( wire5025 ) ;
 assign wire19867 = ( wire19709 ) | ( wire19710 ) | ( wire19864 ) | ( wire19865 ) ;
 assign wire19868 = ( wire19702 ) | ( wire19867 ) | ( n_n41  &  wire1446 ) ;
 assign wire19869 = ( wire19738 ) | ( wire19739 ) | ( wire19757 ) | ( wire19758 ) ;
 assign wire19871 = ( n_n301 ) | ( n_n304 ) | ( wire19813 ) | ( wire19861 ) ;
 assign wire19874 = ( wire166 ) | ( wire235 ) | ( wire283 ) ;
 assign wire19875 = ( n_n34  &  n_n58 ) | ( n_n36  &  n_n56 ) ;
 assign wire19876 = ( n_n36  &  n_n54 ) | ( n_n34  &  n_n54 ) | ( n_n36  &  n_n52 ) | ( n_n34  &  n_n52 ) ;
 assign wire19878 = ( wire1914 ) | ( wire19875 ) | ( wire19876 ) ;
 assign wire19879 = ( (~ i_9_)  &  (~ i_10_)  &  i_11_  &  wire728 ) | ( i_9_  &  (~ i_10_)  &  (~ i_11_)  &  wire728 ) ;
 assign wire19880 = ( n_n33  &  n_n52 ) | ( n_n31  &  wire335 ) ;
 assign wire19882 = ( n_n199  &  wire726 ) | ( n_n199  &  wire720 ) | ( n_n199  &  wire727 ) ;
 assign wire19884 = ( wire1907 ) | ( wire1910 ) | ( wire1912 ) | ( wire19880 ) ;
 assign wire19886 = ( n_n36  &  wire1778 ) | ( n_n36  &  wire1777 ) | ( n_n34  &  wire1777 ) ;
 assign wire19887 = ( n_n36  &  wire127 ) | ( n_n34  &  wire1780 ) ;
 assign wire19888 = ( wire726  &  n_n149 ) | ( n_n216  &  wire728 ) ;
 assign wire19890 = ( wire556 ) | ( n_n34  &  wire156 ) | ( n_n34  &  wire1570 ) ;
 assign wire19891 = ( wire542 ) | ( wire1906 ) | ( wire19886 ) | ( wire19887 ) ;
 assign wire19893 = ( wire1908 ) | ( wire1916 ) | ( wire19878 ) | ( wire19884 ) ;
 assign wire19895 = ( wire726  &  n_n177 ) | ( n_n177  &  wire720 ) | ( n_n177  &  wire727 ) ;
 assign wire19898 = ( wire520 ) | ( n_n30  &  wire1311 ) | ( n_n30  &  wire1482 ) ;
 assign wire19899 = ( wire726  &  n_n191 ) | ( n_n191  &  wire720 ) | ( n_n191  &  wire727 ) ;
 assign wire19901 = ( i_9_  &  i_10_  &  i_11_  &  wire726 ) | ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_)  &  wire726 ) ;
 assign wire19904 = ( wire507 ) | ( wire510 ) | ( wire513 ) ;
 assign wire19905 = ( wire726  &  n_n149 ) | ( wire720  &  n_n149 ) | ( n_n149  &  wire727 ) ;
 assign wire19907 = ( wire499 ) | ( wire552 ) | ( n_n31  &  wire1090 ) ;
 assign wire19909 = ( wire508 ) | ( wire516 ) | ( wire19898 ) | ( wire19904 ) ;
 assign wire19910 = ( n_n5144 ) | ( n_n18  &  n_n159  &  n_n218 ) ;
 assign wire19911 = ( wire19910 ) | ( n_n3  &  wire185 ) ;
 assign wire19912 = ( wire2099 ) | ( wire19695 ) | ( wire19698 ) | ( wire19911 ) ;
 assign wire19913 = ( wire19890 ) | ( wire19891 ) | ( wire19893 ) | ( wire19912 ) ;
 assign wire19914 = ( wire501 ) | ( wire19907 ) | ( wire19909 ) | ( wire19913 ) ;
 assign wire19916 = ( wire95 ) | ( wire729  &  n_n191 ) | ( wire729  &  n_n156 ) ;
 assign wire19917 = ( n_n5144 ) | ( n_n162  &  n_n18  &  n_n219 ) ;
 assign wire19920 = ( n_n7253 ) | ( wire389 ) | ( wire706 ) | ( wire19917 ) ;
 assign wire19922 = ( wire454 ) | ( wire19920 ) | ( wire742  &  wire779 ) ;
 assign wire19923 = ( n_n5144 ) | ( n_n157  &  n_n219  &  n_n111 ) ;
 assign wire19925 = ( wire388 ) | ( wire267  &  wire781 ) ;
 assign wire19926 = ( n_n3389 ) | ( wire19923 ) | ( n_n135  &  wire783 ) ;
 assign wire19928 = ( wire467 ) | ( wire19925 ) | ( wire19926 ) ;
 assign wire19929 = ( i_7_  &  (~ i_6_)  &  n_n48  &  n_n219 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n48  &  n_n219 ) ;
 assign wire19930 = ( i_7_  &  (~ i_6_)  &  n_n219  &  n_n218 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n219  &  n_n218 ) ;
 assign wire19933 = ( n_n7264 ) | ( n_n7262 ) | ( wire19930 ) ;
 assign wire19935 = ( wire95 ) | ( wire729  &  n_n191 ) | ( wire729  &  n_n156 ) ;
 assign wire19938 = ( wire551 ) | ( n_n191  &  wire725  &  wire18833 ) ;
 assign wire19939 = ( n_n7242 ) | ( wire462 ) | ( n_n59  &  wire751 ) ;
 assign wire19941 = ( n_n7260 ) | ( wire439 ) | ( wire19938 ) | ( wire19939 ) ;
 assign wire19943 = ( n_n5144 ) | ( n_n18  &  n_n159  &  n_n218 ) ;
 assign wire19944 = ( wire19943 ) | ( wire77  &  n_n3 ) ;
 assign wire19946 = ( wire707 ) | ( wire138 ) | ( wire19944 ) ;


endmodule

