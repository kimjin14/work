`include "FPGA/define.v"

module fpga_top (
	input fpga_clk,
	input fpga_rst,
	inout [7:0]io_0_1_wire,
	inout [7:0]io_0_2_wire,
	inout [7:0]io_0_3_wire,
	inout [7:0]io_0_4_wire,
	inout [7:0]io_0_5_wire,
	inout [7:0]io_0_6_wire,
	inout [7:0]io_0_7_wire,
	inout [7:0]io_0_8_wire,
	inout [7:0]io_0_9_wire,
	inout [7:0]io_1_0_wire,
	inout [7:0]io_1_10_wire,
	inout [7:0]io_2_0_wire,
	inout [7:0]io_2_10_wire,
	inout [7:0]io_3_0_wire,
	inout [7:0]io_3_10_wire,
	inout [7:0]io_4_0_wire,
	inout [7:0]io_4_10_wire,
	inout [7:0]io_5_0_wire,
	inout [7:0]io_5_10_wire,
	inout [7:0]io_6_0_wire,
	inout [7:0]io_6_10_wire,
	inout [7:0]io_7_0_wire,
	inout [7:0]io_7_10_wire,
	inout [7:0]io_8_0_wire,
	inout [7:0]io_8_10_wire,
	inout [7:0]io_9_0_wire,
	inout [7:0]io_9_10_wire,
	inout [7:0]io_10_1_wire,
	inout [7:0]io_10_2_wire,
	inout [7:0]io_10_3_wire,
	inout [7:0]io_10_4_wire,
	inout [7:0]io_10_5_wire,
	inout [7:0]io_10_6_wire,
	inout [7:0]io_10_7_wire,
	inout [7:0]io_10_8_wire,
	inout [7:0]io_10_9_wire,
	input config_rst,
	input config_clk,
	input config_in
);

wire n24; //IPIN -1 (0,1) #0
wire n25; //OPIN -1 (0,1) #1
wire n26; //IPIN -1 (0,1) #2
wire n27; //IPIN -1 (0,1) #3
wire n28; //OPIN -1 (0,1) #4
wire n29; //IPIN -1 (0,1) #5
wire n30; //IPIN -1 (0,1) #6
wire n31; //OPIN -1 (0,1) #7
wire n32; //IPIN -1 (0,1) #8
wire n33; //IPIN -1 (0,1) #9
wire n34; //OPIN -1 (0,1) #10
wire n35; //IPIN -1 (0,1) #11
wire n36; //IPIN -1 (0,1) #12
wire n37; //OPIN -1 (0,1) #13
wire n38; //IPIN -1 (0,1) #14
wire n39; //IPIN -1 (0,1) #15
wire n40; //OPIN -1 (0,1) #16
wire n41; //IPIN -1 (0,1) #17
wire n42; //IPIN -1 (0,1) #18
wire n43; //OPIN -1 (0,1) #19
wire n44; //IPIN -1 (0,1) #20
wire n45; //IPIN -1 (0,1) #21
wire n46; //OPIN -1 (0,1) #22
wire n47; //IPIN -1 (0,1) #23
wire n72; //IPIN -1 (0,2) #0
wire n73; //OPIN -1 (0,2) #1
wire n74; //IPIN -1 (0,2) #2
wire n75; //IPIN -1 (0,2) #3
wire n76; //OPIN -1 (0,2) #4
wire n77; //IPIN -1 (0,2) #5
wire n78; //IPIN -1 (0,2) #6
wire n79; //OPIN -1 (0,2) #7
wire n80; //IPIN -1 (0,2) #8
wire n81; //IPIN -1 (0,2) #9
wire n82; //OPIN -1 (0,2) #10
wire n83; //IPIN -1 (0,2) #11
wire n84; //IPIN -1 (0,2) #12
wire n85; //OPIN -1 (0,2) #13
wire n86; //IPIN -1 (0,2) #14
wire n87; //IPIN -1 (0,2) #15
wire n88; //OPIN -1 (0,2) #16
wire n89; //IPIN -1 (0,2) #17
wire n90; //IPIN -1 (0,2) #18
wire n91; //OPIN -1 (0,2) #19
wire n92; //IPIN -1 (0,2) #20
wire n93; //IPIN -1 (0,2) #21
wire n94; //OPIN -1 (0,2) #22
wire n95; //IPIN -1 (0,2) #23
wire n120; //IPIN -1 (0,3) #0
wire n121; //OPIN -1 (0,3) #1
wire n122; //IPIN -1 (0,3) #2
wire n123; //IPIN -1 (0,3) #3
wire n124; //OPIN -1 (0,3) #4
wire n125; //IPIN -1 (0,3) #5
wire n126; //IPIN -1 (0,3) #6
wire n127; //OPIN -1 (0,3) #7
wire n128; //IPIN -1 (0,3) #8
wire n129; //IPIN -1 (0,3) #9
wire n130; //OPIN -1 (0,3) #10
wire n131; //IPIN -1 (0,3) #11
wire n132; //IPIN -1 (0,3) #12
wire n133; //OPIN -1 (0,3) #13
wire n134; //IPIN -1 (0,3) #14
wire n135; //IPIN -1 (0,3) #15
wire n136; //OPIN -1 (0,3) #16
wire n137; //IPIN -1 (0,3) #17
wire n138; //IPIN -1 (0,3) #18
wire n139; //OPIN -1 (0,3) #19
wire n140; //IPIN -1 (0,3) #20
wire n141; //IPIN -1 (0,3) #21
wire n142; //OPIN -1 (0,3) #22
wire n143; //IPIN -1 (0,3) #23
wire n168; //IPIN -1 (0,4) #0
wire n169; //OPIN -1 (0,4) #1
wire n170; //IPIN -1 (0,4) #2
wire n171; //IPIN -1 (0,4) #3
wire n172; //OPIN -1 (0,4) #4
wire n173; //IPIN -1 (0,4) #5
wire n174; //IPIN -1 (0,4) #6
wire n175; //OPIN -1 (0,4) #7
wire n176; //IPIN -1 (0,4) #8
wire n177; //IPIN -1 (0,4) #9
wire n178; //OPIN -1 (0,4) #10
wire n179; //IPIN -1 (0,4) #11
wire n180; //IPIN -1 (0,4) #12
wire n181; //OPIN -1 (0,4) #13
wire n182; //IPIN -1 (0,4) #14
wire n183; //IPIN -1 (0,4) #15
wire n184; //OPIN -1 (0,4) #16
wire n185; //IPIN -1 (0,4) #17
wire n186; //IPIN -1 (0,4) #18
wire n187; //OPIN -1 (0,4) #19
wire n188; //IPIN -1 (0,4) #20
wire n189; //IPIN -1 (0,4) #21
wire n190; //OPIN -1 (0,4) #22
wire n191; //IPIN -1 (0,4) #23
wire n216; //IPIN -1 (0,5) #0
wire n217; //OPIN -1 (0,5) #1
wire n218; //IPIN -1 (0,5) #2
wire n219; //IPIN -1 (0,5) #3
wire n220; //OPIN -1 (0,5) #4
wire n221; //IPIN -1 (0,5) #5
wire n222; //IPIN -1 (0,5) #6
wire n223; //OPIN -1 (0,5) #7
wire n224; //IPIN -1 (0,5) #8
wire n225; //IPIN -1 (0,5) #9
wire n226; //OPIN -1 (0,5) #10
wire n227; //IPIN -1 (0,5) #11
wire n228; //IPIN -1 (0,5) #12
wire n229; //OPIN -1 (0,5) #13
wire n230; //IPIN -1 (0,5) #14
wire n231; //IPIN -1 (0,5) #15
wire n232; //OPIN -1 (0,5) #16
wire n233; //IPIN -1 (0,5) #17
wire n234; //IPIN -1 (0,5) #18
wire n235; //OPIN -1 (0,5) #19
wire n236; //IPIN -1 (0,5) #20
wire n237; //IPIN -1 (0,5) #21
wire n238; //OPIN -1 (0,5) #22
wire n239; //IPIN -1 (0,5) #23
wire n264; //IPIN -1 (0,6) #0
wire n265; //OPIN -1 (0,6) #1
wire n266; //IPIN -1 (0,6) #2
wire n267; //IPIN -1 (0,6) #3
wire n268; //OPIN -1 (0,6) #4
wire n269; //IPIN -1 (0,6) #5
wire n270; //IPIN -1 (0,6) #6
wire n271; //OPIN -1 (0,6) #7
wire n272; //IPIN -1 (0,6) #8
wire n273; //IPIN -1 (0,6) #9
wire n274; //OPIN -1 (0,6) #10
wire n275; //IPIN -1 (0,6) #11
wire n276; //IPIN -1 (0,6) #12
wire n277; //OPIN -1 (0,6) #13
wire n278; //IPIN -1 (0,6) #14
wire n279; //IPIN -1 (0,6) #15
wire n280; //OPIN -1 (0,6) #16
wire n281; //IPIN -1 (0,6) #17
wire n282; //IPIN -1 (0,6) #18
wire n283; //OPIN -1 (0,6) #19
wire n284; //IPIN -1 (0,6) #20
wire n285; //IPIN -1 (0,6) #21
wire n286; //OPIN -1 (0,6) #22
wire n287; //IPIN -1 (0,6) #23
wire n312; //IPIN -1 (0,7) #0
wire n313; //OPIN -1 (0,7) #1
wire n314; //IPIN -1 (0,7) #2
wire n315; //IPIN -1 (0,7) #3
wire n316; //OPIN -1 (0,7) #4
wire n317; //IPIN -1 (0,7) #5
wire n318; //IPIN -1 (0,7) #6
wire n319; //OPIN -1 (0,7) #7
wire n320; //IPIN -1 (0,7) #8
wire n321; //IPIN -1 (0,7) #9
wire n322; //OPIN -1 (0,7) #10
wire n323; //IPIN -1 (0,7) #11
wire n324; //IPIN -1 (0,7) #12
wire n325; //OPIN -1 (0,7) #13
wire n326; //IPIN -1 (0,7) #14
wire n327; //IPIN -1 (0,7) #15
wire n328; //OPIN -1 (0,7) #16
wire n329; //IPIN -1 (0,7) #17
wire n330; //IPIN -1 (0,7) #18
wire n331; //OPIN -1 (0,7) #19
wire n332; //IPIN -1 (0,7) #20
wire n333; //IPIN -1 (0,7) #21
wire n334; //OPIN -1 (0,7) #22
wire n335; //IPIN -1 (0,7) #23
wire n360; //IPIN -1 (0,8) #0
wire n361; //OPIN -1 (0,8) #1
wire n362; //IPIN -1 (0,8) #2
wire n363; //IPIN -1 (0,8) #3
wire n364; //OPIN -1 (0,8) #4
wire n365; //IPIN -1 (0,8) #5
wire n366; //IPIN -1 (0,8) #6
wire n367; //OPIN -1 (0,8) #7
wire n368; //IPIN -1 (0,8) #8
wire n369; //IPIN -1 (0,8) #9
wire n370; //OPIN -1 (0,8) #10
wire n371; //IPIN -1 (0,8) #11
wire n372; //IPIN -1 (0,8) #12
wire n373; //OPIN -1 (0,8) #13
wire n374; //IPIN -1 (0,8) #14
wire n375; //IPIN -1 (0,8) #15
wire n376; //OPIN -1 (0,8) #16
wire n377; //IPIN -1 (0,8) #17
wire n378; //IPIN -1 (0,8) #18
wire n379; //OPIN -1 (0,8) #19
wire n380; //IPIN -1 (0,8) #20
wire n381; //IPIN -1 (0,8) #21
wire n382; //OPIN -1 (0,8) #22
wire n383; //IPIN -1 (0,8) #23
wire n408; //IPIN -1 (0,9) #0
wire n409; //OPIN -1 (0,9) #1
wire n410; //IPIN -1 (0,9) #2
wire n411; //IPIN -1 (0,9) #3
wire n412; //OPIN -1 (0,9) #4
wire n413; //IPIN -1 (0,9) #5
wire n414; //IPIN -1 (0,9) #6
wire n415; //OPIN -1 (0,9) #7
wire n416; //IPIN -1 (0,9) #8
wire n417; //IPIN -1 (0,9) #9
wire n418; //OPIN -1 (0,9) #10
wire n419; //IPIN -1 (0,9) #11
wire n420; //IPIN -1 (0,9) #12
wire n421; //OPIN -1 (0,9) #13
wire n422; //IPIN -1 (0,9) #14
wire n423; //IPIN -1 (0,9) #15
wire n424; //OPIN -1 (0,9) #16
wire n425; //IPIN -1 (0,9) #17
wire n426; //IPIN -1 (0,9) #18
wire n427; //OPIN -1 (0,9) #19
wire n428; //IPIN -1 (0,9) #20
wire n429; //IPIN -1 (0,9) #21
wire n430; //OPIN -1 (0,9) #22
wire n431; //IPIN -1 (0,9) #23
wire n456; //IPIN -1 (1,0) #0
wire n457; //OPIN -1 (1,0) #1
wire n458; //IPIN -1 (1,0) #2
wire n459; //IPIN -1 (1,0) #3
wire n460; //OPIN -1 (1,0) #4
wire n461; //IPIN -1 (1,0) #5
wire n462; //IPIN -1 (1,0) #6
wire n463; //OPIN -1 (1,0) #7
wire n464; //IPIN -1 (1,0) #8
wire n465; //IPIN -1 (1,0) #9
wire n466; //OPIN -1 (1,0) #10
wire n467; //IPIN -1 (1,0) #11
wire n468; //IPIN -1 (1,0) #12
wire n469; //OPIN -1 (1,0) #13
wire n470; //IPIN -1 (1,0) #14
wire n471; //IPIN -1 (1,0) #15
wire n472; //OPIN -1 (1,0) #16
wire n473; //IPIN -1 (1,0) #17
wire n474; //IPIN -1 (1,0) #18
wire n475; //OPIN -1 (1,0) #19
wire n476; //IPIN -1 (1,0) #20
wire n477; //IPIN -1 (1,0) #21
wire n478; //OPIN -1 (1,0) #22
wire n479; //IPIN -1 (1,0) #23
wire n505; //IPIN -1 (1,1) #0
wire n506; //IPIN -1 (1,1) #1
wire n507; //IPIN -1 (1,1) #2
wire n508; //IPIN -1 (1,1) #3
wire n509; //IPIN -1 (1,1) #4
wire n510; //IPIN -1 (1,1) #5
wire n511; //IPIN -1 (1,1) #6
wire n512; //IPIN -1 (1,1) #7
wire n513; //IPIN -1 (1,1) #8
wire n514; //IPIN -1 (1,1) #9
wire n515; //IPIN -1 (1,1) #10
wire n516; //IPIN -1 (1,1) #11
wire n517; //IPIN -1 (1,1) #12
wire n518; //IPIN -1 (1,1) #13
wire n519; //IPIN -1 (1,1) #14
wire n520; //IPIN -1 (1,1) #15
wire n521; //IPIN -1 (1,1) #16
wire n522; //IPIN -1 (1,1) #17
wire n523; //IPIN -1 (1,1) #18
wire n524; //IPIN -1 (1,1) #19
wire n525; //IPIN -1 (1,1) #20
wire n526; //IPIN -1 (1,1) #21
wire n527; //IPIN -1 (1,1) #22
wire n528; //IPIN -1 (1,1) #23
wire n529; //IPIN -1 (1,1) #24
wire n530; //IPIN -1 (1,1) #25
wire n531; //IPIN -1 (1,1) #26
wire n532; //IPIN -1 (1,1) #27
wire n533; //IPIN -1 (1,1) #28
wire n534; //IPIN -1 (1,1) #29
wire n535; //IPIN -1 (1,1) #30
wire n536; //IPIN -1 (1,1) #31
wire n537; //IPIN -1 (1,1) #32
wire n538; //IPIN -1 (1,1) #33
wire n539; //IPIN -1 (1,1) #34
wire n540; //IPIN -1 (1,1) #35
wire n541; //IPIN -1 (1,1) #36
wire n542; //IPIN -1 (1,1) #37
wire n543; //IPIN -1 (1,1) #38
wire n544; //IPIN -1 (1,1) #39
wire n545; //IPIN -1 (1,1) #40
wire n546; //IPIN -1 (1,1) #41
wire n547; //IPIN -1 (1,1) #42
wire n548; //IPIN -1 (1,1) #43
wire n549; //IPIN -1 (1,1) #44
wire n550; //IPIN -1 (1,1) #45
wire n551; //IPIN -1 (1,1) #46
wire n552; //IPIN -1 (1,1) #47
wire n553; //IPIN -1 (1,1) #48
wire n554; //IPIN -1 (1,1) #49
wire n555; //IPIN -1 (1,1) #50
wire n556; //IPIN -1 (1,1) #51
wire n557; //OPIN -1 (1,1) #52
wire n558; //OPIN -1 (1,1) #53
wire n559; //OPIN -1 (1,1) #54
wire n560; //OPIN -1 (1,1) #55
wire n561; //OPIN -1 (1,1) #56
wire n562; //OPIN -1 (1,1) #57
wire n563; //OPIN -1 (1,1) #58
wire n564; //OPIN -1 (1,1) #59
wire n565; //OPIN -1 (1,1) #60
wire n566; //OPIN -1 (1,1) #61
wire n567; //OPIN -1 (1,1) #62
wire n568; //OPIN -1 (1,1) #63
wire n569; //OPIN -1 (1,1) #64
wire n570; //OPIN -1 (1,1) #65
wire n571; //OPIN -1 (1,1) #66
wire n572; //OPIN -1 (1,1) #67
wire n573; //OPIN -1 (1,1) #68
wire n574; //OPIN -1 (1,1) #69
wire n575; //OPIN -1 (1,1) #70
wire n576; //OPIN -1 (1,1) #71
wire n577; //IPIN -1 (1,1) #72
wire n603; //IPIN -1 (1,2) #0
wire n604; //IPIN -1 (1,2) #1
wire n605; //IPIN -1 (1,2) #2
wire n606; //IPIN -1 (1,2) #3
wire n607; //IPIN -1 (1,2) #4
wire n608; //IPIN -1 (1,2) #5
wire n609; //IPIN -1 (1,2) #6
wire n610; //IPIN -1 (1,2) #7
wire n611; //IPIN -1 (1,2) #8
wire n612; //IPIN -1 (1,2) #9
wire n613; //IPIN -1 (1,2) #10
wire n614; //IPIN -1 (1,2) #11
wire n615; //IPIN -1 (1,2) #12
wire n616; //IPIN -1 (1,2) #13
wire n617; //IPIN -1 (1,2) #14
wire n618; //IPIN -1 (1,2) #15
wire n619; //IPIN -1 (1,2) #16
wire n620; //IPIN -1 (1,2) #17
wire n621; //IPIN -1 (1,2) #18
wire n622; //IPIN -1 (1,2) #19
wire n623; //IPIN -1 (1,2) #20
wire n624; //IPIN -1 (1,2) #21
wire n625; //IPIN -1 (1,2) #22
wire n626; //IPIN -1 (1,2) #23
wire n627; //IPIN -1 (1,2) #24
wire n628; //IPIN -1 (1,2) #25
wire n629; //IPIN -1 (1,2) #26
wire n630; //IPIN -1 (1,2) #27
wire n631; //IPIN -1 (1,2) #28
wire n632; //IPIN -1 (1,2) #29
wire n633; //IPIN -1 (1,2) #30
wire n634; //IPIN -1 (1,2) #31
wire n635; //IPIN -1 (1,2) #32
wire n636; //IPIN -1 (1,2) #33
wire n637; //IPIN -1 (1,2) #34
wire n638; //IPIN -1 (1,2) #35
wire n639; //IPIN -1 (1,2) #36
wire n640; //IPIN -1 (1,2) #37
wire n641; //IPIN -1 (1,2) #38
wire n642; //IPIN -1 (1,2) #39
wire n643; //IPIN -1 (1,2) #40
wire n644; //IPIN -1 (1,2) #41
wire n645; //IPIN -1 (1,2) #42
wire n646; //IPIN -1 (1,2) #43
wire n647; //IPIN -1 (1,2) #44
wire n648; //IPIN -1 (1,2) #45
wire n649; //IPIN -1 (1,2) #46
wire n650; //IPIN -1 (1,2) #47
wire n651; //IPIN -1 (1,2) #48
wire n652; //IPIN -1 (1,2) #49
wire n653; //IPIN -1 (1,2) #50
wire n654; //IPIN -1 (1,2) #51
wire n655; //OPIN -1 (1,2) #52
wire n656; //OPIN -1 (1,2) #53
wire n657; //OPIN -1 (1,2) #54
wire n658; //OPIN -1 (1,2) #55
wire n659; //OPIN -1 (1,2) #56
wire n660; //OPIN -1 (1,2) #57
wire n661; //OPIN -1 (1,2) #58
wire n662; //OPIN -1 (1,2) #59
wire n663; //OPIN -1 (1,2) #60
wire n664; //OPIN -1 (1,2) #61
wire n665; //OPIN -1 (1,2) #62
wire n666; //OPIN -1 (1,2) #63
wire n667; //OPIN -1 (1,2) #64
wire n668; //OPIN -1 (1,2) #65
wire n669; //OPIN -1 (1,2) #66
wire n670; //OPIN -1 (1,2) #67
wire n671; //OPIN -1 (1,2) #68
wire n672; //OPIN -1 (1,2) #69
wire n673; //OPIN -1 (1,2) #70
wire n674; //OPIN -1 (1,2) #71
wire n675; //IPIN -1 (1,2) #72
wire n701; //IPIN -1 (1,3) #0
wire n702; //IPIN -1 (1,3) #1
wire n703; //IPIN -1 (1,3) #2
wire n704; //IPIN -1 (1,3) #3
wire n705; //IPIN -1 (1,3) #4
wire n706; //IPIN -1 (1,3) #5
wire n707; //IPIN -1 (1,3) #6
wire n708; //IPIN -1 (1,3) #7
wire n709; //IPIN -1 (1,3) #8
wire n710; //IPIN -1 (1,3) #9
wire n711; //IPIN -1 (1,3) #10
wire n712; //IPIN -1 (1,3) #11
wire n713; //IPIN -1 (1,3) #12
wire n714; //IPIN -1 (1,3) #13
wire n715; //IPIN -1 (1,3) #14
wire n716; //IPIN -1 (1,3) #15
wire n717; //IPIN -1 (1,3) #16
wire n718; //IPIN -1 (1,3) #17
wire n719; //IPIN -1 (1,3) #18
wire n720; //IPIN -1 (1,3) #19
wire n721; //IPIN -1 (1,3) #20
wire n722; //IPIN -1 (1,3) #21
wire n723; //IPIN -1 (1,3) #22
wire n724; //IPIN -1 (1,3) #23
wire n725; //IPIN -1 (1,3) #24
wire n726; //IPIN -1 (1,3) #25
wire n727; //IPIN -1 (1,3) #26
wire n728; //IPIN -1 (1,3) #27
wire n729; //IPIN -1 (1,3) #28
wire n730; //IPIN -1 (1,3) #29
wire n731; //IPIN -1 (1,3) #30
wire n732; //IPIN -1 (1,3) #31
wire n733; //IPIN -1 (1,3) #32
wire n734; //IPIN -1 (1,3) #33
wire n735; //IPIN -1 (1,3) #34
wire n736; //IPIN -1 (1,3) #35
wire n737; //IPIN -1 (1,3) #36
wire n738; //IPIN -1 (1,3) #37
wire n739; //IPIN -1 (1,3) #38
wire n740; //IPIN -1 (1,3) #39
wire n741; //IPIN -1 (1,3) #40
wire n742; //IPIN -1 (1,3) #41
wire n743; //IPIN -1 (1,3) #42
wire n744; //IPIN -1 (1,3) #43
wire n745; //IPIN -1 (1,3) #44
wire n746; //IPIN -1 (1,3) #45
wire n747; //IPIN -1 (1,3) #46
wire n748; //IPIN -1 (1,3) #47
wire n749; //IPIN -1 (1,3) #48
wire n750; //IPIN -1 (1,3) #49
wire n751; //IPIN -1 (1,3) #50
wire n752; //IPIN -1 (1,3) #51
wire n753; //OPIN -1 (1,3) #52
wire n754; //OPIN -1 (1,3) #53
wire n755; //OPIN -1 (1,3) #54
wire n756; //OPIN -1 (1,3) #55
wire n757; //OPIN -1 (1,3) #56
wire n758; //OPIN -1 (1,3) #57
wire n759; //OPIN -1 (1,3) #58
wire n760; //OPIN -1 (1,3) #59
wire n761; //OPIN -1 (1,3) #60
wire n762; //OPIN -1 (1,3) #61
wire n763; //OPIN -1 (1,3) #62
wire n764; //OPIN -1 (1,3) #63
wire n765; //OPIN -1 (1,3) #64
wire n766; //OPIN -1 (1,3) #65
wire n767; //OPIN -1 (1,3) #66
wire n768; //OPIN -1 (1,3) #67
wire n769; //OPIN -1 (1,3) #68
wire n770; //OPIN -1 (1,3) #69
wire n771; //OPIN -1 (1,3) #70
wire n772; //OPIN -1 (1,3) #71
wire n773; //IPIN -1 (1,3) #72
wire n799; //IPIN -1 (1,4) #0
wire n800; //IPIN -1 (1,4) #1
wire n801; //IPIN -1 (1,4) #2
wire n802; //IPIN -1 (1,4) #3
wire n803; //IPIN -1 (1,4) #4
wire n804; //IPIN -1 (1,4) #5
wire n805; //IPIN -1 (1,4) #6
wire n806; //IPIN -1 (1,4) #7
wire n807; //IPIN -1 (1,4) #8
wire n808; //IPIN -1 (1,4) #9
wire n809; //IPIN -1 (1,4) #10
wire n810; //IPIN -1 (1,4) #11
wire n811; //IPIN -1 (1,4) #12
wire n812; //IPIN -1 (1,4) #13
wire n813; //IPIN -1 (1,4) #14
wire n814; //IPIN -1 (1,4) #15
wire n815; //IPIN -1 (1,4) #16
wire n816; //IPIN -1 (1,4) #17
wire n817; //IPIN -1 (1,4) #18
wire n818; //IPIN -1 (1,4) #19
wire n819; //IPIN -1 (1,4) #20
wire n820; //IPIN -1 (1,4) #21
wire n821; //IPIN -1 (1,4) #22
wire n822; //IPIN -1 (1,4) #23
wire n823; //IPIN -1 (1,4) #24
wire n824; //IPIN -1 (1,4) #25
wire n825; //IPIN -1 (1,4) #26
wire n826; //IPIN -1 (1,4) #27
wire n827; //IPIN -1 (1,4) #28
wire n828; //IPIN -1 (1,4) #29
wire n829; //IPIN -1 (1,4) #30
wire n830; //IPIN -1 (1,4) #31
wire n831; //IPIN -1 (1,4) #32
wire n832; //IPIN -1 (1,4) #33
wire n833; //IPIN -1 (1,4) #34
wire n834; //IPIN -1 (1,4) #35
wire n835; //IPIN -1 (1,4) #36
wire n836; //IPIN -1 (1,4) #37
wire n837; //IPIN -1 (1,4) #38
wire n838; //IPIN -1 (1,4) #39
wire n839; //IPIN -1 (1,4) #40
wire n840; //IPIN -1 (1,4) #41
wire n841; //IPIN -1 (1,4) #42
wire n842; //IPIN -1 (1,4) #43
wire n843; //IPIN -1 (1,4) #44
wire n844; //IPIN -1 (1,4) #45
wire n845; //IPIN -1 (1,4) #46
wire n846; //IPIN -1 (1,4) #47
wire n847; //IPIN -1 (1,4) #48
wire n848; //IPIN -1 (1,4) #49
wire n849; //IPIN -1 (1,4) #50
wire n850; //IPIN -1 (1,4) #51
wire n851; //OPIN -1 (1,4) #52
wire n852; //OPIN -1 (1,4) #53
wire n853; //OPIN -1 (1,4) #54
wire n854; //OPIN -1 (1,4) #55
wire n855; //OPIN -1 (1,4) #56
wire n856; //OPIN -1 (1,4) #57
wire n857; //OPIN -1 (1,4) #58
wire n858; //OPIN -1 (1,4) #59
wire n859; //OPIN -1 (1,4) #60
wire n860; //OPIN -1 (1,4) #61
wire n861; //OPIN -1 (1,4) #62
wire n862; //OPIN -1 (1,4) #63
wire n863; //OPIN -1 (1,4) #64
wire n864; //OPIN -1 (1,4) #65
wire n865; //OPIN -1 (1,4) #66
wire n866; //OPIN -1 (1,4) #67
wire n867; //OPIN -1 (1,4) #68
wire n868; //OPIN -1 (1,4) #69
wire n869; //OPIN -1 (1,4) #70
wire n870; //OPIN -1 (1,4) #71
wire n871; //IPIN -1 (1,4) #72
wire n897; //IPIN -1 (1,5) #0
wire n898; //IPIN -1 (1,5) #1
wire n899; //IPIN -1 (1,5) #2
wire n900; //IPIN -1 (1,5) #3
wire n901; //IPIN -1 (1,5) #4
wire n902; //IPIN -1 (1,5) #5
wire n903; //IPIN -1 (1,5) #6
wire n904; //IPIN -1 (1,5) #7
wire n905; //IPIN -1 (1,5) #8
wire n906; //IPIN -1 (1,5) #9
wire n907; //IPIN -1 (1,5) #10
wire n908; //IPIN -1 (1,5) #11
wire n909; //IPIN -1 (1,5) #12
wire n910; //IPIN -1 (1,5) #13
wire n911; //IPIN -1 (1,5) #14
wire n912; //IPIN -1 (1,5) #15
wire n913; //IPIN -1 (1,5) #16
wire n914; //IPIN -1 (1,5) #17
wire n915; //IPIN -1 (1,5) #18
wire n916; //IPIN -1 (1,5) #19
wire n917; //IPIN -1 (1,5) #20
wire n918; //IPIN -1 (1,5) #21
wire n919; //IPIN -1 (1,5) #22
wire n920; //IPIN -1 (1,5) #23
wire n921; //IPIN -1 (1,5) #24
wire n922; //IPIN -1 (1,5) #25
wire n923; //IPIN -1 (1,5) #26
wire n924; //IPIN -1 (1,5) #27
wire n925; //IPIN -1 (1,5) #28
wire n926; //IPIN -1 (1,5) #29
wire n927; //IPIN -1 (1,5) #30
wire n928; //IPIN -1 (1,5) #31
wire n929; //IPIN -1 (1,5) #32
wire n930; //IPIN -1 (1,5) #33
wire n931; //IPIN -1 (1,5) #34
wire n932; //IPIN -1 (1,5) #35
wire n933; //IPIN -1 (1,5) #36
wire n934; //IPIN -1 (1,5) #37
wire n935; //IPIN -1 (1,5) #38
wire n936; //IPIN -1 (1,5) #39
wire n937; //IPIN -1 (1,5) #40
wire n938; //IPIN -1 (1,5) #41
wire n939; //IPIN -1 (1,5) #42
wire n940; //IPIN -1 (1,5) #43
wire n941; //IPIN -1 (1,5) #44
wire n942; //IPIN -1 (1,5) #45
wire n943; //IPIN -1 (1,5) #46
wire n944; //IPIN -1 (1,5) #47
wire n945; //IPIN -1 (1,5) #48
wire n946; //IPIN -1 (1,5) #49
wire n947; //IPIN -1 (1,5) #50
wire n948; //IPIN -1 (1,5) #51
wire n949; //OPIN -1 (1,5) #52
wire n950; //OPIN -1 (1,5) #53
wire n951; //OPIN -1 (1,5) #54
wire n952; //OPIN -1 (1,5) #55
wire n953; //OPIN -1 (1,5) #56
wire n954; //OPIN -1 (1,5) #57
wire n955; //OPIN -1 (1,5) #58
wire n956; //OPIN -1 (1,5) #59
wire n957; //OPIN -1 (1,5) #60
wire n958; //OPIN -1 (1,5) #61
wire n959; //OPIN -1 (1,5) #62
wire n960; //OPIN -1 (1,5) #63
wire n961; //OPIN -1 (1,5) #64
wire n962; //OPIN -1 (1,5) #65
wire n963; //OPIN -1 (1,5) #66
wire n964; //OPIN -1 (1,5) #67
wire n965; //OPIN -1 (1,5) #68
wire n966; //OPIN -1 (1,5) #69
wire n967; //OPIN -1 (1,5) #70
wire n968; //OPIN -1 (1,5) #71
wire n969; //IPIN -1 (1,5) #72
wire n995; //IPIN -1 (1,6) #0
wire n996; //IPIN -1 (1,6) #1
wire n997; //IPIN -1 (1,6) #2
wire n998; //IPIN -1 (1,6) #3
wire n999; //IPIN -1 (1,6) #4
wire n1000; //IPIN -1 (1,6) #5
wire n1001; //IPIN -1 (1,6) #6
wire n1002; //IPIN -1 (1,6) #7
wire n1003; //IPIN -1 (1,6) #8
wire n1004; //IPIN -1 (1,6) #9
wire n1005; //IPIN -1 (1,6) #10
wire n1006; //IPIN -1 (1,6) #11
wire n1007; //IPIN -1 (1,6) #12
wire n1008; //IPIN -1 (1,6) #13
wire n1009; //IPIN -1 (1,6) #14
wire n1010; //IPIN -1 (1,6) #15
wire n1011; //IPIN -1 (1,6) #16
wire n1012; //IPIN -1 (1,6) #17
wire n1013; //IPIN -1 (1,6) #18
wire n1014; //IPIN -1 (1,6) #19
wire n1015; //IPIN -1 (1,6) #20
wire n1016; //IPIN -1 (1,6) #21
wire n1017; //IPIN -1 (1,6) #22
wire n1018; //IPIN -1 (1,6) #23
wire n1019; //IPIN -1 (1,6) #24
wire n1020; //IPIN -1 (1,6) #25
wire n1021; //IPIN -1 (1,6) #26
wire n1022; //IPIN -1 (1,6) #27
wire n1023; //IPIN -1 (1,6) #28
wire n1024; //IPIN -1 (1,6) #29
wire n1025; //IPIN -1 (1,6) #30
wire n1026; //IPIN -1 (1,6) #31
wire n1027; //IPIN -1 (1,6) #32
wire n1028; //IPIN -1 (1,6) #33
wire n1029; //IPIN -1 (1,6) #34
wire n1030; //IPIN -1 (1,6) #35
wire n1031; //IPIN -1 (1,6) #36
wire n1032; //IPIN -1 (1,6) #37
wire n1033; //IPIN -1 (1,6) #38
wire n1034; //IPIN -1 (1,6) #39
wire n1035; //IPIN -1 (1,6) #40
wire n1036; //IPIN -1 (1,6) #41
wire n1037; //IPIN -1 (1,6) #42
wire n1038; //IPIN -1 (1,6) #43
wire n1039; //IPIN -1 (1,6) #44
wire n1040; //IPIN -1 (1,6) #45
wire n1041; //IPIN -1 (1,6) #46
wire n1042; //IPIN -1 (1,6) #47
wire n1043; //IPIN -1 (1,6) #48
wire n1044; //IPIN -1 (1,6) #49
wire n1045; //IPIN -1 (1,6) #50
wire n1046; //IPIN -1 (1,6) #51
wire n1047; //OPIN -1 (1,6) #52
wire n1048; //OPIN -1 (1,6) #53
wire n1049; //OPIN -1 (1,6) #54
wire n1050; //OPIN -1 (1,6) #55
wire n1051; //OPIN -1 (1,6) #56
wire n1052; //OPIN -1 (1,6) #57
wire n1053; //OPIN -1 (1,6) #58
wire n1054; //OPIN -1 (1,6) #59
wire n1055; //OPIN -1 (1,6) #60
wire n1056; //OPIN -1 (1,6) #61
wire n1057; //OPIN -1 (1,6) #62
wire n1058; //OPIN -1 (1,6) #63
wire n1059; //OPIN -1 (1,6) #64
wire n1060; //OPIN -1 (1,6) #65
wire n1061; //OPIN -1 (1,6) #66
wire n1062; //OPIN -1 (1,6) #67
wire n1063; //OPIN -1 (1,6) #68
wire n1064; //OPIN -1 (1,6) #69
wire n1065; //OPIN -1 (1,6) #70
wire n1066; //OPIN -1 (1,6) #71
wire n1067; //IPIN -1 (1,6) #72
wire n1093; //IPIN -1 (1,7) #0
wire n1094; //IPIN -1 (1,7) #1
wire n1095; //IPIN -1 (1,7) #2
wire n1096; //IPIN -1 (1,7) #3
wire n1097; //IPIN -1 (1,7) #4
wire n1098; //IPIN -1 (1,7) #5
wire n1099; //IPIN -1 (1,7) #6
wire n1100; //IPIN -1 (1,7) #7
wire n1101; //IPIN -1 (1,7) #8
wire n1102; //IPIN -1 (1,7) #9
wire n1103; //IPIN -1 (1,7) #10
wire n1104; //IPIN -1 (1,7) #11
wire n1105; //IPIN -1 (1,7) #12
wire n1106; //IPIN -1 (1,7) #13
wire n1107; //IPIN -1 (1,7) #14
wire n1108; //IPIN -1 (1,7) #15
wire n1109; //IPIN -1 (1,7) #16
wire n1110; //IPIN -1 (1,7) #17
wire n1111; //IPIN -1 (1,7) #18
wire n1112; //IPIN -1 (1,7) #19
wire n1113; //IPIN -1 (1,7) #20
wire n1114; //IPIN -1 (1,7) #21
wire n1115; //IPIN -1 (1,7) #22
wire n1116; //IPIN -1 (1,7) #23
wire n1117; //IPIN -1 (1,7) #24
wire n1118; //IPIN -1 (1,7) #25
wire n1119; //IPIN -1 (1,7) #26
wire n1120; //IPIN -1 (1,7) #27
wire n1121; //IPIN -1 (1,7) #28
wire n1122; //IPIN -1 (1,7) #29
wire n1123; //IPIN -1 (1,7) #30
wire n1124; //IPIN -1 (1,7) #31
wire n1125; //IPIN -1 (1,7) #32
wire n1126; //IPIN -1 (1,7) #33
wire n1127; //IPIN -1 (1,7) #34
wire n1128; //IPIN -1 (1,7) #35
wire n1129; //IPIN -1 (1,7) #36
wire n1130; //IPIN -1 (1,7) #37
wire n1131; //IPIN -1 (1,7) #38
wire n1132; //IPIN -1 (1,7) #39
wire n1133; //IPIN -1 (1,7) #40
wire n1134; //IPIN -1 (1,7) #41
wire n1135; //IPIN -1 (1,7) #42
wire n1136; //IPIN -1 (1,7) #43
wire n1137; //IPIN -1 (1,7) #44
wire n1138; //IPIN -1 (1,7) #45
wire n1139; //IPIN -1 (1,7) #46
wire n1140; //IPIN -1 (1,7) #47
wire n1141; //IPIN -1 (1,7) #48
wire n1142; //IPIN -1 (1,7) #49
wire n1143; //IPIN -1 (1,7) #50
wire n1144; //IPIN -1 (1,7) #51
wire n1145; //OPIN -1 (1,7) #52
wire n1146; //OPIN -1 (1,7) #53
wire n1147; //OPIN -1 (1,7) #54
wire n1148; //OPIN -1 (1,7) #55
wire n1149; //OPIN -1 (1,7) #56
wire n1150; //OPIN -1 (1,7) #57
wire n1151; //OPIN -1 (1,7) #58
wire n1152; //OPIN -1 (1,7) #59
wire n1153; //OPIN -1 (1,7) #60
wire n1154; //OPIN -1 (1,7) #61
wire n1155; //OPIN -1 (1,7) #62
wire n1156; //OPIN -1 (1,7) #63
wire n1157; //OPIN -1 (1,7) #64
wire n1158; //OPIN -1 (1,7) #65
wire n1159; //OPIN -1 (1,7) #66
wire n1160; //OPIN -1 (1,7) #67
wire n1161; //OPIN -1 (1,7) #68
wire n1162; //OPIN -1 (1,7) #69
wire n1163; //OPIN -1 (1,7) #70
wire n1164; //OPIN -1 (1,7) #71
wire n1165; //IPIN -1 (1,7) #72
wire n1191; //IPIN -1 (1,8) #0
wire n1192; //IPIN -1 (1,8) #1
wire n1193; //IPIN -1 (1,8) #2
wire n1194; //IPIN -1 (1,8) #3
wire n1195; //IPIN -1 (1,8) #4
wire n1196; //IPIN -1 (1,8) #5
wire n1197; //IPIN -1 (1,8) #6
wire n1198; //IPIN -1 (1,8) #7
wire n1199; //IPIN -1 (1,8) #8
wire n1200; //IPIN -1 (1,8) #9
wire n1201; //IPIN -1 (1,8) #10
wire n1202; //IPIN -1 (1,8) #11
wire n1203; //IPIN -1 (1,8) #12
wire n1204; //IPIN -1 (1,8) #13
wire n1205; //IPIN -1 (1,8) #14
wire n1206; //IPIN -1 (1,8) #15
wire n1207; //IPIN -1 (1,8) #16
wire n1208; //IPIN -1 (1,8) #17
wire n1209; //IPIN -1 (1,8) #18
wire n1210; //IPIN -1 (1,8) #19
wire n1211; //IPIN -1 (1,8) #20
wire n1212; //IPIN -1 (1,8) #21
wire n1213; //IPIN -1 (1,8) #22
wire n1214; //IPIN -1 (1,8) #23
wire n1215; //IPIN -1 (1,8) #24
wire n1216; //IPIN -1 (1,8) #25
wire n1217; //IPIN -1 (1,8) #26
wire n1218; //IPIN -1 (1,8) #27
wire n1219; //IPIN -1 (1,8) #28
wire n1220; //IPIN -1 (1,8) #29
wire n1221; //IPIN -1 (1,8) #30
wire n1222; //IPIN -1 (1,8) #31
wire n1223; //IPIN -1 (1,8) #32
wire n1224; //IPIN -1 (1,8) #33
wire n1225; //IPIN -1 (1,8) #34
wire n1226; //IPIN -1 (1,8) #35
wire n1227; //IPIN -1 (1,8) #36
wire n1228; //IPIN -1 (1,8) #37
wire n1229; //IPIN -1 (1,8) #38
wire n1230; //IPIN -1 (1,8) #39
wire n1231; //IPIN -1 (1,8) #40
wire n1232; //IPIN -1 (1,8) #41
wire n1233; //IPIN -1 (1,8) #42
wire n1234; //IPIN -1 (1,8) #43
wire n1235; //IPIN -1 (1,8) #44
wire n1236; //IPIN -1 (1,8) #45
wire n1237; //IPIN -1 (1,8) #46
wire n1238; //IPIN -1 (1,8) #47
wire n1239; //IPIN -1 (1,8) #48
wire n1240; //IPIN -1 (1,8) #49
wire n1241; //IPIN -1 (1,8) #50
wire n1242; //IPIN -1 (1,8) #51
wire n1243; //OPIN -1 (1,8) #52
wire n1244; //OPIN -1 (1,8) #53
wire n1245; //OPIN -1 (1,8) #54
wire n1246; //OPIN -1 (1,8) #55
wire n1247; //OPIN -1 (1,8) #56
wire n1248; //OPIN -1 (1,8) #57
wire n1249; //OPIN -1 (1,8) #58
wire n1250; //OPIN -1 (1,8) #59
wire n1251; //OPIN -1 (1,8) #60
wire n1252; //OPIN -1 (1,8) #61
wire n1253; //OPIN -1 (1,8) #62
wire n1254; //OPIN -1 (1,8) #63
wire n1255; //OPIN -1 (1,8) #64
wire n1256; //OPIN -1 (1,8) #65
wire n1257; //OPIN -1 (1,8) #66
wire n1258; //OPIN -1 (1,8) #67
wire n1259; //OPIN -1 (1,8) #68
wire n1260; //OPIN -1 (1,8) #69
wire n1261; //OPIN -1 (1,8) #70
wire n1262; //OPIN -1 (1,8) #71
wire n1263; //IPIN -1 (1,8) #72
wire n1289; //IPIN -1 (1,9) #0
wire n1290; //IPIN -1 (1,9) #1
wire n1291; //IPIN -1 (1,9) #2
wire n1292; //IPIN -1 (1,9) #3
wire n1293; //IPIN -1 (1,9) #4
wire n1294; //IPIN -1 (1,9) #5
wire n1295; //IPIN -1 (1,9) #6
wire n1296; //IPIN -1 (1,9) #7
wire n1297; //IPIN -1 (1,9) #8
wire n1298; //IPIN -1 (1,9) #9
wire n1299; //IPIN -1 (1,9) #10
wire n1300; //IPIN -1 (1,9) #11
wire n1301; //IPIN -1 (1,9) #12
wire n1302; //IPIN -1 (1,9) #13
wire n1303; //IPIN -1 (1,9) #14
wire n1304; //IPIN -1 (1,9) #15
wire n1305; //IPIN -1 (1,9) #16
wire n1306; //IPIN -1 (1,9) #17
wire n1307; //IPIN -1 (1,9) #18
wire n1308; //IPIN -1 (1,9) #19
wire n1309; //IPIN -1 (1,9) #20
wire n1310; //IPIN -1 (1,9) #21
wire n1311; //IPIN -1 (1,9) #22
wire n1312; //IPIN -1 (1,9) #23
wire n1313; //IPIN -1 (1,9) #24
wire n1314; //IPIN -1 (1,9) #25
wire n1315; //IPIN -1 (1,9) #26
wire n1316; //IPIN -1 (1,9) #27
wire n1317; //IPIN -1 (1,9) #28
wire n1318; //IPIN -1 (1,9) #29
wire n1319; //IPIN -1 (1,9) #30
wire n1320; //IPIN -1 (1,9) #31
wire n1321; //IPIN -1 (1,9) #32
wire n1322; //IPIN -1 (1,9) #33
wire n1323; //IPIN -1 (1,9) #34
wire n1324; //IPIN -1 (1,9) #35
wire n1325; //IPIN -1 (1,9) #36
wire n1326; //IPIN -1 (1,9) #37
wire n1327; //IPIN -1 (1,9) #38
wire n1328; //IPIN -1 (1,9) #39
wire n1329; //IPIN -1 (1,9) #40
wire n1330; //IPIN -1 (1,9) #41
wire n1331; //IPIN -1 (1,9) #42
wire n1332; //IPIN -1 (1,9) #43
wire n1333; //IPIN -1 (1,9) #44
wire n1334; //IPIN -1 (1,9) #45
wire n1335; //IPIN -1 (1,9) #46
wire n1336; //IPIN -1 (1,9) #47
wire n1337; //IPIN -1 (1,9) #48
wire n1338; //IPIN -1 (1,9) #49
wire n1339; //IPIN -1 (1,9) #50
wire n1340; //IPIN -1 (1,9) #51
wire n1341; //OPIN -1 (1,9) #52
wire n1342; //OPIN -1 (1,9) #53
wire n1343; //OPIN -1 (1,9) #54
wire n1344; //OPIN -1 (1,9) #55
wire n1345; //OPIN -1 (1,9) #56
wire n1346; //OPIN -1 (1,9) #57
wire n1347; //OPIN -1 (1,9) #58
wire n1348; //OPIN -1 (1,9) #59
wire n1349; //OPIN -1 (1,9) #60
wire n1350; //OPIN -1 (1,9) #61
wire n1351; //OPIN -1 (1,9) #62
wire n1352; //OPIN -1 (1,9) #63
wire n1353; //OPIN -1 (1,9) #64
wire n1354; //OPIN -1 (1,9) #65
wire n1355; //OPIN -1 (1,9) #66
wire n1356; //OPIN -1 (1,9) #67
wire n1357; //OPIN -1 (1,9) #68
wire n1358; //OPIN -1 (1,9) #69
wire n1359; //OPIN -1 (1,9) #70
wire n1360; //OPIN -1 (1,9) #71
wire n1361; //IPIN -1 (1,9) #72
wire n1386; //IPIN -1 (1,10) #0
wire n1387; //OPIN -1 (1,10) #1
wire n1388; //IPIN -1 (1,10) #2
wire n1389; //IPIN -1 (1,10) #3
wire n1390; //OPIN -1 (1,10) #4
wire n1391; //IPIN -1 (1,10) #5
wire n1392; //IPIN -1 (1,10) #6
wire n1393; //OPIN -1 (1,10) #7
wire n1394; //IPIN -1 (1,10) #8
wire n1395; //IPIN -1 (1,10) #9
wire n1396; //OPIN -1 (1,10) #10
wire n1397; //IPIN -1 (1,10) #11
wire n1398; //IPIN -1 (1,10) #12
wire n1399; //OPIN -1 (1,10) #13
wire n1400; //IPIN -1 (1,10) #14
wire n1401; //IPIN -1 (1,10) #15
wire n1402; //OPIN -1 (1,10) #16
wire n1403; //IPIN -1 (1,10) #17
wire n1404; //IPIN -1 (1,10) #18
wire n1405; //OPIN -1 (1,10) #19
wire n1406; //IPIN -1 (1,10) #20
wire n1407; //IPIN -1 (1,10) #21
wire n1408; //OPIN -1 (1,10) #22
wire n1409; //IPIN -1 (1,10) #23
wire n1434; //IPIN -1 (2,0) #0
wire n1435; //OPIN -1 (2,0) #1
wire n1436; //IPIN -1 (2,0) #2
wire n1437; //IPIN -1 (2,0) #3
wire n1438; //OPIN -1 (2,0) #4
wire n1439; //IPIN -1 (2,0) #5
wire n1440; //IPIN -1 (2,0) #6
wire n1441; //OPIN -1 (2,0) #7
wire n1442; //IPIN -1 (2,0) #8
wire n1443; //IPIN -1 (2,0) #9
wire n1444; //OPIN -1 (2,0) #10
wire n1445; //IPIN -1 (2,0) #11
wire n1446; //IPIN -1 (2,0) #12
wire n1447; //OPIN -1 (2,0) #13
wire n1448; //IPIN -1 (2,0) #14
wire n1449; //IPIN -1 (2,0) #15
wire n1450; //OPIN -1 (2,0) #16
wire n1451; //IPIN -1 (2,0) #17
wire n1452; //IPIN -1 (2,0) #18
wire n1453; //OPIN -1 (2,0) #19
wire n1454; //IPIN -1 (2,0) #20
wire n1455; //IPIN -1 (2,0) #21
wire n1456; //OPIN -1 (2,0) #22
wire n1457; //IPIN -1 (2,0) #23
wire n1483; //IPIN -1 (2,1) #0
wire n1484; //IPIN -1 (2,1) #1
wire n1485; //IPIN -1 (2,1) #2
wire n1486; //IPIN -1 (2,1) #3
wire n1487; //IPIN -1 (2,1) #4
wire n1488; //IPIN -1 (2,1) #5
wire n1489; //IPIN -1 (2,1) #6
wire n1490; //IPIN -1 (2,1) #7
wire n1491; //IPIN -1 (2,1) #8
wire n1492; //IPIN -1 (2,1) #9
wire n1493; //IPIN -1 (2,1) #10
wire n1494; //IPIN -1 (2,1) #11
wire n1495; //IPIN -1 (2,1) #12
wire n1496; //IPIN -1 (2,1) #13
wire n1497; //IPIN -1 (2,1) #14
wire n1498; //IPIN -1 (2,1) #15
wire n1499; //IPIN -1 (2,1) #16
wire n1500; //IPIN -1 (2,1) #17
wire n1501; //IPIN -1 (2,1) #18
wire n1502; //IPIN -1 (2,1) #19
wire n1503; //IPIN -1 (2,1) #20
wire n1504; //IPIN -1 (2,1) #21
wire n1505; //IPIN -1 (2,1) #22
wire n1506; //IPIN -1 (2,1) #23
wire n1507; //IPIN -1 (2,1) #24
wire n1508; //IPIN -1 (2,1) #25
wire n1509; //IPIN -1 (2,1) #26
wire n1510; //IPIN -1 (2,1) #27
wire n1511; //IPIN -1 (2,1) #28
wire n1512; //IPIN -1 (2,1) #29
wire n1513; //IPIN -1 (2,1) #30
wire n1514; //IPIN -1 (2,1) #31
wire n1515; //IPIN -1 (2,1) #32
wire n1516; //IPIN -1 (2,1) #33
wire n1517; //IPIN -1 (2,1) #34
wire n1518; //IPIN -1 (2,1) #35
wire n1519; //IPIN -1 (2,1) #36
wire n1520; //IPIN -1 (2,1) #37
wire n1521; //IPIN -1 (2,1) #38
wire n1522; //IPIN -1 (2,1) #39
wire n1523; //IPIN -1 (2,1) #40
wire n1524; //IPIN -1 (2,1) #41
wire n1525; //IPIN -1 (2,1) #42
wire n1526; //IPIN -1 (2,1) #43
wire n1527; //IPIN -1 (2,1) #44
wire n1528; //IPIN -1 (2,1) #45
wire n1529; //IPIN -1 (2,1) #46
wire n1530; //IPIN -1 (2,1) #47
wire n1531; //IPIN -1 (2,1) #48
wire n1532; //IPIN -1 (2,1) #49
wire n1533; //IPIN -1 (2,1) #50
wire n1534; //IPIN -1 (2,1) #51
wire n1535; //OPIN -1 (2,1) #52
wire n1536; //OPIN -1 (2,1) #53
wire n1537; //OPIN -1 (2,1) #54
wire n1538; //OPIN -1 (2,1) #55
wire n1539; //OPIN -1 (2,1) #56
wire n1540; //OPIN -1 (2,1) #57
wire n1541; //OPIN -1 (2,1) #58
wire n1542; //OPIN -1 (2,1) #59
wire n1543; //OPIN -1 (2,1) #60
wire n1544; //OPIN -1 (2,1) #61
wire n1545; //OPIN -1 (2,1) #62
wire n1546; //OPIN -1 (2,1) #63
wire n1547; //OPIN -1 (2,1) #64
wire n1548; //OPIN -1 (2,1) #65
wire n1549; //OPIN -1 (2,1) #66
wire n1550; //OPIN -1 (2,1) #67
wire n1551; //OPIN -1 (2,1) #68
wire n1552; //OPIN -1 (2,1) #69
wire n1553; //OPIN -1 (2,1) #70
wire n1554; //OPIN -1 (2,1) #71
wire n1555; //IPIN -1 (2,1) #72
wire n1581; //IPIN -1 (2,2) #0
wire n1582; //IPIN -1 (2,2) #1
wire n1583; //IPIN -1 (2,2) #2
wire n1584; //IPIN -1 (2,2) #3
wire n1585; //IPIN -1 (2,2) #4
wire n1586; //IPIN -1 (2,2) #5
wire n1587; //IPIN -1 (2,2) #6
wire n1588; //IPIN -1 (2,2) #7
wire n1589; //IPIN -1 (2,2) #8
wire n1590; //IPIN -1 (2,2) #9
wire n1591; //IPIN -1 (2,2) #10
wire n1592; //IPIN -1 (2,2) #11
wire n1593; //IPIN -1 (2,2) #12
wire n1594; //IPIN -1 (2,2) #13
wire n1595; //IPIN -1 (2,2) #14
wire n1596; //IPIN -1 (2,2) #15
wire n1597; //IPIN -1 (2,2) #16
wire n1598; //IPIN -1 (2,2) #17
wire n1599; //IPIN -1 (2,2) #18
wire n1600; //IPIN -1 (2,2) #19
wire n1601; //IPIN -1 (2,2) #20
wire n1602; //IPIN -1 (2,2) #21
wire n1603; //IPIN -1 (2,2) #22
wire n1604; //IPIN -1 (2,2) #23
wire n1605; //IPIN -1 (2,2) #24
wire n1606; //IPIN -1 (2,2) #25
wire n1607; //IPIN -1 (2,2) #26
wire n1608; //IPIN -1 (2,2) #27
wire n1609; //IPIN -1 (2,2) #28
wire n1610; //IPIN -1 (2,2) #29
wire n1611; //IPIN -1 (2,2) #30
wire n1612; //IPIN -1 (2,2) #31
wire n1613; //IPIN -1 (2,2) #32
wire n1614; //IPIN -1 (2,2) #33
wire n1615; //IPIN -1 (2,2) #34
wire n1616; //IPIN -1 (2,2) #35
wire n1617; //IPIN -1 (2,2) #36
wire n1618; //IPIN -1 (2,2) #37
wire n1619; //IPIN -1 (2,2) #38
wire n1620; //IPIN -1 (2,2) #39
wire n1621; //IPIN -1 (2,2) #40
wire n1622; //IPIN -1 (2,2) #41
wire n1623; //IPIN -1 (2,2) #42
wire n1624; //IPIN -1 (2,2) #43
wire n1625; //IPIN -1 (2,2) #44
wire n1626; //IPIN -1 (2,2) #45
wire n1627; //IPIN -1 (2,2) #46
wire n1628; //IPIN -1 (2,2) #47
wire n1629; //IPIN -1 (2,2) #48
wire n1630; //IPIN -1 (2,2) #49
wire n1631; //IPIN -1 (2,2) #50
wire n1632; //IPIN -1 (2,2) #51
wire n1633; //OPIN -1 (2,2) #52
wire n1634; //OPIN -1 (2,2) #53
wire n1635; //OPIN -1 (2,2) #54
wire n1636; //OPIN -1 (2,2) #55
wire n1637; //OPIN -1 (2,2) #56
wire n1638; //OPIN -1 (2,2) #57
wire n1639; //OPIN -1 (2,2) #58
wire n1640; //OPIN -1 (2,2) #59
wire n1641; //OPIN -1 (2,2) #60
wire n1642; //OPIN -1 (2,2) #61
wire n1643; //OPIN -1 (2,2) #62
wire n1644; //OPIN -1 (2,2) #63
wire n1645; //OPIN -1 (2,2) #64
wire n1646; //OPIN -1 (2,2) #65
wire n1647; //OPIN -1 (2,2) #66
wire n1648; //OPIN -1 (2,2) #67
wire n1649; //OPIN -1 (2,2) #68
wire n1650; //OPIN -1 (2,2) #69
wire n1651; //OPIN -1 (2,2) #70
wire n1652; //OPIN -1 (2,2) #71
wire n1653; //IPIN -1 (2,2) #72
wire n1679; //IPIN -1 (2,3) #0
wire n1680; //IPIN -1 (2,3) #1
wire n1681; //IPIN -1 (2,3) #2
wire n1682; //IPIN -1 (2,3) #3
wire n1683; //IPIN -1 (2,3) #4
wire n1684; //IPIN -1 (2,3) #5
wire n1685; //IPIN -1 (2,3) #6
wire n1686; //IPIN -1 (2,3) #7
wire n1687; //IPIN -1 (2,3) #8
wire n1688; //IPIN -1 (2,3) #9
wire n1689; //IPIN -1 (2,3) #10
wire n1690; //IPIN -1 (2,3) #11
wire n1691; //IPIN -1 (2,3) #12
wire n1692; //IPIN -1 (2,3) #13
wire n1693; //IPIN -1 (2,3) #14
wire n1694; //IPIN -1 (2,3) #15
wire n1695; //IPIN -1 (2,3) #16
wire n1696; //IPIN -1 (2,3) #17
wire n1697; //IPIN -1 (2,3) #18
wire n1698; //IPIN -1 (2,3) #19
wire n1699; //IPIN -1 (2,3) #20
wire n1700; //IPIN -1 (2,3) #21
wire n1701; //IPIN -1 (2,3) #22
wire n1702; //IPIN -1 (2,3) #23
wire n1703; //IPIN -1 (2,3) #24
wire n1704; //IPIN -1 (2,3) #25
wire n1705; //IPIN -1 (2,3) #26
wire n1706; //IPIN -1 (2,3) #27
wire n1707; //IPIN -1 (2,3) #28
wire n1708; //IPIN -1 (2,3) #29
wire n1709; //IPIN -1 (2,3) #30
wire n1710; //IPIN -1 (2,3) #31
wire n1711; //IPIN -1 (2,3) #32
wire n1712; //IPIN -1 (2,3) #33
wire n1713; //IPIN -1 (2,3) #34
wire n1714; //IPIN -1 (2,3) #35
wire n1715; //IPIN -1 (2,3) #36
wire n1716; //IPIN -1 (2,3) #37
wire n1717; //IPIN -1 (2,3) #38
wire n1718; //IPIN -1 (2,3) #39
wire n1719; //IPIN -1 (2,3) #40
wire n1720; //IPIN -1 (2,3) #41
wire n1721; //IPIN -1 (2,3) #42
wire n1722; //IPIN -1 (2,3) #43
wire n1723; //IPIN -1 (2,3) #44
wire n1724; //IPIN -1 (2,3) #45
wire n1725; //IPIN -1 (2,3) #46
wire n1726; //IPIN -1 (2,3) #47
wire n1727; //IPIN -1 (2,3) #48
wire n1728; //IPIN -1 (2,3) #49
wire n1729; //IPIN -1 (2,3) #50
wire n1730; //IPIN -1 (2,3) #51
wire n1731; //OPIN -1 (2,3) #52
wire n1732; //OPIN -1 (2,3) #53
wire n1733; //OPIN -1 (2,3) #54
wire n1734; //OPIN -1 (2,3) #55
wire n1735; //OPIN -1 (2,3) #56
wire n1736; //OPIN -1 (2,3) #57
wire n1737; //OPIN -1 (2,3) #58
wire n1738; //OPIN -1 (2,3) #59
wire n1739; //OPIN -1 (2,3) #60
wire n1740; //OPIN -1 (2,3) #61
wire n1741; //OPIN -1 (2,3) #62
wire n1742; //OPIN -1 (2,3) #63
wire n1743; //OPIN -1 (2,3) #64
wire n1744; //OPIN -1 (2,3) #65
wire n1745; //OPIN -1 (2,3) #66
wire n1746; //OPIN -1 (2,3) #67
wire n1747; //OPIN -1 (2,3) #68
wire n1748; //OPIN -1 (2,3) #69
wire n1749; //OPIN -1 (2,3) #70
wire n1750; //OPIN -1 (2,3) #71
wire n1751; //IPIN -1 (2,3) #72
wire n1777; //IPIN -1 (2,4) #0
wire n1778; //IPIN -1 (2,4) #1
wire n1779; //IPIN -1 (2,4) #2
wire n1780; //IPIN -1 (2,4) #3
wire n1781; //IPIN -1 (2,4) #4
wire n1782; //IPIN -1 (2,4) #5
wire n1783; //IPIN -1 (2,4) #6
wire n1784; //IPIN -1 (2,4) #7
wire n1785; //IPIN -1 (2,4) #8
wire n1786; //IPIN -1 (2,4) #9
wire n1787; //IPIN -1 (2,4) #10
wire n1788; //IPIN -1 (2,4) #11
wire n1789; //IPIN -1 (2,4) #12
wire n1790; //IPIN -1 (2,4) #13
wire n1791; //IPIN -1 (2,4) #14
wire n1792; //IPIN -1 (2,4) #15
wire n1793; //IPIN -1 (2,4) #16
wire n1794; //IPIN -1 (2,4) #17
wire n1795; //IPIN -1 (2,4) #18
wire n1796; //IPIN -1 (2,4) #19
wire n1797; //IPIN -1 (2,4) #20
wire n1798; //IPIN -1 (2,4) #21
wire n1799; //IPIN -1 (2,4) #22
wire n1800; //IPIN -1 (2,4) #23
wire n1801; //IPIN -1 (2,4) #24
wire n1802; //IPIN -1 (2,4) #25
wire n1803; //IPIN -1 (2,4) #26
wire n1804; //IPIN -1 (2,4) #27
wire n1805; //IPIN -1 (2,4) #28
wire n1806; //IPIN -1 (2,4) #29
wire n1807; //IPIN -1 (2,4) #30
wire n1808; //IPIN -1 (2,4) #31
wire n1809; //IPIN -1 (2,4) #32
wire n1810; //IPIN -1 (2,4) #33
wire n1811; //IPIN -1 (2,4) #34
wire n1812; //IPIN -1 (2,4) #35
wire n1813; //IPIN -1 (2,4) #36
wire n1814; //IPIN -1 (2,4) #37
wire n1815; //IPIN -1 (2,4) #38
wire n1816; //IPIN -1 (2,4) #39
wire n1817; //IPIN -1 (2,4) #40
wire n1818; //IPIN -1 (2,4) #41
wire n1819; //IPIN -1 (2,4) #42
wire n1820; //IPIN -1 (2,4) #43
wire n1821; //IPIN -1 (2,4) #44
wire n1822; //IPIN -1 (2,4) #45
wire n1823; //IPIN -1 (2,4) #46
wire n1824; //IPIN -1 (2,4) #47
wire n1825; //IPIN -1 (2,4) #48
wire n1826; //IPIN -1 (2,4) #49
wire n1827; //IPIN -1 (2,4) #50
wire n1828; //IPIN -1 (2,4) #51
wire n1829; //OPIN -1 (2,4) #52
wire n1830; //OPIN -1 (2,4) #53
wire n1831; //OPIN -1 (2,4) #54
wire n1832; //OPIN -1 (2,4) #55
wire n1833; //OPIN -1 (2,4) #56
wire n1834; //OPIN -1 (2,4) #57
wire n1835; //OPIN -1 (2,4) #58
wire n1836; //OPIN -1 (2,4) #59
wire n1837; //OPIN -1 (2,4) #60
wire n1838; //OPIN -1 (2,4) #61
wire n1839; //OPIN -1 (2,4) #62
wire n1840; //OPIN -1 (2,4) #63
wire n1841; //OPIN -1 (2,4) #64
wire n1842; //OPIN -1 (2,4) #65
wire n1843; //OPIN -1 (2,4) #66
wire n1844; //OPIN -1 (2,4) #67
wire n1845; //OPIN -1 (2,4) #68
wire n1846; //OPIN -1 (2,4) #69
wire n1847; //OPIN -1 (2,4) #70
wire n1848; //OPIN -1 (2,4) #71
wire n1849; //IPIN -1 (2,4) #72
wire n1875; //IPIN -1 (2,5) #0
wire n1876; //IPIN -1 (2,5) #1
wire n1877; //IPIN -1 (2,5) #2
wire n1878; //IPIN -1 (2,5) #3
wire n1879; //IPIN -1 (2,5) #4
wire n1880; //IPIN -1 (2,5) #5
wire n1881; //IPIN -1 (2,5) #6
wire n1882; //IPIN -1 (2,5) #7
wire n1883; //IPIN -1 (2,5) #8
wire n1884; //IPIN -1 (2,5) #9
wire n1885; //IPIN -1 (2,5) #10
wire n1886; //IPIN -1 (2,5) #11
wire n1887; //IPIN -1 (2,5) #12
wire n1888; //IPIN -1 (2,5) #13
wire n1889; //IPIN -1 (2,5) #14
wire n1890; //IPIN -1 (2,5) #15
wire n1891; //IPIN -1 (2,5) #16
wire n1892; //IPIN -1 (2,5) #17
wire n1893; //IPIN -1 (2,5) #18
wire n1894; //IPIN -1 (2,5) #19
wire n1895; //IPIN -1 (2,5) #20
wire n1896; //IPIN -1 (2,5) #21
wire n1897; //IPIN -1 (2,5) #22
wire n1898; //IPIN -1 (2,5) #23
wire n1899; //IPIN -1 (2,5) #24
wire n1900; //IPIN -1 (2,5) #25
wire n1901; //IPIN -1 (2,5) #26
wire n1902; //IPIN -1 (2,5) #27
wire n1903; //IPIN -1 (2,5) #28
wire n1904; //IPIN -1 (2,5) #29
wire n1905; //IPIN -1 (2,5) #30
wire n1906; //IPIN -1 (2,5) #31
wire n1907; //IPIN -1 (2,5) #32
wire n1908; //IPIN -1 (2,5) #33
wire n1909; //IPIN -1 (2,5) #34
wire n1910; //IPIN -1 (2,5) #35
wire n1911; //IPIN -1 (2,5) #36
wire n1912; //IPIN -1 (2,5) #37
wire n1913; //IPIN -1 (2,5) #38
wire n1914; //IPIN -1 (2,5) #39
wire n1915; //IPIN -1 (2,5) #40
wire n1916; //IPIN -1 (2,5) #41
wire n1917; //IPIN -1 (2,5) #42
wire n1918; //IPIN -1 (2,5) #43
wire n1919; //IPIN -1 (2,5) #44
wire n1920; //IPIN -1 (2,5) #45
wire n1921; //IPIN -1 (2,5) #46
wire n1922; //IPIN -1 (2,5) #47
wire n1923; //IPIN -1 (2,5) #48
wire n1924; //IPIN -1 (2,5) #49
wire n1925; //IPIN -1 (2,5) #50
wire n1926; //IPIN -1 (2,5) #51
wire n1927; //OPIN -1 (2,5) #52
wire n1928; //OPIN -1 (2,5) #53
wire n1929; //OPIN -1 (2,5) #54
wire n1930; //OPIN -1 (2,5) #55
wire n1931; //OPIN -1 (2,5) #56
wire n1932; //OPIN -1 (2,5) #57
wire n1933; //OPIN -1 (2,5) #58
wire n1934; //OPIN -1 (2,5) #59
wire n1935; //OPIN -1 (2,5) #60
wire n1936; //OPIN -1 (2,5) #61
wire n1937; //OPIN -1 (2,5) #62
wire n1938; //OPIN -1 (2,5) #63
wire n1939; //OPIN -1 (2,5) #64
wire n1940; //OPIN -1 (2,5) #65
wire n1941; //OPIN -1 (2,5) #66
wire n1942; //OPIN -1 (2,5) #67
wire n1943; //OPIN -1 (2,5) #68
wire n1944; //OPIN -1 (2,5) #69
wire n1945; //OPIN -1 (2,5) #70
wire n1946; //OPIN -1 (2,5) #71
wire n1947; //IPIN -1 (2,5) #72
wire n1973; //IPIN -1 (2,6) #0
wire n1974; //IPIN -1 (2,6) #1
wire n1975; //IPIN -1 (2,6) #2
wire n1976; //IPIN -1 (2,6) #3
wire n1977; //IPIN -1 (2,6) #4
wire n1978; //IPIN -1 (2,6) #5
wire n1979; //IPIN -1 (2,6) #6
wire n1980; //IPIN -1 (2,6) #7
wire n1981; //IPIN -1 (2,6) #8
wire n1982; //IPIN -1 (2,6) #9
wire n1983; //IPIN -1 (2,6) #10
wire n1984; //IPIN -1 (2,6) #11
wire n1985; //IPIN -1 (2,6) #12
wire n1986; //IPIN -1 (2,6) #13
wire n1987; //IPIN -1 (2,6) #14
wire n1988; //IPIN -1 (2,6) #15
wire n1989; //IPIN -1 (2,6) #16
wire n1990; //IPIN -1 (2,6) #17
wire n1991; //IPIN -1 (2,6) #18
wire n1992; //IPIN -1 (2,6) #19
wire n1993; //IPIN -1 (2,6) #20
wire n1994; //IPIN -1 (2,6) #21
wire n1995; //IPIN -1 (2,6) #22
wire n1996; //IPIN -1 (2,6) #23
wire n1997; //IPIN -1 (2,6) #24
wire n1998; //IPIN -1 (2,6) #25
wire n1999; //IPIN -1 (2,6) #26
wire n2000; //IPIN -1 (2,6) #27
wire n2001; //IPIN -1 (2,6) #28
wire n2002; //IPIN -1 (2,6) #29
wire n2003; //IPIN -1 (2,6) #30
wire n2004; //IPIN -1 (2,6) #31
wire n2005; //IPIN -1 (2,6) #32
wire n2006; //IPIN -1 (2,6) #33
wire n2007; //IPIN -1 (2,6) #34
wire n2008; //IPIN -1 (2,6) #35
wire n2009; //IPIN -1 (2,6) #36
wire n2010; //IPIN -1 (2,6) #37
wire n2011; //IPIN -1 (2,6) #38
wire n2012; //IPIN -1 (2,6) #39
wire n2013; //IPIN -1 (2,6) #40
wire n2014; //IPIN -1 (2,6) #41
wire n2015; //IPIN -1 (2,6) #42
wire n2016; //IPIN -1 (2,6) #43
wire n2017; //IPIN -1 (2,6) #44
wire n2018; //IPIN -1 (2,6) #45
wire n2019; //IPIN -1 (2,6) #46
wire n2020; //IPIN -1 (2,6) #47
wire n2021; //IPIN -1 (2,6) #48
wire n2022; //IPIN -1 (2,6) #49
wire n2023; //IPIN -1 (2,6) #50
wire n2024; //IPIN -1 (2,6) #51
wire n2025; //OPIN -1 (2,6) #52
wire n2026; //OPIN -1 (2,6) #53
wire n2027; //OPIN -1 (2,6) #54
wire n2028; //OPIN -1 (2,6) #55
wire n2029; //OPIN -1 (2,6) #56
wire n2030; //OPIN -1 (2,6) #57
wire n2031; //OPIN -1 (2,6) #58
wire n2032; //OPIN -1 (2,6) #59
wire n2033; //OPIN -1 (2,6) #60
wire n2034; //OPIN -1 (2,6) #61
wire n2035; //OPIN -1 (2,6) #62
wire n2036; //OPIN -1 (2,6) #63
wire n2037; //OPIN -1 (2,6) #64
wire n2038; //OPIN -1 (2,6) #65
wire n2039; //OPIN -1 (2,6) #66
wire n2040; //OPIN -1 (2,6) #67
wire n2041; //OPIN -1 (2,6) #68
wire n2042; //OPIN -1 (2,6) #69
wire n2043; //OPIN -1 (2,6) #70
wire n2044; //OPIN -1 (2,6) #71
wire n2045; //IPIN -1 (2,6) #72
wire n2071; //IPIN -1 (2,7) #0
wire n2072; //IPIN -1 (2,7) #1
wire n2073; //IPIN -1 (2,7) #2
wire n2074; //IPIN -1 (2,7) #3
wire n2075; //IPIN -1 (2,7) #4
wire n2076; //IPIN -1 (2,7) #5
wire n2077; //IPIN -1 (2,7) #6
wire n2078; //IPIN -1 (2,7) #7
wire n2079; //IPIN -1 (2,7) #8
wire n2080; //IPIN -1 (2,7) #9
wire n2081; //IPIN -1 (2,7) #10
wire n2082; //IPIN -1 (2,7) #11
wire n2083; //IPIN -1 (2,7) #12
wire n2084; //IPIN -1 (2,7) #13
wire n2085; //IPIN -1 (2,7) #14
wire n2086; //IPIN -1 (2,7) #15
wire n2087; //IPIN -1 (2,7) #16
wire n2088; //IPIN -1 (2,7) #17
wire n2089; //IPIN -1 (2,7) #18
wire n2090; //IPIN -1 (2,7) #19
wire n2091; //IPIN -1 (2,7) #20
wire n2092; //IPIN -1 (2,7) #21
wire n2093; //IPIN -1 (2,7) #22
wire n2094; //IPIN -1 (2,7) #23
wire n2095; //IPIN -1 (2,7) #24
wire n2096; //IPIN -1 (2,7) #25
wire n2097; //IPIN -1 (2,7) #26
wire n2098; //IPIN -1 (2,7) #27
wire n2099; //IPIN -1 (2,7) #28
wire n2100; //IPIN -1 (2,7) #29
wire n2101; //IPIN -1 (2,7) #30
wire n2102; //IPIN -1 (2,7) #31
wire n2103; //IPIN -1 (2,7) #32
wire n2104; //IPIN -1 (2,7) #33
wire n2105; //IPIN -1 (2,7) #34
wire n2106; //IPIN -1 (2,7) #35
wire n2107; //IPIN -1 (2,7) #36
wire n2108; //IPIN -1 (2,7) #37
wire n2109; //IPIN -1 (2,7) #38
wire n2110; //IPIN -1 (2,7) #39
wire n2111; //IPIN -1 (2,7) #40
wire n2112; //IPIN -1 (2,7) #41
wire n2113; //IPIN -1 (2,7) #42
wire n2114; //IPIN -1 (2,7) #43
wire n2115; //IPIN -1 (2,7) #44
wire n2116; //IPIN -1 (2,7) #45
wire n2117; //IPIN -1 (2,7) #46
wire n2118; //IPIN -1 (2,7) #47
wire n2119; //IPIN -1 (2,7) #48
wire n2120; //IPIN -1 (2,7) #49
wire n2121; //IPIN -1 (2,7) #50
wire n2122; //IPIN -1 (2,7) #51
wire n2123; //OPIN -1 (2,7) #52
wire n2124; //OPIN -1 (2,7) #53
wire n2125; //OPIN -1 (2,7) #54
wire n2126; //OPIN -1 (2,7) #55
wire n2127; //OPIN -1 (2,7) #56
wire n2128; //OPIN -1 (2,7) #57
wire n2129; //OPIN -1 (2,7) #58
wire n2130; //OPIN -1 (2,7) #59
wire n2131; //OPIN -1 (2,7) #60
wire n2132; //OPIN -1 (2,7) #61
wire n2133; //OPIN -1 (2,7) #62
wire n2134; //OPIN -1 (2,7) #63
wire n2135; //OPIN -1 (2,7) #64
wire n2136; //OPIN -1 (2,7) #65
wire n2137; //OPIN -1 (2,7) #66
wire n2138; //OPIN -1 (2,7) #67
wire n2139; //OPIN -1 (2,7) #68
wire n2140; //OPIN -1 (2,7) #69
wire n2141; //OPIN -1 (2,7) #70
wire n2142; //OPIN -1 (2,7) #71
wire n2143; //IPIN -1 (2,7) #72
wire n2169; //IPIN -1 (2,8) #0
wire n2170; //IPIN -1 (2,8) #1
wire n2171; //IPIN -1 (2,8) #2
wire n2172; //IPIN -1 (2,8) #3
wire n2173; //IPIN -1 (2,8) #4
wire n2174; //IPIN -1 (2,8) #5
wire n2175; //IPIN -1 (2,8) #6
wire n2176; //IPIN -1 (2,8) #7
wire n2177; //IPIN -1 (2,8) #8
wire n2178; //IPIN -1 (2,8) #9
wire n2179; //IPIN -1 (2,8) #10
wire n2180; //IPIN -1 (2,8) #11
wire n2181; //IPIN -1 (2,8) #12
wire n2182; //IPIN -1 (2,8) #13
wire n2183; //IPIN -1 (2,8) #14
wire n2184; //IPIN -1 (2,8) #15
wire n2185; //IPIN -1 (2,8) #16
wire n2186; //IPIN -1 (2,8) #17
wire n2187; //IPIN -1 (2,8) #18
wire n2188; //IPIN -1 (2,8) #19
wire n2189; //IPIN -1 (2,8) #20
wire n2190; //IPIN -1 (2,8) #21
wire n2191; //IPIN -1 (2,8) #22
wire n2192; //IPIN -1 (2,8) #23
wire n2193; //IPIN -1 (2,8) #24
wire n2194; //IPIN -1 (2,8) #25
wire n2195; //IPIN -1 (2,8) #26
wire n2196; //IPIN -1 (2,8) #27
wire n2197; //IPIN -1 (2,8) #28
wire n2198; //IPIN -1 (2,8) #29
wire n2199; //IPIN -1 (2,8) #30
wire n2200; //IPIN -1 (2,8) #31
wire n2201; //IPIN -1 (2,8) #32
wire n2202; //IPIN -1 (2,8) #33
wire n2203; //IPIN -1 (2,8) #34
wire n2204; //IPIN -1 (2,8) #35
wire n2205; //IPIN -1 (2,8) #36
wire n2206; //IPIN -1 (2,8) #37
wire n2207; //IPIN -1 (2,8) #38
wire n2208; //IPIN -1 (2,8) #39
wire n2209; //IPIN -1 (2,8) #40
wire n2210; //IPIN -1 (2,8) #41
wire n2211; //IPIN -1 (2,8) #42
wire n2212; //IPIN -1 (2,8) #43
wire n2213; //IPIN -1 (2,8) #44
wire n2214; //IPIN -1 (2,8) #45
wire n2215; //IPIN -1 (2,8) #46
wire n2216; //IPIN -1 (2,8) #47
wire n2217; //IPIN -1 (2,8) #48
wire n2218; //IPIN -1 (2,8) #49
wire n2219; //IPIN -1 (2,8) #50
wire n2220; //IPIN -1 (2,8) #51
wire n2221; //OPIN -1 (2,8) #52
wire n2222; //OPIN -1 (2,8) #53
wire n2223; //OPIN -1 (2,8) #54
wire n2224; //OPIN -1 (2,8) #55
wire n2225; //OPIN -1 (2,8) #56
wire n2226; //OPIN -1 (2,8) #57
wire n2227; //OPIN -1 (2,8) #58
wire n2228; //OPIN -1 (2,8) #59
wire n2229; //OPIN -1 (2,8) #60
wire n2230; //OPIN -1 (2,8) #61
wire n2231; //OPIN -1 (2,8) #62
wire n2232; //OPIN -1 (2,8) #63
wire n2233; //OPIN -1 (2,8) #64
wire n2234; //OPIN -1 (2,8) #65
wire n2235; //OPIN -1 (2,8) #66
wire n2236; //OPIN -1 (2,8) #67
wire n2237; //OPIN -1 (2,8) #68
wire n2238; //OPIN -1 (2,8) #69
wire n2239; //OPIN -1 (2,8) #70
wire n2240; //OPIN -1 (2,8) #71
wire n2241; //IPIN -1 (2,8) #72
wire n2267; //IPIN -1 (2,9) #0
wire n2268; //IPIN -1 (2,9) #1
wire n2269; //IPIN -1 (2,9) #2
wire n2270; //IPIN -1 (2,9) #3
wire n2271; //IPIN -1 (2,9) #4
wire n2272; //IPIN -1 (2,9) #5
wire n2273; //IPIN -1 (2,9) #6
wire n2274; //IPIN -1 (2,9) #7
wire n2275; //IPIN -1 (2,9) #8
wire n2276; //IPIN -1 (2,9) #9
wire n2277; //IPIN -1 (2,9) #10
wire n2278; //IPIN -1 (2,9) #11
wire n2279; //IPIN -1 (2,9) #12
wire n2280; //IPIN -1 (2,9) #13
wire n2281; //IPIN -1 (2,9) #14
wire n2282; //IPIN -1 (2,9) #15
wire n2283; //IPIN -1 (2,9) #16
wire n2284; //IPIN -1 (2,9) #17
wire n2285; //IPIN -1 (2,9) #18
wire n2286; //IPIN -1 (2,9) #19
wire n2287; //IPIN -1 (2,9) #20
wire n2288; //IPIN -1 (2,9) #21
wire n2289; //IPIN -1 (2,9) #22
wire n2290; //IPIN -1 (2,9) #23
wire n2291; //IPIN -1 (2,9) #24
wire n2292; //IPIN -1 (2,9) #25
wire n2293; //IPIN -1 (2,9) #26
wire n2294; //IPIN -1 (2,9) #27
wire n2295; //IPIN -1 (2,9) #28
wire n2296; //IPIN -1 (2,9) #29
wire n2297; //IPIN -1 (2,9) #30
wire n2298; //IPIN -1 (2,9) #31
wire n2299; //IPIN -1 (2,9) #32
wire n2300; //IPIN -1 (2,9) #33
wire n2301; //IPIN -1 (2,9) #34
wire n2302; //IPIN -1 (2,9) #35
wire n2303; //IPIN -1 (2,9) #36
wire n2304; //IPIN -1 (2,9) #37
wire n2305; //IPIN -1 (2,9) #38
wire n2306; //IPIN -1 (2,9) #39
wire n2307; //IPIN -1 (2,9) #40
wire n2308; //IPIN -1 (2,9) #41
wire n2309; //IPIN -1 (2,9) #42
wire n2310; //IPIN -1 (2,9) #43
wire n2311; //IPIN -1 (2,9) #44
wire n2312; //IPIN -1 (2,9) #45
wire n2313; //IPIN -1 (2,9) #46
wire n2314; //IPIN -1 (2,9) #47
wire n2315; //IPIN -1 (2,9) #48
wire n2316; //IPIN -1 (2,9) #49
wire n2317; //IPIN -1 (2,9) #50
wire n2318; //IPIN -1 (2,9) #51
wire n2319; //OPIN -1 (2,9) #52
wire n2320; //OPIN -1 (2,9) #53
wire n2321; //OPIN -1 (2,9) #54
wire n2322; //OPIN -1 (2,9) #55
wire n2323; //OPIN -1 (2,9) #56
wire n2324; //OPIN -1 (2,9) #57
wire n2325; //OPIN -1 (2,9) #58
wire n2326; //OPIN -1 (2,9) #59
wire n2327; //OPIN -1 (2,9) #60
wire n2328; //OPIN -1 (2,9) #61
wire n2329; //OPIN -1 (2,9) #62
wire n2330; //OPIN -1 (2,9) #63
wire n2331; //OPIN -1 (2,9) #64
wire n2332; //OPIN -1 (2,9) #65
wire n2333; //OPIN -1 (2,9) #66
wire n2334; //OPIN -1 (2,9) #67
wire n2335; //OPIN -1 (2,9) #68
wire n2336; //OPIN -1 (2,9) #69
wire n2337; //OPIN -1 (2,9) #70
wire n2338; //OPIN -1 (2,9) #71
wire n2339; //IPIN -1 (2,9) #72
wire n2364; //IPIN -1 (2,10) #0
wire n2365; //OPIN -1 (2,10) #1
wire n2366; //IPIN -1 (2,10) #2
wire n2367; //IPIN -1 (2,10) #3
wire n2368; //OPIN -1 (2,10) #4
wire n2369; //IPIN -1 (2,10) #5
wire n2370; //IPIN -1 (2,10) #6
wire n2371; //OPIN -1 (2,10) #7
wire n2372; //IPIN -1 (2,10) #8
wire n2373; //IPIN -1 (2,10) #9
wire n2374; //OPIN -1 (2,10) #10
wire n2375; //IPIN -1 (2,10) #11
wire n2376; //IPIN -1 (2,10) #12
wire n2377; //OPIN -1 (2,10) #13
wire n2378; //IPIN -1 (2,10) #14
wire n2379; //IPIN -1 (2,10) #15
wire n2380; //OPIN -1 (2,10) #16
wire n2381; //IPIN -1 (2,10) #17
wire n2382; //IPIN -1 (2,10) #18
wire n2383; //OPIN -1 (2,10) #19
wire n2384; //IPIN -1 (2,10) #20
wire n2385; //IPIN -1 (2,10) #21
wire n2386; //OPIN -1 (2,10) #22
wire n2387; //IPIN -1 (2,10) #23
wire n2412; //IPIN -1 (3,0) #0
wire n2413; //OPIN -1 (3,0) #1
wire n2414; //IPIN -1 (3,0) #2
wire n2415; //IPIN -1 (3,0) #3
wire n2416; //OPIN -1 (3,0) #4
wire n2417; //IPIN -1 (3,0) #5
wire n2418; //IPIN -1 (3,0) #6
wire n2419; //OPIN -1 (3,0) #7
wire n2420; //IPIN -1 (3,0) #8
wire n2421; //IPIN -1 (3,0) #9
wire n2422; //OPIN -1 (3,0) #10
wire n2423; //IPIN -1 (3,0) #11
wire n2424; //IPIN -1 (3,0) #12
wire n2425; //OPIN -1 (3,0) #13
wire n2426; //IPIN -1 (3,0) #14
wire n2427; //IPIN -1 (3,0) #15
wire n2428; //OPIN -1 (3,0) #16
wire n2429; //IPIN -1 (3,0) #17
wire n2430; //IPIN -1 (3,0) #18
wire n2431; //OPIN -1 (3,0) #19
wire n2432; //IPIN -1 (3,0) #20
wire n2433; //IPIN -1 (3,0) #21
wire n2434; //OPIN -1 (3,0) #22
wire n2435; //IPIN -1 (3,0) #23
wire n2461; //IPIN -1 (3,1) #0
wire n2462; //IPIN -1 (3,1) #1
wire n2463; //IPIN -1 (3,1) #2
wire n2464; //IPIN -1 (3,1) #3
wire n2465; //IPIN -1 (3,1) #4
wire n2466; //IPIN -1 (3,1) #5
wire n2467; //IPIN -1 (3,1) #6
wire n2468; //IPIN -1 (3,1) #7
wire n2469; //IPIN -1 (3,1) #8
wire n2470; //IPIN -1 (3,1) #9
wire n2471; //IPIN -1 (3,1) #10
wire n2472; //IPIN -1 (3,1) #11
wire n2473; //IPIN -1 (3,1) #12
wire n2474; //IPIN -1 (3,1) #13
wire n2475; //IPIN -1 (3,1) #14
wire n2476; //IPIN -1 (3,1) #15
wire n2477; //IPIN -1 (3,1) #16
wire n2478; //IPIN -1 (3,1) #17
wire n2479; //IPIN -1 (3,1) #18
wire n2480; //IPIN -1 (3,1) #19
wire n2481; //IPIN -1 (3,1) #20
wire n2482; //IPIN -1 (3,1) #21
wire n2483; //IPIN -1 (3,1) #22
wire n2484; //IPIN -1 (3,1) #23
wire n2485; //IPIN -1 (3,1) #24
wire n2486; //IPIN -1 (3,1) #25
wire n2487; //IPIN -1 (3,1) #26
wire n2488; //IPIN -1 (3,1) #27
wire n2489; //IPIN -1 (3,1) #28
wire n2490; //IPIN -1 (3,1) #29
wire n2491; //IPIN -1 (3,1) #30
wire n2492; //IPIN -1 (3,1) #31
wire n2493; //IPIN -1 (3,1) #32
wire n2494; //IPIN -1 (3,1) #33
wire n2495; //IPIN -1 (3,1) #34
wire n2496; //IPIN -1 (3,1) #35
wire n2497; //IPIN -1 (3,1) #36
wire n2498; //IPIN -1 (3,1) #37
wire n2499; //IPIN -1 (3,1) #38
wire n2500; //IPIN -1 (3,1) #39
wire n2501; //IPIN -1 (3,1) #40
wire n2502; //IPIN -1 (3,1) #41
wire n2503; //IPIN -1 (3,1) #42
wire n2504; //IPIN -1 (3,1) #43
wire n2505; //IPIN -1 (3,1) #44
wire n2506; //IPIN -1 (3,1) #45
wire n2507; //IPIN -1 (3,1) #46
wire n2508; //IPIN -1 (3,1) #47
wire n2509; //IPIN -1 (3,1) #48
wire n2510; //IPIN -1 (3,1) #49
wire n2511; //IPIN -1 (3,1) #50
wire n2512; //IPIN -1 (3,1) #51
wire n2513; //OPIN -1 (3,1) #52
wire n2514; //OPIN -1 (3,1) #53
wire n2515; //OPIN -1 (3,1) #54
wire n2516; //OPIN -1 (3,1) #55
wire n2517; //OPIN -1 (3,1) #56
wire n2518; //OPIN -1 (3,1) #57
wire n2519; //OPIN -1 (3,1) #58
wire n2520; //OPIN -1 (3,1) #59
wire n2521; //OPIN -1 (3,1) #60
wire n2522; //OPIN -1 (3,1) #61
wire n2523; //OPIN -1 (3,1) #62
wire n2524; //OPIN -1 (3,1) #63
wire n2525; //OPIN -1 (3,1) #64
wire n2526; //OPIN -1 (3,1) #65
wire n2527; //OPIN -1 (3,1) #66
wire n2528; //OPIN -1 (3,1) #67
wire n2529; //OPIN -1 (3,1) #68
wire n2530; //OPIN -1 (3,1) #69
wire n2531; //OPIN -1 (3,1) #70
wire n2532; //OPIN -1 (3,1) #71
wire n2533; //IPIN -1 (3,1) #72
wire n2559; //IPIN -1 (3,2) #0
wire n2560; //IPIN -1 (3,2) #1
wire n2561; //IPIN -1 (3,2) #2
wire n2562; //IPIN -1 (3,2) #3
wire n2563; //IPIN -1 (3,2) #4
wire n2564; //IPIN -1 (3,2) #5
wire n2565; //IPIN -1 (3,2) #6
wire n2566; //IPIN -1 (3,2) #7
wire n2567; //IPIN -1 (3,2) #8
wire n2568; //IPIN -1 (3,2) #9
wire n2569; //IPIN -1 (3,2) #10
wire n2570; //IPIN -1 (3,2) #11
wire n2571; //IPIN -1 (3,2) #12
wire n2572; //IPIN -1 (3,2) #13
wire n2573; //IPIN -1 (3,2) #14
wire n2574; //IPIN -1 (3,2) #15
wire n2575; //IPIN -1 (3,2) #16
wire n2576; //IPIN -1 (3,2) #17
wire n2577; //IPIN -1 (3,2) #18
wire n2578; //IPIN -1 (3,2) #19
wire n2579; //IPIN -1 (3,2) #20
wire n2580; //IPIN -1 (3,2) #21
wire n2581; //IPIN -1 (3,2) #22
wire n2582; //IPIN -1 (3,2) #23
wire n2583; //IPIN -1 (3,2) #24
wire n2584; //IPIN -1 (3,2) #25
wire n2585; //IPIN -1 (3,2) #26
wire n2586; //IPIN -1 (3,2) #27
wire n2587; //IPIN -1 (3,2) #28
wire n2588; //IPIN -1 (3,2) #29
wire n2589; //IPIN -1 (3,2) #30
wire n2590; //IPIN -1 (3,2) #31
wire n2591; //IPIN -1 (3,2) #32
wire n2592; //IPIN -1 (3,2) #33
wire n2593; //IPIN -1 (3,2) #34
wire n2594; //IPIN -1 (3,2) #35
wire n2595; //IPIN -1 (3,2) #36
wire n2596; //IPIN -1 (3,2) #37
wire n2597; //IPIN -1 (3,2) #38
wire n2598; //IPIN -1 (3,2) #39
wire n2599; //IPIN -1 (3,2) #40
wire n2600; //IPIN -1 (3,2) #41
wire n2601; //IPIN -1 (3,2) #42
wire n2602; //IPIN -1 (3,2) #43
wire n2603; //IPIN -1 (3,2) #44
wire n2604; //IPIN -1 (3,2) #45
wire n2605; //IPIN -1 (3,2) #46
wire n2606; //IPIN -1 (3,2) #47
wire n2607; //IPIN -1 (3,2) #48
wire n2608; //IPIN -1 (3,2) #49
wire n2609; //IPIN -1 (3,2) #50
wire n2610; //IPIN -1 (3,2) #51
wire n2611; //OPIN -1 (3,2) #52
wire n2612; //OPIN -1 (3,2) #53
wire n2613; //OPIN -1 (3,2) #54
wire n2614; //OPIN -1 (3,2) #55
wire n2615; //OPIN -1 (3,2) #56
wire n2616; //OPIN -1 (3,2) #57
wire n2617; //OPIN -1 (3,2) #58
wire n2618; //OPIN -1 (3,2) #59
wire n2619; //OPIN -1 (3,2) #60
wire n2620; //OPIN -1 (3,2) #61
wire n2621; //OPIN -1 (3,2) #62
wire n2622; //OPIN -1 (3,2) #63
wire n2623; //OPIN -1 (3,2) #64
wire n2624; //OPIN -1 (3,2) #65
wire n2625; //OPIN -1 (3,2) #66
wire n2626; //OPIN -1 (3,2) #67
wire n2627; //OPIN -1 (3,2) #68
wire n2628; //OPIN -1 (3,2) #69
wire n2629; //OPIN -1 (3,2) #70
wire n2630; //OPIN -1 (3,2) #71
wire n2631; //IPIN -1 (3,2) #72
wire n2657; //IPIN -1 (3,3) #0
wire n2658; //IPIN -1 (3,3) #1
wire n2659; //IPIN -1 (3,3) #2
wire n2660; //IPIN -1 (3,3) #3
wire n2661; //IPIN -1 (3,3) #4
wire n2662; //IPIN -1 (3,3) #5
wire n2663; //IPIN -1 (3,3) #6
wire n2664; //IPIN -1 (3,3) #7
wire n2665; //IPIN -1 (3,3) #8
wire n2666; //IPIN -1 (3,3) #9
wire n2667; //IPIN -1 (3,3) #10
wire n2668; //IPIN -1 (3,3) #11
wire n2669; //IPIN -1 (3,3) #12
wire n2670; //IPIN -1 (3,3) #13
wire n2671; //IPIN -1 (3,3) #14
wire n2672; //IPIN -1 (3,3) #15
wire n2673; //IPIN -1 (3,3) #16
wire n2674; //IPIN -1 (3,3) #17
wire n2675; //IPIN -1 (3,3) #18
wire n2676; //IPIN -1 (3,3) #19
wire n2677; //IPIN -1 (3,3) #20
wire n2678; //IPIN -1 (3,3) #21
wire n2679; //IPIN -1 (3,3) #22
wire n2680; //IPIN -1 (3,3) #23
wire n2681; //IPIN -1 (3,3) #24
wire n2682; //IPIN -1 (3,3) #25
wire n2683; //IPIN -1 (3,3) #26
wire n2684; //IPIN -1 (3,3) #27
wire n2685; //IPIN -1 (3,3) #28
wire n2686; //IPIN -1 (3,3) #29
wire n2687; //IPIN -1 (3,3) #30
wire n2688; //IPIN -1 (3,3) #31
wire n2689; //IPIN -1 (3,3) #32
wire n2690; //IPIN -1 (3,3) #33
wire n2691; //IPIN -1 (3,3) #34
wire n2692; //IPIN -1 (3,3) #35
wire n2693; //IPIN -1 (3,3) #36
wire n2694; //IPIN -1 (3,3) #37
wire n2695; //IPIN -1 (3,3) #38
wire n2696; //IPIN -1 (3,3) #39
wire n2697; //IPIN -1 (3,3) #40
wire n2698; //IPIN -1 (3,3) #41
wire n2699; //IPIN -1 (3,3) #42
wire n2700; //IPIN -1 (3,3) #43
wire n2701; //IPIN -1 (3,3) #44
wire n2702; //IPIN -1 (3,3) #45
wire n2703; //IPIN -1 (3,3) #46
wire n2704; //IPIN -1 (3,3) #47
wire n2705; //IPIN -1 (3,3) #48
wire n2706; //IPIN -1 (3,3) #49
wire n2707; //IPIN -1 (3,3) #50
wire n2708; //IPIN -1 (3,3) #51
wire n2709; //OPIN -1 (3,3) #52
wire n2710; //OPIN -1 (3,3) #53
wire n2711; //OPIN -1 (3,3) #54
wire n2712; //OPIN -1 (3,3) #55
wire n2713; //OPIN -1 (3,3) #56
wire n2714; //OPIN -1 (3,3) #57
wire n2715; //OPIN -1 (3,3) #58
wire n2716; //OPIN -1 (3,3) #59
wire n2717; //OPIN -1 (3,3) #60
wire n2718; //OPIN -1 (3,3) #61
wire n2719; //OPIN -1 (3,3) #62
wire n2720; //OPIN -1 (3,3) #63
wire n2721; //OPIN -1 (3,3) #64
wire n2722; //OPIN -1 (3,3) #65
wire n2723; //OPIN -1 (3,3) #66
wire n2724; //OPIN -1 (3,3) #67
wire n2725; //OPIN -1 (3,3) #68
wire n2726; //OPIN -1 (3,3) #69
wire n2727; //OPIN -1 (3,3) #70
wire n2728; //OPIN -1 (3,3) #71
wire n2729; //IPIN -1 (3,3) #72
wire n2755; //IPIN -1 (3,4) #0
wire n2756; //IPIN -1 (3,4) #1
wire n2757; //IPIN -1 (3,4) #2
wire n2758; //IPIN -1 (3,4) #3
wire n2759; //IPIN -1 (3,4) #4
wire n2760; //IPIN -1 (3,4) #5
wire n2761; //IPIN -1 (3,4) #6
wire n2762; //IPIN -1 (3,4) #7
wire n2763; //IPIN -1 (3,4) #8
wire n2764; //IPIN -1 (3,4) #9
wire n2765; //IPIN -1 (3,4) #10
wire n2766; //IPIN -1 (3,4) #11
wire n2767; //IPIN -1 (3,4) #12
wire n2768; //IPIN -1 (3,4) #13
wire n2769; //IPIN -1 (3,4) #14
wire n2770; //IPIN -1 (3,4) #15
wire n2771; //IPIN -1 (3,4) #16
wire n2772; //IPIN -1 (3,4) #17
wire n2773; //IPIN -1 (3,4) #18
wire n2774; //IPIN -1 (3,4) #19
wire n2775; //IPIN -1 (3,4) #20
wire n2776; //IPIN -1 (3,4) #21
wire n2777; //IPIN -1 (3,4) #22
wire n2778; //IPIN -1 (3,4) #23
wire n2779; //IPIN -1 (3,4) #24
wire n2780; //IPIN -1 (3,4) #25
wire n2781; //IPIN -1 (3,4) #26
wire n2782; //IPIN -1 (3,4) #27
wire n2783; //IPIN -1 (3,4) #28
wire n2784; //IPIN -1 (3,4) #29
wire n2785; //IPIN -1 (3,4) #30
wire n2786; //IPIN -1 (3,4) #31
wire n2787; //IPIN -1 (3,4) #32
wire n2788; //IPIN -1 (3,4) #33
wire n2789; //IPIN -1 (3,4) #34
wire n2790; //IPIN -1 (3,4) #35
wire n2791; //IPIN -1 (3,4) #36
wire n2792; //IPIN -1 (3,4) #37
wire n2793; //IPIN -1 (3,4) #38
wire n2794; //IPIN -1 (3,4) #39
wire n2795; //IPIN -1 (3,4) #40
wire n2796; //IPIN -1 (3,4) #41
wire n2797; //IPIN -1 (3,4) #42
wire n2798; //IPIN -1 (3,4) #43
wire n2799; //IPIN -1 (3,4) #44
wire n2800; //IPIN -1 (3,4) #45
wire n2801; //IPIN -1 (3,4) #46
wire n2802; //IPIN -1 (3,4) #47
wire n2803; //IPIN -1 (3,4) #48
wire n2804; //IPIN -1 (3,4) #49
wire n2805; //IPIN -1 (3,4) #50
wire n2806; //IPIN -1 (3,4) #51
wire n2807; //OPIN -1 (3,4) #52
wire n2808; //OPIN -1 (3,4) #53
wire n2809; //OPIN -1 (3,4) #54
wire n2810; //OPIN -1 (3,4) #55
wire n2811; //OPIN -1 (3,4) #56
wire n2812; //OPIN -1 (3,4) #57
wire n2813; //OPIN -1 (3,4) #58
wire n2814; //OPIN -1 (3,4) #59
wire n2815; //OPIN -1 (3,4) #60
wire n2816; //OPIN -1 (3,4) #61
wire n2817; //OPIN -1 (3,4) #62
wire n2818; //OPIN -1 (3,4) #63
wire n2819; //OPIN -1 (3,4) #64
wire n2820; //OPIN -1 (3,4) #65
wire n2821; //OPIN -1 (3,4) #66
wire n2822; //OPIN -1 (3,4) #67
wire n2823; //OPIN -1 (3,4) #68
wire n2824; //OPIN -1 (3,4) #69
wire n2825; //OPIN -1 (3,4) #70
wire n2826; //OPIN -1 (3,4) #71
wire n2827; //IPIN -1 (3,4) #72
wire n2853; //IPIN -1 (3,5) #0
wire n2854; //IPIN -1 (3,5) #1
wire n2855; //IPIN -1 (3,5) #2
wire n2856; //IPIN -1 (3,5) #3
wire n2857; //IPIN -1 (3,5) #4
wire n2858; //IPIN -1 (3,5) #5
wire n2859; //IPIN -1 (3,5) #6
wire n2860; //IPIN -1 (3,5) #7
wire n2861; //IPIN -1 (3,5) #8
wire n2862; //IPIN -1 (3,5) #9
wire n2863; //IPIN -1 (3,5) #10
wire n2864; //IPIN -1 (3,5) #11
wire n2865; //IPIN -1 (3,5) #12
wire n2866; //IPIN -1 (3,5) #13
wire n2867; //IPIN -1 (3,5) #14
wire n2868; //IPIN -1 (3,5) #15
wire n2869; //IPIN -1 (3,5) #16
wire n2870; //IPIN -1 (3,5) #17
wire n2871; //IPIN -1 (3,5) #18
wire n2872; //IPIN -1 (3,5) #19
wire n2873; //IPIN -1 (3,5) #20
wire n2874; //IPIN -1 (3,5) #21
wire n2875; //IPIN -1 (3,5) #22
wire n2876; //IPIN -1 (3,5) #23
wire n2877; //IPIN -1 (3,5) #24
wire n2878; //IPIN -1 (3,5) #25
wire n2879; //IPIN -1 (3,5) #26
wire n2880; //IPIN -1 (3,5) #27
wire n2881; //IPIN -1 (3,5) #28
wire n2882; //IPIN -1 (3,5) #29
wire n2883; //IPIN -1 (3,5) #30
wire n2884; //IPIN -1 (3,5) #31
wire n2885; //IPIN -1 (3,5) #32
wire n2886; //IPIN -1 (3,5) #33
wire n2887; //IPIN -1 (3,5) #34
wire n2888; //IPIN -1 (3,5) #35
wire n2889; //IPIN -1 (3,5) #36
wire n2890; //IPIN -1 (3,5) #37
wire n2891; //IPIN -1 (3,5) #38
wire n2892; //IPIN -1 (3,5) #39
wire n2893; //IPIN -1 (3,5) #40
wire n2894; //IPIN -1 (3,5) #41
wire n2895; //IPIN -1 (3,5) #42
wire n2896; //IPIN -1 (3,5) #43
wire n2897; //IPIN -1 (3,5) #44
wire n2898; //IPIN -1 (3,5) #45
wire n2899; //IPIN -1 (3,5) #46
wire n2900; //IPIN -1 (3,5) #47
wire n2901; //IPIN -1 (3,5) #48
wire n2902; //IPIN -1 (3,5) #49
wire n2903; //IPIN -1 (3,5) #50
wire n2904; //IPIN -1 (3,5) #51
wire n2905; //OPIN -1 (3,5) #52
wire n2906; //OPIN -1 (3,5) #53
wire n2907; //OPIN -1 (3,5) #54
wire n2908; //OPIN -1 (3,5) #55
wire n2909; //OPIN -1 (3,5) #56
wire n2910; //OPIN -1 (3,5) #57
wire n2911; //OPIN -1 (3,5) #58
wire n2912; //OPIN -1 (3,5) #59
wire n2913; //OPIN -1 (3,5) #60
wire n2914; //OPIN -1 (3,5) #61
wire n2915; //OPIN -1 (3,5) #62
wire n2916; //OPIN -1 (3,5) #63
wire n2917; //OPIN -1 (3,5) #64
wire n2918; //OPIN -1 (3,5) #65
wire n2919; //OPIN -1 (3,5) #66
wire n2920; //OPIN -1 (3,5) #67
wire n2921; //OPIN -1 (3,5) #68
wire n2922; //OPIN -1 (3,5) #69
wire n2923; //OPIN -1 (3,5) #70
wire n2924; //OPIN -1 (3,5) #71
wire n2925; //IPIN -1 (3,5) #72
wire n2951; //IPIN -1 (3,6) #0
wire n2952; //IPIN -1 (3,6) #1
wire n2953; //IPIN -1 (3,6) #2
wire n2954; //IPIN -1 (3,6) #3
wire n2955; //IPIN -1 (3,6) #4
wire n2956; //IPIN -1 (3,6) #5
wire n2957; //IPIN -1 (3,6) #6
wire n2958; //IPIN -1 (3,6) #7
wire n2959; //IPIN -1 (3,6) #8
wire n2960; //IPIN -1 (3,6) #9
wire n2961; //IPIN -1 (3,6) #10
wire n2962; //IPIN -1 (3,6) #11
wire n2963; //IPIN -1 (3,6) #12
wire n2964; //IPIN -1 (3,6) #13
wire n2965; //IPIN -1 (3,6) #14
wire n2966; //IPIN -1 (3,6) #15
wire n2967; //IPIN -1 (3,6) #16
wire n2968; //IPIN -1 (3,6) #17
wire n2969; //IPIN -1 (3,6) #18
wire n2970; //IPIN -1 (3,6) #19
wire n2971; //IPIN -1 (3,6) #20
wire n2972; //IPIN -1 (3,6) #21
wire n2973; //IPIN -1 (3,6) #22
wire n2974; //IPIN -1 (3,6) #23
wire n2975; //IPIN -1 (3,6) #24
wire n2976; //IPIN -1 (3,6) #25
wire n2977; //IPIN -1 (3,6) #26
wire n2978; //IPIN -1 (3,6) #27
wire n2979; //IPIN -1 (3,6) #28
wire n2980; //IPIN -1 (3,6) #29
wire n2981; //IPIN -1 (3,6) #30
wire n2982; //IPIN -1 (3,6) #31
wire n2983; //IPIN -1 (3,6) #32
wire n2984; //IPIN -1 (3,6) #33
wire n2985; //IPIN -1 (3,6) #34
wire n2986; //IPIN -1 (3,6) #35
wire n2987; //IPIN -1 (3,6) #36
wire n2988; //IPIN -1 (3,6) #37
wire n2989; //IPIN -1 (3,6) #38
wire n2990; //IPIN -1 (3,6) #39
wire n2991; //IPIN -1 (3,6) #40
wire n2992; //IPIN -1 (3,6) #41
wire n2993; //IPIN -1 (3,6) #42
wire n2994; //IPIN -1 (3,6) #43
wire n2995; //IPIN -1 (3,6) #44
wire n2996; //IPIN -1 (3,6) #45
wire n2997; //IPIN -1 (3,6) #46
wire n2998; //IPIN -1 (3,6) #47
wire n2999; //IPIN -1 (3,6) #48
wire n3000; //IPIN -1 (3,6) #49
wire n3001; //IPIN -1 (3,6) #50
wire n3002; //IPIN -1 (3,6) #51
wire n3003; //OPIN -1 (3,6) #52
wire n3004; //OPIN -1 (3,6) #53
wire n3005; //OPIN -1 (3,6) #54
wire n3006; //OPIN -1 (3,6) #55
wire n3007; //OPIN -1 (3,6) #56
wire n3008; //OPIN -1 (3,6) #57
wire n3009; //OPIN -1 (3,6) #58
wire n3010; //OPIN -1 (3,6) #59
wire n3011; //OPIN -1 (3,6) #60
wire n3012; //OPIN -1 (3,6) #61
wire n3013; //OPIN -1 (3,6) #62
wire n3014; //OPIN -1 (3,6) #63
wire n3015; //OPIN -1 (3,6) #64
wire n3016; //OPIN -1 (3,6) #65
wire n3017; //OPIN -1 (3,6) #66
wire n3018; //OPIN -1 (3,6) #67
wire n3019; //OPIN -1 (3,6) #68
wire n3020; //OPIN -1 (3,6) #69
wire n3021; //OPIN -1 (3,6) #70
wire n3022; //OPIN -1 (3,6) #71
wire n3023; //IPIN -1 (3,6) #72
wire n3049; //IPIN -1 (3,7) #0
wire n3050; //IPIN -1 (3,7) #1
wire n3051; //IPIN -1 (3,7) #2
wire n3052; //IPIN -1 (3,7) #3
wire n3053; //IPIN -1 (3,7) #4
wire n3054; //IPIN -1 (3,7) #5
wire n3055; //IPIN -1 (3,7) #6
wire n3056; //IPIN -1 (3,7) #7
wire n3057; //IPIN -1 (3,7) #8
wire n3058; //IPIN -1 (3,7) #9
wire n3059; //IPIN -1 (3,7) #10
wire n3060; //IPIN -1 (3,7) #11
wire n3061; //IPIN -1 (3,7) #12
wire n3062; //IPIN -1 (3,7) #13
wire n3063; //IPIN -1 (3,7) #14
wire n3064; //IPIN -1 (3,7) #15
wire n3065; //IPIN -1 (3,7) #16
wire n3066; //IPIN -1 (3,7) #17
wire n3067; //IPIN -1 (3,7) #18
wire n3068; //IPIN -1 (3,7) #19
wire n3069; //IPIN -1 (3,7) #20
wire n3070; //IPIN -1 (3,7) #21
wire n3071; //IPIN -1 (3,7) #22
wire n3072; //IPIN -1 (3,7) #23
wire n3073; //IPIN -1 (3,7) #24
wire n3074; //IPIN -1 (3,7) #25
wire n3075; //IPIN -1 (3,7) #26
wire n3076; //IPIN -1 (3,7) #27
wire n3077; //IPIN -1 (3,7) #28
wire n3078; //IPIN -1 (3,7) #29
wire n3079; //IPIN -1 (3,7) #30
wire n3080; //IPIN -1 (3,7) #31
wire n3081; //IPIN -1 (3,7) #32
wire n3082; //IPIN -1 (3,7) #33
wire n3083; //IPIN -1 (3,7) #34
wire n3084; //IPIN -1 (3,7) #35
wire n3085; //IPIN -1 (3,7) #36
wire n3086; //IPIN -1 (3,7) #37
wire n3087; //IPIN -1 (3,7) #38
wire n3088; //IPIN -1 (3,7) #39
wire n3089; //IPIN -1 (3,7) #40
wire n3090; //IPIN -1 (3,7) #41
wire n3091; //IPIN -1 (3,7) #42
wire n3092; //IPIN -1 (3,7) #43
wire n3093; //IPIN -1 (3,7) #44
wire n3094; //IPIN -1 (3,7) #45
wire n3095; //IPIN -1 (3,7) #46
wire n3096; //IPIN -1 (3,7) #47
wire n3097; //IPIN -1 (3,7) #48
wire n3098; //IPIN -1 (3,7) #49
wire n3099; //IPIN -1 (3,7) #50
wire n3100; //IPIN -1 (3,7) #51
wire n3101; //OPIN -1 (3,7) #52
wire n3102; //OPIN -1 (3,7) #53
wire n3103; //OPIN -1 (3,7) #54
wire n3104; //OPIN -1 (3,7) #55
wire n3105; //OPIN -1 (3,7) #56
wire n3106; //OPIN -1 (3,7) #57
wire n3107; //OPIN -1 (3,7) #58
wire n3108; //OPIN -1 (3,7) #59
wire n3109; //OPIN -1 (3,7) #60
wire n3110; //OPIN -1 (3,7) #61
wire n3111; //OPIN -1 (3,7) #62
wire n3112; //OPIN -1 (3,7) #63
wire n3113; //OPIN -1 (3,7) #64
wire n3114; //OPIN -1 (3,7) #65
wire n3115; //OPIN -1 (3,7) #66
wire n3116; //OPIN -1 (3,7) #67
wire n3117; //OPIN -1 (3,7) #68
wire n3118; //OPIN -1 (3,7) #69
wire n3119; //OPIN -1 (3,7) #70
wire n3120; //OPIN -1 (3,7) #71
wire n3121; //IPIN -1 (3,7) #72
wire n3147; //IPIN -1 (3,8) #0
wire n3148; //IPIN -1 (3,8) #1
wire n3149; //IPIN -1 (3,8) #2
wire n3150; //IPIN -1 (3,8) #3
wire n3151; //IPIN -1 (3,8) #4
wire n3152; //IPIN -1 (3,8) #5
wire n3153; //IPIN -1 (3,8) #6
wire n3154; //IPIN -1 (3,8) #7
wire n3155; //IPIN -1 (3,8) #8
wire n3156; //IPIN -1 (3,8) #9
wire n3157; //IPIN -1 (3,8) #10
wire n3158; //IPIN -1 (3,8) #11
wire n3159; //IPIN -1 (3,8) #12
wire n3160; //IPIN -1 (3,8) #13
wire n3161; //IPIN -1 (3,8) #14
wire n3162; //IPIN -1 (3,8) #15
wire n3163; //IPIN -1 (3,8) #16
wire n3164; //IPIN -1 (3,8) #17
wire n3165; //IPIN -1 (3,8) #18
wire n3166; //IPIN -1 (3,8) #19
wire n3167; //IPIN -1 (3,8) #20
wire n3168; //IPIN -1 (3,8) #21
wire n3169; //IPIN -1 (3,8) #22
wire n3170; //IPIN -1 (3,8) #23
wire n3171; //IPIN -1 (3,8) #24
wire n3172; //IPIN -1 (3,8) #25
wire n3173; //IPIN -1 (3,8) #26
wire n3174; //IPIN -1 (3,8) #27
wire n3175; //IPIN -1 (3,8) #28
wire n3176; //IPIN -1 (3,8) #29
wire n3177; //IPIN -1 (3,8) #30
wire n3178; //IPIN -1 (3,8) #31
wire n3179; //IPIN -1 (3,8) #32
wire n3180; //IPIN -1 (3,8) #33
wire n3181; //IPIN -1 (3,8) #34
wire n3182; //IPIN -1 (3,8) #35
wire n3183; //IPIN -1 (3,8) #36
wire n3184; //IPIN -1 (3,8) #37
wire n3185; //IPIN -1 (3,8) #38
wire n3186; //IPIN -1 (3,8) #39
wire n3187; //IPIN -1 (3,8) #40
wire n3188; //IPIN -1 (3,8) #41
wire n3189; //IPIN -1 (3,8) #42
wire n3190; //IPIN -1 (3,8) #43
wire n3191; //IPIN -1 (3,8) #44
wire n3192; //IPIN -1 (3,8) #45
wire n3193; //IPIN -1 (3,8) #46
wire n3194; //IPIN -1 (3,8) #47
wire n3195; //IPIN -1 (3,8) #48
wire n3196; //IPIN -1 (3,8) #49
wire n3197; //IPIN -1 (3,8) #50
wire n3198; //IPIN -1 (3,8) #51
wire n3199; //OPIN -1 (3,8) #52
wire n3200; //OPIN -1 (3,8) #53
wire n3201; //OPIN -1 (3,8) #54
wire n3202; //OPIN -1 (3,8) #55
wire n3203; //OPIN -1 (3,8) #56
wire n3204; //OPIN -1 (3,8) #57
wire n3205; //OPIN -1 (3,8) #58
wire n3206; //OPIN -1 (3,8) #59
wire n3207; //OPIN -1 (3,8) #60
wire n3208; //OPIN -1 (3,8) #61
wire n3209; //OPIN -1 (3,8) #62
wire n3210; //OPIN -1 (3,8) #63
wire n3211; //OPIN -1 (3,8) #64
wire n3212; //OPIN -1 (3,8) #65
wire n3213; //OPIN -1 (3,8) #66
wire n3214; //OPIN -1 (3,8) #67
wire n3215; //OPIN -1 (3,8) #68
wire n3216; //OPIN -1 (3,8) #69
wire n3217; //OPIN -1 (3,8) #70
wire n3218; //OPIN -1 (3,8) #71
wire n3219; //IPIN -1 (3,8) #72
wire n3245; //IPIN -1 (3,9) #0
wire n3246; //IPIN -1 (3,9) #1
wire n3247; //IPIN -1 (3,9) #2
wire n3248; //IPIN -1 (3,9) #3
wire n3249; //IPIN -1 (3,9) #4
wire n3250; //IPIN -1 (3,9) #5
wire n3251; //IPIN -1 (3,9) #6
wire n3252; //IPIN -1 (3,9) #7
wire n3253; //IPIN -1 (3,9) #8
wire n3254; //IPIN -1 (3,9) #9
wire n3255; //IPIN -1 (3,9) #10
wire n3256; //IPIN -1 (3,9) #11
wire n3257; //IPIN -1 (3,9) #12
wire n3258; //IPIN -1 (3,9) #13
wire n3259; //IPIN -1 (3,9) #14
wire n3260; //IPIN -1 (3,9) #15
wire n3261; //IPIN -1 (3,9) #16
wire n3262; //IPIN -1 (3,9) #17
wire n3263; //IPIN -1 (3,9) #18
wire n3264; //IPIN -1 (3,9) #19
wire n3265; //IPIN -1 (3,9) #20
wire n3266; //IPIN -1 (3,9) #21
wire n3267; //IPIN -1 (3,9) #22
wire n3268; //IPIN -1 (3,9) #23
wire n3269; //IPIN -1 (3,9) #24
wire n3270; //IPIN -1 (3,9) #25
wire n3271; //IPIN -1 (3,9) #26
wire n3272; //IPIN -1 (3,9) #27
wire n3273; //IPIN -1 (3,9) #28
wire n3274; //IPIN -1 (3,9) #29
wire n3275; //IPIN -1 (3,9) #30
wire n3276; //IPIN -1 (3,9) #31
wire n3277; //IPIN -1 (3,9) #32
wire n3278; //IPIN -1 (3,9) #33
wire n3279; //IPIN -1 (3,9) #34
wire n3280; //IPIN -1 (3,9) #35
wire n3281; //IPIN -1 (3,9) #36
wire n3282; //IPIN -1 (3,9) #37
wire n3283; //IPIN -1 (3,9) #38
wire n3284; //IPIN -1 (3,9) #39
wire n3285; //IPIN -1 (3,9) #40
wire n3286; //IPIN -1 (3,9) #41
wire n3287; //IPIN -1 (3,9) #42
wire n3288; //IPIN -1 (3,9) #43
wire n3289; //IPIN -1 (3,9) #44
wire n3290; //IPIN -1 (3,9) #45
wire n3291; //IPIN -1 (3,9) #46
wire n3292; //IPIN -1 (3,9) #47
wire n3293; //IPIN -1 (3,9) #48
wire n3294; //IPIN -1 (3,9) #49
wire n3295; //IPIN -1 (3,9) #50
wire n3296; //IPIN -1 (3,9) #51
wire n3297; //OPIN -1 (3,9) #52
wire n3298; //OPIN -1 (3,9) #53
wire n3299; //OPIN -1 (3,9) #54
wire n3300; //OPIN -1 (3,9) #55
wire n3301; //OPIN -1 (3,9) #56
wire n3302; //OPIN -1 (3,9) #57
wire n3303; //OPIN -1 (3,9) #58
wire n3304; //OPIN -1 (3,9) #59
wire n3305; //OPIN -1 (3,9) #60
wire n3306; //OPIN -1 (3,9) #61
wire n3307; //OPIN -1 (3,9) #62
wire n3308; //OPIN -1 (3,9) #63
wire n3309; //OPIN -1 (3,9) #64
wire n3310; //OPIN -1 (3,9) #65
wire n3311; //OPIN -1 (3,9) #66
wire n3312; //OPIN -1 (3,9) #67
wire n3313; //OPIN -1 (3,9) #68
wire n3314; //OPIN -1 (3,9) #69
wire n3315; //OPIN -1 (3,9) #70
wire n3316; //OPIN -1 (3,9) #71
wire n3317; //IPIN -1 (3,9) #72
wire n3342; //IPIN -1 (3,10) #0
wire n3343; //OPIN -1 (3,10) #1
wire n3344; //IPIN -1 (3,10) #2
wire n3345; //IPIN -1 (3,10) #3
wire n3346; //OPIN -1 (3,10) #4
wire n3347; //IPIN -1 (3,10) #5
wire n3348; //IPIN -1 (3,10) #6
wire n3349; //OPIN -1 (3,10) #7
wire n3350; //IPIN -1 (3,10) #8
wire n3351; //IPIN -1 (3,10) #9
wire n3352; //OPIN -1 (3,10) #10
wire n3353; //IPIN -1 (3,10) #11
wire n3354; //IPIN -1 (3,10) #12
wire n3355; //OPIN -1 (3,10) #13
wire n3356; //IPIN -1 (3,10) #14
wire n3357; //IPIN -1 (3,10) #15
wire n3358; //OPIN -1 (3,10) #16
wire n3359; //IPIN -1 (3,10) #17
wire n3360; //IPIN -1 (3,10) #18
wire n3361; //OPIN -1 (3,10) #19
wire n3362; //IPIN -1 (3,10) #20
wire n3363; //IPIN -1 (3,10) #21
wire n3364; //OPIN -1 (3,10) #22
wire n3365; //IPIN -1 (3,10) #23
wire n3390; //IPIN -1 (4,0) #0
wire n3391; //OPIN -1 (4,0) #1
wire n3392; //IPIN -1 (4,0) #2
wire n3393; //IPIN -1 (4,0) #3
wire n3394; //OPIN -1 (4,0) #4
wire n3395; //IPIN -1 (4,0) #5
wire n3396; //IPIN -1 (4,0) #6
wire n3397; //OPIN -1 (4,0) #7
wire n3398; //IPIN -1 (4,0) #8
wire n3399; //IPIN -1 (4,0) #9
wire n3400; //OPIN -1 (4,0) #10
wire n3401; //IPIN -1 (4,0) #11
wire n3402; //IPIN -1 (4,0) #12
wire n3403; //OPIN -1 (4,0) #13
wire n3404; //IPIN -1 (4,0) #14
wire n3405; //IPIN -1 (4,0) #15
wire n3406; //OPIN -1 (4,0) #16
wire n3407; //IPIN -1 (4,0) #17
wire n3408; //IPIN -1 (4,0) #18
wire n3409; //OPIN -1 (4,0) #19
wire n3410; //IPIN -1 (4,0) #20
wire n3411; //IPIN -1 (4,0) #21
wire n3412; //OPIN -1 (4,0) #22
wire n3413; //IPIN -1 (4,0) #23
wire n3439; //IPIN -1 (4,1) #0
wire n3440; //IPIN -1 (4,1) #1
wire n3441; //IPIN -1 (4,1) #2
wire n3442; //IPIN -1 (4,1) #3
wire n3443; //IPIN -1 (4,1) #4
wire n3444; //IPIN -1 (4,1) #5
wire n3445; //IPIN -1 (4,1) #6
wire n3446; //IPIN -1 (4,1) #7
wire n3447; //IPIN -1 (4,1) #8
wire n3448; //IPIN -1 (4,1) #9
wire n3449; //IPIN -1 (4,1) #10
wire n3450; //IPIN -1 (4,1) #11
wire n3451; //IPIN -1 (4,1) #12
wire n3452; //IPIN -1 (4,1) #13
wire n3453; //IPIN -1 (4,1) #14
wire n3454; //IPIN -1 (4,1) #15
wire n3455; //IPIN -1 (4,1) #16
wire n3456; //IPIN -1 (4,1) #17
wire n3457; //IPIN -1 (4,1) #18
wire n3458; //IPIN -1 (4,1) #19
wire n3459; //IPIN -1 (4,1) #20
wire n3460; //IPIN -1 (4,1) #21
wire n3461; //IPIN -1 (4,1) #22
wire n3462; //IPIN -1 (4,1) #23
wire n3463; //IPIN -1 (4,1) #24
wire n3464; //IPIN -1 (4,1) #25
wire n3465; //IPIN -1 (4,1) #26
wire n3466; //IPIN -1 (4,1) #27
wire n3467; //IPIN -1 (4,1) #28
wire n3468; //IPIN -1 (4,1) #29
wire n3469; //IPIN -1 (4,1) #30
wire n3470; //IPIN -1 (4,1) #31
wire n3471; //IPIN -1 (4,1) #32
wire n3472; //IPIN -1 (4,1) #33
wire n3473; //IPIN -1 (4,1) #34
wire n3474; //IPIN -1 (4,1) #35
wire n3475; //IPIN -1 (4,1) #36
wire n3476; //IPIN -1 (4,1) #37
wire n3477; //IPIN -1 (4,1) #38
wire n3478; //IPIN -1 (4,1) #39
wire n3479; //IPIN -1 (4,1) #40
wire n3480; //IPIN -1 (4,1) #41
wire n3481; //IPIN -1 (4,1) #42
wire n3482; //IPIN -1 (4,1) #43
wire n3483; //IPIN -1 (4,1) #44
wire n3484; //IPIN -1 (4,1) #45
wire n3485; //IPIN -1 (4,1) #46
wire n3486; //IPIN -1 (4,1) #47
wire n3487; //IPIN -1 (4,1) #48
wire n3488; //IPIN -1 (4,1) #49
wire n3489; //IPIN -1 (4,1) #50
wire n3490; //IPIN -1 (4,1) #51
wire n3491; //OPIN -1 (4,1) #52
wire n3492; //OPIN -1 (4,1) #53
wire n3493; //OPIN -1 (4,1) #54
wire n3494; //OPIN -1 (4,1) #55
wire n3495; //OPIN -1 (4,1) #56
wire n3496; //OPIN -1 (4,1) #57
wire n3497; //OPIN -1 (4,1) #58
wire n3498; //OPIN -1 (4,1) #59
wire n3499; //OPIN -1 (4,1) #60
wire n3500; //OPIN -1 (4,1) #61
wire n3501; //OPIN -1 (4,1) #62
wire n3502; //OPIN -1 (4,1) #63
wire n3503; //OPIN -1 (4,1) #64
wire n3504; //OPIN -1 (4,1) #65
wire n3505; //OPIN -1 (4,1) #66
wire n3506; //OPIN -1 (4,1) #67
wire n3507; //OPIN -1 (4,1) #68
wire n3508; //OPIN -1 (4,1) #69
wire n3509; //OPIN -1 (4,1) #70
wire n3510; //OPIN -1 (4,1) #71
wire n3511; //IPIN -1 (4,1) #72
wire n3537; //IPIN -1 (4,2) #0
wire n3538; //IPIN -1 (4,2) #1
wire n3539; //IPIN -1 (4,2) #2
wire n3540; //IPIN -1 (4,2) #3
wire n3541; //IPIN -1 (4,2) #4
wire n3542; //IPIN -1 (4,2) #5
wire n3543; //IPIN -1 (4,2) #6
wire n3544; //IPIN -1 (4,2) #7
wire n3545; //IPIN -1 (4,2) #8
wire n3546; //IPIN -1 (4,2) #9
wire n3547; //IPIN -1 (4,2) #10
wire n3548; //IPIN -1 (4,2) #11
wire n3549; //IPIN -1 (4,2) #12
wire n3550; //IPIN -1 (4,2) #13
wire n3551; //IPIN -1 (4,2) #14
wire n3552; //IPIN -1 (4,2) #15
wire n3553; //IPIN -1 (4,2) #16
wire n3554; //IPIN -1 (4,2) #17
wire n3555; //IPIN -1 (4,2) #18
wire n3556; //IPIN -1 (4,2) #19
wire n3557; //IPIN -1 (4,2) #20
wire n3558; //IPIN -1 (4,2) #21
wire n3559; //IPIN -1 (4,2) #22
wire n3560; //IPIN -1 (4,2) #23
wire n3561; //IPIN -1 (4,2) #24
wire n3562; //IPIN -1 (4,2) #25
wire n3563; //IPIN -1 (4,2) #26
wire n3564; //IPIN -1 (4,2) #27
wire n3565; //IPIN -1 (4,2) #28
wire n3566; //IPIN -1 (4,2) #29
wire n3567; //IPIN -1 (4,2) #30
wire n3568; //IPIN -1 (4,2) #31
wire n3569; //IPIN -1 (4,2) #32
wire n3570; //IPIN -1 (4,2) #33
wire n3571; //IPIN -1 (4,2) #34
wire n3572; //IPIN -1 (4,2) #35
wire n3573; //IPIN -1 (4,2) #36
wire n3574; //IPIN -1 (4,2) #37
wire n3575; //IPIN -1 (4,2) #38
wire n3576; //IPIN -1 (4,2) #39
wire n3577; //IPIN -1 (4,2) #40
wire n3578; //IPIN -1 (4,2) #41
wire n3579; //IPIN -1 (4,2) #42
wire n3580; //IPIN -1 (4,2) #43
wire n3581; //IPIN -1 (4,2) #44
wire n3582; //IPIN -1 (4,2) #45
wire n3583; //IPIN -1 (4,2) #46
wire n3584; //IPIN -1 (4,2) #47
wire n3585; //IPIN -1 (4,2) #48
wire n3586; //IPIN -1 (4,2) #49
wire n3587; //IPIN -1 (4,2) #50
wire n3588; //IPIN -1 (4,2) #51
wire n3589; //OPIN -1 (4,2) #52
wire n3590; //OPIN -1 (4,2) #53
wire n3591; //OPIN -1 (4,2) #54
wire n3592; //OPIN -1 (4,2) #55
wire n3593; //OPIN -1 (4,2) #56
wire n3594; //OPIN -1 (4,2) #57
wire n3595; //OPIN -1 (4,2) #58
wire n3596; //OPIN -1 (4,2) #59
wire n3597; //OPIN -1 (4,2) #60
wire n3598; //OPIN -1 (4,2) #61
wire n3599; //OPIN -1 (4,2) #62
wire n3600; //OPIN -1 (4,2) #63
wire n3601; //OPIN -1 (4,2) #64
wire n3602; //OPIN -1 (4,2) #65
wire n3603; //OPIN -1 (4,2) #66
wire n3604; //OPIN -1 (4,2) #67
wire n3605; //OPIN -1 (4,2) #68
wire n3606; //OPIN -1 (4,2) #69
wire n3607; //OPIN -1 (4,2) #70
wire n3608; //OPIN -1 (4,2) #71
wire n3609; //IPIN -1 (4,2) #72
wire n3635; //IPIN -1 (4,3) #0
wire n3636; //IPIN -1 (4,3) #1
wire n3637; //IPIN -1 (4,3) #2
wire n3638; //IPIN -1 (4,3) #3
wire n3639; //IPIN -1 (4,3) #4
wire n3640; //IPIN -1 (4,3) #5
wire n3641; //IPIN -1 (4,3) #6
wire n3642; //IPIN -1 (4,3) #7
wire n3643; //IPIN -1 (4,3) #8
wire n3644; //IPIN -1 (4,3) #9
wire n3645; //IPIN -1 (4,3) #10
wire n3646; //IPIN -1 (4,3) #11
wire n3647; //IPIN -1 (4,3) #12
wire n3648; //IPIN -1 (4,3) #13
wire n3649; //IPIN -1 (4,3) #14
wire n3650; //IPIN -1 (4,3) #15
wire n3651; //IPIN -1 (4,3) #16
wire n3652; //IPIN -1 (4,3) #17
wire n3653; //IPIN -1 (4,3) #18
wire n3654; //IPIN -1 (4,3) #19
wire n3655; //IPIN -1 (4,3) #20
wire n3656; //IPIN -1 (4,3) #21
wire n3657; //IPIN -1 (4,3) #22
wire n3658; //IPIN -1 (4,3) #23
wire n3659; //IPIN -1 (4,3) #24
wire n3660; //IPIN -1 (4,3) #25
wire n3661; //IPIN -1 (4,3) #26
wire n3662; //IPIN -1 (4,3) #27
wire n3663; //IPIN -1 (4,3) #28
wire n3664; //IPIN -1 (4,3) #29
wire n3665; //IPIN -1 (4,3) #30
wire n3666; //IPIN -1 (4,3) #31
wire n3667; //IPIN -1 (4,3) #32
wire n3668; //IPIN -1 (4,3) #33
wire n3669; //IPIN -1 (4,3) #34
wire n3670; //IPIN -1 (4,3) #35
wire n3671; //IPIN -1 (4,3) #36
wire n3672; //IPIN -1 (4,3) #37
wire n3673; //IPIN -1 (4,3) #38
wire n3674; //IPIN -1 (4,3) #39
wire n3675; //IPIN -1 (4,3) #40
wire n3676; //IPIN -1 (4,3) #41
wire n3677; //IPIN -1 (4,3) #42
wire n3678; //IPIN -1 (4,3) #43
wire n3679; //IPIN -1 (4,3) #44
wire n3680; //IPIN -1 (4,3) #45
wire n3681; //IPIN -1 (4,3) #46
wire n3682; //IPIN -1 (4,3) #47
wire n3683; //IPIN -1 (4,3) #48
wire n3684; //IPIN -1 (4,3) #49
wire n3685; //IPIN -1 (4,3) #50
wire n3686; //IPIN -1 (4,3) #51
wire n3687; //OPIN -1 (4,3) #52
wire n3688; //OPIN -1 (4,3) #53
wire n3689; //OPIN -1 (4,3) #54
wire n3690; //OPIN -1 (4,3) #55
wire n3691; //OPIN -1 (4,3) #56
wire n3692; //OPIN -1 (4,3) #57
wire n3693; //OPIN -1 (4,3) #58
wire n3694; //OPIN -1 (4,3) #59
wire n3695; //OPIN -1 (4,3) #60
wire n3696; //OPIN -1 (4,3) #61
wire n3697; //OPIN -1 (4,3) #62
wire n3698; //OPIN -1 (4,3) #63
wire n3699; //OPIN -1 (4,3) #64
wire n3700; //OPIN -1 (4,3) #65
wire n3701; //OPIN -1 (4,3) #66
wire n3702; //OPIN -1 (4,3) #67
wire n3703; //OPIN -1 (4,3) #68
wire n3704; //OPIN -1 (4,3) #69
wire n3705; //OPIN -1 (4,3) #70
wire n3706; //OPIN -1 (4,3) #71
wire n3707; //IPIN -1 (4,3) #72
wire n3733; //IPIN -1 (4,4) #0
wire n3734; //IPIN -1 (4,4) #1
wire n3735; //IPIN -1 (4,4) #2
wire n3736; //IPIN -1 (4,4) #3
wire n3737; //IPIN -1 (4,4) #4
wire n3738; //IPIN -1 (4,4) #5
wire n3739; //IPIN -1 (4,4) #6
wire n3740; //IPIN -1 (4,4) #7
wire n3741; //IPIN -1 (4,4) #8
wire n3742; //IPIN -1 (4,4) #9
wire n3743; //IPIN -1 (4,4) #10
wire n3744; //IPIN -1 (4,4) #11
wire n3745; //IPIN -1 (4,4) #12
wire n3746; //IPIN -1 (4,4) #13
wire n3747; //IPIN -1 (4,4) #14
wire n3748; //IPIN -1 (4,4) #15
wire n3749; //IPIN -1 (4,4) #16
wire n3750; //IPIN -1 (4,4) #17
wire n3751; //IPIN -1 (4,4) #18
wire n3752; //IPIN -1 (4,4) #19
wire n3753; //IPIN -1 (4,4) #20
wire n3754; //IPIN -1 (4,4) #21
wire n3755; //IPIN -1 (4,4) #22
wire n3756; //IPIN -1 (4,4) #23
wire n3757; //IPIN -1 (4,4) #24
wire n3758; //IPIN -1 (4,4) #25
wire n3759; //IPIN -1 (4,4) #26
wire n3760; //IPIN -1 (4,4) #27
wire n3761; //IPIN -1 (4,4) #28
wire n3762; //IPIN -1 (4,4) #29
wire n3763; //IPIN -1 (4,4) #30
wire n3764; //IPIN -1 (4,4) #31
wire n3765; //IPIN -1 (4,4) #32
wire n3766; //IPIN -1 (4,4) #33
wire n3767; //IPIN -1 (4,4) #34
wire n3768; //IPIN -1 (4,4) #35
wire n3769; //IPIN -1 (4,4) #36
wire n3770; //IPIN -1 (4,4) #37
wire n3771; //IPIN -1 (4,4) #38
wire n3772; //IPIN -1 (4,4) #39
wire n3773; //IPIN -1 (4,4) #40
wire n3774; //IPIN -1 (4,4) #41
wire n3775; //IPIN -1 (4,4) #42
wire n3776; //IPIN -1 (4,4) #43
wire n3777; //IPIN -1 (4,4) #44
wire n3778; //IPIN -1 (4,4) #45
wire n3779; //IPIN -1 (4,4) #46
wire n3780; //IPIN -1 (4,4) #47
wire n3781; //IPIN -1 (4,4) #48
wire n3782; //IPIN -1 (4,4) #49
wire n3783; //IPIN -1 (4,4) #50
wire n3784; //IPIN -1 (4,4) #51
wire n3785; //OPIN -1 (4,4) #52
wire n3786; //OPIN -1 (4,4) #53
wire n3787; //OPIN -1 (4,4) #54
wire n3788; //OPIN -1 (4,4) #55
wire n3789; //OPIN -1 (4,4) #56
wire n3790; //OPIN -1 (4,4) #57
wire n3791; //OPIN -1 (4,4) #58
wire n3792; //OPIN -1 (4,4) #59
wire n3793; //OPIN -1 (4,4) #60
wire n3794; //OPIN -1 (4,4) #61
wire n3795; //OPIN -1 (4,4) #62
wire n3796; //OPIN -1 (4,4) #63
wire n3797; //OPIN -1 (4,4) #64
wire n3798; //OPIN -1 (4,4) #65
wire n3799; //OPIN -1 (4,4) #66
wire n3800; //OPIN -1 (4,4) #67
wire n3801; //OPIN -1 (4,4) #68
wire n3802; //OPIN -1 (4,4) #69
wire n3803; //OPIN -1 (4,4) #70
wire n3804; //OPIN -1 (4,4) #71
wire n3805; //IPIN -1 (4,4) #72
wire n3831; //IPIN -1 (4,5) #0
wire n3832; //IPIN -1 (4,5) #1
wire n3833; //IPIN -1 (4,5) #2
wire n3834; //IPIN -1 (4,5) #3
wire n3835; //IPIN -1 (4,5) #4
wire n3836; //IPIN -1 (4,5) #5
wire n3837; //IPIN -1 (4,5) #6
wire n3838; //IPIN -1 (4,5) #7
wire n3839; //IPIN -1 (4,5) #8
wire n3840; //IPIN -1 (4,5) #9
wire n3841; //IPIN -1 (4,5) #10
wire n3842; //IPIN -1 (4,5) #11
wire n3843; //IPIN -1 (4,5) #12
wire n3844; //IPIN -1 (4,5) #13
wire n3845; //IPIN -1 (4,5) #14
wire n3846; //IPIN -1 (4,5) #15
wire n3847; //IPIN -1 (4,5) #16
wire n3848; //IPIN -1 (4,5) #17
wire n3849; //IPIN -1 (4,5) #18
wire n3850; //IPIN -1 (4,5) #19
wire n3851; //IPIN -1 (4,5) #20
wire n3852; //IPIN -1 (4,5) #21
wire n3853; //IPIN -1 (4,5) #22
wire n3854; //IPIN -1 (4,5) #23
wire n3855; //IPIN -1 (4,5) #24
wire n3856; //IPIN -1 (4,5) #25
wire n3857; //IPIN -1 (4,5) #26
wire n3858; //IPIN -1 (4,5) #27
wire n3859; //IPIN -1 (4,5) #28
wire n3860; //IPIN -1 (4,5) #29
wire n3861; //IPIN -1 (4,5) #30
wire n3862; //IPIN -1 (4,5) #31
wire n3863; //IPIN -1 (4,5) #32
wire n3864; //IPIN -1 (4,5) #33
wire n3865; //IPIN -1 (4,5) #34
wire n3866; //IPIN -1 (4,5) #35
wire n3867; //IPIN -1 (4,5) #36
wire n3868; //IPIN -1 (4,5) #37
wire n3869; //IPIN -1 (4,5) #38
wire n3870; //IPIN -1 (4,5) #39
wire n3871; //IPIN -1 (4,5) #40
wire n3872; //IPIN -1 (4,5) #41
wire n3873; //IPIN -1 (4,5) #42
wire n3874; //IPIN -1 (4,5) #43
wire n3875; //IPIN -1 (4,5) #44
wire n3876; //IPIN -1 (4,5) #45
wire n3877; //IPIN -1 (4,5) #46
wire n3878; //IPIN -1 (4,5) #47
wire n3879; //IPIN -1 (4,5) #48
wire n3880; //IPIN -1 (4,5) #49
wire n3881; //IPIN -1 (4,5) #50
wire n3882; //IPIN -1 (4,5) #51
wire n3883; //OPIN -1 (4,5) #52
wire n3884; //OPIN -1 (4,5) #53
wire n3885; //OPIN -1 (4,5) #54
wire n3886; //OPIN -1 (4,5) #55
wire n3887; //OPIN -1 (4,5) #56
wire n3888; //OPIN -1 (4,5) #57
wire n3889; //OPIN -1 (4,5) #58
wire n3890; //OPIN -1 (4,5) #59
wire n3891; //OPIN -1 (4,5) #60
wire n3892; //OPIN -1 (4,5) #61
wire n3893; //OPIN -1 (4,5) #62
wire n3894; //OPIN -1 (4,5) #63
wire n3895; //OPIN -1 (4,5) #64
wire n3896; //OPIN -1 (4,5) #65
wire n3897; //OPIN -1 (4,5) #66
wire n3898; //OPIN -1 (4,5) #67
wire n3899; //OPIN -1 (4,5) #68
wire n3900; //OPIN -1 (4,5) #69
wire n3901; //OPIN -1 (4,5) #70
wire n3902; //OPIN -1 (4,5) #71
wire n3903; //IPIN -1 (4,5) #72
wire n3929; //IPIN -1 (4,6) #0
wire n3930; //IPIN -1 (4,6) #1
wire n3931; //IPIN -1 (4,6) #2
wire n3932; //IPIN -1 (4,6) #3
wire n3933; //IPIN -1 (4,6) #4
wire n3934; //IPIN -1 (4,6) #5
wire n3935; //IPIN -1 (4,6) #6
wire n3936; //IPIN -1 (4,6) #7
wire n3937; //IPIN -1 (4,6) #8
wire n3938; //IPIN -1 (4,6) #9
wire n3939; //IPIN -1 (4,6) #10
wire n3940; //IPIN -1 (4,6) #11
wire n3941; //IPIN -1 (4,6) #12
wire n3942; //IPIN -1 (4,6) #13
wire n3943; //IPIN -1 (4,6) #14
wire n3944; //IPIN -1 (4,6) #15
wire n3945; //IPIN -1 (4,6) #16
wire n3946; //IPIN -1 (4,6) #17
wire n3947; //IPIN -1 (4,6) #18
wire n3948; //IPIN -1 (4,6) #19
wire n3949; //IPIN -1 (4,6) #20
wire n3950; //IPIN -1 (4,6) #21
wire n3951; //IPIN -1 (4,6) #22
wire n3952; //IPIN -1 (4,6) #23
wire n3953; //IPIN -1 (4,6) #24
wire n3954; //IPIN -1 (4,6) #25
wire n3955; //IPIN -1 (4,6) #26
wire n3956; //IPIN -1 (4,6) #27
wire n3957; //IPIN -1 (4,6) #28
wire n3958; //IPIN -1 (4,6) #29
wire n3959; //IPIN -1 (4,6) #30
wire n3960; //IPIN -1 (4,6) #31
wire n3961; //IPIN -1 (4,6) #32
wire n3962; //IPIN -1 (4,6) #33
wire n3963; //IPIN -1 (4,6) #34
wire n3964; //IPIN -1 (4,6) #35
wire n3965; //IPIN -1 (4,6) #36
wire n3966; //IPIN -1 (4,6) #37
wire n3967; //IPIN -1 (4,6) #38
wire n3968; //IPIN -1 (4,6) #39
wire n3969; //IPIN -1 (4,6) #40
wire n3970; //IPIN -1 (4,6) #41
wire n3971; //IPIN -1 (4,6) #42
wire n3972; //IPIN -1 (4,6) #43
wire n3973; //IPIN -1 (4,6) #44
wire n3974; //IPIN -1 (4,6) #45
wire n3975; //IPIN -1 (4,6) #46
wire n3976; //IPIN -1 (4,6) #47
wire n3977; //IPIN -1 (4,6) #48
wire n3978; //IPIN -1 (4,6) #49
wire n3979; //IPIN -1 (4,6) #50
wire n3980; //IPIN -1 (4,6) #51
wire n3981; //OPIN -1 (4,6) #52
wire n3982; //OPIN -1 (4,6) #53
wire n3983; //OPIN -1 (4,6) #54
wire n3984; //OPIN -1 (4,6) #55
wire n3985; //OPIN -1 (4,6) #56
wire n3986; //OPIN -1 (4,6) #57
wire n3987; //OPIN -1 (4,6) #58
wire n3988; //OPIN -1 (4,6) #59
wire n3989; //OPIN -1 (4,6) #60
wire n3990; //OPIN -1 (4,6) #61
wire n3991; //OPIN -1 (4,6) #62
wire n3992; //OPIN -1 (4,6) #63
wire n3993; //OPIN -1 (4,6) #64
wire n3994; //OPIN -1 (4,6) #65
wire n3995; //OPIN -1 (4,6) #66
wire n3996; //OPIN -1 (4,6) #67
wire n3997; //OPIN -1 (4,6) #68
wire n3998; //OPIN -1 (4,6) #69
wire n3999; //OPIN -1 (4,6) #70
wire n4000; //OPIN -1 (4,6) #71
wire n4001; //IPIN -1 (4,6) #72
wire n4027; //IPIN -1 (4,7) #0
wire n4028; //IPIN -1 (4,7) #1
wire n4029; //IPIN -1 (4,7) #2
wire n4030; //IPIN -1 (4,7) #3
wire n4031; //IPIN -1 (4,7) #4
wire n4032; //IPIN -1 (4,7) #5
wire n4033; //IPIN -1 (4,7) #6
wire n4034; //IPIN -1 (4,7) #7
wire n4035; //IPIN -1 (4,7) #8
wire n4036; //IPIN -1 (4,7) #9
wire n4037; //IPIN -1 (4,7) #10
wire n4038; //IPIN -1 (4,7) #11
wire n4039; //IPIN -1 (4,7) #12
wire n4040; //IPIN -1 (4,7) #13
wire n4041; //IPIN -1 (4,7) #14
wire n4042; //IPIN -1 (4,7) #15
wire n4043; //IPIN -1 (4,7) #16
wire n4044; //IPIN -1 (4,7) #17
wire n4045; //IPIN -1 (4,7) #18
wire n4046; //IPIN -1 (4,7) #19
wire n4047; //IPIN -1 (4,7) #20
wire n4048; //IPIN -1 (4,7) #21
wire n4049; //IPIN -1 (4,7) #22
wire n4050; //IPIN -1 (4,7) #23
wire n4051; //IPIN -1 (4,7) #24
wire n4052; //IPIN -1 (4,7) #25
wire n4053; //IPIN -1 (4,7) #26
wire n4054; //IPIN -1 (4,7) #27
wire n4055; //IPIN -1 (4,7) #28
wire n4056; //IPIN -1 (4,7) #29
wire n4057; //IPIN -1 (4,7) #30
wire n4058; //IPIN -1 (4,7) #31
wire n4059; //IPIN -1 (4,7) #32
wire n4060; //IPIN -1 (4,7) #33
wire n4061; //IPIN -1 (4,7) #34
wire n4062; //IPIN -1 (4,7) #35
wire n4063; //IPIN -1 (4,7) #36
wire n4064; //IPIN -1 (4,7) #37
wire n4065; //IPIN -1 (4,7) #38
wire n4066; //IPIN -1 (4,7) #39
wire n4067; //IPIN -1 (4,7) #40
wire n4068; //IPIN -1 (4,7) #41
wire n4069; //IPIN -1 (4,7) #42
wire n4070; //IPIN -1 (4,7) #43
wire n4071; //IPIN -1 (4,7) #44
wire n4072; //IPIN -1 (4,7) #45
wire n4073; //IPIN -1 (4,7) #46
wire n4074; //IPIN -1 (4,7) #47
wire n4075; //IPIN -1 (4,7) #48
wire n4076; //IPIN -1 (4,7) #49
wire n4077; //IPIN -1 (4,7) #50
wire n4078; //IPIN -1 (4,7) #51
wire n4079; //OPIN -1 (4,7) #52
wire n4080; //OPIN -1 (4,7) #53
wire n4081; //OPIN -1 (4,7) #54
wire n4082; //OPIN -1 (4,7) #55
wire n4083; //OPIN -1 (4,7) #56
wire n4084; //OPIN -1 (4,7) #57
wire n4085; //OPIN -1 (4,7) #58
wire n4086; //OPIN -1 (4,7) #59
wire n4087; //OPIN -1 (4,7) #60
wire n4088; //OPIN -1 (4,7) #61
wire n4089; //OPIN -1 (4,7) #62
wire n4090; //OPIN -1 (4,7) #63
wire n4091; //OPIN -1 (4,7) #64
wire n4092; //OPIN -1 (4,7) #65
wire n4093; //OPIN -1 (4,7) #66
wire n4094; //OPIN -1 (4,7) #67
wire n4095; //OPIN -1 (4,7) #68
wire n4096; //OPIN -1 (4,7) #69
wire n4097; //OPIN -1 (4,7) #70
wire n4098; //OPIN -1 (4,7) #71
wire n4099; //IPIN -1 (4,7) #72
wire n4125; //IPIN -1 (4,8) #0
wire n4126; //IPIN -1 (4,8) #1
wire n4127; //IPIN -1 (4,8) #2
wire n4128; //IPIN -1 (4,8) #3
wire n4129; //IPIN -1 (4,8) #4
wire n4130; //IPIN -1 (4,8) #5
wire n4131; //IPIN -1 (4,8) #6
wire n4132; //IPIN -1 (4,8) #7
wire n4133; //IPIN -1 (4,8) #8
wire n4134; //IPIN -1 (4,8) #9
wire n4135; //IPIN -1 (4,8) #10
wire n4136; //IPIN -1 (4,8) #11
wire n4137; //IPIN -1 (4,8) #12
wire n4138; //IPIN -1 (4,8) #13
wire n4139; //IPIN -1 (4,8) #14
wire n4140; //IPIN -1 (4,8) #15
wire n4141; //IPIN -1 (4,8) #16
wire n4142; //IPIN -1 (4,8) #17
wire n4143; //IPIN -1 (4,8) #18
wire n4144; //IPIN -1 (4,8) #19
wire n4145; //IPIN -1 (4,8) #20
wire n4146; //IPIN -1 (4,8) #21
wire n4147; //IPIN -1 (4,8) #22
wire n4148; //IPIN -1 (4,8) #23
wire n4149; //IPIN -1 (4,8) #24
wire n4150; //IPIN -1 (4,8) #25
wire n4151; //IPIN -1 (4,8) #26
wire n4152; //IPIN -1 (4,8) #27
wire n4153; //IPIN -1 (4,8) #28
wire n4154; //IPIN -1 (4,8) #29
wire n4155; //IPIN -1 (4,8) #30
wire n4156; //IPIN -1 (4,8) #31
wire n4157; //IPIN -1 (4,8) #32
wire n4158; //IPIN -1 (4,8) #33
wire n4159; //IPIN -1 (4,8) #34
wire n4160; //IPIN -1 (4,8) #35
wire n4161; //IPIN -1 (4,8) #36
wire n4162; //IPIN -1 (4,8) #37
wire n4163; //IPIN -1 (4,8) #38
wire n4164; //IPIN -1 (4,8) #39
wire n4165; //IPIN -1 (4,8) #40
wire n4166; //IPIN -1 (4,8) #41
wire n4167; //IPIN -1 (4,8) #42
wire n4168; //IPIN -1 (4,8) #43
wire n4169; //IPIN -1 (4,8) #44
wire n4170; //IPIN -1 (4,8) #45
wire n4171; //IPIN -1 (4,8) #46
wire n4172; //IPIN -1 (4,8) #47
wire n4173; //IPIN -1 (4,8) #48
wire n4174; //IPIN -1 (4,8) #49
wire n4175; //IPIN -1 (4,8) #50
wire n4176; //IPIN -1 (4,8) #51
wire n4177; //OPIN -1 (4,8) #52
wire n4178; //OPIN -1 (4,8) #53
wire n4179; //OPIN -1 (4,8) #54
wire n4180; //OPIN -1 (4,8) #55
wire n4181; //OPIN -1 (4,8) #56
wire n4182; //OPIN -1 (4,8) #57
wire n4183; //OPIN -1 (4,8) #58
wire n4184; //OPIN -1 (4,8) #59
wire n4185; //OPIN -1 (4,8) #60
wire n4186; //OPIN -1 (4,8) #61
wire n4187; //OPIN -1 (4,8) #62
wire n4188; //OPIN -1 (4,8) #63
wire n4189; //OPIN -1 (4,8) #64
wire n4190; //OPIN -1 (4,8) #65
wire n4191; //OPIN -1 (4,8) #66
wire n4192; //OPIN -1 (4,8) #67
wire n4193; //OPIN -1 (4,8) #68
wire n4194; //OPIN -1 (4,8) #69
wire n4195; //OPIN -1 (4,8) #70
wire n4196; //OPIN -1 (4,8) #71
wire n4197; //IPIN -1 (4,8) #72
wire n4223; //IPIN -1 (4,9) #0
wire n4224; //IPIN -1 (4,9) #1
wire n4225; //IPIN -1 (4,9) #2
wire n4226; //IPIN -1 (4,9) #3
wire n4227; //IPIN -1 (4,9) #4
wire n4228; //IPIN -1 (4,9) #5
wire n4229; //IPIN -1 (4,9) #6
wire n4230; //IPIN -1 (4,9) #7
wire n4231; //IPIN -1 (4,9) #8
wire n4232; //IPIN -1 (4,9) #9
wire n4233; //IPIN -1 (4,9) #10
wire n4234; //IPIN -1 (4,9) #11
wire n4235; //IPIN -1 (4,9) #12
wire n4236; //IPIN -1 (4,9) #13
wire n4237; //IPIN -1 (4,9) #14
wire n4238; //IPIN -1 (4,9) #15
wire n4239; //IPIN -1 (4,9) #16
wire n4240; //IPIN -1 (4,9) #17
wire n4241; //IPIN -1 (4,9) #18
wire n4242; //IPIN -1 (4,9) #19
wire n4243; //IPIN -1 (4,9) #20
wire n4244; //IPIN -1 (4,9) #21
wire n4245; //IPIN -1 (4,9) #22
wire n4246; //IPIN -1 (4,9) #23
wire n4247; //IPIN -1 (4,9) #24
wire n4248; //IPIN -1 (4,9) #25
wire n4249; //IPIN -1 (4,9) #26
wire n4250; //IPIN -1 (4,9) #27
wire n4251; //IPIN -1 (4,9) #28
wire n4252; //IPIN -1 (4,9) #29
wire n4253; //IPIN -1 (4,9) #30
wire n4254; //IPIN -1 (4,9) #31
wire n4255; //IPIN -1 (4,9) #32
wire n4256; //IPIN -1 (4,9) #33
wire n4257; //IPIN -1 (4,9) #34
wire n4258; //IPIN -1 (4,9) #35
wire n4259; //IPIN -1 (4,9) #36
wire n4260; //IPIN -1 (4,9) #37
wire n4261; //IPIN -1 (4,9) #38
wire n4262; //IPIN -1 (4,9) #39
wire n4263; //IPIN -1 (4,9) #40
wire n4264; //IPIN -1 (4,9) #41
wire n4265; //IPIN -1 (4,9) #42
wire n4266; //IPIN -1 (4,9) #43
wire n4267; //IPIN -1 (4,9) #44
wire n4268; //IPIN -1 (4,9) #45
wire n4269; //IPIN -1 (4,9) #46
wire n4270; //IPIN -1 (4,9) #47
wire n4271; //IPIN -1 (4,9) #48
wire n4272; //IPIN -1 (4,9) #49
wire n4273; //IPIN -1 (4,9) #50
wire n4274; //IPIN -1 (4,9) #51
wire n4275; //OPIN -1 (4,9) #52
wire n4276; //OPIN -1 (4,9) #53
wire n4277; //OPIN -1 (4,9) #54
wire n4278; //OPIN -1 (4,9) #55
wire n4279; //OPIN -1 (4,9) #56
wire n4280; //OPIN -1 (4,9) #57
wire n4281; //OPIN -1 (4,9) #58
wire n4282; //OPIN -1 (4,9) #59
wire n4283; //OPIN -1 (4,9) #60
wire n4284; //OPIN -1 (4,9) #61
wire n4285; //OPIN -1 (4,9) #62
wire n4286; //OPIN -1 (4,9) #63
wire n4287; //OPIN -1 (4,9) #64
wire n4288; //OPIN -1 (4,9) #65
wire n4289; //OPIN -1 (4,9) #66
wire n4290; //OPIN -1 (4,9) #67
wire n4291; //OPIN -1 (4,9) #68
wire n4292; //OPIN -1 (4,9) #69
wire n4293; //OPIN -1 (4,9) #70
wire n4294; //OPIN -1 (4,9) #71
wire n4295; //IPIN -1 (4,9) #72
wire n4320; //IPIN -1 (4,10) #0
wire n4321; //OPIN -1 (4,10) #1
wire n4322; //IPIN -1 (4,10) #2
wire n4323; //IPIN -1 (4,10) #3
wire n4324; //OPIN -1 (4,10) #4
wire n4325; //IPIN -1 (4,10) #5
wire n4326; //IPIN -1 (4,10) #6
wire n4327; //OPIN -1 (4,10) #7
wire n4328; //IPIN -1 (4,10) #8
wire n4329; //IPIN -1 (4,10) #9
wire n4330; //OPIN -1 (4,10) #10
wire n4331; //IPIN -1 (4,10) #11
wire n4332; //IPIN -1 (4,10) #12
wire n4333; //OPIN -1 (4,10) #13
wire n4334; //IPIN -1 (4,10) #14
wire n4335; //IPIN -1 (4,10) #15
wire n4336; //OPIN -1 (4,10) #16
wire n4337; //IPIN -1 (4,10) #17
wire n4338; //IPIN -1 (4,10) #18
wire n4339; //OPIN -1 (4,10) #19
wire n4340; //IPIN -1 (4,10) #20
wire n4341; //IPIN -1 (4,10) #21
wire n4342; //OPIN -1 (4,10) #22
wire n4343; //IPIN -1 (4,10) #23
wire n4368; //IPIN -1 (5,0) #0
wire n4369; //OPIN -1 (5,0) #1
wire n4370; //IPIN -1 (5,0) #2
wire n4371; //IPIN -1 (5,0) #3
wire n4372; //OPIN -1 (5,0) #4
wire n4373; //IPIN -1 (5,0) #5
wire n4374; //IPIN -1 (5,0) #6
wire n4375; //OPIN -1 (5,0) #7
wire n4376; //IPIN -1 (5,0) #8
wire n4377; //IPIN -1 (5,0) #9
wire n4378; //OPIN -1 (5,0) #10
wire n4379; //IPIN -1 (5,0) #11
wire n4380; //IPIN -1 (5,0) #12
wire n4381; //OPIN -1 (5,0) #13
wire n4382; //IPIN -1 (5,0) #14
wire n4383; //IPIN -1 (5,0) #15
wire n4384; //OPIN -1 (5,0) #16
wire n4385; //IPIN -1 (5,0) #17
wire n4386; //IPIN -1 (5,0) #18
wire n4387; //OPIN -1 (5,0) #19
wire n4388; //IPIN -1 (5,0) #20
wire n4389; //IPIN -1 (5,0) #21
wire n4390; //OPIN -1 (5,0) #22
wire n4391; //IPIN -1 (5,0) #23
wire n4417; //IPIN -1 (5,1) #0
wire n4418; //IPIN -1 (5,1) #1
wire n4419; //IPIN -1 (5,1) #2
wire n4420; //IPIN -1 (5,1) #3
wire n4421; //IPIN -1 (5,1) #4
wire n4422; //IPIN -1 (5,1) #5
wire n4423; //IPIN -1 (5,1) #6
wire n4424; //IPIN -1 (5,1) #7
wire n4425; //IPIN -1 (5,1) #8
wire n4426; //IPIN -1 (5,1) #9
wire n4427; //IPIN -1 (5,1) #10
wire n4428; //IPIN -1 (5,1) #11
wire n4429; //IPIN -1 (5,1) #12
wire n4430; //IPIN -1 (5,1) #13
wire n4431; //IPIN -1 (5,1) #14
wire n4432; //IPIN -1 (5,1) #15
wire n4433; //IPIN -1 (5,1) #16
wire n4434; //IPIN -1 (5,1) #17
wire n4435; //IPIN -1 (5,1) #18
wire n4436; //IPIN -1 (5,1) #19
wire n4437; //IPIN -1 (5,1) #20
wire n4438; //IPIN -1 (5,1) #21
wire n4439; //IPIN -1 (5,1) #22
wire n4440; //IPIN -1 (5,1) #23
wire n4441; //IPIN -1 (5,1) #24
wire n4442; //IPIN -1 (5,1) #25
wire n4443; //IPIN -1 (5,1) #26
wire n4444; //IPIN -1 (5,1) #27
wire n4445; //IPIN -1 (5,1) #28
wire n4446; //IPIN -1 (5,1) #29
wire n4447; //IPIN -1 (5,1) #30
wire n4448; //IPIN -1 (5,1) #31
wire n4449; //IPIN -1 (5,1) #32
wire n4450; //IPIN -1 (5,1) #33
wire n4451; //IPIN -1 (5,1) #34
wire n4452; //IPIN -1 (5,1) #35
wire n4453; //IPIN -1 (5,1) #36
wire n4454; //IPIN -1 (5,1) #37
wire n4455; //IPIN -1 (5,1) #38
wire n4456; //IPIN -1 (5,1) #39
wire n4457; //IPIN -1 (5,1) #40
wire n4458; //IPIN -1 (5,1) #41
wire n4459; //IPIN -1 (5,1) #42
wire n4460; //IPIN -1 (5,1) #43
wire n4461; //IPIN -1 (5,1) #44
wire n4462; //IPIN -1 (5,1) #45
wire n4463; //IPIN -1 (5,1) #46
wire n4464; //IPIN -1 (5,1) #47
wire n4465; //IPIN -1 (5,1) #48
wire n4466; //IPIN -1 (5,1) #49
wire n4467; //IPIN -1 (5,1) #50
wire n4468; //IPIN -1 (5,1) #51
wire n4469; //OPIN -1 (5,1) #52
wire n4470; //OPIN -1 (5,1) #53
wire n4471; //OPIN -1 (5,1) #54
wire n4472; //OPIN -1 (5,1) #55
wire n4473; //OPIN -1 (5,1) #56
wire n4474; //OPIN -1 (5,1) #57
wire n4475; //OPIN -1 (5,1) #58
wire n4476; //OPIN -1 (5,1) #59
wire n4477; //OPIN -1 (5,1) #60
wire n4478; //OPIN -1 (5,1) #61
wire n4479; //OPIN -1 (5,1) #62
wire n4480; //OPIN -1 (5,1) #63
wire n4481; //OPIN -1 (5,1) #64
wire n4482; //OPIN -1 (5,1) #65
wire n4483; //OPIN -1 (5,1) #66
wire n4484; //OPIN -1 (5,1) #67
wire n4485; //OPIN -1 (5,1) #68
wire n4486; //OPIN -1 (5,1) #69
wire n4487; //OPIN -1 (5,1) #70
wire n4488; //OPIN -1 (5,1) #71
wire n4489; //IPIN -1 (5,1) #72
wire n4515; //IPIN -1 (5,2) #0
wire n4516; //IPIN -1 (5,2) #1
wire n4517; //IPIN -1 (5,2) #2
wire n4518; //IPIN -1 (5,2) #3
wire n4519; //IPIN -1 (5,2) #4
wire n4520; //IPIN -1 (5,2) #5
wire n4521; //IPIN -1 (5,2) #6
wire n4522; //IPIN -1 (5,2) #7
wire n4523; //IPIN -1 (5,2) #8
wire n4524; //IPIN -1 (5,2) #9
wire n4525; //IPIN -1 (5,2) #10
wire n4526; //IPIN -1 (5,2) #11
wire n4527; //IPIN -1 (5,2) #12
wire n4528; //IPIN -1 (5,2) #13
wire n4529; //IPIN -1 (5,2) #14
wire n4530; //IPIN -1 (5,2) #15
wire n4531; //IPIN -1 (5,2) #16
wire n4532; //IPIN -1 (5,2) #17
wire n4533; //IPIN -1 (5,2) #18
wire n4534; //IPIN -1 (5,2) #19
wire n4535; //IPIN -1 (5,2) #20
wire n4536; //IPIN -1 (5,2) #21
wire n4537; //IPIN -1 (5,2) #22
wire n4538; //IPIN -1 (5,2) #23
wire n4539; //IPIN -1 (5,2) #24
wire n4540; //IPIN -1 (5,2) #25
wire n4541; //IPIN -1 (5,2) #26
wire n4542; //IPIN -1 (5,2) #27
wire n4543; //IPIN -1 (5,2) #28
wire n4544; //IPIN -1 (5,2) #29
wire n4545; //IPIN -1 (5,2) #30
wire n4546; //IPIN -1 (5,2) #31
wire n4547; //IPIN -1 (5,2) #32
wire n4548; //IPIN -1 (5,2) #33
wire n4549; //IPIN -1 (5,2) #34
wire n4550; //IPIN -1 (5,2) #35
wire n4551; //IPIN -1 (5,2) #36
wire n4552; //IPIN -1 (5,2) #37
wire n4553; //IPIN -1 (5,2) #38
wire n4554; //IPIN -1 (5,2) #39
wire n4555; //IPIN -1 (5,2) #40
wire n4556; //IPIN -1 (5,2) #41
wire n4557; //IPIN -1 (5,2) #42
wire n4558; //IPIN -1 (5,2) #43
wire n4559; //IPIN -1 (5,2) #44
wire n4560; //IPIN -1 (5,2) #45
wire n4561; //IPIN -1 (5,2) #46
wire n4562; //IPIN -1 (5,2) #47
wire n4563; //IPIN -1 (5,2) #48
wire n4564; //IPIN -1 (5,2) #49
wire n4565; //IPIN -1 (5,2) #50
wire n4566; //IPIN -1 (5,2) #51
wire n4567; //OPIN -1 (5,2) #52
wire n4568; //OPIN -1 (5,2) #53
wire n4569; //OPIN -1 (5,2) #54
wire n4570; //OPIN -1 (5,2) #55
wire n4571; //OPIN -1 (5,2) #56
wire n4572; //OPIN -1 (5,2) #57
wire n4573; //OPIN -1 (5,2) #58
wire n4574; //OPIN -1 (5,2) #59
wire n4575; //OPIN -1 (5,2) #60
wire n4576; //OPIN -1 (5,2) #61
wire n4577; //OPIN -1 (5,2) #62
wire n4578; //OPIN -1 (5,2) #63
wire n4579; //OPIN -1 (5,2) #64
wire n4580; //OPIN -1 (5,2) #65
wire n4581; //OPIN -1 (5,2) #66
wire n4582; //OPIN -1 (5,2) #67
wire n4583; //OPIN -1 (5,2) #68
wire n4584; //OPIN -1 (5,2) #69
wire n4585; //OPIN -1 (5,2) #70
wire n4586; //OPIN -1 (5,2) #71
wire n4587; //IPIN -1 (5,2) #72
wire n4613; //IPIN -1 (5,3) #0
wire n4614; //IPIN -1 (5,3) #1
wire n4615; //IPIN -1 (5,3) #2
wire n4616; //IPIN -1 (5,3) #3
wire n4617; //IPIN -1 (5,3) #4
wire n4618; //IPIN -1 (5,3) #5
wire n4619; //IPIN -1 (5,3) #6
wire n4620; //IPIN -1 (5,3) #7
wire n4621; //IPIN -1 (5,3) #8
wire n4622; //IPIN -1 (5,3) #9
wire n4623; //IPIN -1 (5,3) #10
wire n4624; //IPIN -1 (5,3) #11
wire n4625; //IPIN -1 (5,3) #12
wire n4626; //IPIN -1 (5,3) #13
wire n4627; //IPIN -1 (5,3) #14
wire n4628; //IPIN -1 (5,3) #15
wire n4629; //IPIN -1 (5,3) #16
wire n4630; //IPIN -1 (5,3) #17
wire n4631; //IPIN -1 (5,3) #18
wire n4632; //IPIN -1 (5,3) #19
wire n4633; //IPIN -1 (5,3) #20
wire n4634; //IPIN -1 (5,3) #21
wire n4635; //IPIN -1 (5,3) #22
wire n4636; //IPIN -1 (5,3) #23
wire n4637; //IPIN -1 (5,3) #24
wire n4638; //IPIN -1 (5,3) #25
wire n4639; //IPIN -1 (5,3) #26
wire n4640; //IPIN -1 (5,3) #27
wire n4641; //IPIN -1 (5,3) #28
wire n4642; //IPIN -1 (5,3) #29
wire n4643; //IPIN -1 (5,3) #30
wire n4644; //IPIN -1 (5,3) #31
wire n4645; //IPIN -1 (5,3) #32
wire n4646; //IPIN -1 (5,3) #33
wire n4647; //IPIN -1 (5,3) #34
wire n4648; //IPIN -1 (5,3) #35
wire n4649; //IPIN -1 (5,3) #36
wire n4650; //IPIN -1 (5,3) #37
wire n4651; //IPIN -1 (5,3) #38
wire n4652; //IPIN -1 (5,3) #39
wire n4653; //IPIN -1 (5,3) #40
wire n4654; //IPIN -1 (5,3) #41
wire n4655; //IPIN -1 (5,3) #42
wire n4656; //IPIN -1 (5,3) #43
wire n4657; //IPIN -1 (5,3) #44
wire n4658; //IPIN -1 (5,3) #45
wire n4659; //IPIN -1 (5,3) #46
wire n4660; //IPIN -1 (5,3) #47
wire n4661; //IPIN -1 (5,3) #48
wire n4662; //IPIN -1 (5,3) #49
wire n4663; //IPIN -1 (5,3) #50
wire n4664; //IPIN -1 (5,3) #51
wire n4665; //OPIN -1 (5,3) #52
wire n4666; //OPIN -1 (5,3) #53
wire n4667; //OPIN -1 (5,3) #54
wire n4668; //OPIN -1 (5,3) #55
wire n4669; //OPIN -1 (5,3) #56
wire n4670; //OPIN -1 (5,3) #57
wire n4671; //OPIN -1 (5,3) #58
wire n4672; //OPIN -1 (5,3) #59
wire n4673; //OPIN -1 (5,3) #60
wire n4674; //OPIN -1 (5,3) #61
wire n4675; //OPIN -1 (5,3) #62
wire n4676; //OPIN -1 (5,3) #63
wire n4677; //OPIN -1 (5,3) #64
wire n4678; //OPIN -1 (5,3) #65
wire n4679; //OPIN -1 (5,3) #66
wire n4680; //OPIN -1 (5,3) #67
wire n4681; //OPIN -1 (5,3) #68
wire n4682; //OPIN -1 (5,3) #69
wire n4683; //OPIN -1 (5,3) #70
wire n4684; //OPIN -1 (5,3) #71
wire n4685; //IPIN -1 (5,3) #72
wire n4711; //IPIN -1 (5,4) #0
wire n4712; //IPIN -1 (5,4) #1
wire n4713; //IPIN -1 (5,4) #2
wire n4714; //IPIN -1 (5,4) #3
wire n4715; //IPIN -1 (5,4) #4
wire n4716; //IPIN -1 (5,4) #5
wire n4717; //IPIN -1 (5,4) #6
wire n4718; //IPIN -1 (5,4) #7
wire n4719; //IPIN -1 (5,4) #8
wire n4720; //IPIN -1 (5,4) #9
wire n4721; //IPIN -1 (5,4) #10
wire n4722; //IPIN -1 (5,4) #11
wire n4723; //IPIN -1 (5,4) #12
wire n4724; //IPIN -1 (5,4) #13
wire n4725; //IPIN -1 (5,4) #14
wire n4726; //IPIN -1 (5,4) #15
wire n4727; //IPIN -1 (5,4) #16
wire n4728; //IPIN -1 (5,4) #17
wire n4729; //IPIN -1 (5,4) #18
wire n4730; //IPIN -1 (5,4) #19
wire n4731; //IPIN -1 (5,4) #20
wire n4732; //IPIN -1 (5,4) #21
wire n4733; //IPIN -1 (5,4) #22
wire n4734; //IPIN -1 (5,4) #23
wire n4735; //IPIN -1 (5,4) #24
wire n4736; //IPIN -1 (5,4) #25
wire n4737; //IPIN -1 (5,4) #26
wire n4738; //IPIN -1 (5,4) #27
wire n4739; //IPIN -1 (5,4) #28
wire n4740; //IPIN -1 (5,4) #29
wire n4741; //IPIN -1 (5,4) #30
wire n4742; //IPIN -1 (5,4) #31
wire n4743; //IPIN -1 (5,4) #32
wire n4744; //IPIN -1 (5,4) #33
wire n4745; //IPIN -1 (5,4) #34
wire n4746; //IPIN -1 (5,4) #35
wire n4747; //IPIN -1 (5,4) #36
wire n4748; //IPIN -1 (5,4) #37
wire n4749; //IPIN -1 (5,4) #38
wire n4750; //IPIN -1 (5,4) #39
wire n4751; //IPIN -1 (5,4) #40
wire n4752; //IPIN -1 (5,4) #41
wire n4753; //IPIN -1 (5,4) #42
wire n4754; //IPIN -1 (5,4) #43
wire n4755; //IPIN -1 (5,4) #44
wire n4756; //IPIN -1 (5,4) #45
wire n4757; //IPIN -1 (5,4) #46
wire n4758; //IPIN -1 (5,4) #47
wire n4759; //IPIN -1 (5,4) #48
wire n4760; //IPIN -1 (5,4) #49
wire n4761; //IPIN -1 (5,4) #50
wire n4762; //IPIN -1 (5,4) #51
wire n4763; //OPIN -1 (5,4) #52
wire n4764; //OPIN -1 (5,4) #53
wire n4765; //OPIN -1 (5,4) #54
wire n4766; //OPIN -1 (5,4) #55
wire n4767; //OPIN -1 (5,4) #56
wire n4768; //OPIN -1 (5,4) #57
wire n4769; //OPIN -1 (5,4) #58
wire n4770; //OPIN -1 (5,4) #59
wire n4771; //OPIN -1 (5,4) #60
wire n4772; //OPIN -1 (5,4) #61
wire n4773; //OPIN -1 (5,4) #62
wire n4774; //OPIN -1 (5,4) #63
wire n4775; //OPIN -1 (5,4) #64
wire n4776; //OPIN -1 (5,4) #65
wire n4777; //OPIN -1 (5,4) #66
wire n4778; //OPIN -1 (5,4) #67
wire n4779; //OPIN -1 (5,4) #68
wire n4780; //OPIN -1 (5,4) #69
wire n4781; //OPIN -1 (5,4) #70
wire n4782; //OPIN -1 (5,4) #71
wire n4783; //IPIN -1 (5,4) #72
wire n4809; //IPIN -1 (5,5) #0
wire n4810; //IPIN -1 (5,5) #1
wire n4811; //IPIN -1 (5,5) #2
wire n4812; //IPIN -1 (5,5) #3
wire n4813; //IPIN -1 (5,5) #4
wire n4814; //IPIN -1 (5,5) #5
wire n4815; //IPIN -1 (5,5) #6
wire n4816; //IPIN -1 (5,5) #7
wire n4817; //IPIN -1 (5,5) #8
wire n4818; //IPIN -1 (5,5) #9
wire n4819; //IPIN -1 (5,5) #10
wire n4820; //IPIN -1 (5,5) #11
wire n4821; //IPIN -1 (5,5) #12
wire n4822; //IPIN -1 (5,5) #13
wire n4823; //IPIN -1 (5,5) #14
wire n4824; //IPIN -1 (5,5) #15
wire n4825; //IPIN -1 (5,5) #16
wire n4826; //IPIN -1 (5,5) #17
wire n4827; //IPIN -1 (5,5) #18
wire n4828; //IPIN -1 (5,5) #19
wire n4829; //IPIN -1 (5,5) #20
wire n4830; //IPIN -1 (5,5) #21
wire n4831; //IPIN -1 (5,5) #22
wire n4832; //IPIN -1 (5,5) #23
wire n4833; //IPIN -1 (5,5) #24
wire n4834; //IPIN -1 (5,5) #25
wire n4835; //IPIN -1 (5,5) #26
wire n4836; //IPIN -1 (5,5) #27
wire n4837; //IPIN -1 (5,5) #28
wire n4838; //IPIN -1 (5,5) #29
wire n4839; //IPIN -1 (5,5) #30
wire n4840; //IPIN -1 (5,5) #31
wire n4841; //IPIN -1 (5,5) #32
wire n4842; //IPIN -1 (5,5) #33
wire n4843; //IPIN -1 (5,5) #34
wire n4844; //IPIN -1 (5,5) #35
wire n4845; //IPIN -1 (5,5) #36
wire n4846; //IPIN -1 (5,5) #37
wire n4847; //IPIN -1 (5,5) #38
wire n4848; //IPIN -1 (5,5) #39
wire n4849; //IPIN -1 (5,5) #40
wire n4850; //IPIN -1 (5,5) #41
wire n4851; //IPIN -1 (5,5) #42
wire n4852; //IPIN -1 (5,5) #43
wire n4853; //IPIN -1 (5,5) #44
wire n4854; //IPIN -1 (5,5) #45
wire n4855; //IPIN -1 (5,5) #46
wire n4856; //IPIN -1 (5,5) #47
wire n4857; //IPIN -1 (5,5) #48
wire n4858; //IPIN -1 (5,5) #49
wire n4859; //IPIN -1 (5,5) #50
wire n4860; //IPIN -1 (5,5) #51
wire n4861; //OPIN -1 (5,5) #52
wire n4862; //OPIN -1 (5,5) #53
wire n4863; //OPIN -1 (5,5) #54
wire n4864; //OPIN -1 (5,5) #55
wire n4865; //OPIN -1 (5,5) #56
wire n4866; //OPIN -1 (5,5) #57
wire n4867; //OPIN -1 (5,5) #58
wire n4868; //OPIN -1 (5,5) #59
wire n4869; //OPIN -1 (5,5) #60
wire n4870; //OPIN -1 (5,5) #61
wire n4871; //OPIN -1 (5,5) #62
wire n4872; //OPIN -1 (5,5) #63
wire n4873; //OPIN -1 (5,5) #64
wire n4874; //OPIN -1 (5,5) #65
wire n4875; //OPIN -1 (5,5) #66
wire n4876; //OPIN -1 (5,5) #67
wire n4877; //OPIN -1 (5,5) #68
wire n4878; //OPIN -1 (5,5) #69
wire n4879; //OPIN -1 (5,5) #70
wire n4880; //OPIN -1 (5,5) #71
wire n4881; //IPIN -1 (5,5) #72
wire n4907; //IPIN -1 (5,6) #0
wire n4908; //IPIN -1 (5,6) #1
wire n4909; //IPIN -1 (5,6) #2
wire n4910; //IPIN -1 (5,6) #3
wire n4911; //IPIN -1 (5,6) #4
wire n4912; //IPIN -1 (5,6) #5
wire n4913; //IPIN -1 (5,6) #6
wire n4914; //IPIN -1 (5,6) #7
wire n4915; //IPIN -1 (5,6) #8
wire n4916; //IPIN -1 (5,6) #9
wire n4917; //IPIN -1 (5,6) #10
wire n4918; //IPIN -1 (5,6) #11
wire n4919; //IPIN -1 (5,6) #12
wire n4920; //IPIN -1 (5,6) #13
wire n4921; //IPIN -1 (5,6) #14
wire n4922; //IPIN -1 (5,6) #15
wire n4923; //IPIN -1 (5,6) #16
wire n4924; //IPIN -1 (5,6) #17
wire n4925; //IPIN -1 (5,6) #18
wire n4926; //IPIN -1 (5,6) #19
wire n4927; //IPIN -1 (5,6) #20
wire n4928; //IPIN -1 (5,6) #21
wire n4929; //IPIN -1 (5,6) #22
wire n4930; //IPIN -1 (5,6) #23
wire n4931; //IPIN -1 (5,6) #24
wire n4932; //IPIN -1 (5,6) #25
wire n4933; //IPIN -1 (5,6) #26
wire n4934; //IPIN -1 (5,6) #27
wire n4935; //IPIN -1 (5,6) #28
wire n4936; //IPIN -1 (5,6) #29
wire n4937; //IPIN -1 (5,6) #30
wire n4938; //IPIN -1 (5,6) #31
wire n4939; //IPIN -1 (5,6) #32
wire n4940; //IPIN -1 (5,6) #33
wire n4941; //IPIN -1 (5,6) #34
wire n4942; //IPIN -1 (5,6) #35
wire n4943; //IPIN -1 (5,6) #36
wire n4944; //IPIN -1 (5,6) #37
wire n4945; //IPIN -1 (5,6) #38
wire n4946; //IPIN -1 (5,6) #39
wire n4947; //IPIN -1 (5,6) #40
wire n4948; //IPIN -1 (5,6) #41
wire n4949; //IPIN -1 (5,6) #42
wire n4950; //IPIN -1 (5,6) #43
wire n4951; //IPIN -1 (5,6) #44
wire n4952; //IPIN -1 (5,6) #45
wire n4953; //IPIN -1 (5,6) #46
wire n4954; //IPIN -1 (5,6) #47
wire n4955; //IPIN -1 (5,6) #48
wire n4956; //IPIN -1 (5,6) #49
wire n4957; //IPIN -1 (5,6) #50
wire n4958; //IPIN -1 (5,6) #51
wire n4959; //OPIN -1 (5,6) #52
wire n4960; //OPIN -1 (5,6) #53
wire n4961; //OPIN -1 (5,6) #54
wire n4962; //OPIN -1 (5,6) #55
wire n4963; //OPIN -1 (5,6) #56
wire n4964; //OPIN -1 (5,6) #57
wire n4965; //OPIN -1 (5,6) #58
wire n4966; //OPIN -1 (5,6) #59
wire n4967; //OPIN -1 (5,6) #60
wire n4968; //OPIN -1 (5,6) #61
wire n4969; //OPIN -1 (5,6) #62
wire n4970; //OPIN -1 (5,6) #63
wire n4971; //OPIN -1 (5,6) #64
wire n4972; //OPIN -1 (5,6) #65
wire n4973; //OPIN -1 (5,6) #66
wire n4974; //OPIN -1 (5,6) #67
wire n4975; //OPIN -1 (5,6) #68
wire n4976; //OPIN -1 (5,6) #69
wire n4977; //OPIN -1 (5,6) #70
wire n4978; //OPIN -1 (5,6) #71
wire n4979; //IPIN -1 (5,6) #72
wire n5005; //IPIN -1 (5,7) #0
wire n5006; //IPIN -1 (5,7) #1
wire n5007; //IPIN -1 (5,7) #2
wire n5008; //IPIN -1 (5,7) #3
wire n5009; //IPIN -1 (5,7) #4
wire n5010; //IPIN -1 (5,7) #5
wire n5011; //IPIN -1 (5,7) #6
wire n5012; //IPIN -1 (5,7) #7
wire n5013; //IPIN -1 (5,7) #8
wire n5014; //IPIN -1 (5,7) #9
wire n5015; //IPIN -1 (5,7) #10
wire n5016; //IPIN -1 (5,7) #11
wire n5017; //IPIN -1 (5,7) #12
wire n5018; //IPIN -1 (5,7) #13
wire n5019; //IPIN -1 (5,7) #14
wire n5020; //IPIN -1 (5,7) #15
wire n5021; //IPIN -1 (5,7) #16
wire n5022; //IPIN -1 (5,7) #17
wire n5023; //IPIN -1 (5,7) #18
wire n5024; //IPIN -1 (5,7) #19
wire n5025; //IPIN -1 (5,7) #20
wire n5026; //IPIN -1 (5,7) #21
wire n5027; //IPIN -1 (5,7) #22
wire n5028; //IPIN -1 (5,7) #23
wire n5029; //IPIN -1 (5,7) #24
wire n5030; //IPIN -1 (5,7) #25
wire n5031; //IPIN -1 (5,7) #26
wire n5032; //IPIN -1 (5,7) #27
wire n5033; //IPIN -1 (5,7) #28
wire n5034; //IPIN -1 (5,7) #29
wire n5035; //IPIN -1 (5,7) #30
wire n5036; //IPIN -1 (5,7) #31
wire n5037; //IPIN -1 (5,7) #32
wire n5038; //IPIN -1 (5,7) #33
wire n5039; //IPIN -1 (5,7) #34
wire n5040; //IPIN -1 (5,7) #35
wire n5041; //IPIN -1 (5,7) #36
wire n5042; //IPIN -1 (5,7) #37
wire n5043; //IPIN -1 (5,7) #38
wire n5044; //IPIN -1 (5,7) #39
wire n5045; //IPIN -1 (5,7) #40
wire n5046; //IPIN -1 (5,7) #41
wire n5047; //IPIN -1 (5,7) #42
wire n5048; //IPIN -1 (5,7) #43
wire n5049; //IPIN -1 (5,7) #44
wire n5050; //IPIN -1 (5,7) #45
wire n5051; //IPIN -1 (5,7) #46
wire n5052; //IPIN -1 (5,7) #47
wire n5053; //IPIN -1 (5,7) #48
wire n5054; //IPIN -1 (5,7) #49
wire n5055; //IPIN -1 (5,7) #50
wire n5056; //IPIN -1 (5,7) #51
wire n5057; //OPIN -1 (5,7) #52
wire n5058; //OPIN -1 (5,7) #53
wire n5059; //OPIN -1 (5,7) #54
wire n5060; //OPIN -1 (5,7) #55
wire n5061; //OPIN -1 (5,7) #56
wire n5062; //OPIN -1 (5,7) #57
wire n5063; //OPIN -1 (5,7) #58
wire n5064; //OPIN -1 (5,7) #59
wire n5065; //OPIN -1 (5,7) #60
wire n5066; //OPIN -1 (5,7) #61
wire n5067; //OPIN -1 (5,7) #62
wire n5068; //OPIN -1 (5,7) #63
wire n5069; //OPIN -1 (5,7) #64
wire n5070; //OPIN -1 (5,7) #65
wire n5071; //OPIN -1 (5,7) #66
wire n5072; //OPIN -1 (5,7) #67
wire n5073; //OPIN -1 (5,7) #68
wire n5074; //OPIN -1 (5,7) #69
wire n5075; //OPIN -1 (5,7) #70
wire n5076; //OPIN -1 (5,7) #71
wire n5077; //IPIN -1 (5,7) #72
wire n5103; //IPIN -1 (5,8) #0
wire n5104; //IPIN -1 (5,8) #1
wire n5105; //IPIN -1 (5,8) #2
wire n5106; //IPIN -1 (5,8) #3
wire n5107; //IPIN -1 (5,8) #4
wire n5108; //IPIN -1 (5,8) #5
wire n5109; //IPIN -1 (5,8) #6
wire n5110; //IPIN -1 (5,8) #7
wire n5111; //IPIN -1 (5,8) #8
wire n5112; //IPIN -1 (5,8) #9
wire n5113; //IPIN -1 (5,8) #10
wire n5114; //IPIN -1 (5,8) #11
wire n5115; //IPIN -1 (5,8) #12
wire n5116; //IPIN -1 (5,8) #13
wire n5117; //IPIN -1 (5,8) #14
wire n5118; //IPIN -1 (5,8) #15
wire n5119; //IPIN -1 (5,8) #16
wire n5120; //IPIN -1 (5,8) #17
wire n5121; //IPIN -1 (5,8) #18
wire n5122; //IPIN -1 (5,8) #19
wire n5123; //IPIN -1 (5,8) #20
wire n5124; //IPIN -1 (5,8) #21
wire n5125; //IPIN -1 (5,8) #22
wire n5126; //IPIN -1 (5,8) #23
wire n5127; //IPIN -1 (5,8) #24
wire n5128; //IPIN -1 (5,8) #25
wire n5129; //IPIN -1 (5,8) #26
wire n5130; //IPIN -1 (5,8) #27
wire n5131; //IPIN -1 (5,8) #28
wire n5132; //IPIN -1 (5,8) #29
wire n5133; //IPIN -1 (5,8) #30
wire n5134; //IPIN -1 (5,8) #31
wire n5135; //IPIN -1 (5,8) #32
wire n5136; //IPIN -1 (5,8) #33
wire n5137; //IPIN -1 (5,8) #34
wire n5138; //IPIN -1 (5,8) #35
wire n5139; //IPIN -1 (5,8) #36
wire n5140; //IPIN -1 (5,8) #37
wire n5141; //IPIN -1 (5,8) #38
wire n5142; //IPIN -1 (5,8) #39
wire n5143; //IPIN -1 (5,8) #40
wire n5144; //IPIN -1 (5,8) #41
wire n5145; //IPIN -1 (5,8) #42
wire n5146; //IPIN -1 (5,8) #43
wire n5147; //IPIN -1 (5,8) #44
wire n5148; //IPIN -1 (5,8) #45
wire n5149; //IPIN -1 (5,8) #46
wire n5150; //IPIN -1 (5,8) #47
wire n5151; //IPIN -1 (5,8) #48
wire n5152; //IPIN -1 (5,8) #49
wire n5153; //IPIN -1 (5,8) #50
wire n5154; //IPIN -1 (5,8) #51
wire n5155; //OPIN -1 (5,8) #52
wire n5156; //OPIN -1 (5,8) #53
wire n5157; //OPIN -1 (5,8) #54
wire n5158; //OPIN -1 (5,8) #55
wire n5159; //OPIN -1 (5,8) #56
wire n5160; //OPIN -1 (5,8) #57
wire n5161; //OPIN -1 (5,8) #58
wire n5162; //OPIN -1 (5,8) #59
wire n5163; //OPIN -1 (5,8) #60
wire n5164; //OPIN -1 (5,8) #61
wire n5165; //OPIN -1 (5,8) #62
wire n5166; //OPIN -1 (5,8) #63
wire n5167; //OPIN -1 (5,8) #64
wire n5168; //OPIN -1 (5,8) #65
wire n5169; //OPIN -1 (5,8) #66
wire n5170; //OPIN -1 (5,8) #67
wire n5171; //OPIN -1 (5,8) #68
wire n5172; //OPIN -1 (5,8) #69
wire n5173; //OPIN -1 (5,8) #70
wire n5174; //OPIN -1 (5,8) #71
wire n5175; //IPIN -1 (5,8) #72
wire n5201; //IPIN -1 (5,9) #0
wire n5202; //IPIN -1 (5,9) #1
wire n5203; //IPIN -1 (5,9) #2
wire n5204; //IPIN -1 (5,9) #3
wire n5205; //IPIN -1 (5,9) #4
wire n5206; //IPIN -1 (5,9) #5
wire n5207; //IPIN -1 (5,9) #6
wire n5208; //IPIN -1 (5,9) #7
wire n5209; //IPIN -1 (5,9) #8
wire n5210; //IPIN -1 (5,9) #9
wire n5211; //IPIN -1 (5,9) #10
wire n5212; //IPIN -1 (5,9) #11
wire n5213; //IPIN -1 (5,9) #12
wire n5214; //IPIN -1 (5,9) #13
wire n5215; //IPIN -1 (5,9) #14
wire n5216; //IPIN -1 (5,9) #15
wire n5217; //IPIN -1 (5,9) #16
wire n5218; //IPIN -1 (5,9) #17
wire n5219; //IPIN -1 (5,9) #18
wire n5220; //IPIN -1 (5,9) #19
wire n5221; //IPIN -1 (5,9) #20
wire n5222; //IPIN -1 (5,9) #21
wire n5223; //IPIN -1 (5,9) #22
wire n5224; //IPIN -1 (5,9) #23
wire n5225; //IPIN -1 (5,9) #24
wire n5226; //IPIN -1 (5,9) #25
wire n5227; //IPIN -1 (5,9) #26
wire n5228; //IPIN -1 (5,9) #27
wire n5229; //IPIN -1 (5,9) #28
wire n5230; //IPIN -1 (5,9) #29
wire n5231; //IPIN -1 (5,9) #30
wire n5232; //IPIN -1 (5,9) #31
wire n5233; //IPIN -1 (5,9) #32
wire n5234; //IPIN -1 (5,9) #33
wire n5235; //IPIN -1 (5,9) #34
wire n5236; //IPIN -1 (5,9) #35
wire n5237; //IPIN -1 (5,9) #36
wire n5238; //IPIN -1 (5,9) #37
wire n5239; //IPIN -1 (5,9) #38
wire n5240; //IPIN -1 (5,9) #39
wire n5241; //IPIN -1 (5,9) #40
wire n5242; //IPIN -1 (5,9) #41
wire n5243; //IPIN -1 (5,9) #42
wire n5244; //IPIN -1 (5,9) #43
wire n5245; //IPIN -1 (5,9) #44
wire n5246; //IPIN -1 (5,9) #45
wire n5247; //IPIN -1 (5,9) #46
wire n5248; //IPIN -1 (5,9) #47
wire n5249; //IPIN -1 (5,9) #48
wire n5250; //IPIN -1 (5,9) #49
wire n5251; //IPIN -1 (5,9) #50
wire n5252; //IPIN -1 (5,9) #51
wire n5253; //OPIN -1 (5,9) #52
wire n5254; //OPIN -1 (5,9) #53
wire n5255; //OPIN -1 (5,9) #54
wire n5256; //OPIN -1 (5,9) #55
wire n5257; //OPIN -1 (5,9) #56
wire n5258; //OPIN -1 (5,9) #57
wire n5259; //OPIN -1 (5,9) #58
wire n5260; //OPIN -1 (5,9) #59
wire n5261; //OPIN -1 (5,9) #60
wire n5262; //OPIN -1 (5,9) #61
wire n5263; //OPIN -1 (5,9) #62
wire n5264; //OPIN -1 (5,9) #63
wire n5265; //OPIN -1 (5,9) #64
wire n5266; //OPIN -1 (5,9) #65
wire n5267; //OPIN -1 (5,9) #66
wire n5268; //OPIN -1 (5,9) #67
wire n5269; //OPIN -1 (5,9) #68
wire n5270; //OPIN -1 (5,9) #69
wire n5271; //OPIN -1 (5,9) #70
wire n5272; //OPIN -1 (5,9) #71
wire n5273; //IPIN -1 (5,9) #72
wire n5298; //IPIN -1 (5,10) #0
wire n5299; //OPIN -1 (5,10) #1
wire n5300; //IPIN -1 (5,10) #2
wire n5301; //IPIN -1 (5,10) #3
wire n5302; //OPIN -1 (5,10) #4
wire n5303; //IPIN -1 (5,10) #5
wire n5304; //IPIN -1 (5,10) #6
wire n5305; //OPIN -1 (5,10) #7
wire n5306; //IPIN -1 (5,10) #8
wire n5307; //IPIN -1 (5,10) #9
wire n5308; //OPIN -1 (5,10) #10
wire n5309; //IPIN -1 (5,10) #11
wire n5310; //IPIN -1 (5,10) #12
wire n5311; //OPIN -1 (5,10) #13
wire n5312; //IPIN -1 (5,10) #14
wire n5313; //IPIN -1 (5,10) #15
wire n5314; //OPIN -1 (5,10) #16
wire n5315; //IPIN -1 (5,10) #17
wire n5316; //IPIN -1 (5,10) #18
wire n5317; //OPIN -1 (5,10) #19
wire n5318; //IPIN -1 (5,10) #20
wire n5319; //IPIN -1 (5,10) #21
wire n5320; //OPIN -1 (5,10) #22
wire n5321; //IPIN -1 (5,10) #23
wire n5346; //IPIN -1 (6,0) #0
wire n5347; //OPIN -1 (6,0) #1
wire n5348; //IPIN -1 (6,0) #2
wire n5349; //IPIN -1 (6,0) #3
wire n5350; //OPIN -1 (6,0) #4
wire n5351; //IPIN -1 (6,0) #5
wire n5352; //IPIN -1 (6,0) #6
wire n5353; //OPIN -1 (6,0) #7
wire n5354; //IPIN -1 (6,0) #8
wire n5355; //IPIN -1 (6,0) #9
wire n5356; //OPIN -1 (6,0) #10
wire n5357; //IPIN -1 (6,0) #11
wire n5358; //IPIN -1 (6,0) #12
wire n5359; //OPIN -1 (6,0) #13
wire n5360; //IPIN -1 (6,0) #14
wire n5361; //IPIN -1 (6,0) #15
wire n5362; //OPIN -1 (6,0) #16
wire n5363; //IPIN -1 (6,0) #17
wire n5364; //IPIN -1 (6,0) #18
wire n5365; //OPIN -1 (6,0) #19
wire n5366; //IPIN -1 (6,0) #20
wire n5367; //IPIN -1 (6,0) #21
wire n5368; //OPIN -1 (6,0) #22
wire n5369; //IPIN -1 (6,0) #23
wire n5395; //IPIN -1 (6,1) #0
wire n5396; //IPIN -1 (6,1) #1
wire n5397; //IPIN -1 (6,1) #2
wire n5398; //IPIN -1 (6,1) #3
wire n5399; //IPIN -1 (6,1) #4
wire n5400; //IPIN -1 (6,1) #5
wire n5401; //IPIN -1 (6,1) #6
wire n5402; //IPIN -1 (6,1) #7
wire n5403; //IPIN -1 (6,1) #8
wire n5404; //IPIN -1 (6,1) #9
wire n5405; //IPIN -1 (6,1) #10
wire n5406; //IPIN -1 (6,1) #11
wire n5407; //IPIN -1 (6,1) #12
wire n5408; //IPIN -1 (6,1) #13
wire n5409; //IPIN -1 (6,1) #14
wire n5410; //IPIN -1 (6,1) #15
wire n5411; //IPIN -1 (6,1) #16
wire n5412; //IPIN -1 (6,1) #17
wire n5413; //IPIN -1 (6,1) #18
wire n5414; //IPIN -1 (6,1) #19
wire n5415; //IPIN -1 (6,1) #20
wire n5416; //IPIN -1 (6,1) #21
wire n5417; //IPIN -1 (6,1) #22
wire n5418; //IPIN -1 (6,1) #23
wire n5419; //IPIN -1 (6,1) #24
wire n5420; //IPIN -1 (6,1) #25
wire n5421; //IPIN -1 (6,1) #26
wire n5422; //IPIN -1 (6,1) #27
wire n5423; //IPIN -1 (6,1) #28
wire n5424; //IPIN -1 (6,1) #29
wire n5425; //IPIN -1 (6,1) #30
wire n5426; //IPIN -1 (6,1) #31
wire n5427; //IPIN -1 (6,1) #32
wire n5428; //IPIN -1 (6,1) #33
wire n5429; //IPIN -1 (6,1) #34
wire n5430; //IPIN -1 (6,1) #35
wire n5431; //IPIN -1 (6,1) #36
wire n5432; //IPIN -1 (6,1) #37
wire n5433; //IPIN -1 (6,1) #38
wire n5434; //IPIN -1 (6,1) #39
wire n5435; //IPIN -1 (6,1) #40
wire n5436; //IPIN -1 (6,1) #41
wire n5437; //IPIN -1 (6,1) #42
wire n5438; //IPIN -1 (6,1) #43
wire n5439; //IPIN -1 (6,1) #44
wire n5440; //IPIN -1 (6,1) #45
wire n5441; //IPIN -1 (6,1) #46
wire n5442; //IPIN -1 (6,1) #47
wire n5443; //IPIN -1 (6,1) #48
wire n5444; //IPIN -1 (6,1) #49
wire n5445; //IPIN -1 (6,1) #50
wire n5446; //IPIN -1 (6,1) #51
wire n5447; //OPIN -1 (6,1) #52
wire n5448; //OPIN -1 (6,1) #53
wire n5449; //OPIN -1 (6,1) #54
wire n5450; //OPIN -1 (6,1) #55
wire n5451; //OPIN -1 (6,1) #56
wire n5452; //OPIN -1 (6,1) #57
wire n5453; //OPIN -1 (6,1) #58
wire n5454; //OPIN -1 (6,1) #59
wire n5455; //OPIN -1 (6,1) #60
wire n5456; //OPIN -1 (6,1) #61
wire n5457; //OPIN -1 (6,1) #62
wire n5458; //OPIN -1 (6,1) #63
wire n5459; //OPIN -1 (6,1) #64
wire n5460; //OPIN -1 (6,1) #65
wire n5461; //OPIN -1 (6,1) #66
wire n5462; //OPIN -1 (6,1) #67
wire n5463; //OPIN -1 (6,1) #68
wire n5464; //OPIN -1 (6,1) #69
wire n5465; //OPIN -1 (6,1) #70
wire n5466; //OPIN -1 (6,1) #71
wire n5467; //IPIN -1 (6,1) #72
wire n5493; //IPIN -1 (6,2) #0
wire n5494; //IPIN -1 (6,2) #1
wire n5495; //IPIN -1 (6,2) #2
wire n5496; //IPIN -1 (6,2) #3
wire n5497; //IPIN -1 (6,2) #4
wire n5498; //IPIN -1 (6,2) #5
wire n5499; //IPIN -1 (6,2) #6
wire n5500; //IPIN -1 (6,2) #7
wire n5501; //IPIN -1 (6,2) #8
wire n5502; //IPIN -1 (6,2) #9
wire n5503; //IPIN -1 (6,2) #10
wire n5504; //IPIN -1 (6,2) #11
wire n5505; //IPIN -1 (6,2) #12
wire n5506; //IPIN -1 (6,2) #13
wire n5507; //IPIN -1 (6,2) #14
wire n5508; //IPIN -1 (6,2) #15
wire n5509; //IPIN -1 (6,2) #16
wire n5510; //IPIN -1 (6,2) #17
wire n5511; //IPIN -1 (6,2) #18
wire n5512; //IPIN -1 (6,2) #19
wire n5513; //IPIN -1 (6,2) #20
wire n5514; //IPIN -1 (6,2) #21
wire n5515; //IPIN -1 (6,2) #22
wire n5516; //IPIN -1 (6,2) #23
wire n5517; //IPIN -1 (6,2) #24
wire n5518; //IPIN -1 (6,2) #25
wire n5519; //IPIN -1 (6,2) #26
wire n5520; //IPIN -1 (6,2) #27
wire n5521; //IPIN -1 (6,2) #28
wire n5522; //IPIN -1 (6,2) #29
wire n5523; //IPIN -1 (6,2) #30
wire n5524; //IPIN -1 (6,2) #31
wire n5525; //IPIN -1 (6,2) #32
wire n5526; //IPIN -1 (6,2) #33
wire n5527; //IPIN -1 (6,2) #34
wire n5528; //IPIN -1 (6,2) #35
wire n5529; //IPIN -1 (6,2) #36
wire n5530; //IPIN -1 (6,2) #37
wire n5531; //IPIN -1 (6,2) #38
wire n5532; //IPIN -1 (6,2) #39
wire n5533; //IPIN -1 (6,2) #40
wire n5534; //IPIN -1 (6,2) #41
wire n5535; //IPIN -1 (6,2) #42
wire n5536; //IPIN -1 (6,2) #43
wire n5537; //IPIN -1 (6,2) #44
wire n5538; //IPIN -1 (6,2) #45
wire n5539; //IPIN -1 (6,2) #46
wire n5540; //IPIN -1 (6,2) #47
wire n5541; //IPIN -1 (6,2) #48
wire n5542; //IPIN -1 (6,2) #49
wire n5543; //IPIN -1 (6,2) #50
wire n5544; //IPIN -1 (6,2) #51
wire n5545; //OPIN -1 (6,2) #52
wire n5546; //OPIN -1 (6,2) #53
wire n5547; //OPIN -1 (6,2) #54
wire n5548; //OPIN -1 (6,2) #55
wire n5549; //OPIN -1 (6,2) #56
wire n5550; //OPIN -1 (6,2) #57
wire n5551; //OPIN -1 (6,2) #58
wire n5552; //OPIN -1 (6,2) #59
wire n5553; //OPIN -1 (6,2) #60
wire n5554; //OPIN -1 (6,2) #61
wire n5555; //OPIN -1 (6,2) #62
wire n5556; //OPIN -1 (6,2) #63
wire n5557; //OPIN -1 (6,2) #64
wire n5558; //OPIN -1 (6,2) #65
wire n5559; //OPIN -1 (6,2) #66
wire n5560; //OPIN -1 (6,2) #67
wire n5561; //OPIN -1 (6,2) #68
wire n5562; //OPIN -1 (6,2) #69
wire n5563; //OPIN -1 (6,2) #70
wire n5564; //OPIN -1 (6,2) #71
wire n5565; //IPIN -1 (6,2) #72
wire n5591; //IPIN -1 (6,3) #0
wire n5592; //IPIN -1 (6,3) #1
wire n5593; //IPIN -1 (6,3) #2
wire n5594; //IPIN -1 (6,3) #3
wire n5595; //IPIN -1 (6,3) #4
wire n5596; //IPIN -1 (6,3) #5
wire n5597; //IPIN -1 (6,3) #6
wire n5598; //IPIN -1 (6,3) #7
wire n5599; //IPIN -1 (6,3) #8
wire n5600; //IPIN -1 (6,3) #9
wire n5601; //IPIN -1 (6,3) #10
wire n5602; //IPIN -1 (6,3) #11
wire n5603; //IPIN -1 (6,3) #12
wire n5604; //IPIN -1 (6,3) #13
wire n5605; //IPIN -1 (6,3) #14
wire n5606; //IPIN -1 (6,3) #15
wire n5607; //IPIN -1 (6,3) #16
wire n5608; //IPIN -1 (6,3) #17
wire n5609; //IPIN -1 (6,3) #18
wire n5610; //IPIN -1 (6,3) #19
wire n5611; //IPIN -1 (6,3) #20
wire n5612; //IPIN -1 (6,3) #21
wire n5613; //IPIN -1 (6,3) #22
wire n5614; //IPIN -1 (6,3) #23
wire n5615; //IPIN -1 (6,3) #24
wire n5616; //IPIN -1 (6,3) #25
wire n5617; //IPIN -1 (6,3) #26
wire n5618; //IPIN -1 (6,3) #27
wire n5619; //IPIN -1 (6,3) #28
wire n5620; //IPIN -1 (6,3) #29
wire n5621; //IPIN -1 (6,3) #30
wire n5622; //IPIN -1 (6,3) #31
wire n5623; //IPIN -1 (6,3) #32
wire n5624; //IPIN -1 (6,3) #33
wire n5625; //IPIN -1 (6,3) #34
wire n5626; //IPIN -1 (6,3) #35
wire n5627; //IPIN -1 (6,3) #36
wire n5628; //IPIN -1 (6,3) #37
wire n5629; //IPIN -1 (6,3) #38
wire n5630; //IPIN -1 (6,3) #39
wire n5631; //IPIN -1 (6,3) #40
wire n5632; //IPIN -1 (6,3) #41
wire n5633; //IPIN -1 (6,3) #42
wire n5634; //IPIN -1 (6,3) #43
wire n5635; //IPIN -1 (6,3) #44
wire n5636; //IPIN -1 (6,3) #45
wire n5637; //IPIN -1 (6,3) #46
wire n5638; //IPIN -1 (6,3) #47
wire n5639; //IPIN -1 (6,3) #48
wire n5640; //IPIN -1 (6,3) #49
wire n5641; //IPIN -1 (6,3) #50
wire n5642; //IPIN -1 (6,3) #51
wire n5643; //OPIN -1 (6,3) #52
wire n5644; //OPIN -1 (6,3) #53
wire n5645; //OPIN -1 (6,3) #54
wire n5646; //OPIN -1 (6,3) #55
wire n5647; //OPIN -1 (6,3) #56
wire n5648; //OPIN -1 (6,3) #57
wire n5649; //OPIN -1 (6,3) #58
wire n5650; //OPIN -1 (6,3) #59
wire n5651; //OPIN -1 (6,3) #60
wire n5652; //OPIN -1 (6,3) #61
wire n5653; //OPIN -1 (6,3) #62
wire n5654; //OPIN -1 (6,3) #63
wire n5655; //OPIN -1 (6,3) #64
wire n5656; //OPIN -1 (6,3) #65
wire n5657; //OPIN -1 (6,3) #66
wire n5658; //OPIN -1 (6,3) #67
wire n5659; //OPIN -1 (6,3) #68
wire n5660; //OPIN -1 (6,3) #69
wire n5661; //OPIN -1 (6,3) #70
wire n5662; //OPIN -1 (6,3) #71
wire n5663; //IPIN -1 (6,3) #72
wire n5689; //IPIN -1 (6,4) #0
wire n5690; //IPIN -1 (6,4) #1
wire n5691; //IPIN -1 (6,4) #2
wire n5692; //IPIN -1 (6,4) #3
wire n5693; //IPIN -1 (6,4) #4
wire n5694; //IPIN -1 (6,4) #5
wire n5695; //IPIN -1 (6,4) #6
wire n5696; //IPIN -1 (6,4) #7
wire n5697; //IPIN -1 (6,4) #8
wire n5698; //IPIN -1 (6,4) #9
wire n5699; //IPIN -1 (6,4) #10
wire n5700; //IPIN -1 (6,4) #11
wire n5701; //IPIN -1 (6,4) #12
wire n5702; //IPIN -1 (6,4) #13
wire n5703; //IPIN -1 (6,4) #14
wire n5704; //IPIN -1 (6,4) #15
wire n5705; //IPIN -1 (6,4) #16
wire n5706; //IPIN -1 (6,4) #17
wire n5707; //IPIN -1 (6,4) #18
wire n5708; //IPIN -1 (6,4) #19
wire n5709; //IPIN -1 (6,4) #20
wire n5710; //IPIN -1 (6,4) #21
wire n5711; //IPIN -1 (6,4) #22
wire n5712; //IPIN -1 (6,4) #23
wire n5713; //IPIN -1 (6,4) #24
wire n5714; //IPIN -1 (6,4) #25
wire n5715; //IPIN -1 (6,4) #26
wire n5716; //IPIN -1 (6,4) #27
wire n5717; //IPIN -1 (6,4) #28
wire n5718; //IPIN -1 (6,4) #29
wire n5719; //IPIN -1 (6,4) #30
wire n5720; //IPIN -1 (6,4) #31
wire n5721; //IPIN -1 (6,4) #32
wire n5722; //IPIN -1 (6,4) #33
wire n5723; //IPIN -1 (6,4) #34
wire n5724; //IPIN -1 (6,4) #35
wire n5725; //IPIN -1 (6,4) #36
wire n5726; //IPIN -1 (6,4) #37
wire n5727; //IPIN -1 (6,4) #38
wire n5728; //IPIN -1 (6,4) #39
wire n5729; //IPIN -1 (6,4) #40
wire n5730; //IPIN -1 (6,4) #41
wire n5731; //IPIN -1 (6,4) #42
wire n5732; //IPIN -1 (6,4) #43
wire n5733; //IPIN -1 (6,4) #44
wire n5734; //IPIN -1 (6,4) #45
wire n5735; //IPIN -1 (6,4) #46
wire n5736; //IPIN -1 (6,4) #47
wire n5737; //IPIN -1 (6,4) #48
wire n5738; //IPIN -1 (6,4) #49
wire n5739; //IPIN -1 (6,4) #50
wire n5740; //IPIN -1 (6,4) #51
wire n5741; //OPIN -1 (6,4) #52
wire n5742; //OPIN -1 (6,4) #53
wire n5743; //OPIN -1 (6,4) #54
wire n5744; //OPIN -1 (6,4) #55
wire n5745; //OPIN -1 (6,4) #56
wire n5746; //OPIN -1 (6,4) #57
wire n5747; //OPIN -1 (6,4) #58
wire n5748; //OPIN -1 (6,4) #59
wire n5749; //OPIN -1 (6,4) #60
wire n5750; //OPIN -1 (6,4) #61
wire n5751; //OPIN -1 (6,4) #62
wire n5752; //OPIN -1 (6,4) #63
wire n5753; //OPIN -1 (6,4) #64
wire n5754; //OPIN -1 (6,4) #65
wire n5755; //OPIN -1 (6,4) #66
wire n5756; //OPIN -1 (6,4) #67
wire n5757; //OPIN -1 (6,4) #68
wire n5758; //OPIN -1 (6,4) #69
wire n5759; //OPIN -1 (6,4) #70
wire n5760; //OPIN -1 (6,4) #71
wire n5761; //IPIN -1 (6,4) #72
wire n5787; //IPIN -1 (6,5) #0
wire n5788; //IPIN -1 (6,5) #1
wire n5789; //IPIN -1 (6,5) #2
wire n5790; //IPIN -1 (6,5) #3
wire n5791; //IPIN -1 (6,5) #4
wire n5792; //IPIN -1 (6,5) #5
wire n5793; //IPIN -1 (6,5) #6
wire n5794; //IPIN -1 (6,5) #7
wire n5795; //IPIN -1 (6,5) #8
wire n5796; //IPIN -1 (6,5) #9
wire n5797; //IPIN -1 (6,5) #10
wire n5798; //IPIN -1 (6,5) #11
wire n5799; //IPIN -1 (6,5) #12
wire n5800; //IPIN -1 (6,5) #13
wire n5801; //IPIN -1 (6,5) #14
wire n5802; //IPIN -1 (6,5) #15
wire n5803; //IPIN -1 (6,5) #16
wire n5804; //IPIN -1 (6,5) #17
wire n5805; //IPIN -1 (6,5) #18
wire n5806; //IPIN -1 (6,5) #19
wire n5807; //IPIN -1 (6,5) #20
wire n5808; //IPIN -1 (6,5) #21
wire n5809; //IPIN -1 (6,5) #22
wire n5810; //IPIN -1 (6,5) #23
wire n5811; //IPIN -1 (6,5) #24
wire n5812; //IPIN -1 (6,5) #25
wire n5813; //IPIN -1 (6,5) #26
wire n5814; //IPIN -1 (6,5) #27
wire n5815; //IPIN -1 (6,5) #28
wire n5816; //IPIN -1 (6,5) #29
wire n5817; //IPIN -1 (6,5) #30
wire n5818; //IPIN -1 (6,5) #31
wire n5819; //IPIN -1 (6,5) #32
wire n5820; //IPIN -1 (6,5) #33
wire n5821; //IPIN -1 (6,5) #34
wire n5822; //IPIN -1 (6,5) #35
wire n5823; //IPIN -1 (6,5) #36
wire n5824; //IPIN -1 (6,5) #37
wire n5825; //IPIN -1 (6,5) #38
wire n5826; //IPIN -1 (6,5) #39
wire n5827; //IPIN -1 (6,5) #40
wire n5828; //IPIN -1 (6,5) #41
wire n5829; //IPIN -1 (6,5) #42
wire n5830; //IPIN -1 (6,5) #43
wire n5831; //IPIN -1 (6,5) #44
wire n5832; //IPIN -1 (6,5) #45
wire n5833; //IPIN -1 (6,5) #46
wire n5834; //IPIN -1 (6,5) #47
wire n5835; //IPIN -1 (6,5) #48
wire n5836; //IPIN -1 (6,5) #49
wire n5837; //IPIN -1 (6,5) #50
wire n5838; //IPIN -1 (6,5) #51
wire n5839; //OPIN -1 (6,5) #52
wire n5840; //OPIN -1 (6,5) #53
wire n5841; //OPIN -1 (6,5) #54
wire n5842; //OPIN -1 (6,5) #55
wire n5843; //OPIN -1 (6,5) #56
wire n5844; //OPIN -1 (6,5) #57
wire n5845; //OPIN -1 (6,5) #58
wire n5846; //OPIN -1 (6,5) #59
wire n5847; //OPIN -1 (6,5) #60
wire n5848; //OPIN -1 (6,5) #61
wire n5849; //OPIN -1 (6,5) #62
wire n5850; //OPIN -1 (6,5) #63
wire n5851; //OPIN -1 (6,5) #64
wire n5852; //OPIN -1 (6,5) #65
wire n5853; //OPIN -1 (6,5) #66
wire n5854; //OPIN -1 (6,5) #67
wire n5855; //OPIN -1 (6,5) #68
wire n5856; //OPIN -1 (6,5) #69
wire n5857; //OPIN -1 (6,5) #70
wire n5858; //OPIN -1 (6,5) #71
wire n5859; //IPIN -1 (6,5) #72
wire n5885; //IPIN -1 (6,6) #0
wire n5886; //IPIN -1 (6,6) #1
wire n5887; //IPIN -1 (6,6) #2
wire n5888; //IPIN -1 (6,6) #3
wire n5889; //IPIN -1 (6,6) #4
wire n5890; //IPIN -1 (6,6) #5
wire n5891; //IPIN -1 (6,6) #6
wire n5892; //IPIN -1 (6,6) #7
wire n5893; //IPIN -1 (6,6) #8
wire n5894; //IPIN -1 (6,6) #9
wire n5895; //IPIN -1 (6,6) #10
wire n5896; //IPIN -1 (6,6) #11
wire n5897; //IPIN -1 (6,6) #12
wire n5898; //IPIN -1 (6,6) #13
wire n5899; //IPIN -1 (6,6) #14
wire n5900; //IPIN -1 (6,6) #15
wire n5901; //IPIN -1 (6,6) #16
wire n5902; //IPIN -1 (6,6) #17
wire n5903; //IPIN -1 (6,6) #18
wire n5904; //IPIN -1 (6,6) #19
wire n5905; //IPIN -1 (6,6) #20
wire n5906; //IPIN -1 (6,6) #21
wire n5907; //IPIN -1 (6,6) #22
wire n5908; //IPIN -1 (6,6) #23
wire n5909; //IPIN -1 (6,6) #24
wire n5910; //IPIN -1 (6,6) #25
wire n5911; //IPIN -1 (6,6) #26
wire n5912; //IPIN -1 (6,6) #27
wire n5913; //IPIN -1 (6,6) #28
wire n5914; //IPIN -1 (6,6) #29
wire n5915; //IPIN -1 (6,6) #30
wire n5916; //IPIN -1 (6,6) #31
wire n5917; //IPIN -1 (6,6) #32
wire n5918; //IPIN -1 (6,6) #33
wire n5919; //IPIN -1 (6,6) #34
wire n5920; //IPIN -1 (6,6) #35
wire n5921; //IPIN -1 (6,6) #36
wire n5922; //IPIN -1 (6,6) #37
wire n5923; //IPIN -1 (6,6) #38
wire n5924; //IPIN -1 (6,6) #39
wire n5925; //IPIN -1 (6,6) #40
wire n5926; //IPIN -1 (6,6) #41
wire n5927; //IPIN -1 (6,6) #42
wire n5928; //IPIN -1 (6,6) #43
wire n5929; //IPIN -1 (6,6) #44
wire n5930; //IPIN -1 (6,6) #45
wire n5931; //IPIN -1 (6,6) #46
wire n5932; //IPIN -1 (6,6) #47
wire n5933; //IPIN -1 (6,6) #48
wire n5934; //IPIN -1 (6,6) #49
wire n5935; //IPIN -1 (6,6) #50
wire n5936; //IPIN -1 (6,6) #51
wire n5937; //OPIN -1 (6,6) #52
wire n5938; //OPIN -1 (6,6) #53
wire n5939; //OPIN -1 (6,6) #54
wire n5940; //OPIN -1 (6,6) #55
wire n5941; //OPIN -1 (6,6) #56
wire n5942; //OPIN -1 (6,6) #57
wire n5943; //OPIN -1 (6,6) #58
wire n5944; //OPIN -1 (6,6) #59
wire n5945; //OPIN -1 (6,6) #60
wire n5946; //OPIN -1 (6,6) #61
wire n5947; //OPIN -1 (6,6) #62
wire n5948; //OPIN -1 (6,6) #63
wire n5949; //OPIN -1 (6,6) #64
wire n5950; //OPIN -1 (6,6) #65
wire n5951; //OPIN -1 (6,6) #66
wire n5952; //OPIN -1 (6,6) #67
wire n5953; //OPIN -1 (6,6) #68
wire n5954; //OPIN -1 (6,6) #69
wire n5955; //OPIN -1 (6,6) #70
wire n5956; //OPIN -1 (6,6) #71
wire n5957; //IPIN -1 (6,6) #72
wire n5983; //IPIN -1 (6,7) #0
wire n5984; //IPIN -1 (6,7) #1
wire n5985; //IPIN -1 (6,7) #2
wire n5986; //IPIN -1 (6,7) #3
wire n5987; //IPIN -1 (6,7) #4
wire n5988; //IPIN -1 (6,7) #5
wire n5989; //IPIN -1 (6,7) #6
wire n5990; //IPIN -1 (6,7) #7
wire n5991; //IPIN -1 (6,7) #8
wire n5992; //IPIN -1 (6,7) #9
wire n5993; //IPIN -1 (6,7) #10
wire n5994; //IPIN -1 (6,7) #11
wire n5995; //IPIN -1 (6,7) #12
wire n5996; //IPIN -1 (6,7) #13
wire n5997; //IPIN -1 (6,7) #14
wire n5998; //IPIN -1 (6,7) #15
wire n5999; //IPIN -1 (6,7) #16
wire n6000; //IPIN -1 (6,7) #17
wire n6001; //IPIN -1 (6,7) #18
wire n6002; //IPIN -1 (6,7) #19
wire n6003; //IPIN -1 (6,7) #20
wire n6004; //IPIN -1 (6,7) #21
wire n6005; //IPIN -1 (6,7) #22
wire n6006; //IPIN -1 (6,7) #23
wire n6007; //IPIN -1 (6,7) #24
wire n6008; //IPIN -1 (6,7) #25
wire n6009; //IPIN -1 (6,7) #26
wire n6010; //IPIN -1 (6,7) #27
wire n6011; //IPIN -1 (6,7) #28
wire n6012; //IPIN -1 (6,7) #29
wire n6013; //IPIN -1 (6,7) #30
wire n6014; //IPIN -1 (6,7) #31
wire n6015; //IPIN -1 (6,7) #32
wire n6016; //IPIN -1 (6,7) #33
wire n6017; //IPIN -1 (6,7) #34
wire n6018; //IPIN -1 (6,7) #35
wire n6019; //IPIN -1 (6,7) #36
wire n6020; //IPIN -1 (6,7) #37
wire n6021; //IPIN -1 (6,7) #38
wire n6022; //IPIN -1 (6,7) #39
wire n6023; //IPIN -1 (6,7) #40
wire n6024; //IPIN -1 (6,7) #41
wire n6025; //IPIN -1 (6,7) #42
wire n6026; //IPIN -1 (6,7) #43
wire n6027; //IPIN -1 (6,7) #44
wire n6028; //IPIN -1 (6,7) #45
wire n6029; //IPIN -1 (6,7) #46
wire n6030; //IPIN -1 (6,7) #47
wire n6031; //IPIN -1 (6,7) #48
wire n6032; //IPIN -1 (6,7) #49
wire n6033; //IPIN -1 (6,7) #50
wire n6034; //IPIN -1 (6,7) #51
wire n6035; //OPIN -1 (6,7) #52
wire n6036; //OPIN -1 (6,7) #53
wire n6037; //OPIN -1 (6,7) #54
wire n6038; //OPIN -1 (6,7) #55
wire n6039; //OPIN -1 (6,7) #56
wire n6040; //OPIN -1 (6,7) #57
wire n6041; //OPIN -1 (6,7) #58
wire n6042; //OPIN -1 (6,7) #59
wire n6043; //OPIN -1 (6,7) #60
wire n6044; //OPIN -1 (6,7) #61
wire n6045; //OPIN -1 (6,7) #62
wire n6046; //OPIN -1 (6,7) #63
wire n6047; //OPIN -1 (6,7) #64
wire n6048; //OPIN -1 (6,7) #65
wire n6049; //OPIN -1 (6,7) #66
wire n6050; //OPIN -1 (6,7) #67
wire n6051; //OPIN -1 (6,7) #68
wire n6052; //OPIN -1 (6,7) #69
wire n6053; //OPIN -1 (6,7) #70
wire n6054; //OPIN -1 (6,7) #71
wire n6055; //IPIN -1 (6,7) #72
wire n6081; //IPIN -1 (6,8) #0
wire n6082; //IPIN -1 (6,8) #1
wire n6083; //IPIN -1 (6,8) #2
wire n6084; //IPIN -1 (6,8) #3
wire n6085; //IPIN -1 (6,8) #4
wire n6086; //IPIN -1 (6,8) #5
wire n6087; //IPIN -1 (6,8) #6
wire n6088; //IPIN -1 (6,8) #7
wire n6089; //IPIN -1 (6,8) #8
wire n6090; //IPIN -1 (6,8) #9
wire n6091; //IPIN -1 (6,8) #10
wire n6092; //IPIN -1 (6,8) #11
wire n6093; //IPIN -1 (6,8) #12
wire n6094; //IPIN -1 (6,8) #13
wire n6095; //IPIN -1 (6,8) #14
wire n6096; //IPIN -1 (6,8) #15
wire n6097; //IPIN -1 (6,8) #16
wire n6098; //IPIN -1 (6,8) #17
wire n6099; //IPIN -1 (6,8) #18
wire n6100; //IPIN -1 (6,8) #19
wire n6101; //IPIN -1 (6,8) #20
wire n6102; //IPIN -1 (6,8) #21
wire n6103; //IPIN -1 (6,8) #22
wire n6104; //IPIN -1 (6,8) #23
wire n6105; //IPIN -1 (6,8) #24
wire n6106; //IPIN -1 (6,8) #25
wire n6107; //IPIN -1 (6,8) #26
wire n6108; //IPIN -1 (6,8) #27
wire n6109; //IPIN -1 (6,8) #28
wire n6110; //IPIN -1 (6,8) #29
wire n6111; //IPIN -1 (6,8) #30
wire n6112; //IPIN -1 (6,8) #31
wire n6113; //IPIN -1 (6,8) #32
wire n6114; //IPIN -1 (6,8) #33
wire n6115; //IPIN -1 (6,8) #34
wire n6116; //IPIN -1 (6,8) #35
wire n6117; //IPIN -1 (6,8) #36
wire n6118; //IPIN -1 (6,8) #37
wire n6119; //IPIN -1 (6,8) #38
wire n6120; //IPIN -1 (6,8) #39
wire n6121; //IPIN -1 (6,8) #40
wire n6122; //IPIN -1 (6,8) #41
wire n6123; //IPIN -1 (6,8) #42
wire n6124; //IPIN -1 (6,8) #43
wire n6125; //IPIN -1 (6,8) #44
wire n6126; //IPIN -1 (6,8) #45
wire n6127; //IPIN -1 (6,8) #46
wire n6128; //IPIN -1 (6,8) #47
wire n6129; //IPIN -1 (6,8) #48
wire n6130; //IPIN -1 (6,8) #49
wire n6131; //IPIN -1 (6,8) #50
wire n6132; //IPIN -1 (6,8) #51
wire n6133; //OPIN -1 (6,8) #52
wire n6134; //OPIN -1 (6,8) #53
wire n6135; //OPIN -1 (6,8) #54
wire n6136; //OPIN -1 (6,8) #55
wire n6137; //OPIN -1 (6,8) #56
wire n6138; //OPIN -1 (6,8) #57
wire n6139; //OPIN -1 (6,8) #58
wire n6140; //OPIN -1 (6,8) #59
wire n6141; //OPIN -1 (6,8) #60
wire n6142; //OPIN -1 (6,8) #61
wire n6143; //OPIN -1 (6,8) #62
wire n6144; //OPIN -1 (6,8) #63
wire n6145; //OPIN -1 (6,8) #64
wire n6146; //OPIN -1 (6,8) #65
wire n6147; //OPIN -1 (6,8) #66
wire n6148; //OPIN -1 (6,8) #67
wire n6149; //OPIN -1 (6,8) #68
wire n6150; //OPIN -1 (6,8) #69
wire n6151; //OPIN -1 (6,8) #70
wire n6152; //OPIN -1 (6,8) #71
wire n6153; //IPIN -1 (6,8) #72
wire n6179; //IPIN -1 (6,9) #0
wire n6180; //IPIN -1 (6,9) #1
wire n6181; //IPIN -1 (6,9) #2
wire n6182; //IPIN -1 (6,9) #3
wire n6183; //IPIN -1 (6,9) #4
wire n6184; //IPIN -1 (6,9) #5
wire n6185; //IPIN -1 (6,9) #6
wire n6186; //IPIN -1 (6,9) #7
wire n6187; //IPIN -1 (6,9) #8
wire n6188; //IPIN -1 (6,9) #9
wire n6189; //IPIN -1 (6,9) #10
wire n6190; //IPIN -1 (6,9) #11
wire n6191; //IPIN -1 (6,9) #12
wire n6192; //IPIN -1 (6,9) #13
wire n6193; //IPIN -1 (6,9) #14
wire n6194; //IPIN -1 (6,9) #15
wire n6195; //IPIN -1 (6,9) #16
wire n6196; //IPIN -1 (6,9) #17
wire n6197; //IPIN -1 (6,9) #18
wire n6198; //IPIN -1 (6,9) #19
wire n6199; //IPIN -1 (6,9) #20
wire n6200; //IPIN -1 (6,9) #21
wire n6201; //IPIN -1 (6,9) #22
wire n6202; //IPIN -1 (6,9) #23
wire n6203; //IPIN -1 (6,9) #24
wire n6204; //IPIN -1 (6,9) #25
wire n6205; //IPIN -1 (6,9) #26
wire n6206; //IPIN -1 (6,9) #27
wire n6207; //IPIN -1 (6,9) #28
wire n6208; //IPIN -1 (6,9) #29
wire n6209; //IPIN -1 (6,9) #30
wire n6210; //IPIN -1 (6,9) #31
wire n6211; //IPIN -1 (6,9) #32
wire n6212; //IPIN -1 (6,9) #33
wire n6213; //IPIN -1 (6,9) #34
wire n6214; //IPIN -1 (6,9) #35
wire n6215; //IPIN -1 (6,9) #36
wire n6216; //IPIN -1 (6,9) #37
wire n6217; //IPIN -1 (6,9) #38
wire n6218; //IPIN -1 (6,9) #39
wire n6219; //IPIN -1 (6,9) #40
wire n6220; //IPIN -1 (6,9) #41
wire n6221; //IPIN -1 (6,9) #42
wire n6222; //IPIN -1 (6,9) #43
wire n6223; //IPIN -1 (6,9) #44
wire n6224; //IPIN -1 (6,9) #45
wire n6225; //IPIN -1 (6,9) #46
wire n6226; //IPIN -1 (6,9) #47
wire n6227; //IPIN -1 (6,9) #48
wire n6228; //IPIN -1 (6,9) #49
wire n6229; //IPIN -1 (6,9) #50
wire n6230; //IPIN -1 (6,9) #51
wire n6231; //OPIN -1 (6,9) #52
wire n6232; //OPIN -1 (6,9) #53
wire n6233; //OPIN -1 (6,9) #54
wire n6234; //OPIN -1 (6,9) #55
wire n6235; //OPIN -1 (6,9) #56
wire n6236; //OPIN -1 (6,9) #57
wire n6237; //OPIN -1 (6,9) #58
wire n6238; //OPIN -1 (6,9) #59
wire n6239; //OPIN -1 (6,9) #60
wire n6240; //OPIN -1 (6,9) #61
wire n6241; //OPIN -1 (6,9) #62
wire n6242; //OPIN -1 (6,9) #63
wire n6243; //OPIN -1 (6,9) #64
wire n6244; //OPIN -1 (6,9) #65
wire n6245; //OPIN -1 (6,9) #66
wire n6246; //OPIN -1 (6,9) #67
wire n6247; //OPIN -1 (6,9) #68
wire n6248; //OPIN -1 (6,9) #69
wire n6249; //OPIN -1 (6,9) #70
wire n6250; //OPIN -1 (6,9) #71
wire n6251; //IPIN -1 (6,9) #72
wire n6276; //IPIN -1 (6,10) #0
wire n6277; //OPIN -1 (6,10) #1
wire n6278; //IPIN -1 (6,10) #2
wire n6279; //IPIN -1 (6,10) #3
wire n6280; //OPIN -1 (6,10) #4
wire n6281; //IPIN -1 (6,10) #5
wire n6282; //IPIN -1 (6,10) #6
wire n6283; //OPIN -1 (6,10) #7
wire n6284; //IPIN -1 (6,10) #8
wire n6285; //IPIN -1 (6,10) #9
wire n6286; //OPIN -1 (6,10) #10
wire n6287; //IPIN -1 (6,10) #11
wire n6288; //IPIN -1 (6,10) #12
wire n6289; //OPIN -1 (6,10) #13
wire n6290; //IPIN -1 (6,10) #14
wire n6291; //IPIN -1 (6,10) #15
wire n6292; //OPIN -1 (6,10) #16
wire n6293; //IPIN -1 (6,10) #17
wire n6294; //IPIN -1 (6,10) #18
wire n6295; //OPIN -1 (6,10) #19
wire n6296; //IPIN -1 (6,10) #20
wire n6297; //IPIN -1 (6,10) #21
wire n6298; //OPIN -1 (6,10) #22
wire n6299; //IPIN -1 (6,10) #23
wire n6324; //IPIN -1 (7,0) #0
wire n6325; //OPIN -1 (7,0) #1
wire n6326; //IPIN -1 (7,0) #2
wire n6327; //IPIN -1 (7,0) #3
wire n6328; //OPIN -1 (7,0) #4
wire n6329; //IPIN -1 (7,0) #5
wire n6330; //IPIN -1 (7,0) #6
wire n6331; //OPIN -1 (7,0) #7
wire n6332; //IPIN -1 (7,0) #8
wire n6333; //IPIN -1 (7,0) #9
wire n6334; //OPIN -1 (7,0) #10
wire n6335; //IPIN -1 (7,0) #11
wire n6336; //IPIN -1 (7,0) #12
wire n6337; //OPIN -1 (7,0) #13
wire n6338; //IPIN -1 (7,0) #14
wire n6339; //IPIN -1 (7,0) #15
wire n6340; //OPIN -1 (7,0) #16
wire n6341; //IPIN -1 (7,0) #17
wire n6342; //IPIN -1 (7,0) #18
wire n6343; //OPIN -1 (7,0) #19
wire n6344; //IPIN -1 (7,0) #20
wire n6345; //IPIN -1 (7,0) #21
wire n6346; //OPIN -1 (7,0) #22
wire n6347; //IPIN -1 (7,0) #23
wire n6373; //IPIN -1 (7,1) #0
wire n6374; //IPIN -1 (7,1) #1
wire n6375; //IPIN -1 (7,1) #2
wire n6376; //IPIN -1 (7,1) #3
wire n6377; //IPIN -1 (7,1) #4
wire n6378; //IPIN -1 (7,1) #5
wire n6379; //IPIN -1 (7,1) #6
wire n6380; //IPIN -1 (7,1) #7
wire n6381; //IPIN -1 (7,1) #8
wire n6382; //IPIN -1 (7,1) #9
wire n6383; //IPIN -1 (7,1) #10
wire n6384; //IPIN -1 (7,1) #11
wire n6385; //IPIN -1 (7,1) #12
wire n6386; //IPIN -1 (7,1) #13
wire n6387; //IPIN -1 (7,1) #14
wire n6388; //IPIN -1 (7,1) #15
wire n6389; //IPIN -1 (7,1) #16
wire n6390; //IPIN -1 (7,1) #17
wire n6391; //IPIN -1 (7,1) #18
wire n6392; //IPIN -1 (7,1) #19
wire n6393; //IPIN -1 (7,1) #20
wire n6394; //IPIN -1 (7,1) #21
wire n6395; //IPIN -1 (7,1) #22
wire n6396; //IPIN -1 (7,1) #23
wire n6397; //IPIN -1 (7,1) #24
wire n6398; //IPIN -1 (7,1) #25
wire n6399; //IPIN -1 (7,1) #26
wire n6400; //IPIN -1 (7,1) #27
wire n6401; //IPIN -1 (7,1) #28
wire n6402; //IPIN -1 (7,1) #29
wire n6403; //IPIN -1 (7,1) #30
wire n6404; //IPIN -1 (7,1) #31
wire n6405; //IPIN -1 (7,1) #32
wire n6406; //IPIN -1 (7,1) #33
wire n6407; //IPIN -1 (7,1) #34
wire n6408; //IPIN -1 (7,1) #35
wire n6409; //IPIN -1 (7,1) #36
wire n6410; //IPIN -1 (7,1) #37
wire n6411; //IPIN -1 (7,1) #38
wire n6412; //IPIN -1 (7,1) #39
wire n6413; //IPIN -1 (7,1) #40
wire n6414; //IPIN -1 (7,1) #41
wire n6415; //IPIN -1 (7,1) #42
wire n6416; //IPIN -1 (7,1) #43
wire n6417; //IPIN -1 (7,1) #44
wire n6418; //IPIN -1 (7,1) #45
wire n6419; //IPIN -1 (7,1) #46
wire n6420; //IPIN -1 (7,1) #47
wire n6421; //IPIN -1 (7,1) #48
wire n6422; //IPIN -1 (7,1) #49
wire n6423; //IPIN -1 (7,1) #50
wire n6424; //IPIN -1 (7,1) #51
wire n6425; //OPIN -1 (7,1) #52
wire n6426; //OPIN -1 (7,1) #53
wire n6427; //OPIN -1 (7,1) #54
wire n6428; //OPIN -1 (7,1) #55
wire n6429; //OPIN -1 (7,1) #56
wire n6430; //OPIN -1 (7,1) #57
wire n6431; //OPIN -1 (7,1) #58
wire n6432; //OPIN -1 (7,1) #59
wire n6433; //OPIN -1 (7,1) #60
wire n6434; //OPIN -1 (7,1) #61
wire n6435; //OPIN -1 (7,1) #62
wire n6436; //OPIN -1 (7,1) #63
wire n6437; //OPIN -1 (7,1) #64
wire n6438; //OPIN -1 (7,1) #65
wire n6439; //OPIN -1 (7,1) #66
wire n6440; //OPIN -1 (7,1) #67
wire n6441; //OPIN -1 (7,1) #68
wire n6442; //OPIN -1 (7,1) #69
wire n6443; //OPIN -1 (7,1) #70
wire n6444; //OPIN -1 (7,1) #71
wire n6445; //IPIN -1 (7,1) #72
wire n6471; //IPIN -1 (7,2) #0
wire n6472; //IPIN -1 (7,2) #1
wire n6473; //IPIN -1 (7,2) #2
wire n6474; //IPIN -1 (7,2) #3
wire n6475; //IPIN -1 (7,2) #4
wire n6476; //IPIN -1 (7,2) #5
wire n6477; //IPIN -1 (7,2) #6
wire n6478; //IPIN -1 (7,2) #7
wire n6479; //IPIN -1 (7,2) #8
wire n6480; //IPIN -1 (7,2) #9
wire n6481; //IPIN -1 (7,2) #10
wire n6482; //IPIN -1 (7,2) #11
wire n6483; //IPIN -1 (7,2) #12
wire n6484; //IPIN -1 (7,2) #13
wire n6485; //IPIN -1 (7,2) #14
wire n6486; //IPIN -1 (7,2) #15
wire n6487; //IPIN -1 (7,2) #16
wire n6488; //IPIN -1 (7,2) #17
wire n6489; //IPIN -1 (7,2) #18
wire n6490; //IPIN -1 (7,2) #19
wire n6491; //IPIN -1 (7,2) #20
wire n6492; //IPIN -1 (7,2) #21
wire n6493; //IPIN -1 (7,2) #22
wire n6494; //IPIN -1 (7,2) #23
wire n6495; //IPIN -1 (7,2) #24
wire n6496; //IPIN -1 (7,2) #25
wire n6497; //IPIN -1 (7,2) #26
wire n6498; //IPIN -1 (7,2) #27
wire n6499; //IPIN -1 (7,2) #28
wire n6500; //IPIN -1 (7,2) #29
wire n6501; //IPIN -1 (7,2) #30
wire n6502; //IPIN -1 (7,2) #31
wire n6503; //IPIN -1 (7,2) #32
wire n6504; //IPIN -1 (7,2) #33
wire n6505; //IPIN -1 (7,2) #34
wire n6506; //IPIN -1 (7,2) #35
wire n6507; //IPIN -1 (7,2) #36
wire n6508; //IPIN -1 (7,2) #37
wire n6509; //IPIN -1 (7,2) #38
wire n6510; //IPIN -1 (7,2) #39
wire n6511; //IPIN -1 (7,2) #40
wire n6512; //IPIN -1 (7,2) #41
wire n6513; //IPIN -1 (7,2) #42
wire n6514; //IPIN -1 (7,2) #43
wire n6515; //IPIN -1 (7,2) #44
wire n6516; //IPIN -1 (7,2) #45
wire n6517; //IPIN -1 (7,2) #46
wire n6518; //IPIN -1 (7,2) #47
wire n6519; //IPIN -1 (7,2) #48
wire n6520; //IPIN -1 (7,2) #49
wire n6521; //IPIN -1 (7,2) #50
wire n6522; //IPIN -1 (7,2) #51
wire n6523; //OPIN -1 (7,2) #52
wire n6524; //OPIN -1 (7,2) #53
wire n6525; //OPIN -1 (7,2) #54
wire n6526; //OPIN -1 (7,2) #55
wire n6527; //OPIN -1 (7,2) #56
wire n6528; //OPIN -1 (7,2) #57
wire n6529; //OPIN -1 (7,2) #58
wire n6530; //OPIN -1 (7,2) #59
wire n6531; //OPIN -1 (7,2) #60
wire n6532; //OPIN -1 (7,2) #61
wire n6533; //OPIN -1 (7,2) #62
wire n6534; //OPIN -1 (7,2) #63
wire n6535; //OPIN -1 (7,2) #64
wire n6536; //OPIN -1 (7,2) #65
wire n6537; //OPIN -1 (7,2) #66
wire n6538; //OPIN -1 (7,2) #67
wire n6539; //OPIN -1 (7,2) #68
wire n6540; //OPIN -1 (7,2) #69
wire n6541; //OPIN -1 (7,2) #70
wire n6542; //OPIN -1 (7,2) #71
wire n6543; //IPIN -1 (7,2) #72
wire n6569; //IPIN -1 (7,3) #0
wire n6570; //IPIN -1 (7,3) #1
wire n6571; //IPIN -1 (7,3) #2
wire n6572; //IPIN -1 (7,3) #3
wire n6573; //IPIN -1 (7,3) #4
wire n6574; //IPIN -1 (7,3) #5
wire n6575; //IPIN -1 (7,3) #6
wire n6576; //IPIN -1 (7,3) #7
wire n6577; //IPIN -1 (7,3) #8
wire n6578; //IPIN -1 (7,3) #9
wire n6579; //IPIN -1 (7,3) #10
wire n6580; //IPIN -1 (7,3) #11
wire n6581; //IPIN -1 (7,3) #12
wire n6582; //IPIN -1 (7,3) #13
wire n6583; //IPIN -1 (7,3) #14
wire n6584; //IPIN -1 (7,3) #15
wire n6585; //IPIN -1 (7,3) #16
wire n6586; //IPIN -1 (7,3) #17
wire n6587; //IPIN -1 (7,3) #18
wire n6588; //IPIN -1 (7,3) #19
wire n6589; //IPIN -1 (7,3) #20
wire n6590; //IPIN -1 (7,3) #21
wire n6591; //IPIN -1 (7,3) #22
wire n6592; //IPIN -1 (7,3) #23
wire n6593; //IPIN -1 (7,3) #24
wire n6594; //IPIN -1 (7,3) #25
wire n6595; //IPIN -1 (7,3) #26
wire n6596; //IPIN -1 (7,3) #27
wire n6597; //IPIN -1 (7,3) #28
wire n6598; //IPIN -1 (7,3) #29
wire n6599; //IPIN -1 (7,3) #30
wire n6600; //IPIN -1 (7,3) #31
wire n6601; //IPIN -1 (7,3) #32
wire n6602; //IPIN -1 (7,3) #33
wire n6603; //IPIN -1 (7,3) #34
wire n6604; //IPIN -1 (7,3) #35
wire n6605; //IPIN -1 (7,3) #36
wire n6606; //IPIN -1 (7,3) #37
wire n6607; //IPIN -1 (7,3) #38
wire n6608; //IPIN -1 (7,3) #39
wire n6609; //IPIN -1 (7,3) #40
wire n6610; //IPIN -1 (7,3) #41
wire n6611; //IPIN -1 (7,3) #42
wire n6612; //IPIN -1 (7,3) #43
wire n6613; //IPIN -1 (7,3) #44
wire n6614; //IPIN -1 (7,3) #45
wire n6615; //IPIN -1 (7,3) #46
wire n6616; //IPIN -1 (7,3) #47
wire n6617; //IPIN -1 (7,3) #48
wire n6618; //IPIN -1 (7,3) #49
wire n6619; //IPIN -1 (7,3) #50
wire n6620; //IPIN -1 (7,3) #51
wire n6621; //OPIN -1 (7,3) #52
wire n6622; //OPIN -1 (7,3) #53
wire n6623; //OPIN -1 (7,3) #54
wire n6624; //OPIN -1 (7,3) #55
wire n6625; //OPIN -1 (7,3) #56
wire n6626; //OPIN -1 (7,3) #57
wire n6627; //OPIN -1 (7,3) #58
wire n6628; //OPIN -1 (7,3) #59
wire n6629; //OPIN -1 (7,3) #60
wire n6630; //OPIN -1 (7,3) #61
wire n6631; //OPIN -1 (7,3) #62
wire n6632; //OPIN -1 (7,3) #63
wire n6633; //OPIN -1 (7,3) #64
wire n6634; //OPIN -1 (7,3) #65
wire n6635; //OPIN -1 (7,3) #66
wire n6636; //OPIN -1 (7,3) #67
wire n6637; //OPIN -1 (7,3) #68
wire n6638; //OPIN -1 (7,3) #69
wire n6639; //OPIN -1 (7,3) #70
wire n6640; //OPIN -1 (7,3) #71
wire n6641; //IPIN -1 (7,3) #72
wire n6667; //IPIN -1 (7,4) #0
wire n6668; //IPIN -1 (7,4) #1
wire n6669; //IPIN -1 (7,4) #2
wire n6670; //IPIN -1 (7,4) #3
wire n6671; //IPIN -1 (7,4) #4
wire n6672; //IPIN -1 (7,4) #5
wire n6673; //IPIN -1 (7,4) #6
wire n6674; //IPIN -1 (7,4) #7
wire n6675; //IPIN -1 (7,4) #8
wire n6676; //IPIN -1 (7,4) #9
wire n6677; //IPIN -1 (7,4) #10
wire n6678; //IPIN -1 (7,4) #11
wire n6679; //IPIN -1 (7,4) #12
wire n6680; //IPIN -1 (7,4) #13
wire n6681; //IPIN -1 (7,4) #14
wire n6682; //IPIN -1 (7,4) #15
wire n6683; //IPIN -1 (7,4) #16
wire n6684; //IPIN -1 (7,4) #17
wire n6685; //IPIN -1 (7,4) #18
wire n6686; //IPIN -1 (7,4) #19
wire n6687; //IPIN -1 (7,4) #20
wire n6688; //IPIN -1 (7,4) #21
wire n6689; //IPIN -1 (7,4) #22
wire n6690; //IPIN -1 (7,4) #23
wire n6691; //IPIN -1 (7,4) #24
wire n6692; //IPIN -1 (7,4) #25
wire n6693; //IPIN -1 (7,4) #26
wire n6694; //IPIN -1 (7,4) #27
wire n6695; //IPIN -1 (7,4) #28
wire n6696; //IPIN -1 (7,4) #29
wire n6697; //IPIN -1 (7,4) #30
wire n6698; //IPIN -1 (7,4) #31
wire n6699; //IPIN -1 (7,4) #32
wire n6700; //IPIN -1 (7,4) #33
wire n6701; //IPIN -1 (7,4) #34
wire n6702; //IPIN -1 (7,4) #35
wire n6703; //IPIN -1 (7,4) #36
wire n6704; //IPIN -1 (7,4) #37
wire n6705; //IPIN -1 (7,4) #38
wire n6706; //IPIN -1 (7,4) #39
wire n6707; //IPIN -1 (7,4) #40
wire n6708; //IPIN -1 (7,4) #41
wire n6709; //IPIN -1 (7,4) #42
wire n6710; //IPIN -1 (7,4) #43
wire n6711; //IPIN -1 (7,4) #44
wire n6712; //IPIN -1 (7,4) #45
wire n6713; //IPIN -1 (7,4) #46
wire n6714; //IPIN -1 (7,4) #47
wire n6715; //IPIN -1 (7,4) #48
wire n6716; //IPIN -1 (7,4) #49
wire n6717; //IPIN -1 (7,4) #50
wire n6718; //IPIN -1 (7,4) #51
wire n6719; //OPIN -1 (7,4) #52
wire n6720; //OPIN -1 (7,4) #53
wire n6721; //OPIN -1 (7,4) #54
wire n6722; //OPIN -1 (7,4) #55
wire n6723; //OPIN -1 (7,4) #56
wire n6724; //OPIN -1 (7,4) #57
wire n6725; //OPIN -1 (7,4) #58
wire n6726; //OPIN -1 (7,4) #59
wire n6727; //OPIN -1 (7,4) #60
wire n6728; //OPIN -1 (7,4) #61
wire n6729; //OPIN -1 (7,4) #62
wire n6730; //OPIN -1 (7,4) #63
wire n6731; //OPIN -1 (7,4) #64
wire n6732; //OPIN -1 (7,4) #65
wire n6733; //OPIN -1 (7,4) #66
wire n6734; //OPIN -1 (7,4) #67
wire n6735; //OPIN -1 (7,4) #68
wire n6736; //OPIN -1 (7,4) #69
wire n6737; //OPIN -1 (7,4) #70
wire n6738; //OPIN -1 (7,4) #71
wire n6739; //IPIN -1 (7,4) #72
wire n6765; //IPIN -1 (7,5) #0
wire n6766; //IPIN -1 (7,5) #1
wire n6767; //IPIN -1 (7,5) #2
wire n6768; //IPIN -1 (7,5) #3
wire n6769; //IPIN -1 (7,5) #4
wire n6770; //IPIN -1 (7,5) #5
wire n6771; //IPIN -1 (7,5) #6
wire n6772; //IPIN -1 (7,5) #7
wire n6773; //IPIN -1 (7,5) #8
wire n6774; //IPIN -1 (7,5) #9
wire n6775; //IPIN -1 (7,5) #10
wire n6776; //IPIN -1 (7,5) #11
wire n6777; //IPIN -1 (7,5) #12
wire n6778; //IPIN -1 (7,5) #13
wire n6779; //IPIN -1 (7,5) #14
wire n6780; //IPIN -1 (7,5) #15
wire n6781; //IPIN -1 (7,5) #16
wire n6782; //IPIN -1 (7,5) #17
wire n6783; //IPIN -1 (7,5) #18
wire n6784; //IPIN -1 (7,5) #19
wire n6785; //IPIN -1 (7,5) #20
wire n6786; //IPIN -1 (7,5) #21
wire n6787; //IPIN -1 (7,5) #22
wire n6788; //IPIN -1 (7,5) #23
wire n6789; //IPIN -1 (7,5) #24
wire n6790; //IPIN -1 (7,5) #25
wire n6791; //IPIN -1 (7,5) #26
wire n6792; //IPIN -1 (7,5) #27
wire n6793; //IPIN -1 (7,5) #28
wire n6794; //IPIN -1 (7,5) #29
wire n6795; //IPIN -1 (7,5) #30
wire n6796; //IPIN -1 (7,5) #31
wire n6797; //IPIN -1 (7,5) #32
wire n6798; //IPIN -1 (7,5) #33
wire n6799; //IPIN -1 (7,5) #34
wire n6800; //IPIN -1 (7,5) #35
wire n6801; //IPIN -1 (7,5) #36
wire n6802; //IPIN -1 (7,5) #37
wire n6803; //IPIN -1 (7,5) #38
wire n6804; //IPIN -1 (7,5) #39
wire n6805; //IPIN -1 (7,5) #40
wire n6806; //IPIN -1 (7,5) #41
wire n6807; //IPIN -1 (7,5) #42
wire n6808; //IPIN -1 (7,5) #43
wire n6809; //IPIN -1 (7,5) #44
wire n6810; //IPIN -1 (7,5) #45
wire n6811; //IPIN -1 (7,5) #46
wire n6812; //IPIN -1 (7,5) #47
wire n6813; //IPIN -1 (7,5) #48
wire n6814; //IPIN -1 (7,5) #49
wire n6815; //IPIN -1 (7,5) #50
wire n6816; //IPIN -1 (7,5) #51
wire n6817; //OPIN -1 (7,5) #52
wire n6818; //OPIN -1 (7,5) #53
wire n6819; //OPIN -1 (7,5) #54
wire n6820; //OPIN -1 (7,5) #55
wire n6821; //OPIN -1 (7,5) #56
wire n6822; //OPIN -1 (7,5) #57
wire n6823; //OPIN -1 (7,5) #58
wire n6824; //OPIN -1 (7,5) #59
wire n6825; //OPIN -1 (7,5) #60
wire n6826; //OPIN -1 (7,5) #61
wire n6827; //OPIN -1 (7,5) #62
wire n6828; //OPIN -1 (7,5) #63
wire n6829; //OPIN -1 (7,5) #64
wire n6830; //OPIN -1 (7,5) #65
wire n6831; //OPIN -1 (7,5) #66
wire n6832; //OPIN -1 (7,5) #67
wire n6833; //OPIN -1 (7,5) #68
wire n6834; //OPIN -1 (7,5) #69
wire n6835; //OPIN -1 (7,5) #70
wire n6836; //OPIN -1 (7,5) #71
wire n6837; //IPIN -1 (7,5) #72
wire n6863; //IPIN -1 (7,6) #0
wire n6864; //IPIN -1 (7,6) #1
wire n6865; //IPIN -1 (7,6) #2
wire n6866; //IPIN -1 (7,6) #3
wire n6867; //IPIN -1 (7,6) #4
wire n6868; //IPIN -1 (7,6) #5
wire n6869; //IPIN -1 (7,6) #6
wire n6870; //IPIN -1 (7,6) #7
wire n6871; //IPIN -1 (7,6) #8
wire n6872; //IPIN -1 (7,6) #9
wire n6873; //IPIN -1 (7,6) #10
wire n6874; //IPIN -1 (7,6) #11
wire n6875; //IPIN -1 (7,6) #12
wire n6876; //IPIN -1 (7,6) #13
wire n6877; //IPIN -1 (7,6) #14
wire n6878; //IPIN -1 (7,6) #15
wire n6879; //IPIN -1 (7,6) #16
wire n6880; //IPIN -1 (7,6) #17
wire n6881; //IPIN -1 (7,6) #18
wire n6882; //IPIN -1 (7,6) #19
wire n6883; //IPIN -1 (7,6) #20
wire n6884; //IPIN -1 (7,6) #21
wire n6885; //IPIN -1 (7,6) #22
wire n6886; //IPIN -1 (7,6) #23
wire n6887; //IPIN -1 (7,6) #24
wire n6888; //IPIN -1 (7,6) #25
wire n6889; //IPIN -1 (7,6) #26
wire n6890; //IPIN -1 (7,6) #27
wire n6891; //IPIN -1 (7,6) #28
wire n6892; //IPIN -1 (7,6) #29
wire n6893; //IPIN -1 (7,6) #30
wire n6894; //IPIN -1 (7,6) #31
wire n6895; //IPIN -1 (7,6) #32
wire n6896; //IPIN -1 (7,6) #33
wire n6897; //IPIN -1 (7,6) #34
wire n6898; //IPIN -1 (7,6) #35
wire n6899; //IPIN -1 (7,6) #36
wire n6900; //IPIN -1 (7,6) #37
wire n6901; //IPIN -1 (7,6) #38
wire n6902; //IPIN -1 (7,6) #39
wire n6903; //IPIN -1 (7,6) #40
wire n6904; //IPIN -1 (7,6) #41
wire n6905; //IPIN -1 (7,6) #42
wire n6906; //IPIN -1 (7,6) #43
wire n6907; //IPIN -1 (7,6) #44
wire n6908; //IPIN -1 (7,6) #45
wire n6909; //IPIN -1 (7,6) #46
wire n6910; //IPIN -1 (7,6) #47
wire n6911; //IPIN -1 (7,6) #48
wire n6912; //IPIN -1 (7,6) #49
wire n6913; //IPIN -1 (7,6) #50
wire n6914; //IPIN -1 (7,6) #51
wire n6915; //OPIN -1 (7,6) #52
wire n6916; //OPIN -1 (7,6) #53
wire n6917; //OPIN -1 (7,6) #54
wire n6918; //OPIN -1 (7,6) #55
wire n6919; //OPIN -1 (7,6) #56
wire n6920; //OPIN -1 (7,6) #57
wire n6921; //OPIN -1 (7,6) #58
wire n6922; //OPIN -1 (7,6) #59
wire n6923; //OPIN -1 (7,6) #60
wire n6924; //OPIN -1 (7,6) #61
wire n6925; //OPIN -1 (7,6) #62
wire n6926; //OPIN -1 (7,6) #63
wire n6927; //OPIN -1 (7,6) #64
wire n6928; //OPIN -1 (7,6) #65
wire n6929; //OPIN -1 (7,6) #66
wire n6930; //OPIN -1 (7,6) #67
wire n6931; //OPIN -1 (7,6) #68
wire n6932; //OPIN -1 (7,6) #69
wire n6933; //OPIN -1 (7,6) #70
wire n6934; //OPIN -1 (7,6) #71
wire n6935; //IPIN -1 (7,6) #72
wire n6961; //IPIN -1 (7,7) #0
wire n6962; //IPIN -1 (7,7) #1
wire n6963; //IPIN -1 (7,7) #2
wire n6964; //IPIN -1 (7,7) #3
wire n6965; //IPIN -1 (7,7) #4
wire n6966; //IPIN -1 (7,7) #5
wire n6967; //IPIN -1 (7,7) #6
wire n6968; //IPIN -1 (7,7) #7
wire n6969; //IPIN -1 (7,7) #8
wire n6970; //IPIN -1 (7,7) #9
wire n6971; //IPIN -1 (7,7) #10
wire n6972; //IPIN -1 (7,7) #11
wire n6973; //IPIN -1 (7,7) #12
wire n6974; //IPIN -1 (7,7) #13
wire n6975; //IPIN -1 (7,7) #14
wire n6976; //IPIN -1 (7,7) #15
wire n6977; //IPIN -1 (7,7) #16
wire n6978; //IPIN -1 (7,7) #17
wire n6979; //IPIN -1 (7,7) #18
wire n6980; //IPIN -1 (7,7) #19
wire n6981; //IPIN -1 (7,7) #20
wire n6982; //IPIN -1 (7,7) #21
wire n6983; //IPIN -1 (7,7) #22
wire n6984; //IPIN -1 (7,7) #23
wire n6985; //IPIN -1 (7,7) #24
wire n6986; //IPIN -1 (7,7) #25
wire n6987; //IPIN -1 (7,7) #26
wire n6988; //IPIN -1 (7,7) #27
wire n6989; //IPIN -1 (7,7) #28
wire n6990; //IPIN -1 (7,7) #29
wire n6991; //IPIN -1 (7,7) #30
wire n6992; //IPIN -1 (7,7) #31
wire n6993; //IPIN -1 (7,7) #32
wire n6994; //IPIN -1 (7,7) #33
wire n6995; //IPIN -1 (7,7) #34
wire n6996; //IPIN -1 (7,7) #35
wire n6997; //IPIN -1 (7,7) #36
wire n6998; //IPIN -1 (7,7) #37
wire n6999; //IPIN -1 (7,7) #38
wire n7000; //IPIN -1 (7,7) #39
wire n7001; //IPIN -1 (7,7) #40
wire n7002; //IPIN -1 (7,7) #41
wire n7003; //IPIN -1 (7,7) #42
wire n7004; //IPIN -1 (7,7) #43
wire n7005; //IPIN -1 (7,7) #44
wire n7006; //IPIN -1 (7,7) #45
wire n7007; //IPIN -1 (7,7) #46
wire n7008; //IPIN -1 (7,7) #47
wire n7009; //IPIN -1 (7,7) #48
wire n7010; //IPIN -1 (7,7) #49
wire n7011; //IPIN -1 (7,7) #50
wire n7012; //IPIN -1 (7,7) #51
wire n7013; //OPIN -1 (7,7) #52
wire n7014; //OPIN -1 (7,7) #53
wire n7015; //OPIN -1 (7,7) #54
wire n7016; //OPIN -1 (7,7) #55
wire n7017; //OPIN -1 (7,7) #56
wire n7018; //OPIN -1 (7,7) #57
wire n7019; //OPIN -1 (7,7) #58
wire n7020; //OPIN -1 (7,7) #59
wire n7021; //OPIN -1 (7,7) #60
wire n7022; //OPIN -1 (7,7) #61
wire n7023; //OPIN -1 (7,7) #62
wire n7024; //OPIN -1 (7,7) #63
wire n7025; //OPIN -1 (7,7) #64
wire n7026; //OPIN -1 (7,7) #65
wire n7027; //OPIN -1 (7,7) #66
wire n7028; //OPIN -1 (7,7) #67
wire n7029; //OPIN -1 (7,7) #68
wire n7030; //OPIN -1 (7,7) #69
wire n7031; //OPIN -1 (7,7) #70
wire n7032; //OPIN -1 (7,7) #71
wire n7033; //IPIN -1 (7,7) #72
wire n7059; //IPIN -1 (7,8) #0
wire n7060; //IPIN -1 (7,8) #1
wire n7061; //IPIN -1 (7,8) #2
wire n7062; //IPIN -1 (7,8) #3
wire n7063; //IPIN -1 (7,8) #4
wire n7064; //IPIN -1 (7,8) #5
wire n7065; //IPIN -1 (7,8) #6
wire n7066; //IPIN -1 (7,8) #7
wire n7067; //IPIN -1 (7,8) #8
wire n7068; //IPIN -1 (7,8) #9
wire n7069; //IPIN -1 (7,8) #10
wire n7070; //IPIN -1 (7,8) #11
wire n7071; //IPIN -1 (7,8) #12
wire n7072; //IPIN -1 (7,8) #13
wire n7073; //IPIN -1 (7,8) #14
wire n7074; //IPIN -1 (7,8) #15
wire n7075; //IPIN -1 (7,8) #16
wire n7076; //IPIN -1 (7,8) #17
wire n7077; //IPIN -1 (7,8) #18
wire n7078; //IPIN -1 (7,8) #19
wire n7079; //IPIN -1 (7,8) #20
wire n7080; //IPIN -1 (7,8) #21
wire n7081; //IPIN -1 (7,8) #22
wire n7082; //IPIN -1 (7,8) #23
wire n7083; //IPIN -1 (7,8) #24
wire n7084; //IPIN -1 (7,8) #25
wire n7085; //IPIN -1 (7,8) #26
wire n7086; //IPIN -1 (7,8) #27
wire n7087; //IPIN -1 (7,8) #28
wire n7088; //IPIN -1 (7,8) #29
wire n7089; //IPIN -1 (7,8) #30
wire n7090; //IPIN -1 (7,8) #31
wire n7091; //IPIN -1 (7,8) #32
wire n7092; //IPIN -1 (7,8) #33
wire n7093; //IPIN -1 (7,8) #34
wire n7094; //IPIN -1 (7,8) #35
wire n7095; //IPIN -1 (7,8) #36
wire n7096; //IPIN -1 (7,8) #37
wire n7097; //IPIN -1 (7,8) #38
wire n7098; //IPIN -1 (7,8) #39
wire n7099; //IPIN -1 (7,8) #40
wire n7100; //IPIN -1 (7,8) #41
wire n7101; //IPIN -1 (7,8) #42
wire n7102; //IPIN -1 (7,8) #43
wire n7103; //IPIN -1 (7,8) #44
wire n7104; //IPIN -1 (7,8) #45
wire n7105; //IPIN -1 (7,8) #46
wire n7106; //IPIN -1 (7,8) #47
wire n7107; //IPIN -1 (7,8) #48
wire n7108; //IPIN -1 (7,8) #49
wire n7109; //IPIN -1 (7,8) #50
wire n7110; //IPIN -1 (7,8) #51
wire n7111; //OPIN -1 (7,8) #52
wire n7112; //OPIN -1 (7,8) #53
wire n7113; //OPIN -1 (7,8) #54
wire n7114; //OPIN -1 (7,8) #55
wire n7115; //OPIN -1 (7,8) #56
wire n7116; //OPIN -1 (7,8) #57
wire n7117; //OPIN -1 (7,8) #58
wire n7118; //OPIN -1 (7,8) #59
wire n7119; //OPIN -1 (7,8) #60
wire n7120; //OPIN -1 (7,8) #61
wire n7121; //OPIN -1 (7,8) #62
wire n7122; //OPIN -1 (7,8) #63
wire n7123; //OPIN -1 (7,8) #64
wire n7124; //OPIN -1 (7,8) #65
wire n7125; //OPIN -1 (7,8) #66
wire n7126; //OPIN -1 (7,8) #67
wire n7127; //OPIN -1 (7,8) #68
wire n7128; //OPIN -1 (7,8) #69
wire n7129; //OPIN -1 (7,8) #70
wire n7130; //OPIN -1 (7,8) #71
wire n7131; //IPIN -1 (7,8) #72
wire n7157; //IPIN -1 (7,9) #0
wire n7158; //IPIN -1 (7,9) #1
wire n7159; //IPIN -1 (7,9) #2
wire n7160; //IPIN -1 (7,9) #3
wire n7161; //IPIN -1 (7,9) #4
wire n7162; //IPIN -1 (7,9) #5
wire n7163; //IPIN -1 (7,9) #6
wire n7164; //IPIN -1 (7,9) #7
wire n7165; //IPIN -1 (7,9) #8
wire n7166; //IPIN -1 (7,9) #9
wire n7167; //IPIN -1 (7,9) #10
wire n7168; //IPIN -1 (7,9) #11
wire n7169; //IPIN -1 (7,9) #12
wire n7170; //IPIN -1 (7,9) #13
wire n7171; //IPIN -1 (7,9) #14
wire n7172; //IPIN -1 (7,9) #15
wire n7173; //IPIN -1 (7,9) #16
wire n7174; //IPIN -1 (7,9) #17
wire n7175; //IPIN -1 (7,9) #18
wire n7176; //IPIN -1 (7,9) #19
wire n7177; //IPIN -1 (7,9) #20
wire n7178; //IPIN -1 (7,9) #21
wire n7179; //IPIN -1 (7,9) #22
wire n7180; //IPIN -1 (7,9) #23
wire n7181; //IPIN -1 (7,9) #24
wire n7182; //IPIN -1 (7,9) #25
wire n7183; //IPIN -1 (7,9) #26
wire n7184; //IPIN -1 (7,9) #27
wire n7185; //IPIN -1 (7,9) #28
wire n7186; //IPIN -1 (7,9) #29
wire n7187; //IPIN -1 (7,9) #30
wire n7188; //IPIN -1 (7,9) #31
wire n7189; //IPIN -1 (7,9) #32
wire n7190; //IPIN -1 (7,9) #33
wire n7191; //IPIN -1 (7,9) #34
wire n7192; //IPIN -1 (7,9) #35
wire n7193; //IPIN -1 (7,9) #36
wire n7194; //IPIN -1 (7,9) #37
wire n7195; //IPIN -1 (7,9) #38
wire n7196; //IPIN -1 (7,9) #39
wire n7197; //IPIN -1 (7,9) #40
wire n7198; //IPIN -1 (7,9) #41
wire n7199; //IPIN -1 (7,9) #42
wire n7200; //IPIN -1 (7,9) #43
wire n7201; //IPIN -1 (7,9) #44
wire n7202; //IPIN -1 (7,9) #45
wire n7203; //IPIN -1 (7,9) #46
wire n7204; //IPIN -1 (7,9) #47
wire n7205; //IPIN -1 (7,9) #48
wire n7206; //IPIN -1 (7,9) #49
wire n7207; //IPIN -1 (7,9) #50
wire n7208; //IPIN -1 (7,9) #51
wire n7209; //OPIN -1 (7,9) #52
wire n7210; //OPIN -1 (7,9) #53
wire n7211; //OPIN -1 (7,9) #54
wire n7212; //OPIN -1 (7,9) #55
wire n7213; //OPIN -1 (7,9) #56
wire n7214; //OPIN -1 (7,9) #57
wire n7215; //OPIN -1 (7,9) #58
wire n7216; //OPIN -1 (7,9) #59
wire n7217; //OPIN -1 (7,9) #60
wire n7218; //OPIN -1 (7,9) #61
wire n7219; //OPIN -1 (7,9) #62
wire n7220; //OPIN -1 (7,9) #63
wire n7221; //OPIN -1 (7,9) #64
wire n7222; //OPIN -1 (7,9) #65
wire n7223; //OPIN -1 (7,9) #66
wire n7224; //OPIN -1 (7,9) #67
wire n7225; //OPIN -1 (7,9) #68
wire n7226; //OPIN -1 (7,9) #69
wire n7227; //OPIN -1 (7,9) #70
wire n7228; //OPIN -1 (7,9) #71
wire n7229; //IPIN -1 (7,9) #72
wire n7254; //IPIN -1 (7,10) #0
wire n7255; //OPIN -1 (7,10) #1
wire n7256; //IPIN -1 (7,10) #2
wire n7257; //IPIN -1 (7,10) #3
wire n7258; //OPIN -1 (7,10) #4
wire n7259; //IPIN -1 (7,10) #5
wire n7260; //IPIN -1 (7,10) #6
wire n7261; //OPIN -1 (7,10) #7
wire n7262; //IPIN -1 (7,10) #8
wire n7263; //IPIN -1 (7,10) #9
wire n7264; //OPIN -1 (7,10) #10
wire n7265; //IPIN -1 (7,10) #11
wire n7266; //IPIN -1 (7,10) #12
wire n7267; //OPIN -1 (7,10) #13
wire n7268; //IPIN -1 (7,10) #14
wire n7269; //IPIN -1 (7,10) #15
wire n7270; //OPIN -1 (7,10) #16
wire n7271; //IPIN -1 (7,10) #17
wire n7272; //IPIN -1 (7,10) #18
wire n7273; //OPIN -1 (7,10) #19
wire n7274; //IPIN -1 (7,10) #20
wire n7275; //IPIN -1 (7,10) #21
wire n7276; //OPIN -1 (7,10) #22
wire n7277; //IPIN -1 (7,10) #23
wire n7302; //IPIN -1 (8,0) #0
wire n7303; //OPIN -1 (8,0) #1
wire n7304; //IPIN -1 (8,0) #2
wire n7305; //IPIN -1 (8,0) #3
wire n7306; //OPIN -1 (8,0) #4
wire n7307; //IPIN -1 (8,0) #5
wire n7308; //IPIN -1 (8,0) #6
wire n7309; //OPIN -1 (8,0) #7
wire n7310; //IPIN -1 (8,0) #8
wire n7311; //IPIN -1 (8,0) #9
wire n7312; //OPIN -1 (8,0) #10
wire n7313; //IPIN -1 (8,0) #11
wire n7314; //IPIN -1 (8,0) #12
wire n7315; //OPIN -1 (8,0) #13
wire n7316; //IPIN -1 (8,0) #14
wire n7317; //IPIN -1 (8,0) #15
wire n7318; //OPIN -1 (8,0) #16
wire n7319; //IPIN -1 (8,0) #17
wire n7320; //IPIN -1 (8,0) #18
wire n7321; //OPIN -1 (8,0) #19
wire n7322; //IPIN -1 (8,0) #20
wire n7323; //IPIN -1 (8,0) #21
wire n7324; //OPIN -1 (8,0) #22
wire n7325; //IPIN -1 (8,0) #23
wire n7351; //IPIN -1 (8,1) #0
wire n7352; //IPIN -1 (8,1) #1
wire n7353; //IPIN -1 (8,1) #2
wire n7354; //IPIN -1 (8,1) #3
wire n7355; //IPIN -1 (8,1) #4
wire n7356; //IPIN -1 (8,1) #5
wire n7357; //IPIN -1 (8,1) #6
wire n7358; //IPIN -1 (8,1) #7
wire n7359; //IPIN -1 (8,1) #8
wire n7360; //IPIN -1 (8,1) #9
wire n7361; //IPIN -1 (8,1) #10
wire n7362; //IPIN -1 (8,1) #11
wire n7363; //IPIN -1 (8,1) #12
wire n7364; //IPIN -1 (8,1) #13
wire n7365; //IPIN -1 (8,1) #14
wire n7366; //IPIN -1 (8,1) #15
wire n7367; //IPIN -1 (8,1) #16
wire n7368; //IPIN -1 (8,1) #17
wire n7369; //IPIN -1 (8,1) #18
wire n7370; //IPIN -1 (8,1) #19
wire n7371; //IPIN -1 (8,1) #20
wire n7372; //IPIN -1 (8,1) #21
wire n7373; //IPIN -1 (8,1) #22
wire n7374; //IPIN -1 (8,1) #23
wire n7375; //IPIN -1 (8,1) #24
wire n7376; //IPIN -1 (8,1) #25
wire n7377; //IPIN -1 (8,1) #26
wire n7378; //IPIN -1 (8,1) #27
wire n7379; //IPIN -1 (8,1) #28
wire n7380; //IPIN -1 (8,1) #29
wire n7381; //IPIN -1 (8,1) #30
wire n7382; //IPIN -1 (8,1) #31
wire n7383; //IPIN -1 (8,1) #32
wire n7384; //IPIN -1 (8,1) #33
wire n7385; //IPIN -1 (8,1) #34
wire n7386; //IPIN -1 (8,1) #35
wire n7387; //IPIN -1 (8,1) #36
wire n7388; //IPIN -1 (8,1) #37
wire n7389; //IPIN -1 (8,1) #38
wire n7390; //IPIN -1 (8,1) #39
wire n7391; //IPIN -1 (8,1) #40
wire n7392; //IPIN -1 (8,1) #41
wire n7393; //IPIN -1 (8,1) #42
wire n7394; //IPIN -1 (8,1) #43
wire n7395; //IPIN -1 (8,1) #44
wire n7396; //IPIN -1 (8,1) #45
wire n7397; //IPIN -1 (8,1) #46
wire n7398; //IPIN -1 (8,1) #47
wire n7399; //IPIN -1 (8,1) #48
wire n7400; //IPIN -1 (8,1) #49
wire n7401; //IPIN -1 (8,1) #50
wire n7402; //IPIN -1 (8,1) #51
wire n7403; //OPIN -1 (8,1) #52
wire n7404; //OPIN -1 (8,1) #53
wire n7405; //OPIN -1 (8,1) #54
wire n7406; //OPIN -1 (8,1) #55
wire n7407; //OPIN -1 (8,1) #56
wire n7408; //OPIN -1 (8,1) #57
wire n7409; //OPIN -1 (8,1) #58
wire n7410; //OPIN -1 (8,1) #59
wire n7411; //OPIN -1 (8,1) #60
wire n7412; //OPIN -1 (8,1) #61
wire n7413; //OPIN -1 (8,1) #62
wire n7414; //OPIN -1 (8,1) #63
wire n7415; //OPIN -1 (8,1) #64
wire n7416; //OPIN -1 (8,1) #65
wire n7417; //OPIN -1 (8,1) #66
wire n7418; //OPIN -1 (8,1) #67
wire n7419; //OPIN -1 (8,1) #68
wire n7420; //OPIN -1 (8,1) #69
wire n7421; //OPIN -1 (8,1) #70
wire n7422; //OPIN -1 (8,1) #71
wire n7423; //IPIN -1 (8,1) #72
wire n7449; //IPIN -1 (8,2) #0
wire n7450; //IPIN -1 (8,2) #1
wire n7451; //IPIN -1 (8,2) #2
wire n7452; //IPIN -1 (8,2) #3
wire n7453; //IPIN -1 (8,2) #4
wire n7454; //IPIN -1 (8,2) #5
wire n7455; //IPIN -1 (8,2) #6
wire n7456; //IPIN -1 (8,2) #7
wire n7457; //IPIN -1 (8,2) #8
wire n7458; //IPIN -1 (8,2) #9
wire n7459; //IPIN -1 (8,2) #10
wire n7460; //IPIN -1 (8,2) #11
wire n7461; //IPIN -1 (8,2) #12
wire n7462; //IPIN -1 (8,2) #13
wire n7463; //IPIN -1 (8,2) #14
wire n7464; //IPIN -1 (8,2) #15
wire n7465; //IPIN -1 (8,2) #16
wire n7466; //IPIN -1 (8,2) #17
wire n7467; //IPIN -1 (8,2) #18
wire n7468; //IPIN -1 (8,2) #19
wire n7469; //IPIN -1 (8,2) #20
wire n7470; //IPIN -1 (8,2) #21
wire n7471; //IPIN -1 (8,2) #22
wire n7472; //IPIN -1 (8,2) #23
wire n7473; //IPIN -1 (8,2) #24
wire n7474; //IPIN -1 (8,2) #25
wire n7475; //IPIN -1 (8,2) #26
wire n7476; //IPIN -1 (8,2) #27
wire n7477; //IPIN -1 (8,2) #28
wire n7478; //IPIN -1 (8,2) #29
wire n7479; //IPIN -1 (8,2) #30
wire n7480; //IPIN -1 (8,2) #31
wire n7481; //IPIN -1 (8,2) #32
wire n7482; //IPIN -1 (8,2) #33
wire n7483; //IPIN -1 (8,2) #34
wire n7484; //IPIN -1 (8,2) #35
wire n7485; //IPIN -1 (8,2) #36
wire n7486; //IPIN -1 (8,2) #37
wire n7487; //IPIN -1 (8,2) #38
wire n7488; //IPIN -1 (8,2) #39
wire n7489; //IPIN -1 (8,2) #40
wire n7490; //IPIN -1 (8,2) #41
wire n7491; //IPIN -1 (8,2) #42
wire n7492; //IPIN -1 (8,2) #43
wire n7493; //IPIN -1 (8,2) #44
wire n7494; //IPIN -1 (8,2) #45
wire n7495; //IPIN -1 (8,2) #46
wire n7496; //IPIN -1 (8,2) #47
wire n7497; //IPIN -1 (8,2) #48
wire n7498; //IPIN -1 (8,2) #49
wire n7499; //IPIN -1 (8,2) #50
wire n7500; //IPIN -1 (8,2) #51
wire n7501; //OPIN -1 (8,2) #52
wire n7502; //OPIN -1 (8,2) #53
wire n7503; //OPIN -1 (8,2) #54
wire n7504; //OPIN -1 (8,2) #55
wire n7505; //OPIN -1 (8,2) #56
wire n7506; //OPIN -1 (8,2) #57
wire n7507; //OPIN -1 (8,2) #58
wire n7508; //OPIN -1 (8,2) #59
wire n7509; //OPIN -1 (8,2) #60
wire n7510; //OPIN -1 (8,2) #61
wire n7511; //OPIN -1 (8,2) #62
wire n7512; //OPIN -1 (8,2) #63
wire n7513; //OPIN -1 (8,2) #64
wire n7514; //OPIN -1 (8,2) #65
wire n7515; //OPIN -1 (8,2) #66
wire n7516; //OPIN -1 (8,2) #67
wire n7517; //OPIN -1 (8,2) #68
wire n7518; //OPIN -1 (8,2) #69
wire n7519; //OPIN -1 (8,2) #70
wire n7520; //OPIN -1 (8,2) #71
wire n7521; //IPIN -1 (8,2) #72
wire n7547; //IPIN -1 (8,3) #0
wire n7548; //IPIN -1 (8,3) #1
wire n7549; //IPIN -1 (8,3) #2
wire n7550; //IPIN -1 (8,3) #3
wire n7551; //IPIN -1 (8,3) #4
wire n7552; //IPIN -1 (8,3) #5
wire n7553; //IPIN -1 (8,3) #6
wire n7554; //IPIN -1 (8,3) #7
wire n7555; //IPIN -1 (8,3) #8
wire n7556; //IPIN -1 (8,3) #9
wire n7557; //IPIN -1 (8,3) #10
wire n7558; //IPIN -1 (8,3) #11
wire n7559; //IPIN -1 (8,3) #12
wire n7560; //IPIN -1 (8,3) #13
wire n7561; //IPIN -1 (8,3) #14
wire n7562; //IPIN -1 (8,3) #15
wire n7563; //IPIN -1 (8,3) #16
wire n7564; //IPIN -1 (8,3) #17
wire n7565; //IPIN -1 (8,3) #18
wire n7566; //IPIN -1 (8,3) #19
wire n7567; //IPIN -1 (8,3) #20
wire n7568; //IPIN -1 (8,3) #21
wire n7569; //IPIN -1 (8,3) #22
wire n7570; //IPIN -1 (8,3) #23
wire n7571; //IPIN -1 (8,3) #24
wire n7572; //IPIN -1 (8,3) #25
wire n7573; //IPIN -1 (8,3) #26
wire n7574; //IPIN -1 (8,3) #27
wire n7575; //IPIN -1 (8,3) #28
wire n7576; //IPIN -1 (8,3) #29
wire n7577; //IPIN -1 (8,3) #30
wire n7578; //IPIN -1 (8,3) #31
wire n7579; //IPIN -1 (8,3) #32
wire n7580; //IPIN -1 (8,3) #33
wire n7581; //IPIN -1 (8,3) #34
wire n7582; //IPIN -1 (8,3) #35
wire n7583; //IPIN -1 (8,3) #36
wire n7584; //IPIN -1 (8,3) #37
wire n7585; //IPIN -1 (8,3) #38
wire n7586; //IPIN -1 (8,3) #39
wire n7587; //IPIN -1 (8,3) #40
wire n7588; //IPIN -1 (8,3) #41
wire n7589; //IPIN -1 (8,3) #42
wire n7590; //IPIN -1 (8,3) #43
wire n7591; //IPIN -1 (8,3) #44
wire n7592; //IPIN -1 (8,3) #45
wire n7593; //IPIN -1 (8,3) #46
wire n7594; //IPIN -1 (8,3) #47
wire n7595; //IPIN -1 (8,3) #48
wire n7596; //IPIN -1 (8,3) #49
wire n7597; //IPIN -1 (8,3) #50
wire n7598; //IPIN -1 (8,3) #51
wire n7599; //OPIN -1 (8,3) #52
wire n7600; //OPIN -1 (8,3) #53
wire n7601; //OPIN -1 (8,3) #54
wire n7602; //OPIN -1 (8,3) #55
wire n7603; //OPIN -1 (8,3) #56
wire n7604; //OPIN -1 (8,3) #57
wire n7605; //OPIN -1 (8,3) #58
wire n7606; //OPIN -1 (8,3) #59
wire n7607; //OPIN -1 (8,3) #60
wire n7608; //OPIN -1 (8,3) #61
wire n7609; //OPIN -1 (8,3) #62
wire n7610; //OPIN -1 (8,3) #63
wire n7611; //OPIN -1 (8,3) #64
wire n7612; //OPIN -1 (8,3) #65
wire n7613; //OPIN -1 (8,3) #66
wire n7614; //OPIN -1 (8,3) #67
wire n7615; //OPIN -1 (8,3) #68
wire n7616; //OPIN -1 (8,3) #69
wire n7617; //OPIN -1 (8,3) #70
wire n7618; //OPIN -1 (8,3) #71
wire n7619; //IPIN -1 (8,3) #72
wire n7645; //IPIN -1 (8,4) #0
wire n7646; //IPIN -1 (8,4) #1
wire n7647; //IPIN -1 (8,4) #2
wire n7648; //IPIN -1 (8,4) #3
wire n7649; //IPIN -1 (8,4) #4
wire n7650; //IPIN -1 (8,4) #5
wire n7651; //IPIN -1 (8,4) #6
wire n7652; //IPIN -1 (8,4) #7
wire n7653; //IPIN -1 (8,4) #8
wire n7654; //IPIN -1 (8,4) #9
wire n7655; //IPIN -1 (8,4) #10
wire n7656; //IPIN -1 (8,4) #11
wire n7657; //IPIN -1 (8,4) #12
wire n7658; //IPIN -1 (8,4) #13
wire n7659; //IPIN -1 (8,4) #14
wire n7660; //IPIN -1 (8,4) #15
wire n7661; //IPIN -1 (8,4) #16
wire n7662; //IPIN -1 (8,4) #17
wire n7663; //IPIN -1 (8,4) #18
wire n7664; //IPIN -1 (8,4) #19
wire n7665; //IPIN -1 (8,4) #20
wire n7666; //IPIN -1 (8,4) #21
wire n7667; //IPIN -1 (8,4) #22
wire n7668; //IPIN -1 (8,4) #23
wire n7669; //IPIN -1 (8,4) #24
wire n7670; //IPIN -1 (8,4) #25
wire n7671; //IPIN -1 (8,4) #26
wire n7672; //IPIN -1 (8,4) #27
wire n7673; //IPIN -1 (8,4) #28
wire n7674; //IPIN -1 (8,4) #29
wire n7675; //IPIN -1 (8,4) #30
wire n7676; //IPIN -1 (8,4) #31
wire n7677; //IPIN -1 (8,4) #32
wire n7678; //IPIN -1 (8,4) #33
wire n7679; //IPIN -1 (8,4) #34
wire n7680; //IPIN -1 (8,4) #35
wire n7681; //IPIN -1 (8,4) #36
wire n7682; //IPIN -1 (8,4) #37
wire n7683; //IPIN -1 (8,4) #38
wire n7684; //IPIN -1 (8,4) #39
wire n7685; //IPIN -1 (8,4) #40
wire n7686; //IPIN -1 (8,4) #41
wire n7687; //IPIN -1 (8,4) #42
wire n7688; //IPIN -1 (8,4) #43
wire n7689; //IPIN -1 (8,4) #44
wire n7690; //IPIN -1 (8,4) #45
wire n7691; //IPIN -1 (8,4) #46
wire n7692; //IPIN -1 (8,4) #47
wire n7693; //IPIN -1 (8,4) #48
wire n7694; //IPIN -1 (8,4) #49
wire n7695; //IPIN -1 (8,4) #50
wire n7696; //IPIN -1 (8,4) #51
wire n7697; //OPIN -1 (8,4) #52
wire n7698; //OPIN -1 (8,4) #53
wire n7699; //OPIN -1 (8,4) #54
wire n7700; //OPIN -1 (8,4) #55
wire n7701; //OPIN -1 (8,4) #56
wire n7702; //OPIN -1 (8,4) #57
wire n7703; //OPIN -1 (8,4) #58
wire n7704; //OPIN -1 (8,4) #59
wire n7705; //OPIN -1 (8,4) #60
wire n7706; //OPIN -1 (8,4) #61
wire n7707; //OPIN -1 (8,4) #62
wire n7708; //OPIN -1 (8,4) #63
wire n7709; //OPIN -1 (8,4) #64
wire n7710; //OPIN -1 (8,4) #65
wire n7711; //OPIN -1 (8,4) #66
wire n7712; //OPIN -1 (8,4) #67
wire n7713; //OPIN -1 (8,4) #68
wire n7714; //OPIN -1 (8,4) #69
wire n7715; //OPIN -1 (8,4) #70
wire n7716; //OPIN -1 (8,4) #71
wire n7717; //IPIN -1 (8,4) #72
wire n7743; //IPIN -1 (8,5) #0
wire n7744; //IPIN -1 (8,5) #1
wire n7745; //IPIN -1 (8,5) #2
wire n7746; //IPIN -1 (8,5) #3
wire n7747; //IPIN -1 (8,5) #4
wire n7748; //IPIN -1 (8,5) #5
wire n7749; //IPIN -1 (8,5) #6
wire n7750; //IPIN -1 (8,5) #7
wire n7751; //IPIN -1 (8,5) #8
wire n7752; //IPIN -1 (8,5) #9
wire n7753; //IPIN -1 (8,5) #10
wire n7754; //IPIN -1 (8,5) #11
wire n7755; //IPIN -1 (8,5) #12
wire n7756; //IPIN -1 (8,5) #13
wire n7757; //IPIN -1 (8,5) #14
wire n7758; //IPIN -1 (8,5) #15
wire n7759; //IPIN -1 (8,5) #16
wire n7760; //IPIN -1 (8,5) #17
wire n7761; //IPIN -1 (8,5) #18
wire n7762; //IPIN -1 (8,5) #19
wire n7763; //IPIN -1 (8,5) #20
wire n7764; //IPIN -1 (8,5) #21
wire n7765; //IPIN -1 (8,5) #22
wire n7766; //IPIN -1 (8,5) #23
wire n7767; //IPIN -1 (8,5) #24
wire n7768; //IPIN -1 (8,5) #25
wire n7769; //IPIN -1 (8,5) #26
wire n7770; //IPIN -1 (8,5) #27
wire n7771; //IPIN -1 (8,5) #28
wire n7772; //IPIN -1 (8,5) #29
wire n7773; //IPIN -1 (8,5) #30
wire n7774; //IPIN -1 (8,5) #31
wire n7775; //IPIN -1 (8,5) #32
wire n7776; //IPIN -1 (8,5) #33
wire n7777; //IPIN -1 (8,5) #34
wire n7778; //IPIN -1 (8,5) #35
wire n7779; //IPIN -1 (8,5) #36
wire n7780; //IPIN -1 (8,5) #37
wire n7781; //IPIN -1 (8,5) #38
wire n7782; //IPIN -1 (8,5) #39
wire n7783; //IPIN -1 (8,5) #40
wire n7784; //IPIN -1 (8,5) #41
wire n7785; //IPIN -1 (8,5) #42
wire n7786; //IPIN -1 (8,5) #43
wire n7787; //IPIN -1 (8,5) #44
wire n7788; //IPIN -1 (8,5) #45
wire n7789; //IPIN -1 (8,5) #46
wire n7790; //IPIN -1 (8,5) #47
wire n7791; //IPIN -1 (8,5) #48
wire n7792; //IPIN -1 (8,5) #49
wire n7793; //IPIN -1 (8,5) #50
wire n7794; //IPIN -1 (8,5) #51
wire n7795; //OPIN -1 (8,5) #52
wire n7796; //OPIN -1 (8,5) #53
wire n7797; //OPIN -1 (8,5) #54
wire n7798; //OPIN -1 (8,5) #55
wire n7799; //OPIN -1 (8,5) #56
wire n7800; //OPIN -1 (8,5) #57
wire n7801; //OPIN -1 (8,5) #58
wire n7802; //OPIN -1 (8,5) #59
wire n7803; //OPIN -1 (8,5) #60
wire n7804; //OPIN -1 (8,5) #61
wire n7805; //OPIN -1 (8,5) #62
wire n7806; //OPIN -1 (8,5) #63
wire n7807; //OPIN -1 (8,5) #64
wire n7808; //OPIN -1 (8,5) #65
wire n7809; //OPIN -1 (8,5) #66
wire n7810; //OPIN -1 (8,5) #67
wire n7811; //OPIN -1 (8,5) #68
wire n7812; //OPIN -1 (8,5) #69
wire n7813; //OPIN -1 (8,5) #70
wire n7814; //OPIN -1 (8,5) #71
wire n7815; //IPIN -1 (8,5) #72
wire n7841; //IPIN -1 (8,6) #0
wire n7842; //IPIN -1 (8,6) #1
wire n7843; //IPIN -1 (8,6) #2
wire n7844; //IPIN -1 (8,6) #3
wire n7845; //IPIN -1 (8,6) #4
wire n7846; //IPIN -1 (8,6) #5
wire n7847; //IPIN -1 (8,6) #6
wire n7848; //IPIN -1 (8,6) #7
wire n7849; //IPIN -1 (8,6) #8
wire n7850; //IPIN -1 (8,6) #9
wire n7851; //IPIN -1 (8,6) #10
wire n7852; //IPIN -1 (8,6) #11
wire n7853; //IPIN -1 (8,6) #12
wire n7854; //IPIN -1 (8,6) #13
wire n7855; //IPIN -1 (8,6) #14
wire n7856; //IPIN -1 (8,6) #15
wire n7857; //IPIN -1 (8,6) #16
wire n7858; //IPIN -1 (8,6) #17
wire n7859; //IPIN -1 (8,6) #18
wire n7860; //IPIN -1 (8,6) #19
wire n7861; //IPIN -1 (8,6) #20
wire n7862; //IPIN -1 (8,6) #21
wire n7863; //IPIN -1 (8,6) #22
wire n7864; //IPIN -1 (8,6) #23
wire n7865; //IPIN -1 (8,6) #24
wire n7866; //IPIN -1 (8,6) #25
wire n7867; //IPIN -1 (8,6) #26
wire n7868; //IPIN -1 (8,6) #27
wire n7869; //IPIN -1 (8,6) #28
wire n7870; //IPIN -1 (8,6) #29
wire n7871; //IPIN -1 (8,6) #30
wire n7872; //IPIN -1 (8,6) #31
wire n7873; //IPIN -1 (8,6) #32
wire n7874; //IPIN -1 (8,6) #33
wire n7875; //IPIN -1 (8,6) #34
wire n7876; //IPIN -1 (8,6) #35
wire n7877; //IPIN -1 (8,6) #36
wire n7878; //IPIN -1 (8,6) #37
wire n7879; //IPIN -1 (8,6) #38
wire n7880; //IPIN -1 (8,6) #39
wire n7881; //IPIN -1 (8,6) #40
wire n7882; //IPIN -1 (8,6) #41
wire n7883; //IPIN -1 (8,6) #42
wire n7884; //IPIN -1 (8,6) #43
wire n7885; //IPIN -1 (8,6) #44
wire n7886; //IPIN -1 (8,6) #45
wire n7887; //IPIN -1 (8,6) #46
wire n7888; //IPIN -1 (8,6) #47
wire n7889; //IPIN -1 (8,6) #48
wire n7890; //IPIN -1 (8,6) #49
wire n7891; //IPIN -1 (8,6) #50
wire n7892; //IPIN -1 (8,6) #51
wire n7893; //OPIN -1 (8,6) #52
wire n7894; //OPIN -1 (8,6) #53
wire n7895; //OPIN -1 (8,6) #54
wire n7896; //OPIN -1 (8,6) #55
wire n7897; //OPIN -1 (8,6) #56
wire n7898; //OPIN -1 (8,6) #57
wire n7899; //OPIN -1 (8,6) #58
wire n7900; //OPIN -1 (8,6) #59
wire n7901; //OPIN -1 (8,6) #60
wire n7902; //OPIN -1 (8,6) #61
wire n7903; //OPIN -1 (8,6) #62
wire n7904; //OPIN -1 (8,6) #63
wire n7905; //OPIN -1 (8,6) #64
wire n7906; //OPIN -1 (8,6) #65
wire n7907; //OPIN -1 (8,6) #66
wire n7908; //OPIN -1 (8,6) #67
wire n7909; //OPIN -1 (8,6) #68
wire n7910; //OPIN -1 (8,6) #69
wire n7911; //OPIN -1 (8,6) #70
wire n7912; //OPIN -1 (8,6) #71
wire n7913; //IPIN -1 (8,6) #72
wire n7939; //IPIN -1 (8,7) #0
wire n7940; //IPIN -1 (8,7) #1
wire n7941; //IPIN -1 (8,7) #2
wire n7942; //IPIN -1 (8,7) #3
wire n7943; //IPIN -1 (8,7) #4
wire n7944; //IPIN -1 (8,7) #5
wire n7945; //IPIN -1 (8,7) #6
wire n7946; //IPIN -1 (8,7) #7
wire n7947; //IPIN -1 (8,7) #8
wire n7948; //IPIN -1 (8,7) #9
wire n7949; //IPIN -1 (8,7) #10
wire n7950; //IPIN -1 (8,7) #11
wire n7951; //IPIN -1 (8,7) #12
wire n7952; //IPIN -1 (8,7) #13
wire n7953; //IPIN -1 (8,7) #14
wire n7954; //IPIN -1 (8,7) #15
wire n7955; //IPIN -1 (8,7) #16
wire n7956; //IPIN -1 (8,7) #17
wire n7957; //IPIN -1 (8,7) #18
wire n7958; //IPIN -1 (8,7) #19
wire n7959; //IPIN -1 (8,7) #20
wire n7960; //IPIN -1 (8,7) #21
wire n7961; //IPIN -1 (8,7) #22
wire n7962; //IPIN -1 (8,7) #23
wire n7963; //IPIN -1 (8,7) #24
wire n7964; //IPIN -1 (8,7) #25
wire n7965; //IPIN -1 (8,7) #26
wire n7966; //IPIN -1 (8,7) #27
wire n7967; //IPIN -1 (8,7) #28
wire n7968; //IPIN -1 (8,7) #29
wire n7969; //IPIN -1 (8,7) #30
wire n7970; //IPIN -1 (8,7) #31
wire n7971; //IPIN -1 (8,7) #32
wire n7972; //IPIN -1 (8,7) #33
wire n7973; //IPIN -1 (8,7) #34
wire n7974; //IPIN -1 (8,7) #35
wire n7975; //IPIN -1 (8,7) #36
wire n7976; //IPIN -1 (8,7) #37
wire n7977; //IPIN -1 (8,7) #38
wire n7978; //IPIN -1 (8,7) #39
wire n7979; //IPIN -1 (8,7) #40
wire n7980; //IPIN -1 (8,7) #41
wire n7981; //IPIN -1 (8,7) #42
wire n7982; //IPIN -1 (8,7) #43
wire n7983; //IPIN -1 (8,7) #44
wire n7984; //IPIN -1 (8,7) #45
wire n7985; //IPIN -1 (8,7) #46
wire n7986; //IPIN -1 (8,7) #47
wire n7987; //IPIN -1 (8,7) #48
wire n7988; //IPIN -1 (8,7) #49
wire n7989; //IPIN -1 (8,7) #50
wire n7990; //IPIN -1 (8,7) #51
wire n7991; //OPIN -1 (8,7) #52
wire n7992; //OPIN -1 (8,7) #53
wire n7993; //OPIN -1 (8,7) #54
wire n7994; //OPIN -1 (8,7) #55
wire n7995; //OPIN -1 (8,7) #56
wire n7996; //OPIN -1 (8,7) #57
wire n7997; //OPIN -1 (8,7) #58
wire n7998; //OPIN -1 (8,7) #59
wire n7999; //OPIN -1 (8,7) #60
wire n8000; //OPIN -1 (8,7) #61
wire n8001; //OPIN -1 (8,7) #62
wire n8002; //OPIN -1 (8,7) #63
wire n8003; //OPIN -1 (8,7) #64
wire n8004; //OPIN -1 (8,7) #65
wire n8005; //OPIN -1 (8,7) #66
wire n8006; //OPIN -1 (8,7) #67
wire n8007; //OPIN -1 (8,7) #68
wire n8008; //OPIN -1 (8,7) #69
wire n8009; //OPIN -1 (8,7) #70
wire n8010; //OPIN -1 (8,7) #71
wire n8011; //IPIN -1 (8,7) #72
wire n8037; //IPIN -1 (8,8) #0
wire n8038; //IPIN -1 (8,8) #1
wire n8039; //IPIN -1 (8,8) #2
wire n8040; //IPIN -1 (8,8) #3
wire n8041; //IPIN -1 (8,8) #4
wire n8042; //IPIN -1 (8,8) #5
wire n8043; //IPIN -1 (8,8) #6
wire n8044; //IPIN -1 (8,8) #7
wire n8045; //IPIN -1 (8,8) #8
wire n8046; //IPIN -1 (8,8) #9
wire n8047; //IPIN -1 (8,8) #10
wire n8048; //IPIN -1 (8,8) #11
wire n8049; //IPIN -1 (8,8) #12
wire n8050; //IPIN -1 (8,8) #13
wire n8051; //IPIN -1 (8,8) #14
wire n8052; //IPIN -1 (8,8) #15
wire n8053; //IPIN -1 (8,8) #16
wire n8054; //IPIN -1 (8,8) #17
wire n8055; //IPIN -1 (8,8) #18
wire n8056; //IPIN -1 (8,8) #19
wire n8057; //IPIN -1 (8,8) #20
wire n8058; //IPIN -1 (8,8) #21
wire n8059; //IPIN -1 (8,8) #22
wire n8060; //IPIN -1 (8,8) #23
wire n8061; //IPIN -1 (8,8) #24
wire n8062; //IPIN -1 (8,8) #25
wire n8063; //IPIN -1 (8,8) #26
wire n8064; //IPIN -1 (8,8) #27
wire n8065; //IPIN -1 (8,8) #28
wire n8066; //IPIN -1 (8,8) #29
wire n8067; //IPIN -1 (8,8) #30
wire n8068; //IPIN -1 (8,8) #31
wire n8069; //IPIN -1 (8,8) #32
wire n8070; //IPIN -1 (8,8) #33
wire n8071; //IPIN -1 (8,8) #34
wire n8072; //IPIN -1 (8,8) #35
wire n8073; //IPIN -1 (8,8) #36
wire n8074; //IPIN -1 (8,8) #37
wire n8075; //IPIN -1 (8,8) #38
wire n8076; //IPIN -1 (8,8) #39
wire n8077; //IPIN -1 (8,8) #40
wire n8078; //IPIN -1 (8,8) #41
wire n8079; //IPIN -1 (8,8) #42
wire n8080; //IPIN -1 (8,8) #43
wire n8081; //IPIN -1 (8,8) #44
wire n8082; //IPIN -1 (8,8) #45
wire n8083; //IPIN -1 (8,8) #46
wire n8084; //IPIN -1 (8,8) #47
wire n8085; //IPIN -1 (8,8) #48
wire n8086; //IPIN -1 (8,8) #49
wire n8087; //IPIN -1 (8,8) #50
wire n8088; //IPIN -1 (8,8) #51
wire n8089; //OPIN -1 (8,8) #52
wire n8090; //OPIN -1 (8,8) #53
wire n8091; //OPIN -1 (8,8) #54
wire n8092; //OPIN -1 (8,8) #55
wire n8093; //OPIN -1 (8,8) #56
wire n8094; //OPIN -1 (8,8) #57
wire n8095; //OPIN -1 (8,8) #58
wire n8096; //OPIN -1 (8,8) #59
wire n8097; //OPIN -1 (8,8) #60
wire n8098; //OPIN -1 (8,8) #61
wire n8099; //OPIN -1 (8,8) #62
wire n8100; //OPIN -1 (8,8) #63
wire n8101; //OPIN -1 (8,8) #64
wire n8102; //OPIN -1 (8,8) #65
wire n8103; //OPIN -1 (8,8) #66
wire n8104; //OPIN -1 (8,8) #67
wire n8105; //OPIN -1 (8,8) #68
wire n8106; //OPIN -1 (8,8) #69
wire n8107; //OPIN -1 (8,8) #70
wire n8108; //OPIN -1 (8,8) #71
wire n8109; //IPIN -1 (8,8) #72
wire n8135; //IPIN -1 (8,9) #0
wire n8136; //IPIN -1 (8,9) #1
wire n8137; //IPIN -1 (8,9) #2
wire n8138; //IPIN -1 (8,9) #3
wire n8139; //IPIN -1 (8,9) #4
wire n8140; //IPIN -1 (8,9) #5
wire n8141; //IPIN -1 (8,9) #6
wire n8142; //IPIN -1 (8,9) #7
wire n8143; //IPIN -1 (8,9) #8
wire n8144; //IPIN -1 (8,9) #9
wire n8145; //IPIN -1 (8,9) #10
wire n8146; //IPIN -1 (8,9) #11
wire n8147; //IPIN -1 (8,9) #12
wire n8148; //IPIN -1 (8,9) #13
wire n8149; //IPIN -1 (8,9) #14
wire n8150; //IPIN -1 (8,9) #15
wire n8151; //IPIN -1 (8,9) #16
wire n8152; //IPIN -1 (8,9) #17
wire n8153; //IPIN -1 (8,9) #18
wire n8154; //IPIN -1 (8,9) #19
wire n8155; //IPIN -1 (8,9) #20
wire n8156; //IPIN -1 (8,9) #21
wire n8157; //IPIN -1 (8,9) #22
wire n8158; //IPIN -1 (8,9) #23
wire n8159; //IPIN -1 (8,9) #24
wire n8160; //IPIN -1 (8,9) #25
wire n8161; //IPIN -1 (8,9) #26
wire n8162; //IPIN -1 (8,9) #27
wire n8163; //IPIN -1 (8,9) #28
wire n8164; //IPIN -1 (8,9) #29
wire n8165; //IPIN -1 (8,9) #30
wire n8166; //IPIN -1 (8,9) #31
wire n8167; //IPIN -1 (8,9) #32
wire n8168; //IPIN -1 (8,9) #33
wire n8169; //IPIN -1 (8,9) #34
wire n8170; //IPIN -1 (8,9) #35
wire n8171; //IPIN -1 (8,9) #36
wire n8172; //IPIN -1 (8,9) #37
wire n8173; //IPIN -1 (8,9) #38
wire n8174; //IPIN -1 (8,9) #39
wire n8175; //IPIN -1 (8,9) #40
wire n8176; //IPIN -1 (8,9) #41
wire n8177; //IPIN -1 (8,9) #42
wire n8178; //IPIN -1 (8,9) #43
wire n8179; //IPIN -1 (8,9) #44
wire n8180; //IPIN -1 (8,9) #45
wire n8181; //IPIN -1 (8,9) #46
wire n8182; //IPIN -1 (8,9) #47
wire n8183; //IPIN -1 (8,9) #48
wire n8184; //IPIN -1 (8,9) #49
wire n8185; //IPIN -1 (8,9) #50
wire n8186; //IPIN -1 (8,9) #51
wire n8187; //OPIN -1 (8,9) #52
wire n8188; //OPIN -1 (8,9) #53
wire n8189; //OPIN -1 (8,9) #54
wire n8190; //OPIN -1 (8,9) #55
wire n8191; //OPIN -1 (8,9) #56
wire n8192; //OPIN -1 (8,9) #57
wire n8193; //OPIN -1 (8,9) #58
wire n8194; //OPIN -1 (8,9) #59
wire n8195; //OPIN -1 (8,9) #60
wire n8196; //OPIN -1 (8,9) #61
wire n8197; //OPIN -1 (8,9) #62
wire n8198; //OPIN -1 (8,9) #63
wire n8199; //OPIN -1 (8,9) #64
wire n8200; //OPIN -1 (8,9) #65
wire n8201; //OPIN -1 (8,9) #66
wire n8202; //OPIN -1 (8,9) #67
wire n8203; //OPIN -1 (8,9) #68
wire n8204; //OPIN -1 (8,9) #69
wire n8205; //OPIN -1 (8,9) #70
wire n8206; //OPIN -1 (8,9) #71
wire n8207; //IPIN -1 (8,9) #72
wire n8232; //IPIN -1 (8,10) #0
wire n8233; //OPIN -1 (8,10) #1
wire n8234; //IPIN -1 (8,10) #2
wire n8235; //IPIN -1 (8,10) #3
wire n8236; //OPIN -1 (8,10) #4
wire n8237; //IPIN -1 (8,10) #5
wire n8238; //IPIN -1 (8,10) #6
wire n8239; //OPIN -1 (8,10) #7
wire n8240; //IPIN -1 (8,10) #8
wire n8241; //IPIN -1 (8,10) #9
wire n8242; //OPIN -1 (8,10) #10
wire n8243; //IPIN -1 (8,10) #11
wire n8244; //IPIN -1 (8,10) #12
wire n8245; //OPIN -1 (8,10) #13
wire n8246; //IPIN -1 (8,10) #14
wire n8247; //IPIN -1 (8,10) #15
wire n8248; //OPIN -1 (8,10) #16
wire n8249; //IPIN -1 (8,10) #17
wire n8250; //IPIN -1 (8,10) #18
wire n8251; //OPIN -1 (8,10) #19
wire n8252; //IPIN -1 (8,10) #20
wire n8253; //IPIN -1 (8,10) #21
wire n8254; //OPIN -1 (8,10) #22
wire n8255; //IPIN -1 (8,10) #23
wire n8280; //IPIN -1 (9,0) #0
wire n8281; //OPIN -1 (9,0) #1
wire n8282; //IPIN -1 (9,0) #2
wire n8283; //IPIN -1 (9,0) #3
wire n8284; //OPIN -1 (9,0) #4
wire n8285; //IPIN -1 (9,0) #5
wire n8286; //IPIN -1 (9,0) #6
wire n8287; //OPIN -1 (9,0) #7
wire n8288; //IPIN -1 (9,0) #8
wire n8289; //IPIN -1 (9,0) #9
wire n8290; //OPIN -1 (9,0) #10
wire n8291; //IPIN -1 (9,0) #11
wire n8292; //IPIN -1 (9,0) #12
wire n8293; //OPIN -1 (9,0) #13
wire n8294; //IPIN -1 (9,0) #14
wire n8295; //IPIN -1 (9,0) #15
wire n8296; //OPIN -1 (9,0) #16
wire n8297; //IPIN -1 (9,0) #17
wire n8298; //IPIN -1 (9,0) #18
wire n8299; //OPIN -1 (9,0) #19
wire n8300; //IPIN -1 (9,0) #20
wire n8301; //IPIN -1 (9,0) #21
wire n8302; //OPIN -1 (9,0) #22
wire n8303; //IPIN -1 (9,0) #23
wire n8329; //IPIN -1 (9,1) #0
wire n8330; //IPIN -1 (9,1) #1
wire n8331; //IPIN -1 (9,1) #2
wire n8332; //IPIN -1 (9,1) #3
wire n8333; //IPIN -1 (9,1) #4
wire n8334; //IPIN -1 (9,1) #5
wire n8335; //IPIN -1 (9,1) #6
wire n8336; //IPIN -1 (9,1) #7
wire n8337; //IPIN -1 (9,1) #8
wire n8338; //IPIN -1 (9,1) #9
wire n8339; //IPIN -1 (9,1) #10
wire n8340; //IPIN -1 (9,1) #11
wire n8341; //IPIN -1 (9,1) #12
wire n8342; //IPIN -1 (9,1) #13
wire n8343; //IPIN -1 (9,1) #14
wire n8344; //IPIN -1 (9,1) #15
wire n8345; //IPIN -1 (9,1) #16
wire n8346; //IPIN -1 (9,1) #17
wire n8347; //IPIN -1 (9,1) #18
wire n8348; //IPIN -1 (9,1) #19
wire n8349; //IPIN -1 (9,1) #20
wire n8350; //IPIN -1 (9,1) #21
wire n8351; //IPIN -1 (9,1) #22
wire n8352; //IPIN -1 (9,1) #23
wire n8353; //IPIN -1 (9,1) #24
wire n8354; //IPIN -1 (9,1) #25
wire n8355; //IPIN -1 (9,1) #26
wire n8356; //IPIN -1 (9,1) #27
wire n8357; //IPIN -1 (9,1) #28
wire n8358; //IPIN -1 (9,1) #29
wire n8359; //IPIN -1 (9,1) #30
wire n8360; //IPIN -1 (9,1) #31
wire n8361; //IPIN -1 (9,1) #32
wire n8362; //IPIN -1 (9,1) #33
wire n8363; //IPIN -1 (9,1) #34
wire n8364; //IPIN -1 (9,1) #35
wire n8365; //IPIN -1 (9,1) #36
wire n8366; //IPIN -1 (9,1) #37
wire n8367; //IPIN -1 (9,1) #38
wire n8368; //IPIN -1 (9,1) #39
wire n8369; //IPIN -1 (9,1) #40
wire n8370; //IPIN -1 (9,1) #41
wire n8371; //IPIN -1 (9,1) #42
wire n8372; //IPIN -1 (9,1) #43
wire n8373; //IPIN -1 (9,1) #44
wire n8374; //IPIN -1 (9,1) #45
wire n8375; //IPIN -1 (9,1) #46
wire n8376; //IPIN -1 (9,1) #47
wire n8377; //IPIN -1 (9,1) #48
wire n8378; //IPIN -1 (9,1) #49
wire n8379; //IPIN -1 (9,1) #50
wire n8380; //IPIN -1 (9,1) #51
wire n8381; //OPIN -1 (9,1) #52
wire n8382; //OPIN -1 (9,1) #53
wire n8383; //OPIN -1 (9,1) #54
wire n8384; //OPIN -1 (9,1) #55
wire n8385; //OPIN -1 (9,1) #56
wire n8386; //OPIN -1 (9,1) #57
wire n8387; //OPIN -1 (9,1) #58
wire n8388; //OPIN -1 (9,1) #59
wire n8389; //OPIN -1 (9,1) #60
wire n8390; //OPIN -1 (9,1) #61
wire n8391; //OPIN -1 (9,1) #62
wire n8392; //OPIN -1 (9,1) #63
wire n8393; //OPIN -1 (9,1) #64
wire n8394; //OPIN -1 (9,1) #65
wire n8395; //OPIN -1 (9,1) #66
wire n8396; //OPIN -1 (9,1) #67
wire n8397; //OPIN -1 (9,1) #68
wire n8398; //OPIN -1 (9,1) #69
wire n8399; //OPIN -1 (9,1) #70
wire n8400; //OPIN -1 (9,1) #71
wire n8401; //IPIN -1 (9,1) #72
wire n8427; //IPIN -1 (9,2) #0
wire n8428; //IPIN -1 (9,2) #1
wire n8429; //IPIN -1 (9,2) #2
wire n8430; //IPIN -1 (9,2) #3
wire n8431; //IPIN -1 (9,2) #4
wire n8432; //IPIN -1 (9,2) #5
wire n8433; //IPIN -1 (9,2) #6
wire n8434; //IPIN -1 (9,2) #7
wire n8435; //IPIN -1 (9,2) #8
wire n8436; //IPIN -1 (9,2) #9
wire n8437; //IPIN -1 (9,2) #10
wire n8438; //IPIN -1 (9,2) #11
wire n8439; //IPIN -1 (9,2) #12
wire n8440; //IPIN -1 (9,2) #13
wire n8441; //IPIN -1 (9,2) #14
wire n8442; //IPIN -1 (9,2) #15
wire n8443; //IPIN -1 (9,2) #16
wire n8444; //IPIN -1 (9,2) #17
wire n8445; //IPIN -1 (9,2) #18
wire n8446; //IPIN -1 (9,2) #19
wire n8447; //IPIN -1 (9,2) #20
wire n8448; //IPIN -1 (9,2) #21
wire n8449; //IPIN -1 (9,2) #22
wire n8450; //IPIN -1 (9,2) #23
wire n8451; //IPIN -1 (9,2) #24
wire n8452; //IPIN -1 (9,2) #25
wire n8453; //IPIN -1 (9,2) #26
wire n8454; //IPIN -1 (9,2) #27
wire n8455; //IPIN -1 (9,2) #28
wire n8456; //IPIN -1 (9,2) #29
wire n8457; //IPIN -1 (9,2) #30
wire n8458; //IPIN -1 (9,2) #31
wire n8459; //IPIN -1 (9,2) #32
wire n8460; //IPIN -1 (9,2) #33
wire n8461; //IPIN -1 (9,2) #34
wire n8462; //IPIN -1 (9,2) #35
wire n8463; //IPIN -1 (9,2) #36
wire n8464; //IPIN -1 (9,2) #37
wire n8465; //IPIN -1 (9,2) #38
wire n8466; //IPIN -1 (9,2) #39
wire n8467; //IPIN -1 (9,2) #40
wire n8468; //IPIN -1 (9,2) #41
wire n8469; //IPIN -1 (9,2) #42
wire n8470; //IPIN -1 (9,2) #43
wire n8471; //IPIN -1 (9,2) #44
wire n8472; //IPIN -1 (9,2) #45
wire n8473; //IPIN -1 (9,2) #46
wire n8474; //IPIN -1 (9,2) #47
wire n8475; //IPIN -1 (9,2) #48
wire n8476; //IPIN -1 (9,2) #49
wire n8477; //IPIN -1 (9,2) #50
wire n8478; //IPIN -1 (9,2) #51
wire n8479; //OPIN -1 (9,2) #52
wire n8480; //OPIN -1 (9,2) #53
wire n8481; //OPIN -1 (9,2) #54
wire n8482; //OPIN -1 (9,2) #55
wire n8483; //OPIN -1 (9,2) #56
wire n8484; //OPIN -1 (9,2) #57
wire n8485; //OPIN -1 (9,2) #58
wire n8486; //OPIN -1 (9,2) #59
wire n8487; //OPIN -1 (9,2) #60
wire n8488; //OPIN -1 (9,2) #61
wire n8489; //OPIN -1 (9,2) #62
wire n8490; //OPIN -1 (9,2) #63
wire n8491; //OPIN -1 (9,2) #64
wire n8492; //OPIN -1 (9,2) #65
wire n8493; //OPIN -1 (9,2) #66
wire n8494; //OPIN -1 (9,2) #67
wire n8495; //OPIN -1 (9,2) #68
wire n8496; //OPIN -1 (9,2) #69
wire n8497; //OPIN -1 (9,2) #70
wire n8498; //OPIN -1 (9,2) #71
wire n8499; //IPIN -1 (9,2) #72
wire n8525; //IPIN -1 (9,3) #0
wire n8526; //IPIN -1 (9,3) #1
wire n8527; //IPIN -1 (9,3) #2
wire n8528; //IPIN -1 (9,3) #3
wire n8529; //IPIN -1 (9,3) #4
wire n8530; //IPIN -1 (9,3) #5
wire n8531; //IPIN -1 (9,3) #6
wire n8532; //IPIN -1 (9,3) #7
wire n8533; //IPIN -1 (9,3) #8
wire n8534; //IPIN -1 (9,3) #9
wire n8535; //IPIN -1 (9,3) #10
wire n8536; //IPIN -1 (9,3) #11
wire n8537; //IPIN -1 (9,3) #12
wire n8538; //IPIN -1 (9,3) #13
wire n8539; //IPIN -1 (9,3) #14
wire n8540; //IPIN -1 (9,3) #15
wire n8541; //IPIN -1 (9,3) #16
wire n8542; //IPIN -1 (9,3) #17
wire n8543; //IPIN -1 (9,3) #18
wire n8544; //IPIN -1 (9,3) #19
wire n8545; //IPIN -1 (9,3) #20
wire n8546; //IPIN -1 (9,3) #21
wire n8547; //IPIN -1 (9,3) #22
wire n8548; //IPIN -1 (9,3) #23
wire n8549; //IPIN -1 (9,3) #24
wire n8550; //IPIN -1 (9,3) #25
wire n8551; //IPIN -1 (9,3) #26
wire n8552; //IPIN -1 (9,3) #27
wire n8553; //IPIN -1 (9,3) #28
wire n8554; //IPIN -1 (9,3) #29
wire n8555; //IPIN -1 (9,3) #30
wire n8556; //IPIN -1 (9,3) #31
wire n8557; //IPIN -1 (9,3) #32
wire n8558; //IPIN -1 (9,3) #33
wire n8559; //IPIN -1 (9,3) #34
wire n8560; //IPIN -1 (9,3) #35
wire n8561; //IPIN -1 (9,3) #36
wire n8562; //IPIN -1 (9,3) #37
wire n8563; //IPIN -1 (9,3) #38
wire n8564; //IPIN -1 (9,3) #39
wire n8565; //IPIN -1 (9,3) #40
wire n8566; //IPIN -1 (9,3) #41
wire n8567; //IPIN -1 (9,3) #42
wire n8568; //IPIN -1 (9,3) #43
wire n8569; //IPIN -1 (9,3) #44
wire n8570; //IPIN -1 (9,3) #45
wire n8571; //IPIN -1 (9,3) #46
wire n8572; //IPIN -1 (9,3) #47
wire n8573; //IPIN -1 (9,3) #48
wire n8574; //IPIN -1 (9,3) #49
wire n8575; //IPIN -1 (9,3) #50
wire n8576; //IPIN -1 (9,3) #51
wire n8577; //OPIN -1 (9,3) #52
wire n8578; //OPIN -1 (9,3) #53
wire n8579; //OPIN -1 (9,3) #54
wire n8580; //OPIN -1 (9,3) #55
wire n8581; //OPIN -1 (9,3) #56
wire n8582; //OPIN -1 (9,3) #57
wire n8583; //OPIN -1 (9,3) #58
wire n8584; //OPIN -1 (9,3) #59
wire n8585; //OPIN -1 (9,3) #60
wire n8586; //OPIN -1 (9,3) #61
wire n8587; //OPIN -1 (9,3) #62
wire n8588; //OPIN -1 (9,3) #63
wire n8589; //OPIN -1 (9,3) #64
wire n8590; //OPIN -1 (9,3) #65
wire n8591; //OPIN -1 (9,3) #66
wire n8592; //OPIN -1 (9,3) #67
wire n8593; //OPIN -1 (9,3) #68
wire n8594; //OPIN -1 (9,3) #69
wire n8595; //OPIN -1 (9,3) #70
wire n8596; //OPIN -1 (9,3) #71
wire n8597; //IPIN -1 (9,3) #72
wire n8623; //IPIN -1 (9,4) #0
wire n8624; //IPIN -1 (9,4) #1
wire n8625; //IPIN -1 (9,4) #2
wire n8626; //IPIN -1 (9,4) #3
wire n8627; //IPIN -1 (9,4) #4
wire n8628; //IPIN -1 (9,4) #5
wire n8629; //IPIN -1 (9,4) #6
wire n8630; //IPIN -1 (9,4) #7
wire n8631; //IPIN -1 (9,4) #8
wire n8632; //IPIN -1 (9,4) #9
wire n8633; //IPIN -1 (9,4) #10
wire n8634; //IPIN -1 (9,4) #11
wire n8635; //IPIN -1 (9,4) #12
wire n8636; //IPIN -1 (9,4) #13
wire n8637; //IPIN -1 (9,4) #14
wire n8638; //IPIN -1 (9,4) #15
wire n8639; //IPIN -1 (9,4) #16
wire n8640; //IPIN -1 (9,4) #17
wire n8641; //IPIN -1 (9,4) #18
wire n8642; //IPIN -1 (9,4) #19
wire n8643; //IPIN -1 (9,4) #20
wire n8644; //IPIN -1 (9,4) #21
wire n8645; //IPIN -1 (9,4) #22
wire n8646; //IPIN -1 (9,4) #23
wire n8647; //IPIN -1 (9,4) #24
wire n8648; //IPIN -1 (9,4) #25
wire n8649; //IPIN -1 (9,4) #26
wire n8650; //IPIN -1 (9,4) #27
wire n8651; //IPIN -1 (9,4) #28
wire n8652; //IPIN -1 (9,4) #29
wire n8653; //IPIN -1 (9,4) #30
wire n8654; //IPIN -1 (9,4) #31
wire n8655; //IPIN -1 (9,4) #32
wire n8656; //IPIN -1 (9,4) #33
wire n8657; //IPIN -1 (9,4) #34
wire n8658; //IPIN -1 (9,4) #35
wire n8659; //IPIN -1 (9,4) #36
wire n8660; //IPIN -1 (9,4) #37
wire n8661; //IPIN -1 (9,4) #38
wire n8662; //IPIN -1 (9,4) #39
wire n8663; //IPIN -1 (9,4) #40
wire n8664; //IPIN -1 (9,4) #41
wire n8665; //IPIN -1 (9,4) #42
wire n8666; //IPIN -1 (9,4) #43
wire n8667; //IPIN -1 (9,4) #44
wire n8668; //IPIN -1 (9,4) #45
wire n8669; //IPIN -1 (9,4) #46
wire n8670; //IPIN -1 (9,4) #47
wire n8671; //IPIN -1 (9,4) #48
wire n8672; //IPIN -1 (9,4) #49
wire n8673; //IPIN -1 (9,4) #50
wire n8674; //IPIN -1 (9,4) #51
wire n8675; //OPIN -1 (9,4) #52
wire n8676; //OPIN -1 (9,4) #53
wire n8677; //OPIN -1 (9,4) #54
wire n8678; //OPIN -1 (9,4) #55
wire n8679; //OPIN -1 (9,4) #56
wire n8680; //OPIN -1 (9,4) #57
wire n8681; //OPIN -1 (9,4) #58
wire n8682; //OPIN -1 (9,4) #59
wire n8683; //OPIN -1 (9,4) #60
wire n8684; //OPIN -1 (9,4) #61
wire n8685; //OPIN -1 (9,4) #62
wire n8686; //OPIN -1 (9,4) #63
wire n8687; //OPIN -1 (9,4) #64
wire n8688; //OPIN -1 (9,4) #65
wire n8689; //OPIN -1 (9,4) #66
wire n8690; //OPIN -1 (9,4) #67
wire n8691; //OPIN -1 (9,4) #68
wire n8692; //OPIN -1 (9,4) #69
wire n8693; //OPIN -1 (9,4) #70
wire n8694; //OPIN -1 (9,4) #71
wire n8695; //IPIN -1 (9,4) #72
wire n8721; //IPIN -1 (9,5) #0
wire n8722; //IPIN -1 (9,5) #1
wire n8723; //IPIN -1 (9,5) #2
wire n8724; //IPIN -1 (9,5) #3
wire n8725; //IPIN -1 (9,5) #4
wire n8726; //IPIN -1 (9,5) #5
wire n8727; //IPIN -1 (9,5) #6
wire n8728; //IPIN -1 (9,5) #7
wire n8729; //IPIN -1 (9,5) #8
wire n8730; //IPIN -1 (9,5) #9
wire n8731; //IPIN -1 (9,5) #10
wire n8732; //IPIN -1 (9,5) #11
wire n8733; //IPIN -1 (9,5) #12
wire n8734; //IPIN -1 (9,5) #13
wire n8735; //IPIN -1 (9,5) #14
wire n8736; //IPIN -1 (9,5) #15
wire n8737; //IPIN -1 (9,5) #16
wire n8738; //IPIN -1 (9,5) #17
wire n8739; //IPIN -1 (9,5) #18
wire n8740; //IPIN -1 (9,5) #19
wire n8741; //IPIN -1 (9,5) #20
wire n8742; //IPIN -1 (9,5) #21
wire n8743; //IPIN -1 (9,5) #22
wire n8744; //IPIN -1 (9,5) #23
wire n8745; //IPIN -1 (9,5) #24
wire n8746; //IPIN -1 (9,5) #25
wire n8747; //IPIN -1 (9,5) #26
wire n8748; //IPIN -1 (9,5) #27
wire n8749; //IPIN -1 (9,5) #28
wire n8750; //IPIN -1 (9,5) #29
wire n8751; //IPIN -1 (9,5) #30
wire n8752; //IPIN -1 (9,5) #31
wire n8753; //IPIN -1 (9,5) #32
wire n8754; //IPIN -1 (9,5) #33
wire n8755; //IPIN -1 (9,5) #34
wire n8756; //IPIN -1 (9,5) #35
wire n8757; //IPIN -1 (9,5) #36
wire n8758; //IPIN -1 (9,5) #37
wire n8759; //IPIN -1 (9,5) #38
wire n8760; //IPIN -1 (9,5) #39
wire n8761; //IPIN -1 (9,5) #40
wire n8762; //IPIN -1 (9,5) #41
wire n8763; //IPIN -1 (9,5) #42
wire n8764; //IPIN -1 (9,5) #43
wire n8765; //IPIN -1 (9,5) #44
wire n8766; //IPIN -1 (9,5) #45
wire n8767; //IPIN -1 (9,5) #46
wire n8768; //IPIN -1 (9,5) #47
wire n8769; //IPIN -1 (9,5) #48
wire n8770; //IPIN -1 (9,5) #49
wire n8771; //IPIN -1 (9,5) #50
wire n8772; //IPIN -1 (9,5) #51
wire n8773; //OPIN -1 (9,5) #52
wire n8774; //OPIN -1 (9,5) #53
wire n8775; //OPIN -1 (9,5) #54
wire n8776; //OPIN -1 (9,5) #55
wire n8777; //OPIN -1 (9,5) #56
wire n8778; //OPIN -1 (9,5) #57
wire n8779; //OPIN -1 (9,5) #58
wire n8780; //OPIN -1 (9,5) #59
wire n8781; //OPIN -1 (9,5) #60
wire n8782; //OPIN -1 (9,5) #61
wire n8783; //OPIN -1 (9,5) #62
wire n8784; //OPIN -1 (9,5) #63
wire n8785; //OPIN -1 (9,5) #64
wire n8786; //OPIN -1 (9,5) #65
wire n8787; //OPIN -1 (9,5) #66
wire n8788; //OPIN -1 (9,5) #67
wire n8789; //OPIN -1 (9,5) #68
wire n8790; //OPIN -1 (9,5) #69
wire n8791; //OPIN -1 (9,5) #70
wire n8792; //OPIN -1 (9,5) #71
wire n8793; //IPIN -1 (9,5) #72
wire n8819; //IPIN -1 (9,6) #0
wire n8820; //IPIN -1 (9,6) #1
wire n8821; //IPIN -1 (9,6) #2
wire n8822; //IPIN -1 (9,6) #3
wire n8823; //IPIN -1 (9,6) #4
wire n8824; //IPIN -1 (9,6) #5
wire n8825; //IPIN -1 (9,6) #6
wire n8826; //IPIN -1 (9,6) #7
wire n8827; //IPIN -1 (9,6) #8
wire n8828; //IPIN -1 (9,6) #9
wire n8829; //IPIN -1 (9,6) #10
wire n8830; //IPIN -1 (9,6) #11
wire n8831; //IPIN -1 (9,6) #12
wire n8832; //IPIN -1 (9,6) #13
wire n8833; //IPIN -1 (9,6) #14
wire n8834; //IPIN -1 (9,6) #15
wire n8835; //IPIN -1 (9,6) #16
wire n8836; //IPIN -1 (9,6) #17
wire n8837; //IPIN -1 (9,6) #18
wire n8838; //IPIN -1 (9,6) #19
wire n8839; //IPIN -1 (9,6) #20
wire n8840; //IPIN -1 (9,6) #21
wire n8841; //IPIN -1 (9,6) #22
wire n8842; //IPIN -1 (9,6) #23
wire n8843; //IPIN -1 (9,6) #24
wire n8844; //IPIN -1 (9,6) #25
wire n8845; //IPIN -1 (9,6) #26
wire n8846; //IPIN -1 (9,6) #27
wire n8847; //IPIN -1 (9,6) #28
wire n8848; //IPIN -1 (9,6) #29
wire n8849; //IPIN -1 (9,6) #30
wire n8850; //IPIN -1 (9,6) #31
wire n8851; //IPIN -1 (9,6) #32
wire n8852; //IPIN -1 (9,6) #33
wire n8853; //IPIN -1 (9,6) #34
wire n8854; //IPIN -1 (9,6) #35
wire n8855; //IPIN -1 (9,6) #36
wire n8856; //IPIN -1 (9,6) #37
wire n8857; //IPIN -1 (9,6) #38
wire n8858; //IPIN -1 (9,6) #39
wire n8859; //IPIN -1 (9,6) #40
wire n8860; //IPIN -1 (9,6) #41
wire n8861; //IPIN -1 (9,6) #42
wire n8862; //IPIN -1 (9,6) #43
wire n8863; //IPIN -1 (9,6) #44
wire n8864; //IPIN -1 (9,6) #45
wire n8865; //IPIN -1 (9,6) #46
wire n8866; //IPIN -1 (9,6) #47
wire n8867; //IPIN -1 (9,6) #48
wire n8868; //IPIN -1 (9,6) #49
wire n8869; //IPIN -1 (9,6) #50
wire n8870; //IPIN -1 (9,6) #51
wire n8871; //OPIN -1 (9,6) #52
wire n8872; //OPIN -1 (9,6) #53
wire n8873; //OPIN -1 (9,6) #54
wire n8874; //OPIN -1 (9,6) #55
wire n8875; //OPIN -1 (9,6) #56
wire n8876; //OPIN -1 (9,6) #57
wire n8877; //OPIN -1 (9,6) #58
wire n8878; //OPIN -1 (9,6) #59
wire n8879; //OPIN -1 (9,6) #60
wire n8880; //OPIN -1 (9,6) #61
wire n8881; //OPIN -1 (9,6) #62
wire n8882; //OPIN -1 (9,6) #63
wire n8883; //OPIN -1 (9,6) #64
wire n8884; //OPIN -1 (9,6) #65
wire n8885; //OPIN -1 (9,6) #66
wire n8886; //OPIN -1 (9,6) #67
wire n8887; //OPIN -1 (9,6) #68
wire n8888; //OPIN -1 (9,6) #69
wire n8889; //OPIN -1 (9,6) #70
wire n8890; //OPIN -1 (9,6) #71
wire n8891; //IPIN -1 (9,6) #72
wire n8917; //IPIN -1 (9,7) #0
wire n8918; //IPIN -1 (9,7) #1
wire n8919; //IPIN -1 (9,7) #2
wire n8920; //IPIN -1 (9,7) #3
wire n8921; //IPIN -1 (9,7) #4
wire n8922; //IPIN -1 (9,7) #5
wire n8923; //IPIN -1 (9,7) #6
wire n8924; //IPIN -1 (9,7) #7
wire n8925; //IPIN -1 (9,7) #8
wire n8926; //IPIN -1 (9,7) #9
wire n8927; //IPIN -1 (9,7) #10
wire n8928; //IPIN -1 (9,7) #11
wire n8929; //IPIN -1 (9,7) #12
wire n8930; //IPIN -1 (9,7) #13
wire n8931; //IPIN -1 (9,7) #14
wire n8932; //IPIN -1 (9,7) #15
wire n8933; //IPIN -1 (9,7) #16
wire n8934; //IPIN -1 (9,7) #17
wire n8935; //IPIN -1 (9,7) #18
wire n8936; //IPIN -1 (9,7) #19
wire n8937; //IPIN -1 (9,7) #20
wire n8938; //IPIN -1 (9,7) #21
wire n8939; //IPIN -1 (9,7) #22
wire n8940; //IPIN -1 (9,7) #23
wire n8941; //IPIN -1 (9,7) #24
wire n8942; //IPIN -1 (9,7) #25
wire n8943; //IPIN -1 (9,7) #26
wire n8944; //IPIN -1 (9,7) #27
wire n8945; //IPIN -1 (9,7) #28
wire n8946; //IPIN -1 (9,7) #29
wire n8947; //IPIN -1 (9,7) #30
wire n8948; //IPIN -1 (9,7) #31
wire n8949; //IPIN -1 (9,7) #32
wire n8950; //IPIN -1 (9,7) #33
wire n8951; //IPIN -1 (9,7) #34
wire n8952; //IPIN -1 (9,7) #35
wire n8953; //IPIN -1 (9,7) #36
wire n8954; //IPIN -1 (9,7) #37
wire n8955; //IPIN -1 (9,7) #38
wire n8956; //IPIN -1 (9,7) #39
wire n8957; //IPIN -1 (9,7) #40
wire n8958; //IPIN -1 (9,7) #41
wire n8959; //IPIN -1 (9,7) #42
wire n8960; //IPIN -1 (9,7) #43
wire n8961; //IPIN -1 (9,7) #44
wire n8962; //IPIN -1 (9,7) #45
wire n8963; //IPIN -1 (9,7) #46
wire n8964; //IPIN -1 (9,7) #47
wire n8965; //IPIN -1 (9,7) #48
wire n8966; //IPIN -1 (9,7) #49
wire n8967; //IPIN -1 (9,7) #50
wire n8968; //IPIN -1 (9,7) #51
wire n8969; //OPIN -1 (9,7) #52
wire n8970; //OPIN -1 (9,7) #53
wire n8971; //OPIN -1 (9,7) #54
wire n8972; //OPIN -1 (9,7) #55
wire n8973; //OPIN -1 (9,7) #56
wire n8974; //OPIN -1 (9,7) #57
wire n8975; //OPIN -1 (9,7) #58
wire n8976; //OPIN -1 (9,7) #59
wire n8977; //OPIN -1 (9,7) #60
wire n8978; //OPIN -1 (9,7) #61
wire n8979; //OPIN -1 (9,7) #62
wire n8980; //OPIN -1 (9,7) #63
wire n8981; //OPIN -1 (9,7) #64
wire n8982; //OPIN -1 (9,7) #65
wire n8983; //OPIN -1 (9,7) #66
wire n8984; //OPIN -1 (9,7) #67
wire n8985; //OPIN -1 (9,7) #68
wire n8986; //OPIN -1 (9,7) #69
wire n8987; //OPIN -1 (9,7) #70
wire n8988; //OPIN -1 (9,7) #71
wire n8989; //IPIN -1 (9,7) #72
wire n9015; //IPIN -1 (9,8) #0
wire n9016; //IPIN -1 (9,8) #1
wire n9017; //IPIN -1 (9,8) #2
wire n9018; //IPIN -1 (9,8) #3
wire n9019; //IPIN -1 (9,8) #4
wire n9020; //IPIN -1 (9,8) #5
wire n9021; //IPIN -1 (9,8) #6
wire n9022; //IPIN -1 (9,8) #7
wire n9023; //IPIN -1 (9,8) #8
wire n9024; //IPIN -1 (9,8) #9
wire n9025; //IPIN -1 (9,8) #10
wire n9026; //IPIN -1 (9,8) #11
wire n9027; //IPIN -1 (9,8) #12
wire n9028; //IPIN -1 (9,8) #13
wire n9029; //IPIN -1 (9,8) #14
wire n9030; //IPIN -1 (9,8) #15
wire n9031; //IPIN -1 (9,8) #16
wire n9032; //IPIN -1 (9,8) #17
wire n9033; //IPIN -1 (9,8) #18
wire n9034; //IPIN -1 (9,8) #19
wire n9035; //IPIN -1 (9,8) #20
wire n9036; //IPIN -1 (9,8) #21
wire n9037; //IPIN -1 (9,8) #22
wire n9038; //IPIN -1 (9,8) #23
wire n9039; //IPIN -1 (9,8) #24
wire n9040; //IPIN -1 (9,8) #25
wire n9041; //IPIN -1 (9,8) #26
wire n9042; //IPIN -1 (9,8) #27
wire n9043; //IPIN -1 (9,8) #28
wire n9044; //IPIN -1 (9,8) #29
wire n9045; //IPIN -1 (9,8) #30
wire n9046; //IPIN -1 (9,8) #31
wire n9047; //IPIN -1 (9,8) #32
wire n9048; //IPIN -1 (9,8) #33
wire n9049; //IPIN -1 (9,8) #34
wire n9050; //IPIN -1 (9,8) #35
wire n9051; //IPIN -1 (9,8) #36
wire n9052; //IPIN -1 (9,8) #37
wire n9053; //IPIN -1 (9,8) #38
wire n9054; //IPIN -1 (9,8) #39
wire n9055; //IPIN -1 (9,8) #40
wire n9056; //IPIN -1 (9,8) #41
wire n9057; //IPIN -1 (9,8) #42
wire n9058; //IPIN -1 (9,8) #43
wire n9059; //IPIN -1 (9,8) #44
wire n9060; //IPIN -1 (9,8) #45
wire n9061; //IPIN -1 (9,8) #46
wire n9062; //IPIN -1 (9,8) #47
wire n9063; //IPIN -1 (9,8) #48
wire n9064; //IPIN -1 (9,8) #49
wire n9065; //IPIN -1 (9,8) #50
wire n9066; //IPIN -1 (9,8) #51
wire n9067; //OPIN -1 (9,8) #52
wire n9068; //OPIN -1 (9,8) #53
wire n9069; //OPIN -1 (9,8) #54
wire n9070; //OPIN -1 (9,8) #55
wire n9071; //OPIN -1 (9,8) #56
wire n9072; //OPIN -1 (9,8) #57
wire n9073; //OPIN -1 (9,8) #58
wire n9074; //OPIN -1 (9,8) #59
wire n9075; //OPIN -1 (9,8) #60
wire n9076; //OPIN -1 (9,8) #61
wire n9077; //OPIN -1 (9,8) #62
wire n9078; //OPIN -1 (9,8) #63
wire n9079; //OPIN -1 (9,8) #64
wire n9080; //OPIN -1 (9,8) #65
wire n9081; //OPIN -1 (9,8) #66
wire n9082; //OPIN -1 (9,8) #67
wire n9083; //OPIN -1 (9,8) #68
wire n9084; //OPIN -1 (9,8) #69
wire n9085; //OPIN -1 (9,8) #70
wire n9086; //OPIN -1 (9,8) #71
wire n9087; //IPIN -1 (9,8) #72
wire n9113; //IPIN -1 (9,9) #0
wire n9114; //IPIN -1 (9,9) #1
wire n9115; //IPIN -1 (9,9) #2
wire n9116; //IPIN -1 (9,9) #3
wire n9117; //IPIN -1 (9,9) #4
wire n9118; //IPIN -1 (9,9) #5
wire n9119; //IPIN -1 (9,9) #6
wire n9120; //IPIN -1 (9,9) #7
wire n9121; //IPIN -1 (9,9) #8
wire n9122; //IPIN -1 (9,9) #9
wire n9123; //IPIN -1 (9,9) #10
wire n9124; //IPIN -1 (9,9) #11
wire n9125; //IPIN -1 (9,9) #12
wire n9126; //IPIN -1 (9,9) #13
wire n9127; //IPIN -1 (9,9) #14
wire n9128; //IPIN -1 (9,9) #15
wire n9129; //IPIN -1 (9,9) #16
wire n9130; //IPIN -1 (9,9) #17
wire n9131; //IPIN -1 (9,9) #18
wire n9132; //IPIN -1 (9,9) #19
wire n9133; //IPIN -1 (9,9) #20
wire n9134; //IPIN -1 (9,9) #21
wire n9135; //IPIN -1 (9,9) #22
wire n9136; //IPIN -1 (9,9) #23
wire n9137; //IPIN -1 (9,9) #24
wire n9138; //IPIN -1 (9,9) #25
wire n9139; //IPIN -1 (9,9) #26
wire n9140; //IPIN -1 (9,9) #27
wire n9141; //IPIN -1 (9,9) #28
wire n9142; //IPIN -1 (9,9) #29
wire n9143; //IPIN -1 (9,9) #30
wire n9144; //IPIN -1 (9,9) #31
wire n9145; //IPIN -1 (9,9) #32
wire n9146; //IPIN -1 (9,9) #33
wire n9147; //IPIN -1 (9,9) #34
wire n9148; //IPIN -1 (9,9) #35
wire n9149; //IPIN -1 (9,9) #36
wire n9150; //IPIN -1 (9,9) #37
wire n9151; //IPIN -1 (9,9) #38
wire n9152; //IPIN -1 (9,9) #39
wire n9153; //IPIN -1 (9,9) #40
wire n9154; //IPIN -1 (9,9) #41
wire n9155; //IPIN -1 (9,9) #42
wire n9156; //IPIN -1 (9,9) #43
wire n9157; //IPIN -1 (9,9) #44
wire n9158; //IPIN -1 (9,9) #45
wire n9159; //IPIN -1 (9,9) #46
wire n9160; //IPIN -1 (9,9) #47
wire n9161; //IPIN -1 (9,9) #48
wire n9162; //IPIN -1 (9,9) #49
wire n9163; //IPIN -1 (9,9) #50
wire n9164; //IPIN -1 (9,9) #51
wire n9165; //OPIN -1 (9,9) #52
wire n9166; //OPIN -1 (9,9) #53
wire n9167; //OPIN -1 (9,9) #54
wire n9168; //OPIN -1 (9,9) #55
wire n9169; //OPIN -1 (9,9) #56
wire n9170; //OPIN -1 (9,9) #57
wire n9171; //OPIN -1 (9,9) #58
wire n9172; //OPIN -1 (9,9) #59
wire n9173; //OPIN -1 (9,9) #60
wire n9174; //OPIN -1 (9,9) #61
wire n9175; //OPIN -1 (9,9) #62
wire n9176; //OPIN -1 (9,9) #63
wire n9177; //OPIN -1 (9,9) #64
wire n9178; //OPIN -1 (9,9) #65
wire n9179; //OPIN -1 (9,9) #66
wire n9180; //OPIN -1 (9,9) #67
wire n9181; //OPIN -1 (9,9) #68
wire n9182; //OPIN -1 (9,9) #69
wire n9183; //OPIN -1 (9,9) #70
wire n9184; //OPIN -1 (9,9) #71
wire n9185; //IPIN -1 (9,9) #72
wire n9210; //IPIN -1 (9,10) #0
wire n9211; //OPIN -1 (9,10) #1
wire n9212; //IPIN -1 (9,10) #2
wire n9213; //IPIN -1 (9,10) #3
wire n9214; //OPIN -1 (9,10) #4
wire n9215; //IPIN -1 (9,10) #5
wire n9216; //IPIN -1 (9,10) #6
wire n9217; //OPIN -1 (9,10) #7
wire n9218; //IPIN -1 (9,10) #8
wire n9219; //IPIN -1 (9,10) #9
wire n9220; //OPIN -1 (9,10) #10
wire n9221; //IPIN -1 (9,10) #11
wire n9222; //IPIN -1 (9,10) #12
wire n9223; //OPIN -1 (9,10) #13
wire n9224; //IPIN -1 (9,10) #14
wire n9225; //IPIN -1 (9,10) #15
wire n9226; //OPIN -1 (9,10) #16
wire n9227; //IPIN -1 (9,10) #17
wire n9228; //IPIN -1 (9,10) #18
wire n9229; //OPIN -1 (9,10) #19
wire n9230; //IPIN -1 (9,10) #20
wire n9231; //IPIN -1 (9,10) #21
wire n9232; //OPIN -1 (9,10) #22
wire n9233; //IPIN -1 (9,10) #23
wire n9258; //IPIN -1 (10,1) #0
wire n9259; //OPIN -1 (10,1) #1
wire n9260; //IPIN -1 (10,1) #2
wire n9261; //IPIN -1 (10,1) #3
wire n9262; //OPIN -1 (10,1) #4
wire n9263; //IPIN -1 (10,1) #5
wire n9264; //IPIN -1 (10,1) #6
wire n9265; //OPIN -1 (10,1) #7
wire n9266; //IPIN -1 (10,1) #8
wire n9267; //IPIN -1 (10,1) #9
wire n9268; //OPIN -1 (10,1) #10
wire n9269; //IPIN -1 (10,1) #11
wire n9270; //IPIN -1 (10,1) #12
wire n9271; //OPIN -1 (10,1) #13
wire n9272; //IPIN -1 (10,1) #14
wire n9273; //IPIN -1 (10,1) #15
wire n9274; //OPIN -1 (10,1) #16
wire n9275; //IPIN -1 (10,1) #17
wire n9276; //IPIN -1 (10,1) #18
wire n9277; //OPIN -1 (10,1) #19
wire n9278; //IPIN -1 (10,1) #20
wire n9279; //IPIN -1 (10,1) #21
wire n9280; //OPIN -1 (10,1) #22
wire n9281; //IPIN -1 (10,1) #23
wire n9306; //IPIN -1 (10,2) #0
wire n9307; //OPIN -1 (10,2) #1
wire n9308; //IPIN -1 (10,2) #2
wire n9309; //IPIN -1 (10,2) #3
wire n9310; //OPIN -1 (10,2) #4
wire n9311; //IPIN -1 (10,2) #5
wire n9312; //IPIN -1 (10,2) #6
wire n9313; //OPIN -1 (10,2) #7
wire n9314; //IPIN -1 (10,2) #8
wire n9315; //IPIN -1 (10,2) #9
wire n9316; //OPIN -1 (10,2) #10
wire n9317; //IPIN -1 (10,2) #11
wire n9318; //IPIN -1 (10,2) #12
wire n9319; //OPIN -1 (10,2) #13
wire n9320; //IPIN -1 (10,2) #14
wire n9321; //IPIN -1 (10,2) #15
wire n9322; //OPIN -1 (10,2) #16
wire n9323; //IPIN -1 (10,2) #17
wire n9324; //IPIN -1 (10,2) #18
wire n9325; //OPIN -1 (10,2) #19
wire n9326; //IPIN -1 (10,2) #20
wire n9327; //IPIN -1 (10,2) #21
wire n9328; //OPIN -1 (10,2) #22
wire n9329; //IPIN -1 (10,2) #23
wire n9354; //IPIN -1 (10,3) #0
wire n9355; //OPIN -1 (10,3) #1
wire n9356; //IPIN -1 (10,3) #2
wire n9357; //IPIN -1 (10,3) #3
wire n9358; //OPIN -1 (10,3) #4
wire n9359; //IPIN -1 (10,3) #5
wire n9360; //IPIN -1 (10,3) #6
wire n9361; //OPIN -1 (10,3) #7
wire n9362; //IPIN -1 (10,3) #8
wire n9363; //IPIN -1 (10,3) #9
wire n9364; //OPIN -1 (10,3) #10
wire n9365; //IPIN -1 (10,3) #11
wire n9366; //IPIN -1 (10,3) #12
wire n9367; //OPIN -1 (10,3) #13
wire n9368; //IPIN -1 (10,3) #14
wire n9369; //IPIN -1 (10,3) #15
wire n9370; //OPIN -1 (10,3) #16
wire n9371; //IPIN -1 (10,3) #17
wire n9372; //IPIN -1 (10,3) #18
wire n9373; //OPIN -1 (10,3) #19
wire n9374; //IPIN -1 (10,3) #20
wire n9375; //IPIN -1 (10,3) #21
wire n9376; //OPIN -1 (10,3) #22
wire n9377; //IPIN -1 (10,3) #23
wire n9402; //IPIN -1 (10,4) #0
wire n9403; //OPIN -1 (10,4) #1
wire n9404; //IPIN -1 (10,4) #2
wire n9405; //IPIN -1 (10,4) #3
wire n9406; //OPIN -1 (10,4) #4
wire n9407; //IPIN -1 (10,4) #5
wire n9408; //IPIN -1 (10,4) #6
wire n9409; //OPIN -1 (10,4) #7
wire n9410; //IPIN -1 (10,4) #8
wire n9411; //IPIN -1 (10,4) #9
wire n9412; //OPIN -1 (10,4) #10
wire n9413; //IPIN -1 (10,4) #11
wire n9414; //IPIN -1 (10,4) #12
wire n9415; //OPIN -1 (10,4) #13
wire n9416; //IPIN -1 (10,4) #14
wire n9417; //IPIN -1 (10,4) #15
wire n9418; //OPIN -1 (10,4) #16
wire n9419; //IPIN -1 (10,4) #17
wire n9420; //IPIN -1 (10,4) #18
wire n9421; //OPIN -1 (10,4) #19
wire n9422; //IPIN -1 (10,4) #20
wire n9423; //IPIN -1 (10,4) #21
wire n9424; //OPIN -1 (10,4) #22
wire n9425; //IPIN -1 (10,4) #23
wire n9450; //IPIN -1 (10,5) #0
wire n9451; //OPIN -1 (10,5) #1
wire n9452; //IPIN -1 (10,5) #2
wire n9453; //IPIN -1 (10,5) #3
wire n9454; //OPIN -1 (10,5) #4
wire n9455; //IPIN -1 (10,5) #5
wire n9456; //IPIN -1 (10,5) #6
wire n9457; //OPIN -1 (10,5) #7
wire n9458; //IPIN -1 (10,5) #8
wire n9459; //IPIN -1 (10,5) #9
wire n9460; //OPIN -1 (10,5) #10
wire n9461; //IPIN -1 (10,5) #11
wire n9462; //IPIN -1 (10,5) #12
wire n9463; //OPIN -1 (10,5) #13
wire n9464; //IPIN -1 (10,5) #14
wire n9465; //IPIN -1 (10,5) #15
wire n9466; //OPIN -1 (10,5) #16
wire n9467; //IPIN -1 (10,5) #17
wire n9468; //IPIN -1 (10,5) #18
wire n9469; //OPIN -1 (10,5) #19
wire n9470; //IPIN -1 (10,5) #20
wire n9471; //IPIN -1 (10,5) #21
wire n9472; //OPIN -1 (10,5) #22
wire n9473; //IPIN -1 (10,5) #23
wire n9498; //IPIN -1 (10,6) #0
wire n9499; //OPIN -1 (10,6) #1
wire n9500; //IPIN -1 (10,6) #2
wire n9501; //IPIN -1 (10,6) #3
wire n9502; //OPIN -1 (10,6) #4
wire n9503; //IPIN -1 (10,6) #5
wire n9504; //IPIN -1 (10,6) #6
wire n9505; //OPIN -1 (10,6) #7
wire n9506; //IPIN -1 (10,6) #8
wire n9507; //IPIN -1 (10,6) #9
wire n9508; //OPIN -1 (10,6) #10
wire n9509; //IPIN -1 (10,6) #11
wire n9510; //IPIN -1 (10,6) #12
wire n9511; //OPIN -1 (10,6) #13
wire n9512; //IPIN -1 (10,6) #14
wire n9513; //IPIN -1 (10,6) #15
wire n9514; //OPIN -1 (10,6) #16
wire n9515; //IPIN -1 (10,6) #17
wire n9516; //IPIN -1 (10,6) #18
wire n9517; //OPIN -1 (10,6) #19
wire n9518; //IPIN -1 (10,6) #20
wire n9519; //IPIN -1 (10,6) #21
wire n9520; //OPIN -1 (10,6) #22
wire n9521; //IPIN -1 (10,6) #23
wire n9546; //IPIN -1 (10,7) #0
wire n9547; //OPIN -1 (10,7) #1
wire n9548; //IPIN -1 (10,7) #2
wire n9549; //IPIN -1 (10,7) #3
wire n9550; //OPIN -1 (10,7) #4
wire n9551; //IPIN -1 (10,7) #5
wire n9552; //IPIN -1 (10,7) #6
wire n9553; //OPIN -1 (10,7) #7
wire n9554; //IPIN -1 (10,7) #8
wire n9555; //IPIN -1 (10,7) #9
wire n9556; //OPIN -1 (10,7) #10
wire n9557; //IPIN -1 (10,7) #11
wire n9558; //IPIN -1 (10,7) #12
wire n9559; //OPIN -1 (10,7) #13
wire n9560; //IPIN -1 (10,7) #14
wire n9561; //IPIN -1 (10,7) #15
wire n9562; //OPIN -1 (10,7) #16
wire n9563; //IPIN -1 (10,7) #17
wire n9564; //IPIN -1 (10,7) #18
wire n9565; //OPIN -1 (10,7) #19
wire n9566; //IPIN -1 (10,7) #20
wire n9567; //IPIN -1 (10,7) #21
wire n9568; //OPIN -1 (10,7) #22
wire n9569; //IPIN -1 (10,7) #23
wire n9594; //IPIN -1 (10,8) #0
wire n9595; //OPIN -1 (10,8) #1
wire n9596; //IPIN -1 (10,8) #2
wire n9597; //IPIN -1 (10,8) #3
wire n9598; //OPIN -1 (10,8) #4
wire n9599; //IPIN -1 (10,8) #5
wire n9600; //IPIN -1 (10,8) #6
wire n9601; //OPIN -1 (10,8) #7
wire n9602; //IPIN -1 (10,8) #8
wire n9603; //IPIN -1 (10,8) #9
wire n9604; //OPIN -1 (10,8) #10
wire n9605; //IPIN -1 (10,8) #11
wire n9606; //IPIN -1 (10,8) #12
wire n9607; //OPIN -1 (10,8) #13
wire n9608; //IPIN -1 (10,8) #14
wire n9609; //IPIN -1 (10,8) #15
wire n9610; //OPIN -1 (10,8) #16
wire n9611; //IPIN -1 (10,8) #17
wire n9612; //IPIN -1 (10,8) #18
wire n9613; //OPIN -1 (10,8) #19
wire n9614; //IPIN -1 (10,8) #20
wire n9615; //IPIN -1 (10,8) #21
wire n9616; //OPIN -1 (10,8) #22
wire n9617; //IPIN -1 (10,8) #23
wire n9642; //IPIN -1 (10,9) #0
wire n9643; //OPIN -1 (10,9) #1
wire n9644; //IPIN -1 (10,9) #2
wire n9645; //IPIN -1 (10,9) #3
wire n9646; //OPIN -1 (10,9) #4
wire n9647; //IPIN -1 (10,9) #5
wire n9648; //IPIN -1 (10,9) #6
wire n9649; //OPIN -1 (10,9) #7
wire n9650; //IPIN -1 (10,9) #8
wire n9651; //IPIN -1 (10,9) #9
wire n9652; //OPIN -1 (10,9) #10
wire n9653; //IPIN -1 (10,9) #11
wire n9654; //IPIN -1 (10,9) #12
wire n9655; //OPIN -1 (10,9) #13
wire n9656; //IPIN -1 (10,9) #14
wire n9657; //IPIN -1 (10,9) #15
wire n9658; //OPIN -1 (10,9) #16
wire n9659; //IPIN -1 (10,9) #17
wire n9660; //IPIN -1 (10,9) #18
wire n9661; //OPIN -1 (10,9) #19
wire n9662; //IPIN -1 (10,9) #20
wire n9663; //IPIN -1 (10,9) #21
wire n9664; //OPIN -1 (10,9) #22
wire n9665; //IPIN -1 (10,9) #23
wire n9666; //CHANX 4 (1,0) #0
wire n9666_0;
wire n9666_1;
buffer_wire buffer_9666_1 (.in(n9666_0), .out(n9666_1));
wire n9667; //CHANX 4 (1,0) #1
wire n9667_0;
wire n9667_1;
buffer_wire buffer_9667_1 (.in(n9667_0), .out(n9667_1));
wire n9668; //CHANX 1 (1,0) #2
wire n9668_0;
wire n9669; //CHANX 1 (1,0) #3
wire n9669_0;
wire n9670; //CHANX 2 (1,0) #4
wire n9670_0;
wire n9671; //CHANX 2 (1,0) #5
wire n9671_0;
wire n9672; //CHANX 3 (1,0) #6
wire n9672_0;
wire n9673; //CHANX 3 (1,0) #7
wire n9673_0;
wire n9674; //CHANX 4 (1,0) #8
wire n9674_0;
wire n9674_1;
buffer_wire buffer_9674_1 (.in(n9674_0), .out(n9674_1));
wire n9675; //CHANX 4 (1,0) #9
wire n9675_0;
wire n9675_1;
buffer_wire buffer_9675_1 (.in(n9675_0), .out(n9675_1));
wire n9676; //CHANX 1 (1,0) #10
wire n9676_0;
wire n9677; //CHANX 1 (1,0) #11
wire n9677_0;
wire n9678; //CHANX 2 (1,0) #12
wire n9678_0;
wire n9679; //CHANX 2 (1,0) #13
wire n9679_0;
wire n9680; //CHANX 3 (1,0) #14
wire n9680_0;
wire n9681; //CHANX 3 (1,0) #15
wire n9681_0;
wire n9682; //CHANX 4 (1,0) #16
wire n9682_0;
wire n9682_1;
buffer_wire buffer_9682_1 (.in(n9682_0), .out(n9682_1));
wire n9683; //CHANX 4 (1,0) #17
wire n9683_0;
wire n9683_1;
buffer_wire buffer_9683_1 (.in(n9683_0), .out(n9683_1));
wire n9684; //CHANX 1 (1,0) #18
wire n9684_0;
wire n9685; //CHANX 1 (1,0) #19
wire n9685_0;
wire n9686; //CHANX 2 (1,0) #20
wire n9686_0;
wire n9687; //CHANX 2 (1,0) #21
wire n9687_0;
wire n9688; //CHANX 3 (1,0) #22
wire n9688_0;
wire n9689; //CHANX 3 (1,0) #23
wire n9689_0;
wire n9690; //CHANX 4 (1,0) #24
wire n9690_0;
wire n9690_1;
buffer_wire buffer_9690_1 (.in(n9690_0), .out(n9690_1));
wire n9691; //CHANX 4 (1,0) #25
wire n9691_0;
wire n9691_1;
buffer_wire buffer_9691_1 (.in(n9691_0), .out(n9691_1));
wire n9692; //CHANX 1 (1,0) #26
wire n9692_0;
wire n9693; //CHANX 1 (1,0) #27
wire n9693_0;
wire n9694; //CHANX 2 (1,0) #28
wire n9694_0;
wire n9695; //CHANX 2 (1,0) #29
wire n9695_0;
wire n9696; //CHANX 3 (1,0) #30
wire n9696_0;
wire n9697; //CHANX 3 (1,0) #31
wire n9697_0;
wire n9698; //CHANX 4 (1,0) #32
wire n9698_0;
wire n9698_1;
buffer_wire buffer_9698_1 (.in(n9698_0), .out(n9698_1));
wire n9699; //CHANX 4 (1,0) #33
wire n9699_0;
wire n9699_1;
buffer_wire buffer_9699_1 (.in(n9699_0), .out(n9699_1));
wire n9700; //CHANX 1 (1,0) #34
wire n9700_0;
wire n9701; //CHANX 1 (1,0) #35
wire n9701_0;
wire n9702; //CHANX 2 (1,0) #36
wire n9702_0;
wire n9703; //CHANX 2 (1,0) #37
wire n9703_0;
wire n9704; //CHANX 3 (1,0) #38
wire n9704_0;
wire n9705; //CHANX 3 (1,0) #39
wire n9705_0;
wire n9706; //CHANX 4 (1,0) #40
wire n9706_0;
wire n9706_1;
buffer_wire buffer_9706_1 (.in(n9706_0), .out(n9706_1));
wire n9707; //CHANX 4 (1,0) #41
wire n9707_0;
wire n9707_1;
buffer_wire buffer_9707_1 (.in(n9707_0), .out(n9707_1));
wire n9708; //CHANX 1 (1,0) #42
wire n9708_0;
wire n9709; //CHANX 1 (1,0) #43
wire n9709_0;
wire n9710; //CHANX 2 (1,0) #44
wire n9710_0;
wire n9711; //CHANX 2 (1,0) #45
wire n9711_0;
wire n9712; //CHANX 3 (1,0) #46
wire n9712_0;
wire n9713; //CHANX 3 (1,0) #47
wire n9713_0;
wire n9714; //CHANX 4 (1,0) #48
wire n9714_0;
wire n9714_1;
buffer_wire buffer_9714_1 (.in(n9714_0), .out(n9714_1));
wire n9715; //CHANX 4 (1,0) #49
wire n9715_0;
wire n9715_1;
buffer_wire buffer_9715_1 (.in(n9715_0), .out(n9715_1));
wire n9716; //CHANX 1 (1,0) #50
wire n9716_0;
wire n9717; //CHANX 1 (1,0) #51
wire n9717_0;
wire n9718; //CHANX 2 (1,0) #52
wire n9718_0;
wire n9719; //CHANX 2 (1,0) #53
wire n9719_0;
wire n9720; //CHANX 3 (1,0) #54
wire n9720_0;
wire n9721; //CHANX 3 (1,0) #55
wire n9721_0;
wire n9722; //CHANX 4 (1,0) #56
wire n9722_0;
wire n9722_1;
buffer_wire buffer_9722_1 (.in(n9722_0), .out(n9722_1));
wire n9723; //CHANX 4 (1,0) #57
wire n9723_0;
wire n9723_1;
buffer_wire buffer_9723_1 (.in(n9723_0), .out(n9723_1));
wire n9724; //CHANX 1 (1,0) #58
wire n9724_0;
wire n9725; //CHANX 1 (1,0) #59
wire n9725_0;
wire n9726; //CHANX 2 (1,0) #60
wire n9726_0;
wire n9727; //CHANX 2 (1,0) #61
wire n9727_0;
wire n9728; //CHANX 3 (1,0) #62
wire n9728_0;
wire n9729; //CHANX 3 (1,0) #63
wire n9729_0;
wire n9730; //CHANX 4 (1,0) #64
wire n9730_0;
wire n9730_1;
buffer_wire buffer_9730_1 (.in(n9730_0), .out(n9730_1));
wire n9731; //CHANX 4 (1,0) #65
wire n9731_0;
wire n9731_1;
buffer_wire buffer_9731_1 (.in(n9731_0), .out(n9731_1));
wire n9732; //CHANX 1 (1,0) #66
wire n9732_0;
wire n9733; //CHANX 1 (1,0) #67
wire n9733_0;
wire n9734; //CHANX 2 (1,0) #68
wire n9734_0;
wire n9735; //CHANX 2 (1,0) #69
wire n9735_0;
wire n9736; //CHANX 3 (1,0) #70
wire n9736_0;
wire n9737; //CHANX 3 (1,0) #71
wire n9737_0;
wire n9738; //CHANX 4 (1,0) #72
wire n9738_0;
wire n9738_1;
buffer_wire buffer_9738_1 (.in(n9738_0), .out(n9738_1));
wire n9739; //CHANX 4 (1,0) #73
wire n9739_0;
wire n9739_1;
buffer_wire buffer_9739_1 (.in(n9739_0), .out(n9739_1));
wire n9740; //CHANX 1 (1,0) #74
wire n9740_0;
wire n9741; //CHANX 1 (1,0) #75
wire n9741_0;
wire n9742; //CHANX 2 (1,0) #76
wire n9742_0;
wire n9743; //CHANX 2 (1,0) #77
wire n9743_0;
wire n9744; //CHANX 3 (1,0) #78
wire n9744_0;
wire n9745; //CHANX 3 (1,0) #79
wire n9745_0;
wire n9746; //CHANX 8 (1,0) #80
wire n9746_0;
wire n9746_1;
wire n9746_2;
buffer_wire buffer_9746_2 (.in(n9746_1), .out(n9746_2));
buffer_wire buffer_9746_1 (.in(n9746_0), .out(n9746_1));
wire n9747; //CHANX 8 (1,0) #81
wire n9747_0;
wire n9747_1;
wire n9747_2;
buffer_wire buffer_9747_2 (.in(n9747_1), .out(n9747_2));
buffer_wire buffer_9747_1 (.in(n9747_0), .out(n9747_1));
wire n9748; //CHANX 9 (1,0) #82
wire n9748_0;
wire n9748_1;
wire n9748_2;
buffer_wire buffer_9748_2 (.in(n9748_1), .out(n9748_2));
buffer_wire buffer_9748_1 (.in(n9748_0), .out(n9748_1));
wire n9749; //CHANX 9 (1,0) #83
wire n9749_0;
wire n9749_1;
wire n9749_2;
buffer_wire buffer_9749_2 (.in(n9749_1), .out(n9749_2));
buffer_wire buffer_9749_1 (.in(n9749_0), .out(n9749_1));
wire n9750; //CHANX 9 (1,0) #84
wire n9750_0;
wire n9750_1;
wire n9750_2;
buffer_wire buffer_9750_2 (.in(n9750_1), .out(n9750_2));
buffer_wire buffer_9750_1 (.in(n9750_0), .out(n9750_1));
wire n9751; //CHANX 9 (1,0) #85
wire n9751_0;
wire n9751_1;
wire n9751_2;
buffer_wire buffer_9751_2 (.in(n9751_1), .out(n9751_2));
buffer_wire buffer_9751_1 (.in(n9751_0), .out(n9751_1));
wire n9752; //CHANX 9 (1,0) #86
wire n9752_0;
wire n9752_1;
wire n9752_2;
buffer_wire buffer_9752_2 (.in(n9752_1), .out(n9752_2));
buffer_wire buffer_9752_1 (.in(n9752_0), .out(n9752_1));
wire n9753; //CHANX 9 (1,0) #87
wire n9753_0;
wire n9753_1;
wire n9753_2;
buffer_wire buffer_9753_2 (.in(n9753_1), .out(n9753_2));
buffer_wire buffer_9753_1 (.in(n9753_0), .out(n9753_1));
wire n9754; //CHANX 9 (1,0) #88
wire n9754_0;
wire n9754_1;
wire n9754_2;
buffer_wire buffer_9754_2 (.in(n9754_1), .out(n9754_2));
buffer_wire buffer_9754_1 (.in(n9754_0), .out(n9754_1));
wire n9755; //CHANX 9 (1,0) #89
wire n9755_0;
wire n9755_1;
wire n9755_2;
buffer_wire buffer_9755_2 (.in(n9755_1), .out(n9755_2));
buffer_wire buffer_9755_1 (.in(n9755_0), .out(n9755_1));
wire n9756; //CHANX 9 (1,0) #90
wire n9756_0;
wire n9756_1;
wire n9756_2;
buffer_wire buffer_9756_2 (.in(n9756_1), .out(n9756_2));
buffer_wire buffer_9756_1 (.in(n9756_0), .out(n9756_1));
wire n9757; //CHANX 9 (1,0) #91
wire n9757_0;
wire n9757_1;
wire n9757_2;
buffer_wire buffer_9757_2 (.in(n9757_1), .out(n9757_2));
buffer_wire buffer_9757_1 (.in(n9757_0), .out(n9757_1));
wire n9758; //CHANX 4 (2,0) #2
wire n9758_0;
wire n9758_1;
buffer_wire buffer_9758_1 (.in(n9758_0), .out(n9758_1));
wire n9759; //CHANX 4 (2,0) #3
wire n9759_0;
wire n9759_1;
buffer_wire buffer_9759_1 (.in(n9759_0), .out(n9759_1));
wire n9760; //CHANX 4 (2,0) #10
wire n9760_0;
wire n9760_1;
buffer_wire buffer_9760_1 (.in(n9760_0), .out(n9760_1));
wire n9761; //CHANX 4 (2,0) #11
wire n9761_0;
wire n9761_1;
buffer_wire buffer_9761_1 (.in(n9761_0), .out(n9761_1));
wire n9762; //CHANX 4 (2,0) #18
wire n9762_0;
wire n9762_1;
buffer_wire buffer_9762_1 (.in(n9762_0), .out(n9762_1));
wire n9763; //CHANX 4 (2,0) #19
wire n9763_0;
wire n9763_1;
buffer_wire buffer_9763_1 (.in(n9763_0), .out(n9763_1));
wire n9764; //CHANX 4 (2,0) #26
wire n9764_0;
wire n9764_1;
buffer_wire buffer_9764_1 (.in(n9764_0), .out(n9764_1));
wire n9765; //CHANX 4 (2,0) #27
wire n9765_0;
wire n9765_1;
buffer_wire buffer_9765_1 (.in(n9765_0), .out(n9765_1));
wire n9766; //CHANX 4 (2,0) #34
wire n9766_0;
wire n9766_1;
buffer_wire buffer_9766_1 (.in(n9766_0), .out(n9766_1));
wire n9767; //CHANX 4 (2,0) #35
wire n9767_0;
wire n9767_1;
buffer_wire buffer_9767_1 (.in(n9767_0), .out(n9767_1));
wire n9768; //CHANX 4 (2,0) #42
wire n9768_0;
wire n9768_1;
buffer_wire buffer_9768_1 (.in(n9768_0), .out(n9768_1));
wire n9769; //CHANX 4 (2,0) #43
wire n9769_0;
wire n9769_1;
buffer_wire buffer_9769_1 (.in(n9769_0), .out(n9769_1));
wire n9770; //CHANX 4 (2,0) #50
wire n9770_0;
wire n9770_1;
buffer_wire buffer_9770_1 (.in(n9770_0), .out(n9770_1));
wire n9771; //CHANX 4 (2,0) #51
wire n9771_0;
wire n9771_1;
buffer_wire buffer_9771_1 (.in(n9771_0), .out(n9771_1));
wire n9772; //CHANX 4 (2,0) #58
wire n9772_0;
wire n9772_1;
buffer_wire buffer_9772_1 (.in(n9772_0), .out(n9772_1));
wire n9773; //CHANX 4 (2,0) #59
wire n9773_0;
wire n9773_1;
buffer_wire buffer_9773_1 (.in(n9773_0), .out(n9773_1));
wire n9774; //CHANX 4 (2,0) #66
wire n9774_0;
wire n9774_1;
buffer_wire buffer_9774_1 (.in(n9774_0), .out(n9774_1));
wire n9775; //CHANX 4 (2,0) #67
wire n9775_0;
wire n9775_1;
buffer_wire buffer_9775_1 (.in(n9775_0), .out(n9775_1));
wire n9776; //CHANX 4 (2,0) #74
wire n9776_0;
wire n9776_1;
buffer_wire buffer_9776_1 (.in(n9776_0), .out(n9776_1));
wire n9777; //CHANX 4 (2,0) #75
wire n9777_0;
wire n9777_1;
buffer_wire buffer_9777_1 (.in(n9777_0), .out(n9777_1));
wire n9778; //CHANX 4 (3,0) #4
wire n9778_0;
wire n9778_1;
buffer_wire buffer_9778_1 (.in(n9778_0), .out(n9778_1));
wire n9779; //CHANX 4 (3,0) #5
wire n9779_0;
wire n9779_1;
buffer_wire buffer_9779_1 (.in(n9779_0), .out(n9779_1));
wire n9780; //CHANX 4 (3,0) #12
wire n9780_0;
wire n9780_1;
buffer_wire buffer_9780_1 (.in(n9780_0), .out(n9780_1));
wire n9781; //CHANX 4 (3,0) #13
wire n9781_0;
wire n9781_1;
buffer_wire buffer_9781_1 (.in(n9781_0), .out(n9781_1));
wire n9782; //CHANX 4 (3,0) #20
wire n9782_0;
wire n9782_1;
buffer_wire buffer_9782_1 (.in(n9782_0), .out(n9782_1));
wire n9783; //CHANX 4 (3,0) #21
wire n9783_0;
wire n9783_1;
buffer_wire buffer_9783_1 (.in(n9783_0), .out(n9783_1));
wire n9784; //CHANX 4 (3,0) #28
wire n9784_0;
wire n9784_1;
buffer_wire buffer_9784_1 (.in(n9784_0), .out(n9784_1));
wire n9785; //CHANX 4 (3,0) #29
wire n9785_0;
wire n9785_1;
buffer_wire buffer_9785_1 (.in(n9785_0), .out(n9785_1));
wire n9786; //CHANX 4 (3,0) #36
wire n9786_0;
wire n9786_1;
buffer_wire buffer_9786_1 (.in(n9786_0), .out(n9786_1));
wire n9787; //CHANX 4 (3,0) #37
wire n9787_0;
wire n9787_1;
buffer_wire buffer_9787_1 (.in(n9787_0), .out(n9787_1));
wire n9788; //CHANX 4 (3,0) #44
wire n9788_0;
wire n9788_1;
buffer_wire buffer_9788_1 (.in(n9788_0), .out(n9788_1));
wire n9789; //CHANX 4 (3,0) #45
wire n9789_0;
wire n9789_1;
buffer_wire buffer_9789_1 (.in(n9789_0), .out(n9789_1));
wire n9790; //CHANX 4 (3,0) #52
wire n9790_0;
wire n9790_1;
buffer_wire buffer_9790_1 (.in(n9790_0), .out(n9790_1));
wire n9791; //CHANX 4 (3,0) #53
wire n9791_0;
wire n9791_1;
buffer_wire buffer_9791_1 (.in(n9791_0), .out(n9791_1));
wire n9792; //CHANX 4 (3,0) #60
wire n9792_0;
wire n9792_1;
buffer_wire buffer_9792_1 (.in(n9792_0), .out(n9792_1));
wire n9793; //CHANX 4 (3,0) #61
wire n9793_0;
wire n9793_1;
buffer_wire buffer_9793_1 (.in(n9793_0), .out(n9793_1));
wire n9794; //CHANX 4 (3,0) #68
wire n9794_0;
wire n9794_1;
buffer_wire buffer_9794_1 (.in(n9794_0), .out(n9794_1));
wire n9795; //CHANX 4 (3,0) #69
wire n9795_0;
wire n9795_1;
buffer_wire buffer_9795_1 (.in(n9795_0), .out(n9795_1));
wire n9796; //CHANX 4 (3,0) #76
wire n9796_0;
wire n9796_1;
buffer_wire buffer_9796_1 (.in(n9796_0), .out(n9796_1));
wire n9797; //CHANX 4 (3,0) #77
wire n9797_0;
wire n9797_1;
buffer_wire buffer_9797_1 (.in(n9797_0), .out(n9797_1));
wire n9798; //CHANX 4 (4,0) #6
wire n9798_0;
wire n9798_1;
buffer_wire buffer_9798_1 (.in(n9798_0), .out(n9798_1));
wire n9799; //CHANX 4 (4,0) #7
wire n9799_0;
wire n9799_1;
buffer_wire buffer_9799_1 (.in(n9799_0), .out(n9799_1));
wire n9800; //CHANX 4 (4,0) #14
wire n9800_0;
wire n9800_1;
buffer_wire buffer_9800_1 (.in(n9800_0), .out(n9800_1));
wire n9801; //CHANX 4 (4,0) #15
wire n9801_0;
wire n9801_1;
buffer_wire buffer_9801_1 (.in(n9801_0), .out(n9801_1));
wire n9802; //CHANX 4 (4,0) #22
wire n9802_0;
wire n9802_1;
buffer_wire buffer_9802_1 (.in(n9802_0), .out(n9802_1));
wire n9803; //CHANX 4 (4,0) #23
wire n9803_0;
wire n9803_1;
buffer_wire buffer_9803_1 (.in(n9803_0), .out(n9803_1));
wire n9804; //CHANX 4 (4,0) #30
wire n9804_0;
wire n9804_1;
buffer_wire buffer_9804_1 (.in(n9804_0), .out(n9804_1));
wire n9805; //CHANX 4 (4,0) #31
wire n9805_0;
wire n9805_1;
buffer_wire buffer_9805_1 (.in(n9805_0), .out(n9805_1));
wire n9806; //CHANX 4 (4,0) #38
wire n9806_0;
wire n9806_1;
buffer_wire buffer_9806_1 (.in(n9806_0), .out(n9806_1));
wire n9807; //CHANX 4 (4,0) #39
wire n9807_0;
wire n9807_1;
buffer_wire buffer_9807_1 (.in(n9807_0), .out(n9807_1));
wire n9808; //CHANX 4 (4,0) #46
wire n9808_0;
wire n9808_1;
buffer_wire buffer_9808_1 (.in(n9808_0), .out(n9808_1));
wire n9809; //CHANX 4 (4,0) #47
wire n9809_0;
wire n9809_1;
buffer_wire buffer_9809_1 (.in(n9809_0), .out(n9809_1));
wire n9810; //CHANX 4 (4,0) #54
wire n9810_0;
wire n9810_1;
buffer_wire buffer_9810_1 (.in(n9810_0), .out(n9810_1));
wire n9811; //CHANX 4 (4,0) #55
wire n9811_0;
wire n9811_1;
buffer_wire buffer_9811_1 (.in(n9811_0), .out(n9811_1));
wire n9812; //CHANX 4 (4,0) #62
wire n9812_0;
wire n9812_1;
buffer_wire buffer_9812_1 (.in(n9812_0), .out(n9812_1));
wire n9813; //CHANX 4 (4,0) #63
wire n9813_0;
wire n9813_1;
buffer_wire buffer_9813_1 (.in(n9813_0), .out(n9813_1));
wire n9814; //CHANX 4 (4,0) #70
wire n9814_0;
wire n9814_1;
buffer_wire buffer_9814_1 (.in(n9814_0), .out(n9814_1));
wire n9815; //CHANX 4 (4,0) #71
wire n9815_0;
wire n9815_1;
buffer_wire buffer_9815_1 (.in(n9815_0), .out(n9815_1));
wire n9816; //CHANX 4 (4,0) #78
wire n9816_0;
wire n9816_1;
buffer_wire buffer_9816_1 (.in(n9816_0), .out(n9816_1));
wire n9817; //CHANX 4 (4,0) #79
wire n9817_0;
wire n9817_1;
buffer_wire buffer_9817_1 (.in(n9817_0), .out(n9817_1));
wire n9818; //CHANX 4 (5,0) #0
wire n9818_0;
wire n9818_1;
buffer_wire buffer_9818_1 (.in(n9818_0), .out(n9818_1));
wire n9819; //CHANX 4 (5,0) #1
wire n9819_0;
wire n9819_1;
buffer_wire buffer_9819_1 (.in(n9819_0), .out(n9819_1));
wire n9820; //CHANX 4 (5,0) #8
wire n9820_0;
wire n9820_1;
buffer_wire buffer_9820_1 (.in(n9820_0), .out(n9820_1));
wire n9821; //CHANX 4 (5,0) #9
wire n9821_0;
wire n9821_1;
buffer_wire buffer_9821_1 (.in(n9821_0), .out(n9821_1));
wire n9822; //CHANX 4 (5,0) #16
wire n9822_0;
wire n9822_1;
buffer_wire buffer_9822_1 (.in(n9822_0), .out(n9822_1));
wire n9823; //CHANX 4 (5,0) #17
wire n9823_0;
wire n9823_1;
buffer_wire buffer_9823_1 (.in(n9823_0), .out(n9823_1));
wire n9824; //CHANX 4 (5,0) #24
wire n9824_0;
wire n9824_1;
buffer_wire buffer_9824_1 (.in(n9824_0), .out(n9824_1));
wire n9825; //CHANX 4 (5,0) #25
wire n9825_0;
wire n9825_1;
buffer_wire buffer_9825_1 (.in(n9825_0), .out(n9825_1));
wire n9826; //CHANX 4 (5,0) #32
wire n9826_0;
wire n9826_1;
buffer_wire buffer_9826_1 (.in(n9826_0), .out(n9826_1));
wire n9827; //CHANX 4 (5,0) #33
wire n9827_0;
wire n9827_1;
buffer_wire buffer_9827_1 (.in(n9827_0), .out(n9827_1));
wire n9828; //CHANX 4 (5,0) #40
wire n9828_0;
wire n9828_1;
buffer_wire buffer_9828_1 (.in(n9828_0), .out(n9828_1));
wire n9829; //CHANX 4 (5,0) #41
wire n9829_0;
wire n9829_1;
buffer_wire buffer_9829_1 (.in(n9829_0), .out(n9829_1));
wire n9830; //CHANX 4 (5,0) #48
wire n9830_0;
wire n9830_1;
buffer_wire buffer_9830_1 (.in(n9830_0), .out(n9830_1));
wire n9831; //CHANX 4 (5,0) #49
wire n9831_0;
wire n9831_1;
buffer_wire buffer_9831_1 (.in(n9831_0), .out(n9831_1));
wire n9832; //CHANX 4 (5,0) #56
wire n9832_0;
wire n9832_1;
buffer_wire buffer_9832_1 (.in(n9832_0), .out(n9832_1));
wire n9833; //CHANX 4 (5,0) #57
wire n9833_0;
wire n9833_1;
buffer_wire buffer_9833_1 (.in(n9833_0), .out(n9833_1));
wire n9834; //CHANX 4 (5,0) #64
wire n9834_0;
wire n9834_1;
buffer_wire buffer_9834_1 (.in(n9834_0), .out(n9834_1));
wire n9835; //CHANX 4 (5,0) #65
wire n9835_0;
wire n9835_1;
buffer_wire buffer_9835_1 (.in(n9835_0), .out(n9835_1));
wire n9836; //CHANX 4 (5,0) #72
wire n9836_0;
wire n9836_1;
buffer_wire buffer_9836_1 (.in(n9836_0), .out(n9836_1));
wire n9837; //CHANX 4 (5,0) #73
wire n9837_0;
wire n9837_1;
buffer_wire buffer_9837_1 (.in(n9837_0), .out(n9837_1));
wire n9838; //CHANX 4 (6,0) #2
wire n9838_0;
wire n9838_1;
buffer_wire buffer_9838_1 (.in(n9838_0), .out(n9838_1));
wire n9839; //CHANX 4 (6,0) #3
wire n9839_0;
wire n9839_1;
buffer_wire buffer_9839_1 (.in(n9839_0), .out(n9839_1));
wire n9840; //CHANX 4 (6,0) #10
wire n9840_0;
wire n9840_1;
buffer_wire buffer_9840_1 (.in(n9840_0), .out(n9840_1));
wire n9841; //CHANX 4 (6,0) #11
wire n9841_0;
wire n9841_1;
buffer_wire buffer_9841_1 (.in(n9841_0), .out(n9841_1));
wire n9842; //CHANX 4 (6,0) #18
wire n9842_0;
wire n9842_1;
buffer_wire buffer_9842_1 (.in(n9842_0), .out(n9842_1));
wire n9843; //CHANX 4 (6,0) #19
wire n9843_0;
wire n9843_1;
buffer_wire buffer_9843_1 (.in(n9843_0), .out(n9843_1));
wire n9844; //CHANX 4 (6,0) #26
wire n9844_0;
wire n9844_1;
buffer_wire buffer_9844_1 (.in(n9844_0), .out(n9844_1));
wire n9845; //CHANX 4 (6,0) #27
wire n9845_0;
wire n9845_1;
buffer_wire buffer_9845_1 (.in(n9845_0), .out(n9845_1));
wire n9846; //CHANX 4 (6,0) #34
wire n9846_0;
wire n9846_1;
buffer_wire buffer_9846_1 (.in(n9846_0), .out(n9846_1));
wire n9847; //CHANX 4 (6,0) #35
wire n9847_0;
wire n9847_1;
buffer_wire buffer_9847_1 (.in(n9847_0), .out(n9847_1));
wire n9848; //CHANX 4 (6,0) #42
wire n9848_0;
wire n9848_1;
buffer_wire buffer_9848_1 (.in(n9848_0), .out(n9848_1));
wire n9849; //CHANX 4 (6,0) #43
wire n9849_0;
wire n9849_1;
buffer_wire buffer_9849_1 (.in(n9849_0), .out(n9849_1));
wire n9850; //CHANX 4 (6,0) #50
wire n9850_0;
wire n9850_1;
buffer_wire buffer_9850_1 (.in(n9850_0), .out(n9850_1));
wire n9851; //CHANX 4 (6,0) #51
wire n9851_0;
wire n9851_1;
buffer_wire buffer_9851_1 (.in(n9851_0), .out(n9851_1));
wire n9852; //CHANX 4 (6,0) #58
wire n9852_0;
wire n9852_1;
buffer_wire buffer_9852_1 (.in(n9852_0), .out(n9852_1));
wire n9853; //CHANX 4 (6,0) #59
wire n9853_0;
wire n9853_1;
buffer_wire buffer_9853_1 (.in(n9853_0), .out(n9853_1));
wire n9854; //CHANX 4 (6,0) #66
wire n9854_0;
wire n9854_1;
buffer_wire buffer_9854_1 (.in(n9854_0), .out(n9854_1));
wire n9855; //CHANX 4 (6,0) #67
wire n9855_0;
wire n9855_1;
buffer_wire buffer_9855_1 (.in(n9855_0), .out(n9855_1));
wire n9856; //CHANX 4 (6,0) #74
wire n9856_0;
wire n9856_1;
buffer_wire buffer_9856_1 (.in(n9856_0), .out(n9856_1));
wire n9857; //CHANX 4 (6,0) #75
wire n9857_0;
wire n9857_1;
buffer_wire buffer_9857_1 (.in(n9857_0), .out(n9857_1));
wire n9858; //CHANX 3 (7,0) #4
wire n9858_0;
wire n9859; //CHANX 3 (7,0) #5
wire n9859_0;
wire n9860; //CHANX 3 (7,0) #12
wire n9860_0;
wire n9861; //CHANX 3 (7,0) #13
wire n9861_0;
wire n9862; //CHANX 3 (7,0) #20
wire n9862_0;
wire n9863; //CHANX 3 (7,0) #21
wire n9863_0;
wire n9864; //CHANX 3 (7,0) #28
wire n9864_0;
wire n9865; //CHANX 3 (7,0) #29
wire n9865_0;
wire n9866; //CHANX 3 (7,0) #36
wire n9866_0;
wire n9867; //CHANX 3 (7,0) #37
wire n9867_0;
wire n9868; //CHANX 3 (7,0) #44
wire n9868_0;
wire n9869; //CHANX 3 (7,0) #45
wire n9869_0;
wire n9870; //CHANX 3 (7,0) #52
wire n9870_0;
wire n9871; //CHANX 3 (7,0) #53
wire n9871_0;
wire n9872; //CHANX 3 (7,0) #60
wire n9872_0;
wire n9873; //CHANX 3 (7,0) #61
wire n9873_0;
wire n9874; //CHANX 3 (7,0) #68
wire n9874_0;
wire n9875; //CHANX 3 (7,0) #69
wire n9875_0;
wire n9876; //CHANX 3 (7,0) #76
wire n9876_0;
wire n9877; //CHANX 3 (7,0) #77
wire n9877_0;
wire n9878; //CHANX 2 (8,0) #6
wire n9878_0;
wire n9879; //CHANX 2 (8,0) #7
wire n9879_0;
wire n9880; //CHANX 2 (8,0) #14
wire n9880_0;
wire n9881; //CHANX 2 (8,0) #15
wire n9881_0;
wire n9882; //CHANX 2 (8,0) #22
wire n9882_0;
wire n9883; //CHANX 2 (8,0) #23
wire n9883_0;
wire n9884; //CHANX 2 (8,0) #30
wire n9884_0;
wire n9885; //CHANX 2 (8,0) #31
wire n9885_0;
wire n9886; //CHANX 2 (8,0) #38
wire n9886_0;
wire n9887; //CHANX 2 (8,0) #39
wire n9887_0;
wire n9888; //CHANX 2 (8,0) #46
wire n9888_0;
wire n9889; //CHANX 2 (8,0) #47
wire n9889_0;
wire n9890; //CHANX 2 (8,0) #54
wire n9890_0;
wire n9891; //CHANX 2 (8,0) #55
wire n9891_0;
wire n9892; //CHANX 2 (8,0) #62
wire n9892_0;
wire n9893; //CHANX 2 (8,0) #63
wire n9893_0;
wire n9894; //CHANX 2 (8,0) #70
wire n9894_0;
wire n9895; //CHANX 2 (8,0) #71
wire n9895_0;
wire n9896; //CHANX 2 (8,0) #78
wire n9896_0;
wire n9897; //CHANX 2 (8,0) #79
wire n9897_0;
wire n9898; //CHANX 1 (9,0) #0
wire n9898_0;
wire n9899; //CHANX 1 (9,0) #1
wire n9899_0;
wire n9900; //CHANX 1 (9,0) #8
wire n9900_0;
wire n9901; //CHANX 1 (9,0) #9
wire n9901_0;
wire n9902; //CHANX 1 (9,0) #16
wire n9902_0;
wire n9903; //CHANX 1 (9,0) #17
wire n9903_0;
wire n9904; //CHANX 1 (9,0) #24
wire n9904_0;
wire n9905; //CHANX 1 (9,0) #25
wire n9905_0;
wire n9906; //CHANX 1 (9,0) #32
wire n9906_0;
wire n9907; //CHANX 1 (9,0) #33
wire n9907_0;
wire n9908; //CHANX 1 (9,0) #40
wire n9908_0;
wire n9909; //CHANX 1 (9,0) #41
wire n9909_0;
wire n9910; //CHANX 1 (9,0) #48
wire n9910_0;
wire n9911; //CHANX 1 (9,0) #49
wire n9911_0;
wire n9912; //CHANX 1 (9,0) #56
wire n9912_0;
wire n9913; //CHANX 1 (9,0) #57
wire n9913_0;
wire n9914; //CHANX 1 (9,0) #64
wire n9914_0;
wire n9915; //CHANX 1 (9,0) #65
wire n9915_0;
wire n9916; //CHANX 1 (9,0) #72
wire n9916_0;
wire n9917; //CHANX 1 (9,0) #73
wire n9917_0;
wire n9918; //CHANX 1 (9,0) #80
wire n9918_0;
wire n9919; //CHANX 1 (9,0) #81
wire n9919_0;
wire n9920; //CHANX 3 (1,1) #0
wire n9920_0;
wire n9921; //CHANX 3 (1,1) #1
wire n9921_0;
wire n9922; //CHANX 4 (1,1) #2
wire n9922_0;
wire n9922_1;
buffer_wire buffer_9922_1 (.in(n9922_0), .out(n9922_1));
wire n9923; //CHANX 4 (1,1) #3
wire n9923_0;
wire n9923_1;
buffer_wire buffer_9923_1 (.in(n9923_0), .out(n9923_1));
wire n9924; //CHANX 1 (1,1) #4
wire n9924_0;
wire n9925; //CHANX 1 (1,1) #5
wire n9925_0;
wire n9926; //CHANX 2 (1,1) #6
wire n9926_0;
wire n9927; //CHANX 2 (1,1) #7
wire n9927_0;
wire n9928; //CHANX 3 (1,1) #8
wire n9928_0;
wire n9929; //CHANX 3 (1,1) #9
wire n9929_0;
wire n9930; //CHANX 4 (1,1) #10
wire n9930_0;
wire n9930_1;
buffer_wire buffer_9930_1 (.in(n9930_0), .out(n9930_1));
wire n9931; //CHANX 4 (1,1) #11
wire n9931_0;
wire n9931_1;
buffer_wire buffer_9931_1 (.in(n9931_0), .out(n9931_1));
wire n9932; //CHANX 1 (1,1) #12
wire n9932_0;
wire n9933; //CHANX 1 (1,1) #13
wire n9933_0;
wire n9934; //CHANX 2 (1,1) #14
wire n9934_0;
wire n9935; //CHANX 2 (1,1) #15
wire n9935_0;
wire n9936; //CHANX 3 (1,1) #16
wire n9936_0;
wire n9937; //CHANX 3 (1,1) #17
wire n9937_0;
wire n9938; //CHANX 4 (1,1) #18
wire n9938_0;
wire n9938_1;
buffer_wire buffer_9938_1 (.in(n9938_0), .out(n9938_1));
wire n9939; //CHANX 4 (1,1) #19
wire n9939_0;
wire n9939_1;
buffer_wire buffer_9939_1 (.in(n9939_0), .out(n9939_1));
wire n9940; //CHANX 1 (1,1) #20
wire n9940_0;
wire n9941; //CHANX 1 (1,1) #21
wire n9941_0;
wire n9942; //CHANX 2 (1,1) #22
wire n9942_0;
wire n9943; //CHANX 2 (1,1) #23
wire n9943_0;
wire n9944; //CHANX 3 (1,1) #24
wire n9944_0;
wire n9945; //CHANX 3 (1,1) #25
wire n9945_0;
wire n9946; //CHANX 4 (1,1) #26
wire n9946_0;
wire n9946_1;
buffer_wire buffer_9946_1 (.in(n9946_0), .out(n9946_1));
wire n9947; //CHANX 4 (1,1) #27
wire n9947_0;
wire n9947_1;
buffer_wire buffer_9947_1 (.in(n9947_0), .out(n9947_1));
wire n9948; //CHANX 1 (1,1) #28
wire n9948_0;
wire n9949; //CHANX 1 (1,1) #29
wire n9949_0;
wire n9950; //CHANX 2 (1,1) #30
wire n9950_0;
wire n9951; //CHANX 2 (1,1) #31
wire n9951_0;
wire n9952; //CHANX 3 (1,1) #32
wire n9952_0;
wire n9953; //CHANX 3 (1,1) #33
wire n9953_0;
wire n9954; //CHANX 4 (1,1) #34
wire n9954_0;
wire n9954_1;
buffer_wire buffer_9954_1 (.in(n9954_0), .out(n9954_1));
wire n9955; //CHANX 4 (1,1) #35
wire n9955_0;
wire n9955_1;
buffer_wire buffer_9955_1 (.in(n9955_0), .out(n9955_1));
wire n9956; //CHANX 1 (1,1) #36
wire n9956_0;
wire n9957; //CHANX 1 (1,1) #37
wire n9957_0;
wire n9958; //CHANX 2 (1,1) #38
wire n9958_0;
wire n9959; //CHANX 2 (1,1) #39
wire n9959_0;
wire n9960; //CHANX 3 (1,1) #40
wire n9960_0;
wire n9961; //CHANX 3 (1,1) #41
wire n9961_0;
wire n9962; //CHANX 4 (1,1) #42
wire n9962_0;
wire n9962_1;
buffer_wire buffer_9962_1 (.in(n9962_0), .out(n9962_1));
wire n9963; //CHANX 4 (1,1) #43
wire n9963_0;
wire n9963_1;
buffer_wire buffer_9963_1 (.in(n9963_0), .out(n9963_1));
wire n9964; //CHANX 1 (1,1) #44
wire n9964_0;
wire n9965; //CHANX 1 (1,1) #45
wire n9965_0;
wire n9966; //CHANX 2 (1,1) #46
wire n9966_0;
wire n9967; //CHANX 2 (1,1) #47
wire n9967_0;
wire n9968; //CHANX 3 (1,1) #48
wire n9968_0;
wire n9969; //CHANX 3 (1,1) #49
wire n9969_0;
wire n9970; //CHANX 4 (1,1) #50
wire n9970_0;
wire n9970_1;
buffer_wire buffer_9970_1 (.in(n9970_0), .out(n9970_1));
wire n9971; //CHANX 4 (1,1) #51
wire n9971_0;
wire n9971_1;
buffer_wire buffer_9971_1 (.in(n9971_0), .out(n9971_1));
wire n9972; //CHANX 1 (1,1) #52
wire n9972_0;
wire n9973; //CHANX 1 (1,1) #53
wire n9973_0;
wire n9974; //CHANX 2 (1,1) #54
wire n9974_0;
wire n9975; //CHANX 2 (1,1) #55
wire n9975_0;
wire n9976; //CHANX 3 (1,1) #56
wire n9976_0;
wire n9977; //CHANX 3 (1,1) #57
wire n9977_0;
wire n9978; //CHANX 4 (1,1) #58
wire n9978_0;
wire n9978_1;
buffer_wire buffer_9978_1 (.in(n9978_0), .out(n9978_1));
wire n9979; //CHANX 4 (1,1) #59
wire n9979_0;
wire n9979_1;
buffer_wire buffer_9979_1 (.in(n9979_0), .out(n9979_1));
wire n9980; //CHANX 1 (1,1) #60
wire n9980_0;
wire n9981; //CHANX 1 (1,1) #61
wire n9981_0;
wire n9982; //CHANX 2 (1,1) #62
wire n9982_0;
wire n9983; //CHANX 2 (1,1) #63
wire n9983_0;
wire n9984; //CHANX 3 (1,1) #64
wire n9984_0;
wire n9985; //CHANX 3 (1,1) #65
wire n9985_0;
wire n9986; //CHANX 4 (1,1) #66
wire n9986_0;
wire n9986_1;
buffer_wire buffer_9986_1 (.in(n9986_0), .out(n9986_1));
wire n9987; //CHANX 4 (1,1) #67
wire n9987_0;
wire n9987_1;
buffer_wire buffer_9987_1 (.in(n9987_0), .out(n9987_1));
wire n9988; //CHANX 1 (1,1) #68
wire n9988_0;
wire n9989; //CHANX 1 (1,1) #69
wire n9989_0;
wire n9990; //CHANX 2 (1,1) #70
wire n9990_0;
wire n9991; //CHANX 2 (1,1) #71
wire n9991_0;
wire n9992; //CHANX 3 (1,1) #72
wire n9992_0;
wire n9993; //CHANX 3 (1,1) #73
wire n9993_0;
wire n9994; //CHANX 4 (1,1) #74
wire n9994_0;
wire n9994_1;
buffer_wire buffer_9994_1 (.in(n9994_0), .out(n9994_1));
wire n9995; //CHANX 4 (1,1) #75
wire n9995_0;
wire n9995_1;
buffer_wire buffer_9995_1 (.in(n9995_0), .out(n9995_1));
wire n9996; //CHANX 1 (1,1) #76
wire n9996_0;
wire n9997; //CHANX 1 (1,1) #77
wire n9997_0;
wire n9998; //CHANX 2 (1,1) #78
wire n9998_0;
wire n9999; //CHANX 2 (1,1) #79
wire n9999_0;
wire n10000; //CHANX 7 (1,1) #80
wire n10000_0;
wire n10000_1;
wire n10000_2;
buffer_wire buffer_10000_2 (.in(n10000_1), .out(n10000_2));
buffer_wire buffer_10000_1 (.in(n10000_0), .out(n10000_1));
wire n10001; //CHANX 7 (1,1) #81
wire n10001_0;
wire n10001_1;
wire n10001_2;
buffer_wire buffer_10001_2 (.in(n10001_1), .out(n10001_2));
buffer_wire buffer_10001_1 (.in(n10001_0), .out(n10001_1));
wire n10002; //CHANX 8 (1,1) #82
wire n10002_0;
wire n10002_1;
wire n10002_2;
buffer_wire buffer_10002_2 (.in(n10002_1), .out(n10002_2));
buffer_wire buffer_10002_1 (.in(n10002_0), .out(n10002_1));
wire n10003; //CHANX 8 (1,1) #83
wire n10003_0;
wire n10003_1;
wire n10003_2;
buffer_wire buffer_10003_2 (.in(n10003_1), .out(n10003_2));
buffer_wire buffer_10003_1 (.in(n10003_0), .out(n10003_1));
wire n10004; //CHANX 9 (1,1) #84
wire n10004_0;
wire n10004_1;
wire n10004_2;
buffer_wire buffer_10004_2 (.in(n10004_1), .out(n10004_2));
buffer_wire buffer_10004_1 (.in(n10004_0), .out(n10004_1));
wire n10005; //CHANX 9 (1,1) #85
wire n10005_0;
wire n10005_1;
wire n10005_2;
buffer_wire buffer_10005_2 (.in(n10005_1), .out(n10005_2));
buffer_wire buffer_10005_1 (.in(n10005_0), .out(n10005_1));
wire n10006; //CHANX 9 (1,1) #86
wire n10006_0;
wire n10006_1;
wire n10006_2;
buffer_wire buffer_10006_2 (.in(n10006_1), .out(n10006_2));
buffer_wire buffer_10006_1 (.in(n10006_0), .out(n10006_1));
wire n10007; //CHANX 9 (1,1) #87
wire n10007_0;
wire n10007_1;
wire n10007_2;
buffer_wire buffer_10007_2 (.in(n10007_1), .out(n10007_2));
buffer_wire buffer_10007_1 (.in(n10007_0), .out(n10007_1));
wire n10008; //CHANX 9 (1,1) #88
wire n10008_0;
wire n10008_1;
wire n10008_2;
buffer_wire buffer_10008_2 (.in(n10008_1), .out(n10008_2));
buffer_wire buffer_10008_1 (.in(n10008_0), .out(n10008_1));
wire n10009; //CHANX 9 (1,1) #89
wire n10009_0;
wire n10009_1;
wire n10009_2;
buffer_wire buffer_10009_2 (.in(n10009_1), .out(n10009_2));
buffer_wire buffer_10009_1 (.in(n10009_0), .out(n10009_1));
wire n10010; //CHANX 9 (1,1) #90
wire n10010_0;
wire n10010_1;
wire n10010_2;
buffer_wire buffer_10010_2 (.in(n10010_1), .out(n10010_2));
buffer_wire buffer_10010_1 (.in(n10010_0), .out(n10010_1));
wire n10011; //CHANX 9 (1,1) #91
wire n10011_0;
wire n10011_1;
wire n10011_2;
buffer_wire buffer_10011_2 (.in(n10011_1), .out(n10011_2));
buffer_wire buffer_10011_1 (.in(n10011_0), .out(n10011_1));
wire n10012; //CHANX 4 (2,1) #4
wire n10012_0;
wire n10012_1;
buffer_wire buffer_10012_1 (.in(n10012_0), .out(n10012_1));
wire n10013; //CHANX 4 (2,1) #5
wire n10013_0;
wire n10013_1;
buffer_wire buffer_10013_1 (.in(n10013_0), .out(n10013_1));
wire n10014; //CHANX 4 (2,1) #12
wire n10014_0;
wire n10014_1;
buffer_wire buffer_10014_1 (.in(n10014_0), .out(n10014_1));
wire n10015; //CHANX 4 (2,1) #13
wire n10015_0;
wire n10015_1;
buffer_wire buffer_10015_1 (.in(n10015_0), .out(n10015_1));
wire n10016; //CHANX 4 (2,1) #20
wire n10016_0;
wire n10016_1;
buffer_wire buffer_10016_1 (.in(n10016_0), .out(n10016_1));
wire n10017; //CHANX 4 (2,1) #21
wire n10017_0;
wire n10017_1;
buffer_wire buffer_10017_1 (.in(n10017_0), .out(n10017_1));
wire n10018; //CHANX 4 (2,1) #28
wire n10018_0;
wire n10018_1;
buffer_wire buffer_10018_1 (.in(n10018_0), .out(n10018_1));
wire n10019; //CHANX 4 (2,1) #29
wire n10019_0;
wire n10019_1;
buffer_wire buffer_10019_1 (.in(n10019_0), .out(n10019_1));
wire n10020; //CHANX 4 (2,1) #36
wire n10020_0;
wire n10020_1;
buffer_wire buffer_10020_1 (.in(n10020_0), .out(n10020_1));
wire n10021; //CHANX 4 (2,1) #37
wire n10021_0;
wire n10021_1;
buffer_wire buffer_10021_1 (.in(n10021_0), .out(n10021_1));
wire n10022; //CHANX 4 (2,1) #44
wire n10022_0;
wire n10022_1;
buffer_wire buffer_10022_1 (.in(n10022_0), .out(n10022_1));
wire n10023; //CHANX 4 (2,1) #45
wire n10023_0;
wire n10023_1;
buffer_wire buffer_10023_1 (.in(n10023_0), .out(n10023_1));
wire n10024; //CHANX 4 (2,1) #52
wire n10024_0;
wire n10024_1;
buffer_wire buffer_10024_1 (.in(n10024_0), .out(n10024_1));
wire n10025; //CHANX 4 (2,1) #53
wire n10025_0;
wire n10025_1;
buffer_wire buffer_10025_1 (.in(n10025_0), .out(n10025_1));
wire n10026; //CHANX 4 (2,1) #60
wire n10026_0;
wire n10026_1;
buffer_wire buffer_10026_1 (.in(n10026_0), .out(n10026_1));
wire n10027; //CHANX 4 (2,1) #61
wire n10027_0;
wire n10027_1;
buffer_wire buffer_10027_1 (.in(n10027_0), .out(n10027_1));
wire n10028; //CHANX 4 (2,1) #68
wire n10028_0;
wire n10028_1;
buffer_wire buffer_10028_1 (.in(n10028_0), .out(n10028_1));
wire n10029; //CHANX 4 (2,1) #69
wire n10029_0;
wire n10029_1;
buffer_wire buffer_10029_1 (.in(n10029_0), .out(n10029_1));
wire n10030; //CHANX 4 (2,1) #76
wire n10030_0;
wire n10030_1;
buffer_wire buffer_10030_1 (.in(n10030_0), .out(n10030_1));
wire n10031; //CHANX 4 (2,1) #77
wire n10031_0;
wire n10031_1;
buffer_wire buffer_10031_1 (.in(n10031_0), .out(n10031_1));
wire n10032; //CHANX 4 (3,1) #6
wire n10032_0;
wire n10032_1;
buffer_wire buffer_10032_1 (.in(n10032_0), .out(n10032_1));
wire n10033; //CHANX 4 (3,1) #7
wire n10033_0;
wire n10033_1;
buffer_wire buffer_10033_1 (.in(n10033_0), .out(n10033_1));
wire n10034; //CHANX 4 (3,1) #14
wire n10034_0;
wire n10034_1;
buffer_wire buffer_10034_1 (.in(n10034_0), .out(n10034_1));
wire n10035; //CHANX 4 (3,1) #15
wire n10035_0;
wire n10035_1;
buffer_wire buffer_10035_1 (.in(n10035_0), .out(n10035_1));
wire n10036; //CHANX 4 (3,1) #22
wire n10036_0;
wire n10036_1;
buffer_wire buffer_10036_1 (.in(n10036_0), .out(n10036_1));
wire n10037; //CHANX 4 (3,1) #23
wire n10037_0;
wire n10037_1;
buffer_wire buffer_10037_1 (.in(n10037_0), .out(n10037_1));
wire n10038; //CHANX 4 (3,1) #30
wire n10038_0;
wire n10038_1;
buffer_wire buffer_10038_1 (.in(n10038_0), .out(n10038_1));
wire n10039; //CHANX 4 (3,1) #31
wire n10039_0;
wire n10039_1;
buffer_wire buffer_10039_1 (.in(n10039_0), .out(n10039_1));
wire n10040; //CHANX 4 (3,1) #38
wire n10040_0;
wire n10040_1;
buffer_wire buffer_10040_1 (.in(n10040_0), .out(n10040_1));
wire n10041; //CHANX 4 (3,1) #39
wire n10041_0;
wire n10041_1;
buffer_wire buffer_10041_1 (.in(n10041_0), .out(n10041_1));
wire n10042; //CHANX 4 (3,1) #46
wire n10042_0;
wire n10042_1;
buffer_wire buffer_10042_1 (.in(n10042_0), .out(n10042_1));
wire n10043; //CHANX 4 (3,1) #47
wire n10043_0;
wire n10043_1;
buffer_wire buffer_10043_1 (.in(n10043_0), .out(n10043_1));
wire n10044; //CHANX 4 (3,1) #54
wire n10044_0;
wire n10044_1;
buffer_wire buffer_10044_1 (.in(n10044_0), .out(n10044_1));
wire n10045; //CHANX 4 (3,1) #55
wire n10045_0;
wire n10045_1;
buffer_wire buffer_10045_1 (.in(n10045_0), .out(n10045_1));
wire n10046; //CHANX 4 (3,1) #62
wire n10046_0;
wire n10046_1;
buffer_wire buffer_10046_1 (.in(n10046_0), .out(n10046_1));
wire n10047; //CHANX 4 (3,1) #63
wire n10047_0;
wire n10047_1;
buffer_wire buffer_10047_1 (.in(n10047_0), .out(n10047_1));
wire n10048; //CHANX 4 (3,1) #70
wire n10048_0;
wire n10048_1;
buffer_wire buffer_10048_1 (.in(n10048_0), .out(n10048_1));
wire n10049; //CHANX 4 (3,1) #71
wire n10049_0;
wire n10049_1;
buffer_wire buffer_10049_1 (.in(n10049_0), .out(n10049_1));
wire n10050; //CHANX 4 (3,1) #78
wire n10050_0;
wire n10050_1;
buffer_wire buffer_10050_1 (.in(n10050_0), .out(n10050_1));
wire n10051; //CHANX 4 (3,1) #79
wire n10051_0;
wire n10051_1;
buffer_wire buffer_10051_1 (.in(n10051_0), .out(n10051_1));
wire n10052; //CHANX 4 (4,1) #0
wire n10052_0;
wire n10052_1;
buffer_wire buffer_10052_1 (.in(n10052_0), .out(n10052_1));
wire n10053; //CHANX 4 (4,1) #1
wire n10053_0;
wire n10053_1;
buffer_wire buffer_10053_1 (.in(n10053_0), .out(n10053_1));
wire n10054; //CHANX 4 (4,1) #8
wire n10054_0;
wire n10054_1;
buffer_wire buffer_10054_1 (.in(n10054_0), .out(n10054_1));
wire n10055; //CHANX 4 (4,1) #9
wire n10055_0;
wire n10055_1;
buffer_wire buffer_10055_1 (.in(n10055_0), .out(n10055_1));
wire n10056; //CHANX 4 (4,1) #16
wire n10056_0;
wire n10056_1;
buffer_wire buffer_10056_1 (.in(n10056_0), .out(n10056_1));
wire n10057; //CHANX 4 (4,1) #17
wire n10057_0;
wire n10057_1;
buffer_wire buffer_10057_1 (.in(n10057_0), .out(n10057_1));
wire n10058; //CHANX 4 (4,1) #24
wire n10058_0;
wire n10058_1;
buffer_wire buffer_10058_1 (.in(n10058_0), .out(n10058_1));
wire n10059; //CHANX 4 (4,1) #25
wire n10059_0;
wire n10059_1;
buffer_wire buffer_10059_1 (.in(n10059_0), .out(n10059_1));
wire n10060; //CHANX 4 (4,1) #32
wire n10060_0;
wire n10060_1;
buffer_wire buffer_10060_1 (.in(n10060_0), .out(n10060_1));
wire n10061; //CHANX 4 (4,1) #33
wire n10061_0;
wire n10061_1;
buffer_wire buffer_10061_1 (.in(n10061_0), .out(n10061_1));
wire n10062; //CHANX 4 (4,1) #40
wire n10062_0;
wire n10062_1;
buffer_wire buffer_10062_1 (.in(n10062_0), .out(n10062_1));
wire n10063; //CHANX 4 (4,1) #41
wire n10063_0;
wire n10063_1;
buffer_wire buffer_10063_1 (.in(n10063_0), .out(n10063_1));
wire n10064; //CHANX 4 (4,1) #48
wire n10064_0;
wire n10064_1;
buffer_wire buffer_10064_1 (.in(n10064_0), .out(n10064_1));
wire n10065; //CHANX 4 (4,1) #49
wire n10065_0;
wire n10065_1;
buffer_wire buffer_10065_1 (.in(n10065_0), .out(n10065_1));
wire n10066; //CHANX 4 (4,1) #56
wire n10066_0;
wire n10066_1;
buffer_wire buffer_10066_1 (.in(n10066_0), .out(n10066_1));
wire n10067; //CHANX 4 (4,1) #57
wire n10067_0;
wire n10067_1;
buffer_wire buffer_10067_1 (.in(n10067_0), .out(n10067_1));
wire n10068; //CHANX 4 (4,1) #64
wire n10068_0;
wire n10068_1;
buffer_wire buffer_10068_1 (.in(n10068_0), .out(n10068_1));
wire n10069; //CHANX 4 (4,1) #65
wire n10069_0;
wire n10069_1;
buffer_wire buffer_10069_1 (.in(n10069_0), .out(n10069_1));
wire n10070; //CHANX 4 (4,1) #72
wire n10070_0;
wire n10070_1;
buffer_wire buffer_10070_1 (.in(n10070_0), .out(n10070_1));
wire n10071; //CHANX 4 (4,1) #73
wire n10071_0;
wire n10071_1;
buffer_wire buffer_10071_1 (.in(n10071_0), .out(n10071_1));
wire n10072; //CHANX 4 (5,1) #2
wire n10072_0;
wire n10072_1;
buffer_wire buffer_10072_1 (.in(n10072_0), .out(n10072_1));
wire n10073; //CHANX 4 (5,1) #3
wire n10073_0;
wire n10073_1;
buffer_wire buffer_10073_1 (.in(n10073_0), .out(n10073_1));
wire n10074; //CHANX 4 (5,1) #10
wire n10074_0;
wire n10074_1;
buffer_wire buffer_10074_1 (.in(n10074_0), .out(n10074_1));
wire n10075; //CHANX 4 (5,1) #11
wire n10075_0;
wire n10075_1;
buffer_wire buffer_10075_1 (.in(n10075_0), .out(n10075_1));
wire n10076; //CHANX 4 (5,1) #18
wire n10076_0;
wire n10076_1;
buffer_wire buffer_10076_1 (.in(n10076_0), .out(n10076_1));
wire n10077; //CHANX 4 (5,1) #19
wire n10077_0;
wire n10077_1;
buffer_wire buffer_10077_1 (.in(n10077_0), .out(n10077_1));
wire n10078; //CHANX 4 (5,1) #26
wire n10078_0;
wire n10078_1;
buffer_wire buffer_10078_1 (.in(n10078_0), .out(n10078_1));
wire n10079; //CHANX 4 (5,1) #27
wire n10079_0;
wire n10079_1;
buffer_wire buffer_10079_1 (.in(n10079_0), .out(n10079_1));
wire n10080; //CHANX 4 (5,1) #34
wire n10080_0;
wire n10080_1;
buffer_wire buffer_10080_1 (.in(n10080_0), .out(n10080_1));
wire n10081; //CHANX 4 (5,1) #35
wire n10081_0;
wire n10081_1;
buffer_wire buffer_10081_1 (.in(n10081_0), .out(n10081_1));
wire n10082; //CHANX 4 (5,1) #42
wire n10082_0;
wire n10082_1;
buffer_wire buffer_10082_1 (.in(n10082_0), .out(n10082_1));
wire n10083; //CHANX 4 (5,1) #43
wire n10083_0;
wire n10083_1;
buffer_wire buffer_10083_1 (.in(n10083_0), .out(n10083_1));
wire n10084; //CHANX 4 (5,1) #50
wire n10084_0;
wire n10084_1;
buffer_wire buffer_10084_1 (.in(n10084_0), .out(n10084_1));
wire n10085; //CHANX 4 (5,1) #51
wire n10085_0;
wire n10085_1;
buffer_wire buffer_10085_1 (.in(n10085_0), .out(n10085_1));
wire n10086; //CHANX 4 (5,1) #58
wire n10086_0;
wire n10086_1;
buffer_wire buffer_10086_1 (.in(n10086_0), .out(n10086_1));
wire n10087; //CHANX 4 (5,1) #59
wire n10087_0;
wire n10087_1;
buffer_wire buffer_10087_1 (.in(n10087_0), .out(n10087_1));
wire n10088; //CHANX 4 (5,1) #66
wire n10088_0;
wire n10088_1;
buffer_wire buffer_10088_1 (.in(n10088_0), .out(n10088_1));
wire n10089; //CHANX 4 (5,1) #67
wire n10089_0;
wire n10089_1;
buffer_wire buffer_10089_1 (.in(n10089_0), .out(n10089_1));
wire n10090; //CHANX 4 (5,1) #74
wire n10090_0;
wire n10090_1;
buffer_wire buffer_10090_1 (.in(n10090_0), .out(n10090_1));
wire n10091; //CHANX 4 (5,1) #75
wire n10091_0;
wire n10091_1;
buffer_wire buffer_10091_1 (.in(n10091_0), .out(n10091_1));
wire n10092; //CHANX 4 (6,1) #4
wire n10092_0;
wire n10092_1;
buffer_wire buffer_10092_1 (.in(n10092_0), .out(n10092_1));
wire n10093; //CHANX 4 (6,1) #5
wire n10093_0;
wire n10093_1;
buffer_wire buffer_10093_1 (.in(n10093_0), .out(n10093_1));
wire n10094; //CHANX 4 (6,1) #12
wire n10094_0;
wire n10094_1;
buffer_wire buffer_10094_1 (.in(n10094_0), .out(n10094_1));
wire n10095; //CHANX 4 (6,1) #13
wire n10095_0;
wire n10095_1;
buffer_wire buffer_10095_1 (.in(n10095_0), .out(n10095_1));
wire n10096; //CHANX 4 (6,1) #20
wire n10096_0;
wire n10096_1;
buffer_wire buffer_10096_1 (.in(n10096_0), .out(n10096_1));
wire n10097; //CHANX 4 (6,1) #21
wire n10097_0;
wire n10097_1;
buffer_wire buffer_10097_1 (.in(n10097_0), .out(n10097_1));
wire n10098; //CHANX 4 (6,1) #28
wire n10098_0;
wire n10098_1;
buffer_wire buffer_10098_1 (.in(n10098_0), .out(n10098_1));
wire n10099; //CHANX 4 (6,1) #29
wire n10099_0;
wire n10099_1;
buffer_wire buffer_10099_1 (.in(n10099_0), .out(n10099_1));
wire n10100; //CHANX 4 (6,1) #36
wire n10100_0;
wire n10100_1;
buffer_wire buffer_10100_1 (.in(n10100_0), .out(n10100_1));
wire n10101; //CHANX 4 (6,1) #37
wire n10101_0;
wire n10101_1;
buffer_wire buffer_10101_1 (.in(n10101_0), .out(n10101_1));
wire n10102; //CHANX 4 (6,1) #44
wire n10102_0;
wire n10102_1;
buffer_wire buffer_10102_1 (.in(n10102_0), .out(n10102_1));
wire n10103; //CHANX 4 (6,1) #45
wire n10103_0;
wire n10103_1;
buffer_wire buffer_10103_1 (.in(n10103_0), .out(n10103_1));
wire n10104; //CHANX 4 (6,1) #52
wire n10104_0;
wire n10104_1;
buffer_wire buffer_10104_1 (.in(n10104_0), .out(n10104_1));
wire n10105; //CHANX 4 (6,1) #53
wire n10105_0;
wire n10105_1;
buffer_wire buffer_10105_1 (.in(n10105_0), .out(n10105_1));
wire n10106; //CHANX 4 (6,1) #60
wire n10106_0;
wire n10106_1;
buffer_wire buffer_10106_1 (.in(n10106_0), .out(n10106_1));
wire n10107; //CHANX 4 (6,1) #61
wire n10107_0;
wire n10107_1;
buffer_wire buffer_10107_1 (.in(n10107_0), .out(n10107_1));
wire n10108; //CHANX 4 (6,1) #68
wire n10108_0;
wire n10108_1;
buffer_wire buffer_10108_1 (.in(n10108_0), .out(n10108_1));
wire n10109; //CHANX 4 (6,1) #69
wire n10109_0;
wire n10109_1;
buffer_wire buffer_10109_1 (.in(n10109_0), .out(n10109_1));
wire n10110; //CHANX 4 (6,1) #76
wire n10110_0;
wire n10110_1;
buffer_wire buffer_10110_1 (.in(n10110_0), .out(n10110_1));
wire n10111; //CHANX 4 (6,1) #77
wire n10111_0;
wire n10111_1;
buffer_wire buffer_10111_1 (.in(n10111_0), .out(n10111_1));
wire n10112; //CHANX 3 (7,1) #6
wire n10112_0;
wire n10113; //CHANX 3 (7,1) #7
wire n10113_0;
wire n10114; //CHANX 3 (7,1) #14
wire n10114_0;
wire n10115; //CHANX 3 (7,1) #15
wire n10115_0;
wire n10116; //CHANX 3 (7,1) #22
wire n10116_0;
wire n10117; //CHANX 3 (7,1) #23
wire n10117_0;
wire n10118; //CHANX 3 (7,1) #30
wire n10118_0;
wire n10119; //CHANX 3 (7,1) #31
wire n10119_0;
wire n10120; //CHANX 3 (7,1) #38
wire n10120_0;
wire n10121; //CHANX 3 (7,1) #39
wire n10121_0;
wire n10122; //CHANX 3 (7,1) #46
wire n10122_0;
wire n10123; //CHANX 3 (7,1) #47
wire n10123_0;
wire n10124; //CHANX 3 (7,1) #54
wire n10124_0;
wire n10125; //CHANX 3 (7,1) #55
wire n10125_0;
wire n10126; //CHANX 3 (7,1) #62
wire n10126_0;
wire n10127; //CHANX 3 (7,1) #63
wire n10127_0;
wire n10128; //CHANX 3 (7,1) #70
wire n10128_0;
wire n10129; //CHANX 3 (7,1) #71
wire n10129_0;
wire n10130; //CHANX 3 (7,1) #78
wire n10130_0;
wire n10131; //CHANX 3 (7,1) #79
wire n10131_0;
wire n10132; //CHANX 2 (8,1) #0
wire n10132_0;
wire n10133; //CHANX 2 (8,1) #1
wire n10133_0;
wire n10134; //CHANX 2 (8,1) #8
wire n10134_0;
wire n10135; //CHANX 2 (8,1) #9
wire n10135_0;
wire n10136; //CHANX 2 (8,1) #16
wire n10136_0;
wire n10137; //CHANX 2 (8,1) #17
wire n10137_0;
wire n10138; //CHANX 2 (8,1) #24
wire n10138_0;
wire n10139; //CHANX 2 (8,1) #25
wire n10139_0;
wire n10140; //CHANX 2 (8,1) #32
wire n10140_0;
wire n10141; //CHANX 2 (8,1) #33
wire n10141_0;
wire n10142; //CHANX 2 (8,1) #40
wire n10142_0;
wire n10143; //CHANX 2 (8,1) #41
wire n10143_0;
wire n10144; //CHANX 2 (8,1) #48
wire n10144_0;
wire n10145; //CHANX 2 (8,1) #49
wire n10145_0;
wire n10146; //CHANX 2 (8,1) #56
wire n10146_0;
wire n10147; //CHANX 2 (8,1) #57
wire n10147_0;
wire n10148; //CHANX 2 (8,1) #64
wire n10148_0;
wire n10149; //CHANX 2 (8,1) #65
wire n10149_0;
wire n10150; //CHANX 2 (8,1) #72
wire n10150_0;
wire n10151; //CHANX 2 (8,1) #73
wire n10151_0;
wire n10152; //CHANX 2 (8,1) #80
wire n10152_0;
wire n10153; //CHANX 2 (8,1) #81
wire n10153_0;
wire n10154; //CHANX 1 (9,1) #2
wire n10154_0;
wire n10155; //CHANX 1 (9,1) #3
wire n10155_0;
wire n10156; //CHANX 1 (9,1) #10
wire n10156_0;
wire n10157; //CHANX 1 (9,1) #11
wire n10157_0;
wire n10158; //CHANX 1 (9,1) #18
wire n10158_0;
wire n10159; //CHANX 1 (9,1) #19
wire n10159_0;
wire n10160; //CHANX 1 (9,1) #26
wire n10160_0;
wire n10161; //CHANX 1 (9,1) #27
wire n10161_0;
wire n10162; //CHANX 1 (9,1) #34
wire n10162_0;
wire n10163; //CHANX 1 (9,1) #35
wire n10163_0;
wire n10164; //CHANX 1 (9,1) #42
wire n10164_0;
wire n10165; //CHANX 1 (9,1) #43
wire n10165_0;
wire n10166; //CHANX 1 (9,1) #50
wire n10166_0;
wire n10167; //CHANX 1 (9,1) #51
wire n10167_0;
wire n10168; //CHANX 1 (9,1) #58
wire n10168_0;
wire n10169; //CHANX 1 (9,1) #59
wire n10169_0;
wire n10170; //CHANX 1 (9,1) #66
wire n10170_0;
wire n10171; //CHANX 1 (9,1) #67
wire n10171_0;
wire n10172; //CHANX 1 (9,1) #74
wire n10172_0;
wire n10173; //CHANX 1 (9,1) #75
wire n10173_0;
wire n10174; //CHANX 1 (9,1) #82
wire n10174_0;
wire n10175; //CHANX 1 (9,1) #83
wire n10175_0;
wire n10176; //CHANX 2 (1,2) #0
wire n10176_0;
wire n10177; //CHANX 2 (1,2) #1
wire n10177_0;
wire n10178; //CHANX 3 (1,2) #2
wire n10178_0;
wire n10179; //CHANX 3 (1,2) #3
wire n10179_0;
wire n10180; //CHANX 4 (1,2) #4
wire n10180_0;
wire n10180_1;
buffer_wire buffer_10180_1 (.in(n10180_0), .out(n10180_1));
wire n10181; //CHANX 4 (1,2) #5
wire n10181_0;
wire n10181_1;
buffer_wire buffer_10181_1 (.in(n10181_0), .out(n10181_1));
wire n10182; //CHANX 1 (1,2) #6
wire n10182_0;
wire n10183; //CHANX 1 (1,2) #7
wire n10183_0;
wire n10184; //CHANX 2 (1,2) #8
wire n10184_0;
wire n10185; //CHANX 2 (1,2) #9
wire n10185_0;
wire n10186; //CHANX 3 (1,2) #10
wire n10186_0;
wire n10187; //CHANX 3 (1,2) #11
wire n10187_0;
wire n10188; //CHANX 4 (1,2) #12
wire n10188_0;
wire n10188_1;
buffer_wire buffer_10188_1 (.in(n10188_0), .out(n10188_1));
wire n10189; //CHANX 4 (1,2) #13
wire n10189_0;
wire n10189_1;
buffer_wire buffer_10189_1 (.in(n10189_0), .out(n10189_1));
wire n10190; //CHANX 1 (1,2) #14
wire n10190_0;
wire n10191; //CHANX 1 (1,2) #15
wire n10191_0;
wire n10192; //CHANX 2 (1,2) #16
wire n10192_0;
wire n10193; //CHANX 2 (1,2) #17
wire n10193_0;
wire n10194; //CHANX 3 (1,2) #18
wire n10194_0;
wire n10195; //CHANX 3 (1,2) #19
wire n10195_0;
wire n10196; //CHANX 4 (1,2) #20
wire n10196_0;
wire n10196_1;
buffer_wire buffer_10196_1 (.in(n10196_0), .out(n10196_1));
wire n10197; //CHANX 4 (1,2) #21
wire n10197_0;
wire n10197_1;
buffer_wire buffer_10197_1 (.in(n10197_0), .out(n10197_1));
wire n10198; //CHANX 1 (1,2) #22
wire n10198_0;
wire n10199; //CHANX 1 (1,2) #23
wire n10199_0;
wire n10200; //CHANX 2 (1,2) #24
wire n10200_0;
wire n10201; //CHANX 2 (1,2) #25
wire n10201_0;
wire n10202; //CHANX 3 (1,2) #26
wire n10202_0;
wire n10203; //CHANX 3 (1,2) #27
wire n10203_0;
wire n10204; //CHANX 4 (1,2) #28
wire n10204_0;
wire n10204_1;
buffer_wire buffer_10204_1 (.in(n10204_0), .out(n10204_1));
wire n10205; //CHANX 4 (1,2) #29
wire n10205_0;
wire n10205_1;
buffer_wire buffer_10205_1 (.in(n10205_0), .out(n10205_1));
wire n10206; //CHANX 1 (1,2) #30
wire n10206_0;
wire n10207; //CHANX 1 (1,2) #31
wire n10207_0;
wire n10208; //CHANX 2 (1,2) #32
wire n10208_0;
wire n10209; //CHANX 2 (1,2) #33
wire n10209_0;
wire n10210; //CHANX 3 (1,2) #34
wire n10210_0;
wire n10211; //CHANX 3 (1,2) #35
wire n10211_0;
wire n10212; //CHANX 4 (1,2) #36
wire n10212_0;
wire n10212_1;
buffer_wire buffer_10212_1 (.in(n10212_0), .out(n10212_1));
wire n10213; //CHANX 4 (1,2) #37
wire n10213_0;
wire n10213_1;
buffer_wire buffer_10213_1 (.in(n10213_0), .out(n10213_1));
wire n10214; //CHANX 1 (1,2) #38
wire n10214_0;
wire n10215; //CHANX 1 (1,2) #39
wire n10215_0;
wire n10216; //CHANX 2 (1,2) #40
wire n10216_0;
wire n10217; //CHANX 2 (1,2) #41
wire n10217_0;
wire n10218; //CHANX 3 (1,2) #42
wire n10218_0;
wire n10219; //CHANX 3 (1,2) #43
wire n10219_0;
wire n10220; //CHANX 4 (1,2) #44
wire n10220_0;
wire n10220_1;
buffer_wire buffer_10220_1 (.in(n10220_0), .out(n10220_1));
wire n10221; //CHANX 4 (1,2) #45
wire n10221_0;
wire n10221_1;
buffer_wire buffer_10221_1 (.in(n10221_0), .out(n10221_1));
wire n10222; //CHANX 1 (1,2) #46
wire n10222_0;
wire n10223; //CHANX 1 (1,2) #47
wire n10223_0;
wire n10224; //CHANX 2 (1,2) #48
wire n10224_0;
wire n10225; //CHANX 2 (1,2) #49
wire n10225_0;
wire n10226; //CHANX 3 (1,2) #50
wire n10226_0;
wire n10227; //CHANX 3 (1,2) #51
wire n10227_0;
wire n10228; //CHANX 4 (1,2) #52
wire n10228_0;
wire n10228_1;
buffer_wire buffer_10228_1 (.in(n10228_0), .out(n10228_1));
wire n10229; //CHANX 4 (1,2) #53
wire n10229_0;
wire n10229_1;
buffer_wire buffer_10229_1 (.in(n10229_0), .out(n10229_1));
wire n10230; //CHANX 1 (1,2) #54
wire n10230_0;
wire n10231; //CHANX 1 (1,2) #55
wire n10231_0;
wire n10232; //CHANX 2 (1,2) #56
wire n10232_0;
wire n10233; //CHANX 2 (1,2) #57
wire n10233_0;
wire n10234; //CHANX 3 (1,2) #58
wire n10234_0;
wire n10235; //CHANX 3 (1,2) #59
wire n10235_0;
wire n10236; //CHANX 4 (1,2) #60
wire n10236_0;
wire n10236_1;
buffer_wire buffer_10236_1 (.in(n10236_0), .out(n10236_1));
wire n10237; //CHANX 4 (1,2) #61
wire n10237_0;
wire n10237_1;
buffer_wire buffer_10237_1 (.in(n10237_0), .out(n10237_1));
wire n10238; //CHANX 1 (1,2) #62
wire n10238_0;
wire n10239; //CHANX 1 (1,2) #63
wire n10239_0;
wire n10240; //CHANX 2 (1,2) #64
wire n10240_0;
wire n10241; //CHANX 2 (1,2) #65
wire n10241_0;
wire n10242; //CHANX 3 (1,2) #66
wire n10242_0;
wire n10243; //CHANX 3 (1,2) #67
wire n10243_0;
wire n10244; //CHANX 4 (1,2) #68
wire n10244_0;
wire n10244_1;
buffer_wire buffer_10244_1 (.in(n10244_0), .out(n10244_1));
wire n10245; //CHANX 4 (1,2) #69
wire n10245_0;
wire n10245_1;
buffer_wire buffer_10245_1 (.in(n10245_0), .out(n10245_1));
wire n10246; //CHANX 1 (1,2) #70
wire n10246_0;
wire n10247; //CHANX 1 (1,2) #71
wire n10247_0;
wire n10248; //CHANX 2 (1,2) #72
wire n10248_0;
wire n10249; //CHANX 2 (1,2) #73
wire n10249_0;
wire n10250; //CHANX 3 (1,2) #74
wire n10250_0;
wire n10251; //CHANX 3 (1,2) #75
wire n10251_0;
wire n10252; //CHANX 4 (1,2) #76
wire n10252_0;
wire n10252_1;
buffer_wire buffer_10252_1 (.in(n10252_0), .out(n10252_1));
wire n10253; //CHANX 4 (1,2) #77
wire n10253_0;
wire n10253_1;
buffer_wire buffer_10253_1 (.in(n10253_0), .out(n10253_1));
wire n10254; //CHANX 1 (1,2) #78
wire n10254_0;
wire n10255; //CHANX 1 (1,2) #79
wire n10255_0;
wire n10256; //CHANX 6 (1,2) #80
wire n10256_0;
wire n10256_1;
buffer_wire buffer_10256_1 (.in(n10256_0), .out(n10256_1));
wire n10257; //CHANX 6 (1,2) #81
wire n10257_0;
wire n10257_1;
buffer_wire buffer_10257_1 (.in(n10257_0), .out(n10257_1));
wire n10258; //CHANX 7 (1,2) #82
wire n10258_0;
wire n10258_1;
wire n10258_2;
buffer_wire buffer_10258_2 (.in(n10258_1), .out(n10258_2));
buffer_wire buffer_10258_1 (.in(n10258_0), .out(n10258_1));
wire n10259; //CHANX 7 (1,2) #83
wire n10259_0;
wire n10259_1;
wire n10259_2;
buffer_wire buffer_10259_2 (.in(n10259_1), .out(n10259_2));
buffer_wire buffer_10259_1 (.in(n10259_0), .out(n10259_1));
wire n10260; //CHANX 8 (1,2) #84
wire n10260_0;
wire n10260_1;
wire n10260_2;
buffer_wire buffer_10260_2 (.in(n10260_1), .out(n10260_2));
buffer_wire buffer_10260_1 (.in(n10260_0), .out(n10260_1));
wire n10261; //CHANX 8 (1,2) #85
wire n10261_0;
wire n10261_1;
wire n10261_2;
buffer_wire buffer_10261_2 (.in(n10261_1), .out(n10261_2));
buffer_wire buffer_10261_1 (.in(n10261_0), .out(n10261_1));
wire n10262; //CHANX 9 (1,2) #86
wire n10262_0;
wire n10262_1;
wire n10262_2;
buffer_wire buffer_10262_2 (.in(n10262_1), .out(n10262_2));
buffer_wire buffer_10262_1 (.in(n10262_0), .out(n10262_1));
wire n10263; //CHANX 9 (1,2) #87
wire n10263_0;
wire n10263_1;
wire n10263_2;
buffer_wire buffer_10263_2 (.in(n10263_1), .out(n10263_2));
buffer_wire buffer_10263_1 (.in(n10263_0), .out(n10263_1));
wire n10264; //CHANX 9 (1,2) #88
wire n10264_0;
wire n10264_1;
wire n10264_2;
buffer_wire buffer_10264_2 (.in(n10264_1), .out(n10264_2));
buffer_wire buffer_10264_1 (.in(n10264_0), .out(n10264_1));
wire n10265; //CHANX 9 (1,2) #89
wire n10265_0;
wire n10265_1;
wire n10265_2;
buffer_wire buffer_10265_2 (.in(n10265_1), .out(n10265_2));
buffer_wire buffer_10265_1 (.in(n10265_0), .out(n10265_1));
wire n10266; //CHANX 9 (1,2) #90
wire n10266_0;
wire n10266_1;
wire n10266_2;
buffer_wire buffer_10266_2 (.in(n10266_1), .out(n10266_2));
buffer_wire buffer_10266_1 (.in(n10266_0), .out(n10266_1));
wire n10267; //CHANX 9 (1,2) #91
wire n10267_0;
wire n10267_1;
wire n10267_2;
buffer_wire buffer_10267_2 (.in(n10267_1), .out(n10267_2));
buffer_wire buffer_10267_1 (.in(n10267_0), .out(n10267_1));
wire n10268; //CHANX 4 (2,2) #6
wire n10268_0;
wire n10268_1;
buffer_wire buffer_10268_1 (.in(n10268_0), .out(n10268_1));
wire n10269; //CHANX 4 (2,2) #7
wire n10269_0;
wire n10269_1;
buffer_wire buffer_10269_1 (.in(n10269_0), .out(n10269_1));
wire n10270; //CHANX 4 (2,2) #14
wire n10270_0;
wire n10270_1;
buffer_wire buffer_10270_1 (.in(n10270_0), .out(n10270_1));
wire n10271; //CHANX 4 (2,2) #15
wire n10271_0;
wire n10271_1;
buffer_wire buffer_10271_1 (.in(n10271_0), .out(n10271_1));
wire n10272; //CHANX 4 (2,2) #22
wire n10272_0;
wire n10272_1;
buffer_wire buffer_10272_1 (.in(n10272_0), .out(n10272_1));
wire n10273; //CHANX 4 (2,2) #23
wire n10273_0;
wire n10273_1;
buffer_wire buffer_10273_1 (.in(n10273_0), .out(n10273_1));
wire n10274; //CHANX 4 (2,2) #30
wire n10274_0;
wire n10274_1;
buffer_wire buffer_10274_1 (.in(n10274_0), .out(n10274_1));
wire n10275; //CHANX 4 (2,2) #31
wire n10275_0;
wire n10275_1;
buffer_wire buffer_10275_1 (.in(n10275_0), .out(n10275_1));
wire n10276; //CHANX 4 (2,2) #38
wire n10276_0;
wire n10276_1;
buffer_wire buffer_10276_1 (.in(n10276_0), .out(n10276_1));
wire n10277; //CHANX 4 (2,2) #39
wire n10277_0;
wire n10277_1;
buffer_wire buffer_10277_1 (.in(n10277_0), .out(n10277_1));
wire n10278; //CHANX 4 (2,2) #46
wire n10278_0;
wire n10278_1;
buffer_wire buffer_10278_1 (.in(n10278_0), .out(n10278_1));
wire n10279; //CHANX 4 (2,2) #47
wire n10279_0;
wire n10279_1;
buffer_wire buffer_10279_1 (.in(n10279_0), .out(n10279_1));
wire n10280; //CHANX 4 (2,2) #54
wire n10280_0;
wire n10280_1;
buffer_wire buffer_10280_1 (.in(n10280_0), .out(n10280_1));
wire n10281; //CHANX 4 (2,2) #55
wire n10281_0;
wire n10281_1;
buffer_wire buffer_10281_1 (.in(n10281_0), .out(n10281_1));
wire n10282; //CHANX 4 (2,2) #62
wire n10282_0;
wire n10282_1;
buffer_wire buffer_10282_1 (.in(n10282_0), .out(n10282_1));
wire n10283; //CHANX 4 (2,2) #63
wire n10283_0;
wire n10283_1;
buffer_wire buffer_10283_1 (.in(n10283_0), .out(n10283_1));
wire n10284; //CHANX 4 (2,2) #70
wire n10284_0;
wire n10284_1;
buffer_wire buffer_10284_1 (.in(n10284_0), .out(n10284_1));
wire n10285; //CHANX 4 (2,2) #71
wire n10285_0;
wire n10285_1;
buffer_wire buffer_10285_1 (.in(n10285_0), .out(n10285_1));
wire n10286; //CHANX 4 (2,2) #78
wire n10286_0;
wire n10286_1;
buffer_wire buffer_10286_1 (.in(n10286_0), .out(n10286_1));
wire n10287; //CHANX 4 (2,2) #79
wire n10287_0;
wire n10287_1;
buffer_wire buffer_10287_1 (.in(n10287_0), .out(n10287_1));
wire n10288; //CHANX 4 (3,2) #0
wire n10288_0;
wire n10288_1;
buffer_wire buffer_10288_1 (.in(n10288_0), .out(n10288_1));
wire n10289; //CHANX 4 (3,2) #1
wire n10289_0;
wire n10289_1;
buffer_wire buffer_10289_1 (.in(n10289_0), .out(n10289_1));
wire n10290; //CHANX 4 (3,2) #8
wire n10290_0;
wire n10290_1;
buffer_wire buffer_10290_1 (.in(n10290_0), .out(n10290_1));
wire n10291; //CHANX 4 (3,2) #9
wire n10291_0;
wire n10291_1;
buffer_wire buffer_10291_1 (.in(n10291_0), .out(n10291_1));
wire n10292; //CHANX 4 (3,2) #16
wire n10292_0;
wire n10292_1;
buffer_wire buffer_10292_1 (.in(n10292_0), .out(n10292_1));
wire n10293; //CHANX 4 (3,2) #17
wire n10293_0;
wire n10293_1;
buffer_wire buffer_10293_1 (.in(n10293_0), .out(n10293_1));
wire n10294; //CHANX 4 (3,2) #24
wire n10294_0;
wire n10294_1;
buffer_wire buffer_10294_1 (.in(n10294_0), .out(n10294_1));
wire n10295; //CHANX 4 (3,2) #25
wire n10295_0;
wire n10295_1;
buffer_wire buffer_10295_1 (.in(n10295_0), .out(n10295_1));
wire n10296; //CHANX 4 (3,2) #32
wire n10296_0;
wire n10296_1;
buffer_wire buffer_10296_1 (.in(n10296_0), .out(n10296_1));
wire n10297; //CHANX 4 (3,2) #33
wire n10297_0;
wire n10297_1;
buffer_wire buffer_10297_1 (.in(n10297_0), .out(n10297_1));
wire n10298; //CHANX 4 (3,2) #40
wire n10298_0;
wire n10298_1;
buffer_wire buffer_10298_1 (.in(n10298_0), .out(n10298_1));
wire n10299; //CHANX 4 (3,2) #41
wire n10299_0;
wire n10299_1;
buffer_wire buffer_10299_1 (.in(n10299_0), .out(n10299_1));
wire n10300; //CHANX 4 (3,2) #48
wire n10300_0;
wire n10300_1;
buffer_wire buffer_10300_1 (.in(n10300_0), .out(n10300_1));
wire n10301; //CHANX 4 (3,2) #49
wire n10301_0;
wire n10301_1;
buffer_wire buffer_10301_1 (.in(n10301_0), .out(n10301_1));
wire n10302; //CHANX 4 (3,2) #56
wire n10302_0;
wire n10302_1;
buffer_wire buffer_10302_1 (.in(n10302_0), .out(n10302_1));
wire n10303; //CHANX 4 (3,2) #57
wire n10303_0;
wire n10303_1;
buffer_wire buffer_10303_1 (.in(n10303_0), .out(n10303_1));
wire n10304; //CHANX 4 (3,2) #64
wire n10304_0;
wire n10304_1;
buffer_wire buffer_10304_1 (.in(n10304_0), .out(n10304_1));
wire n10305; //CHANX 4 (3,2) #65
wire n10305_0;
wire n10305_1;
buffer_wire buffer_10305_1 (.in(n10305_0), .out(n10305_1));
wire n10306; //CHANX 4 (3,2) #72
wire n10306_0;
wire n10306_1;
buffer_wire buffer_10306_1 (.in(n10306_0), .out(n10306_1));
wire n10307; //CHANX 4 (3,2) #73
wire n10307_0;
wire n10307_1;
buffer_wire buffer_10307_1 (.in(n10307_0), .out(n10307_1));
wire n10308; //CHANX 4 (4,2) #2
wire n10308_0;
wire n10308_1;
buffer_wire buffer_10308_1 (.in(n10308_0), .out(n10308_1));
wire n10309; //CHANX 4 (4,2) #3
wire n10309_0;
wire n10309_1;
buffer_wire buffer_10309_1 (.in(n10309_0), .out(n10309_1));
wire n10310; //CHANX 4 (4,2) #10
wire n10310_0;
wire n10310_1;
buffer_wire buffer_10310_1 (.in(n10310_0), .out(n10310_1));
wire n10311; //CHANX 4 (4,2) #11
wire n10311_0;
wire n10311_1;
buffer_wire buffer_10311_1 (.in(n10311_0), .out(n10311_1));
wire n10312; //CHANX 4 (4,2) #18
wire n10312_0;
wire n10312_1;
buffer_wire buffer_10312_1 (.in(n10312_0), .out(n10312_1));
wire n10313; //CHANX 4 (4,2) #19
wire n10313_0;
wire n10313_1;
buffer_wire buffer_10313_1 (.in(n10313_0), .out(n10313_1));
wire n10314; //CHANX 4 (4,2) #26
wire n10314_0;
wire n10314_1;
buffer_wire buffer_10314_1 (.in(n10314_0), .out(n10314_1));
wire n10315; //CHANX 4 (4,2) #27
wire n10315_0;
wire n10315_1;
buffer_wire buffer_10315_1 (.in(n10315_0), .out(n10315_1));
wire n10316; //CHANX 4 (4,2) #34
wire n10316_0;
wire n10316_1;
buffer_wire buffer_10316_1 (.in(n10316_0), .out(n10316_1));
wire n10317; //CHANX 4 (4,2) #35
wire n10317_0;
wire n10317_1;
buffer_wire buffer_10317_1 (.in(n10317_0), .out(n10317_1));
wire n10318; //CHANX 4 (4,2) #42
wire n10318_0;
wire n10318_1;
buffer_wire buffer_10318_1 (.in(n10318_0), .out(n10318_1));
wire n10319; //CHANX 4 (4,2) #43
wire n10319_0;
wire n10319_1;
buffer_wire buffer_10319_1 (.in(n10319_0), .out(n10319_1));
wire n10320; //CHANX 4 (4,2) #50
wire n10320_0;
wire n10320_1;
buffer_wire buffer_10320_1 (.in(n10320_0), .out(n10320_1));
wire n10321; //CHANX 4 (4,2) #51
wire n10321_0;
wire n10321_1;
buffer_wire buffer_10321_1 (.in(n10321_0), .out(n10321_1));
wire n10322; //CHANX 4 (4,2) #58
wire n10322_0;
wire n10322_1;
buffer_wire buffer_10322_1 (.in(n10322_0), .out(n10322_1));
wire n10323; //CHANX 4 (4,2) #59
wire n10323_0;
wire n10323_1;
buffer_wire buffer_10323_1 (.in(n10323_0), .out(n10323_1));
wire n10324; //CHANX 4 (4,2) #66
wire n10324_0;
wire n10324_1;
buffer_wire buffer_10324_1 (.in(n10324_0), .out(n10324_1));
wire n10325; //CHANX 4 (4,2) #67
wire n10325_0;
wire n10325_1;
buffer_wire buffer_10325_1 (.in(n10325_0), .out(n10325_1));
wire n10326; //CHANX 4 (4,2) #74
wire n10326_0;
wire n10326_1;
buffer_wire buffer_10326_1 (.in(n10326_0), .out(n10326_1));
wire n10327; //CHANX 4 (4,2) #75
wire n10327_0;
wire n10327_1;
buffer_wire buffer_10327_1 (.in(n10327_0), .out(n10327_1));
wire n10328; //CHANX 4 (5,2) #4
wire n10328_0;
wire n10328_1;
buffer_wire buffer_10328_1 (.in(n10328_0), .out(n10328_1));
wire n10329; //CHANX 4 (5,2) #5
wire n10329_0;
wire n10329_1;
buffer_wire buffer_10329_1 (.in(n10329_0), .out(n10329_1));
wire n10330; //CHANX 4 (5,2) #12
wire n10330_0;
wire n10330_1;
buffer_wire buffer_10330_1 (.in(n10330_0), .out(n10330_1));
wire n10331; //CHANX 4 (5,2) #13
wire n10331_0;
wire n10331_1;
buffer_wire buffer_10331_1 (.in(n10331_0), .out(n10331_1));
wire n10332; //CHANX 4 (5,2) #20
wire n10332_0;
wire n10332_1;
buffer_wire buffer_10332_1 (.in(n10332_0), .out(n10332_1));
wire n10333; //CHANX 4 (5,2) #21
wire n10333_0;
wire n10333_1;
buffer_wire buffer_10333_1 (.in(n10333_0), .out(n10333_1));
wire n10334; //CHANX 4 (5,2) #28
wire n10334_0;
wire n10334_1;
buffer_wire buffer_10334_1 (.in(n10334_0), .out(n10334_1));
wire n10335; //CHANX 4 (5,2) #29
wire n10335_0;
wire n10335_1;
buffer_wire buffer_10335_1 (.in(n10335_0), .out(n10335_1));
wire n10336; //CHANX 4 (5,2) #36
wire n10336_0;
wire n10336_1;
buffer_wire buffer_10336_1 (.in(n10336_0), .out(n10336_1));
wire n10337; //CHANX 4 (5,2) #37
wire n10337_0;
wire n10337_1;
buffer_wire buffer_10337_1 (.in(n10337_0), .out(n10337_1));
wire n10338; //CHANX 4 (5,2) #44
wire n10338_0;
wire n10338_1;
buffer_wire buffer_10338_1 (.in(n10338_0), .out(n10338_1));
wire n10339; //CHANX 4 (5,2) #45
wire n10339_0;
wire n10339_1;
buffer_wire buffer_10339_1 (.in(n10339_0), .out(n10339_1));
wire n10340; //CHANX 4 (5,2) #52
wire n10340_0;
wire n10340_1;
buffer_wire buffer_10340_1 (.in(n10340_0), .out(n10340_1));
wire n10341; //CHANX 4 (5,2) #53
wire n10341_0;
wire n10341_1;
buffer_wire buffer_10341_1 (.in(n10341_0), .out(n10341_1));
wire n10342; //CHANX 4 (5,2) #60
wire n10342_0;
wire n10342_1;
buffer_wire buffer_10342_1 (.in(n10342_0), .out(n10342_1));
wire n10343; //CHANX 4 (5,2) #61
wire n10343_0;
wire n10343_1;
buffer_wire buffer_10343_1 (.in(n10343_0), .out(n10343_1));
wire n10344; //CHANX 4 (5,2) #68
wire n10344_0;
wire n10344_1;
buffer_wire buffer_10344_1 (.in(n10344_0), .out(n10344_1));
wire n10345; //CHANX 4 (5,2) #69
wire n10345_0;
wire n10345_1;
buffer_wire buffer_10345_1 (.in(n10345_0), .out(n10345_1));
wire n10346; //CHANX 4 (5,2) #76
wire n10346_0;
wire n10346_1;
buffer_wire buffer_10346_1 (.in(n10346_0), .out(n10346_1));
wire n10347; //CHANX 4 (5,2) #77
wire n10347_0;
wire n10347_1;
buffer_wire buffer_10347_1 (.in(n10347_0), .out(n10347_1));
wire n10348; //CHANX 4 (6,2) #6
wire n10348_0;
wire n10348_1;
buffer_wire buffer_10348_1 (.in(n10348_0), .out(n10348_1));
wire n10349; //CHANX 4 (6,2) #7
wire n10349_0;
wire n10349_1;
buffer_wire buffer_10349_1 (.in(n10349_0), .out(n10349_1));
wire n10350; //CHANX 4 (6,2) #14
wire n10350_0;
wire n10350_1;
buffer_wire buffer_10350_1 (.in(n10350_0), .out(n10350_1));
wire n10351; //CHANX 4 (6,2) #15
wire n10351_0;
wire n10351_1;
buffer_wire buffer_10351_1 (.in(n10351_0), .out(n10351_1));
wire n10352; //CHANX 4 (6,2) #22
wire n10352_0;
wire n10352_1;
buffer_wire buffer_10352_1 (.in(n10352_0), .out(n10352_1));
wire n10353; //CHANX 4 (6,2) #23
wire n10353_0;
wire n10353_1;
buffer_wire buffer_10353_1 (.in(n10353_0), .out(n10353_1));
wire n10354; //CHANX 4 (6,2) #30
wire n10354_0;
wire n10354_1;
buffer_wire buffer_10354_1 (.in(n10354_0), .out(n10354_1));
wire n10355; //CHANX 4 (6,2) #31
wire n10355_0;
wire n10355_1;
buffer_wire buffer_10355_1 (.in(n10355_0), .out(n10355_1));
wire n10356; //CHANX 4 (6,2) #38
wire n10356_0;
wire n10356_1;
buffer_wire buffer_10356_1 (.in(n10356_0), .out(n10356_1));
wire n10357; //CHANX 4 (6,2) #39
wire n10357_0;
wire n10357_1;
buffer_wire buffer_10357_1 (.in(n10357_0), .out(n10357_1));
wire n10358; //CHANX 4 (6,2) #46
wire n10358_0;
wire n10358_1;
buffer_wire buffer_10358_1 (.in(n10358_0), .out(n10358_1));
wire n10359; //CHANX 4 (6,2) #47
wire n10359_0;
wire n10359_1;
buffer_wire buffer_10359_1 (.in(n10359_0), .out(n10359_1));
wire n10360; //CHANX 4 (6,2) #54
wire n10360_0;
wire n10360_1;
buffer_wire buffer_10360_1 (.in(n10360_0), .out(n10360_1));
wire n10361; //CHANX 4 (6,2) #55
wire n10361_0;
wire n10361_1;
buffer_wire buffer_10361_1 (.in(n10361_0), .out(n10361_1));
wire n10362; //CHANX 4 (6,2) #62
wire n10362_0;
wire n10362_1;
buffer_wire buffer_10362_1 (.in(n10362_0), .out(n10362_1));
wire n10363; //CHANX 4 (6,2) #63
wire n10363_0;
wire n10363_1;
buffer_wire buffer_10363_1 (.in(n10363_0), .out(n10363_1));
wire n10364; //CHANX 4 (6,2) #70
wire n10364_0;
wire n10364_1;
buffer_wire buffer_10364_1 (.in(n10364_0), .out(n10364_1));
wire n10365; //CHANX 4 (6,2) #71
wire n10365_0;
wire n10365_1;
buffer_wire buffer_10365_1 (.in(n10365_0), .out(n10365_1));
wire n10366; //CHANX 4 (6,2) #78
wire n10366_0;
wire n10366_1;
buffer_wire buffer_10366_1 (.in(n10366_0), .out(n10366_1));
wire n10367; //CHANX 4 (6,2) #79
wire n10367_0;
wire n10367_1;
buffer_wire buffer_10367_1 (.in(n10367_0), .out(n10367_1));
wire n10368; //CHANX 3 (7,2) #0
wire n10368_0;
wire n10369; //CHANX 3 (7,2) #1
wire n10369_0;
wire n10370; //CHANX 3 (7,2) #8
wire n10370_0;
wire n10371; //CHANX 3 (7,2) #9
wire n10371_0;
wire n10372; //CHANX 3 (7,2) #16
wire n10372_0;
wire n10373; //CHANX 3 (7,2) #17
wire n10373_0;
wire n10374; //CHANX 3 (7,2) #24
wire n10374_0;
wire n10375; //CHANX 3 (7,2) #25
wire n10375_0;
wire n10376; //CHANX 3 (7,2) #32
wire n10376_0;
wire n10377; //CHANX 3 (7,2) #33
wire n10377_0;
wire n10378; //CHANX 3 (7,2) #40
wire n10378_0;
wire n10379; //CHANX 3 (7,2) #41
wire n10379_0;
wire n10380; //CHANX 3 (7,2) #48
wire n10380_0;
wire n10381; //CHANX 3 (7,2) #49
wire n10381_0;
wire n10382; //CHANX 3 (7,2) #56
wire n10382_0;
wire n10383; //CHANX 3 (7,2) #57
wire n10383_0;
wire n10384; //CHANX 3 (7,2) #64
wire n10384_0;
wire n10385; //CHANX 3 (7,2) #65
wire n10385_0;
wire n10386; //CHANX 3 (7,2) #72
wire n10386_0;
wire n10387; //CHANX 3 (7,2) #73
wire n10387_0;
wire n10388; //CHANX 3 (7,2) #80
wire n10388_0;
wire n10389; //CHANX 3 (7,2) #81
wire n10389_0;
wire n10390; //CHANX 2 (8,2) #2
wire n10390_0;
wire n10391; //CHANX 2 (8,2) #3
wire n10391_0;
wire n10392; //CHANX 2 (8,2) #10
wire n10392_0;
wire n10393; //CHANX 2 (8,2) #11
wire n10393_0;
wire n10394; //CHANX 2 (8,2) #18
wire n10394_0;
wire n10395; //CHANX 2 (8,2) #19
wire n10395_0;
wire n10396; //CHANX 2 (8,2) #26
wire n10396_0;
wire n10397; //CHANX 2 (8,2) #27
wire n10397_0;
wire n10398; //CHANX 2 (8,2) #34
wire n10398_0;
wire n10399; //CHANX 2 (8,2) #35
wire n10399_0;
wire n10400; //CHANX 2 (8,2) #42
wire n10400_0;
wire n10401; //CHANX 2 (8,2) #43
wire n10401_0;
wire n10402; //CHANX 2 (8,2) #50
wire n10402_0;
wire n10403; //CHANX 2 (8,2) #51
wire n10403_0;
wire n10404; //CHANX 2 (8,2) #58
wire n10404_0;
wire n10405; //CHANX 2 (8,2) #59
wire n10405_0;
wire n10406; //CHANX 2 (8,2) #66
wire n10406_0;
wire n10407; //CHANX 2 (8,2) #67
wire n10407_0;
wire n10408; //CHANX 2 (8,2) #74
wire n10408_0;
wire n10409; //CHANX 2 (8,2) #75
wire n10409_0;
wire n10410; //CHANX 2 (8,2) #82
wire n10410_0;
wire n10411; //CHANX 2 (8,2) #83
wire n10411_0;
wire n10412; //CHANX 1 (9,2) #4
wire n10412_0;
wire n10413; //CHANX 1 (9,2) #5
wire n10413_0;
wire n10414; //CHANX 1 (9,2) #12
wire n10414_0;
wire n10415; //CHANX 1 (9,2) #13
wire n10415_0;
wire n10416; //CHANX 1 (9,2) #20
wire n10416_0;
wire n10417; //CHANX 1 (9,2) #21
wire n10417_0;
wire n10418; //CHANX 1 (9,2) #28
wire n10418_0;
wire n10419; //CHANX 1 (9,2) #29
wire n10419_0;
wire n10420; //CHANX 1 (9,2) #36
wire n10420_0;
wire n10421; //CHANX 1 (9,2) #37
wire n10421_0;
wire n10422; //CHANX 1 (9,2) #44
wire n10422_0;
wire n10423; //CHANX 1 (9,2) #45
wire n10423_0;
wire n10424; //CHANX 1 (9,2) #52
wire n10424_0;
wire n10425; //CHANX 1 (9,2) #53
wire n10425_0;
wire n10426; //CHANX 1 (9,2) #60
wire n10426_0;
wire n10427; //CHANX 1 (9,2) #61
wire n10427_0;
wire n10428; //CHANX 1 (9,2) #68
wire n10428_0;
wire n10429; //CHANX 1 (9,2) #69
wire n10429_0;
wire n10430; //CHANX 1 (9,2) #76
wire n10430_0;
wire n10431; //CHANX 1 (9,2) #77
wire n10431_0;
wire n10432; //CHANX 1 (9,2) #84
wire n10432_0;
wire n10433; //CHANX 1 (9,2) #85
wire n10433_0;
wire n10434; //CHANX 1 (1,3) #0
wire n10434_0;
wire n10435; //CHANX 1 (1,3) #1
wire n10435_0;
wire n10436; //CHANX 2 (1,3) #2
wire n10436_0;
wire n10437; //CHANX 2 (1,3) #3
wire n10437_0;
wire n10438; //CHANX 3 (1,3) #4
wire n10438_0;
wire n10439; //CHANX 3 (1,3) #5
wire n10439_0;
wire n10440; //CHANX 4 (1,3) #6
wire n10440_0;
wire n10440_1;
buffer_wire buffer_10440_1 (.in(n10440_0), .out(n10440_1));
wire n10441; //CHANX 4 (1,3) #7
wire n10441_0;
wire n10441_1;
buffer_wire buffer_10441_1 (.in(n10441_0), .out(n10441_1));
wire n10442; //CHANX 1 (1,3) #8
wire n10442_0;
wire n10443; //CHANX 1 (1,3) #9
wire n10443_0;
wire n10444; //CHANX 2 (1,3) #10
wire n10444_0;
wire n10445; //CHANX 2 (1,3) #11
wire n10445_0;
wire n10446; //CHANX 3 (1,3) #12
wire n10446_0;
wire n10447; //CHANX 3 (1,3) #13
wire n10447_0;
wire n10448; //CHANX 4 (1,3) #14
wire n10448_0;
wire n10448_1;
buffer_wire buffer_10448_1 (.in(n10448_0), .out(n10448_1));
wire n10449; //CHANX 4 (1,3) #15
wire n10449_0;
wire n10449_1;
buffer_wire buffer_10449_1 (.in(n10449_0), .out(n10449_1));
wire n10450; //CHANX 1 (1,3) #16
wire n10450_0;
wire n10451; //CHANX 1 (1,3) #17
wire n10451_0;
wire n10452; //CHANX 2 (1,3) #18
wire n10452_0;
wire n10453; //CHANX 2 (1,3) #19
wire n10453_0;
wire n10454; //CHANX 3 (1,3) #20
wire n10454_0;
wire n10455; //CHANX 3 (1,3) #21
wire n10455_0;
wire n10456; //CHANX 4 (1,3) #22
wire n10456_0;
wire n10456_1;
buffer_wire buffer_10456_1 (.in(n10456_0), .out(n10456_1));
wire n10457; //CHANX 4 (1,3) #23
wire n10457_0;
wire n10457_1;
buffer_wire buffer_10457_1 (.in(n10457_0), .out(n10457_1));
wire n10458; //CHANX 1 (1,3) #24
wire n10458_0;
wire n10459; //CHANX 1 (1,3) #25
wire n10459_0;
wire n10460; //CHANX 2 (1,3) #26
wire n10460_0;
wire n10461; //CHANX 2 (1,3) #27
wire n10461_0;
wire n10462; //CHANX 3 (1,3) #28
wire n10462_0;
wire n10463; //CHANX 3 (1,3) #29
wire n10463_0;
wire n10464; //CHANX 4 (1,3) #30
wire n10464_0;
wire n10464_1;
buffer_wire buffer_10464_1 (.in(n10464_0), .out(n10464_1));
wire n10465; //CHANX 4 (1,3) #31
wire n10465_0;
wire n10465_1;
buffer_wire buffer_10465_1 (.in(n10465_0), .out(n10465_1));
wire n10466; //CHANX 1 (1,3) #32
wire n10466_0;
wire n10467; //CHANX 1 (1,3) #33
wire n10467_0;
wire n10468; //CHANX 2 (1,3) #34
wire n10468_0;
wire n10469; //CHANX 2 (1,3) #35
wire n10469_0;
wire n10470; //CHANX 3 (1,3) #36
wire n10470_0;
wire n10471; //CHANX 3 (1,3) #37
wire n10471_0;
wire n10472; //CHANX 4 (1,3) #38
wire n10472_0;
wire n10472_1;
buffer_wire buffer_10472_1 (.in(n10472_0), .out(n10472_1));
wire n10473; //CHANX 4 (1,3) #39
wire n10473_0;
wire n10473_1;
buffer_wire buffer_10473_1 (.in(n10473_0), .out(n10473_1));
wire n10474; //CHANX 1 (1,3) #40
wire n10474_0;
wire n10475; //CHANX 1 (1,3) #41
wire n10475_0;
wire n10476; //CHANX 2 (1,3) #42
wire n10476_0;
wire n10477; //CHANX 2 (1,3) #43
wire n10477_0;
wire n10478; //CHANX 3 (1,3) #44
wire n10478_0;
wire n10479; //CHANX 3 (1,3) #45
wire n10479_0;
wire n10480; //CHANX 4 (1,3) #46
wire n10480_0;
wire n10480_1;
buffer_wire buffer_10480_1 (.in(n10480_0), .out(n10480_1));
wire n10481; //CHANX 4 (1,3) #47
wire n10481_0;
wire n10481_1;
buffer_wire buffer_10481_1 (.in(n10481_0), .out(n10481_1));
wire n10482; //CHANX 1 (1,3) #48
wire n10482_0;
wire n10483; //CHANX 1 (1,3) #49
wire n10483_0;
wire n10484; //CHANX 2 (1,3) #50
wire n10484_0;
wire n10485; //CHANX 2 (1,3) #51
wire n10485_0;
wire n10486; //CHANX 3 (1,3) #52
wire n10486_0;
wire n10487; //CHANX 3 (1,3) #53
wire n10487_0;
wire n10488; //CHANX 4 (1,3) #54
wire n10488_0;
wire n10488_1;
buffer_wire buffer_10488_1 (.in(n10488_0), .out(n10488_1));
wire n10489; //CHANX 4 (1,3) #55
wire n10489_0;
wire n10489_1;
buffer_wire buffer_10489_1 (.in(n10489_0), .out(n10489_1));
wire n10490; //CHANX 1 (1,3) #56
wire n10490_0;
wire n10491; //CHANX 1 (1,3) #57
wire n10491_0;
wire n10492; //CHANX 2 (1,3) #58
wire n10492_0;
wire n10493; //CHANX 2 (1,3) #59
wire n10493_0;
wire n10494; //CHANX 3 (1,3) #60
wire n10494_0;
wire n10495; //CHANX 3 (1,3) #61
wire n10495_0;
wire n10496; //CHANX 4 (1,3) #62
wire n10496_0;
wire n10496_1;
buffer_wire buffer_10496_1 (.in(n10496_0), .out(n10496_1));
wire n10497; //CHANX 4 (1,3) #63
wire n10497_0;
wire n10497_1;
buffer_wire buffer_10497_1 (.in(n10497_0), .out(n10497_1));
wire n10498; //CHANX 1 (1,3) #64
wire n10498_0;
wire n10499; //CHANX 1 (1,3) #65
wire n10499_0;
wire n10500; //CHANX 2 (1,3) #66
wire n10500_0;
wire n10501; //CHANX 2 (1,3) #67
wire n10501_0;
wire n10502; //CHANX 3 (1,3) #68
wire n10502_0;
wire n10503; //CHANX 3 (1,3) #69
wire n10503_0;
wire n10504; //CHANX 4 (1,3) #70
wire n10504_0;
wire n10504_1;
buffer_wire buffer_10504_1 (.in(n10504_0), .out(n10504_1));
wire n10505; //CHANX 4 (1,3) #71
wire n10505_0;
wire n10505_1;
buffer_wire buffer_10505_1 (.in(n10505_0), .out(n10505_1));
wire n10506; //CHANX 1 (1,3) #72
wire n10506_0;
wire n10507; //CHANX 1 (1,3) #73
wire n10507_0;
wire n10508; //CHANX 2 (1,3) #74
wire n10508_0;
wire n10509; //CHANX 2 (1,3) #75
wire n10509_0;
wire n10510; //CHANX 3 (1,3) #76
wire n10510_0;
wire n10511; //CHANX 3 (1,3) #77
wire n10511_0;
wire n10512; //CHANX 4 (1,3) #78
wire n10512_0;
wire n10512_1;
buffer_wire buffer_10512_1 (.in(n10512_0), .out(n10512_1));
wire n10513; //CHANX 4 (1,3) #79
wire n10513_0;
wire n10513_1;
buffer_wire buffer_10513_1 (.in(n10513_0), .out(n10513_1));
wire n10514; //CHANX 5 (1,3) #80
wire n10514_0;
wire n10514_1;
buffer_wire buffer_10514_1 (.in(n10514_0), .out(n10514_1));
wire n10515; //CHANX 5 (1,3) #81
wire n10515_0;
wire n10515_1;
buffer_wire buffer_10515_1 (.in(n10515_0), .out(n10515_1));
wire n10516; //CHANX 6 (1,3) #82
wire n10516_0;
wire n10516_1;
buffer_wire buffer_10516_1 (.in(n10516_0), .out(n10516_1));
wire n10517; //CHANX 6 (1,3) #83
wire n10517_0;
wire n10517_1;
buffer_wire buffer_10517_1 (.in(n10517_0), .out(n10517_1));
wire n10518; //CHANX 7 (1,3) #84
wire n10518_0;
wire n10518_1;
wire n10518_2;
buffer_wire buffer_10518_2 (.in(n10518_1), .out(n10518_2));
buffer_wire buffer_10518_1 (.in(n10518_0), .out(n10518_1));
wire n10519; //CHANX 7 (1,3) #85
wire n10519_0;
wire n10519_1;
wire n10519_2;
buffer_wire buffer_10519_2 (.in(n10519_1), .out(n10519_2));
buffer_wire buffer_10519_1 (.in(n10519_0), .out(n10519_1));
wire n10520; //CHANX 8 (1,3) #86
wire n10520_0;
wire n10520_1;
wire n10520_2;
buffer_wire buffer_10520_2 (.in(n10520_1), .out(n10520_2));
buffer_wire buffer_10520_1 (.in(n10520_0), .out(n10520_1));
wire n10521; //CHANX 8 (1,3) #87
wire n10521_0;
wire n10521_1;
wire n10521_2;
buffer_wire buffer_10521_2 (.in(n10521_1), .out(n10521_2));
buffer_wire buffer_10521_1 (.in(n10521_0), .out(n10521_1));
wire n10522; //CHANX 9 (1,3) #88
wire n10522_0;
wire n10522_1;
wire n10522_2;
buffer_wire buffer_10522_2 (.in(n10522_1), .out(n10522_2));
buffer_wire buffer_10522_1 (.in(n10522_0), .out(n10522_1));
wire n10523; //CHANX 9 (1,3) #89
wire n10523_0;
wire n10523_1;
wire n10523_2;
buffer_wire buffer_10523_2 (.in(n10523_1), .out(n10523_2));
buffer_wire buffer_10523_1 (.in(n10523_0), .out(n10523_1));
wire n10524; //CHANX 9 (1,3) #90
wire n10524_0;
wire n10524_1;
wire n10524_2;
buffer_wire buffer_10524_2 (.in(n10524_1), .out(n10524_2));
buffer_wire buffer_10524_1 (.in(n10524_0), .out(n10524_1));
wire n10525; //CHANX 9 (1,3) #91
wire n10525_0;
wire n10525_1;
wire n10525_2;
buffer_wire buffer_10525_2 (.in(n10525_1), .out(n10525_2));
buffer_wire buffer_10525_1 (.in(n10525_0), .out(n10525_1));
wire n10526; //CHANX 4 (2,3) #0
wire n10526_0;
wire n10526_1;
buffer_wire buffer_10526_1 (.in(n10526_0), .out(n10526_1));
wire n10527; //CHANX 4 (2,3) #1
wire n10527_0;
wire n10527_1;
buffer_wire buffer_10527_1 (.in(n10527_0), .out(n10527_1));
wire n10528; //CHANX 4 (2,3) #8
wire n10528_0;
wire n10528_1;
buffer_wire buffer_10528_1 (.in(n10528_0), .out(n10528_1));
wire n10529; //CHANX 4 (2,3) #9
wire n10529_0;
wire n10529_1;
buffer_wire buffer_10529_1 (.in(n10529_0), .out(n10529_1));
wire n10530; //CHANX 4 (2,3) #16
wire n10530_0;
wire n10530_1;
buffer_wire buffer_10530_1 (.in(n10530_0), .out(n10530_1));
wire n10531; //CHANX 4 (2,3) #17
wire n10531_0;
wire n10531_1;
buffer_wire buffer_10531_1 (.in(n10531_0), .out(n10531_1));
wire n10532; //CHANX 4 (2,3) #24
wire n10532_0;
wire n10532_1;
buffer_wire buffer_10532_1 (.in(n10532_0), .out(n10532_1));
wire n10533; //CHANX 4 (2,3) #25
wire n10533_0;
wire n10533_1;
buffer_wire buffer_10533_1 (.in(n10533_0), .out(n10533_1));
wire n10534; //CHANX 4 (2,3) #32
wire n10534_0;
wire n10534_1;
buffer_wire buffer_10534_1 (.in(n10534_0), .out(n10534_1));
wire n10535; //CHANX 4 (2,3) #33
wire n10535_0;
wire n10535_1;
buffer_wire buffer_10535_1 (.in(n10535_0), .out(n10535_1));
wire n10536; //CHANX 4 (2,3) #40
wire n10536_0;
wire n10536_1;
buffer_wire buffer_10536_1 (.in(n10536_0), .out(n10536_1));
wire n10537; //CHANX 4 (2,3) #41
wire n10537_0;
wire n10537_1;
buffer_wire buffer_10537_1 (.in(n10537_0), .out(n10537_1));
wire n10538; //CHANX 4 (2,3) #48
wire n10538_0;
wire n10538_1;
buffer_wire buffer_10538_1 (.in(n10538_0), .out(n10538_1));
wire n10539; //CHANX 4 (2,3) #49
wire n10539_0;
wire n10539_1;
buffer_wire buffer_10539_1 (.in(n10539_0), .out(n10539_1));
wire n10540; //CHANX 4 (2,3) #56
wire n10540_0;
wire n10540_1;
buffer_wire buffer_10540_1 (.in(n10540_0), .out(n10540_1));
wire n10541; //CHANX 4 (2,3) #57
wire n10541_0;
wire n10541_1;
buffer_wire buffer_10541_1 (.in(n10541_0), .out(n10541_1));
wire n10542; //CHANX 4 (2,3) #64
wire n10542_0;
wire n10542_1;
buffer_wire buffer_10542_1 (.in(n10542_0), .out(n10542_1));
wire n10543; //CHANX 4 (2,3) #65
wire n10543_0;
wire n10543_1;
buffer_wire buffer_10543_1 (.in(n10543_0), .out(n10543_1));
wire n10544; //CHANX 4 (2,3) #72
wire n10544_0;
wire n10544_1;
buffer_wire buffer_10544_1 (.in(n10544_0), .out(n10544_1));
wire n10545; //CHANX 4 (2,3) #73
wire n10545_0;
wire n10545_1;
buffer_wire buffer_10545_1 (.in(n10545_0), .out(n10545_1));
wire n10546; //CHANX 4 (3,3) #2
wire n10546_0;
wire n10546_1;
buffer_wire buffer_10546_1 (.in(n10546_0), .out(n10546_1));
wire n10547; //CHANX 4 (3,3) #3
wire n10547_0;
wire n10547_1;
buffer_wire buffer_10547_1 (.in(n10547_0), .out(n10547_1));
wire n10548; //CHANX 4 (3,3) #10
wire n10548_0;
wire n10548_1;
buffer_wire buffer_10548_1 (.in(n10548_0), .out(n10548_1));
wire n10549; //CHANX 4 (3,3) #11
wire n10549_0;
wire n10549_1;
buffer_wire buffer_10549_1 (.in(n10549_0), .out(n10549_1));
wire n10550; //CHANX 4 (3,3) #18
wire n10550_0;
wire n10550_1;
buffer_wire buffer_10550_1 (.in(n10550_0), .out(n10550_1));
wire n10551; //CHANX 4 (3,3) #19
wire n10551_0;
wire n10551_1;
buffer_wire buffer_10551_1 (.in(n10551_0), .out(n10551_1));
wire n10552; //CHANX 4 (3,3) #26
wire n10552_0;
wire n10552_1;
buffer_wire buffer_10552_1 (.in(n10552_0), .out(n10552_1));
wire n10553; //CHANX 4 (3,3) #27
wire n10553_0;
wire n10553_1;
buffer_wire buffer_10553_1 (.in(n10553_0), .out(n10553_1));
wire n10554; //CHANX 4 (3,3) #34
wire n10554_0;
wire n10554_1;
buffer_wire buffer_10554_1 (.in(n10554_0), .out(n10554_1));
wire n10555; //CHANX 4 (3,3) #35
wire n10555_0;
wire n10555_1;
buffer_wire buffer_10555_1 (.in(n10555_0), .out(n10555_1));
wire n10556; //CHANX 4 (3,3) #42
wire n10556_0;
wire n10556_1;
buffer_wire buffer_10556_1 (.in(n10556_0), .out(n10556_1));
wire n10557; //CHANX 4 (3,3) #43
wire n10557_0;
wire n10557_1;
buffer_wire buffer_10557_1 (.in(n10557_0), .out(n10557_1));
wire n10558; //CHANX 4 (3,3) #50
wire n10558_0;
wire n10558_1;
buffer_wire buffer_10558_1 (.in(n10558_0), .out(n10558_1));
wire n10559; //CHANX 4 (3,3) #51
wire n10559_0;
wire n10559_1;
buffer_wire buffer_10559_1 (.in(n10559_0), .out(n10559_1));
wire n10560; //CHANX 4 (3,3) #58
wire n10560_0;
wire n10560_1;
buffer_wire buffer_10560_1 (.in(n10560_0), .out(n10560_1));
wire n10561; //CHANX 4 (3,3) #59
wire n10561_0;
wire n10561_1;
buffer_wire buffer_10561_1 (.in(n10561_0), .out(n10561_1));
wire n10562; //CHANX 4 (3,3) #66
wire n10562_0;
wire n10562_1;
buffer_wire buffer_10562_1 (.in(n10562_0), .out(n10562_1));
wire n10563; //CHANX 4 (3,3) #67
wire n10563_0;
wire n10563_1;
buffer_wire buffer_10563_1 (.in(n10563_0), .out(n10563_1));
wire n10564; //CHANX 4 (3,3) #74
wire n10564_0;
wire n10564_1;
buffer_wire buffer_10564_1 (.in(n10564_0), .out(n10564_1));
wire n10565; //CHANX 4 (3,3) #75
wire n10565_0;
wire n10565_1;
buffer_wire buffer_10565_1 (.in(n10565_0), .out(n10565_1));
wire n10566; //CHANX 4 (4,3) #4
wire n10566_0;
wire n10566_1;
buffer_wire buffer_10566_1 (.in(n10566_0), .out(n10566_1));
wire n10567; //CHANX 4 (4,3) #5
wire n10567_0;
wire n10567_1;
buffer_wire buffer_10567_1 (.in(n10567_0), .out(n10567_1));
wire n10568; //CHANX 4 (4,3) #12
wire n10568_0;
wire n10568_1;
buffer_wire buffer_10568_1 (.in(n10568_0), .out(n10568_1));
wire n10569; //CHANX 4 (4,3) #13
wire n10569_0;
wire n10569_1;
buffer_wire buffer_10569_1 (.in(n10569_0), .out(n10569_1));
wire n10570; //CHANX 4 (4,3) #20
wire n10570_0;
wire n10570_1;
buffer_wire buffer_10570_1 (.in(n10570_0), .out(n10570_1));
wire n10571; //CHANX 4 (4,3) #21
wire n10571_0;
wire n10571_1;
buffer_wire buffer_10571_1 (.in(n10571_0), .out(n10571_1));
wire n10572; //CHANX 4 (4,3) #28
wire n10572_0;
wire n10572_1;
buffer_wire buffer_10572_1 (.in(n10572_0), .out(n10572_1));
wire n10573; //CHANX 4 (4,3) #29
wire n10573_0;
wire n10573_1;
buffer_wire buffer_10573_1 (.in(n10573_0), .out(n10573_1));
wire n10574; //CHANX 4 (4,3) #36
wire n10574_0;
wire n10574_1;
buffer_wire buffer_10574_1 (.in(n10574_0), .out(n10574_1));
wire n10575; //CHANX 4 (4,3) #37
wire n10575_0;
wire n10575_1;
buffer_wire buffer_10575_1 (.in(n10575_0), .out(n10575_1));
wire n10576; //CHANX 4 (4,3) #44
wire n10576_0;
wire n10576_1;
buffer_wire buffer_10576_1 (.in(n10576_0), .out(n10576_1));
wire n10577; //CHANX 4 (4,3) #45
wire n10577_0;
wire n10577_1;
buffer_wire buffer_10577_1 (.in(n10577_0), .out(n10577_1));
wire n10578; //CHANX 4 (4,3) #52
wire n10578_0;
wire n10578_1;
buffer_wire buffer_10578_1 (.in(n10578_0), .out(n10578_1));
wire n10579; //CHANX 4 (4,3) #53
wire n10579_0;
wire n10579_1;
buffer_wire buffer_10579_1 (.in(n10579_0), .out(n10579_1));
wire n10580; //CHANX 4 (4,3) #60
wire n10580_0;
wire n10580_1;
buffer_wire buffer_10580_1 (.in(n10580_0), .out(n10580_1));
wire n10581; //CHANX 4 (4,3) #61
wire n10581_0;
wire n10581_1;
buffer_wire buffer_10581_1 (.in(n10581_0), .out(n10581_1));
wire n10582; //CHANX 4 (4,3) #68
wire n10582_0;
wire n10582_1;
buffer_wire buffer_10582_1 (.in(n10582_0), .out(n10582_1));
wire n10583; //CHANX 4 (4,3) #69
wire n10583_0;
wire n10583_1;
buffer_wire buffer_10583_1 (.in(n10583_0), .out(n10583_1));
wire n10584; //CHANX 4 (4,3) #76
wire n10584_0;
wire n10584_1;
buffer_wire buffer_10584_1 (.in(n10584_0), .out(n10584_1));
wire n10585; //CHANX 4 (4,3) #77
wire n10585_0;
wire n10585_1;
buffer_wire buffer_10585_1 (.in(n10585_0), .out(n10585_1));
wire n10586; //CHANX 4 (5,3) #6
wire n10586_0;
wire n10586_1;
buffer_wire buffer_10586_1 (.in(n10586_0), .out(n10586_1));
wire n10587; //CHANX 4 (5,3) #7
wire n10587_0;
wire n10587_1;
buffer_wire buffer_10587_1 (.in(n10587_0), .out(n10587_1));
wire n10588; //CHANX 4 (5,3) #14
wire n10588_0;
wire n10588_1;
buffer_wire buffer_10588_1 (.in(n10588_0), .out(n10588_1));
wire n10589; //CHANX 4 (5,3) #15
wire n10589_0;
wire n10589_1;
buffer_wire buffer_10589_1 (.in(n10589_0), .out(n10589_1));
wire n10590; //CHANX 4 (5,3) #22
wire n10590_0;
wire n10590_1;
buffer_wire buffer_10590_1 (.in(n10590_0), .out(n10590_1));
wire n10591; //CHANX 4 (5,3) #23
wire n10591_0;
wire n10591_1;
buffer_wire buffer_10591_1 (.in(n10591_0), .out(n10591_1));
wire n10592; //CHANX 4 (5,3) #30
wire n10592_0;
wire n10592_1;
buffer_wire buffer_10592_1 (.in(n10592_0), .out(n10592_1));
wire n10593; //CHANX 4 (5,3) #31
wire n10593_0;
wire n10593_1;
buffer_wire buffer_10593_1 (.in(n10593_0), .out(n10593_1));
wire n10594; //CHANX 4 (5,3) #38
wire n10594_0;
wire n10594_1;
buffer_wire buffer_10594_1 (.in(n10594_0), .out(n10594_1));
wire n10595; //CHANX 4 (5,3) #39
wire n10595_0;
wire n10595_1;
buffer_wire buffer_10595_1 (.in(n10595_0), .out(n10595_1));
wire n10596; //CHANX 4 (5,3) #46
wire n10596_0;
wire n10596_1;
buffer_wire buffer_10596_1 (.in(n10596_0), .out(n10596_1));
wire n10597; //CHANX 4 (5,3) #47
wire n10597_0;
wire n10597_1;
buffer_wire buffer_10597_1 (.in(n10597_0), .out(n10597_1));
wire n10598; //CHANX 4 (5,3) #54
wire n10598_0;
wire n10598_1;
buffer_wire buffer_10598_1 (.in(n10598_0), .out(n10598_1));
wire n10599; //CHANX 4 (5,3) #55
wire n10599_0;
wire n10599_1;
buffer_wire buffer_10599_1 (.in(n10599_0), .out(n10599_1));
wire n10600; //CHANX 4 (5,3) #62
wire n10600_0;
wire n10600_1;
buffer_wire buffer_10600_1 (.in(n10600_0), .out(n10600_1));
wire n10601; //CHANX 4 (5,3) #63
wire n10601_0;
wire n10601_1;
buffer_wire buffer_10601_1 (.in(n10601_0), .out(n10601_1));
wire n10602; //CHANX 4 (5,3) #70
wire n10602_0;
wire n10602_1;
buffer_wire buffer_10602_1 (.in(n10602_0), .out(n10602_1));
wire n10603; //CHANX 4 (5,3) #71
wire n10603_0;
wire n10603_1;
buffer_wire buffer_10603_1 (.in(n10603_0), .out(n10603_1));
wire n10604; //CHANX 4 (5,3) #78
wire n10604_0;
wire n10604_1;
buffer_wire buffer_10604_1 (.in(n10604_0), .out(n10604_1));
wire n10605; //CHANX 4 (5,3) #79
wire n10605_0;
wire n10605_1;
buffer_wire buffer_10605_1 (.in(n10605_0), .out(n10605_1));
wire n10606; //CHANX 4 (6,3) #0
wire n10606_0;
wire n10606_1;
buffer_wire buffer_10606_1 (.in(n10606_0), .out(n10606_1));
wire n10607; //CHANX 4 (6,3) #1
wire n10607_0;
wire n10607_1;
buffer_wire buffer_10607_1 (.in(n10607_0), .out(n10607_1));
wire n10608; //CHANX 4 (6,3) #8
wire n10608_0;
wire n10608_1;
buffer_wire buffer_10608_1 (.in(n10608_0), .out(n10608_1));
wire n10609; //CHANX 4 (6,3) #9
wire n10609_0;
wire n10609_1;
buffer_wire buffer_10609_1 (.in(n10609_0), .out(n10609_1));
wire n10610; //CHANX 4 (6,3) #16
wire n10610_0;
wire n10610_1;
buffer_wire buffer_10610_1 (.in(n10610_0), .out(n10610_1));
wire n10611; //CHANX 4 (6,3) #17
wire n10611_0;
wire n10611_1;
buffer_wire buffer_10611_1 (.in(n10611_0), .out(n10611_1));
wire n10612; //CHANX 4 (6,3) #24
wire n10612_0;
wire n10612_1;
buffer_wire buffer_10612_1 (.in(n10612_0), .out(n10612_1));
wire n10613; //CHANX 4 (6,3) #25
wire n10613_0;
wire n10613_1;
buffer_wire buffer_10613_1 (.in(n10613_0), .out(n10613_1));
wire n10614; //CHANX 4 (6,3) #32
wire n10614_0;
wire n10614_1;
buffer_wire buffer_10614_1 (.in(n10614_0), .out(n10614_1));
wire n10615; //CHANX 4 (6,3) #33
wire n10615_0;
wire n10615_1;
buffer_wire buffer_10615_1 (.in(n10615_0), .out(n10615_1));
wire n10616; //CHANX 4 (6,3) #40
wire n10616_0;
wire n10616_1;
buffer_wire buffer_10616_1 (.in(n10616_0), .out(n10616_1));
wire n10617; //CHANX 4 (6,3) #41
wire n10617_0;
wire n10617_1;
buffer_wire buffer_10617_1 (.in(n10617_0), .out(n10617_1));
wire n10618; //CHANX 4 (6,3) #48
wire n10618_0;
wire n10618_1;
buffer_wire buffer_10618_1 (.in(n10618_0), .out(n10618_1));
wire n10619; //CHANX 4 (6,3) #49
wire n10619_0;
wire n10619_1;
buffer_wire buffer_10619_1 (.in(n10619_0), .out(n10619_1));
wire n10620; //CHANX 4 (6,3) #56
wire n10620_0;
wire n10620_1;
buffer_wire buffer_10620_1 (.in(n10620_0), .out(n10620_1));
wire n10621; //CHANX 4 (6,3) #57
wire n10621_0;
wire n10621_1;
buffer_wire buffer_10621_1 (.in(n10621_0), .out(n10621_1));
wire n10622; //CHANX 4 (6,3) #64
wire n10622_0;
wire n10622_1;
buffer_wire buffer_10622_1 (.in(n10622_0), .out(n10622_1));
wire n10623; //CHANX 4 (6,3) #65
wire n10623_0;
wire n10623_1;
buffer_wire buffer_10623_1 (.in(n10623_0), .out(n10623_1));
wire n10624; //CHANX 4 (6,3) #72
wire n10624_0;
wire n10624_1;
buffer_wire buffer_10624_1 (.in(n10624_0), .out(n10624_1));
wire n10625; //CHANX 4 (6,3) #73
wire n10625_0;
wire n10625_1;
buffer_wire buffer_10625_1 (.in(n10625_0), .out(n10625_1));
wire n10626; //CHANX 4 (6,3) #80
wire n10626_0;
wire n10626_1;
buffer_wire buffer_10626_1 (.in(n10626_0), .out(n10626_1));
wire n10627; //CHANX 4 (6,3) #81
wire n10627_0;
wire n10627_1;
buffer_wire buffer_10627_1 (.in(n10627_0), .out(n10627_1));
wire n10628; //CHANX 3 (7,3) #2
wire n10628_0;
wire n10629; //CHANX 3 (7,3) #3
wire n10629_0;
wire n10630; //CHANX 3 (7,3) #10
wire n10630_0;
wire n10631; //CHANX 3 (7,3) #11
wire n10631_0;
wire n10632; //CHANX 3 (7,3) #18
wire n10632_0;
wire n10633; //CHANX 3 (7,3) #19
wire n10633_0;
wire n10634; //CHANX 3 (7,3) #26
wire n10634_0;
wire n10635; //CHANX 3 (7,3) #27
wire n10635_0;
wire n10636; //CHANX 3 (7,3) #34
wire n10636_0;
wire n10637; //CHANX 3 (7,3) #35
wire n10637_0;
wire n10638; //CHANX 3 (7,3) #42
wire n10638_0;
wire n10639; //CHANX 3 (7,3) #43
wire n10639_0;
wire n10640; //CHANX 3 (7,3) #50
wire n10640_0;
wire n10641; //CHANX 3 (7,3) #51
wire n10641_0;
wire n10642; //CHANX 3 (7,3) #58
wire n10642_0;
wire n10643; //CHANX 3 (7,3) #59
wire n10643_0;
wire n10644; //CHANX 3 (7,3) #66
wire n10644_0;
wire n10645; //CHANX 3 (7,3) #67
wire n10645_0;
wire n10646; //CHANX 3 (7,3) #74
wire n10646_0;
wire n10647; //CHANX 3 (7,3) #75
wire n10647_0;
wire n10648; //CHANX 3 (7,3) #82
wire n10648_0;
wire n10649; //CHANX 3 (7,3) #83
wire n10649_0;
wire n10650; //CHANX 2 (8,3) #4
wire n10650_0;
wire n10651; //CHANX 2 (8,3) #5
wire n10651_0;
wire n10652; //CHANX 2 (8,3) #12
wire n10652_0;
wire n10653; //CHANX 2 (8,3) #13
wire n10653_0;
wire n10654; //CHANX 2 (8,3) #20
wire n10654_0;
wire n10655; //CHANX 2 (8,3) #21
wire n10655_0;
wire n10656; //CHANX 2 (8,3) #28
wire n10656_0;
wire n10657; //CHANX 2 (8,3) #29
wire n10657_0;
wire n10658; //CHANX 2 (8,3) #36
wire n10658_0;
wire n10659; //CHANX 2 (8,3) #37
wire n10659_0;
wire n10660; //CHANX 2 (8,3) #44
wire n10660_0;
wire n10661; //CHANX 2 (8,3) #45
wire n10661_0;
wire n10662; //CHANX 2 (8,3) #52
wire n10662_0;
wire n10663; //CHANX 2 (8,3) #53
wire n10663_0;
wire n10664; //CHANX 2 (8,3) #60
wire n10664_0;
wire n10665; //CHANX 2 (8,3) #61
wire n10665_0;
wire n10666; //CHANX 2 (8,3) #68
wire n10666_0;
wire n10667; //CHANX 2 (8,3) #69
wire n10667_0;
wire n10668; //CHANX 2 (8,3) #76
wire n10668_0;
wire n10669; //CHANX 2 (8,3) #77
wire n10669_0;
wire n10670; //CHANX 2 (8,3) #84
wire n10670_0;
wire n10671; //CHANX 2 (8,3) #85
wire n10671_0;
wire n10672; //CHANX 1 (9,3) #6
wire n10672_0;
wire n10673; //CHANX 1 (9,3) #7
wire n10673_0;
wire n10674; //CHANX 1 (9,3) #14
wire n10674_0;
wire n10675; //CHANX 1 (9,3) #15
wire n10675_0;
wire n10676; //CHANX 1 (9,3) #22
wire n10676_0;
wire n10677; //CHANX 1 (9,3) #23
wire n10677_0;
wire n10678; //CHANX 1 (9,3) #30
wire n10678_0;
wire n10679; //CHANX 1 (9,3) #31
wire n10679_0;
wire n10680; //CHANX 1 (9,3) #38
wire n10680_0;
wire n10681; //CHANX 1 (9,3) #39
wire n10681_0;
wire n10682; //CHANX 1 (9,3) #46
wire n10682_0;
wire n10683; //CHANX 1 (9,3) #47
wire n10683_0;
wire n10684; //CHANX 1 (9,3) #54
wire n10684_0;
wire n10685; //CHANX 1 (9,3) #55
wire n10685_0;
wire n10686; //CHANX 1 (9,3) #62
wire n10686_0;
wire n10687; //CHANX 1 (9,3) #63
wire n10687_0;
wire n10688; //CHANX 1 (9,3) #70
wire n10688_0;
wire n10689; //CHANX 1 (9,3) #71
wire n10689_0;
wire n10690; //CHANX 1 (9,3) #78
wire n10690_0;
wire n10691; //CHANX 1 (9,3) #79
wire n10691_0;
wire n10692; //CHANX 1 (9,3) #86
wire n10692_0;
wire n10693; //CHANX 1 (9,3) #87
wire n10693_0;
wire n10694; //CHANX 4 (1,4) #0
wire n10694_0;
wire n10694_1;
buffer_wire buffer_10694_1 (.in(n10694_0), .out(n10694_1));
wire n10695; //CHANX 4 (1,4) #1
wire n10695_0;
wire n10695_1;
buffer_wire buffer_10695_1 (.in(n10695_0), .out(n10695_1));
wire n10696; //CHANX 1 (1,4) #2
wire n10696_0;
wire n10697; //CHANX 1 (1,4) #3
wire n10697_0;
wire n10698; //CHANX 2 (1,4) #4
wire n10698_0;
wire n10699; //CHANX 2 (1,4) #5
wire n10699_0;
wire n10700; //CHANX 3 (1,4) #6
wire n10700_0;
wire n10701; //CHANX 3 (1,4) #7
wire n10701_0;
wire n10702; //CHANX 4 (1,4) #8
wire n10702_0;
wire n10702_1;
buffer_wire buffer_10702_1 (.in(n10702_0), .out(n10702_1));
wire n10703; //CHANX 4 (1,4) #9
wire n10703_0;
wire n10703_1;
buffer_wire buffer_10703_1 (.in(n10703_0), .out(n10703_1));
wire n10704; //CHANX 1 (1,4) #10
wire n10704_0;
wire n10705; //CHANX 1 (1,4) #11
wire n10705_0;
wire n10706; //CHANX 2 (1,4) #12
wire n10706_0;
wire n10707; //CHANX 2 (1,4) #13
wire n10707_0;
wire n10708; //CHANX 3 (1,4) #14
wire n10708_0;
wire n10709; //CHANX 3 (1,4) #15
wire n10709_0;
wire n10710; //CHANX 4 (1,4) #16
wire n10710_0;
wire n10710_1;
buffer_wire buffer_10710_1 (.in(n10710_0), .out(n10710_1));
wire n10711; //CHANX 4 (1,4) #17
wire n10711_0;
wire n10711_1;
buffer_wire buffer_10711_1 (.in(n10711_0), .out(n10711_1));
wire n10712; //CHANX 1 (1,4) #18
wire n10712_0;
wire n10713; //CHANX 1 (1,4) #19
wire n10713_0;
wire n10714; //CHANX 2 (1,4) #20
wire n10714_0;
wire n10715; //CHANX 2 (1,4) #21
wire n10715_0;
wire n10716; //CHANX 3 (1,4) #22
wire n10716_0;
wire n10717; //CHANX 3 (1,4) #23
wire n10717_0;
wire n10718; //CHANX 4 (1,4) #24
wire n10718_0;
wire n10718_1;
buffer_wire buffer_10718_1 (.in(n10718_0), .out(n10718_1));
wire n10719; //CHANX 4 (1,4) #25
wire n10719_0;
wire n10719_1;
buffer_wire buffer_10719_1 (.in(n10719_0), .out(n10719_1));
wire n10720; //CHANX 1 (1,4) #26
wire n10720_0;
wire n10721; //CHANX 1 (1,4) #27
wire n10721_0;
wire n10722; //CHANX 2 (1,4) #28
wire n10722_0;
wire n10723; //CHANX 2 (1,4) #29
wire n10723_0;
wire n10724; //CHANX 3 (1,4) #30
wire n10724_0;
wire n10725; //CHANX 3 (1,4) #31
wire n10725_0;
wire n10726; //CHANX 4 (1,4) #32
wire n10726_0;
wire n10726_1;
buffer_wire buffer_10726_1 (.in(n10726_0), .out(n10726_1));
wire n10727; //CHANX 4 (1,4) #33
wire n10727_0;
wire n10727_1;
buffer_wire buffer_10727_1 (.in(n10727_0), .out(n10727_1));
wire n10728; //CHANX 1 (1,4) #34
wire n10728_0;
wire n10729; //CHANX 1 (1,4) #35
wire n10729_0;
wire n10730; //CHANX 2 (1,4) #36
wire n10730_0;
wire n10731; //CHANX 2 (1,4) #37
wire n10731_0;
wire n10732; //CHANX 3 (1,4) #38
wire n10732_0;
wire n10733; //CHANX 3 (1,4) #39
wire n10733_0;
wire n10734; //CHANX 4 (1,4) #40
wire n10734_0;
wire n10734_1;
buffer_wire buffer_10734_1 (.in(n10734_0), .out(n10734_1));
wire n10735; //CHANX 4 (1,4) #41
wire n10735_0;
wire n10735_1;
buffer_wire buffer_10735_1 (.in(n10735_0), .out(n10735_1));
wire n10736; //CHANX 1 (1,4) #42
wire n10736_0;
wire n10737; //CHANX 1 (1,4) #43
wire n10737_0;
wire n10738; //CHANX 2 (1,4) #44
wire n10738_0;
wire n10739; //CHANX 2 (1,4) #45
wire n10739_0;
wire n10740; //CHANX 3 (1,4) #46
wire n10740_0;
wire n10741; //CHANX 3 (1,4) #47
wire n10741_0;
wire n10742; //CHANX 4 (1,4) #48
wire n10742_0;
wire n10742_1;
buffer_wire buffer_10742_1 (.in(n10742_0), .out(n10742_1));
wire n10743; //CHANX 4 (1,4) #49
wire n10743_0;
wire n10743_1;
buffer_wire buffer_10743_1 (.in(n10743_0), .out(n10743_1));
wire n10744; //CHANX 1 (1,4) #50
wire n10744_0;
wire n10745; //CHANX 1 (1,4) #51
wire n10745_0;
wire n10746; //CHANX 2 (1,4) #52
wire n10746_0;
wire n10747; //CHANX 2 (1,4) #53
wire n10747_0;
wire n10748; //CHANX 3 (1,4) #54
wire n10748_0;
wire n10749; //CHANX 3 (1,4) #55
wire n10749_0;
wire n10750; //CHANX 4 (1,4) #56
wire n10750_0;
wire n10750_1;
buffer_wire buffer_10750_1 (.in(n10750_0), .out(n10750_1));
wire n10751; //CHANX 4 (1,4) #57
wire n10751_0;
wire n10751_1;
buffer_wire buffer_10751_1 (.in(n10751_0), .out(n10751_1));
wire n10752; //CHANX 1 (1,4) #58
wire n10752_0;
wire n10753; //CHANX 1 (1,4) #59
wire n10753_0;
wire n10754; //CHANX 2 (1,4) #60
wire n10754_0;
wire n10755; //CHANX 2 (1,4) #61
wire n10755_0;
wire n10756; //CHANX 3 (1,4) #62
wire n10756_0;
wire n10757; //CHANX 3 (1,4) #63
wire n10757_0;
wire n10758; //CHANX 4 (1,4) #64
wire n10758_0;
wire n10758_1;
buffer_wire buffer_10758_1 (.in(n10758_0), .out(n10758_1));
wire n10759; //CHANX 4 (1,4) #65
wire n10759_0;
wire n10759_1;
buffer_wire buffer_10759_1 (.in(n10759_0), .out(n10759_1));
wire n10760; //CHANX 1 (1,4) #66
wire n10760_0;
wire n10761; //CHANX 1 (1,4) #67
wire n10761_0;
wire n10762; //CHANX 2 (1,4) #68
wire n10762_0;
wire n10763; //CHANX 2 (1,4) #69
wire n10763_0;
wire n10764; //CHANX 3 (1,4) #70
wire n10764_0;
wire n10765; //CHANX 3 (1,4) #71
wire n10765_0;
wire n10766; //CHANX 4 (1,4) #72
wire n10766_0;
wire n10766_1;
buffer_wire buffer_10766_1 (.in(n10766_0), .out(n10766_1));
wire n10767; //CHANX 4 (1,4) #73
wire n10767_0;
wire n10767_1;
buffer_wire buffer_10767_1 (.in(n10767_0), .out(n10767_1));
wire n10768; //CHANX 1 (1,4) #74
wire n10768_0;
wire n10769; //CHANX 1 (1,4) #75
wire n10769_0;
wire n10770; //CHANX 2 (1,4) #76
wire n10770_0;
wire n10771; //CHANX 2 (1,4) #77
wire n10771_0;
wire n10772; //CHANX 3 (1,4) #78
wire n10772_0;
wire n10773; //CHANX 3 (1,4) #79
wire n10773_0;
wire n10774; //CHANX 4 (1,4) #80
wire n10774_0;
wire n10774_1;
buffer_wire buffer_10774_1 (.in(n10774_0), .out(n10774_1));
wire n10775; //CHANX 4 (1,4) #81
wire n10775_0;
wire n10775_1;
buffer_wire buffer_10775_1 (.in(n10775_0), .out(n10775_1));
wire n10776; //CHANX 5 (1,4) #82
wire n10776_0;
wire n10776_1;
buffer_wire buffer_10776_1 (.in(n10776_0), .out(n10776_1));
wire n10777; //CHANX 5 (1,4) #83
wire n10777_0;
wire n10777_1;
buffer_wire buffer_10777_1 (.in(n10777_0), .out(n10777_1));
wire n10778; //CHANX 6 (1,4) #84
wire n10778_0;
wire n10778_1;
buffer_wire buffer_10778_1 (.in(n10778_0), .out(n10778_1));
wire n10779; //CHANX 6 (1,4) #85
wire n10779_0;
wire n10779_1;
buffer_wire buffer_10779_1 (.in(n10779_0), .out(n10779_1));
wire n10780; //CHANX 7 (1,4) #86
wire n10780_0;
wire n10780_1;
wire n10780_2;
buffer_wire buffer_10780_2 (.in(n10780_1), .out(n10780_2));
buffer_wire buffer_10780_1 (.in(n10780_0), .out(n10780_1));
wire n10781; //CHANX 7 (1,4) #87
wire n10781_0;
wire n10781_1;
wire n10781_2;
buffer_wire buffer_10781_2 (.in(n10781_1), .out(n10781_2));
buffer_wire buffer_10781_1 (.in(n10781_0), .out(n10781_1));
wire n10782; //CHANX 8 (1,4) #88
wire n10782_0;
wire n10782_1;
wire n10782_2;
buffer_wire buffer_10782_2 (.in(n10782_1), .out(n10782_2));
buffer_wire buffer_10782_1 (.in(n10782_0), .out(n10782_1));
wire n10783; //CHANX 8 (1,4) #89
wire n10783_0;
wire n10783_1;
wire n10783_2;
buffer_wire buffer_10783_2 (.in(n10783_1), .out(n10783_2));
buffer_wire buffer_10783_1 (.in(n10783_0), .out(n10783_1));
wire n10784; //CHANX 9 (1,4) #90
wire n10784_0;
wire n10784_1;
wire n10784_2;
buffer_wire buffer_10784_2 (.in(n10784_1), .out(n10784_2));
buffer_wire buffer_10784_1 (.in(n10784_0), .out(n10784_1));
wire n10785; //CHANX 9 (1,4) #91
wire n10785_0;
wire n10785_1;
wire n10785_2;
buffer_wire buffer_10785_2 (.in(n10785_1), .out(n10785_2));
buffer_wire buffer_10785_1 (.in(n10785_0), .out(n10785_1));
wire n10786; //CHANX 4 (2,4) #2
wire n10786_0;
wire n10786_1;
buffer_wire buffer_10786_1 (.in(n10786_0), .out(n10786_1));
wire n10787; //CHANX 4 (2,4) #3
wire n10787_0;
wire n10787_1;
buffer_wire buffer_10787_1 (.in(n10787_0), .out(n10787_1));
wire n10788; //CHANX 4 (2,4) #10
wire n10788_0;
wire n10788_1;
buffer_wire buffer_10788_1 (.in(n10788_0), .out(n10788_1));
wire n10789; //CHANX 4 (2,4) #11
wire n10789_0;
wire n10789_1;
buffer_wire buffer_10789_1 (.in(n10789_0), .out(n10789_1));
wire n10790; //CHANX 4 (2,4) #18
wire n10790_0;
wire n10790_1;
buffer_wire buffer_10790_1 (.in(n10790_0), .out(n10790_1));
wire n10791; //CHANX 4 (2,4) #19
wire n10791_0;
wire n10791_1;
buffer_wire buffer_10791_1 (.in(n10791_0), .out(n10791_1));
wire n10792; //CHANX 4 (2,4) #26
wire n10792_0;
wire n10792_1;
buffer_wire buffer_10792_1 (.in(n10792_0), .out(n10792_1));
wire n10793; //CHANX 4 (2,4) #27
wire n10793_0;
wire n10793_1;
buffer_wire buffer_10793_1 (.in(n10793_0), .out(n10793_1));
wire n10794; //CHANX 4 (2,4) #34
wire n10794_0;
wire n10794_1;
buffer_wire buffer_10794_1 (.in(n10794_0), .out(n10794_1));
wire n10795; //CHANX 4 (2,4) #35
wire n10795_0;
wire n10795_1;
buffer_wire buffer_10795_1 (.in(n10795_0), .out(n10795_1));
wire n10796; //CHANX 4 (2,4) #42
wire n10796_0;
wire n10796_1;
buffer_wire buffer_10796_1 (.in(n10796_0), .out(n10796_1));
wire n10797; //CHANX 4 (2,4) #43
wire n10797_0;
wire n10797_1;
buffer_wire buffer_10797_1 (.in(n10797_0), .out(n10797_1));
wire n10798; //CHANX 4 (2,4) #50
wire n10798_0;
wire n10798_1;
buffer_wire buffer_10798_1 (.in(n10798_0), .out(n10798_1));
wire n10799; //CHANX 4 (2,4) #51
wire n10799_0;
wire n10799_1;
buffer_wire buffer_10799_1 (.in(n10799_0), .out(n10799_1));
wire n10800; //CHANX 4 (2,4) #58
wire n10800_0;
wire n10800_1;
buffer_wire buffer_10800_1 (.in(n10800_0), .out(n10800_1));
wire n10801; //CHANX 4 (2,4) #59
wire n10801_0;
wire n10801_1;
buffer_wire buffer_10801_1 (.in(n10801_0), .out(n10801_1));
wire n10802; //CHANX 4 (2,4) #66
wire n10802_0;
wire n10802_1;
buffer_wire buffer_10802_1 (.in(n10802_0), .out(n10802_1));
wire n10803; //CHANX 4 (2,4) #67
wire n10803_0;
wire n10803_1;
buffer_wire buffer_10803_1 (.in(n10803_0), .out(n10803_1));
wire n10804; //CHANX 4 (2,4) #74
wire n10804_0;
wire n10804_1;
buffer_wire buffer_10804_1 (.in(n10804_0), .out(n10804_1));
wire n10805; //CHANX 4 (2,4) #75
wire n10805_0;
wire n10805_1;
buffer_wire buffer_10805_1 (.in(n10805_0), .out(n10805_1));
wire n10806; //CHANX 4 (3,4) #4
wire n10806_0;
wire n10806_1;
buffer_wire buffer_10806_1 (.in(n10806_0), .out(n10806_1));
wire n10807; //CHANX 4 (3,4) #5
wire n10807_0;
wire n10807_1;
buffer_wire buffer_10807_1 (.in(n10807_0), .out(n10807_1));
wire n10808; //CHANX 4 (3,4) #12
wire n10808_0;
wire n10808_1;
buffer_wire buffer_10808_1 (.in(n10808_0), .out(n10808_1));
wire n10809; //CHANX 4 (3,4) #13
wire n10809_0;
wire n10809_1;
buffer_wire buffer_10809_1 (.in(n10809_0), .out(n10809_1));
wire n10810; //CHANX 4 (3,4) #20
wire n10810_0;
wire n10810_1;
buffer_wire buffer_10810_1 (.in(n10810_0), .out(n10810_1));
wire n10811; //CHANX 4 (3,4) #21
wire n10811_0;
wire n10811_1;
buffer_wire buffer_10811_1 (.in(n10811_0), .out(n10811_1));
wire n10812; //CHANX 4 (3,4) #28
wire n10812_0;
wire n10812_1;
buffer_wire buffer_10812_1 (.in(n10812_0), .out(n10812_1));
wire n10813; //CHANX 4 (3,4) #29
wire n10813_0;
wire n10813_1;
buffer_wire buffer_10813_1 (.in(n10813_0), .out(n10813_1));
wire n10814; //CHANX 4 (3,4) #36
wire n10814_0;
wire n10814_1;
buffer_wire buffer_10814_1 (.in(n10814_0), .out(n10814_1));
wire n10815; //CHANX 4 (3,4) #37
wire n10815_0;
wire n10815_1;
buffer_wire buffer_10815_1 (.in(n10815_0), .out(n10815_1));
wire n10816; //CHANX 4 (3,4) #44
wire n10816_0;
wire n10816_1;
buffer_wire buffer_10816_1 (.in(n10816_0), .out(n10816_1));
wire n10817; //CHANX 4 (3,4) #45
wire n10817_0;
wire n10817_1;
buffer_wire buffer_10817_1 (.in(n10817_0), .out(n10817_1));
wire n10818; //CHANX 4 (3,4) #52
wire n10818_0;
wire n10818_1;
buffer_wire buffer_10818_1 (.in(n10818_0), .out(n10818_1));
wire n10819; //CHANX 4 (3,4) #53
wire n10819_0;
wire n10819_1;
buffer_wire buffer_10819_1 (.in(n10819_0), .out(n10819_1));
wire n10820; //CHANX 4 (3,4) #60
wire n10820_0;
wire n10820_1;
buffer_wire buffer_10820_1 (.in(n10820_0), .out(n10820_1));
wire n10821; //CHANX 4 (3,4) #61
wire n10821_0;
wire n10821_1;
buffer_wire buffer_10821_1 (.in(n10821_0), .out(n10821_1));
wire n10822; //CHANX 4 (3,4) #68
wire n10822_0;
wire n10822_1;
buffer_wire buffer_10822_1 (.in(n10822_0), .out(n10822_1));
wire n10823; //CHANX 4 (3,4) #69
wire n10823_0;
wire n10823_1;
buffer_wire buffer_10823_1 (.in(n10823_0), .out(n10823_1));
wire n10824; //CHANX 4 (3,4) #76
wire n10824_0;
wire n10824_1;
buffer_wire buffer_10824_1 (.in(n10824_0), .out(n10824_1));
wire n10825; //CHANX 4 (3,4) #77
wire n10825_0;
wire n10825_1;
buffer_wire buffer_10825_1 (.in(n10825_0), .out(n10825_1));
wire n10826; //CHANX 4 (4,4) #6
wire n10826_0;
wire n10826_1;
buffer_wire buffer_10826_1 (.in(n10826_0), .out(n10826_1));
wire n10827; //CHANX 4 (4,4) #7
wire n10827_0;
wire n10827_1;
buffer_wire buffer_10827_1 (.in(n10827_0), .out(n10827_1));
wire n10828; //CHANX 4 (4,4) #14
wire n10828_0;
wire n10828_1;
buffer_wire buffer_10828_1 (.in(n10828_0), .out(n10828_1));
wire n10829; //CHANX 4 (4,4) #15
wire n10829_0;
wire n10829_1;
buffer_wire buffer_10829_1 (.in(n10829_0), .out(n10829_1));
wire n10830; //CHANX 4 (4,4) #22
wire n10830_0;
wire n10830_1;
buffer_wire buffer_10830_1 (.in(n10830_0), .out(n10830_1));
wire n10831; //CHANX 4 (4,4) #23
wire n10831_0;
wire n10831_1;
buffer_wire buffer_10831_1 (.in(n10831_0), .out(n10831_1));
wire n10832; //CHANX 4 (4,4) #30
wire n10832_0;
wire n10832_1;
buffer_wire buffer_10832_1 (.in(n10832_0), .out(n10832_1));
wire n10833; //CHANX 4 (4,4) #31
wire n10833_0;
wire n10833_1;
buffer_wire buffer_10833_1 (.in(n10833_0), .out(n10833_1));
wire n10834; //CHANX 4 (4,4) #38
wire n10834_0;
wire n10834_1;
buffer_wire buffer_10834_1 (.in(n10834_0), .out(n10834_1));
wire n10835; //CHANX 4 (4,4) #39
wire n10835_0;
wire n10835_1;
buffer_wire buffer_10835_1 (.in(n10835_0), .out(n10835_1));
wire n10836; //CHANX 4 (4,4) #46
wire n10836_0;
wire n10836_1;
buffer_wire buffer_10836_1 (.in(n10836_0), .out(n10836_1));
wire n10837; //CHANX 4 (4,4) #47
wire n10837_0;
wire n10837_1;
buffer_wire buffer_10837_1 (.in(n10837_0), .out(n10837_1));
wire n10838; //CHANX 4 (4,4) #54
wire n10838_0;
wire n10838_1;
buffer_wire buffer_10838_1 (.in(n10838_0), .out(n10838_1));
wire n10839; //CHANX 4 (4,4) #55
wire n10839_0;
wire n10839_1;
buffer_wire buffer_10839_1 (.in(n10839_0), .out(n10839_1));
wire n10840; //CHANX 4 (4,4) #62
wire n10840_0;
wire n10840_1;
buffer_wire buffer_10840_1 (.in(n10840_0), .out(n10840_1));
wire n10841; //CHANX 4 (4,4) #63
wire n10841_0;
wire n10841_1;
buffer_wire buffer_10841_1 (.in(n10841_0), .out(n10841_1));
wire n10842; //CHANX 4 (4,4) #70
wire n10842_0;
wire n10842_1;
buffer_wire buffer_10842_1 (.in(n10842_0), .out(n10842_1));
wire n10843; //CHANX 4 (4,4) #71
wire n10843_0;
wire n10843_1;
buffer_wire buffer_10843_1 (.in(n10843_0), .out(n10843_1));
wire n10844; //CHANX 4 (4,4) #78
wire n10844_0;
wire n10844_1;
buffer_wire buffer_10844_1 (.in(n10844_0), .out(n10844_1));
wire n10845; //CHANX 4 (4,4) #79
wire n10845_0;
wire n10845_1;
buffer_wire buffer_10845_1 (.in(n10845_0), .out(n10845_1));
wire n10846; //CHANX 4 (5,4) #0
wire n10846_0;
wire n10846_1;
buffer_wire buffer_10846_1 (.in(n10846_0), .out(n10846_1));
wire n10847; //CHANX 4 (5,4) #1
wire n10847_0;
wire n10847_1;
buffer_wire buffer_10847_1 (.in(n10847_0), .out(n10847_1));
wire n10848; //CHANX 4 (5,4) #8
wire n10848_0;
wire n10848_1;
buffer_wire buffer_10848_1 (.in(n10848_0), .out(n10848_1));
wire n10849; //CHANX 4 (5,4) #9
wire n10849_0;
wire n10849_1;
buffer_wire buffer_10849_1 (.in(n10849_0), .out(n10849_1));
wire n10850; //CHANX 4 (5,4) #16
wire n10850_0;
wire n10850_1;
buffer_wire buffer_10850_1 (.in(n10850_0), .out(n10850_1));
wire n10851; //CHANX 4 (5,4) #17
wire n10851_0;
wire n10851_1;
buffer_wire buffer_10851_1 (.in(n10851_0), .out(n10851_1));
wire n10852; //CHANX 4 (5,4) #24
wire n10852_0;
wire n10852_1;
buffer_wire buffer_10852_1 (.in(n10852_0), .out(n10852_1));
wire n10853; //CHANX 4 (5,4) #25
wire n10853_0;
wire n10853_1;
buffer_wire buffer_10853_1 (.in(n10853_0), .out(n10853_1));
wire n10854; //CHANX 4 (5,4) #32
wire n10854_0;
wire n10854_1;
buffer_wire buffer_10854_1 (.in(n10854_0), .out(n10854_1));
wire n10855; //CHANX 4 (5,4) #33
wire n10855_0;
wire n10855_1;
buffer_wire buffer_10855_1 (.in(n10855_0), .out(n10855_1));
wire n10856; //CHANX 4 (5,4) #40
wire n10856_0;
wire n10856_1;
buffer_wire buffer_10856_1 (.in(n10856_0), .out(n10856_1));
wire n10857; //CHANX 4 (5,4) #41
wire n10857_0;
wire n10857_1;
buffer_wire buffer_10857_1 (.in(n10857_0), .out(n10857_1));
wire n10858; //CHANX 4 (5,4) #48
wire n10858_0;
wire n10858_1;
buffer_wire buffer_10858_1 (.in(n10858_0), .out(n10858_1));
wire n10859; //CHANX 4 (5,4) #49
wire n10859_0;
wire n10859_1;
buffer_wire buffer_10859_1 (.in(n10859_0), .out(n10859_1));
wire n10860; //CHANX 4 (5,4) #56
wire n10860_0;
wire n10860_1;
buffer_wire buffer_10860_1 (.in(n10860_0), .out(n10860_1));
wire n10861; //CHANX 4 (5,4) #57
wire n10861_0;
wire n10861_1;
buffer_wire buffer_10861_1 (.in(n10861_0), .out(n10861_1));
wire n10862; //CHANX 4 (5,4) #64
wire n10862_0;
wire n10862_1;
buffer_wire buffer_10862_1 (.in(n10862_0), .out(n10862_1));
wire n10863; //CHANX 4 (5,4) #65
wire n10863_0;
wire n10863_1;
buffer_wire buffer_10863_1 (.in(n10863_0), .out(n10863_1));
wire n10864; //CHANX 4 (5,4) #72
wire n10864_0;
wire n10864_1;
buffer_wire buffer_10864_1 (.in(n10864_0), .out(n10864_1));
wire n10865; //CHANX 4 (5,4) #73
wire n10865_0;
wire n10865_1;
buffer_wire buffer_10865_1 (.in(n10865_0), .out(n10865_1));
wire n10866; //CHANX 5 (5,4) #80
wire n10866_0;
wire n10866_1;
buffer_wire buffer_10866_1 (.in(n10866_0), .out(n10866_1));
wire n10867; //CHANX 5 (5,4) #81
wire n10867_0;
wire n10867_1;
buffer_wire buffer_10867_1 (.in(n10867_0), .out(n10867_1));
wire n10868; //CHANX 4 (6,4) #2
wire n10868_0;
wire n10868_1;
buffer_wire buffer_10868_1 (.in(n10868_0), .out(n10868_1));
wire n10869; //CHANX 4 (6,4) #3
wire n10869_0;
wire n10869_1;
buffer_wire buffer_10869_1 (.in(n10869_0), .out(n10869_1));
wire n10870; //CHANX 4 (6,4) #10
wire n10870_0;
wire n10870_1;
buffer_wire buffer_10870_1 (.in(n10870_0), .out(n10870_1));
wire n10871; //CHANX 4 (6,4) #11
wire n10871_0;
wire n10871_1;
buffer_wire buffer_10871_1 (.in(n10871_0), .out(n10871_1));
wire n10872; //CHANX 4 (6,4) #18
wire n10872_0;
wire n10872_1;
buffer_wire buffer_10872_1 (.in(n10872_0), .out(n10872_1));
wire n10873; //CHANX 4 (6,4) #19
wire n10873_0;
wire n10873_1;
buffer_wire buffer_10873_1 (.in(n10873_0), .out(n10873_1));
wire n10874; //CHANX 4 (6,4) #26
wire n10874_0;
wire n10874_1;
buffer_wire buffer_10874_1 (.in(n10874_0), .out(n10874_1));
wire n10875; //CHANX 4 (6,4) #27
wire n10875_0;
wire n10875_1;
buffer_wire buffer_10875_1 (.in(n10875_0), .out(n10875_1));
wire n10876; //CHANX 4 (6,4) #34
wire n10876_0;
wire n10876_1;
buffer_wire buffer_10876_1 (.in(n10876_0), .out(n10876_1));
wire n10877; //CHANX 4 (6,4) #35
wire n10877_0;
wire n10877_1;
buffer_wire buffer_10877_1 (.in(n10877_0), .out(n10877_1));
wire n10878; //CHANX 4 (6,4) #42
wire n10878_0;
wire n10878_1;
buffer_wire buffer_10878_1 (.in(n10878_0), .out(n10878_1));
wire n10879; //CHANX 4 (6,4) #43
wire n10879_0;
wire n10879_1;
buffer_wire buffer_10879_1 (.in(n10879_0), .out(n10879_1));
wire n10880; //CHANX 4 (6,4) #50
wire n10880_0;
wire n10880_1;
buffer_wire buffer_10880_1 (.in(n10880_0), .out(n10880_1));
wire n10881; //CHANX 4 (6,4) #51
wire n10881_0;
wire n10881_1;
buffer_wire buffer_10881_1 (.in(n10881_0), .out(n10881_1));
wire n10882; //CHANX 4 (6,4) #58
wire n10882_0;
wire n10882_1;
buffer_wire buffer_10882_1 (.in(n10882_0), .out(n10882_1));
wire n10883; //CHANX 4 (6,4) #59
wire n10883_0;
wire n10883_1;
buffer_wire buffer_10883_1 (.in(n10883_0), .out(n10883_1));
wire n10884; //CHANX 4 (6,4) #66
wire n10884_0;
wire n10884_1;
buffer_wire buffer_10884_1 (.in(n10884_0), .out(n10884_1));
wire n10885; //CHANX 4 (6,4) #67
wire n10885_0;
wire n10885_1;
buffer_wire buffer_10885_1 (.in(n10885_0), .out(n10885_1));
wire n10886; //CHANX 4 (6,4) #74
wire n10886_0;
wire n10886_1;
buffer_wire buffer_10886_1 (.in(n10886_0), .out(n10886_1));
wire n10887; //CHANX 4 (6,4) #75
wire n10887_0;
wire n10887_1;
buffer_wire buffer_10887_1 (.in(n10887_0), .out(n10887_1));
wire n10888; //CHANX 4 (6,4) #82
wire n10888_0;
wire n10888_1;
buffer_wire buffer_10888_1 (.in(n10888_0), .out(n10888_1));
wire n10889; //CHANX 4 (6,4) #83
wire n10889_0;
wire n10889_1;
buffer_wire buffer_10889_1 (.in(n10889_0), .out(n10889_1));
wire n10890; //CHANX 3 (7,4) #4
wire n10890_0;
wire n10891; //CHANX 3 (7,4) #5
wire n10891_0;
wire n10892; //CHANX 3 (7,4) #12
wire n10892_0;
wire n10893; //CHANX 3 (7,4) #13
wire n10893_0;
wire n10894; //CHANX 3 (7,4) #20
wire n10894_0;
wire n10895; //CHANX 3 (7,4) #21
wire n10895_0;
wire n10896; //CHANX 3 (7,4) #28
wire n10896_0;
wire n10897; //CHANX 3 (7,4) #29
wire n10897_0;
wire n10898; //CHANX 3 (7,4) #36
wire n10898_0;
wire n10899; //CHANX 3 (7,4) #37
wire n10899_0;
wire n10900; //CHANX 3 (7,4) #44
wire n10900_0;
wire n10901; //CHANX 3 (7,4) #45
wire n10901_0;
wire n10902; //CHANX 3 (7,4) #52
wire n10902_0;
wire n10903; //CHANX 3 (7,4) #53
wire n10903_0;
wire n10904; //CHANX 3 (7,4) #60
wire n10904_0;
wire n10905; //CHANX 3 (7,4) #61
wire n10905_0;
wire n10906; //CHANX 3 (7,4) #68
wire n10906_0;
wire n10907; //CHANX 3 (7,4) #69
wire n10907_0;
wire n10908; //CHANX 3 (7,4) #76
wire n10908_0;
wire n10909; //CHANX 3 (7,4) #77
wire n10909_0;
wire n10910; //CHANX 3 (7,4) #84
wire n10910_0;
wire n10911; //CHANX 3 (7,4) #85
wire n10911_0;
wire n10912; //CHANX 2 (8,4) #6
wire n10912_0;
wire n10913; //CHANX 2 (8,4) #7
wire n10913_0;
wire n10914; //CHANX 2 (8,4) #14
wire n10914_0;
wire n10915; //CHANX 2 (8,4) #15
wire n10915_0;
wire n10916; //CHANX 2 (8,4) #22
wire n10916_0;
wire n10917; //CHANX 2 (8,4) #23
wire n10917_0;
wire n10918; //CHANX 2 (8,4) #30
wire n10918_0;
wire n10919; //CHANX 2 (8,4) #31
wire n10919_0;
wire n10920; //CHANX 2 (8,4) #38
wire n10920_0;
wire n10921; //CHANX 2 (8,4) #39
wire n10921_0;
wire n10922; //CHANX 2 (8,4) #46
wire n10922_0;
wire n10923; //CHANX 2 (8,4) #47
wire n10923_0;
wire n10924; //CHANX 2 (8,4) #54
wire n10924_0;
wire n10925; //CHANX 2 (8,4) #55
wire n10925_0;
wire n10926; //CHANX 2 (8,4) #62
wire n10926_0;
wire n10927; //CHANX 2 (8,4) #63
wire n10927_0;
wire n10928; //CHANX 2 (8,4) #70
wire n10928_0;
wire n10929; //CHANX 2 (8,4) #71
wire n10929_0;
wire n10930; //CHANX 2 (8,4) #78
wire n10930_0;
wire n10931; //CHANX 2 (8,4) #79
wire n10931_0;
wire n10932; //CHANX 2 (8,4) #86
wire n10932_0;
wire n10933; //CHANX 2 (8,4) #87
wire n10933_0;
wire n10934; //CHANX 1 (9,4) #0
wire n10934_0;
wire n10935; //CHANX 1 (9,4) #1
wire n10935_0;
wire n10936; //CHANX 1 (9,4) #8
wire n10936_0;
wire n10937; //CHANX 1 (9,4) #9
wire n10937_0;
wire n10938; //CHANX 1 (9,4) #16
wire n10938_0;
wire n10939; //CHANX 1 (9,4) #17
wire n10939_0;
wire n10940; //CHANX 1 (9,4) #24
wire n10940_0;
wire n10941; //CHANX 1 (9,4) #25
wire n10941_0;
wire n10942; //CHANX 1 (9,4) #32
wire n10942_0;
wire n10943; //CHANX 1 (9,4) #33
wire n10943_0;
wire n10944; //CHANX 1 (9,4) #40
wire n10944_0;
wire n10945; //CHANX 1 (9,4) #41
wire n10945_0;
wire n10946; //CHANX 1 (9,4) #48
wire n10946_0;
wire n10947; //CHANX 1 (9,4) #49
wire n10947_0;
wire n10948; //CHANX 1 (9,4) #56
wire n10948_0;
wire n10949; //CHANX 1 (9,4) #57
wire n10949_0;
wire n10950; //CHANX 1 (9,4) #64
wire n10950_0;
wire n10951; //CHANX 1 (9,4) #65
wire n10951_0;
wire n10952; //CHANX 1 (9,4) #72
wire n10952_0;
wire n10953; //CHANX 1 (9,4) #73
wire n10953_0;
wire n10954; //CHANX 1 (9,4) #88
wire n10954_0;
wire n10955; //CHANX 1 (9,4) #89
wire n10955_0;
wire n10956; //CHANX 3 (1,5) #0
wire n10956_0;
wire n10957; //CHANX 3 (1,5) #1
wire n10957_0;
wire n10958; //CHANX 4 (1,5) #2
wire n10958_0;
wire n10958_1;
buffer_wire buffer_10958_1 (.in(n10958_0), .out(n10958_1));
wire n10959; //CHANX 4 (1,5) #3
wire n10959_0;
wire n10959_1;
buffer_wire buffer_10959_1 (.in(n10959_0), .out(n10959_1));
wire n10960; //CHANX 1 (1,5) #4
wire n10960_0;
wire n10961; //CHANX 1 (1,5) #5
wire n10961_0;
wire n10962; //CHANX 2 (1,5) #6
wire n10962_0;
wire n10963; //CHANX 2 (1,5) #7
wire n10963_0;
wire n10964; //CHANX 3 (1,5) #8
wire n10964_0;
wire n10965; //CHANX 3 (1,5) #9
wire n10965_0;
wire n10966; //CHANX 4 (1,5) #10
wire n10966_0;
wire n10966_1;
buffer_wire buffer_10966_1 (.in(n10966_0), .out(n10966_1));
wire n10967; //CHANX 4 (1,5) #11
wire n10967_0;
wire n10967_1;
buffer_wire buffer_10967_1 (.in(n10967_0), .out(n10967_1));
wire n10968; //CHANX 1 (1,5) #12
wire n10968_0;
wire n10969; //CHANX 1 (1,5) #13
wire n10969_0;
wire n10970; //CHANX 2 (1,5) #14
wire n10970_0;
wire n10971; //CHANX 2 (1,5) #15
wire n10971_0;
wire n10972; //CHANX 3 (1,5) #16
wire n10972_0;
wire n10973; //CHANX 3 (1,5) #17
wire n10973_0;
wire n10974; //CHANX 4 (1,5) #18
wire n10974_0;
wire n10974_1;
buffer_wire buffer_10974_1 (.in(n10974_0), .out(n10974_1));
wire n10975; //CHANX 4 (1,5) #19
wire n10975_0;
wire n10975_1;
buffer_wire buffer_10975_1 (.in(n10975_0), .out(n10975_1));
wire n10976; //CHANX 1 (1,5) #20
wire n10976_0;
wire n10977; //CHANX 1 (1,5) #21
wire n10977_0;
wire n10978; //CHANX 2 (1,5) #22
wire n10978_0;
wire n10979; //CHANX 2 (1,5) #23
wire n10979_0;
wire n10980; //CHANX 3 (1,5) #24
wire n10980_0;
wire n10981; //CHANX 3 (1,5) #25
wire n10981_0;
wire n10982; //CHANX 4 (1,5) #26
wire n10982_0;
wire n10982_1;
buffer_wire buffer_10982_1 (.in(n10982_0), .out(n10982_1));
wire n10983; //CHANX 4 (1,5) #27
wire n10983_0;
wire n10983_1;
buffer_wire buffer_10983_1 (.in(n10983_0), .out(n10983_1));
wire n10984; //CHANX 1 (1,5) #28
wire n10984_0;
wire n10985; //CHANX 1 (1,5) #29
wire n10985_0;
wire n10986; //CHANX 2 (1,5) #30
wire n10986_0;
wire n10987; //CHANX 2 (1,5) #31
wire n10987_0;
wire n10988; //CHANX 3 (1,5) #32
wire n10988_0;
wire n10989; //CHANX 3 (1,5) #33
wire n10989_0;
wire n10990; //CHANX 4 (1,5) #34
wire n10990_0;
wire n10990_1;
buffer_wire buffer_10990_1 (.in(n10990_0), .out(n10990_1));
wire n10991; //CHANX 4 (1,5) #35
wire n10991_0;
wire n10991_1;
buffer_wire buffer_10991_1 (.in(n10991_0), .out(n10991_1));
wire n10992; //CHANX 1 (1,5) #36
wire n10992_0;
wire n10993; //CHANX 1 (1,5) #37
wire n10993_0;
wire n10994; //CHANX 2 (1,5) #38
wire n10994_0;
wire n10995; //CHANX 2 (1,5) #39
wire n10995_0;
wire n10996; //CHANX 3 (1,5) #40
wire n10996_0;
wire n10997; //CHANX 3 (1,5) #41
wire n10997_0;
wire n10998; //CHANX 4 (1,5) #42
wire n10998_0;
wire n10998_1;
buffer_wire buffer_10998_1 (.in(n10998_0), .out(n10998_1));
wire n10999; //CHANX 4 (1,5) #43
wire n10999_0;
wire n10999_1;
buffer_wire buffer_10999_1 (.in(n10999_0), .out(n10999_1));
wire n11000; //CHANX 1 (1,5) #44
wire n11000_0;
wire n11001; //CHANX 1 (1,5) #45
wire n11001_0;
wire n11002; //CHANX 2 (1,5) #46
wire n11002_0;
wire n11003; //CHANX 2 (1,5) #47
wire n11003_0;
wire n11004; //CHANX 3 (1,5) #48
wire n11004_0;
wire n11005; //CHANX 3 (1,5) #49
wire n11005_0;
wire n11006; //CHANX 4 (1,5) #50
wire n11006_0;
wire n11006_1;
buffer_wire buffer_11006_1 (.in(n11006_0), .out(n11006_1));
wire n11007; //CHANX 4 (1,5) #51
wire n11007_0;
wire n11007_1;
buffer_wire buffer_11007_1 (.in(n11007_0), .out(n11007_1));
wire n11008; //CHANX 1 (1,5) #52
wire n11008_0;
wire n11009; //CHANX 1 (1,5) #53
wire n11009_0;
wire n11010; //CHANX 2 (1,5) #54
wire n11010_0;
wire n11011; //CHANX 2 (1,5) #55
wire n11011_0;
wire n11012; //CHANX 3 (1,5) #56
wire n11012_0;
wire n11013; //CHANX 3 (1,5) #57
wire n11013_0;
wire n11014; //CHANX 4 (1,5) #58
wire n11014_0;
wire n11014_1;
buffer_wire buffer_11014_1 (.in(n11014_0), .out(n11014_1));
wire n11015; //CHANX 4 (1,5) #59
wire n11015_0;
wire n11015_1;
buffer_wire buffer_11015_1 (.in(n11015_0), .out(n11015_1));
wire n11016; //CHANX 1 (1,5) #60
wire n11016_0;
wire n11017; //CHANX 1 (1,5) #61
wire n11017_0;
wire n11018; //CHANX 2 (1,5) #62
wire n11018_0;
wire n11019; //CHANX 2 (1,5) #63
wire n11019_0;
wire n11020; //CHANX 3 (1,5) #64
wire n11020_0;
wire n11021; //CHANX 3 (1,5) #65
wire n11021_0;
wire n11022; //CHANX 4 (1,5) #66
wire n11022_0;
wire n11022_1;
buffer_wire buffer_11022_1 (.in(n11022_0), .out(n11022_1));
wire n11023; //CHANX 4 (1,5) #67
wire n11023_0;
wire n11023_1;
buffer_wire buffer_11023_1 (.in(n11023_0), .out(n11023_1));
wire n11024; //CHANX 1 (1,5) #68
wire n11024_0;
wire n11025; //CHANX 1 (1,5) #69
wire n11025_0;
wire n11026; //CHANX 2 (1,5) #70
wire n11026_0;
wire n11027; //CHANX 2 (1,5) #71
wire n11027_0;
wire n11028; //CHANX 3 (1,5) #72
wire n11028_0;
wire n11029; //CHANX 3 (1,5) #73
wire n11029_0;
wire n11030; //CHANX 4 (1,5) #74
wire n11030_0;
wire n11030_1;
buffer_wire buffer_11030_1 (.in(n11030_0), .out(n11030_1));
wire n11031; //CHANX 4 (1,5) #75
wire n11031_0;
wire n11031_1;
buffer_wire buffer_11031_1 (.in(n11031_0), .out(n11031_1));
wire n11032; //CHANX 1 (1,5) #76
wire n11032_0;
wire n11033; //CHANX 1 (1,5) #77
wire n11033_0;
wire n11034; //CHANX 2 (1,5) #78
wire n11034_0;
wire n11035; //CHANX 2 (1,5) #79
wire n11035_0;
wire n11036; //CHANX 3 (1,5) #80
wire n11036_0;
wire n11037; //CHANX 3 (1,5) #81
wire n11037_0;
wire n11038; //CHANX 4 (1,5) #82
wire n11038_0;
wire n11038_1;
buffer_wire buffer_11038_1 (.in(n11038_0), .out(n11038_1));
wire n11039; //CHANX 4 (1,5) #83
wire n11039_0;
wire n11039_1;
buffer_wire buffer_11039_1 (.in(n11039_0), .out(n11039_1));
wire n11040; //CHANX 5 (1,5) #84
wire n11040_0;
wire n11040_1;
buffer_wire buffer_11040_1 (.in(n11040_0), .out(n11040_1));
wire n11041; //CHANX 5 (1,5) #85
wire n11041_0;
wire n11041_1;
buffer_wire buffer_11041_1 (.in(n11041_0), .out(n11041_1));
wire n11042; //CHANX 6 (1,5) #86
wire n11042_0;
wire n11042_1;
buffer_wire buffer_11042_1 (.in(n11042_0), .out(n11042_1));
wire n11043; //CHANX 6 (1,5) #87
wire n11043_0;
wire n11043_1;
buffer_wire buffer_11043_1 (.in(n11043_0), .out(n11043_1));
wire n11044; //CHANX 7 (1,5) #88
wire n11044_0;
wire n11044_1;
wire n11044_2;
buffer_wire buffer_11044_2 (.in(n11044_1), .out(n11044_2));
buffer_wire buffer_11044_1 (.in(n11044_0), .out(n11044_1));
wire n11045; //CHANX 7 (1,5) #89
wire n11045_0;
wire n11045_1;
wire n11045_2;
buffer_wire buffer_11045_2 (.in(n11045_1), .out(n11045_2));
buffer_wire buffer_11045_1 (.in(n11045_0), .out(n11045_1));
wire n11046; //CHANX 8 (1,5) #90
wire n11046_0;
wire n11046_1;
wire n11046_2;
buffer_wire buffer_11046_2 (.in(n11046_1), .out(n11046_2));
buffer_wire buffer_11046_1 (.in(n11046_0), .out(n11046_1));
wire n11047; //CHANX 8 (1,5) #91
wire n11047_0;
wire n11047_1;
wire n11047_2;
buffer_wire buffer_11047_2 (.in(n11047_1), .out(n11047_2));
buffer_wire buffer_11047_1 (.in(n11047_0), .out(n11047_1));
wire n11048; //CHANX 4 (2,5) #4
wire n11048_0;
wire n11048_1;
buffer_wire buffer_11048_1 (.in(n11048_0), .out(n11048_1));
wire n11049; //CHANX 4 (2,5) #5
wire n11049_0;
wire n11049_1;
buffer_wire buffer_11049_1 (.in(n11049_0), .out(n11049_1));
wire n11050; //CHANX 4 (2,5) #12
wire n11050_0;
wire n11050_1;
buffer_wire buffer_11050_1 (.in(n11050_0), .out(n11050_1));
wire n11051; //CHANX 4 (2,5) #13
wire n11051_0;
wire n11051_1;
buffer_wire buffer_11051_1 (.in(n11051_0), .out(n11051_1));
wire n11052; //CHANX 4 (2,5) #20
wire n11052_0;
wire n11052_1;
buffer_wire buffer_11052_1 (.in(n11052_0), .out(n11052_1));
wire n11053; //CHANX 4 (2,5) #21
wire n11053_0;
wire n11053_1;
buffer_wire buffer_11053_1 (.in(n11053_0), .out(n11053_1));
wire n11054; //CHANX 4 (2,5) #28
wire n11054_0;
wire n11054_1;
buffer_wire buffer_11054_1 (.in(n11054_0), .out(n11054_1));
wire n11055; //CHANX 4 (2,5) #29
wire n11055_0;
wire n11055_1;
buffer_wire buffer_11055_1 (.in(n11055_0), .out(n11055_1));
wire n11056; //CHANX 4 (2,5) #36
wire n11056_0;
wire n11056_1;
buffer_wire buffer_11056_1 (.in(n11056_0), .out(n11056_1));
wire n11057; //CHANX 4 (2,5) #37
wire n11057_0;
wire n11057_1;
buffer_wire buffer_11057_1 (.in(n11057_0), .out(n11057_1));
wire n11058; //CHANX 4 (2,5) #44
wire n11058_0;
wire n11058_1;
buffer_wire buffer_11058_1 (.in(n11058_0), .out(n11058_1));
wire n11059; //CHANX 4 (2,5) #45
wire n11059_0;
wire n11059_1;
buffer_wire buffer_11059_1 (.in(n11059_0), .out(n11059_1));
wire n11060; //CHANX 4 (2,5) #52
wire n11060_0;
wire n11060_1;
buffer_wire buffer_11060_1 (.in(n11060_0), .out(n11060_1));
wire n11061; //CHANX 4 (2,5) #53
wire n11061_0;
wire n11061_1;
buffer_wire buffer_11061_1 (.in(n11061_0), .out(n11061_1));
wire n11062; //CHANX 4 (2,5) #60
wire n11062_0;
wire n11062_1;
buffer_wire buffer_11062_1 (.in(n11062_0), .out(n11062_1));
wire n11063; //CHANX 4 (2,5) #61
wire n11063_0;
wire n11063_1;
buffer_wire buffer_11063_1 (.in(n11063_0), .out(n11063_1));
wire n11064; //CHANX 4 (2,5) #68
wire n11064_0;
wire n11064_1;
buffer_wire buffer_11064_1 (.in(n11064_0), .out(n11064_1));
wire n11065; //CHANX 4 (2,5) #69
wire n11065_0;
wire n11065_1;
buffer_wire buffer_11065_1 (.in(n11065_0), .out(n11065_1));
wire n11066; //CHANX 4 (2,5) #76
wire n11066_0;
wire n11066_1;
buffer_wire buffer_11066_1 (.in(n11066_0), .out(n11066_1));
wire n11067; //CHANX 4 (2,5) #77
wire n11067_0;
wire n11067_1;
buffer_wire buffer_11067_1 (.in(n11067_0), .out(n11067_1));
wire n11068; //CHANX 4 (3,5) #6
wire n11068_0;
wire n11068_1;
buffer_wire buffer_11068_1 (.in(n11068_0), .out(n11068_1));
wire n11069; //CHANX 4 (3,5) #7
wire n11069_0;
wire n11069_1;
buffer_wire buffer_11069_1 (.in(n11069_0), .out(n11069_1));
wire n11070; //CHANX 4 (3,5) #14
wire n11070_0;
wire n11070_1;
buffer_wire buffer_11070_1 (.in(n11070_0), .out(n11070_1));
wire n11071; //CHANX 4 (3,5) #15
wire n11071_0;
wire n11071_1;
buffer_wire buffer_11071_1 (.in(n11071_0), .out(n11071_1));
wire n11072; //CHANX 4 (3,5) #22
wire n11072_0;
wire n11072_1;
buffer_wire buffer_11072_1 (.in(n11072_0), .out(n11072_1));
wire n11073; //CHANX 4 (3,5) #23
wire n11073_0;
wire n11073_1;
buffer_wire buffer_11073_1 (.in(n11073_0), .out(n11073_1));
wire n11074; //CHANX 4 (3,5) #30
wire n11074_0;
wire n11074_1;
buffer_wire buffer_11074_1 (.in(n11074_0), .out(n11074_1));
wire n11075; //CHANX 4 (3,5) #31
wire n11075_0;
wire n11075_1;
buffer_wire buffer_11075_1 (.in(n11075_0), .out(n11075_1));
wire n11076; //CHANX 4 (3,5) #38
wire n11076_0;
wire n11076_1;
buffer_wire buffer_11076_1 (.in(n11076_0), .out(n11076_1));
wire n11077; //CHANX 4 (3,5) #39
wire n11077_0;
wire n11077_1;
buffer_wire buffer_11077_1 (.in(n11077_0), .out(n11077_1));
wire n11078; //CHANX 4 (3,5) #46
wire n11078_0;
wire n11078_1;
buffer_wire buffer_11078_1 (.in(n11078_0), .out(n11078_1));
wire n11079; //CHANX 4 (3,5) #47
wire n11079_0;
wire n11079_1;
buffer_wire buffer_11079_1 (.in(n11079_0), .out(n11079_1));
wire n11080; //CHANX 4 (3,5) #54
wire n11080_0;
wire n11080_1;
buffer_wire buffer_11080_1 (.in(n11080_0), .out(n11080_1));
wire n11081; //CHANX 4 (3,5) #55
wire n11081_0;
wire n11081_1;
buffer_wire buffer_11081_1 (.in(n11081_0), .out(n11081_1));
wire n11082; //CHANX 4 (3,5) #62
wire n11082_0;
wire n11082_1;
buffer_wire buffer_11082_1 (.in(n11082_0), .out(n11082_1));
wire n11083; //CHANX 4 (3,5) #63
wire n11083_0;
wire n11083_1;
buffer_wire buffer_11083_1 (.in(n11083_0), .out(n11083_1));
wire n11084; //CHANX 4 (3,5) #70
wire n11084_0;
wire n11084_1;
buffer_wire buffer_11084_1 (.in(n11084_0), .out(n11084_1));
wire n11085; //CHANX 4 (3,5) #71
wire n11085_0;
wire n11085_1;
buffer_wire buffer_11085_1 (.in(n11085_0), .out(n11085_1));
wire n11086; //CHANX 4 (3,5) #78
wire n11086_0;
wire n11086_1;
buffer_wire buffer_11086_1 (.in(n11086_0), .out(n11086_1));
wire n11087; //CHANX 4 (3,5) #79
wire n11087_0;
wire n11087_1;
buffer_wire buffer_11087_1 (.in(n11087_0), .out(n11087_1));
wire n11088; //CHANX 4 (4,5) #0
wire n11088_0;
wire n11088_1;
buffer_wire buffer_11088_1 (.in(n11088_0), .out(n11088_1));
wire n11089; //CHANX 4 (4,5) #1
wire n11089_0;
wire n11089_1;
buffer_wire buffer_11089_1 (.in(n11089_0), .out(n11089_1));
wire n11090; //CHANX 4 (4,5) #8
wire n11090_0;
wire n11090_1;
buffer_wire buffer_11090_1 (.in(n11090_0), .out(n11090_1));
wire n11091; //CHANX 4 (4,5) #9
wire n11091_0;
wire n11091_1;
buffer_wire buffer_11091_1 (.in(n11091_0), .out(n11091_1));
wire n11092; //CHANX 4 (4,5) #16
wire n11092_0;
wire n11092_1;
buffer_wire buffer_11092_1 (.in(n11092_0), .out(n11092_1));
wire n11093; //CHANX 4 (4,5) #17
wire n11093_0;
wire n11093_1;
buffer_wire buffer_11093_1 (.in(n11093_0), .out(n11093_1));
wire n11094; //CHANX 4 (4,5) #24
wire n11094_0;
wire n11094_1;
buffer_wire buffer_11094_1 (.in(n11094_0), .out(n11094_1));
wire n11095; //CHANX 4 (4,5) #25
wire n11095_0;
wire n11095_1;
buffer_wire buffer_11095_1 (.in(n11095_0), .out(n11095_1));
wire n11096; //CHANX 4 (4,5) #32
wire n11096_0;
wire n11096_1;
buffer_wire buffer_11096_1 (.in(n11096_0), .out(n11096_1));
wire n11097; //CHANX 4 (4,5) #33
wire n11097_0;
wire n11097_1;
buffer_wire buffer_11097_1 (.in(n11097_0), .out(n11097_1));
wire n11098; //CHANX 4 (4,5) #40
wire n11098_0;
wire n11098_1;
buffer_wire buffer_11098_1 (.in(n11098_0), .out(n11098_1));
wire n11099; //CHANX 4 (4,5) #41
wire n11099_0;
wire n11099_1;
buffer_wire buffer_11099_1 (.in(n11099_0), .out(n11099_1));
wire n11100; //CHANX 4 (4,5) #48
wire n11100_0;
wire n11100_1;
buffer_wire buffer_11100_1 (.in(n11100_0), .out(n11100_1));
wire n11101; //CHANX 4 (4,5) #49
wire n11101_0;
wire n11101_1;
buffer_wire buffer_11101_1 (.in(n11101_0), .out(n11101_1));
wire n11102; //CHANX 4 (4,5) #56
wire n11102_0;
wire n11102_1;
buffer_wire buffer_11102_1 (.in(n11102_0), .out(n11102_1));
wire n11103; //CHANX 4 (4,5) #57
wire n11103_0;
wire n11103_1;
buffer_wire buffer_11103_1 (.in(n11103_0), .out(n11103_1));
wire n11104; //CHANX 4 (4,5) #64
wire n11104_0;
wire n11104_1;
buffer_wire buffer_11104_1 (.in(n11104_0), .out(n11104_1));
wire n11105; //CHANX 4 (4,5) #65
wire n11105_0;
wire n11105_1;
buffer_wire buffer_11105_1 (.in(n11105_0), .out(n11105_1));
wire n11106; //CHANX 4 (4,5) #72
wire n11106_0;
wire n11106_1;
buffer_wire buffer_11106_1 (.in(n11106_0), .out(n11106_1));
wire n11107; //CHANX 4 (4,5) #73
wire n11107_0;
wire n11107_1;
buffer_wire buffer_11107_1 (.in(n11107_0), .out(n11107_1));
wire n11108; //CHANX 6 (4,5) #80
wire n11108_0;
wire n11108_1;
buffer_wire buffer_11108_1 (.in(n11108_0), .out(n11108_1));
wire n11109; //CHANX 6 (4,5) #81
wire n11109_0;
wire n11109_1;
buffer_wire buffer_11109_1 (.in(n11109_0), .out(n11109_1));
wire n11110; //CHANX 4 (5,5) #2
wire n11110_0;
wire n11110_1;
buffer_wire buffer_11110_1 (.in(n11110_0), .out(n11110_1));
wire n11111; //CHANX 4 (5,5) #3
wire n11111_0;
wire n11111_1;
buffer_wire buffer_11111_1 (.in(n11111_0), .out(n11111_1));
wire n11112; //CHANX 4 (5,5) #10
wire n11112_0;
wire n11112_1;
buffer_wire buffer_11112_1 (.in(n11112_0), .out(n11112_1));
wire n11113; //CHANX 4 (5,5) #11
wire n11113_0;
wire n11113_1;
buffer_wire buffer_11113_1 (.in(n11113_0), .out(n11113_1));
wire n11114; //CHANX 4 (5,5) #18
wire n11114_0;
wire n11114_1;
buffer_wire buffer_11114_1 (.in(n11114_0), .out(n11114_1));
wire n11115; //CHANX 4 (5,5) #19
wire n11115_0;
wire n11115_1;
buffer_wire buffer_11115_1 (.in(n11115_0), .out(n11115_1));
wire n11116; //CHANX 4 (5,5) #26
wire n11116_0;
wire n11116_1;
buffer_wire buffer_11116_1 (.in(n11116_0), .out(n11116_1));
wire n11117; //CHANX 4 (5,5) #27
wire n11117_0;
wire n11117_1;
buffer_wire buffer_11117_1 (.in(n11117_0), .out(n11117_1));
wire n11118; //CHANX 4 (5,5) #34
wire n11118_0;
wire n11118_1;
buffer_wire buffer_11118_1 (.in(n11118_0), .out(n11118_1));
wire n11119; //CHANX 4 (5,5) #35
wire n11119_0;
wire n11119_1;
buffer_wire buffer_11119_1 (.in(n11119_0), .out(n11119_1));
wire n11120; //CHANX 4 (5,5) #42
wire n11120_0;
wire n11120_1;
buffer_wire buffer_11120_1 (.in(n11120_0), .out(n11120_1));
wire n11121; //CHANX 4 (5,5) #43
wire n11121_0;
wire n11121_1;
buffer_wire buffer_11121_1 (.in(n11121_0), .out(n11121_1));
wire n11122; //CHANX 4 (5,5) #50
wire n11122_0;
wire n11122_1;
buffer_wire buffer_11122_1 (.in(n11122_0), .out(n11122_1));
wire n11123; //CHANX 4 (5,5) #51
wire n11123_0;
wire n11123_1;
buffer_wire buffer_11123_1 (.in(n11123_0), .out(n11123_1));
wire n11124; //CHANX 4 (5,5) #58
wire n11124_0;
wire n11124_1;
buffer_wire buffer_11124_1 (.in(n11124_0), .out(n11124_1));
wire n11125; //CHANX 4 (5,5) #59
wire n11125_0;
wire n11125_1;
buffer_wire buffer_11125_1 (.in(n11125_0), .out(n11125_1));
wire n11126; //CHANX 4 (5,5) #66
wire n11126_0;
wire n11126_1;
buffer_wire buffer_11126_1 (.in(n11126_0), .out(n11126_1));
wire n11127; //CHANX 4 (5,5) #67
wire n11127_0;
wire n11127_1;
buffer_wire buffer_11127_1 (.in(n11127_0), .out(n11127_1));
wire n11128; //CHANX 4 (5,5) #74
wire n11128_0;
wire n11128_1;
buffer_wire buffer_11128_1 (.in(n11128_0), .out(n11128_1));
wire n11129; //CHANX 4 (5,5) #75
wire n11129_0;
wire n11129_1;
buffer_wire buffer_11129_1 (.in(n11129_0), .out(n11129_1));
wire n11130; //CHANX 5 (5,5) #82
wire n11130_0;
wire n11130_1;
buffer_wire buffer_11130_1 (.in(n11130_0), .out(n11130_1));
wire n11131; //CHANX 5 (5,5) #83
wire n11131_0;
wire n11131_1;
buffer_wire buffer_11131_1 (.in(n11131_0), .out(n11131_1));
wire n11132; //CHANX 4 (6,5) #4
wire n11132_0;
wire n11132_1;
buffer_wire buffer_11132_1 (.in(n11132_0), .out(n11132_1));
wire n11133; //CHANX 4 (6,5) #5
wire n11133_0;
wire n11133_1;
buffer_wire buffer_11133_1 (.in(n11133_0), .out(n11133_1));
wire n11134; //CHANX 4 (6,5) #12
wire n11134_0;
wire n11134_1;
buffer_wire buffer_11134_1 (.in(n11134_0), .out(n11134_1));
wire n11135; //CHANX 4 (6,5) #13
wire n11135_0;
wire n11135_1;
buffer_wire buffer_11135_1 (.in(n11135_0), .out(n11135_1));
wire n11136; //CHANX 4 (6,5) #20
wire n11136_0;
wire n11136_1;
buffer_wire buffer_11136_1 (.in(n11136_0), .out(n11136_1));
wire n11137; //CHANX 4 (6,5) #21
wire n11137_0;
wire n11137_1;
buffer_wire buffer_11137_1 (.in(n11137_0), .out(n11137_1));
wire n11138; //CHANX 4 (6,5) #28
wire n11138_0;
wire n11138_1;
buffer_wire buffer_11138_1 (.in(n11138_0), .out(n11138_1));
wire n11139; //CHANX 4 (6,5) #29
wire n11139_0;
wire n11139_1;
buffer_wire buffer_11139_1 (.in(n11139_0), .out(n11139_1));
wire n11140; //CHANX 4 (6,5) #36
wire n11140_0;
wire n11140_1;
buffer_wire buffer_11140_1 (.in(n11140_0), .out(n11140_1));
wire n11141; //CHANX 4 (6,5) #37
wire n11141_0;
wire n11141_1;
buffer_wire buffer_11141_1 (.in(n11141_0), .out(n11141_1));
wire n11142; //CHANX 4 (6,5) #44
wire n11142_0;
wire n11142_1;
buffer_wire buffer_11142_1 (.in(n11142_0), .out(n11142_1));
wire n11143; //CHANX 4 (6,5) #45
wire n11143_0;
wire n11143_1;
buffer_wire buffer_11143_1 (.in(n11143_0), .out(n11143_1));
wire n11144; //CHANX 4 (6,5) #52
wire n11144_0;
wire n11144_1;
buffer_wire buffer_11144_1 (.in(n11144_0), .out(n11144_1));
wire n11145; //CHANX 4 (6,5) #53
wire n11145_0;
wire n11145_1;
buffer_wire buffer_11145_1 (.in(n11145_0), .out(n11145_1));
wire n11146; //CHANX 4 (6,5) #60
wire n11146_0;
wire n11146_1;
buffer_wire buffer_11146_1 (.in(n11146_0), .out(n11146_1));
wire n11147; //CHANX 4 (6,5) #61
wire n11147_0;
wire n11147_1;
buffer_wire buffer_11147_1 (.in(n11147_0), .out(n11147_1));
wire n11148; //CHANX 4 (6,5) #68
wire n11148_0;
wire n11148_1;
buffer_wire buffer_11148_1 (.in(n11148_0), .out(n11148_1));
wire n11149; //CHANX 4 (6,5) #69
wire n11149_0;
wire n11149_1;
buffer_wire buffer_11149_1 (.in(n11149_0), .out(n11149_1));
wire n11150; //CHANX 4 (6,5) #76
wire n11150_0;
wire n11150_1;
buffer_wire buffer_11150_1 (.in(n11150_0), .out(n11150_1));
wire n11151; //CHANX 4 (6,5) #77
wire n11151_0;
wire n11151_1;
buffer_wire buffer_11151_1 (.in(n11151_0), .out(n11151_1));
wire n11152; //CHANX 4 (6,5) #84
wire n11152_0;
wire n11152_1;
buffer_wire buffer_11152_1 (.in(n11152_0), .out(n11152_1));
wire n11153; //CHANX 4 (6,5) #85
wire n11153_0;
wire n11153_1;
buffer_wire buffer_11153_1 (.in(n11153_0), .out(n11153_1));
wire n11154; //CHANX 3 (7,5) #6
wire n11154_0;
wire n11155; //CHANX 3 (7,5) #7
wire n11155_0;
wire n11156; //CHANX 3 (7,5) #14
wire n11156_0;
wire n11157; //CHANX 3 (7,5) #15
wire n11157_0;
wire n11158; //CHANX 3 (7,5) #22
wire n11158_0;
wire n11159; //CHANX 3 (7,5) #23
wire n11159_0;
wire n11160; //CHANX 3 (7,5) #30
wire n11160_0;
wire n11161; //CHANX 3 (7,5) #31
wire n11161_0;
wire n11162; //CHANX 3 (7,5) #38
wire n11162_0;
wire n11163; //CHANX 3 (7,5) #39
wire n11163_0;
wire n11164; //CHANX 3 (7,5) #46
wire n11164_0;
wire n11165; //CHANX 3 (7,5) #47
wire n11165_0;
wire n11166; //CHANX 3 (7,5) #54
wire n11166_0;
wire n11167; //CHANX 3 (7,5) #55
wire n11167_0;
wire n11168; //CHANX 3 (7,5) #62
wire n11168_0;
wire n11169; //CHANX 3 (7,5) #63
wire n11169_0;
wire n11170; //CHANX 3 (7,5) #70
wire n11170_0;
wire n11171; //CHANX 3 (7,5) #71
wire n11171_0;
wire n11172; //CHANX 3 (7,5) #78
wire n11172_0;
wire n11173; //CHANX 3 (7,5) #79
wire n11173_0;
wire n11174; //CHANX 3 (7,5) #86
wire n11174_0;
wire n11175; //CHANX 3 (7,5) #87
wire n11175_0;
wire n11176; //CHANX 2 (8,5) #0
wire n11176_0;
wire n11177; //CHANX 2 (8,5) #1
wire n11177_0;
wire n11178; //CHANX 2 (8,5) #8
wire n11178_0;
wire n11179; //CHANX 2 (8,5) #9
wire n11179_0;
wire n11180; //CHANX 2 (8,5) #16
wire n11180_0;
wire n11181; //CHANX 2 (8,5) #17
wire n11181_0;
wire n11182; //CHANX 2 (8,5) #24
wire n11182_0;
wire n11183; //CHANX 2 (8,5) #25
wire n11183_0;
wire n11184; //CHANX 2 (8,5) #32
wire n11184_0;
wire n11185; //CHANX 2 (8,5) #33
wire n11185_0;
wire n11186; //CHANX 2 (8,5) #40
wire n11186_0;
wire n11187; //CHANX 2 (8,5) #41
wire n11187_0;
wire n11188; //CHANX 2 (8,5) #48
wire n11188_0;
wire n11189; //CHANX 2 (8,5) #49
wire n11189_0;
wire n11190; //CHANX 2 (8,5) #56
wire n11190_0;
wire n11191; //CHANX 2 (8,5) #57
wire n11191_0;
wire n11192; //CHANX 2 (8,5) #64
wire n11192_0;
wire n11193; //CHANX 2 (8,5) #65
wire n11193_0;
wire n11194; //CHANX 2 (8,5) #72
wire n11194_0;
wire n11195; //CHANX 2 (8,5) #73
wire n11195_0;
wire n11196; //CHANX 2 (8,5) #88
wire n11196_0;
wire n11197; //CHANX 2 (8,5) #89
wire n11197_0;
wire n11198; //CHANX 1 (9,5) #2
wire n11198_0;
wire n11199; //CHANX 1 (9,5) #3
wire n11199_0;
wire n11200; //CHANX 1 (9,5) #10
wire n11200_0;
wire n11201; //CHANX 1 (9,5) #11
wire n11201_0;
wire n11202; //CHANX 1 (9,5) #18
wire n11202_0;
wire n11203; //CHANX 1 (9,5) #19
wire n11203_0;
wire n11204; //CHANX 1 (9,5) #26
wire n11204_0;
wire n11205; //CHANX 1 (9,5) #27
wire n11205_0;
wire n11206; //CHANX 1 (9,5) #34
wire n11206_0;
wire n11207; //CHANX 1 (9,5) #35
wire n11207_0;
wire n11208; //CHANX 1 (9,5) #42
wire n11208_0;
wire n11209; //CHANX 1 (9,5) #43
wire n11209_0;
wire n11210; //CHANX 1 (9,5) #50
wire n11210_0;
wire n11211; //CHANX 1 (9,5) #51
wire n11211_0;
wire n11212; //CHANX 1 (9,5) #58
wire n11212_0;
wire n11213; //CHANX 1 (9,5) #59
wire n11213_0;
wire n11214; //CHANX 1 (9,5) #66
wire n11214_0;
wire n11215; //CHANX 1 (9,5) #67
wire n11215_0;
wire n11216; //CHANX 1 (9,5) #74
wire n11216_0;
wire n11217; //CHANX 1 (9,5) #75
wire n11217_0;
wire n11218; //CHANX 1 (9,5) #90
wire n11218_0;
wire n11219; //CHANX 1 (9,5) #91
wire n11219_0;
wire n11220; //CHANX 2 (1,6) #0
wire n11220_0;
wire n11221; //CHANX 2 (1,6) #1
wire n11221_0;
wire n11222; //CHANX 3 (1,6) #2
wire n11222_0;
wire n11223; //CHANX 3 (1,6) #3
wire n11223_0;
wire n11224; //CHANX 4 (1,6) #4
wire n11224_0;
wire n11224_1;
buffer_wire buffer_11224_1 (.in(n11224_0), .out(n11224_1));
wire n11225; //CHANX 4 (1,6) #5
wire n11225_0;
wire n11225_1;
buffer_wire buffer_11225_1 (.in(n11225_0), .out(n11225_1));
wire n11226; //CHANX 1 (1,6) #6
wire n11226_0;
wire n11227; //CHANX 1 (1,6) #7
wire n11227_0;
wire n11228; //CHANX 2 (1,6) #8
wire n11228_0;
wire n11229; //CHANX 2 (1,6) #9
wire n11229_0;
wire n11230; //CHANX 3 (1,6) #10
wire n11230_0;
wire n11231; //CHANX 3 (1,6) #11
wire n11231_0;
wire n11232; //CHANX 4 (1,6) #12
wire n11232_0;
wire n11232_1;
buffer_wire buffer_11232_1 (.in(n11232_0), .out(n11232_1));
wire n11233; //CHANX 4 (1,6) #13
wire n11233_0;
wire n11233_1;
buffer_wire buffer_11233_1 (.in(n11233_0), .out(n11233_1));
wire n11234; //CHANX 1 (1,6) #14
wire n11234_0;
wire n11235; //CHANX 1 (1,6) #15
wire n11235_0;
wire n11236; //CHANX 2 (1,6) #16
wire n11236_0;
wire n11237; //CHANX 2 (1,6) #17
wire n11237_0;
wire n11238; //CHANX 3 (1,6) #18
wire n11238_0;
wire n11239; //CHANX 3 (1,6) #19
wire n11239_0;
wire n11240; //CHANX 4 (1,6) #20
wire n11240_0;
wire n11240_1;
buffer_wire buffer_11240_1 (.in(n11240_0), .out(n11240_1));
wire n11241; //CHANX 4 (1,6) #21
wire n11241_0;
wire n11241_1;
buffer_wire buffer_11241_1 (.in(n11241_0), .out(n11241_1));
wire n11242; //CHANX 1 (1,6) #22
wire n11242_0;
wire n11243; //CHANX 1 (1,6) #23
wire n11243_0;
wire n11244; //CHANX 2 (1,6) #24
wire n11244_0;
wire n11245; //CHANX 2 (1,6) #25
wire n11245_0;
wire n11246; //CHANX 3 (1,6) #26
wire n11246_0;
wire n11247; //CHANX 3 (1,6) #27
wire n11247_0;
wire n11248; //CHANX 4 (1,6) #28
wire n11248_0;
wire n11248_1;
buffer_wire buffer_11248_1 (.in(n11248_0), .out(n11248_1));
wire n11249; //CHANX 4 (1,6) #29
wire n11249_0;
wire n11249_1;
buffer_wire buffer_11249_1 (.in(n11249_0), .out(n11249_1));
wire n11250; //CHANX 1 (1,6) #30
wire n11250_0;
wire n11251; //CHANX 1 (1,6) #31
wire n11251_0;
wire n11252; //CHANX 2 (1,6) #32
wire n11252_0;
wire n11253; //CHANX 2 (1,6) #33
wire n11253_0;
wire n11254; //CHANX 3 (1,6) #34
wire n11254_0;
wire n11255; //CHANX 3 (1,6) #35
wire n11255_0;
wire n11256; //CHANX 4 (1,6) #36
wire n11256_0;
wire n11256_1;
buffer_wire buffer_11256_1 (.in(n11256_0), .out(n11256_1));
wire n11257; //CHANX 4 (1,6) #37
wire n11257_0;
wire n11257_1;
buffer_wire buffer_11257_1 (.in(n11257_0), .out(n11257_1));
wire n11258; //CHANX 1 (1,6) #38
wire n11258_0;
wire n11259; //CHANX 1 (1,6) #39
wire n11259_0;
wire n11260; //CHANX 2 (1,6) #40
wire n11260_0;
wire n11261; //CHANX 2 (1,6) #41
wire n11261_0;
wire n11262; //CHANX 3 (1,6) #42
wire n11262_0;
wire n11263; //CHANX 3 (1,6) #43
wire n11263_0;
wire n11264; //CHANX 4 (1,6) #44
wire n11264_0;
wire n11264_1;
buffer_wire buffer_11264_1 (.in(n11264_0), .out(n11264_1));
wire n11265; //CHANX 4 (1,6) #45
wire n11265_0;
wire n11265_1;
buffer_wire buffer_11265_1 (.in(n11265_0), .out(n11265_1));
wire n11266; //CHANX 1 (1,6) #46
wire n11266_0;
wire n11267; //CHANX 1 (1,6) #47
wire n11267_0;
wire n11268; //CHANX 2 (1,6) #48
wire n11268_0;
wire n11269; //CHANX 2 (1,6) #49
wire n11269_0;
wire n11270; //CHANX 3 (1,6) #50
wire n11270_0;
wire n11271; //CHANX 3 (1,6) #51
wire n11271_0;
wire n11272; //CHANX 4 (1,6) #52
wire n11272_0;
wire n11272_1;
buffer_wire buffer_11272_1 (.in(n11272_0), .out(n11272_1));
wire n11273; //CHANX 4 (1,6) #53
wire n11273_0;
wire n11273_1;
buffer_wire buffer_11273_1 (.in(n11273_0), .out(n11273_1));
wire n11274; //CHANX 1 (1,6) #54
wire n11274_0;
wire n11275; //CHANX 1 (1,6) #55
wire n11275_0;
wire n11276; //CHANX 2 (1,6) #56
wire n11276_0;
wire n11277; //CHANX 2 (1,6) #57
wire n11277_0;
wire n11278; //CHANX 3 (1,6) #58
wire n11278_0;
wire n11279; //CHANX 3 (1,6) #59
wire n11279_0;
wire n11280; //CHANX 4 (1,6) #60
wire n11280_0;
wire n11280_1;
buffer_wire buffer_11280_1 (.in(n11280_0), .out(n11280_1));
wire n11281; //CHANX 4 (1,6) #61
wire n11281_0;
wire n11281_1;
buffer_wire buffer_11281_1 (.in(n11281_0), .out(n11281_1));
wire n11282; //CHANX 1 (1,6) #62
wire n11282_0;
wire n11283; //CHANX 1 (1,6) #63
wire n11283_0;
wire n11284; //CHANX 2 (1,6) #64
wire n11284_0;
wire n11285; //CHANX 2 (1,6) #65
wire n11285_0;
wire n11286; //CHANX 3 (1,6) #66
wire n11286_0;
wire n11287; //CHANX 3 (1,6) #67
wire n11287_0;
wire n11288; //CHANX 4 (1,6) #68
wire n11288_0;
wire n11288_1;
buffer_wire buffer_11288_1 (.in(n11288_0), .out(n11288_1));
wire n11289; //CHANX 4 (1,6) #69
wire n11289_0;
wire n11289_1;
buffer_wire buffer_11289_1 (.in(n11289_0), .out(n11289_1));
wire n11290; //CHANX 1 (1,6) #70
wire n11290_0;
wire n11291; //CHANX 1 (1,6) #71
wire n11291_0;
wire n11292; //CHANX 2 (1,6) #72
wire n11292_0;
wire n11293; //CHANX 2 (1,6) #73
wire n11293_0;
wire n11294; //CHANX 3 (1,6) #74
wire n11294_0;
wire n11295; //CHANX 3 (1,6) #75
wire n11295_0;
wire n11296; //CHANX 4 (1,6) #76
wire n11296_0;
wire n11296_1;
buffer_wire buffer_11296_1 (.in(n11296_0), .out(n11296_1));
wire n11297; //CHANX 4 (1,6) #77
wire n11297_0;
wire n11297_1;
buffer_wire buffer_11297_1 (.in(n11297_0), .out(n11297_1));
wire n11298; //CHANX 1 (1,6) #78
wire n11298_0;
wire n11299; //CHANX 1 (1,6) #79
wire n11299_0;
wire n11300; //CHANX 2 (1,6) #80
wire n11300_0;
wire n11301; //CHANX 2 (1,6) #81
wire n11301_0;
wire n11302; //CHANX 3 (1,6) #82
wire n11302_0;
wire n11303; //CHANX 3 (1,6) #83
wire n11303_0;
wire n11304; //CHANX 4 (1,6) #84
wire n11304_0;
wire n11304_1;
buffer_wire buffer_11304_1 (.in(n11304_0), .out(n11304_1));
wire n11305; //CHANX 4 (1,6) #85
wire n11305_0;
wire n11305_1;
buffer_wire buffer_11305_1 (.in(n11305_0), .out(n11305_1));
wire n11306; //CHANX 5 (1,6) #86
wire n11306_0;
wire n11306_1;
buffer_wire buffer_11306_1 (.in(n11306_0), .out(n11306_1));
wire n11307; //CHANX 5 (1,6) #87
wire n11307_0;
wire n11307_1;
buffer_wire buffer_11307_1 (.in(n11307_0), .out(n11307_1));
wire n11308; //CHANX 6 (1,6) #88
wire n11308_0;
wire n11308_1;
buffer_wire buffer_11308_1 (.in(n11308_0), .out(n11308_1));
wire n11309; //CHANX 6 (1,6) #89
wire n11309_0;
wire n11309_1;
buffer_wire buffer_11309_1 (.in(n11309_0), .out(n11309_1));
wire n11310; //CHANX 7 (1,6) #90
wire n11310_0;
wire n11310_1;
wire n11310_2;
buffer_wire buffer_11310_2 (.in(n11310_1), .out(n11310_2));
buffer_wire buffer_11310_1 (.in(n11310_0), .out(n11310_1));
wire n11311; //CHANX 7 (1,6) #91
wire n11311_0;
wire n11311_1;
wire n11311_2;
buffer_wire buffer_11311_2 (.in(n11311_1), .out(n11311_2));
buffer_wire buffer_11311_1 (.in(n11311_0), .out(n11311_1));
wire n11312; //CHANX 4 (2,6) #6
wire n11312_0;
wire n11312_1;
buffer_wire buffer_11312_1 (.in(n11312_0), .out(n11312_1));
wire n11313; //CHANX 4 (2,6) #7
wire n11313_0;
wire n11313_1;
buffer_wire buffer_11313_1 (.in(n11313_0), .out(n11313_1));
wire n11314; //CHANX 4 (2,6) #14
wire n11314_0;
wire n11314_1;
buffer_wire buffer_11314_1 (.in(n11314_0), .out(n11314_1));
wire n11315; //CHANX 4 (2,6) #15
wire n11315_0;
wire n11315_1;
buffer_wire buffer_11315_1 (.in(n11315_0), .out(n11315_1));
wire n11316; //CHANX 4 (2,6) #22
wire n11316_0;
wire n11316_1;
buffer_wire buffer_11316_1 (.in(n11316_0), .out(n11316_1));
wire n11317; //CHANX 4 (2,6) #23
wire n11317_0;
wire n11317_1;
buffer_wire buffer_11317_1 (.in(n11317_0), .out(n11317_1));
wire n11318; //CHANX 4 (2,6) #30
wire n11318_0;
wire n11318_1;
buffer_wire buffer_11318_1 (.in(n11318_0), .out(n11318_1));
wire n11319; //CHANX 4 (2,6) #31
wire n11319_0;
wire n11319_1;
buffer_wire buffer_11319_1 (.in(n11319_0), .out(n11319_1));
wire n11320; //CHANX 4 (2,6) #38
wire n11320_0;
wire n11320_1;
buffer_wire buffer_11320_1 (.in(n11320_0), .out(n11320_1));
wire n11321; //CHANX 4 (2,6) #39
wire n11321_0;
wire n11321_1;
buffer_wire buffer_11321_1 (.in(n11321_0), .out(n11321_1));
wire n11322; //CHANX 4 (2,6) #46
wire n11322_0;
wire n11322_1;
buffer_wire buffer_11322_1 (.in(n11322_0), .out(n11322_1));
wire n11323; //CHANX 4 (2,6) #47
wire n11323_0;
wire n11323_1;
buffer_wire buffer_11323_1 (.in(n11323_0), .out(n11323_1));
wire n11324; //CHANX 4 (2,6) #54
wire n11324_0;
wire n11324_1;
buffer_wire buffer_11324_1 (.in(n11324_0), .out(n11324_1));
wire n11325; //CHANX 4 (2,6) #55
wire n11325_0;
wire n11325_1;
buffer_wire buffer_11325_1 (.in(n11325_0), .out(n11325_1));
wire n11326; //CHANX 4 (2,6) #62
wire n11326_0;
wire n11326_1;
buffer_wire buffer_11326_1 (.in(n11326_0), .out(n11326_1));
wire n11327; //CHANX 4 (2,6) #63
wire n11327_0;
wire n11327_1;
buffer_wire buffer_11327_1 (.in(n11327_0), .out(n11327_1));
wire n11328; //CHANX 4 (2,6) #70
wire n11328_0;
wire n11328_1;
buffer_wire buffer_11328_1 (.in(n11328_0), .out(n11328_1));
wire n11329; //CHANX 4 (2,6) #71
wire n11329_0;
wire n11329_1;
buffer_wire buffer_11329_1 (.in(n11329_0), .out(n11329_1));
wire n11330; //CHANX 4 (2,6) #78
wire n11330_0;
wire n11330_1;
buffer_wire buffer_11330_1 (.in(n11330_0), .out(n11330_1));
wire n11331; //CHANX 4 (2,6) #79
wire n11331_0;
wire n11331_1;
buffer_wire buffer_11331_1 (.in(n11331_0), .out(n11331_1));
wire n11332; //CHANX 4 (3,6) #0
wire n11332_0;
wire n11332_1;
buffer_wire buffer_11332_1 (.in(n11332_0), .out(n11332_1));
wire n11333; //CHANX 4 (3,6) #1
wire n11333_0;
wire n11333_1;
buffer_wire buffer_11333_1 (.in(n11333_0), .out(n11333_1));
wire n11334; //CHANX 4 (3,6) #8
wire n11334_0;
wire n11334_1;
buffer_wire buffer_11334_1 (.in(n11334_0), .out(n11334_1));
wire n11335; //CHANX 4 (3,6) #9
wire n11335_0;
wire n11335_1;
buffer_wire buffer_11335_1 (.in(n11335_0), .out(n11335_1));
wire n11336; //CHANX 4 (3,6) #16
wire n11336_0;
wire n11336_1;
buffer_wire buffer_11336_1 (.in(n11336_0), .out(n11336_1));
wire n11337; //CHANX 4 (3,6) #17
wire n11337_0;
wire n11337_1;
buffer_wire buffer_11337_1 (.in(n11337_0), .out(n11337_1));
wire n11338; //CHANX 4 (3,6) #24
wire n11338_0;
wire n11338_1;
buffer_wire buffer_11338_1 (.in(n11338_0), .out(n11338_1));
wire n11339; //CHANX 4 (3,6) #25
wire n11339_0;
wire n11339_1;
buffer_wire buffer_11339_1 (.in(n11339_0), .out(n11339_1));
wire n11340; //CHANX 4 (3,6) #32
wire n11340_0;
wire n11340_1;
buffer_wire buffer_11340_1 (.in(n11340_0), .out(n11340_1));
wire n11341; //CHANX 4 (3,6) #33
wire n11341_0;
wire n11341_1;
buffer_wire buffer_11341_1 (.in(n11341_0), .out(n11341_1));
wire n11342; //CHANX 4 (3,6) #40
wire n11342_0;
wire n11342_1;
buffer_wire buffer_11342_1 (.in(n11342_0), .out(n11342_1));
wire n11343; //CHANX 4 (3,6) #41
wire n11343_0;
wire n11343_1;
buffer_wire buffer_11343_1 (.in(n11343_0), .out(n11343_1));
wire n11344; //CHANX 4 (3,6) #48
wire n11344_0;
wire n11344_1;
buffer_wire buffer_11344_1 (.in(n11344_0), .out(n11344_1));
wire n11345; //CHANX 4 (3,6) #49
wire n11345_0;
wire n11345_1;
buffer_wire buffer_11345_1 (.in(n11345_0), .out(n11345_1));
wire n11346; //CHANX 4 (3,6) #56
wire n11346_0;
wire n11346_1;
buffer_wire buffer_11346_1 (.in(n11346_0), .out(n11346_1));
wire n11347; //CHANX 4 (3,6) #57
wire n11347_0;
wire n11347_1;
buffer_wire buffer_11347_1 (.in(n11347_0), .out(n11347_1));
wire n11348; //CHANX 4 (3,6) #64
wire n11348_0;
wire n11348_1;
buffer_wire buffer_11348_1 (.in(n11348_0), .out(n11348_1));
wire n11349; //CHANX 4 (3,6) #65
wire n11349_0;
wire n11349_1;
buffer_wire buffer_11349_1 (.in(n11349_0), .out(n11349_1));
wire n11350; //CHANX 4 (3,6) #72
wire n11350_0;
wire n11350_1;
buffer_wire buffer_11350_1 (.in(n11350_0), .out(n11350_1));
wire n11351; //CHANX 4 (3,6) #73
wire n11351_0;
wire n11351_1;
buffer_wire buffer_11351_1 (.in(n11351_0), .out(n11351_1));
wire n11352; //CHANX 7 (3,6) #80
wire n11352_0;
wire n11352_1;
wire n11352_2;
buffer_wire buffer_11352_2 (.in(n11352_1), .out(n11352_2));
buffer_wire buffer_11352_1 (.in(n11352_0), .out(n11352_1));
wire n11353; //CHANX 7 (3,6) #81
wire n11353_0;
wire n11353_1;
wire n11353_2;
buffer_wire buffer_11353_2 (.in(n11353_1), .out(n11353_2));
buffer_wire buffer_11353_1 (.in(n11353_0), .out(n11353_1));
wire n11354; //CHANX 4 (4,6) #2
wire n11354_0;
wire n11354_1;
buffer_wire buffer_11354_1 (.in(n11354_0), .out(n11354_1));
wire n11355; //CHANX 4 (4,6) #3
wire n11355_0;
wire n11355_1;
buffer_wire buffer_11355_1 (.in(n11355_0), .out(n11355_1));
wire n11356; //CHANX 4 (4,6) #10
wire n11356_0;
wire n11356_1;
buffer_wire buffer_11356_1 (.in(n11356_0), .out(n11356_1));
wire n11357; //CHANX 4 (4,6) #11
wire n11357_0;
wire n11357_1;
buffer_wire buffer_11357_1 (.in(n11357_0), .out(n11357_1));
wire n11358; //CHANX 4 (4,6) #18
wire n11358_0;
wire n11358_1;
buffer_wire buffer_11358_1 (.in(n11358_0), .out(n11358_1));
wire n11359; //CHANX 4 (4,6) #19
wire n11359_0;
wire n11359_1;
buffer_wire buffer_11359_1 (.in(n11359_0), .out(n11359_1));
wire n11360; //CHANX 4 (4,6) #26
wire n11360_0;
wire n11360_1;
buffer_wire buffer_11360_1 (.in(n11360_0), .out(n11360_1));
wire n11361; //CHANX 4 (4,6) #27
wire n11361_0;
wire n11361_1;
buffer_wire buffer_11361_1 (.in(n11361_0), .out(n11361_1));
wire n11362; //CHANX 4 (4,6) #34
wire n11362_0;
wire n11362_1;
buffer_wire buffer_11362_1 (.in(n11362_0), .out(n11362_1));
wire n11363; //CHANX 4 (4,6) #35
wire n11363_0;
wire n11363_1;
buffer_wire buffer_11363_1 (.in(n11363_0), .out(n11363_1));
wire n11364; //CHANX 4 (4,6) #42
wire n11364_0;
wire n11364_1;
buffer_wire buffer_11364_1 (.in(n11364_0), .out(n11364_1));
wire n11365; //CHANX 4 (4,6) #43
wire n11365_0;
wire n11365_1;
buffer_wire buffer_11365_1 (.in(n11365_0), .out(n11365_1));
wire n11366; //CHANX 4 (4,6) #50
wire n11366_0;
wire n11366_1;
buffer_wire buffer_11366_1 (.in(n11366_0), .out(n11366_1));
wire n11367; //CHANX 4 (4,6) #51
wire n11367_0;
wire n11367_1;
buffer_wire buffer_11367_1 (.in(n11367_0), .out(n11367_1));
wire n11368; //CHANX 4 (4,6) #58
wire n11368_0;
wire n11368_1;
buffer_wire buffer_11368_1 (.in(n11368_0), .out(n11368_1));
wire n11369; //CHANX 4 (4,6) #59
wire n11369_0;
wire n11369_1;
buffer_wire buffer_11369_1 (.in(n11369_0), .out(n11369_1));
wire n11370; //CHANX 4 (4,6) #66
wire n11370_0;
wire n11370_1;
buffer_wire buffer_11370_1 (.in(n11370_0), .out(n11370_1));
wire n11371; //CHANX 4 (4,6) #67
wire n11371_0;
wire n11371_1;
buffer_wire buffer_11371_1 (.in(n11371_0), .out(n11371_1));
wire n11372; //CHANX 4 (4,6) #74
wire n11372_0;
wire n11372_1;
buffer_wire buffer_11372_1 (.in(n11372_0), .out(n11372_1));
wire n11373; //CHANX 4 (4,6) #75
wire n11373_0;
wire n11373_1;
buffer_wire buffer_11373_1 (.in(n11373_0), .out(n11373_1));
wire n11374; //CHANX 6 (4,6) #82
wire n11374_0;
wire n11374_1;
buffer_wire buffer_11374_1 (.in(n11374_0), .out(n11374_1));
wire n11375; //CHANX 6 (4,6) #83
wire n11375_0;
wire n11375_1;
buffer_wire buffer_11375_1 (.in(n11375_0), .out(n11375_1));
wire n11376; //CHANX 4 (5,6) #4
wire n11376_0;
wire n11376_1;
buffer_wire buffer_11376_1 (.in(n11376_0), .out(n11376_1));
wire n11377; //CHANX 4 (5,6) #5
wire n11377_0;
wire n11377_1;
buffer_wire buffer_11377_1 (.in(n11377_0), .out(n11377_1));
wire n11378; //CHANX 4 (5,6) #12
wire n11378_0;
wire n11378_1;
buffer_wire buffer_11378_1 (.in(n11378_0), .out(n11378_1));
wire n11379; //CHANX 4 (5,6) #13
wire n11379_0;
wire n11379_1;
buffer_wire buffer_11379_1 (.in(n11379_0), .out(n11379_1));
wire n11380; //CHANX 4 (5,6) #20
wire n11380_0;
wire n11380_1;
buffer_wire buffer_11380_1 (.in(n11380_0), .out(n11380_1));
wire n11381; //CHANX 4 (5,6) #21
wire n11381_0;
wire n11381_1;
buffer_wire buffer_11381_1 (.in(n11381_0), .out(n11381_1));
wire n11382; //CHANX 4 (5,6) #28
wire n11382_0;
wire n11382_1;
buffer_wire buffer_11382_1 (.in(n11382_0), .out(n11382_1));
wire n11383; //CHANX 4 (5,6) #29
wire n11383_0;
wire n11383_1;
buffer_wire buffer_11383_1 (.in(n11383_0), .out(n11383_1));
wire n11384; //CHANX 4 (5,6) #36
wire n11384_0;
wire n11384_1;
buffer_wire buffer_11384_1 (.in(n11384_0), .out(n11384_1));
wire n11385; //CHANX 4 (5,6) #37
wire n11385_0;
wire n11385_1;
buffer_wire buffer_11385_1 (.in(n11385_0), .out(n11385_1));
wire n11386; //CHANX 4 (5,6) #44
wire n11386_0;
wire n11386_1;
buffer_wire buffer_11386_1 (.in(n11386_0), .out(n11386_1));
wire n11387; //CHANX 4 (5,6) #45
wire n11387_0;
wire n11387_1;
buffer_wire buffer_11387_1 (.in(n11387_0), .out(n11387_1));
wire n11388; //CHANX 4 (5,6) #52
wire n11388_0;
wire n11388_1;
buffer_wire buffer_11388_1 (.in(n11388_0), .out(n11388_1));
wire n11389; //CHANX 4 (5,6) #53
wire n11389_0;
wire n11389_1;
buffer_wire buffer_11389_1 (.in(n11389_0), .out(n11389_1));
wire n11390; //CHANX 4 (5,6) #60
wire n11390_0;
wire n11390_1;
buffer_wire buffer_11390_1 (.in(n11390_0), .out(n11390_1));
wire n11391; //CHANX 4 (5,6) #61
wire n11391_0;
wire n11391_1;
buffer_wire buffer_11391_1 (.in(n11391_0), .out(n11391_1));
wire n11392; //CHANX 4 (5,6) #68
wire n11392_0;
wire n11392_1;
buffer_wire buffer_11392_1 (.in(n11392_0), .out(n11392_1));
wire n11393; //CHANX 4 (5,6) #69
wire n11393_0;
wire n11393_1;
buffer_wire buffer_11393_1 (.in(n11393_0), .out(n11393_1));
wire n11394; //CHANX 4 (5,6) #76
wire n11394_0;
wire n11394_1;
buffer_wire buffer_11394_1 (.in(n11394_0), .out(n11394_1));
wire n11395; //CHANX 4 (5,6) #77
wire n11395_0;
wire n11395_1;
buffer_wire buffer_11395_1 (.in(n11395_0), .out(n11395_1));
wire n11396; //CHANX 5 (5,6) #84
wire n11396_0;
wire n11396_1;
buffer_wire buffer_11396_1 (.in(n11396_0), .out(n11396_1));
wire n11397; //CHANX 5 (5,6) #85
wire n11397_0;
wire n11397_1;
buffer_wire buffer_11397_1 (.in(n11397_0), .out(n11397_1));
wire n11398; //CHANX 4 (6,6) #6
wire n11398_0;
wire n11398_1;
buffer_wire buffer_11398_1 (.in(n11398_0), .out(n11398_1));
wire n11399; //CHANX 4 (6,6) #7
wire n11399_0;
wire n11399_1;
buffer_wire buffer_11399_1 (.in(n11399_0), .out(n11399_1));
wire n11400; //CHANX 4 (6,6) #14
wire n11400_0;
wire n11400_1;
buffer_wire buffer_11400_1 (.in(n11400_0), .out(n11400_1));
wire n11401; //CHANX 4 (6,6) #15
wire n11401_0;
wire n11401_1;
buffer_wire buffer_11401_1 (.in(n11401_0), .out(n11401_1));
wire n11402; //CHANX 4 (6,6) #22
wire n11402_0;
wire n11402_1;
buffer_wire buffer_11402_1 (.in(n11402_0), .out(n11402_1));
wire n11403; //CHANX 4 (6,6) #23
wire n11403_0;
wire n11403_1;
buffer_wire buffer_11403_1 (.in(n11403_0), .out(n11403_1));
wire n11404; //CHANX 4 (6,6) #30
wire n11404_0;
wire n11404_1;
buffer_wire buffer_11404_1 (.in(n11404_0), .out(n11404_1));
wire n11405; //CHANX 4 (6,6) #31
wire n11405_0;
wire n11405_1;
buffer_wire buffer_11405_1 (.in(n11405_0), .out(n11405_1));
wire n11406; //CHANX 4 (6,6) #38
wire n11406_0;
wire n11406_1;
buffer_wire buffer_11406_1 (.in(n11406_0), .out(n11406_1));
wire n11407; //CHANX 4 (6,6) #39
wire n11407_0;
wire n11407_1;
buffer_wire buffer_11407_1 (.in(n11407_0), .out(n11407_1));
wire n11408; //CHANX 4 (6,6) #46
wire n11408_0;
wire n11408_1;
buffer_wire buffer_11408_1 (.in(n11408_0), .out(n11408_1));
wire n11409; //CHANX 4 (6,6) #47
wire n11409_0;
wire n11409_1;
buffer_wire buffer_11409_1 (.in(n11409_0), .out(n11409_1));
wire n11410; //CHANX 4 (6,6) #54
wire n11410_0;
wire n11410_1;
buffer_wire buffer_11410_1 (.in(n11410_0), .out(n11410_1));
wire n11411; //CHANX 4 (6,6) #55
wire n11411_0;
wire n11411_1;
buffer_wire buffer_11411_1 (.in(n11411_0), .out(n11411_1));
wire n11412; //CHANX 4 (6,6) #62
wire n11412_0;
wire n11412_1;
buffer_wire buffer_11412_1 (.in(n11412_0), .out(n11412_1));
wire n11413; //CHANX 4 (6,6) #63
wire n11413_0;
wire n11413_1;
buffer_wire buffer_11413_1 (.in(n11413_0), .out(n11413_1));
wire n11414; //CHANX 4 (6,6) #70
wire n11414_0;
wire n11414_1;
buffer_wire buffer_11414_1 (.in(n11414_0), .out(n11414_1));
wire n11415; //CHANX 4 (6,6) #71
wire n11415_0;
wire n11415_1;
buffer_wire buffer_11415_1 (.in(n11415_0), .out(n11415_1));
wire n11416; //CHANX 4 (6,6) #78
wire n11416_0;
wire n11416_1;
buffer_wire buffer_11416_1 (.in(n11416_0), .out(n11416_1));
wire n11417; //CHANX 4 (6,6) #79
wire n11417_0;
wire n11417_1;
buffer_wire buffer_11417_1 (.in(n11417_0), .out(n11417_1));
wire n11418; //CHANX 4 (6,6) #86
wire n11418_0;
wire n11418_1;
buffer_wire buffer_11418_1 (.in(n11418_0), .out(n11418_1));
wire n11419; //CHANX 4 (6,6) #87
wire n11419_0;
wire n11419_1;
buffer_wire buffer_11419_1 (.in(n11419_0), .out(n11419_1));
wire n11420; //CHANX 3 (7,6) #0
wire n11420_0;
wire n11421; //CHANX 3 (7,6) #1
wire n11421_0;
wire n11422; //CHANX 3 (7,6) #8
wire n11422_0;
wire n11423; //CHANX 3 (7,6) #9
wire n11423_0;
wire n11424; //CHANX 3 (7,6) #16
wire n11424_0;
wire n11425; //CHANX 3 (7,6) #17
wire n11425_0;
wire n11426; //CHANX 3 (7,6) #24
wire n11426_0;
wire n11427; //CHANX 3 (7,6) #25
wire n11427_0;
wire n11428; //CHANX 3 (7,6) #32
wire n11428_0;
wire n11429; //CHANX 3 (7,6) #33
wire n11429_0;
wire n11430; //CHANX 3 (7,6) #40
wire n11430_0;
wire n11431; //CHANX 3 (7,6) #41
wire n11431_0;
wire n11432; //CHANX 3 (7,6) #48
wire n11432_0;
wire n11433; //CHANX 3 (7,6) #49
wire n11433_0;
wire n11434; //CHANX 3 (7,6) #56
wire n11434_0;
wire n11435; //CHANX 3 (7,6) #57
wire n11435_0;
wire n11436; //CHANX 3 (7,6) #64
wire n11436_0;
wire n11437; //CHANX 3 (7,6) #65
wire n11437_0;
wire n11438; //CHANX 3 (7,6) #72
wire n11438_0;
wire n11439; //CHANX 3 (7,6) #73
wire n11439_0;
wire n11440; //CHANX 3 (7,6) #88
wire n11440_0;
wire n11441; //CHANX 3 (7,6) #89
wire n11441_0;
wire n11442; //CHANX 2 (8,6) #2
wire n11442_0;
wire n11443; //CHANX 2 (8,6) #3
wire n11443_0;
wire n11444; //CHANX 2 (8,6) #10
wire n11444_0;
wire n11445; //CHANX 2 (8,6) #11
wire n11445_0;
wire n11446; //CHANX 2 (8,6) #18
wire n11446_0;
wire n11447; //CHANX 2 (8,6) #19
wire n11447_0;
wire n11448; //CHANX 2 (8,6) #26
wire n11448_0;
wire n11449; //CHANX 2 (8,6) #27
wire n11449_0;
wire n11450; //CHANX 2 (8,6) #34
wire n11450_0;
wire n11451; //CHANX 2 (8,6) #35
wire n11451_0;
wire n11452; //CHANX 2 (8,6) #42
wire n11452_0;
wire n11453; //CHANX 2 (8,6) #43
wire n11453_0;
wire n11454; //CHANX 2 (8,6) #50
wire n11454_0;
wire n11455; //CHANX 2 (8,6) #51
wire n11455_0;
wire n11456; //CHANX 2 (8,6) #58
wire n11456_0;
wire n11457; //CHANX 2 (8,6) #59
wire n11457_0;
wire n11458; //CHANX 2 (8,6) #66
wire n11458_0;
wire n11459; //CHANX 2 (8,6) #67
wire n11459_0;
wire n11460; //CHANX 2 (8,6) #74
wire n11460_0;
wire n11461; //CHANX 2 (8,6) #75
wire n11461_0;
wire n11462; //CHANX 2 (8,6) #90
wire n11462_0;
wire n11463; //CHANX 2 (8,6) #91
wire n11463_0;
wire n11464; //CHANX 1 (9,6) #4
wire n11464_0;
wire n11465; //CHANX 1 (9,6) #5
wire n11465_0;
wire n11466; //CHANX 1 (9,6) #12
wire n11466_0;
wire n11467; //CHANX 1 (9,6) #13
wire n11467_0;
wire n11468; //CHANX 1 (9,6) #20
wire n11468_0;
wire n11469; //CHANX 1 (9,6) #21
wire n11469_0;
wire n11470; //CHANX 1 (9,6) #28
wire n11470_0;
wire n11471; //CHANX 1 (9,6) #29
wire n11471_0;
wire n11472; //CHANX 1 (9,6) #36
wire n11472_0;
wire n11473; //CHANX 1 (9,6) #37
wire n11473_0;
wire n11474; //CHANX 1 (9,6) #44
wire n11474_0;
wire n11475; //CHANX 1 (9,6) #45
wire n11475_0;
wire n11476; //CHANX 1 (9,6) #52
wire n11476_0;
wire n11477; //CHANX 1 (9,6) #53
wire n11477_0;
wire n11478; //CHANX 1 (9,6) #60
wire n11478_0;
wire n11479; //CHANX 1 (9,6) #61
wire n11479_0;
wire n11480; //CHANX 1 (9,6) #68
wire n11480_0;
wire n11481; //CHANX 1 (9,6) #69
wire n11481_0;
wire n11482; //CHANX 1 (9,6) #76
wire n11482_0;
wire n11483; //CHANX 1 (9,6) #77
wire n11483_0;
wire n11484; //CHANX 1 (1,7) #0
wire n11484_0;
wire n11485; //CHANX 1 (1,7) #1
wire n11485_0;
wire n11486; //CHANX 2 (1,7) #2
wire n11486_0;
wire n11487; //CHANX 2 (1,7) #3
wire n11487_0;
wire n11488; //CHANX 3 (1,7) #4
wire n11488_0;
wire n11489; //CHANX 3 (1,7) #5
wire n11489_0;
wire n11490; //CHANX 4 (1,7) #6
wire n11490_0;
wire n11490_1;
buffer_wire buffer_11490_1 (.in(n11490_0), .out(n11490_1));
wire n11491; //CHANX 4 (1,7) #7
wire n11491_0;
wire n11491_1;
buffer_wire buffer_11491_1 (.in(n11491_0), .out(n11491_1));
wire n11492; //CHANX 1 (1,7) #8
wire n11492_0;
wire n11493; //CHANX 1 (1,7) #9
wire n11493_0;
wire n11494; //CHANX 2 (1,7) #10
wire n11494_0;
wire n11495; //CHANX 2 (1,7) #11
wire n11495_0;
wire n11496; //CHANX 3 (1,7) #12
wire n11496_0;
wire n11497; //CHANX 3 (1,7) #13
wire n11497_0;
wire n11498; //CHANX 4 (1,7) #14
wire n11498_0;
wire n11498_1;
buffer_wire buffer_11498_1 (.in(n11498_0), .out(n11498_1));
wire n11499; //CHANX 4 (1,7) #15
wire n11499_0;
wire n11499_1;
buffer_wire buffer_11499_1 (.in(n11499_0), .out(n11499_1));
wire n11500; //CHANX 1 (1,7) #16
wire n11500_0;
wire n11501; //CHANX 1 (1,7) #17
wire n11501_0;
wire n11502; //CHANX 2 (1,7) #18
wire n11502_0;
wire n11503; //CHANX 2 (1,7) #19
wire n11503_0;
wire n11504; //CHANX 3 (1,7) #20
wire n11504_0;
wire n11505; //CHANX 3 (1,7) #21
wire n11505_0;
wire n11506; //CHANX 4 (1,7) #22
wire n11506_0;
wire n11506_1;
buffer_wire buffer_11506_1 (.in(n11506_0), .out(n11506_1));
wire n11507; //CHANX 4 (1,7) #23
wire n11507_0;
wire n11507_1;
buffer_wire buffer_11507_1 (.in(n11507_0), .out(n11507_1));
wire n11508; //CHANX 1 (1,7) #24
wire n11508_0;
wire n11509; //CHANX 1 (1,7) #25
wire n11509_0;
wire n11510; //CHANX 2 (1,7) #26
wire n11510_0;
wire n11511; //CHANX 2 (1,7) #27
wire n11511_0;
wire n11512; //CHANX 3 (1,7) #28
wire n11512_0;
wire n11513; //CHANX 3 (1,7) #29
wire n11513_0;
wire n11514; //CHANX 4 (1,7) #30
wire n11514_0;
wire n11514_1;
buffer_wire buffer_11514_1 (.in(n11514_0), .out(n11514_1));
wire n11515; //CHANX 4 (1,7) #31
wire n11515_0;
wire n11515_1;
buffer_wire buffer_11515_1 (.in(n11515_0), .out(n11515_1));
wire n11516; //CHANX 1 (1,7) #32
wire n11516_0;
wire n11517; //CHANX 1 (1,7) #33
wire n11517_0;
wire n11518; //CHANX 2 (1,7) #34
wire n11518_0;
wire n11519; //CHANX 2 (1,7) #35
wire n11519_0;
wire n11520; //CHANX 3 (1,7) #36
wire n11520_0;
wire n11521; //CHANX 3 (1,7) #37
wire n11521_0;
wire n11522; //CHANX 4 (1,7) #38
wire n11522_0;
wire n11522_1;
buffer_wire buffer_11522_1 (.in(n11522_0), .out(n11522_1));
wire n11523; //CHANX 4 (1,7) #39
wire n11523_0;
wire n11523_1;
buffer_wire buffer_11523_1 (.in(n11523_0), .out(n11523_1));
wire n11524; //CHANX 1 (1,7) #40
wire n11524_0;
wire n11525; //CHANX 1 (1,7) #41
wire n11525_0;
wire n11526; //CHANX 2 (1,7) #42
wire n11526_0;
wire n11527; //CHANX 2 (1,7) #43
wire n11527_0;
wire n11528; //CHANX 3 (1,7) #44
wire n11528_0;
wire n11529; //CHANX 3 (1,7) #45
wire n11529_0;
wire n11530; //CHANX 4 (1,7) #46
wire n11530_0;
wire n11530_1;
buffer_wire buffer_11530_1 (.in(n11530_0), .out(n11530_1));
wire n11531; //CHANX 4 (1,7) #47
wire n11531_0;
wire n11531_1;
buffer_wire buffer_11531_1 (.in(n11531_0), .out(n11531_1));
wire n11532; //CHANX 1 (1,7) #48
wire n11532_0;
wire n11533; //CHANX 1 (1,7) #49
wire n11533_0;
wire n11534; //CHANX 2 (1,7) #50
wire n11534_0;
wire n11535; //CHANX 2 (1,7) #51
wire n11535_0;
wire n11536; //CHANX 3 (1,7) #52
wire n11536_0;
wire n11537; //CHANX 3 (1,7) #53
wire n11537_0;
wire n11538; //CHANX 4 (1,7) #54
wire n11538_0;
wire n11538_1;
buffer_wire buffer_11538_1 (.in(n11538_0), .out(n11538_1));
wire n11539; //CHANX 4 (1,7) #55
wire n11539_0;
wire n11539_1;
buffer_wire buffer_11539_1 (.in(n11539_0), .out(n11539_1));
wire n11540; //CHANX 1 (1,7) #56
wire n11540_0;
wire n11541; //CHANX 1 (1,7) #57
wire n11541_0;
wire n11542; //CHANX 2 (1,7) #58
wire n11542_0;
wire n11543; //CHANX 2 (1,7) #59
wire n11543_0;
wire n11544; //CHANX 3 (1,7) #60
wire n11544_0;
wire n11545; //CHANX 3 (1,7) #61
wire n11545_0;
wire n11546; //CHANX 4 (1,7) #62
wire n11546_0;
wire n11546_1;
buffer_wire buffer_11546_1 (.in(n11546_0), .out(n11546_1));
wire n11547; //CHANX 4 (1,7) #63
wire n11547_0;
wire n11547_1;
buffer_wire buffer_11547_1 (.in(n11547_0), .out(n11547_1));
wire n11548; //CHANX 1 (1,7) #64
wire n11548_0;
wire n11549; //CHANX 1 (1,7) #65
wire n11549_0;
wire n11550; //CHANX 2 (1,7) #66
wire n11550_0;
wire n11551; //CHANX 2 (1,7) #67
wire n11551_0;
wire n11552; //CHANX 3 (1,7) #68
wire n11552_0;
wire n11553; //CHANX 3 (1,7) #69
wire n11553_0;
wire n11554; //CHANX 4 (1,7) #70
wire n11554_0;
wire n11554_1;
buffer_wire buffer_11554_1 (.in(n11554_0), .out(n11554_1));
wire n11555; //CHANX 4 (1,7) #71
wire n11555_0;
wire n11555_1;
buffer_wire buffer_11555_1 (.in(n11555_0), .out(n11555_1));
wire n11556; //CHANX 1 (1,7) #72
wire n11556_0;
wire n11557; //CHANX 1 (1,7) #73
wire n11557_0;
wire n11558; //CHANX 2 (1,7) #74
wire n11558_0;
wire n11559; //CHANX 2 (1,7) #75
wire n11559_0;
wire n11560; //CHANX 3 (1,7) #76
wire n11560_0;
wire n11561; //CHANX 3 (1,7) #77
wire n11561_0;
wire n11562; //CHANX 4 (1,7) #78
wire n11562_0;
wire n11562_1;
buffer_wire buffer_11562_1 (.in(n11562_0), .out(n11562_1));
wire n11563; //CHANX 4 (1,7) #79
wire n11563_0;
wire n11563_1;
buffer_wire buffer_11563_1 (.in(n11563_0), .out(n11563_1));
wire n11564; //CHANX 1 (1,7) #80
wire n11564_0;
wire n11565; //CHANX 1 (1,7) #81
wire n11565_0;
wire n11566; //CHANX 2 (1,7) #82
wire n11566_0;
wire n11567; //CHANX 2 (1,7) #83
wire n11567_0;
wire n11568; //CHANX 3 (1,7) #84
wire n11568_0;
wire n11569; //CHANX 3 (1,7) #85
wire n11569_0;
wire n11570; //CHANX 4 (1,7) #86
wire n11570_0;
wire n11570_1;
buffer_wire buffer_11570_1 (.in(n11570_0), .out(n11570_1));
wire n11571; //CHANX 4 (1,7) #87
wire n11571_0;
wire n11571_1;
buffer_wire buffer_11571_1 (.in(n11571_0), .out(n11571_1));
wire n11572; //CHANX 5 (1,7) #88
wire n11572_0;
wire n11572_1;
buffer_wire buffer_11572_1 (.in(n11572_0), .out(n11572_1));
wire n11573; //CHANX 5 (1,7) #89
wire n11573_0;
wire n11573_1;
buffer_wire buffer_11573_1 (.in(n11573_0), .out(n11573_1));
wire n11574; //CHANX 6 (1,7) #90
wire n11574_0;
wire n11574_1;
buffer_wire buffer_11574_1 (.in(n11574_0), .out(n11574_1));
wire n11575; //CHANX 6 (1,7) #91
wire n11575_0;
wire n11575_1;
buffer_wire buffer_11575_1 (.in(n11575_0), .out(n11575_1));
wire n11576; //CHANX 4 (2,7) #0
wire n11576_0;
wire n11576_1;
buffer_wire buffer_11576_1 (.in(n11576_0), .out(n11576_1));
wire n11577; //CHANX 4 (2,7) #1
wire n11577_0;
wire n11577_1;
buffer_wire buffer_11577_1 (.in(n11577_0), .out(n11577_1));
wire n11578; //CHANX 4 (2,7) #8
wire n11578_0;
wire n11578_1;
buffer_wire buffer_11578_1 (.in(n11578_0), .out(n11578_1));
wire n11579; //CHANX 4 (2,7) #9
wire n11579_0;
wire n11579_1;
buffer_wire buffer_11579_1 (.in(n11579_0), .out(n11579_1));
wire n11580; //CHANX 4 (2,7) #16
wire n11580_0;
wire n11580_1;
buffer_wire buffer_11580_1 (.in(n11580_0), .out(n11580_1));
wire n11581; //CHANX 4 (2,7) #17
wire n11581_0;
wire n11581_1;
buffer_wire buffer_11581_1 (.in(n11581_0), .out(n11581_1));
wire n11582; //CHANX 4 (2,7) #24
wire n11582_0;
wire n11582_1;
buffer_wire buffer_11582_1 (.in(n11582_0), .out(n11582_1));
wire n11583; //CHANX 4 (2,7) #25
wire n11583_0;
wire n11583_1;
buffer_wire buffer_11583_1 (.in(n11583_0), .out(n11583_1));
wire n11584; //CHANX 4 (2,7) #32
wire n11584_0;
wire n11584_1;
buffer_wire buffer_11584_1 (.in(n11584_0), .out(n11584_1));
wire n11585; //CHANX 4 (2,7) #33
wire n11585_0;
wire n11585_1;
buffer_wire buffer_11585_1 (.in(n11585_0), .out(n11585_1));
wire n11586; //CHANX 4 (2,7) #40
wire n11586_0;
wire n11586_1;
buffer_wire buffer_11586_1 (.in(n11586_0), .out(n11586_1));
wire n11587; //CHANX 4 (2,7) #41
wire n11587_0;
wire n11587_1;
buffer_wire buffer_11587_1 (.in(n11587_0), .out(n11587_1));
wire n11588; //CHANX 4 (2,7) #48
wire n11588_0;
wire n11588_1;
buffer_wire buffer_11588_1 (.in(n11588_0), .out(n11588_1));
wire n11589; //CHANX 4 (2,7) #49
wire n11589_0;
wire n11589_1;
buffer_wire buffer_11589_1 (.in(n11589_0), .out(n11589_1));
wire n11590; //CHANX 4 (2,7) #56
wire n11590_0;
wire n11590_1;
buffer_wire buffer_11590_1 (.in(n11590_0), .out(n11590_1));
wire n11591; //CHANX 4 (2,7) #57
wire n11591_0;
wire n11591_1;
buffer_wire buffer_11591_1 (.in(n11591_0), .out(n11591_1));
wire n11592; //CHANX 4 (2,7) #64
wire n11592_0;
wire n11592_1;
buffer_wire buffer_11592_1 (.in(n11592_0), .out(n11592_1));
wire n11593; //CHANX 4 (2,7) #65
wire n11593_0;
wire n11593_1;
buffer_wire buffer_11593_1 (.in(n11593_0), .out(n11593_1));
wire n11594; //CHANX 4 (2,7) #72
wire n11594_0;
wire n11594_1;
buffer_wire buffer_11594_1 (.in(n11594_0), .out(n11594_1));
wire n11595; //CHANX 4 (2,7) #73
wire n11595_0;
wire n11595_1;
buffer_wire buffer_11595_1 (.in(n11595_0), .out(n11595_1));
wire n11596; //CHANX 8 (2,7) #80
wire n11596_0;
wire n11596_1;
wire n11596_2;
buffer_wire buffer_11596_2 (.in(n11596_1), .out(n11596_2));
buffer_wire buffer_11596_1 (.in(n11596_0), .out(n11596_1));
wire n11597; //CHANX 8 (2,7) #81
wire n11597_0;
wire n11597_1;
wire n11597_2;
buffer_wire buffer_11597_2 (.in(n11597_1), .out(n11597_2));
buffer_wire buffer_11597_1 (.in(n11597_0), .out(n11597_1));
wire n11598; //CHANX 4 (3,7) #2
wire n11598_0;
wire n11598_1;
buffer_wire buffer_11598_1 (.in(n11598_0), .out(n11598_1));
wire n11599; //CHANX 4 (3,7) #3
wire n11599_0;
wire n11599_1;
buffer_wire buffer_11599_1 (.in(n11599_0), .out(n11599_1));
wire n11600; //CHANX 4 (3,7) #10
wire n11600_0;
wire n11600_1;
buffer_wire buffer_11600_1 (.in(n11600_0), .out(n11600_1));
wire n11601; //CHANX 4 (3,7) #11
wire n11601_0;
wire n11601_1;
buffer_wire buffer_11601_1 (.in(n11601_0), .out(n11601_1));
wire n11602; //CHANX 4 (3,7) #18
wire n11602_0;
wire n11602_1;
buffer_wire buffer_11602_1 (.in(n11602_0), .out(n11602_1));
wire n11603; //CHANX 4 (3,7) #19
wire n11603_0;
wire n11603_1;
buffer_wire buffer_11603_1 (.in(n11603_0), .out(n11603_1));
wire n11604; //CHANX 4 (3,7) #26
wire n11604_0;
wire n11604_1;
buffer_wire buffer_11604_1 (.in(n11604_0), .out(n11604_1));
wire n11605; //CHANX 4 (3,7) #27
wire n11605_0;
wire n11605_1;
buffer_wire buffer_11605_1 (.in(n11605_0), .out(n11605_1));
wire n11606; //CHANX 4 (3,7) #34
wire n11606_0;
wire n11606_1;
buffer_wire buffer_11606_1 (.in(n11606_0), .out(n11606_1));
wire n11607; //CHANX 4 (3,7) #35
wire n11607_0;
wire n11607_1;
buffer_wire buffer_11607_1 (.in(n11607_0), .out(n11607_1));
wire n11608; //CHANX 4 (3,7) #42
wire n11608_0;
wire n11608_1;
buffer_wire buffer_11608_1 (.in(n11608_0), .out(n11608_1));
wire n11609; //CHANX 4 (3,7) #43
wire n11609_0;
wire n11609_1;
buffer_wire buffer_11609_1 (.in(n11609_0), .out(n11609_1));
wire n11610; //CHANX 4 (3,7) #50
wire n11610_0;
wire n11610_1;
buffer_wire buffer_11610_1 (.in(n11610_0), .out(n11610_1));
wire n11611; //CHANX 4 (3,7) #51
wire n11611_0;
wire n11611_1;
buffer_wire buffer_11611_1 (.in(n11611_0), .out(n11611_1));
wire n11612; //CHANX 4 (3,7) #58
wire n11612_0;
wire n11612_1;
buffer_wire buffer_11612_1 (.in(n11612_0), .out(n11612_1));
wire n11613; //CHANX 4 (3,7) #59
wire n11613_0;
wire n11613_1;
buffer_wire buffer_11613_1 (.in(n11613_0), .out(n11613_1));
wire n11614; //CHANX 4 (3,7) #66
wire n11614_0;
wire n11614_1;
buffer_wire buffer_11614_1 (.in(n11614_0), .out(n11614_1));
wire n11615; //CHANX 4 (3,7) #67
wire n11615_0;
wire n11615_1;
buffer_wire buffer_11615_1 (.in(n11615_0), .out(n11615_1));
wire n11616; //CHANX 4 (3,7) #74
wire n11616_0;
wire n11616_1;
buffer_wire buffer_11616_1 (.in(n11616_0), .out(n11616_1));
wire n11617; //CHANX 4 (3,7) #75
wire n11617_0;
wire n11617_1;
buffer_wire buffer_11617_1 (.in(n11617_0), .out(n11617_1));
wire n11618; //CHANX 7 (3,7) #82
wire n11618_0;
wire n11618_1;
wire n11618_2;
buffer_wire buffer_11618_2 (.in(n11618_1), .out(n11618_2));
buffer_wire buffer_11618_1 (.in(n11618_0), .out(n11618_1));
wire n11619; //CHANX 7 (3,7) #83
wire n11619_0;
wire n11619_1;
wire n11619_2;
buffer_wire buffer_11619_2 (.in(n11619_1), .out(n11619_2));
buffer_wire buffer_11619_1 (.in(n11619_0), .out(n11619_1));
wire n11620; //CHANX 4 (4,7) #4
wire n11620_0;
wire n11620_1;
buffer_wire buffer_11620_1 (.in(n11620_0), .out(n11620_1));
wire n11621; //CHANX 4 (4,7) #5
wire n11621_0;
wire n11621_1;
buffer_wire buffer_11621_1 (.in(n11621_0), .out(n11621_1));
wire n11622; //CHANX 4 (4,7) #12
wire n11622_0;
wire n11622_1;
buffer_wire buffer_11622_1 (.in(n11622_0), .out(n11622_1));
wire n11623; //CHANX 4 (4,7) #13
wire n11623_0;
wire n11623_1;
buffer_wire buffer_11623_1 (.in(n11623_0), .out(n11623_1));
wire n11624; //CHANX 4 (4,7) #20
wire n11624_0;
wire n11624_1;
buffer_wire buffer_11624_1 (.in(n11624_0), .out(n11624_1));
wire n11625; //CHANX 4 (4,7) #21
wire n11625_0;
wire n11625_1;
buffer_wire buffer_11625_1 (.in(n11625_0), .out(n11625_1));
wire n11626; //CHANX 4 (4,7) #28
wire n11626_0;
wire n11626_1;
buffer_wire buffer_11626_1 (.in(n11626_0), .out(n11626_1));
wire n11627; //CHANX 4 (4,7) #29
wire n11627_0;
wire n11627_1;
buffer_wire buffer_11627_1 (.in(n11627_0), .out(n11627_1));
wire n11628; //CHANX 4 (4,7) #36
wire n11628_0;
wire n11628_1;
buffer_wire buffer_11628_1 (.in(n11628_0), .out(n11628_1));
wire n11629; //CHANX 4 (4,7) #37
wire n11629_0;
wire n11629_1;
buffer_wire buffer_11629_1 (.in(n11629_0), .out(n11629_1));
wire n11630; //CHANX 4 (4,7) #44
wire n11630_0;
wire n11630_1;
buffer_wire buffer_11630_1 (.in(n11630_0), .out(n11630_1));
wire n11631; //CHANX 4 (4,7) #45
wire n11631_0;
wire n11631_1;
buffer_wire buffer_11631_1 (.in(n11631_0), .out(n11631_1));
wire n11632; //CHANX 4 (4,7) #52
wire n11632_0;
wire n11632_1;
buffer_wire buffer_11632_1 (.in(n11632_0), .out(n11632_1));
wire n11633; //CHANX 4 (4,7) #53
wire n11633_0;
wire n11633_1;
buffer_wire buffer_11633_1 (.in(n11633_0), .out(n11633_1));
wire n11634; //CHANX 4 (4,7) #60
wire n11634_0;
wire n11634_1;
buffer_wire buffer_11634_1 (.in(n11634_0), .out(n11634_1));
wire n11635; //CHANX 4 (4,7) #61
wire n11635_0;
wire n11635_1;
buffer_wire buffer_11635_1 (.in(n11635_0), .out(n11635_1));
wire n11636; //CHANX 4 (4,7) #68
wire n11636_0;
wire n11636_1;
buffer_wire buffer_11636_1 (.in(n11636_0), .out(n11636_1));
wire n11637; //CHANX 4 (4,7) #69
wire n11637_0;
wire n11637_1;
buffer_wire buffer_11637_1 (.in(n11637_0), .out(n11637_1));
wire n11638; //CHANX 4 (4,7) #76
wire n11638_0;
wire n11638_1;
buffer_wire buffer_11638_1 (.in(n11638_0), .out(n11638_1));
wire n11639; //CHANX 4 (4,7) #77
wire n11639_0;
wire n11639_1;
buffer_wire buffer_11639_1 (.in(n11639_0), .out(n11639_1));
wire n11640; //CHANX 6 (4,7) #84
wire n11640_0;
wire n11640_1;
buffer_wire buffer_11640_1 (.in(n11640_0), .out(n11640_1));
wire n11641; //CHANX 6 (4,7) #85
wire n11641_0;
wire n11641_1;
buffer_wire buffer_11641_1 (.in(n11641_0), .out(n11641_1));
wire n11642; //CHANX 4 (5,7) #6
wire n11642_0;
wire n11642_1;
buffer_wire buffer_11642_1 (.in(n11642_0), .out(n11642_1));
wire n11643; //CHANX 4 (5,7) #7
wire n11643_0;
wire n11643_1;
buffer_wire buffer_11643_1 (.in(n11643_0), .out(n11643_1));
wire n11644; //CHANX 4 (5,7) #14
wire n11644_0;
wire n11644_1;
buffer_wire buffer_11644_1 (.in(n11644_0), .out(n11644_1));
wire n11645; //CHANX 4 (5,7) #15
wire n11645_0;
wire n11645_1;
buffer_wire buffer_11645_1 (.in(n11645_0), .out(n11645_1));
wire n11646; //CHANX 4 (5,7) #22
wire n11646_0;
wire n11646_1;
buffer_wire buffer_11646_1 (.in(n11646_0), .out(n11646_1));
wire n11647; //CHANX 4 (5,7) #23
wire n11647_0;
wire n11647_1;
buffer_wire buffer_11647_1 (.in(n11647_0), .out(n11647_1));
wire n11648; //CHANX 4 (5,7) #30
wire n11648_0;
wire n11648_1;
buffer_wire buffer_11648_1 (.in(n11648_0), .out(n11648_1));
wire n11649; //CHANX 4 (5,7) #31
wire n11649_0;
wire n11649_1;
buffer_wire buffer_11649_1 (.in(n11649_0), .out(n11649_1));
wire n11650; //CHANX 4 (5,7) #38
wire n11650_0;
wire n11650_1;
buffer_wire buffer_11650_1 (.in(n11650_0), .out(n11650_1));
wire n11651; //CHANX 4 (5,7) #39
wire n11651_0;
wire n11651_1;
buffer_wire buffer_11651_1 (.in(n11651_0), .out(n11651_1));
wire n11652; //CHANX 4 (5,7) #46
wire n11652_0;
wire n11652_1;
buffer_wire buffer_11652_1 (.in(n11652_0), .out(n11652_1));
wire n11653; //CHANX 4 (5,7) #47
wire n11653_0;
wire n11653_1;
buffer_wire buffer_11653_1 (.in(n11653_0), .out(n11653_1));
wire n11654; //CHANX 4 (5,7) #54
wire n11654_0;
wire n11654_1;
buffer_wire buffer_11654_1 (.in(n11654_0), .out(n11654_1));
wire n11655; //CHANX 4 (5,7) #55
wire n11655_0;
wire n11655_1;
buffer_wire buffer_11655_1 (.in(n11655_0), .out(n11655_1));
wire n11656; //CHANX 4 (5,7) #62
wire n11656_0;
wire n11656_1;
buffer_wire buffer_11656_1 (.in(n11656_0), .out(n11656_1));
wire n11657; //CHANX 4 (5,7) #63
wire n11657_0;
wire n11657_1;
buffer_wire buffer_11657_1 (.in(n11657_0), .out(n11657_1));
wire n11658; //CHANX 4 (5,7) #70
wire n11658_0;
wire n11658_1;
buffer_wire buffer_11658_1 (.in(n11658_0), .out(n11658_1));
wire n11659; //CHANX 4 (5,7) #71
wire n11659_0;
wire n11659_1;
buffer_wire buffer_11659_1 (.in(n11659_0), .out(n11659_1));
wire n11660; //CHANX 4 (5,7) #78
wire n11660_0;
wire n11660_1;
buffer_wire buffer_11660_1 (.in(n11660_0), .out(n11660_1));
wire n11661; //CHANX 4 (5,7) #79
wire n11661_0;
wire n11661_1;
buffer_wire buffer_11661_1 (.in(n11661_0), .out(n11661_1));
wire n11662; //CHANX 5 (5,7) #86
wire n11662_0;
wire n11662_1;
buffer_wire buffer_11662_1 (.in(n11662_0), .out(n11662_1));
wire n11663; //CHANX 5 (5,7) #87
wire n11663_0;
wire n11663_1;
buffer_wire buffer_11663_1 (.in(n11663_0), .out(n11663_1));
wire n11664; //CHANX 4 (6,7) #0
wire n11664_0;
wire n11664_1;
buffer_wire buffer_11664_1 (.in(n11664_0), .out(n11664_1));
wire n11665; //CHANX 4 (6,7) #1
wire n11665_0;
wire n11665_1;
buffer_wire buffer_11665_1 (.in(n11665_0), .out(n11665_1));
wire n11666; //CHANX 4 (6,7) #8
wire n11666_0;
wire n11666_1;
buffer_wire buffer_11666_1 (.in(n11666_0), .out(n11666_1));
wire n11667; //CHANX 4 (6,7) #9
wire n11667_0;
wire n11667_1;
buffer_wire buffer_11667_1 (.in(n11667_0), .out(n11667_1));
wire n11668; //CHANX 4 (6,7) #16
wire n11668_0;
wire n11668_1;
buffer_wire buffer_11668_1 (.in(n11668_0), .out(n11668_1));
wire n11669; //CHANX 4 (6,7) #17
wire n11669_0;
wire n11669_1;
buffer_wire buffer_11669_1 (.in(n11669_0), .out(n11669_1));
wire n11670; //CHANX 4 (6,7) #24
wire n11670_0;
wire n11670_1;
buffer_wire buffer_11670_1 (.in(n11670_0), .out(n11670_1));
wire n11671; //CHANX 4 (6,7) #25
wire n11671_0;
wire n11671_1;
buffer_wire buffer_11671_1 (.in(n11671_0), .out(n11671_1));
wire n11672; //CHANX 4 (6,7) #32
wire n11672_0;
wire n11672_1;
buffer_wire buffer_11672_1 (.in(n11672_0), .out(n11672_1));
wire n11673; //CHANX 4 (6,7) #33
wire n11673_0;
wire n11673_1;
buffer_wire buffer_11673_1 (.in(n11673_0), .out(n11673_1));
wire n11674; //CHANX 4 (6,7) #40
wire n11674_0;
wire n11674_1;
buffer_wire buffer_11674_1 (.in(n11674_0), .out(n11674_1));
wire n11675; //CHANX 4 (6,7) #41
wire n11675_0;
wire n11675_1;
buffer_wire buffer_11675_1 (.in(n11675_0), .out(n11675_1));
wire n11676; //CHANX 4 (6,7) #48
wire n11676_0;
wire n11676_1;
buffer_wire buffer_11676_1 (.in(n11676_0), .out(n11676_1));
wire n11677; //CHANX 4 (6,7) #49
wire n11677_0;
wire n11677_1;
buffer_wire buffer_11677_1 (.in(n11677_0), .out(n11677_1));
wire n11678; //CHANX 4 (6,7) #56
wire n11678_0;
wire n11678_1;
buffer_wire buffer_11678_1 (.in(n11678_0), .out(n11678_1));
wire n11679; //CHANX 4 (6,7) #57
wire n11679_0;
wire n11679_1;
buffer_wire buffer_11679_1 (.in(n11679_0), .out(n11679_1));
wire n11680; //CHANX 4 (6,7) #64
wire n11680_0;
wire n11680_1;
buffer_wire buffer_11680_1 (.in(n11680_0), .out(n11680_1));
wire n11681; //CHANX 4 (6,7) #65
wire n11681_0;
wire n11681_1;
buffer_wire buffer_11681_1 (.in(n11681_0), .out(n11681_1));
wire n11682; //CHANX 4 (6,7) #72
wire n11682_0;
wire n11682_1;
buffer_wire buffer_11682_1 (.in(n11682_0), .out(n11682_1));
wire n11683; //CHANX 4 (6,7) #73
wire n11683_0;
wire n11683_1;
buffer_wire buffer_11683_1 (.in(n11683_0), .out(n11683_1));
wire n11684; //CHANX 4 (6,7) #88
wire n11684_0;
wire n11684_1;
buffer_wire buffer_11684_1 (.in(n11684_0), .out(n11684_1));
wire n11685; //CHANX 4 (6,7) #89
wire n11685_0;
wire n11685_1;
buffer_wire buffer_11685_1 (.in(n11685_0), .out(n11685_1));
wire n11686; //CHANX 3 (7,7) #2
wire n11686_0;
wire n11687; //CHANX 3 (7,7) #3
wire n11687_0;
wire n11688; //CHANX 3 (7,7) #10
wire n11688_0;
wire n11689; //CHANX 3 (7,7) #11
wire n11689_0;
wire n11690; //CHANX 3 (7,7) #18
wire n11690_0;
wire n11691; //CHANX 3 (7,7) #19
wire n11691_0;
wire n11692; //CHANX 3 (7,7) #26
wire n11692_0;
wire n11693; //CHANX 3 (7,7) #27
wire n11693_0;
wire n11694; //CHANX 3 (7,7) #34
wire n11694_0;
wire n11695; //CHANX 3 (7,7) #35
wire n11695_0;
wire n11696; //CHANX 3 (7,7) #42
wire n11696_0;
wire n11697; //CHANX 3 (7,7) #43
wire n11697_0;
wire n11698; //CHANX 3 (7,7) #50
wire n11698_0;
wire n11699; //CHANX 3 (7,7) #51
wire n11699_0;
wire n11700; //CHANX 3 (7,7) #58
wire n11700_0;
wire n11701; //CHANX 3 (7,7) #59
wire n11701_0;
wire n11702; //CHANX 3 (7,7) #66
wire n11702_0;
wire n11703; //CHANX 3 (7,7) #67
wire n11703_0;
wire n11704; //CHANX 3 (7,7) #74
wire n11704_0;
wire n11705; //CHANX 3 (7,7) #75
wire n11705_0;
wire n11706; //CHANX 3 (7,7) #90
wire n11706_0;
wire n11707; //CHANX 3 (7,7) #91
wire n11707_0;
wire n11708; //CHANX 2 (8,7) #4
wire n11708_0;
wire n11709; //CHANX 2 (8,7) #5
wire n11709_0;
wire n11710; //CHANX 2 (8,7) #12
wire n11710_0;
wire n11711; //CHANX 2 (8,7) #13
wire n11711_0;
wire n11712; //CHANX 2 (8,7) #20
wire n11712_0;
wire n11713; //CHANX 2 (8,7) #21
wire n11713_0;
wire n11714; //CHANX 2 (8,7) #28
wire n11714_0;
wire n11715; //CHANX 2 (8,7) #29
wire n11715_0;
wire n11716; //CHANX 2 (8,7) #36
wire n11716_0;
wire n11717; //CHANX 2 (8,7) #37
wire n11717_0;
wire n11718; //CHANX 2 (8,7) #44
wire n11718_0;
wire n11719; //CHANX 2 (8,7) #45
wire n11719_0;
wire n11720; //CHANX 2 (8,7) #52
wire n11720_0;
wire n11721; //CHANX 2 (8,7) #53
wire n11721_0;
wire n11722; //CHANX 2 (8,7) #60
wire n11722_0;
wire n11723; //CHANX 2 (8,7) #61
wire n11723_0;
wire n11724; //CHANX 2 (8,7) #68
wire n11724_0;
wire n11725; //CHANX 2 (8,7) #69
wire n11725_0;
wire n11726; //CHANX 2 (8,7) #76
wire n11726_0;
wire n11727; //CHANX 2 (8,7) #77
wire n11727_0;
wire n11728; //CHANX 1 (9,7) #6
wire n11728_0;
wire n11729; //CHANX 1 (9,7) #7
wire n11729_0;
wire n11730; //CHANX 1 (9,7) #14
wire n11730_0;
wire n11731; //CHANX 1 (9,7) #15
wire n11731_0;
wire n11732; //CHANX 1 (9,7) #22
wire n11732_0;
wire n11733; //CHANX 1 (9,7) #23
wire n11733_0;
wire n11734; //CHANX 1 (9,7) #30
wire n11734_0;
wire n11735; //CHANX 1 (9,7) #31
wire n11735_0;
wire n11736; //CHANX 1 (9,7) #38
wire n11736_0;
wire n11737; //CHANX 1 (9,7) #39
wire n11737_0;
wire n11738; //CHANX 1 (9,7) #46
wire n11738_0;
wire n11739; //CHANX 1 (9,7) #47
wire n11739_0;
wire n11740; //CHANX 1 (9,7) #54
wire n11740_0;
wire n11741; //CHANX 1 (9,7) #55
wire n11741_0;
wire n11742; //CHANX 1 (9,7) #62
wire n11742_0;
wire n11743; //CHANX 1 (9,7) #63
wire n11743_0;
wire n11744; //CHANX 1 (9,7) #70
wire n11744_0;
wire n11745; //CHANX 1 (9,7) #71
wire n11745_0;
wire n11746; //CHANX 1 (9,7) #78
wire n11746_0;
wire n11747; //CHANX 1 (9,7) #79
wire n11747_0;
wire n11748; //CHANX 4 (1,8) #0
wire n11748_0;
wire n11748_1;
buffer_wire buffer_11748_1 (.in(n11748_0), .out(n11748_1));
wire n11749; //CHANX 4 (1,8) #1
wire n11749_0;
wire n11749_1;
buffer_wire buffer_11749_1 (.in(n11749_0), .out(n11749_1));
wire n11750; //CHANX 1 (1,8) #2
wire n11750_0;
wire n11751; //CHANX 1 (1,8) #3
wire n11751_0;
wire n11752; //CHANX 2 (1,8) #4
wire n11752_0;
wire n11753; //CHANX 2 (1,8) #5
wire n11753_0;
wire n11754; //CHANX 3 (1,8) #6
wire n11754_0;
wire n11755; //CHANX 3 (1,8) #7
wire n11755_0;
wire n11756; //CHANX 4 (1,8) #8
wire n11756_0;
wire n11756_1;
buffer_wire buffer_11756_1 (.in(n11756_0), .out(n11756_1));
wire n11757; //CHANX 4 (1,8) #9
wire n11757_0;
wire n11757_1;
buffer_wire buffer_11757_1 (.in(n11757_0), .out(n11757_1));
wire n11758; //CHANX 1 (1,8) #10
wire n11758_0;
wire n11759; //CHANX 1 (1,8) #11
wire n11759_0;
wire n11760; //CHANX 2 (1,8) #12
wire n11760_0;
wire n11761; //CHANX 2 (1,8) #13
wire n11761_0;
wire n11762; //CHANX 3 (1,8) #14
wire n11762_0;
wire n11763; //CHANX 3 (1,8) #15
wire n11763_0;
wire n11764; //CHANX 4 (1,8) #16
wire n11764_0;
wire n11764_1;
buffer_wire buffer_11764_1 (.in(n11764_0), .out(n11764_1));
wire n11765; //CHANX 4 (1,8) #17
wire n11765_0;
wire n11765_1;
buffer_wire buffer_11765_1 (.in(n11765_0), .out(n11765_1));
wire n11766; //CHANX 1 (1,8) #18
wire n11766_0;
wire n11767; //CHANX 1 (1,8) #19
wire n11767_0;
wire n11768; //CHANX 2 (1,8) #20
wire n11768_0;
wire n11769; //CHANX 2 (1,8) #21
wire n11769_0;
wire n11770; //CHANX 3 (1,8) #22
wire n11770_0;
wire n11771; //CHANX 3 (1,8) #23
wire n11771_0;
wire n11772; //CHANX 4 (1,8) #24
wire n11772_0;
wire n11772_1;
buffer_wire buffer_11772_1 (.in(n11772_0), .out(n11772_1));
wire n11773; //CHANX 4 (1,8) #25
wire n11773_0;
wire n11773_1;
buffer_wire buffer_11773_1 (.in(n11773_0), .out(n11773_1));
wire n11774; //CHANX 1 (1,8) #26
wire n11774_0;
wire n11775; //CHANX 1 (1,8) #27
wire n11775_0;
wire n11776; //CHANX 2 (1,8) #28
wire n11776_0;
wire n11777; //CHANX 2 (1,8) #29
wire n11777_0;
wire n11778; //CHANX 3 (1,8) #30
wire n11778_0;
wire n11779; //CHANX 3 (1,8) #31
wire n11779_0;
wire n11780; //CHANX 4 (1,8) #32
wire n11780_0;
wire n11780_1;
buffer_wire buffer_11780_1 (.in(n11780_0), .out(n11780_1));
wire n11781; //CHANX 4 (1,8) #33
wire n11781_0;
wire n11781_1;
buffer_wire buffer_11781_1 (.in(n11781_0), .out(n11781_1));
wire n11782; //CHANX 1 (1,8) #34
wire n11782_0;
wire n11783; //CHANX 1 (1,8) #35
wire n11783_0;
wire n11784; //CHANX 2 (1,8) #36
wire n11784_0;
wire n11785; //CHANX 2 (1,8) #37
wire n11785_0;
wire n11786; //CHANX 3 (1,8) #38
wire n11786_0;
wire n11787; //CHANX 3 (1,8) #39
wire n11787_0;
wire n11788; //CHANX 4 (1,8) #40
wire n11788_0;
wire n11788_1;
buffer_wire buffer_11788_1 (.in(n11788_0), .out(n11788_1));
wire n11789; //CHANX 4 (1,8) #41
wire n11789_0;
wire n11789_1;
buffer_wire buffer_11789_1 (.in(n11789_0), .out(n11789_1));
wire n11790; //CHANX 1 (1,8) #42
wire n11790_0;
wire n11791; //CHANX 1 (1,8) #43
wire n11791_0;
wire n11792; //CHANX 2 (1,8) #44
wire n11792_0;
wire n11793; //CHANX 2 (1,8) #45
wire n11793_0;
wire n11794; //CHANX 3 (1,8) #46
wire n11794_0;
wire n11795; //CHANX 3 (1,8) #47
wire n11795_0;
wire n11796; //CHANX 4 (1,8) #48
wire n11796_0;
wire n11796_1;
buffer_wire buffer_11796_1 (.in(n11796_0), .out(n11796_1));
wire n11797; //CHANX 4 (1,8) #49
wire n11797_0;
wire n11797_1;
buffer_wire buffer_11797_1 (.in(n11797_0), .out(n11797_1));
wire n11798; //CHANX 1 (1,8) #50
wire n11798_0;
wire n11799; //CHANX 1 (1,8) #51
wire n11799_0;
wire n11800; //CHANX 2 (1,8) #52
wire n11800_0;
wire n11801; //CHANX 2 (1,8) #53
wire n11801_0;
wire n11802; //CHANX 3 (1,8) #54
wire n11802_0;
wire n11803; //CHANX 3 (1,8) #55
wire n11803_0;
wire n11804; //CHANX 4 (1,8) #56
wire n11804_0;
wire n11804_1;
buffer_wire buffer_11804_1 (.in(n11804_0), .out(n11804_1));
wire n11805; //CHANX 4 (1,8) #57
wire n11805_0;
wire n11805_1;
buffer_wire buffer_11805_1 (.in(n11805_0), .out(n11805_1));
wire n11806; //CHANX 1 (1,8) #58
wire n11806_0;
wire n11807; //CHANX 1 (1,8) #59
wire n11807_0;
wire n11808; //CHANX 2 (1,8) #60
wire n11808_0;
wire n11809; //CHANX 2 (1,8) #61
wire n11809_0;
wire n11810; //CHANX 3 (1,8) #62
wire n11810_0;
wire n11811; //CHANX 3 (1,8) #63
wire n11811_0;
wire n11812; //CHANX 4 (1,8) #64
wire n11812_0;
wire n11812_1;
buffer_wire buffer_11812_1 (.in(n11812_0), .out(n11812_1));
wire n11813; //CHANX 4 (1,8) #65
wire n11813_0;
wire n11813_1;
buffer_wire buffer_11813_1 (.in(n11813_0), .out(n11813_1));
wire n11814; //CHANX 1 (1,8) #66
wire n11814_0;
wire n11815; //CHANX 1 (1,8) #67
wire n11815_0;
wire n11816; //CHANX 2 (1,8) #68
wire n11816_0;
wire n11817; //CHANX 2 (1,8) #69
wire n11817_0;
wire n11818; //CHANX 3 (1,8) #70
wire n11818_0;
wire n11819; //CHANX 3 (1,8) #71
wire n11819_0;
wire n11820; //CHANX 4 (1,8) #72
wire n11820_0;
wire n11820_1;
buffer_wire buffer_11820_1 (.in(n11820_0), .out(n11820_1));
wire n11821; //CHANX 4 (1,8) #73
wire n11821_0;
wire n11821_1;
buffer_wire buffer_11821_1 (.in(n11821_0), .out(n11821_1));
wire n11822; //CHANX 1 (1,8) #74
wire n11822_0;
wire n11823; //CHANX 1 (1,8) #75
wire n11823_0;
wire n11824; //CHANX 2 (1,8) #76
wire n11824_0;
wire n11825; //CHANX 2 (1,8) #77
wire n11825_0;
wire n11826; //CHANX 3 (1,8) #78
wire n11826_0;
wire n11827; //CHANX 3 (1,8) #79
wire n11827_0;
wire n11828; //CHANX 9 (1,8) #80
wire n11828_0;
wire n11828_1;
wire n11828_2;
buffer_wire buffer_11828_2 (.in(n11828_1), .out(n11828_2));
buffer_wire buffer_11828_1 (.in(n11828_0), .out(n11828_1));
wire n11829; //CHANX 9 (1,8) #81
wire n11829_0;
wire n11829_1;
wire n11829_2;
buffer_wire buffer_11829_2 (.in(n11829_1), .out(n11829_2));
buffer_wire buffer_11829_1 (.in(n11829_0), .out(n11829_1));
wire n11830; //CHANX 1 (1,8) #82
wire n11830_0;
wire n11831; //CHANX 1 (1,8) #83
wire n11831_0;
wire n11832; //CHANX 2 (1,8) #84
wire n11832_0;
wire n11833; //CHANX 2 (1,8) #85
wire n11833_0;
wire n11834; //CHANX 3 (1,8) #86
wire n11834_0;
wire n11835; //CHANX 3 (1,8) #87
wire n11835_0;
wire n11836; //CHANX 4 (1,8) #88
wire n11836_0;
wire n11836_1;
buffer_wire buffer_11836_1 (.in(n11836_0), .out(n11836_1));
wire n11837; //CHANX 4 (1,8) #89
wire n11837_0;
wire n11837_1;
buffer_wire buffer_11837_1 (.in(n11837_0), .out(n11837_1));
wire n11838; //CHANX 5 (1,8) #90
wire n11838_0;
wire n11838_1;
buffer_wire buffer_11838_1 (.in(n11838_0), .out(n11838_1));
wire n11839; //CHANX 5 (1,8) #91
wire n11839_0;
wire n11839_1;
buffer_wire buffer_11839_1 (.in(n11839_0), .out(n11839_1));
wire n11840; //CHANX 4 (2,8) #2
wire n11840_0;
wire n11840_1;
buffer_wire buffer_11840_1 (.in(n11840_0), .out(n11840_1));
wire n11841; //CHANX 4 (2,8) #3
wire n11841_0;
wire n11841_1;
buffer_wire buffer_11841_1 (.in(n11841_0), .out(n11841_1));
wire n11842; //CHANX 4 (2,8) #10
wire n11842_0;
wire n11842_1;
buffer_wire buffer_11842_1 (.in(n11842_0), .out(n11842_1));
wire n11843; //CHANX 4 (2,8) #11
wire n11843_0;
wire n11843_1;
buffer_wire buffer_11843_1 (.in(n11843_0), .out(n11843_1));
wire n11844; //CHANX 4 (2,8) #18
wire n11844_0;
wire n11844_1;
buffer_wire buffer_11844_1 (.in(n11844_0), .out(n11844_1));
wire n11845; //CHANX 4 (2,8) #19
wire n11845_0;
wire n11845_1;
buffer_wire buffer_11845_1 (.in(n11845_0), .out(n11845_1));
wire n11846; //CHANX 4 (2,8) #26
wire n11846_0;
wire n11846_1;
buffer_wire buffer_11846_1 (.in(n11846_0), .out(n11846_1));
wire n11847; //CHANX 4 (2,8) #27
wire n11847_0;
wire n11847_1;
buffer_wire buffer_11847_1 (.in(n11847_0), .out(n11847_1));
wire n11848; //CHANX 4 (2,8) #34
wire n11848_0;
wire n11848_1;
buffer_wire buffer_11848_1 (.in(n11848_0), .out(n11848_1));
wire n11849; //CHANX 4 (2,8) #35
wire n11849_0;
wire n11849_1;
buffer_wire buffer_11849_1 (.in(n11849_0), .out(n11849_1));
wire n11850; //CHANX 4 (2,8) #42
wire n11850_0;
wire n11850_1;
buffer_wire buffer_11850_1 (.in(n11850_0), .out(n11850_1));
wire n11851; //CHANX 4 (2,8) #43
wire n11851_0;
wire n11851_1;
buffer_wire buffer_11851_1 (.in(n11851_0), .out(n11851_1));
wire n11852; //CHANX 4 (2,8) #50
wire n11852_0;
wire n11852_1;
buffer_wire buffer_11852_1 (.in(n11852_0), .out(n11852_1));
wire n11853; //CHANX 4 (2,8) #51
wire n11853_0;
wire n11853_1;
buffer_wire buffer_11853_1 (.in(n11853_0), .out(n11853_1));
wire n11854; //CHANX 4 (2,8) #58
wire n11854_0;
wire n11854_1;
buffer_wire buffer_11854_1 (.in(n11854_0), .out(n11854_1));
wire n11855; //CHANX 4 (2,8) #59
wire n11855_0;
wire n11855_1;
buffer_wire buffer_11855_1 (.in(n11855_0), .out(n11855_1));
wire n11856; //CHANX 4 (2,8) #66
wire n11856_0;
wire n11856_1;
buffer_wire buffer_11856_1 (.in(n11856_0), .out(n11856_1));
wire n11857; //CHANX 4 (2,8) #67
wire n11857_0;
wire n11857_1;
buffer_wire buffer_11857_1 (.in(n11857_0), .out(n11857_1));
wire n11858; //CHANX 4 (2,8) #74
wire n11858_0;
wire n11858_1;
buffer_wire buffer_11858_1 (.in(n11858_0), .out(n11858_1));
wire n11859; //CHANX 4 (2,8) #75
wire n11859_0;
wire n11859_1;
buffer_wire buffer_11859_1 (.in(n11859_0), .out(n11859_1));
wire n11860; //CHANX 8 (2,8) #82
wire n11860_0;
wire n11860_1;
wire n11860_2;
buffer_wire buffer_11860_2 (.in(n11860_1), .out(n11860_2));
buffer_wire buffer_11860_1 (.in(n11860_0), .out(n11860_1));
wire n11861; //CHANX 8 (2,8) #83
wire n11861_0;
wire n11861_1;
wire n11861_2;
buffer_wire buffer_11861_2 (.in(n11861_1), .out(n11861_2));
buffer_wire buffer_11861_1 (.in(n11861_0), .out(n11861_1));
wire n11862; //CHANX 4 (3,8) #4
wire n11862_0;
wire n11862_1;
buffer_wire buffer_11862_1 (.in(n11862_0), .out(n11862_1));
wire n11863; //CHANX 4 (3,8) #5
wire n11863_0;
wire n11863_1;
buffer_wire buffer_11863_1 (.in(n11863_0), .out(n11863_1));
wire n11864; //CHANX 4 (3,8) #12
wire n11864_0;
wire n11864_1;
buffer_wire buffer_11864_1 (.in(n11864_0), .out(n11864_1));
wire n11865; //CHANX 4 (3,8) #13
wire n11865_0;
wire n11865_1;
buffer_wire buffer_11865_1 (.in(n11865_0), .out(n11865_1));
wire n11866; //CHANX 4 (3,8) #20
wire n11866_0;
wire n11866_1;
buffer_wire buffer_11866_1 (.in(n11866_0), .out(n11866_1));
wire n11867; //CHANX 4 (3,8) #21
wire n11867_0;
wire n11867_1;
buffer_wire buffer_11867_1 (.in(n11867_0), .out(n11867_1));
wire n11868; //CHANX 4 (3,8) #28
wire n11868_0;
wire n11868_1;
buffer_wire buffer_11868_1 (.in(n11868_0), .out(n11868_1));
wire n11869; //CHANX 4 (3,8) #29
wire n11869_0;
wire n11869_1;
buffer_wire buffer_11869_1 (.in(n11869_0), .out(n11869_1));
wire n11870; //CHANX 4 (3,8) #36
wire n11870_0;
wire n11870_1;
buffer_wire buffer_11870_1 (.in(n11870_0), .out(n11870_1));
wire n11871; //CHANX 4 (3,8) #37
wire n11871_0;
wire n11871_1;
buffer_wire buffer_11871_1 (.in(n11871_0), .out(n11871_1));
wire n11872; //CHANX 4 (3,8) #44
wire n11872_0;
wire n11872_1;
buffer_wire buffer_11872_1 (.in(n11872_0), .out(n11872_1));
wire n11873; //CHANX 4 (3,8) #45
wire n11873_0;
wire n11873_1;
buffer_wire buffer_11873_1 (.in(n11873_0), .out(n11873_1));
wire n11874; //CHANX 4 (3,8) #52
wire n11874_0;
wire n11874_1;
buffer_wire buffer_11874_1 (.in(n11874_0), .out(n11874_1));
wire n11875; //CHANX 4 (3,8) #53
wire n11875_0;
wire n11875_1;
buffer_wire buffer_11875_1 (.in(n11875_0), .out(n11875_1));
wire n11876; //CHANX 4 (3,8) #60
wire n11876_0;
wire n11876_1;
buffer_wire buffer_11876_1 (.in(n11876_0), .out(n11876_1));
wire n11877; //CHANX 4 (3,8) #61
wire n11877_0;
wire n11877_1;
buffer_wire buffer_11877_1 (.in(n11877_0), .out(n11877_1));
wire n11878; //CHANX 4 (3,8) #68
wire n11878_0;
wire n11878_1;
buffer_wire buffer_11878_1 (.in(n11878_0), .out(n11878_1));
wire n11879; //CHANX 4 (3,8) #69
wire n11879_0;
wire n11879_1;
buffer_wire buffer_11879_1 (.in(n11879_0), .out(n11879_1));
wire n11880; //CHANX 4 (3,8) #76
wire n11880_0;
wire n11880_1;
buffer_wire buffer_11880_1 (.in(n11880_0), .out(n11880_1));
wire n11881; //CHANX 4 (3,8) #77
wire n11881_0;
wire n11881_1;
buffer_wire buffer_11881_1 (.in(n11881_0), .out(n11881_1));
wire n11882; //CHANX 7 (3,8) #84
wire n11882_0;
wire n11882_1;
wire n11882_2;
buffer_wire buffer_11882_2 (.in(n11882_1), .out(n11882_2));
buffer_wire buffer_11882_1 (.in(n11882_0), .out(n11882_1));
wire n11883; //CHANX 7 (3,8) #85
wire n11883_0;
wire n11883_1;
wire n11883_2;
buffer_wire buffer_11883_2 (.in(n11883_1), .out(n11883_2));
buffer_wire buffer_11883_1 (.in(n11883_0), .out(n11883_1));
wire n11884; //CHANX 4 (4,8) #6
wire n11884_0;
wire n11884_1;
buffer_wire buffer_11884_1 (.in(n11884_0), .out(n11884_1));
wire n11885; //CHANX 4 (4,8) #7
wire n11885_0;
wire n11885_1;
buffer_wire buffer_11885_1 (.in(n11885_0), .out(n11885_1));
wire n11886; //CHANX 4 (4,8) #14
wire n11886_0;
wire n11886_1;
buffer_wire buffer_11886_1 (.in(n11886_0), .out(n11886_1));
wire n11887; //CHANX 4 (4,8) #15
wire n11887_0;
wire n11887_1;
buffer_wire buffer_11887_1 (.in(n11887_0), .out(n11887_1));
wire n11888; //CHANX 4 (4,8) #22
wire n11888_0;
wire n11888_1;
buffer_wire buffer_11888_1 (.in(n11888_0), .out(n11888_1));
wire n11889; //CHANX 4 (4,8) #23
wire n11889_0;
wire n11889_1;
buffer_wire buffer_11889_1 (.in(n11889_0), .out(n11889_1));
wire n11890; //CHANX 4 (4,8) #30
wire n11890_0;
wire n11890_1;
buffer_wire buffer_11890_1 (.in(n11890_0), .out(n11890_1));
wire n11891; //CHANX 4 (4,8) #31
wire n11891_0;
wire n11891_1;
buffer_wire buffer_11891_1 (.in(n11891_0), .out(n11891_1));
wire n11892; //CHANX 4 (4,8) #38
wire n11892_0;
wire n11892_1;
buffer_wire buffer_11892_1 (.in(n11892_0), .out(n11892_1));
wire n11893; //CHANX 4 (4,8) #39
wire n11893_0;
wire n11893_1;
buffer_wire buffer_11893_1 (.in(n11893_0), .out(n11893_1));
wire n11894; //CHANX 4 (4,8) #46
wire n11894_0;
wire n11894_1;
buffer_wire buffer_11894_1 (.in(n11894_0), .out(n11894_1));
wire n11895; //CHANX 4 (4,8) #47
wire n11895_0;
wire n11895_1;
buffer_wire buffer_11895_1 (.in(n11895_0), .out(n11895_1));
wire n11896; //CHANX 4 (4,8) #54
wire n11896_0;
wire n11896_1;
buffer_wire buffer_11896_1 (.in(n11896_0), .out(n11896_1));
wire n11897; //CHANX 4 (4,8) #55
wire n11897_0;
wire n11897_1;
buffer_wire buffer_11897_1 (.in(n11897_0), .out(n11897_1));
wire n11898; //CHANX 4 (4,8) #62
wire n11898_0;
wire n11898_1;
buffer_wire buffer_11898_1 (.in(n11898_0), .out(n11898_1));
wire n11899; //CHANX 4 (4,8) #63
wire n11899_0;
wire n11899_1;
buffer_wire buffer_11899_1 (.in(n11899_0), .out(n11899_1));
wire n11900; //CHANX 4 (4,8) #70
wire n11900_0;
wire n11900_1;
buffer_wire buffer_11900_1 (.in(n11900_0), .out(n11900_1));
wire n11901; //CHANX 4 (4,8) #71
wire n11901_0;
wire n11901_1;
buffer_wire buffer_11901_1 (.in(n11901_0), .out(n11901_1));
wire n11902; //CHANX 4 (4,8) #78
wire n11902_0;
wire n11902_1;
buffer_wire buffer_11902_1 (.in(n11902_0), .out(n11902_1));
wire n11903; //CHANX 4 (4,8) #79
wire n11903_0;
wire n11903_1;
buffer_wire buffer_11903_1 (.in(n11903_0), .out(n11903_1));
wire n11904; //CHANX 6 (4,8) #86
wire n11904_0;
wire n11904_1;
buffer_wire buffer_11904_1 (.in(n11904_0), .out(n11904_1));
wire n11905; //CHANX 6 (4,8) #87
wire n11905_0;
wire n11905_1;
buffer_wire buffer_11905_1 (.in(n11905_0), .out(n11905_1));
wire n11906; //CHANX 4 (5,8) #0
wire n11906_0;
wire n11906_1;
buffer_wire buffer_11906_1 (.in(n11906_0), .out(n11906_1));
wire n11907; //CHANX 4 (5,8) #1
wire n11907_0;
wire n11907_1;
buffer_wire buffer_11907_1 (.in(n11907_0), .out(n11907_1));
wire n11908; //CHANX 4 (5,8) #8
wire n11908_0;
wire n11908_1;
buffer_wire buffer_11908_1 (.in(n11908_0), .out(n11908_1));
wire n11909; //CHANX 4 (5,8) #9
wire n11909_0;
wire n11909_1;
buffer_wire buffer_11909_1 (.in(n11909_0), .out(n11909_1));
wire n11910; //CHANX 4 (5,8) #16
wire n11910_0;
wire n11910_1;
buffer_wire buffer_11910_1 (.in(n11910_0), .out(n11910_1));
wire n11911; //CHANX 4 (5,8) #17
wire n11911_0;
wire n11911_1;
buffer_wire buffer_11911_1 (.in(n11911_0), .out(n11911_1));
wire n11912; //CHANX 4 (5,8) #24
wire n11912_0;
wire n11912_1;
buffer_wire buffer_11912_1 (.in(n11912_0), .out(n11912_1));
wire n11913; //CHANX 4 (5,8) #25
wire n11913_0;
wire n11913_1;
buffer_wire buffer_11913_1 (.in(n11913_0), .out(n11913_1));
wire n11914; //CHANX 4 (5,8) #32
wire n11914_0;
wire n11914_1;
buffer_wire buffer_11914_1 (.in(n11914_0), .out(n11914_1));
wire n11915; //CHANX 4 (5,8) #33
wire n11915_0;
wire n11915_1;
buffer_wire buffer_11915_1 (.in(n11915_0), .out(n11915_1));
wire n11916; //CHANX 4 (5,8) #40
wire n11916_0;
wire n11916_1;
buffer_wire buffer_11916_1 (.in(n11916_0), .out(n11916_1));
wire n11917; //CHANX 4 (5,8) #41
wire n11917_0;
wire n11917_1;
buffer_wire buffer_11917_1 (.in(n11917_0), .out(n11917_1));
wire n11918; //CHANX 4 (5,8) #48
wire n11918_0;
wire n11918_1;
buffer_wire buffer_11918_1 (.in(n11918_0), .out(n11918_1));
wire n11919; //CHANX 4 (5,8) #49
wire n11919_0;
wire n11919_1;
buffer_wire buffer_11919_1 (.in(n11919_0), .out(n11919_1));
wire n11920; //CHANX 4 (5,8) #56
wire n11920_0;
wire n11920_1;
buffer_wire buffer_11920_1 (.in(n11920_0), .out(n11920_1));
wire n11921; //CHANX 4 (5,8) #57
wire n11921_0;
wire n11921_1;
buffer_wire buffer_11921_1 (.in(n11921_0), .out(n11921_1));
wire n11922; //CHANX 4 (5,8) #64
wire n11922_0;
wire n11922_1;
buffer_wire buffer_11922_1 (.in(n11922_0), .out(n11922_1));
wire n11923; //CHANX 4 (5,8) #65
wire n11923_0;
wire n11923_1;
buffer_wire buffer_11923_1 (.in(n11923_0), .out(n11923_1));
wire n11924; //CHANX 4 (5,8) #72
wire n11924_0;
wire n11924_1;
buffer_wire buffer_11924_1 (.in(n11924_0), .out(n11924_1));
wire n11925; //CHANX 4 (5,8) #73
wire n11925_0;
wire n11925_1;
buffer_wire buffer_11925_1 (.in(n11925_0), .out(n11925_1));
wire n11926; //CHANX 5 (5,8) #88
wire n11926_0;
wire n11926_1;
buffer_wire buffer_11926_1 (.in(n11926_0), .out(n11926_1));
wire n11927; //CHANX 5 (5,8) #89
wire n11927_0;
wire n11927_1;
buffer_wire buffer_11927_1 (.in(n11927_0), .out(n11927_1));
wire n11928; //CHANX 4 (6,8) #2
wire n11928_0;
wire n11928_1;
buffer_wire buffer_11928_1 (.in(n11928_0), .out(n11928_1));
wire n11929; //CHANX 4 (6,8) #3
wire n11929_0;
wire n11929_1;
buffer_wire buffer_11929_1 (.in(n11929_0), .out(n11929_1));
wire n11930; //CHANX 4 (6,8) #10
wire n11930_0;
wire n11930_1;
buffer_wire buffer_11930_1 (.in(n11930_0), .out(n11930_1));
wire n11931; //CHANX 4 (6,8) #11
wire n11931_0;
wire n11931_1;
buffer_wire buffer_11931_1 (.in(n11931_0), .out(n11931_1));
wire n11932; //CHANX 4 (6,8) #18
wire n11932_0;
wire n11932_1;
buffer_wire buffer_11932_1 (.in(n11932_0), .out(n11932_1));
wire n11933; //CHANX 4 (6,8) #19
wire n11933_0;
wire n11933_1;
buffer_wire buffer_11933_1 (.in(n11933_0), .out(n11933_1));
wire n11934; //CHANX 4 (6,8) #26
wire n11934_0;
wire n11934_1;
buffer_wire buffer_11934_1 (.in(n11934_0), .out(n11934_1));
wire n11935; //CHANX 4 (6,8) #27
wire n11935_0;
wire n11935_1;
buffer_wire buffer_11935_1 (.in(n11935_0), .out(n11935_1));
wire n11936; //CHANX 4 (6,8) #34
wire n11936_0;
wire n11936_1;
buffer_wire buffer_11936_1 (.in(n11936_0), .out(n11936_1));
wire n11937; //CHANX 4 (6,8) #35
wire n11937_0;
wire n11937_1;
buffer_wire buffer_11937_1 (.in(n11937_0), .out(n11937_1));
wire n11938; //CHANX 4 (6,8) #42
wire n11938_0;
wire n11938_1;
buffer_wire buffer_11938_1 (.in(n11938_0), .out(n11938_1));
wire n11939; //CHANX 4 (6,8) #43
wire n11939_0;
wire n11939_1;
buffer_wire buffer_11939_1 (.in(n11939_0), .out(n11939_1));
wire n11940; //CHANX 4 (6,8) #50
wire n11940_0;
wire n11940_1;
buffer_wire buffer_11940_1 (.in(n11940_0), .out(n11940_1));
wire n11941; //CHANX 4 (6,8) #51
wire n11941_0;
wire n11941_1;
buffer_wire buffer_11941_1 (.in(n11941_0), .out(n11941_1));
wire n11942; //CHANX 4 (6,8) #58
wire n11942_0;
wire n11942_1;
buffer_wire buffer_11942_1 (.in(n11942_0), .out(n11942_1));
wire n11943; //CHANX 4 (6,8) #59
wire n11943_0;
wire n11943_1;
buffer_wire buffer_11943_1 (.in(n11943_0), .out(n11943_1));
wire n11944; //CHANX 4 (6,8) #66
wire n11944_0;
wire n11944_1;
buffer_wire buffer_11944_1 (.in(n11944_0), .out(n11944_1));
wire n11945; //CHANX 4 (6,8) #67
wire n11945_0;
wire n11945_1;
buffer_wire buffer_11945_1 (.in(n11945_0), .out(n11945_1));
wire n11946; //CHANX 4 (6,8) #74
wire n11946_0;
wire n11946_1;
buffer_wire buffer_11946_1 (.in(n11946_0), .out(n11946_1));
wire n11947; //CHANX 4 (6,8) #75
wire n11947_0;
wire n11947_1;
buffer_wire buffer_11947_1 (.in(n11947_0), .out(n11947_1));
wire n11948; //CHANX 4 (6,8) #90
wire n11948_0;
wire n11948_1;
buffer_wire buffer_11948_1 (.in(n11948_0), .out(n11948_1));
wire n11949; //CHANX 4 (6,8) #91
wire n11949_0;
wire n11949_1;
buffer_wire buffer_11949_1 (.in(n11949_0), .out(n11949_1));
wire n11950; //CHANX 3 (7,8) #4
wire n11950_0;
wire n11951; //CHANX 3 (7,8) #5
wire n11951_0;
wire n11952; //CHANX 3 (7,8) #12
wire n11952_0;
wire n11953; //CHANX 3 (7,8) #13
wire n11953_0;
wire n11954; //CHANX 3 (7,8) #20
wire n11954_0;
wire n11955; //CHANX 3 (7,8) #21
wire n11955_0;
wire n11956; //CHANX 3 (7,8) #28
wire n11956_0;
wire n11957; //CHANX 3 (7,8) #29
wire n11957_0;
wire n11958; //CHANX 3 (7,8) #36
wire n11958_0;
wire n11959; //CHANX 3 (7,8) #37
wire n11959_0;
wire n11960; //CHANX 3 (7,8) #44
wire n11960_0;
wire n11961; //CHANX 3 (7,8) #45
wire n11961_0;
wire n11962; //CHANX 3 (7,8) #52
wire n11962_0;
wire n11963; //CHANX 3 (7,8) #53
wire n11963_0;
wire n11964; //CHANX 3 (7,8) #60
wire n11964_0;
wire n11965; //CHANX 3 (7,8) #61
wire n11965_0;
wire n11966; //CHANX 3 (7,8) #68
wire n11966_0;
wire n11967; //CHANX 3 (7,8) #69
wire n11967_0;
wire n11968; //CHANX 3 (7,8) #76
wire n11968_0;
wire n11969; //CHANX 3 (7,8) #77
wire n11969_0;
wire n11970; //CHANX 2 (8,8) #6
wire n11970_0;
wire n11971; //CHANX 2 (8,8) #7
wire n11971_0;
wire n11972; //CHANX 2 (8,8) #14
wire n11972_0;
wire n11973; //CHANX 2 (8,8) #15
wire n11973_0;
wire n11974; //CHANX 2 (8,8) #22
wire n11974_0;
wire n11975; //CHANX 2 (8,8) #23
wire n11975_0;
wire n11976; //CHANX 2 (8,8) #30
wire n11976_0;
wire n11977; //CHANX 2 (8,8) #31
wire n11977_0;
wire n11978; //CHANX 2 (8,8) #38
wire n11978_0;
wire n11979; //CHANX 2 (8,8) #39
wire n11979_0;
wire n11980; //CHANX 2 (8,8) #46
wire n11980_0;
wire n11981; //CHANX 2 (8,8) #47
wire n11981_0;
wire n11982; //CHANX 2 (8,8) #54
wire n11982_0;
wire n11983; //CHANX 2 (8,8) #55
wire n11983_0;
wire n11984; //CHANX 2 (8,8) #62
wire n11984_0;
wire n11985; //CHANX 2 (8,8) #63
wire n11985_0;
wire n11986; //CHANX 2 (8,8) #70
wire n11986_0;
wire n11987; //CHANX 2 (8,8) #71
wire n11987_0;
wire n11988; //CHANX 2 (8,8) #78
wire n11988_0;
wire n11989; //CHANX 2 (8,8) #79
wire n11989_0;
wire n11990; //CHANX 1 (9,8) #0
wire n11990_0;
wire n11991; //CHANX 1 (9,8) #1
wire n11991_0;
wire n11992; //CHANX 1 (9,8) #8
wire n11992_0;
wire n11993; //CHANX 1 (9,8) #9
wire n11993_0;
wire n11994; //CHANX 1 (9,8) #16
wire n11994_0;
wire n11995; //CHANX 1 (9,8) #17
wire n11995_0;
wire n11996; //CHANX 1 (9,8) #24
wire n11996_0;
wire n11997; //CHANX 1 (9,8) #25
wire n11997_0;
wire n11998; //CHANX 1 (9,8) #32
wire n11998_0;
wire n11999; //CHANX 1 (9,8) #33
wire n11999_0;
wire n12000; //CHANX 1 (9,8) #40
wire n12000_0;
wire n12001; //CHANX 1 (9,8) #41
wire n12001_0;
wire n12002; //CHANX 1 (9,8) #48
wire n12002_0;
wire n12003; //CHANX 1 (9,8) #49
wire n12003_0;
wire n12004; //CHANX 1 (9,8) #56
wire n12004_0;
wire n12005; //CHANX 1 (9,8) #57
wire n12005_0;
wire n12006; //CHANX 1 (9,8) #64
wire n12006_0;
wire n12007; //CHANX 1 (9,8) #65
wire n12007_0;
wire n12008; //CHANX 1 (9,8) #72
wire n12008_0;
wire n12009; //CHANX 1 (9,8) #73
wire n12009_0;
wire n12010; //CHANX 3 (1,9) #0
wire n12010_0;
wire n12011; //CHANX 3 (1,9) #1
wire n12011_0;
wire n12012; //CHANX 4 (1,9) #2
wire n12012_0;
wire n12012_1;
buffer_wire buffer_12012_1 (.in(n12012_0), .out(n12012_1));
wire n12013; //CHANX 4 (1,9) #3
wire n12013_0;
wire n12013_1;
buffer_wire buffer_12013_1 (.in(n12013_0), .out(n12013_1));
wire n12014; //CHANX 1 (1,9) #4
wire n12014_0;
wire n12015; //CHANX 1 (1,9) #5
wire n12015_0;
wire n12016; //CHANX 2 (1,9) #6
wire n12016_0;
wire n12017; //CHANX 2 (1,9) #7
wire n12017_0;
wire n12018; //CHANX 3 (1,9) #8
wire n12018_0;
wire n12019; //CHANX 3 (1,9) #9
wire n12019_0;
wire n12020; //CHANX 4 (1,9) #10
wire n12020_0;
wire n12020_1;
buffer_wire buffer_12020_1 (.in(n12020_0), .out(n12020_1));
wire n12021; //CHANX 4 (1,9) #11
wire n12021_0;
wire n12021_1;
buffer_wire buffer_12021_1 (.in(n12021_0), .out(n12021_1));
wire n12022; //CHANX 1 (1,9) #12
wire n12022_0;
wire n12023; //CHANX 1 (1,9) #13
wire n12023_0;
wire n12024; //CHANX 2 (1,9) #14
wire n12024_0;
wire n12025; //CHANX 2 (1,9) #15
wire n12025_0;
wire n12026; //CHANX 3 (1,9) #16
wire n12026_0;
wire n12027; //CHANX 3 (1,9) #17
wire n12027_0;
wire n12028; //CHANX 4 (1,9) #18
wire n12028_0;
wire n12028_1;
buffer_wire buffer_12028_1 (.in(n12028_0), .out(n12028_1));
wire n12029; //CHANX 4 (1,9) #19
wire n12029_0;
wire n12029_1;
buffer_wire buffer_12029_1 (.in(n12029_0), .out(n12029_1));
wire n12030; //CHANX 1 (1,9) #20
wire n12030_0;
wire n12031; //CHANX 1 (1,9) #21
wire n12031_0;
wire n12032; //CHANX 2 (1,9) #22
wire n12032_0;
wire n12033; //CHANX 2 (1,9) #23
wire n12033_0;
wire n12034; //CHANX 3 (1,9) #24
wire n12034_0;
wire n12035; //CHANX 3 (1,9) #25
wire n12035_0;
wire n12036; //CHANX 4 (1,9) #26
wire n12036_0;
wire n12036_1;
buffer_wire buffer_12036_1 (.in(n12036_0), .out(n12036_1));
wire n12037; //CHANX 4 (1,9) #27
wire n12037_0;
wire n12037_1;
buffer_wire buffer_12037_1 (.in(n12037_0), .out(n12037_1));
wire n12038; //CHANX 1 (1,9) #28
wire n12038_0;
wire n12039; //CHANX 1 (1,9) #29
wire n12039_0;
wire n12040; //CHANX 2 (1,9) #30
wire n12040_0;
wire n12041; //CHANX 2 (1,9) #31
wire n12041_0;
wire n12042; //CHANX 3 (1,9) #32
wire n12042_0;
wire n12043; //CHANX 3 (1,9) #33
wire n12043_0;
wire n12044; //CHANX 4 (1,9) #34
wire n12044_0;
wire n12044_1;
buffer_wire buffer_12044_1 (.in(n12044_0), .out(n12044_1));
wire n12045; //CHANX 4 (1,9) #35
wire n12045_0;
wire n12045_1;
buffer_wire buffer_12045_1 (.in(n12045_0), .out(n12045_1));
wire n12046; //CHANX 1 (1,9) #36
wire n12046_0;
wire n12047; //CHANX 1 (1,9) #37
wire n12047_0;
wire n12048; //CHANX 2 (1,9) #38
wire n12048_0;
wire n12049; //CHANX 2 (1,9) #39
wire n12049_0;
wire n12050; //CHANX 3 (1,9) #40
wire n12050_0;
wire n12051; //CHANX 3 (1,9) #41
wire n12051_0;
wire n12052; //CHANX 4 (1,9) #42
wire n12052_0;
wire n12052_1;
buffer_wire buffer_12052_1 (.in(n12052_0), .out(n12052_1));
wire n12053; //CHANX 4 (1,9) #43
wire n12053_0;
wire n12053_1;
buffer_wire buffer_12053_1 (.in(n12053_0), .out(n12053_1));
wire n12054; //CHANX 1 (1,9) #44
wire n12054_0;
wire n12055; //CHANX 1 (1,9) #45
wire n12055_0;
wire n12056; //CHANX 2 (1,9) #46
wire n12056_0;
wire n12057; //CHANX 2 (1,9) #47
wire n12057_0;
wire n12058; //CHANX 3 (1,9) #48
wire n12058_0;
wire n12059; //CHANX 3 (1,9) #49
wire n12059_0;
wire n12060; //CHANX 4 (1,9) #50
wire n12060_0;
wire n12060_1;
buffer_wire buffer_12060_1 (.in(n12060_0), .out(n12060_1));
wire n12061; //CHANX 4 (1,9) #51
wire n12061_0;
wire n12061_1;
buffer_wire buffer_12061_1 (.in(n12061_0), .out(n12061_1));
wire n12062; //CHANX 1 (1,9) #52
wire n12062_0;
wire n12063; //CHANX 1 (1,9) #53
wire n12063_0;
wire n12064; //CHANX 2 (1,9) #54
wire n12064_0;
wire n12065; //CHANX 2 (1,9) #55
wire n12065_0;
wire n12066; //CHANX 3 (1,9) #56
wire n12066_0;
wire n12067; //CHANX 3 (1,9) #57
wire n12067_0;
wire n12068; //CHANX 4 (1,9) #58
wire n12068_0;
wire n12068_1;
buffer_wire buffer_12068_1 (.in(n12068_0), .out(n12068_1));
wire n12069; //CHANX 4 (1,9) #59
wire n12069_0;
wire n12069_1;
buffer_wire buffer_12069_1 (.in(n12069_0), .out(n12069_1));
wire n12070; //CHANX 1 (1,9) #60
wire n12070_0;
wire n12071; //CHANX 1 (1,9) #61
wire n12071_0;
wire n12072; //CHANX 2 (1,9) #62
wire n12072_0;
wire n12073; //CHANX 2 (1,9) #63
wire n12073_0;
wire n12074; //CHANX 3 (1,9) #64
wire n12074_0;
wire n12075; //CHANX 3 (1,9) #65
wire n12075_0;
wire n12076; //CHANX 4 (1,9) #66
wire n12076_0;
wire n12076_1;
buffer_wire buffer_12076_1 (.in(n12076_0), .out(n12076_1));
wire n12077; //CHANX 4 (1,9) #67
wire n12077_0;
wire n12077_1;
buffer_wire buffer_12077_1 (.in(n12077_0), .out(n12077_1));
wire n12078; //CHANX 1 (1,9) #68
wire n12078_0;
wire n12079; //CHANX 1 (1,9) #69
wire n12079_0;
wire n12080; //CHANX 2 (1,9) #70
wire n12080_0;
wire n12081; //CHANX 2 (1,9) #71
wire n12081_0;
wire n12082; //CHANX 3 (1,9) #72
wire n12082_0;
wire n12083; //CHANX 3 (1,9) #73
wire n12083_0;
wire n12084; //CHANX 4 (1,9) #74
wire n12084_0;
wire n12084_1;
buffer_wire buffer_12084_1 (.in(n12084_0), .out(n12084_1));
wire n12085; //CHANX 4 (1,9) #75
wire n12085_0;
wire n12085_1;
buffer_wire buffer_12085_1 (.in(n12085_0), .out(n12085_1));
wire n12086; //CHANX 1 (1,9) #76
wire n12086_0;
wire n12087; //CHANX 1 (1,9) #77
wire n12087_0;
wire n12088; //CHANX 2 (1,9) #78
wire n12088_0;
wire n12089; //CHANX 2 (1,9) #79
wire n12089_0;
wire n12090; //CHANX 9 (1,9) #80
wire n12090_0;
wire n12090_1;
wire n12090_2;
buffer_wire buffer_12090_2 (.in(n12090_1), .out(n12090_2));
buffer_wire buffer_12090_1 (.in(n12090_0), .out(n12090_1));
wire n12091; //CHANX 9 (1,9) #81
wire n12091_0;
wire n12091_1;
wire n12091_2;
buffer_wire buffer_12091_2 (.in(n12091_1), .out(n12091_2));
buffer_wire buffer_12091_1 (.in(n12091_0), .out(n12091_1));
wire n12092; //CHANX 9 (1,9) #82
wire n12092_0;
wire n12092_1;
wire n12092_2;
buffer_wire buffer_12092_2 (.in(n12092_1), .out(n12092_2));
buffer_wire buffer_12092_1 (.in(n12092_0), .out(n12092_1));
wire n12093; //CHANX 9 (1,9) #83
wire n12093_0;
wire n12093_1;
wire n12093_2;
buffer_wire buffer_12093_2 (.in(n12093_1), .out(n12093_2));
buffer_wire buffer_12093_1 (.in(n12093_0), .out(n12093_1));
wire n12094; //CHANX 1 (1,9) #84
wire n12094_0;
wire n12095; //CHANX 1 (1,9) #85
wire n12095_0;
wire n12096; //CHANX 2 (1,9) #86
wire n12096_0;
wire n12097; //CHANX 2 (1,9) #87
wire n12097_0;
wire n12098; //CHANX 3 (1,9) #88
wire n12098_0;
wire n12099; //CHANX 3 (1,9) #89
wire n12099_0;
wire n12100; //CHANX 4 (1,9) #90
wire n12100_0;
wire n12100_1;
buffer_wire buffer_12100_1 (.in(n12100_0), .out(n12100_1));
wire n12101; //CHANX 4 (1,9) #91
wire n12101_0;
wire n12101_1;
buffer_wire buffer_12101_1 (.in(n12101_0), .out(n12101_1));
wire n12102; //CHANX 4 (2,9) #4
wire n12102_0;
wire n12102_1;
buffer_wire buffer_12102_1 (.in(n12102_0), .out(n12102_1));
wire n12103; //CHANX 4 (2,9) #5
wire n12103_0;
wire n12103_1;
buffer_wire buffer_12103_1 (.in(n12103_0), .out(n12103_1));
wire n12104; //CHANX 4 (2,9) #12
wire n12104_0;
wire n12104_1;
buffer_wire buffer_12104_1 (.in(n12104_0), .out(n12104_1));
wire n12105; //CHANX 4 (2,9) #13
wire n12105_0;
wire n12105_1;
buffer_wire buffer_12105_1 (.in(n12105_0), .out(n12105_1));
wire n12106; //CHANX 4 (2,9) #20
wire n12106_0;
wire n12106_1;
buffer_wire buffer_12106_1 (.in(n12106_0), .out(n12106_1));
wire n12107; //CHANX 4 (2,9) #21
wire n12107_0;
wire n12107_1;
buffer_wire buffer_12107_1 (.in(n12107_0), .out(n12107_1));
wire n12108; //CHANX 4 (2,9) #28
wire n12108_0;
wire n12108_1;
buffer_wire buffer_12108_1 (.in(n12108_0), .out(n12108_1));
wire n12109; //CHANX 4 (2,9) #29
wire n12109_0;
wire n12109_1;
buffer_wire buffer_12109_1 (.in(n12109_0), .out(n12109_1));
wire n12110; //CHANX 4 (2,9) #36
wire n12110_0;
wire n12110_1;
buffer_wire buffer_12110_1 (.in(n12110_0), .out(n12110_1));
wire n12111; //CHANX 4 (2,9) #37
wire n12111_0;
wire n12111_1;
buffer_wire buffer_12111_1 (.in(n12111_0), .out(n12111_1));
wire n12112; //CHANX 4 (2,9) #44
wire n12112_0;
wire n12112_1;
buffer_wire buffer_12112_1 (.in(n12112_0), .out(n12112_1));
wire n12113; //CHANX 4 (2,9) #45
wire n12113_0;
wire n12113_1;
buffer_wire buffer_12113_1 (.in(n12113_0), .out(n12113_1));
wire n12114; //CHANX 4 (2,9) #52
wire n12114_0;
wire n12114_1;
buffer_wire buffer_12114_1 (.in(n12114_0), .out(n12114_1));
wire n12115; //CHANX 4 (2,9) #53
wire n12115_0;
wire n12115_1;
buffer_wire buffer_12115_1 (.in(n12115_0), .out(n12115_1));
wire n12116; //CHANX 4 (2,9) #60
wire n12116_0;
wire n12116_1;
buffer_wire buffer_12116_1 (.in(n12116_0), .out(n12116_1));
wire n12117; //CHANX 4 (2,9) #61
wire n12117_0;
wire n12117_1;
buffer_wire buffer_12117_1 (.in(n12117_0), .out(n12117_1));
wire n12118; //CHANX 4 (2,9) #68
wire n12118_0;
wire n12118_1;
buffer_wire buffer_12118_1 (.in(n12118_0), .out(n12118_1));
wire n12119; //CHANX 4 (2,9) #69
wire n12119_0;
wire n12119_1;
buffer_wire buffer_12119_1 (.in(n12119_0), .out(n12119_1));
wire n12120; //CHANX 4 (2,9) #76
wire n12120_0;
wire n12120_1;
buffer_wire buffer_12120_1 (.in(n12120_0), .out(n12120_1));
wire n12121; //CHANX 4 (2,9) #77
wire n12121_0;
wire n12121_1;
buffer_wire buffer_12121_1 (.in(n12121_0), .out(n12121_1));
wire n12122; //CHANX 8 (2,9) #84
wire n12122_0;
wire n12122_1;
wire n12122_2;
buffer_wire buffer_12122_2 (.in(n12122_1), .out(n12122_2));
buffer_wire buffer_12122_1 (.in(n12122_0), .out(n12122_1));
wire n12123; //CHANX 8 (2,9) #85
wire n12123_0;
wire n12123_1;
wire n12123_2;
buffer_wire buffer_12123_2 (.in(n12123_1), .out(n12123_2));
buffer_wire buffer_12123_1 (.in(n12123_0), .out(n12123_1));
wire n12124; //CHANX 4 (3,9) #6
wire n12124_0;
wire n12124_1;
buffer_wire buffer_12124_1 (.in(n12124_0), .out(n12124_1));
wire n12125; //CHANX 4 (3,9) #7
wire n12125_0;
wire n12125_1;
buffer_wire buffer_12125_1 (.in(n12125_0), .out(n12125_1));
wire n12126; //CHANX 4 (3,9) #14
wire n12126_0;
wire n12126_1;
buffer_wire buffer_12126_1 (.in(n12126_0), .out(n12126_1));
wire n12127; //CHANX 4 (3,9) #15
wire n12127_0;
wire n12127_1;
buffer_wire buffer_12127_1 (.in(n12127_0), .out(n12127_1));
wire n12128; //CHANX 4 (3,9) #22
wire n12128_0;
wire n12128_1;
buffer_wire buffer_12128_1 (.in(n12128_0), .out(n12128_1));
wire n12129; //CHANX 4 (3,9) #23
wire n12129_0;
wire n12129_1;
buffer_wire buffer_12129_1 (.in(n12129_0), .out(n12129_1));
wire n12130; //CHANX 4 (3,9) #30
wire n12130_0;
wire n12130_1;
buffer_wire buffer_12130_1 (.in(n12130_0), .out(n12130_1));
wire n12131; //CHANX 4 (3,9) #31
wire n12131_0;
wire n12131_1;
buffer_wire buffer_12131_1 (.in(n12131_0), .out(n12131_1));
wire n12132; //CHANX 4 (3,9) #38
wire n12132_0;
wire n12132_1;
buffer_wire buffer_12132_1 (.in(n12132_0), .out(n12132_1));
wire n12133; //CHANX 4 (3,9) #39
wire n12133_0;
wire n12133_1;
buffer_wire buffer_12133_1 (.in(n12133_0), .out(n12133_1));
wire n12134; //CHANX 4 (3,9) #46
wire n12134_0;
wire n12134_1;
buffer_wire buffer_12134_1 (.in(n12134_0), .out(n12134_1));
wire n12135; //CHANX 4 (3,9) #47
wire n12135_0;
wire n12135_1;
buffer_wire buffer_12135_1 (.in(n12135_0), .out(n12135_1));
wire n12136; //CHANX 4 (3,9) #54
wire n12136_0;
wire n12136_1;
buffer_wire buffer_12136_1 (.in(n12136_0), .out(n12136_1));
wire n12137; //CHANX 4 (3,9) #55
wire n12137_0;
wire n12137_1;
buffer_wire buffer_12137_1 (.in(n12137_0), .out(n12137_1));
wire n12138; //CHANX 4 (3,9) #62
wire n12138_0;
wire n12138_1;
buffer_wire buffer_12138_1 (.in(n12138_0), .out(n12138_1));
wire n12139; //CHANX 4 (3,9) #63
wire n12139_0;
wire n12139_1;
buffer_wire buffer_12139_1 (.in(n12139_0), .out(n12139_1));
wire n12140; //CHANX 4 (3,9) #70
wire n12140_0;
wire n12140_1;
buffer_wire buffer_12140_1 (.in(n12140_0), .out(n12140_1));
wire n12141; //CHANX 4 (3,9) #71
wire n12141_0;
wire n12141_1;
buffer_wire buffer_12141_1 (.in(n12141_0), .out(n12141_1));
wire n12142; //CHANX 4 (3,9) #78
wire n12142_0;
wire n12142_1;
buffer_wire buffer_12142_1 (.in(n12142_0), .out(n12142_1));
wire n12143; //CHANX 4 (3,9) #79
wire n12143_0;
wire n12143_1;
buffer_wire buffer_12143_1 (.in(n12143_0), .out(n12143_1));
wire n12144; //CHANX 7 (3,9) #86
wire n12144_0;
wire n12144_1;
wire n12144_2;
buffer_wire buffer_12144_2 (.in(n12144_1), .out(n12144_2));
buffer_wire buffer_12144_1 (.in(n12144_0), .out(n12144_1));
wire n12145; //CHANX 7 (3,9) #87
wire n12145_0;
wire n12145_1;
wire n12145_2;
buffer_wire buffer_12145_2 (.in(n12145_1), .out(n12145_2));
buffer_wire buffer_12145_1 (.in(n12145_0), .out(n12145_1));
wire n12146; //CHANX 4 (4,9) #0
wire n12146_0;
wire n12146_1;
buffer_wire buffer_12146_1 (.in(n12146_0), .out(n12146_1));
wire n12147; //CHANX 4 (4,9) #1
wire n12147_0;
wire n12147_1;
buffer_wire buffer_12147_1 (.in(n12147_0), .out(n12147_1));
wire n12148; //CHANX 4 (4,9) #8
wire n12148_0;
wire n12148_1;
buffer_wire buffer_12148_1 (.in(n12148_0), .out(n12148_1));
wire n12149; //CHANX 4 (4,9) #9
wire n12149_0;
wire n12149_1;
buffer_wire buffer_12149_1 (.in(n12149_0), .out(n12149_1));
wire n12150; //CHANX 4 (4,9) #16
wire n12150_0;
wire n12150_1;
buffer_wire buffer_12150_1 (.in(n12150_0), .out(n12150_1));
wire n12151; //CHANX 4 (4,9) #17
wire n12151_0;
wire n12151_1;
buffer_wire buffer_12151_1 (.in(n12151_0), .out(n12151_1));
wire n12152; //CHANX 4 (4,9) #24
wire n12152_0;
wire n12152_1;
buffer_wire buffer_12152_1 (.in(n12152_0), .out(n12152_1));
wire n12153; //CHANX 4 (4,9) #25
wire n12153_0;
wire n12153_1;
buffer_wire buffer_12153_1 (.in(n12153_0), .out(n12153_1));
wire n12154; //CHANX 4 (4,9) #32
wire n12154_0;
wire n12154_1;
buffer_wire buffer_12154_1 (.in(n12154_0), .out(n12154_1));
wire n12155; //CHANX 4 (4,9) #33
wire n12155_0;
wire n12155_1;
buffer_wire buffer_12155_1 (.in(n12155_0), .out(n12155_1));
wire n12156; //CHANX 4 (4,9) #40
wire n12156_0;
wire n12156_1;
buffer_wire buffer_12156_1 (.in(n12156_0), .out(n12156_1));
wire n12157; //CHANX 4 (4,9) #41
wire n12157_0;
wire n12157_1;
buffer_wire buffer_12157_1 (.in(n12157_0), .out(n12157_1));
wire n12158; //CHANX 4 (4,9) #48
wire n12158_0;
wire n12158_1;
buffer_wire buffer_12158_1 (.in(n12158_0), .out(n12158_1));
wire n12159; //CHANX 4 (4,9) #49
wire n12159_0;
wire n12159_1;
buffer_wire buffer_12159_1 (.in(n12159_0), .out(n12159_1));
wire n12160; //CHANX 4 (4,9) #56
wire n12160_0;
wire n12160_1;
buffer_wire buffer_12160_1 (.in(n12160_0), .out(n12160_1));
wire n12161; //CHANX 4 (4,9) #57
wire n12161_0;
wire n12161_1;
buffer_wire buffer_12161_1 (.in(n12161_0), .out(n12161_1));
wire n12162; //CHANX 4 (4,9) #64
wire n12162_0;
wire n12162_1;
buffer_wire buffer_12162_1 (.in(n12162_0), .out(n12162_1));
wire n12163; //CHANX 4 (4,9) #65
wire n12163_0;
wire n12163_1;
buffer_wire buffer_12163_1 (.in(n12163_0), .out(n12163_1));
wire n12164; //CHANX 4 (4,9) #72
wire n12164_0;
wire n12164_1;
buffer_wire buffer_12164_1 (.in(n12164_0), .out(n12164_1));
wire n12165; //CHANX 4 (4,9) #73
wire n12165_0;
wire n12165_1;
buffer_wire buffer_12165_1 (.in(n12165_0), .out(n12165_1));
wire n12166; //CHANX 6 (4,9) #88
wire n12166_0;
wire n12166_1;
buffer_wire buffer_12166_1 (.in(n12166_0), .out(n12166_1));
wire n12167; //CHANX 6 (4,9) #89
wire n12167_0;
wire n12167_1;
buffer_wire buffer_12167_1 (.in(n12167_0), .out(n12167_1));
wire n12168; //CHANX 4 (5,9) #2
wire n12168_0;
wire n12168_1;
buffer_wire buffer_12168_1 (.in(n12168_0), .out(n12168_1));
wire n12169; //CHANX 4 (5,9) #3
wire n12169_0;
wire n12169_1;
buffer_wire buffer_12169_1 (.in(n12169_0), .out(n12169_1));
wire n12170; //CHANX 4 (5,9) #10
wire n12170_0;
wire n12170_1;
buffer_wire buffer_12170_1 (.in(n12170_0), .out(n12170_1));
wire n12171; //CHANX 4 (5,9) #11
wire n12171_0;
wire n12171_1;
buffer_wire buffer_12171_1 (.in(n12171_0), .out(n12171_1));
wire n12172; //CHANX 4 (5,9) #18
wire n12172_0;
wire n12172_1;
buffer_wire buffer_12172_1 (.in(n12172_0), .out(n12172_1));
wire n12173; //CHANX 4 (5,9) #19
wire n12173_0;
wire n12173_1;
buffer_wire buffer_12173_1 (.in(n12173_0), .out(n12173_1));
wire n12174; //CHANX 4 (5,9) #26
wire n12174_0;
wire n12174_1;
buffer_wire buffer_12174_1 (.in(n12174_0), .out(n12174_1));
wire n12175; //CHANX 4 (5,9) #27
wire n12175_0;
wire n12175_1;
buffer_wire buffer_12175_1 (.in(n12175_0), .out(n12175_1));
wire n12176; //CHANX 4 (5,9) #34
wire n12176_0;
wire n12176_1;
buffer_wire buffer_12176_1 (.in(n12176_0), .out(n12176_1));
wire n12177; //CHANX 4 (5,9) #35
wire n12177_0;
wire n12177_1;
buffer_wire buffer_12177_1 (.in(n12177_0), .out(n12177_1));
wire n12178; //CHANX 4 (5,9) #42
wire n12178_0;
wire n12178_1;
buffer_wire buffer_12178_1 (.in(n12178_0), .out(n12178_1));
wire n12179; //CHANX 4 (5,9) #43
wire n12179_0;
wire n12179_1;
buffer_wire buffer_12179_1 (.in(n12179_0), .out(n12179_1));
wire n12180; //CHANX 4 (5,9) #50
wire n12180_0;
wire n12180_1;
buffer_wire buffer_12180_1 (.in(n12180_0), .out(n12180_1));
wire n12181; //CHANX 4 (5,9) #51
wire n12181_0;
wire n12181_1;
buffer_wire buffer_12181_1 (.in(n12181_0), .out(n12181_1));
wire n12182; //CHANX 4 (5,9) #58
wire n12182_0;
wire n12182_1;
buffer_wire buffer_12182_1 (.in(n12182_0), .out(n12182_1));
wire n12183; //CHANX 4 (5,9) #59
wire n12183_0;
wire n12183_1;
buffer_wire buffer_12183_1 (.in(n12183_0), .out(n12183_1));
wire n12184; //CHANX 4 (5,9) #66
wire n12184_0;
wire n12184_1;
buffer_wire buffer_12184_1 (.in(n12184_0), .out(n12184_1));
wire n12185; //CHANX 4 (5,9) #67
wire n12185_0;
wire n12185_1;
buffer_wire buffer_12185_1 (.in(n12185_0), .out(n12185_1));
wire n12186; //CHANX 4 (5,9) #74
wire n12186_0;
wire n12186_1;
buffer_wire buffer_12186_1 (.in(n12186_0), .out(n12186_1));
wire n12187; //CHANX 4 (5,9) #75
wire n12187_0;
wire n12187_1;
buffer_wire buffer_12187_1 (.in(n12187_0), .out(n12187_1));
wire n12188; //CHANX 5 (5,9) #90
wire n12188_0;
wire n12188_1;
buffer_wire buffer_12188_1 (.in(n12188_0), .out(n12188_1));
wire n12189; //CHANX 5 (5,9) #91
wire n12189_0;
wire n12189_1;
buffer_wire buffer_12189_1 (.in(n12189_0), .out(n12189_1));
wire n12190; //CHANX 4 (6,9) #4
wire n12190_0;
wire n12190_1;
buffer_wire buffer_12190_1 (.in(n12190_0), .out(n12190_1));
wire n12191; //CHANX 4 (6,9) #5
wire n12191_0;
wire n12191_1;
buffer_wire buffer_12191_1 (.in(n12191_0), .out(n12191_1));
wire n12192; //CHANX 4 (6,9) #12
wire n12192_0;
wire n12192_1;
buffer_wire buffer_12192_1 (.in(n12192_0), .out(n12192_1));
wire n12193; //CHANX 4 (6,9) #13
wire n12193_0;
wire n12193_1;
buffer_wire buffer_12193_1 (.in(n12193_0), .out(n12193_1));
wire n12194; //CHANX 4 (6,9) #20
wire n12194_0;
wire n12194_1;
buffer_wire buffer_12194_1 (.in(n12194_0), .out(n12194_1));
wire n12195; //CHANX 4 (6,9) #21
wire n12195_0;
wire n12195_1;
buffer_wire buffer_12195_1 (.in(n12195_0), .out(n12195_1));
wire n12196; //CHANX 4 (6,9) #28
wire n12196_0;
wire n12196_1;
buffer_wire buffer_12196_1 (.in(n12196_0), .out(n12196_1));
wire n12197; //CHANX 4 (6,9) #29
wire n12197_0;
wire n12197_1;
buffer_wire buffer_12197_1 (.in(n12197_0), .out(n12197_1));
wire n12198; //CHANX 4 (6,9) #36
wire n12198_0;
wire n12198_1;
buffer_wire buffer_12198_1 (.in(n12198_0), .out(n12198_1));
wire n12199; //CHANX 4 (6,9) #37
wire n12199_0;
wire n12199_1;
buffer_wire buffer_12199_1 (.in(n12199_0), .out(n12199_1));
wire n12200; //CHANX 4 (6,9) #44
wire n12200_0;
wire n12200_1;
buffer_wire buffer_12200_1 (.in(n12200_0), .out(n12200_1));
wire n12201; //CHANX 4 (6,9) #45
wire n12201_0;
wire n12201_1;
buffer_wire buffer_12201_1 (.in(n12201_0), .out(n12201_1));
wire n12202; //CHANX 4 (6,9) #52
wire n12202_0;
wire n12202_1;
buffer_wire buffer_12202_1 (.in(n12202_0), .out(n12202_1));
wire n12203; //CHANX 4 (6,9) #53
wire n12203_0;
wire n12203_1;
buffer_wire buffer_12203_1 (.in(n12203_0), .out(n12203_1));
wire n12204; //CHANX 4 (6,9) #60
wire n12204_0;
wire n12204_1;
buffer_wire buffer_12204_1 (.in(n12204_0), .out(n12204_1));
wire n12205; //CHANX 4 (6,9) #61
wire n12205_0;
wire n12205_1;
buffer_wire buffer_12205_1 (.in(n12205_0), .out(n12205_1));
wire n12206; //CHANX 4 (6,9) #68
wire n12206_0;
wire n12206_1;
buffer_wire buffer_12206_1 (.in(n12206_0), .out(n12206_1));
wire n12207; //CHANX 4 (6,9) #69
wire n12207_0;
wire n12207_1;
buffer_wire buffer_12207_1 (.in(n12207_0), .out(n12207_1));
wire n12208; //CHANX 4 (6,9) #76
wire n12208_0;
wire n12208_1;
buffer_wire buffer_12208_1 (.in(n12208_0), .out(n12208_1));
wire n12209; //CHANX 4 (6,9) #77
wire n12209_0;
wire n12209_1;
buffer_wire buffer_12209_1 (.in(n12209_0), .out(n12209_1));
wire n12210; //CHANX 3 (7,9) #6
wire n12210_0;
wire n12211; //CHANX 3 (7,9) #7
wire n12211_0;
wire n12212; //CHANX 3 (7,9) #14
wire n12212_0;
wire n12213; //CHANX 3 (7,9) #15
wire n12213_0;
wire n12214; //CHANX 3 (7,9) #22
wire n12214_0;
wire n12215; //CHANX 3 (7,9) #23
wire n12215_0;
wire n12216; //CHANX 3 (7,9) #30
wire n12216_0;
wire n12217; //CHANX 3 (7,9) #31
wire n12217_0;
wire n12218; //CHANX 3 (7,9) #38
wire n12218_0;
wire n12219; //CHANX 3 (7,9) #39
wire n12219_0;
wire n12220; //CHANX 3 (7,9) #46
wire n12220_0;
wire n12221; //CHANX 3 (7,9) #47
wire n12221_0;
wire n12222; //CHANX 3 (7,9) #54
wire n12222_0;
wire n12223; //CHANX 3 (7,9) #55
wire n12223_0;
wire n12224; //CHANX 3 (7,9) #62
wire n12224_0;
wire n12225; //CHANX 3 (7,9) #63
wire n12225_0;
wire n12226; //CHANX 3 (7,9) #70
wire n12226_0;
wire n12227; //CHANX 3 (7,9) #71
wire n12227_0;
wire n12228; //CHANX 3 (7,9) #78
wire n12228_0;
wire n12229; //CHANX 3 (7,9) #79
wire n12229_0;
wire n12230; //CHANX 2 (8,9) #0
wire n12230_0;
wire n12231; //CHANX 2 (8,9) #1
wire n12231_0;
wire n12232; //CHANX 2 (8,9) #8
wire n12232_0;
wire n12233; //CHANX 2 (8,9) #9
wire n12233_0;
wire n12234; //CHANX 2 (8,9) #16
wire n12234_0;
wire n12235; //CHANX 2 (8,9) #17
wire n12235_0;
wire n12236; //CHANX 2 (8,9) #24
wire n12236_0;
wire n12237; //CHANX 2 (8,9) #25
wire n12237_0;
wire n12238; //CHANX 2 (8,9) #32
wire n12238_0;
wire n12239; //CHANX 2 (8,9) #33
wire n12239_0;
wire n12240; //CHANX 2 (8,9) #40
wire n12240_0;
wire n12241; //CHANX 2 (8,9) #41
wire n12241_0;
wire n12242; //CHANX 2 (8,9) #48
wire n12242_0;
wire n12243; //CHANX 2 (8,9) #49
wire n12243_0;
wire n12244; //CHANX 2 (8,9) #56
wire n12244_0;
wire n12245; //CHANX 2 (8,9) #57
wire n12245_0;
wire n12246; //CHANX 2 (8,9) #64
wire n12246_0;
wire n12247; //CHANX 2 (8,9) #65
wire n12247_0;
wire n12248; //CHANX 2 (8,9) #72
wire n12248_0;
wire n12249; //CHANX 2 (8,9) #73
wire n12249_0;
wire n12250; //CHANX 1 (9,9) #2
wire n12250_0;
wire n12251; //CHANX 1 (9,9) #3
wire n12251_0;
wire n12252; //CHANX 1 (9,9) #10
wire n12252_0;
wire n12253; //CHANX 1 (9,9) #11
wire n12253_0;
wire n12254; //CHANX 1 (9,9) #18
wire n12254_0;
wire n12255; //CHANX 1 (9,9) #19
wire n12255_0;
wire n12256; //CHANX 1 (9,9) #26
wire n12256_0;
wire n12257; //CHANX 1 (9,9) #27
wire n12257_0;
wire n12258; //CHANX 1 (9,9) #34
wire n12258_0;
wire n12259; //CHANX 1 (9,9) #35
wire n12259_0;
wire n12260; //CHANX 1 (9,9) #42
wire n12260_0;
wire n12261; //CHANX 1 (9,9) #43
wire n12261_0;
wire n12262; //CHANX 1 (9,9) #50
wire n12262_0;
wire n12263; //CHANX 1 (9,9) #51
wire n12263_0;
wire n12264; //CHANX 1 (9,9) #58
wire n12264_0;
wire n12265; //CHANX 1 (9,9) #59
wire n12265_0;
wire n12266; //CHANX 1 (9,9) #66
wire n12266_0;
wire n12267; //CHANX 1 (9,9) #67
wire n12267_0;
wire n12268; //CHANX 1 (9,9) #74
wire n12268_0;
wire n12269; //CHANX 1 (9,9) #75
wire n12269_0;
wire n12270; //CHANY 4 (0,1) #0
wire n12270_0;
wire n12270_1;
buffer_wire buffer_12270_1 (.in(n12270_0), .out(n12270_1));
wire n12271; //CHANY 4 (0,1) #1
wire n12271_0;
wire n12271_1;
buffer_wire buffer_12271_1 (.in(n12271_0), .out(n12271_1));
wire n12272; //CHANY 1 (0,1) #2
wire n12272_0;
wire n12273; //CHANY 1 (0,1) #3
wire n12273_0;
wire n12274; //CHANY 2 (0,1) #4
wire n12274_0;
wire n12275; //CHANY 2 (0,1) #5
wire n12275_0;
wire n12276; //CHANY 3 (0,1) #6
wire n12276_0;
wire n12277; //CHANY 3 (0,1) #7
wire n12277_0;
wire n12278; //CHANY 4 (0,1) #8
wire n12278_0;
wire n12278_1;
buffer_wire buffer_12278_1 (.in(n12278_0), .out(n12278_1));
wire n12279; //CHANY 4 (0,1) #9
wire n12279_0;
wire n12279_1;
buffer_wire buffer_12279_1 (.in(n12279_0), .out(n12279_1));
wire n12280; //CHANY 1 (0,1) #10
wire n12280_0;
wire n12281; //CHANY 1 (0,1) #11
wire n12281_0;
wire n12282; //CHANY 2 (0,1) #12
wire n12282_0;
wire n12283; //CHANY 2 (0,1) #13
wire n12283_0;
wire n12284; //CHANY 3 (0,1) #14
wire n12284_0;
wire n12285; //CHANY 3 (0,1) #15
wire n12285_0;
wire n12286; //CHANY 4 (0,1) #16
wire n12286_0;
wire n12286_1;
buffer_wire buffer_12286_1 (.in(n12286_0), .out(n12286_1));
wire n12287; //CHANY 4 (0,1) #17
wire n12287_0;
wire n12287_1;
buffer_wire buffer_12287_1 (.in(n12287_0), .out(n12287_1));
wire n12288; //CHANY 1 (0,1) #18
wire n12288_0;
wire n12289; //CHANY 1 (0,1) #19
wire n12289_0;
wire n12290; //CHANY 2 (0,1) #20
wire n12290_0;
wire n12291; //CHANY 2 (0,1) #21
wire n12291_0;
wire n12292; //CHANY 3 (0,1) #22
wire n12292_0;
wire n12293; //CHANY 3 (0,1) #23
wire n12293_0;
wire n12294; //CHANY 4 (0,1) #24
wire n12294_0;
wire n12294_1;
buffer_wire buffer_12294_1 (.in(n12294_0), .out(n12294_1));
wire n12295; //CHANY 4 (0,1) #25
wire n12295_0;
wire n12295_1;
buffer_wire buffer_12295_1 (.in(n12295_0), .out(n12295_1));
wire n12296; //CHANY 1 (0,1) #26
wire n12296_0;
wire n12297; //CHANY 1 (0,1) #27
wire n12297_0;
wire n12298; //CHANY 2 (0,1) #28
wire n12298_0;
wire n12299; //CHANY 2 (0,1) #29
wire n12299_0;
wire n12300; //CHANY 3 (0,1) #30
wire n12300_0;
wire n12301; //CHANY 3 (0,1) #31
wire n12301_0;
wire n12302; //CHANY 4 (0,1) #32
wire n12302_0;
wire n12302_1;
buffer_wire buffer_12302_1 (.in(n12302_0), .out(n12302_1));
wire n12303; //CHANY 4 (0,1) #33
wire n12303_0;
wire n12303_1;
buffer_wire buffer_12303_1 (.in(n12303_0), .out(n12303_1));
wire n12304; //CHANY 1 (0,1) #34
wire n12304_0;
wire n12305; //CHANY 1 (0,1) #35
wire n12305_0;
wire n12306; //CHANY 2 (0,1) #36
wire n12306_0;
wire n12307; //CHANY 2 (0,1) #37
wire n12307_0;
wire n12308; //CHANY 3 (0,1) #38
wire n12308_0;
wire n12309; //CHANY 3 (0,1) #39
wire n12309_0;
wire n12310; //CHANY 4 (0,1) #40
wire n12310_0;
wire n12310_1;
buffer_wire buffer_12310_1 (.in(n12310_0), .out(n12310_1));
wire n12311; //CHANY 4 (0,1) #41
wire n12311_0;
wire n12311_1;
buffer_wire buffer_12311_1 (.in(n12311_0), .out(n12311_1));
wire n12312; //CHANY 1 (0,1) #42
wire n12312_0;
wire n12313; //CHANY 1 (0,1) #43
wire n12313_0;
wire n12314; //CHANY 2 (0,1) #44
wire n12314_0;
wire n12315; //CHANY 2 (0,1) #45
wire n12315_0;
wire n12316; //CHANY 3 (0,1) #46
wire n12316_0;
wire n12317; //CHANY 3 (0,1) #47
wire n12317_0;
wire n12318; //CHANY 4 (0,1) #48
wire n12318_0;
wire n12318_1;
buffer_wire buffer_12318_1 (.in(n12318_0), .out(n12318_1));
wire n12319; //CHANY 4 (0,1) #49
wire n12319_0;
wire n12319_1;
buffer_wire buffer_12319_1 (.in(n12319_0), .out(n12319_1));
wire n12320; //CHANY 1 (0,1) #50
wire n12320_0;
wire n12321; //CHANY 1 (0,1) #51
wire n12321_0;
wire n12322; //CHANY 2 (0,1) #52
wire n12322_0;
wire n12323; //CHANY 2 (0,1) #53
wire n12323_0;
wire n12324; //CHANY 3 (0,1) #54
wire n12324_0;
wire n12325; //CHANY 3 (0,1) #55
wire n12325_0;
wire n12326; //CHANY 4 (0,1) #56
wire n12326_0;
wire n12326_1;
buffer_wire buffer_12326_1 (.in(n12326_0), .out(n12326_1));
wire n12327; //CHANY 4 (0,1) #57
wire n12327_0;
wire n12327_1;
buffer_wire buffer_12327_1 (.in(n12327_0), .out(n12327_1));
wire n12328; //CHANY 1 (0,1) #58
wire n12328_0;
wire n12329; //CHANY 1 (0,1) #59
wire n12329_0;
wire n12330; //CHANY 2 (0,1) #60
wire n12330_0;
wire n12331; //CHANY 2 (0,1) #61
wire n12331_0;
wire n12332; //CHANY 3 (0,1) #62
wire n12332_0;
wire n12333; //CHANY 3 (0,1) #63
wire n12333_0;
wire n12334; //CHANY 4 (0,1) #64
wire n12334_0;
wire n12334_1;
buffer_wire buffer_12334_1 (.in(n12334_0), .out(n12334_1));
wire n12335; //CHANY 4 (0,1) #65
wire n12335_0;
wire n12335_1;
buffer_wire buffer_12335_1 (.in(n12335_0), .out(n12335_1));
wire n12336; //CHANY 1 (0,1) #66
wire n12336_0;
wire n12337; //CHANY 1 (0,1) #67
wire n12337_0;
wire n12338; //CHANY 2 (0,1) #68
wire n12338_0;
wire n12339; //CHANY 2 (0,1) #69
wire n12339_0;
wire n12340; //CHANY 3 (0,1) #70
wire n12340_0;
wire n12341; //CHANY 3 (0,1) #71
wire n12341_0;
wire n12342; //CHANY 4 (0,1) #72
wire n12342_0;
wire n12342_1;
buffer_wire buffer_12342_1 (.in(n12342_0), .out(n12342_1));
wire n12343; //CHANY 4 (0,1) #73
wire n12343_0;
wire n12343_1;
buffer_wire buffer_12343_1 (.in(n12343_0), .out(n12343_1));
wire n12344; //CHANY 1 (0,1) #74
wire n12344_0;
wire n12345; //CHANY 1 (0,1) #75
wire n12345_0;
wire n12346; //CHANY 2 (0,1) #76
wire n12346_0;
wire n12347; //CHANY 2 (0,1) #77
wire n12347_0;
wire n12348; //CHANY 3 (0,1) #78
wire n12348_0;
wire n12349; //CHANY 3 (0,1) #79
wire n12349_0;
wire n12350; //CHANY 8 (0,1) #80
wire n12350_0;
wire n12350_1;
wire n12350_2;
buffer_wire buffer_12350_2 (.in(n12350_1), .out(n12350_2));
buffer_wire buffer_12350_1 (.in(n12350_0), .out(n12350_1));
wire n12351; //CHANY 8 (0,1) #81
wire n12351_0;
wire n12351_1;
wire n12351_2;
buffer_wire buffer_12351_2 (.in(n12351_1), .out(n12351_2));
buffer_wire buffer_12351_1 (.in(n12351_0), .out(n12351_1));
wire n12352; //CHANY 9 (0,1) #82
wire n12352_0;
wire n12352_1;
wire n12352_2;
buffer_wire buffer_12352_2 (.in(n12352_1), .out(n12352_2));
buffer_wire buffer_12352_1 (.in(n12352_0), .out(n12352_1));
wire n12353; //CHANY 9 (0,1) #83
wire n12353_0;
wire n12353_1;
wire n12353_2;
buffer_wire buffer_12353_2 (.in(n12353_1), .out(n12353_2));
buffer_wire buffer_12353_1 (.in(n12353_0), .out(n12353_1));
wire n12354; //CHANY 9 (0,1) #84
wire n12354_0;
wire n12354_1;
wire n12354_2;
buffer_wire buffer_12354_2 (.in(n12354_1), .out(n12354_2));
buffer_wire buffer_12354_1 (.in(n12354_0), .out(n12354_1));
wire n12355; //CHANY 9 (0,1) #85
wire n12355_0;
wire n12355_1;
wire n12355_2;
buffer_wire buffer_12355_2 (.in(n12355_1), .out(n12355_2));
buffer_wire buffer_12355_1 (.in(n12355_0), .out(n12355_1));
wire n12356; //CHANY 9 (0,1) #86
wire n12356_0;
wire n12356_1;
wire n12356_2;
buffer_wire buffer_12356_2 (.in(n12356_1), .out(n12356_2));
buffer_wire buffer_12356_1 (.in(n12356_0), .out(n12356_1));
wire n12357; //CHANY 9 (0,1) #87
wire n12357_0;
wire n12357_1;
wire n12357_2;
buffer_wire buffer_12357_2 (.in(n12357_1), .out(n12357_2));
buffer_wire buffer_12357_1 (.in(n12357_0), .out(n12357_1));
wire n12358; //CHANY 9 (0,1) #88
wire n12358_0;
wire n12358_1;
wire n12358_2;
buffer_wire buffer_12358_2 (.in(n12358_1), .out(n12358_2));
buffer_wire buffer_12358_1 (.in(n12358_0), .out(n12358_1));
wire n12359; //CHANY 9 (0,1) #89
wire n12359_0;
wire n12359_1;
wire n12359_2;
buffer_wire buffer_12359_2 (.in(n12359_1), .out(n12359_2));
buffer_wire buffer_12359_1 (.in(n12359_0), .out(n12359_1));
wire n12360; //CHANY 9 (0,1) #90
wire n12360_0;
wire n12360_1;
wire n12360_2;
buffer_wire buffer_12360_2 (.in(n12360_1), .out(n12360_2));
buffer_wire buffer_12360_1 (.in(n12360_0), .out(n12360_1));
wire n12361; //CHANY 9 (0,1) #91
wire n12361_0;
wire n12361_1;
wire n12361_2;
buffer_wire buffer_12361_2 (.in(n12361_1), .out(n12361_2));
buffer_wire buffer_12361_1 (.in(n12361_0), .out(n12361_1));
wire n12362; //CHANY 4 (0,2) #2
wire n12362_0;
wire n12362_1;
buffer_wire buffer_12362_1 (.in(n12362_0), .out(n12362_1));
wire n12363; //CHANY 4 (0,2) #3
wire n12363_0;
wire n12363_1;
buffer_wire buffer_12363_1 (.in(n12363_0), .out(n12363_1));
wire n12364; //CHANY 4 (0,2) #10
wire n12364_0;
wire n12364_1;
buffer_wire buffer_12364_1 (.in(n12364_0), .out(n12364_1));
wire n12365; //CHANY 4 (0,2) #11
wire n12365_0;
wire n12365_1;
buffer_wire buffer_12365_1 (.in(n12365_0), .out(n12365_1));
wire n12366; //CHANY 4 (0,2) #18
wire n12366_0;
wire n12366_1;
buffer_wire buffer_12366_1 (.in(n12366_0), .out(n12366_1));
wire n12367; //CHANY 4 (0,2) #19
wire n12367_0;
wire n12367_1;
buffer_wire buffer_12367_1 (.in(n12367_0), .out(n12367_1));
wire n12368; //CHANY 4 (0,2) #26
wire n12368_0;
wire n12368_1;
buffer_wire buffer_12368_1 (.in(n12368_0), .out(n12368_1));
wire n12369; //CHANY 4 (0,2) #27
wire n12369_0;
wire n12369_1;
buffer_wire buffer_12369_1 (.in(n12369_0), .out(n12369_1));
wire n12370; //CHANY 4 (0,2) #34
wire n12370_0;
wire n12370_1;
buffer_wire buffer_12370_1 (.in(n12370_0), .out(n12370_1));
wire n12371; //CHANY 4 (0,2) #35
wire n12371_0;
wire n12371_1;
buffer_wire buffer_12371_1 (.in(n12371_0), .out(n12371_1));
wire n12372; //CHANY 4 (0,2) #42
wire n12372_0;
wire n12372_1;
buffer_wire buffer_12372_1 (.in(n12372_0), .out(n12372_1));
wire n12373; //CHANY 4 (0,2) #43
wire n12373_0;
wire n12373_1;
buffer_wire buffer_12373_1 (.in(n12373_0), .out(n12373_1));
wire n12374; //CHANY 4 (0,2) #50
wire n12374_0;
wire n12374_1;
buffer_wire buffer_12374_1 (.in(n12374_0), .out(n12374_1));
wire n12375; //CHANY 4 (0,2) #51
wire n12375_0;
wire n12375_1;
buffer_wire buffer_12375_1 (.in(n12375_0), .out(n12375_1));
wire n12376; //CHANY 4 (0,2) #58
wire n12376_0;
wire n12376_1;
buffer_wire buffer_12376_1 (.in(n12376_0), .out(n12376_1));
wire n12377; //CHANY 4 (0,2) #59
wire n12377_0;
wire n12377_1;
buffer_wire buffer_12377_1 (.in(n12377_0), .out(n12377_1));
wire n12378; //CHANY 4 (0,2) #66
wire n12378_0;
wire n12378_1;
buffer_wire buffer_12378_1 (.in(n12378_0), .out(n12378_1));
wire n12379; //CHANY 4 (0,2) #67
wire n12379_0;
wire n12379_1;
buffer_wire buffer_12379_1 (.in(n12379_0), .out(n12379_1));
wire n12380; //CHANY 4 (0,2) #74
wire n12380_0;
wire n12380_1;
buffer_wire buffer_12380_1 (.in(n12380_0), .out(n12380_1));
wire n12381; //CHANY 4 (0,2) #75
wire n12381_0;
wire n12381_1;
buffer_wire buffer_12381_1 (.in(n12381_0), .out(n12381_1));
wire n12382; //CHANY 4 (0,3) #4
wire n12382_0;
wire n12382_1;
buffer_wire buffer_12382_1 (.in(n12382_0), .out(n12382_1));
wire n12383; //CHANY 4 (0,3) #5
wire n12383_0;
wire n12383_1;
buffer_wire buffer_12383_1 (.in(n12383_0), .out(n12383_1));
wire n12384; //CHANY 4 (0,3) #12
wire n12384_0;
wire n12384_1;
buffer_wire buffer_12384_1 (.in(n12384_0), .out(n12384_1));
wire n12385; //CHANY 4 (0,3) #13
wire n12385_0;
wire n12385_1;
buffer_wire buffer_12385_1 (.in(n12385_0), .out(n12385_1));
wire n12386; //CHANY 4 (0,3) #20
wire n12386_0;
wire n12386_1;
buffer_wire buffer_12386_1 (.in(n12386_0), .out(n12386_1));
wire n12387; //CHANY 4 (0,3) #21
wire n12387_0;
wire n12387_1;
buffer_wire buffer_12387_1 (.in(n12387_0), .out(n12387_1));
wire n12388; //CHANY 4 (0,3) #28
wire n12388_0;
wire n12388_1;
buffer_wire buffer_12388_1 (.in(n12388_0), .out(n12388_1));
wire n12389; //CHANY 4 (0,3) #29
wire n12389_0;
wire n12389_1;
buffer_wire buffer_12389_1 (.in(n12389_0), .out(n12389_1));
wire n12390; //CHANY 4 (0,3) #36
wire n12390_0;
wire n12390_1;
buffer_wire buffer_12390_1 (.in(n12390_0), .out(n12390_1));
wire n12391; //CHANY 4 (0,3) #37
wire n12391_0;
wire n12391_1;
buffer_wire buffer_12391_1 (.in(n12391_0), .out(n12391_1));
wire n12392; //CHANY 4 (0,3) #44
wire n12392_0;
wire n12392_1;
buffer_wire buffer_12392_1 (.in(n12392_0), .out(n12392_1));
wire n12393; //CHANY 4 (0,3) #45
wire n12393_0;
wire n12393_1;
buffer_wire buffer_12393_1 (.in(n12393_0), .out(n12393_1));
wire n12394; //CHANY 4 (0,3) #52
wire n12394_0;
wire n12394_1;
buffer_wire buffer_12394_1 (.in(n12394_0), .out(n12394_1));
wire n12395; //CHANY 4 (0,3) #53
wire n12395_0;
wire n12395_1;
buffer_wire buffer_12395_1 (.in(n12395_0), .out(n12395_1));
wire n12396; //CHANY 4 (0,3) #60
wire n12396_0;
wire n12396_1;
buffer_wire buffer_12396_1 (.in(n12396_0), .out(n12396_1));
wire n12397; //CHANY 4 (0,3) #61
wire n12397_0;
wire n12397_1;
buffer_wire buffer_12397_1 (.in(n12397_0), .out(n12397_1));
wire n12398; //CHANY 4 (0,3) #68
wire n12398_0;
wire n12398_1;
buffer_wire buffer_12398_1 (.in(n12398_0), .out(n12398_1));
wire n12399; //CHANY 4 (0,3) #69
wire n12399_0;
wire n12399_1;
buffer_wire buffer_12399_1 (.in(n12399_0), .out(n12399_1));
wire n12400; //CHANY 4 (0,3) #76
wire n12400_0;
wire n12400_1;
buffer_wire buffer_12400_1 (.in(n12400_0), .out(n12400_1));
wire n12401; //CHANY 4 (0,3) #77
wire n12401_0;
wire n12401_1;
buffer_wire buffer_12401_1 (.in(n12401_0), .out(n12401_1));
wire n12402; //CHANY 4 (0,4) #6
wire n12402_0;
wire n12402_1;
buffer_wire buffer_12402_1 (.in(n12402_0), .out(n12402_1));
wire n12403; //CHANY 4 (0,4) #7
wire n12403_0;
wire n12403_1;
buffer_wire buffer_12403_1 (.in(n12403_0), .out(n12403_1));
wire n12404; //CHANY 4 (0,4) #14
wire n12404_0;
wire n12404_1;
buffer_wire buffer_12404_1 (.in(n12404_0), .out(n12404_1));
wire n12405; //CHANY 4 (0,4) #15
wire n12405_0;
wire n12405_1;
buffer_wire buffer_12405_1 (.in(n12405_0), .out(n12405_1));
wire n12406; //CHANY 4 (0,4) #22
wire n12406_0;
wire n12406_1;
buffer_wire buffer_12406_1 (.in(n12406_0), .out(n12406_1));
wire n12407; //CHANY 4 (0,4) #23
wire n12407_0;
wire n12407_1;
buffer_wire buffer_12407_1 (.in(n12407_0), .out(n12407_1));
wire n12408; //CHANY 4 (0,4) #30
wire n12408_0;
wire n12408_1;
buffer_wire buffer_12408_1 (.in(n12408_0), .out(n12408_1));
wire n12409; //CHANY 4 (0,4) #31
wire n12409_0;
wire n12409_1;
buffer_wire buffer_12409_1 (.in(n12409_0), .out(n12409_1));
wire n12410; //CHANY 4 (0,4) #38
wire n12410_0;
wire n12410_1;
buffer_wire buffer_12410_1 (.in(n12410_0), .out(n12410_1));
wire n12411; //CHANY 4 (0,4) #39
wire n12411_0;
wire n12411_1;
buffer_wire buffer_12411_1 (.in(n12411_0), .out(n12411_1));
wire n12412; //CHANY 4 (0,4) #46
wire n12412_0;
wire n12412_1;
buffer_wire buffer_12412_1 (.in(n12412_0), .out(n12412_1));
wire n12413; //CHANY 4 (0,4) #47
wire n12413_0;
wire n12413_1;
buffer_wire buffer_12413_1 (.in(n12413_0), .out(n12413_1));
wire n12414; //CHANY 4 (0,4) #54
wire n12414_0;
wire n12414_1;
buffer_wire buffer_12414_1 (.in(n12414_0), .out(n12414_1));
wire n12415; //CHANY 4 (0,4) #55
wire n12415_0;
wire n12415_1;
buffer_wire buffer_12415_1 (.in(n12415_0), .out(n12415_1));
wire n12416; //CHANY 4 (0,4) #62
wire n12416_0;
wire n12416_1;
buffer_wire buffer_12416_1 (.in(n12416_0), .out(n12416_1));
wire n12417; //CHANY 4 (0,4) #63
wire n12417_0;
wire n12417_1;
buffer_wire buffer_12417_1 (.in(n12417_0), .out(n12417_1));
wire n12418; //CHANY 4 (0,4) #70
wire n12418_0;
wire n12418_1;
buffer_wire buffer_12418_1 (.in(n12418_0), .out(n12418_1));
wire n12419; //CHANY 4 (0,4) #71
wire n12419_0;
wire n12419_1;
buffer_wire buffer_12419_1 (.in(n12419_0), .out(n12419_1));
wire n12420; //CHANY 4 (0,4) #78
wire n12420_0;
wire n12420_1;
buffer_wire buffer_12420_1 (.in(n12420_0), .out(n12420_1));
wire n12421; //CHANY 4 (0,4) #79
wire n12421_0;
wire n12421_1;
buffer_wire buffer_12421_1 (.in(n12421_0), .out(n12421_1));
wire n12422; //CHANY 4 (0,5) #0
wire n12422_0;
wire n12422_1;
buffer_wire buffer_12422_1 (.in(n12422_0), .out(n12422_1));
wire n12423; //CHANY 4 (0,5) #1
wire n12423_0;
wire n12423_1;
buffer_wire buffer_12423_1 (.in(n12423_0), .out(n12423_1));
wire n12424; //CHANY 4 (0,5) #8
wire n12424_0;
wire n12424_1;
buffer_wire buffer_12424_1 (.in(n12424_0), .out(n12424_1));
wire n12425; //CHANY 4 (0,5) #9
wire n12425_0;
wire n12425_1;
buffer_wire buffer_12425_1 (.in(n12425_0), .out(n12425_1));
wire n12426; //CHANY 4 (0,5) #16
wire n12426_0;
wire n12426_1;
buffer_wire buffer_12426_1 (.in(n12426_0), .out(n12426_1));
wire n12427; //CHANY 4 (0,5) #17
wire n12427_0;
wire n12427_1;
buffer_wire buffer_12427_1 (.in(n12427_0), .out(n12427_1));
wire n12428; //CHANY 4 (0,5) #24
wire n12428_0;
wire n12428_1;
buffer_wire buffer_12428_1 (.in(n12428_0), .out(n12428_1));
wire n12429; //CHANY 4 (0,5) #25
wire n12429_0;
wire n12429_1;
buffer_wire buffer_12429_1 (.in(n12429_0), .out(n12429_1));
wire n12430; //CHANY 4 (0,5) #32
wire n12430_0;
wire n12430_1;
buffer_wire buffer_12430_1 (.in(n12430_0), .out(n12430_1));
wire n12431; //CHANY 4 (0,5) #33
wire n12431_0;
wire n12431_1;
buffer_wire buffer_12431_1 (.in(n12431_0), .out(n12431_1));
wire n12432; //CHANY 4 (0,5) #40
wire n12432_0;
wire n12432_1;
buffer_wire buffer_12432_1 (.in(n12432_0), .out(n12432_1));
wire n12433; //CHANY 4 (0,5) #41
wire n12433_0;
wire n12433_1;
buffer_wire buffer_12433_1 (.in(n12433_0), .out(n12433_1));
wire n12434; //CHANY 4 (0,5) #48
wire n12434_0;
wire n12434_1;
buffer_wire buffer_12434_1 (.in(n12434_0), .out(n12434_1));
wire n12435; //CHANY 4 (0,5) #49
wire n12435_0;
wire n12435_1;
buffer_wire buffer_12435_1 (.in(n12435_0), .out(n12435_1));
wire n12436; //CHANY 4 (0,5) #56
wire n12436_0;
wire n12436_1;
buffer_wire buffer_12436_1 (.in(n12436_0), .out(n12436_1));
wire n12437; //CHANY 4 (0,5) #57
wire n12437_0;
wire n12437_1;
buffer_wire buffer_12437_1 (.in(n12437_0), .out(n12437_1));
wire n12438; //CHANY 4 (0,5) #64
wire n12438_0;
wire n12438_1;
buffer_wire buffer_12438_1 (.in(n12438_0), .out(n12438_1));
wire n12439; //CHANY 4 (0,5) #65
wire n12439_0;
wire n12439_1;
buffer_wire buffer_12439_1 (.in(n12439_0), .out(n12439_1));
wire n12440; //CHANY 4 (0,5) #72
wire n12440_0;
wire n12440_1;
buffer_wire buffer_12440_1 (.in(n12440_0), .out(n12440_1));
wire n12441; //CHANY 4 (0,5) #73
wire n12441_0;
wire n12441_1;
buffer_wire buffer_12441_1 (.in(n12441_0), .out(n12441_1));
wire n12442; //CHANY 4 (0,6) #2
wire n12442_0;
wire n12442_1;
buffer_wire buffer_12442_1 (.in(n12442_0), .out(n12442_1));
wire n12443; //CHANY 4 (0,6) #3
wire n12443_0;
wire n12443_1;
buffer_wire buffer_12443_1 (.in(n12443_0), .out(n12443_1));
wire n12444; //CHANY 4 (0,6) #10
wire n12444_0;
wire n12444_1;
buffer_wire buffer_12444_1 (.in(n12444_0), .out(n12444_1));
wire n12445; //CHANY 4 (0,6) #11
wire n12445_0;
wire n12445_1;
buffer_wire buffer_12445_1 (.in(n12445_0), .out(n12445_1));
wire n12446; //CHANY 4 (0,6) #18
wire n12446_0;
wire n12446_1;
buffer_wire buffer_12446_1 (.in(n12446_0), .out(n12446_1));
wire n12447; //CHANY 4 (0,6) #19
wire n12447_0;
wire n12447_1;
buffer_wire buffer_12447_1 (.in(n12447_0), .out(n12447_1));
wire n12448; //CHANY 4 (0,6) #26
wire n12448_0;
wire n12448_1;
buffer_wire buffer_12448_1 (.in(n12448_0), .out(n12448_1));
wire n12449; //CHANY 4 (0,6) #27
wire n12449_0;
wire n12449_1;
buffer_wire buffer_12449_1 (.in(n12449_0), .out(n12449_1));
wire n12450; //CHANY 4 (0,6) #34
wire n12450_0;
wire n12450_1;
buffer_wire buffer_12450_1 (.in(n12450_0), .out(n12450_1));
wire n12451; //CHANY 4 (0,6) #35
wire n12451_0;
wire n12451_1;
buffer_wire buffer_12451_1 (.in(n12451_0), .out(n12451_1));
wire n12452; //CHANY 4 (0,6) #42
wire n12452_0;
wire n12452_1;
buffer_wire buffer_12452_1 (.in(n12452_0), .out(n12452_1));
wire n12453; //CHANY 4 (0,6) #43
wire n12453_0;
wire n12453_1;
buffer_wire buffer_12453_1 (.in(n12453_0), .out(n12453_1));
wire n12454; //CHANY 4 (0,6) #50
wire n12454_0;
wire n12454_1;
buffer_wire buffer_12454_1 (.in(n12454_0), .out(n12454_1));
wire n12455; //CHANY 4 (0,6) #51
wire n12455_0;
wire n12455_1;
buffer_wire buffer_12455_1 (.in(n12455_0), .out(n12455_1));
wire n12456; //CHANY 4 (0,6) #58
wire n12456_0;
wire n12456_1;
buffer_wire buffer_12456_1 (.in(n12456_0), .out(n12456_1));
wire n12457; //CHANY 4 (0,6) #59
wire n12457_0;
wire n12457_1;
buffer_wire buffer_12457_1 (.in(n12457_0), .out(n12457_1));
wire n12458; //CHANY 4 (0,6) #66
wire n12458_0;
wire n12458_1;
buffer_wire buffer_12458_1 (.in(n12458_0), .out(n12458_1));
wire n12459; //CHANY 4 (0,6) #67
wire n12459_0;
wire n12459_1;
buffer_wire buffer_12459_1 (.in(n12459_0), .out(n12459_1));
wire n12460; //CHANY 4 (0,6) #74
wire n12460_0;
wire n12460_1;
buffer_wire buffer_12460_1 (.in(n12460_0), .out(n12460_1));
wire n12461; //CHANY 4 (0,6) #75
wire n12461_0;
wire n12461_1;
buffer_wire buffer_12461_1 (.in(n12461_0), .out(n12461_1));
wire n12462; //CHANY 3 (0,7) #4
wire n12462_0;
wire n12463; //CHANY 3 (0,7) #5
wire n12463_0;
wire n12464; //CHANY 3 (0,7) #12
wire n12464_0;
wire n12465; //CHANY 3 (0,7) #13
wire n12465_0;
wire n12466; //CHANY 3 (0,7) #20
wire n12466_0;
wire n12467; //CHANY 3 (0,7) #21
wire n12467_0;
wire n12468; //CHANY 3 (0,7) #28
wire n12468_0;
wire n12469; //CHANY 3 (0,7) #29
wire n12469_0;
wire n12470; //CHANY 3 (0,7) #36
wire n12470_0;
wire n12471; //CHANY 3 (0,7) #37
wire n12471_0;
wire n12472; //CHANY 3 (0,7) #44
wire n12472_0;
wire n12473; //CHANY 3 (0,7) #45
wire n12473_0;
wire n12474; //CHANY 3 (0,7) #52
wire n12474_0;
wire n12475; //CHANY 3 (0,7) #53
wire n12475_0;
wire n12476; //CHANY 3 (0,7) #60
wire n12476_0;
wire n12477; //CHANY 3 (0,7) #61
wire n12477_0;
wire n12478; //CHANY 3 (0,7) #68
wire n12478_0;
wire n12479; //CHANY 3 (0,7) #69
wire n12479_0;
wire n12480; //CHANY 3 (0,7) #76
wire n12480_0;
wire n12481; //CHANY 3 (0,7) #77
wire n12481_0;
wire n12482; //CHANY 2 (0,8) #6
wire n12482_0;
wire n12483; //CHANY 2 (0,8) #7
wire n12483_0;
wire n12484; //CHANY 2 (0,8) #14
wire n12484_0;
wire n12485; //CHANY 2 (0,8) #15
wire n12485_0;
wire n12486; //CHANY 2 (0,8) #22
wire n12486_0;
wire n12487; //CHANY 2 (0,8) #23
wire n12487_0;
wire n12488; //CHANY 2 (0,8) #30
wire n12488_0;
wire n12489; //CHANY 2 (0,8) #31
wire n12489_0;
wire n12490; //CHANY 2 (0,8) #38
wire n12490_0;
wire n12491; //CHANY 2 (0,8) #39
wire n12491_0;
wire n12492; //CHANY 2 (0,8) #46
wire n12492_0;
wire n12493; //CHANY 2 (0,8) #47
wire n12493_0;
wire n12494; //CHANY 2 (0,8) #54
wire n12494_0;
wire n12495; //CHANY 2 (0,8) #55
wire n12495_0;
wire n12496; //CHANY 2 (0,8) #62
wire n12496_0;
wire n12497; //CHANY 2 (0,8) #63
wire n12497_0;
wire n12498; //CHANY 2 (0,8) #70
wire n12498_0;
wire n12499; //CHANY 2 (0,8) #71
wire n12499_0;
wire n12500; //CHANY 2 (0,8) #78
wire n12500_0;
wire n12501; //CHANY 2 (0,8) #79
wire n12501_0;
wire n12502; //CHANY 1 (0,9) #0
wire n12502_0;
wire n12503; //CHANY 1 (0,9) #1
wire n12503_0;
wire n12504; //CHANY 1 (0,9) #8
wire n12504_0;
wire n12505; //CHANY 1 (0,9) #9
wire n12505_0;
wire n12506; //CHANY 1 (0,9) #16
wire n12506_0;
wire n12507; //CHANY 1 (0,9) #17
wire n12507_0;
wire n12508; //CHANY 1 (0,9) #24
wire n12508_0;
wire n12509; //CHANY 1 (0,9) #25
wire n12509_0;
wire n12510; //CHANY 1 (0,9) #32
wire n12510_0;
wire n12511; //CHANY 1 (0,9) #33
wire n12511_0;
wire n12512; //CHANY 1 (0,9) #40
wire n12512_0;
wire n12513; //CHANY 1 (0,9) #41
wire n12513_0;
wire n12514; //CHANY 1 (0,9) #48
wire n12514_0;
wire n12515; //CHANY 1 (0,9) #49
wire n12515_0;
wire n12516; //CHANY 1 (0,9) #56
wire n12516_0;
wire n12517; //CHANY 1 (0,9) #57
wire n12517_0;
wire n12518; //CHANY 1 (0,9) #64
wire n12518_0;
wire n12519; //CHANY 1 (0,9) #65
wire n12519_0;
wire n12520; //CHANY 1 (0,9) #72
wire n12520_0;
wire n12521; //CHANY 1 (0,9) #73
wire n12521_0;
wire n12522; //CHANY 1 (0,9) #80
wire n12522_0;
wire n12523; //CHANY 1 (0,9) #81
wire n12523_0;
wire n12524; //CHANY 3 (1,1) #0
wire n12524_0;
wire n12525; //CHANY 3 (1,1) #1
wire n12525_0;
wire n12526; //CHANY 4 (1,1) #2
wire n12526_0;
wire n12526_1;
buffer_wire buffer_12526_1 (.in(n12526_0), .out(n12526_1));
wire n12527; //CHANY 4 (1,1) #3
wire n12527_0;
wire n12527_1;
buffer_wire buffer_12527_1 (.in(n12527_0), .out(n12527_1));
wire n12528; //CHANY 1 (1,1) #4
wire n12528_0;
wire n12529; //CHANY 1 (1,1) #5
wire n12529_0;
wire n12530; //CHANY 2 (1,1) #6
wire n12530_0;
wire n12531; //CHANY 2 (1,1) #7
wire n12531_0;
wire n12532; //CHANY 3 (1,1) #8
wire n12532_0;
wire n12533; //CHANY 3 (1,1) #9
wire n12533_0;
wire n12534; //CHANY 4 (1,1) #10
wire n12534_0;
wire n12534_1;
buffer_wire buffer_12534_1 (.in(n12534_0), .out(n12534_1));
wire n12535; //CHANY 4 (1,1) #11
wire n12535_0;
wire n12535_1;
buffer_wire buffer_12535_1 (.in(n12535_0), .out(n12535_1));
wire n12536; //CHANY 1 (1,1) #12
wire n12536_0;
wire n12537; //CHANY 1 (1,1) #13
wire n12537_0;
wire n12538; //CHANY 2 (1,1) #14
wire n12538_0;
wire n12539; //CHANY 2 (1,1) #15
wire n12539_0;
wire n12540; //CHANY 3 (1,1) #16
wire n12540_0;
wire n12541; //CHANY 3 (1,1) #17
wire n12541_0;
wire n12542; //CHANY 4 (1,1) #18
wire n12542_0;
wire n12542_1;
buffer_wire buffer_12542_1 (.in(n12542_0), .out(n12542_1));
wire n12543; //CHANY 4 (1,1) #19
wire n12543_0;
wire n12543_1;
buffer_wire buffer_12543_1 (.in(n12543_0), .out(n12543_1));
wire n12544; //CHANY 1 (1,1) #20
wire n12544_0;
wire n12545; //CHANY 1 (1,1) #21
wire n12545_0;
wire n12546; //CHANY 2 (1,1) #22
wire n12546_0;
wire n12547; //CHANY 2 (1,1) #23
wire n12547_0;
wire n12548; //CHANY 3 (1,1) #24
wire n12548_0;
wire n12549; //CHANY 3 (1,1) #25
wire n12549_0;
wire n12550; //CHANY 4 (1,1) #26
wire n12550_0;
wire n12550_1;
buffer_wire buffer_12550_1 (.in(n12550_0), .out(n12550_1));
wire n12551; //CHANY 4 (1,1) #27
wire n12551_0;
wire n12551_1;
buffer_wire buffer_12551_1 (.in(n12551_0), .out(n12551_1));
wire n12552; //CHANY 1 (1,1) #28
wire n12552_0;
wire n12553; //CHANY 1 (1,1) #29
wire n12553_0;
wire n12554; //CHANY 2 (1,1) #30
wire n12554_0;
wire n12555; //CHANY 2 (1,1) #31
wire n12555_0;
wire n12556; //CHANY 3 (1,1) #32
wire n12556_0;
wire n12557; //CHANY 3 (1,1) #33
wire n12557_0;
wire n12558; //CHANY 4 (1,1) #34
wire n12558_0;
wire n12558_1;
buffer_wire buffer_12558_1 (.in(n12558_0), .out(n12558_1));
wire n12559; //CHANY 4 (1,1) #35
wire n12559_0;
wire n12559_1;
buffer_wire buffer_12559_1 (.in(n12559_0), .out(n12559_1));
wire n12560; //CHANY 1 (1,1) #36
wire n12560_0;
wire n12561; //CHANY 1 (1,1) #37
wire n12561_0;
wire n12562; //CHANY 2 (1,1) #38
wire n12562_0;
wire n12563; //CHANY 2 (1,1) #39
wire n12563_0;
wire n12564; //CHANY 3 (1,1) #40
wire n12564_0;
wire n12565; //CHANY 3 (1,1) #41
wire n12565_0;
wire n12566; //CHANY 4 (1,1) #42
wire n12566_0;
wire n12566_1;
buffer_wire buffer_12566_1 (.in(n12566_0), .out(n12566_1));
wire n12567; //CHANY 4 (1,1) #43
wire n12567_0;
wire n12567_1;
buffer_wire buffer_12567_1 (.in(n12567_0), .out(n12567_1));
wire n12568; //CHANY 1 (1,1) #44
wire n12568_0;
wire n12569; //CHANY 1 (1,1) #45
wire n12569_0;
wire n12570; //CHANY 2 (1,1) #46
wire n12570_0;
wire n12571; //CHANY 2 (1,1) #47
wire n12571_0;
wire n12572; //CHANY 3 (1,1) #48
wire n12572_0;
wire n12573; //CHANY 3 (1,1) #49
wire n12573_0;
wire n12574; //CHANY 4 (1,1) #50
wire n12574_0;
wire n12574_1;
buffer_wire buffer_12574_1 (.in(n12574_0), .out(n12574_1));
wire n12575; //CHANY 4 (1,1) #51
wire n12575_0;
wire n12575_1;
buffer_wire buffer_12575_1 (.in(n12575_0), .out(n12575_1));
wire n12576; //CHANY 1 (1,1) #52
wire n12576_0;
wire n12577; //CHANY 1 (1,1) #53
wire n12577_0;
wire n12578; //CHANY 2 (1,1) #54
wire n12578_0;
wire n12579; //CHANY 2 (1,1) #55
wire n12579_0;
wire n12580; //CHANY 3 (1,1) #56
wire n12580_0;
wire n12581; //CHANY 3 (1,1) #57
wire n12581_0;
wire n12582; //CHANY 4 (1,1) #58
wire n12582_0;
wire n12582_1;
buffer_wire buffer_12582_1 (.in(n12582_0), .out(n12582_1));
wire n12583; //CHANY 4 (1,1) #59
wire n12583_0;
wire n12583_1;
buffer_wire buffer_12583_1 (.in(n12583_0), .out(n12583_1));
wire n12584; //CHANY 1 (1,1) #60
wire n12584_0;
wire n12585; //CHANY 1 (1,1) #61
wire n12585_0;
wire n12586; //CHANY 2 (1,1) #62
wire n12586_0;
wire n12587; //CHANY 2 (1,1) #63
wire n12587_0;
wire n12588; //CHANY 3 (1,1) #64
wire n12588_0;
wire n12589; //CHANY 3 (1,1) #65
wire n12589_0;
wire n12590; //CHANY 4 (1,1) #66
wire n12590_0;
wire n12590_1;
buffer_wire buffer_12590_1 (.in(n12590_0), .out(n12590_1));
wire n12591; //CHANY 4 (1,1) #67
wire n12591_0;
wire n12591_1;
buffer_wire buffer_12591_1 (.in(n12591_0), .out(n12591_1));
wire n12592; //CHANY 1 (1,1) #68
wire n12592_0;
wire n12593; //CHANY 1 (1,1) #69
wire n12593_0;
wire n12594; //CHANY 2 (1,1) #70
wire n12594_0;
wire n12595; //CHANY 2 (1,1) #71
wire n12595_0;
wire n12596; //CHANY 3 (1,1) #72
wire n12596_0;
wire n12597; //CHANY 3 (1,1) #73
wire n12597_0;
wire n12598; //CHANY 4 (1,1) #74
wire n12598_0;
wire n12598_1;
buffer_wire buffer_12598_1 (.in(n12598_0), .out(n12598_1));
wire n12599; //CHANY 4 (1,1) #75
wire n12599_0;
wire n12599_1;
buffer_wire buffer_12599_1 (.in(n12599_0), .out(n12599_1));
wire n12600; //CHANY 1 (1,1) #76
wire n12600_0;
wire n12601; //CHANY 1 (1,1) #77
wire n12601_0;
wire n12602; //CHANY 2 (1,1) #78
wire n12602_0;
wire n12603; //CHANY 2 (1,1) #79
wire n12603_0;
wire n12604; //CHANY 7 (1,1) #80
wire n12604_0;
wire n12604_1;
wire n12604_2;
buffer_wire buffer_12604_2 (.in(n12604_1), .out(n12604_2));
buffer_wire buffer_12604_1 (.in(n12604_0), .out(n12604_1));
wire n12605; //CHANY 7 (1,1) #81
wire n12605_0;
wire n12605_1;
wire n12605_2;
buffer_wire buffer_12605_2 (.in(n12605_1), .out(n12605_2));
buffer_wire buffer_12605_1 (.in(n12605_0), .out(n12605_1));
wire n12606; //CHANY 8 (1,1) #82
wire n12606_0;
wire n12606_1;
wire n12606_2;
buffer_wire buffer_12606_2 (.in(n12606_1), .out(n12606_2));
buffer_wire buffer_12606_1 (.in(n12606_0), .out(n12606_1));
wire n12607; //CHANY 8 (1,1) #83
wire n12607_0;
wire n12607_1;
wire n12607_2;
buffer_wire buffer_12607_2 (.in(n12607_1), .out(n12607_2));
buffer_wire buffer_12607_1 (.in(n12607_0), .out(n12607_1));
wire n12608; //CHANY 9 (1,1) #84
wire n12608_0;
wire n12608_1;
wire n12608_2;
buffer_wire buffer_12608_2 (.in(n12608_1), .out(n12608_2));
buffer_wire buffer_12608_1 (.in(n12608_0), .out(n12608_1));
wire n12609; //CHANY 9 (1,1) #85
wire n12609_0;
wire n12609_1;
wire n12609_2;
buffer_wire buffer_12609_2 (.in(n12609_1), .out(n12609_2));
buffer_wire buffer_12609_1 (.in(n12609_0), .out(n12609_1));
wire n12610; //CHANY 9 (1,1) #86
wire n12610_0;
wire n12610_1;
wire n12610_2;
buffer_wire buffer_12610_2 (.in(n12610_1), .out(n12610_2));
buffer_wire buffer_12610_1 (.in(n12610_0), .out(n12610_1));
wire n12611; //CHANY 9 (1,1) #87
wire n12611_0;
wire n12611_1;
wire n12611_2;
buffer_wire buffer_12611_2 (.in(n12611_1), .out(n12611_2));
buffer_wire buffer_12611_1 (.in(n12611_0), .out(n12611_1));
wire n12612; //CHANY 9 (1,1) #88
wire n12612_0;
wire n12612_1;
wire n12612_2;
buffer_wire buffer_12612_2 (.in(n12612_1), .out(n12612_2));
buffer_wire buffer_12612_1 (.in(n12612_0), .out(n12612_1));
wire n12613; //CHANY 9 (1,1) #89
wire n12613_0;
wire n12613_1;
wire n12613_2;
buffer_wire buffer_12613_2 (.in(n12613_1), .out(n12613_2));
buffer_wire buffer_12613_1 (.in(n12613_0), .out(n12613_1));
wire n12614; //CHANY 9 (1,1) #90
wire n12614_0;
wire n12614_1;
wire n12614_2;
buffer_wire buffer_12614_2 (.in(n12614_1), .out(n12614_2));
buffer_wire buffer_12614_1 (.in(n12614_0), .out(n12614_1));
wire n12615; //CHANY 9 (1,1) #91
wire n12615_0;
wire n12615_1;
wire n12615_2;
buffer_wire buffer_12615_2 (.in(n12615_1), .out(n12615_2));
buffer_wire buffer_12615_1 (.in(n12615_0), .out(n12615_1));
wire n12616; //CHANY 4 (1,2) #4
wire n12616_0;
wire n12616_1;
buffer_wire buffer_12616_1 (.in(n12616_0), .out(n12616_1));
wire n12617; //CHANY 4 (1,2) #5
wire n12617_0;
wire n12617_1;
buffer_wire buffer_12617_1 (.in(n12617_0), .out(n12617_1));
wire n12618; //CHANY 4 (1,2) #12
wire n12618_0;
wire n12618_1;
buffer_wire buffer_12618_1 (.in(n12618_0), .out(n12618_1));
wire n12619; //CHANY 4 (1,2) #13
wire n12619_0;
wire n12619_1;
buffer_wire buffer_12619_1 (.in(n12619_0), .out(n12619_1));
wire n12620; //CHANY 4 (1,2) #20
wire n12620_0;
wire n12620_1;
buffer_wire buffer_12620_1 (.in(n12620_0), .out(n12620_1));
wire n12621; //CHANY 4 (1,2) #21
wire n12621_0;
wire n12621_1;
buffer_wire buffer_12621_1 (.in(n12621_0), .out(n12621_1));
wire n12622; //CHANY 4 (1,2) #28
wire n12622_0;
wire n12622_1;
buffer_wire buffer_12622_1 (.in(n12622_0), .out(n12622_1));
wire n12623; //CHANY 4 (1,2) #29
wire n12623_0;
wire n12623_1;
buffer_wire buffer_12623_1 (.in(n12623_0), .out(n12623_1));
wire n12624; //CHANY 4 (1,2) #36
wire n12624_0;
wire n12624_1;
buffer_wire buffer_12624_1 (.in(n12624_0), .out(n12624_1));
wire n12625; //CHANY 4 (1,2) #37
wire n12625_0;
wire n12625_1;
buffer_wire buffer_12625_1 (.in(n12625_0), .out(n12625_1));
wire n12626; //CHANY 4 (1,2) #44
wire n12626_0;
wire n12626_1;
buffer_wire buffer_12626_1 (.in(n12626_0), .out(n12626_1));
wire n12627; //CHANY 4 (1,2) #45
wire n12627_0;
wire n12627_1;
buffer_wire buffer_12627_1 (.in(n12627_0), .out(n12627_1));
wire n12628; //CHANY 4 (1,2) #52
wire n12628_0;
wire n12628_1;
buffer_wire buffer_12628_1 (.in(n12628_0), .out(n12628_1));
wire n12629; //CHANY 4 (1,2) #53
wire n12629_0;
wire n12629_1;
buffer_wire buffer_12629_1 (.in(n12629_0), .out(n12629_1));
wire n12630; //CHANY 4 (1,2) #60
wire n12630_0;
wire n12630_1;
buffer_wire buffer_12630_1 (.in(n12630_0), .out(n12630_1));
wire n12631; //CHANY 4 (1,2) #61
wire n12631_0;
wire n12631_1;
buffer_wire buffer_12631_1 (.in(n12631_0), .out(n12631_1));
wire n12632; //CHANY 4 (1,2) #68
wire n12632_0;
wire n12632_1;
buffer_wire buffer_12632_1 (.in(n12632_0), .out(n12632_1));
wire n12633; //CHANY 4 (1,2) #69
wire n12633_0;
wire n12633_1;
buffer_wire buffer_12633_1 (.in(n12633_0), .out(n12633_1));
wire n12634; //CHANY 4 (1,2) #76
wire n12634_0;
wire n12634_1;
buffer_wire buffer_12634_1 (.in(n12634_0), .out(n12634_1));
wire n12635; //CHANY 4 (1,2) #77
wire n12635_0;
wire n12635_1;
buffer_wire buffer_12635_1 (.in(n12635_0), .out(n12635_1));
wire n12636; //CHANY 4 (1,3) #6
wire n12636_0;
wire n12636_1;
buffer_wire buffer_12636_1 (.in(n12636_0), .out(n12636_1));
wire n12637; //CHANY 4 (1,3) #7
wire n12637_0;
wire n12637_1;
buffer_wire buffer_12637_1 (.in(n12637_0), .out(n12637_1));
wire n12638; //CHANY 4 (1,3) #14
wire n12638_0;
wire n12638_1;
buffer_wire buffer_12638_1 (.in(n12638_0), .out(n12638_1));
wire n12639; //CHANY 4 (1,3) #15
wire n12639_0;
wire n12639_1;
buffer_wire buffer_12639_1 (.in(n12639_0), .out(n12639_1));
wire n12640; //CHANY 4 (1,3) #22
wire n12640_0;
wire n12640_1;
buffer_wire buffer_12640_1 (.in(n12640_0), .out(n12640_1));
wire n12641; //CHANY 4 (1,3) #23
wire n12641_0;
wire n12641_1;
buffer_wire buffer_12641_1 (.in(n12641_0), .out(n12641_1));
wire n12642; //CHANY 4 (1,3) #30
wire n12642_0;
wire n12642_1;
buffer_wire buffer_12642_1 (.in(n12642_0), .out(n12642_1));
wire n12643; //CHANY 4 (1,3) #31
wire n12643_0;
wire n12643_1;
buffer_wire buffer_12643_1 (.in(n12643_0), .out(n12643_1));
wire n12644; //CHANY 4 (1,3) #38
wire n12644_0;
wire n12644_1;
buffer_wire buffer_12644_1 (.in(n12644_0), .out(n12644_1));
wire n12645; //CHANY 4 (1,3) #39
wire n12645_0;
wire n12645_1;
buffer_wire buffer_12645_1 (.in(n12645_0), .out(n12645_1));
wire n12646; //CHANY 4 (1,3) #46
wire n12646_0;
wire n12646_1;
buffer_wire buffer_12646_1 (.in(n12646_0), .out(n12646_1));
wire n12647; //CHANY 4 (1,3) #47
wire n12647_0;
wire n12647_1;
buffer_wire buffer_12647_1 (.in(n12647_0), .out(n12647_1));
wire n12648; //CHANY 4 (1,3) #54
wire n12648_0;
wire n12648_1;
buffer_wire buffer_12648_1 (.in(n12648_0), .out(n12648_1));
wire n12649; //CHANY 4 (1,3) #55
wire n12649_0;
wire n12649_1;
buffer_wire buffer_12649_1 (.in(n12649_0), .out(n12649_1));
wire n12650; //CHANY 4 (1,3) #62
wire n12650_0;
wire n12650_1;
buffer_wire buffer_12650_1 (.in(n12650_0), .out(n12650_1));
wire n12651; //CHANY 4 (1,3) #63
wire n12651_0;
wire n12651_1;
buffer_wire buffer_12651_1 (.in(n12651_0), .out(n12651_1));
wire n12652; //CHANY 4 (1,3) #70
wire n12652_0;
wire n12652_1;
buffer_wire buffer_12652_1 (.in(n12652_0), .out(n12652_1));
wire n12653; //CHANY 4 (1,3) #71
wire n12653_0;
wire n12653_1;
buffer_wire buffer_12653_1 (.in(n12653_0), .out(n12653_1));
wire n12654; //CHANY 4 (1,3) #78
wire n12654_0;
wire n12654_1;
buffer_wire buffer_12654_1 (.in(n12654_0), .out(n12654_1));
wire n12655; //CHANY 4 (1,3) #79
wire n12655_0;
wire n12655_1;
buffer_wire buffer_12655_1 (.in(n12655_0), .out(n12655_1));
wire n12656; //CHANY 4 (1,4) #0
wire n12656_0;
wire n12656_1;
buffer_wire buffer_12656_1 (.in(n12656_0), .out(n12656_1));
wire n12657; //CHANY 4 (1,4) #1
wire n12657_0;
wire n12657_1;
buffer_wire buffer_12657_1 (.in(n12657_0), .out(n12657_1));
wire n12658; //CHANY 4 (1,4) #8
wire n12658_0;
wire n12658_1;
buffer_wire buffer_12658_1 (.in(n12658_0), .out(n12658_1));
wire n12659; //CHANY 4 (1,4) #9
wire n12659_0;
wire n12659_1;
buffer_wire buffer_12659_1 (.in(n12659_0), .out(n12659_1));
wire n12660; //CHANY 4 (1,4) #16
wire n12660_0;
wire n12660_1;
buffer_wire buffer_12660_1 (.in(n12660_0), .out(n12660_1));
wire n12661; //CHANY 4 (1,4) #17
wire n12661_0;
wire n12661_1;
buffer_wire buffer_12661_1 (.in(n12661_0), .out(n12661_1));
wire n12662; //CHANY 4 (1,4) #24
wire n12662_0;
wire n12662_1;
buffer_wire buffer_12662_1 (.in(n12662_0), .out(n12662_1));
wire n12663; //CHANY 4 (1,4) #25
wire n12663_0;
wire n12663_1;
buffer_wire buffer_12663_1 (.in(n12663_0), .out(n12663_1));
wire n12664; //CHANY 4 (1,4) #32
wire n12664_0;
wire n12664_1;
buffer_wire buffer_12664_1 (.in(n12664_0), .out(n12664_1));
wire n12665; //CHANY 4 (1,4) #33
wire n12665_0;
wire n12665_1;
buffer_wire buffer_12665_1 (.in(n12665_0), .out(n12665_1));
wire n12666; //CHANY 4 (1,4) #40
wire n12666_0;
wire n12666_1;
buffer_wire buffer_12666_1 (.in(n12666_0), .out(n12666_1));
wire n12667; //CHANY 4 (1,4) #41
wire n12667_0;
wire n12667_1;
buffer_wire buffer_12667_1 (.in(n12667_0), .out(n12667_1));
wire n12668; //CHANY 4 (1,4) #48
wire n12668_0;
wire n12668_1;
buffer_wire buffer_12668_1 (.in(n12668_0), .out(n12668_1));
wire n12669; //CHANY 4 (1,4) #49
wire n12669_0;
wire n12669_1;
buffer_wire buffer_12669_1 (.in(n12669_0), .out(n12669_1));
wire n12670; //CHANY 4 (1,4) #56
wire n12670_0;
wire n12670_1;
buffer_wire buffer_12670_1 (.in(n12670_0), .out(n12670_1));
wire n12671; //CHANY 4 (1,4) #57
wire n12671_0;
wire n12671_1;
buffer_wire buffer_12671_1 (.in(n12671_0), .out(n12671_1));
wire n12672; //CHANY 4 (1,4) #64
wire n12672_0;
wire n12672_1;
buffer_wire buffer_12672_1 (.in(n12672_0), .out(n12672_1));
wire n12673; //CHANY 4 (1,4) #65
wire n12673_0;
wire n12673_1;
buffer_wire buffer_12673_1 (.in(n12673_0), .out(n12673_1));
wire n12674; //CHANY 4 (1,4) #72
wire n12674_0;
wire n12674_1;
buffer_wire buffer_12674_1 (.in(n12674_0), .out(n12674_1));
wire n12675; //CHANY 4 (1,4) #73
wire n12675_0;
wire n12675_1;
buffer_wire buffer_12675_1 (.in(n12675_0), .out(n12675_1));
wire n12676; //CHANY 4 (1,5) #2
wire n12676_0;
wire n12676_1;
buffer_wire buffer_12676_1 (.in(n12676_0), .out(n12676_1));
wire n12677; //CHANY 4 (1,5) #3
wire n12677_0;
wire n12677_1;
buffer_wire buffer_12677_1 (.in(n12677_0), .out(n12677_1));
wire n12678; //CHANY 4 (1,5) #10
wire n12678_0;
wire n12678_1;
buffer_wire buffer_12678_1 (.in(n12678_0), .out(n12678_1));
wire n12679; //CHANY 4 (1,5) #11
wire n12679_0;
wire n12679_1;
buffer_wire buffer_12679_1 (.in(n12679_0), .out(n12679_1));
wire n12680; //CHANY 4 (1,5) #18
wire n12680_0;
wire n12680_1;
buffer_wire buffer_12680_1 (.in(n12680_0), .out(n12680_1));
wire n12681; //CHANY 4 (1,5) #19
wire n12681_0;
wire n12681_1;
buffer_wire buffer_12681_1 (.in(n12681_0), .out(n12681_1));
wire n12682; //CHANY 4 (1,5) #26
wire n12682_0;
wire n12682_1;
buffer_wire buffer_12682_1 (.in(n12682_0), .out(n12682_1));
wire n12683; //CHANY 4 (1,5) #27
wire n12683_0;
wire n12683_1;
buffer_wire buffer_12683_1 (.in(n12683_0), .out(n12683_1));
wire n12684; //CHANY 4 (1,5) #34
wire n12684_0;
wire n12684_1;
buffer_wire buffer_12684_1 (.in(n12684_0), .out(n12684_1));
wire n12685; //CHANY 4 (1,5) #35
wire n12685_0;
wire n12685_1;
buffer_wire buffer_12685_1 (.in(n12685_0), .out(n12685_1));
wire n12686; //CHANY 4 (1,5) #42
wire n12686_0;
wire n12686_1;
buffer_wire buffer_12686_1 (.in(n12686_0), .out(n12686_1));
wire n12687; //CHANY 4 (1,5) #43
wire n12687_0;
wire n12687_1;
buffer_wire buffer_12687_1 (.in(n12687_0), .out(n12687_1));
wire n12688; //CHANY 4 (1,5) #50
wire n12688_0;
wire n12688_1;
buffer_wire buffer_12688_1 (.in(n12688_0), .out(n12688_1));
wire n12689; //CHANY 4 (1,5) #51
wire n12689_0;
wire n12689_1;
buffer_wire buffer_12689_1 (.in(n12689_0), .out(n12689_1));
wire n12690; //CHANY 4 (1,5) #58
wire n12690_0;
wire n12690_1;
buffer_wire buffer_12690_1 (.in(n12690_0), .out(n12690_1));
wire n12691; //CHANY 4 (1,5) #59
wire n12691_0;
wire n12691_1;
buffer_wire buffer_12691_1 (.in(n12691_0), .out(n12691_1));
wire n12692; //CHANY 4 (1,5) #66
wire n12692_0;
wire n12692_1;
buffer_wire buffer_12692_1 (.in(n12692_0), .out(n12692_1));
wire n12693; //CHANY 4 (1,5) #67
wire n12693_0;
wire n12693_1;
buffer_wire buffer_12693_1 (.in(n12693_0), .out(n12693_1));
wire n12694; //CHANY 4 (1,5) #74
wire n12694_0;
wire n12694_1;
buffer_wire buffer_12694_1 (.in(n12694_0), .out(n12694_1));
wire n12695; //CHANY 4 (1,5) #75
wire n12695_0;
wire n12695_1;
buffer_wire buffer_12695_1 (.in(n12695_0), .out(n12695_1));
wire n12696; //CHANY 4 (1,6) #4
wire n12696_0;
wire n12696_1;
buffer_wire buffer_12696_1 (.in(n12696_0), .out(n12696_1));
wire n12697; //CHANY 4 (1,6) #5
wire n12697_0;
wire n12697_1;
buffer_wire buffer_12697_1 (.in(n12697_0), .out(n12697_1));
wire n12698; //CHANY 4 (1,6) #12
wire n12698_0;
wire n12698_1;
buffer_wire buffer_12698_1 (.in(n12698_0), .out(n12698_1));
wire n12699; //CHANY 4 (1,6) #13
wire n12699_0;
wire n12699_1;
buffer_wire buffer_12699_1 (.in(n12699_0), .out(n12699_1));
wire n12700; //CHANY 4 (1,6) #20
wire n12700_0;
wire n12700_1;
buffer_wire buffer_12700_1 (.in(n12700_0), .out(n12700_1));
wire n12701; //CHANY 4 (1,6) #21
wire n12701_0;
wire n12701_1;
buffer_wire buffer_12701_1 (.in(n12701_0), .out(n12701_1));
wire n12702; //CHANY 4 (1,6) #28
wire n12702_0;
wire n12702_1;
buffer_wire buffer_12702_1 (.in(n12702_0), .out(n12702_1));
wire n12703; //CHANY 4 (1,6) #29
wire n12703_0;
wire n12703_1;
buffer_wire buffer_12703_1 (.in(n12703_0), .out(n12703_1));
wire n12704; //CHANY 4 (1,6) #36
wire n12704_0;
wire n12704_1;
buffer_wire buffer_12704_1 (.in(n12704_0), .out(n12704_1));
wire n12705; //CHANY 4 (1,6) #37
wire n12705_0;
wire n12705_1;
buffer_wire buffer_12705_1 (.in(n12705_0), .out(n12705_1));
wire n12706; //CHANY 4 (1,6) #44
wire n12706_0;
wire n12706_1;
buffer_wire buffer_12706_1 (.in(n12706_0), .out(n12706_1));
wire n12707; //CHANY 4 (1,6) #45
wire n12707_0;
wire n12707_1;
buffer_wire buffer_12707_1 (.in(n12707_0), .out(n12707_1));
wire n12708; //CHANY 4 (1,6) #52
wire n12708_0;
wire n12708_1;
buffer_wire buffer_12708_1 (.in(n12708_0), .out(n12708_1));
wire n12709; //CHANY 4 (1,6) #53
wire n12709_0;
wire n12709_1;
buffer_wire buffer_12709_1 (.in(n12709_0), .out(n12709_1));
wire n12710; //CHANY 4 (1,6) #60
wire n12710_0;
wire n12710_1;
buffer_wire buffer_12710_1 (.in(n12710_0), .out(n12710_1));
wire n12711; //CHANY 4 (1,6) #61
wire n12711_0;
wire n12711_1;
buffer_wire buffer_12711_1 (.in(n12711_0), .out(n12711_1));
wire n12712; //CHANY 4 (1,6) #68
wire n12712_0;
wire n12712_1;
buffer_wire buffer_12712_1 (.in(n12712_0), .out(n12712_1));
wire n12713; //CHANY 4 (1,6) #69
wire n12713_0;
wire n12713_1;
buffer_wire buffer_12713_1 (.in(n12713_0), .out(n12713_1));
wire n12714; //CHANY 4 (1,6) #76
wire n12714_0;
wire n12714_1;
buffer_wire buffer_12714_1 (.in(n12714_0), .out(n12714_1));
wire n12715; //CHANY 4 (1,6) #77
wire n12715_0;
wire n12715_1;
buffer_wire buffer_12715_1 (.in(n12715_0), .out(n12715_1));
wire n12716; //CHANY 3 (1,7) #6
wire n12716_0;
wire n12717; //CHANY 3 (1,7) #7
wire n12717_0;
wire n12718; //CHANY 3 (1,7) #14
wire n12718_0;
wire n12719; //CHANY 3 (1,7) #15
wire n12719_0;
wire n12720; //CHANY 3 (1,7) #22
wire n12720_0;
wire n12721; //CHANY 3 (1,7) #23
wire n12721_0;
wire n12722; //CHANY 3 (1,7) #30
wire n12722_0;
wire n12723; //CHANY 3 (1,7) #31
wire n12723_0;
wire n12724; //CHANY 3 (1,7) #38
wire n12724_0;
wire n12725; //CHANY 3 (1,7) #39
wire n12725_0;
wire n12726; //CHANY 3 (1,7) #46
wire n12726_0;
wire n12727; //CHANY 3 (1,7) #47
wire n12727_0;
wire n12728; //CHANY 3 (1,7) #54
wire n12728_0;
wire n12729; //CHANY 3 (1,7) #55
wire n12729_0;
wire n12730; //CHANY 3 (1,7) #62
wire n12730_0;
wire n12731; //CHANY 3 (1,7) #63
wire n12731_0;
wire n12732; //CHANY 3 (1,7) #70
wire n12732_0;
wire n12733; //CHANY 3 (1,7) #71
wire n12733_0;
wire n12734; //CHANY 3 (1,7) #78
wire n12734_0;
wire n12735; //CHANY 3 (1,7) #79
wire n12735_0;
wire n12736; //CHANY 2 (1,8) #0
wire n12736_0;
wire n12737; //CHANY 2 (1,8) #1
wire n12737_0;
wire n12738; //CHANY 2 (1,8) #8
wire n12738_0;
wire n12739; //CHANY 2 (1,8) #9
wire n12739_0;
wire n12740; //CHANY 2 (1,8) #16
wire n12740_0;
wire n12741; //CHANY 2 (1,8) #17
wire n12741_0;
wire n12742; //CHANY 2 (1,8) #24
wire n12742_0;
wire n12743; //CHANY 2 (1,8) #25
wire n12743_0;
wire n12744; //CHANY 2 (1,8) #32
wire n12744_0;
wire n12745; //CHANY 2 (1,8) #33
wire n12745_0;
wire n12746; //CHANY 2 (1,8) #40
wire n12746_0;
wire n12747; //CHANY 2 (1,8) #41
wire n12747_0;
wire n12748; //CHANY 2 (1,8) #48
wire n12748_0;
wire n12749; //CHANY 2 (1,8) #49
wire n12749_0;
wire n12750; //CHANY 2 (1,8) #56
wire n12750_0;
wire n12751; //CHANY 2 (1,8) #57
wire n12751_0;
wire n12752; //CHANY 2 (1,8) #64
wire n12752_0;
wire n12753; //CHANY 2 (1,8) #65
wire n12753_0;
wire n12754; //CHANY 2 (1,8) #72
wire n12754_0;
wire n12755; //CHANY 2 (1,8) #73
wire n12755_0;
wire n12756; //CHANY 2 (1,8) #80
wire n12756_0;
wire n12757; //CHANY 2 (1,8) #81
wire n12757_0;
wire n12758; //CHANY 1 (1,9) #2
wire n12758_0;
wire n12759; //CHANY 1 (1,9) #3
wire n12759_0;
wire n12760; //CHANY 1 (1,9) #10
wire n12760_0;
wire n12761; //CHANY 1 (1,9) #11
wire n12761_0;
wire n12762; //CHANY 1 (1,9) #18
wire n12762_0;
wire n12763; //CHANY 1 (1,9) #19
wire n12763_0;
wire n12764; //CHANY 1 (1,9) #26
wire n12764_0;
wire n12765; //CHANY 1 (1,9) #27
wire n12765_0;
wire n12766; //CHANY 1 (1,9) #34
wire n12766_0;
wire n12767; //CHANY 1 (1,9) #35
wire n12767_0;
wire n12768; //CHANY 1 (1,9) #42
wire n12768_0;
wire n12769; //CHANY 1 (1,9) #43
wire n12769_0;
wire n12770; //CHANY 1 (1,9) #50
wire n12770_0;
wire n12771; //CHANY 1 (1,9) #51
wire n12771_0;
wire n12772; //CHANY 1 (1,9) #58
wire n12772_0;
wire n12773; //CHANY 1 (1,9) #59
wire n12773_0;
wire n12774; //CHANY 1 (1,9) #66
wire n12774_0;
wire n12775; //CHANY 1 (1,9) #67
wire n12775_0;
wire n12776; //CHANY 1 (1,9) #74
wire n12776_0;
wire n12777; //CHANY 1 (1,9) #75
wire n12777_0;
wire n12778; //CHANY 1 (1,9) #82
wire n12778_0;
wire n12779; //CHANY 1 (1,9) #83
wire n12779_0;
wire n12780; //CHANY 2 (2,1) #0
wire n12780_0;
wire n12781; //CHANY 2 (2,1) #1
wire n12781_0;
wire n12782; //CHANY 3 (2,1) #2
wire n12782_0;
wire n12783; //CHANY 3 (2,1) #3
wire n12783_0;
wire n12784; //CHANY 4 (2,1) #4
wire n12784_0;
wire n12784_1;
buffer_wire buffer_12784_1 (.in(n12784_0), .out(n12784_1));
wire n12785; //CHANY 4 (2,1) #5
wire n12785_0;
wire n12785_1;
buffer_wire buffer_12785_1 (.in(n12785_0), .out(n12785_1));
wire n12786; //CHANY 1 (2,1) #6
wire n12786_0;
wire n12787; //CHANY 1 (2,1) #7
wire n12787_0;
wire n12788; //CHANY 2 (2,1) #8
wire n12788_0;
wire n12789; //CHANY 2 (2,1) #9
wire n12789_0;
wire n12790; //CHANY 3 (2,1) #10
wire n12790_0;
wire n12791; //CHANY 3 (2,1) #11
wire n12791_0;
wire n12792; //CHANY 4 (2,1) #12
wire n12792_0;
wire n12792_1;
buffer_wire buffer_12792_1 (.in(n12792_0), .out(n12792_1));
wire n12793; //CHANY 4 (2,1) #13
wire n12793_0;
wire n12793_1;
buffer_wire buffer_12793_1 (.in(n12793_0), .out(n12793_1));
wire n12794; //CHANY 1 (2,1) #14
wire n12794_0;
wire n12795; //CHANY 1 (2,1) #15
wire n12795_0;
wire n12796; //CHANY 2 (2,1) #16
wire n12796_0;
wire n12797; //CHANY 2 (2,1) #17
wire n12797_0;
wire n12798; //CHANY 3 (2,1) #18
wire n12798_0;
wire n12799; //CHANY 3 (2,1) #19
wire n12799_0;
wire n12800; //CHANY 4 (2,1) #20
wire n12800_0;
wire n12800_1;
buffer_wire buffer_12800_1 (.in(n12800_0), .out(n12800_1));
wire n12801; //CHANY 4 (2,1) #21
wire n12801_0;
wire n12801_1;
buffer_wire buffer_12801_1 (.in(n12801_0), .out(n12801_1));
wire n12802; //CHANY 1 (2,1) #22
wire n12802_0;
wire n12803; //CHANY 1 (2,1) #23
wire n12803_0;
wire n12804; //CHANY 2 (2,1) #24
wire n12804_0;
wire n12805; //CHANY 2 (2,1) #25
wire n12805_0;
wire n12806; //CHANY 3 (2,1) #26
wire n12806_0;
wire n12807; //CHANY 3 (2,1) #27
wire n12807_0;
wire n12808; //CHANY 4 (2,1) #28
wire n12808_0;
wire n12808_1;
buffer_wire buffer_12808_1 (.in(n12808_0), .out(n12808_1));
wire n12809; //CHANY 4 (2,1) #29
wire n12809_0;
wire n12809_1;
buffer_wire buffer_12809_1 (.in(n12809_0), .out(n12809_1));
wire n12810; //CHANY 1 (2,1) #30
wire n12810_0;
wire n12811; //CHANY 1 (2,1) #31
wire n12811_0;
wire n12812; //CHANY 2 (2,1) #32
wire n12812_0;
wire n12813; //CHANY 2 (2,1) #33
wire n12813_0;
wire n12814; //CHANY 3 (2,1) #34
wire n12814_0;
wire n12815; //CHANY 3 (2,1) #35
wire n12815_0;
wire n12816; //CHANY 4 (2,1) #36
wire n12816_0;
wire n12816_1;
buffer_wire buffer_12816_1 (.in(n12816_0), .out(n12816_1));
wire n12817; //CHANY 4 (2,1) #37
wire n12817_0;
wire n12817_1;
buffer_wire buffer_12817_1 (.in(n12817_0), .out(n12817_1));
wire n12818; //CHANY 1 (2,1) #38
wire n12818_0;
wire n12819; //CHANY 1 (2,1) #39
wire n12819_0;
wire n12820; //CHANY 2 (2,1) #40
wire n12820_0;
wire n12821; //CHANY 2 (2,1) #41
wire n12821_0;
wire n12822; //CHANY 3 (2,1) #42
wire n12822_0;
wire n12823; //CHANY 3 (2,1) #43
wire n12823_0;
wire n12824; //CHANY 4 (2,1) #44
wire n12824_0;
wire n12824_1;
buffer_wire buffer_12824_1 (.in(n12824_0), .out(n12824_1));
wire n12825; //CHANY 4 (2,1) #45
wire n12825_0;
wire n12825_1;
buffer_wire buffer_12825_1 (.in(n12825_0), .out(n12825_1));
wire n12826; //CHANY 1 (2,1) #46
wire n12826_0;
wire n12827; //CHANY 1 (2,1) #47
wire n12827_0;
wire n12828; //CHANY 2 (2,1) #48
wire n12828_0;
wire n12829; //CHANY 2 (2,1) #49
wire n12829_0;
wire n12830; //CHANY 3 (2,1) #50
wire n12830_0;
wire n12831; //CHANY 3 (2,1) #51
wire n12831_0;
wire n12832; //CHANY 4 (2,1) #52
wire n12832_0;
wire n12832_1;
buffer_wire buffer_12832_1 (.in(n12832_0), .out(n12832_1));
wire n12833; //CHANY 4 (2,1) #53
wire n12833_0;
wire n12833_1;
buffer_wire buffer_12833_1 (.in(n12833_0), .out(n12833_1));
wire n12834; //CHANY 1 (2,1) #54
wire n12834_0;
wire n12835; //CHANY 1 (2,1) #55
wire n12835_0;
wire n12836; //CHANY 2 (2,1) #56
wire n12836_0;
wire n12837; //CHANY 2 (2,1) #57
wire n12837_0;
wire n12838; //CHANY 3 (2,1) #58
wire n12838_0;
wire n12839; //CHANY 3 (2,1) #59
wire n12839_0;
wire n12840; //CHANY 4 (2,1) #60
wire n12840_0;
wire n12840_1;
buffer_wire buffer_12840_1 (.in(n12840_0), .out(n12840_1));
wire n12841; //CHANY 4 (2,1) #61
wire n12841_0;
wire n12841_1;
buffer_wire buffer_12841_1 (.in(n12841_0), .out(n12841_1));
wire n12842; //CHANY 1 (2,1) #62
wire n12842_0;
wire n12843; //CHANY 1 (2,1) #63
wire n12843_0;
wire n12844; //CHANY 2 (2,1) #64
wire n12844_0;
wire n12845; //CHANY 2 (2,1) #65
wire n12845_0;
wire n12846; //CHANY 3 (2,1) #66
wire n12846_0;
wire n12847; //CHANY 3 (2,1) #67
wire n12847_0;
wire n12848; //CHANY 4 (2,1) #68
wire n12848_0;
wire n12848_1;
buffer_wire buffer_12848_1 (.in(n12848_0), .out(n12848_1));
wire n12849; //CHANY 4 (2,1) #69
wire n12849_0;
wire n12849_1;
buffer_wire buffer_12849_1 (.in(n12849_0), .out(n12849_1));
wire n12850; //CHANY 1 (2,1) #70
wire n12850_0;
wire n12851; //CHANY 1 (2,1) #71
wire n12851_0;
wire n12852; //CHANY 2 (2,1) #72
wire n12852_0;
wire n12853; //CHANY 2 (2,1) #73
wire n12853_0;
wire n12854; //CHANY 3 (2,1) #74
wire n12854_0;
wire n12855; //CHANY 3 (2,1) #75
wire n12855_0;
wire n12856; //CHANY 4 (2,1) #76
wire n12856_0;
wire n12856_1;
buffer_wire buffer_12856_1 (.in(n12856_0), .out(n12856_1));
wire n12857; //CHANY 4 (2,1) #77
wire n12857_0;
wire n12857_1;
buffer_wire buffer_12857_1 (.in(n12857_0), .out(n12857_1));
wire n12858; //CHANY 1 (2,1) #78
wire n12858_0;
wire n12859; //CHANY 1 (2,1) #79
wire n12859_0;
wire n12860; //CHANY 6 (2,1) #80
wire n12860_0;
wire n12860_1;
buffer_wire buffer_12860_1 (.in(n12860_0), .out(n12860_1));
wire n12861; //CHANY 6 (2,1) #81
wire n12861_0;
wire n12861_1;
buffer_wire buffer_12861_1 (.in(n12861_0), .out(n12861_1));
wire n12862; //CHANY 7 (2,1) #82
wire n12862_0;
wire n12862_1;
wire n12862_2;
buffer_wire buffer_12862_2 (.in(n12862_1), .out(n12862_2));
buffer_wire buffer_12862_1 (.in(n12862_0), .out(n12862_1));
wire n12863; //CHANY 7 (2,1) #83
wire n12863_0;
wire n12863_1;
wire n12863_2;
buffer_wire buffer_12863_2 (.in(n12863_1), .out(n12863_2));
buffer_wire buffer_12863_1 (.in(n12863_0), .out(n12863_1));
wire n12864; //CHANY 8 (2,1) #84
wire n12864_0;
wire n12864_1;
wire n12864_2;
buffer_wire buffer_12864_2 (.in(n12864_1), .out(n12864_2));
buffer_wire buffer_12864_1 (.in(n12864_0), .out(n12864_1));
wire n12865; //CHANY 8 (2,1) #85
wire n12865_0;
wire n12865_1;
wire n12865_2;
buffer_wire buffer_12865_2 (.in(n12865_1), .out(n12865_2));
buffer_wire buffer_12865_1 (.in(n12865_0), .out(n12865_1));
wire n12866; //CHANY 9 (2,1) #86
wire n12866_0;
wire n12866_1;
wire n12866_2;
buffer_wire buffer_12866_2 (.in(n12866_1), .out(n12866_2));
buffer_wire buffer_12866_1 (.in(n12866_0), .out(n12866_1));
wire n12867; //CHANY 9 (2,1) #87
wire n12867_0;
wire n12867_1;
wire n12867_2;
buffer_wire buffer_12867_2 (.in(n12867_1), .out(n12867_2));
buffer_wire buffer_12867_1 (.in(n12867_0), .out(n12867_1));
wire n12868; //CHANY 9 (2,1) #88
wire n12868_0;
wire n12868_1;
wire n12868_2;
buffer_wire buffer_12868_2 (.in(n12868_1), .out(n12868_2));
buffer_wire buffer_12868_1 (.in(n12868_0), .out(n12868_1));
wire n12869; //CHANY 9 (2,1) #89
wire n12869_0;
wire n12869_1;
wire n12869_2;
buffer_wire buffer_12869_2 (.in(n12869_1), .out(n12869_2));
buffer_wire buffer_12869_1 (.in(n12869_0), .out(n12869_1));
wire n12870; //CHANY 9 (2,1) #90
wire n12870_0;
wire n12870_1;
wire n12870_2;
buffer_wire buffer_12870_2 (.in(n12870_1), .out(n12870_2));
buffer_wire buffer_12870_1 (.in(n12870_0), .out(n12870_1));
wire n12871; //CHANY 9 (2,1) #91
wire n12871_0;
wire n12871_1;
wire n12871_2;
buffer_wire buffer_12871_2 (.in(n12871_1), .out(n12871_2));
buffer_wire buffer_12871_1 (.in(n12871_0), .out(n12871_1));
wire n12872; //CHANY 4 (2,2) #6
wire n12872_0;
wire n12872_1;
buffer_wire buffer_12872_1 (.in(n12872_0), .out(n12872_1));
wire n12873; //CHANY 4 (2,2) #7
wire n12873_0;
wire n12873_1;
buffer_wire buffer_12873_1 (.in(n12873_0), .out(n12873_1));
wire n12874; //CHANY 4 (2,2) #14
wire n12874_0;
wire n12874_1;
buffer_wire buffer_12874_1 (.in(n12874_0), .out(n12874_1));
wire n12875; //CHANY 4 (2,2) #15
wire n12875_0;
wire n12875_1;
buffer_wire buffer_12875_1 (.in(n12875_0), .out(n12875_1));
wire n12876; //CHANY 4 (2,2) #22
wire n12876_0;
wire n12876_1;
buffer_wire buffer_12876_1 (.in(n12876_0), .out(n12876_1));
wire n12877; //CHANY 4 (2,2) #23
wire n12877_0;
wire n12877_1;
buffer_wire buffer_12877_1 (.in(n12877_0), .out(n12877_1));
wire n12878; //CHANY 4 (2,2) #30
wire n12878_0;
wire n12878_1;
buffer_wire buffer_12878_1 (.in(n12878_0), .out(n12878_1));
wire n12879; //CHANY 4 (2,2) #31
wire n12879_0;
wire n12879_1;
buffer_wire buffer_12879_1 (.in(n12879_0), .out(n12879_1));
wire n12880; //CHANY 4 (2,2) #38
wire n12880_0;
wire n12880_1;
buffer_wire buffer_12880_1 (.in(n12880_0), .out(n12880_1));
wire n12881; //CHANY 4 (2,2) #39
wire n12881_0;
wire n12881_1;
buffer_wire buffer_12881_1 (.in(n12881_0), .out(n12881_1));
wire n12882; //CHANY 4 (2,2) #46
wire n12882_0;
wire n12882_1;
buffer_wire buffer_12882_1 (.in(n12882_0), .out(n12882_1));
wire n12883; //CHANY 4 (2,2) #47
wire n12883_0;
wire n12883_1;
buffer_wire buffer_12883_1 (.in(n12883_0), .out(n12883_1));
wire n12884; //CHANY 4 (2,2) #54
wire n12884_0;
wire n12884_1;
buffer_wire buffer_12884_1 (.in(n12884_0), .out(n12884_1));
wire n12885; //CHANY 4 (2,2) #55
wire n12885_0;
wire n12885_1;
buffer_wire buffer_12885_1 (.in(n12885_0), .out(n12885_1));
wire n12886; //CHANY 4 (2,2) #62
wire n12886_0;
wire n12886_1;
buffer_wire buffer_12886_1 (.in(n12886_0), .out(n12886_1));
wire n12887; //CHANY 4 (2,2) #63
wire n12887_0;
wire n12887_1;
buffer_wire buffer_12887_1 (.in(n12887_0), .out(n12887_1));
wire n12888; //CHANY 4 (2,2) #70
wire n12888_0;
wire n12888_1;
buffer_wire buffer_12888_1 (.in(n12888_0), .out(n12888_1));
wire n12889; //CHANY 4 (2,2) #71
wire n12889_0;
wire n12889_1;
buffer_wire buffer_12889_1 (.in(n12889_0), .out(n12889_1));
wire n12890; //CHANY 4 (2,2) #78
wire n12890_0;
wire n12890_1;
buffer_wire buffer_12890_1 (.in(n12890_0), .out(n12890_1));
wire n12891; //CHANY 4 (2,2) #79
wire n12891_0;
wire n12891_1;
buffer_wire buffer_12891_1 (.in(n12891_0), .out(n12891_1));
wire n12892; //CHANY 4 (2,3) #0
wire n12892_0;
wire n12892_1;
buffer_wire buffer_12892_1 (.in(n12892_0), .out(n12892_1));
wire n12893; //CHANY 4 (2,3) #1
wire n12893_0;
wire n12893_1;
buffer_wire buffer_12893_1 (.in(n12893_0), .out(n12893_1));
wire n12894; //CHANY 4 (2,3) #8
wire n12894_0;
wire n12894_1;
buffer_wire buffer_12894_1 (.in(n12894_0), .out(n12894_1));
wire n12895; //CHANY 4 (2,3) #9
wire n12895_0;
wire n12895_1;
buffer_wire buffer_12895_1 (.in(n12895_0), .out(n12895_1));
wire n12896; //CHANY 4 (2,3) #16
wire n12896_0;
wire n12896_1;
buffer_wire buffer_12896_1 (.in(n12896_0), .out(n12896_1));
wire n12897; //CHANY 4 (2,3) #17
wire n12897_0;
wire n12897_1;
buffer_wire buffer_12897_1 (.in(n12897_0), .out(n12897_1));
wire n12898; //CHANY 4 (2,3) #24
wire n12898_0;
wire n12898_1;
buffer_wire buffer_12898_1 (.in(n12898_0), .out(n12898_1));
wire n12899; //CHANY 4 (2,3) #25
wire n12899_0;
wire n12899_1;
buffer_wire buffer_12899_1 (.in(n12899_0), .out(n12899_1));
wire n12900; //CHANY 4 (2,3) #32
wire n12900_0;
wire n12900_1;
buffer_wire buffer_12900_1 (.in(n12900_0), .out(n12900_1));
wire n12901; //CHANY 4 (2,3) #33
wire n12901_0;
wire n12901_1;
buffer_wire buffer_12901_1 (.in(n12901_0), .out(n12901_1));
wire n12902; //CHANY 4 (2,3) #40
wire n12902_0;
wire n12902_1;
buffer_wire buffer_12902_1 (.in(n12902_0), .out(n12902_1));
wire n12903; //CHANY 4 (2,3) #41
wire n12903_0;
wire n12903_1;
buffer_wire buffer_12903_1 (.in(n12903_0), .out(n12903_1));
wire n12904; //CHANY 4 (2,3) #48
wire n12904_0;
wire n12904_1;
buffer_wire buffer_12904_1 (.in(n12904_0), .out(n12904_1));
wire n12905; //CHANY 4 (2,3) #49
wire n12905_0;
wire n12905_1;
buffer_wire buffer_12905_1 (.in(n12905_0), .out(n12905_1));
wire n12906; //CHANY 4 (2,3) #56
wire n12906_0;
wire n12906_1;
buffer_wire buffer_12906_1 (.in(n12906_0), .out(n12906_1));
wire n12907; //CHANY 4 (2,3) #57
wire n12907_0;
wire n12907_1;
buffer_wire buffer_12907_1 (.in(n12907_0), .out(n12907_1));
wire n12908; //CHANY 4 (2,3) #64
wire n12908_0;
wire n12908_1;
buffer_wire buffer_12908_1 (.in(n12908_0), .out(n12908_1));
wire n12909; //CHANY 4 (2,3) #65
wire n12909_0;
wire n12909_1;
buffer_wire buffer_12909_1 (.in(n12909_0), .out(n12909_1));
wire n12910; //CHANY 4 (2,3) #72
wire n12910_0;
wire n12910_1;
buffer_wire buffer_12910_1 (.in(n12910_0), .out(n12910_1));
wire n12911; //CHANY 4 (2,3) #73
wire n12911_0;
wire n12911_1;
buffer_wire buffer_12911_1 (.in(n12911_0), .out(n12911_1));
wire n12912; //CHANY 4 (2,4) #2
wire n12912_0;
wire n12912_1;
buffer_wire buffer_12912_1 (.in(n12912_0), .out(n12912_1));
wire n12913; //CHANY 4 (2,4) #3
wire n12913_0;
wire n12913_1;
buffer_wire buffer_12913_1 (.in(n12913_0), .out(n12913_1));
wire n12914; //CHANY 4 (2,4) #10
wire n12914_0;
wire n12914_1;
buffer_wire buffer_12914_1 (.in(n12914_0), .out(n12914_1));
wire n12915; //CHANY 4 (2,4) #11
wire n12915_0;
wire n12915_1;
buffer_wire buffer_12915_1 (.in(n12915_0), .out(n12915_1));
wire n12916; //CHANY 4 (2,4) #18
wire n12916_0;
wire n12916_1;
buffer_wire buffer_12916_1 (.in(n12916_0), .out(n12916_1));
wire n12917; //CHANY 4 (2,4) #19
wire n12917_0;
wire n12917_1;
buffer_wire buffer_12917_1 (.in(n12917_0), .out(n12917_1));
wire n12918; //CHANY 4 (2,4) #26
wire n12918_0;
wire n12918_1;
buffer_wire buffer_12918_1 (.in(n12918_0), .out(n12918_1));
wire n12919; //CHANY 4 (2,4) #27
wire n12919_0;
wire n12919_1;
buffer_wire buffer_12919_1 (.in(n12919_0), .out(n12919_1));
wire n12920; //CHANY 4 (2,4) #34
wire n12920_0;
wire n12920_1;
buffer_wire buffer_12920_1 (.in(n12920_0), .out(n12920_1));
wire n12921; //CHANY 4 (2,4) #35
wire n12921_0;
wire n12921_1;
buffer_wire buffer_12921_1 (.in(n12921_0), .out(n12921_1));
wire n12922; //CHANY 4 (2,4) #42
wire n12922_0;
wire n12922_1;
buffer_wire buffer_12922_1 (.in(n12922_0), .out(n12922_1));
wire n12923; //CHANY 4 (2,4) #43
wire n12923_0;
wire n12923_1;
buffer_wire buffer_12923_1 (.in(n12923_0), .out(n12923_1));
wire n12924; //CHANY 4 (2,4) #50
wire n12924_0;
wire n12924_1;
buffer_wire buffer_12924_1 (.in(n12924_0), .out(n12924_1));
wire n12925; //CHANY 4 (2,4) #51
wire n12925_0;
wire n12925_1;
buffer_wire buffer_12925_1 (.in(n12925_0), .out(n12925_1));
wire n12926; //CHANY 4 (2,4) #58
wire n12926_0;
wire n12926_1;
buffer_wire buffer_12926_1 (.in(n12926_0), .out(n12926_1));
wire n12927; //CHANY 4 (2,4) #59
wire n12927_0;
wire n12927_1;
buffer_wire buffer_12927_1 (.in(n12927_0), .out(n12927_1));
wire n12928; //CHANY 4 (2,4) #66
wire n12928_0;
wire n12928_1;
buffer_wire buffer_12928_1 (.in(n12928_0), .out(n12928_1));
wire n12929; //CHANY 4 (2,4) #67
wire n12929_0;
wire n12929_1;
buffer_wire buffer_12929_1 (.in(n12929_0), .out(n12929_1));
wire n12930; //CHANY 4 (2,4) #74
wire n12930_0;
wire n12930_1;
buffer_wire buffer_12930_1 (.in(n12930_0), .out(n12930_1));
wire n12931; //CHANY 4 (2,4) #75
wire n12931_0;
wire n12931_1;
buffer_wire buffer_12931_1 (.in(n12931_0), .out(n12931_1));
wire n12932; //CHANY 4 (2,5) #4
wire n12932_0;
wire n12932_1;
buffer_wire buffer_12932_1 (.in(n12932_0), .out(n12932_1));
wire n12933; //CHANY 4 (2,5) #5
wire n12933_0;
wire n12933_1;
buffer_wire buffer_12933_1 (.in(n12933_0), .out(n12933_1));
wire n12934; //CHANY 4 (2,5) #12
wire n12934_0;
wire n12934_1;
buffer_wire buffer_12934_1 (.in(n12934_0), .out(n12934_1));
wire n12935; //CHANY 4 (2,5) #13
wire n12935_0;
wire n12935_1;
buffer_wire buffer_12935_1 (.in(n12935_0), .out(n12935_1));
wire n12936; //CHANY 4 (2,5) #20
wire n12936_0;
wire n12936_1;
buffer_wire buffer_12936_1 (.in(n12936_0), .out(n12936_1));
wire n12937; //CHANY 4 (2,5) #21
wire n12937_0;
wire n12937_1;
buffer_wire buffer_12937_1 (.in(n12937_0), .out(n12937_1));
wire n12938; //CHANY 4 (2,5) #28
wire n12938_0;
wire n12938_1;
buffer_wire buffer_12938_1 (.in(n12938_0), .out(n12938_1));
wire n12939; //CHANY 4 (2,5) #29
wire n12939_0;
wire n12939_1;
buffer_wire buffer_12939_1 (.in(n12939_0), .out(n12939_1));
wire n12940; //CHANY 4 (2,5) #36
wire n12940_0;
wire n12940_1;
buffer_wire buffer_12940_1 (.in(n12940_0), .out(n12940_1));
wire n12941; //CHANY 4 (2,5) #37
wire n12941_0;
wire n12941_1;
buffer_wire buffer_12941_1 (.in(n12941_0), .out(n12941_1));
wire n12942; //CHANY 4 (2,5) #44
wire n12942_0;
wire n12942_1;
buffer_wire buffer_12942_1 (.in(n12942_0), .out(n12942_1));
wire n12943; //CHANY 4 (2,5) #45
wire n12943_0;
wire n12943_1;
buffer_wire buffer_12943_1 (.in(n12943_0), .out(n12943_1));
wire n12944; //CHANY 4 (2,5) #52
wire n12944_0;
wire n12944_1;
buffer_wire buffer_12944_1 (.in(n12944_0), .out(n12944_1));
wire n12945; //CHANY 4 (2,5) #53
wire n12945_0;
wire n12945_1;
buffer_wire buffer_12945_1 (.in(n12945_0), .out(n12945_1));
wire n12946; //CHANY 4 (2,5) #60
wire n12946_0;
wire n12946_1;
buffer_wire buffer_12946_1 (.in(n12946_0), .out(n12946_1));
wire n12947; //CHANY 4 (2,5) #61
wire n12947_0;
wire n12947_1;
buffer_wire buffer_12947_1 (.in(n12947_0), .out(n12947_1));
wire n12948; //CHANY 4 (2,5) #68
wire n12948_0;
wire n12948_1;
buffer_wire buffer_12948_1 (.in(n12948_0), .out(n12948_1));
wire n12949; //CHANY 4 (2,5) #69
wire n12949_0;
wire n12949_1;
buffer_wire buffer_12949_1 (.in(n12949_0), .out(n12949_1));
wire n12950; //CHANY 4 (2,5) #76
wire n12950_0;
wire n12950_1;
buffer_wire buffer_12950_1 (.in(n12950_0), .out(n12950_1));
wire n12951; //CHANY 4 (2,5) #77
wire n12951_0;
wire n12951_1;
buffer_wire buffer_12951_1 (.in(n12951_0), .out(n12951_1));
wire n12952; //CHANY 4 (2,6) #6
wire n12952_0;
wire n12952_1;
buffer_wire buffer_12952_1 (.in(n12952_0), .out(n12952_1));
wire n12953; //CHANY 4 (2,6) #7
wire n12953_0;
wire n12953_1;
buffer_wire buffer_12953_1 (.in(n12953_0), .out(n12953_1));
wire n12954; //CHANY 4 (2,6) #14
wire n12954_0;
wire n12954_1;
buffer_wire buffer_12954_1 (.in(n12954_0), .out(n12954_1));
wire n12955; //CHANY 4 (2,6) #15
wire n12955_0;
wire n12955_1;
buffer_wire buffer_12955_1 (.in(n12955_0), .out(n12955_1));
wire n12956; //CHANY 4 (2,6) #22
wire n12956_0;
wire n12956_1;
buffer_wire buffer_12956_1 (.in(n12956_0), .out(n12956_1));
wire n12957; //CHANY 4 (2,6) #23
wire n12957_0;
wire n12957_1;
buffer_wire buffer_12957_1 (.in(n12957_0), .out(n12957_1));
wire n12958; //CHANY 4 (2,6) #30
wire n12958_0;
wire n12958_1;
buffer_wire buffer_12958_1 (.in(n12958_0), .out(n12958_1));
wire n12959; //CHANY 4 (2,6) #31
wire n12959_0;
wire n12959_1;
buffer_wire buffer_12959_1 (.in(n12959_0), .out(n12959_1));
wire n12960; //CHANY 4 (2,6) #38
wire n12960_0;
wire n12960_1;
buffer_wire buffer_12960_1 (.in(n12960_0), .out(n12960_1));
wire n12961; //CHANY 4 (2,6) #39
wire n12961_0;
wire n12961_1;
buffer_wire buffer_12961_1 (.in(n12961_0), .out(n12961_1));
wire n12962; //CHANY 4 (2,6) #46
wire n12962_0;
wire n12962_1;
buffer_wire buffer_12962_1 (.in(n12962_0), .out(n12962_1));
wire n12963; //CHANY 4 (2,6) #47
wire n12963_0;
wire n12963_1;
buffer_wire buffer_12963_1 (.in(n12963_0), .out(n12963_1));
wire n12964; //CHANY 4 (2,6) #54
wire n12964_0;
wire n12964_1;
buffer_wire buffer_12964_1 (.in(n12964_0), .out(n12964_1));
wire n12965; //CHANY 4 (2,6) #55
wire n12965_0;
wire n12965_1;
buffer_wire buffer_12965_1 (.in(n12965_0), .out(n12965_1));
wire n12966; //CHANY 4 (2,6) #62
wire n12966_0;
wire n12966_1;
buffer_wire buffer_12966_1 (.in(n12966_0), .out(n12966_1));
wire n12967; //CHANY 4 (2,6) #63
wire n12967_0;
wire n12967_1;
buffer_wire buffer_12967_1 (.in(n12967_0), .out(n12967_1));
wire n12968; //CHANY 4 (2,6) #70
wire n12968_0;
wire n12968_1;
buffer_wire buffer_12968_1 (.in(n12968_0), .out(n12968_1));
wire n12969; //CHANY 4 (2,6) #71
wire n12969_0;
wire n12969_1;
buffer_wire buffer_12969_1 (.in(n12969_0), .out(n12969_1));
wire n12970; //CHANY 4 (2,6) #78
wire n12970_0;
wire n12970_1;
buffer_wire buffer_12970_1 (.in(n12970_0), .out(n12970_1));
wire n12971; //CHANY 4 (2,6) #79
wire n12971_0;
wire n12971_1;
buffer_wire buffer_12971_1 (.in(n12971_0), .out(n12971_1));
wire n12972; //CHANY 3 (2,7) #0
wire n12972_0;
wire n12973; //CHANY 3 (2,7) #1
wire n12973_0;
wire n12974; //CHANY 3 (2,7) #8
wire n12974_0;
wire n12975; //CHANY 3 (2,7) #9
wire n12975_0;
wire n12976; //CHANY 3 (2,7) #16
wire n12976_0;
wire n12977; //CHANY 3 (2,7) #17
wire n12977_0;
wire n12978; //CHANY 3 (2,7) #24
wire n12978_0;
wire n12979; //CHANY 3 (2,7) #25
wire n12979_0;
wire n12980; //CHANY 3 (2,7) #32
wire n12980_0;
wire n12981; //CHANY 3 (2,7) #33
wire n12981_0;
wire n12982; //CHANY 3 (2,7) #40
wire n12982_0;
wire n12983; //CHANY 3 (2,7) #41
wire n12983_0;
wire n12984; //CHANY 3 (2,7) #48
wire n12984_0;
wire n12985; //CHANY 3 (2,7) #49
wire n12985_0;
wire n12986; //CHANY 3 (2,7) #56
wire n12986_0;
wire n12987; //CHANY 3 (2,7) #57
wire n12987_0;
wire n12988; //CHANY 3 (2,7) #64
wire n12988_0;
wire n12989; //CHANY 3 (2,7) #65
wire n12989_0;
wire n12990; //CHANY 3 (2,7) #72
wire n12990_0;
wire n12991; //CHANY 3 (2,7) #73
wire n12991_0;
wire n12992; //CHANY 3 (2,7) #80
wire n12992_0;
wire n12993; //CHANY 3 (2,7) #81
wire n12993_0;
wire n12994; //CHANY 2 (2,8) #2
wire n12994_0;
wire n12995; //CHANY 2 (2,8) #3
wire n12995_0;
wire n12996; //CHANY 2 (2,8) #10
wire n12996_0;
wire n12997; //CHANY 2 (2,8) #11
wire n12997_0;
wire n12998; //CHANY 2 (2,8) #18
wire n12998_0;
wire n12999; //CHANY 2 (2,8) #19
wire n12999_0;
wire n13000; //CHANY 2 (2,8) #26
wire n13000_0;
wire n13001; //CHANY 2 (2,8) #27
wire n13001_0;
wire n13002; //CHANY 2 (2,8) #34
wire n13002_0;
wire n13003; //CHANY 2 (2,8) #35
wire n13003_0;
wire n13004; //CHANY 2 (2,8) #42
wire n13004_0;
wire n13005; //CHANY 2 (2,8) #43
wire n13005_0;
wire n13006; //CHANY 2 (2,8) #50
wire n13006_0;
wire n13007; //CHANY 2 (2,8) #51
wire n13007_0;
wire n13008; //CHANY 2 (2,8) #58
wire n13008_0;
wire n13009; //CHANY 2 (2,8) #59
wire n13009_0;
wire n13010; //CHANY 2 (2,8) #66
wire n13010_0;
wire n13011; //CHANY 2 (2,8) #67
wire n13011_0;
wire n13012; //CHANY 2 (2,8) #74
wire n13012_0;
wire n13013; //CHANY 2 (2,8) #75
wire n13013_0;
wire n13014; //CHANY 2 (2,8) #82
wire n13014_0;
wire n13015; //CHANY 2 (2,8) #83
wire n13015_0;
wire n13016; //CHANY 1 (2,9) #4
wire n13016_0;
wire n13017; //CHANY 1 (2,9) #5
wire n13017_0;
wire n13018; //CHANY 1 (2,9) #12
wire n13018_0;
wire n13019; //CHANY 1 (2,9) #13
wire n13019_0;
wire n13020; //CHANY 1 (2,9) #20
wire n13020_0;
wire n13021; //CHANY 1 (2,9) #21
wire n13021_0;
wire n13022; //CHANY 1 (2,9) #28
wire n13022_0;
wire n13023; //CHANY 1 (2,9) #29
wire n13023_0;
wire n13024; //CHANY 1 (2,9) #36
wire n13024_0;
wire n13025; //CHANY 1 (2,9) #37
wire n13025_0;
wire n13026; //CHANY 1 (2,9) #44
wire n13026_0;
wire n13027; //CHANY 1 (2,9) #45
wire n13027_0;
wire n13028; //CHANY 1 (2,9) #52
wire n13028_0;
wire n13029; //CHANY 1 (2,9) #53
wire n13029_0;
wire n13030; //CHANY 1 (2,9) #60
wire n13030_0;
wire n13031; //CHANY 1 (2,9) #61
wire n13031_0;
wire n13032; //CHANY 1 (2,9) #68
wire n13032_0;
wire n13033; //CHANY 1 (2,9) #69
wire n13033_0;
wire n13034; //CHANY 1 (2,9) #76
wire n13034_0;
wire n13035; //CHANY 1 (2,9) #77
wire n13035_0;
wire n13036; //CHANY 1 (2,9) #84
wire n13036_0;
wire n13037; //CHANY 1 (2,9) #85
wire n13037_0;
wire n13038; //CHANY 1 (3,1) #0
wire n13038_0;
wire n13039; //CHANY 1 (3,1) #1
wire n13039_0;
wire n13040; //CHANY 2 (3,1) #2
wire n13040_0;
wire n13041; //CHANY 2 (3,1) #3
wire n13041_0;
wire n13042; //CHANY 3 (3,1) #4
wire n13042_0;
wire n13043; //CHANY 3 (3,1) #5
wire n13043_0;
wire n13044; //CHANY 4 (3,1) #6
wire n13044_0;
wire n13044_1;
buffer_wire buffer_13044_1 (.in(n13044_0), .out(n13044_1));
wire n13045; //CHANY 4 (3,1) #7
wire n13045_0;
wire n13045_1;
buffer_wire buffer_13045_1 (.in(n13045_0), .out(n13045_1));
wire n13046; //CHANY 1 (3,1) #8
wire n13046_0;
wire n13047; //CHANY 1 (3,1) #9
wire n13047_0;
wire n13048; //CHANY 2 (3,1) #10
wire n13048_0;
wire n13049; //CHANY 2 (3,1) #11
wire n13049_0;
wire n13050; //CHANY 3 (3,1) #12
wire n13050_0;
wire n13051; //CHANY 3 (3,1) #13
wire n13051_0;
wire n13052; //CHANY 4 (3,1) #14
wire n13052_0;
wire n13052_1;
buffer_wire buffer_13052_1 (.in(n13052_0), .out(n13052_1));
wire n13053; //CHANY 4 (3,1) #15
wire n13053_0;
wire n13053_1;
buffer_wire buffer_13053_1 (.in(n13053_0), .out(n13053_1));
wire n13054; //CHANY 1 (3,1) #16
wire n13054_0;
wire n13055; //CHANY 1 (3,1) #17
wire n13055_0;
wire n13056; //CHANY 2 (3,1) #18
wire n13056_0;
wire n13057; //CHANY 2 (3,1) #19
wire n13057_0;
wire n13058; //CHANY 3 (3,1) #20
wire n13058_0;
wire n13059; //CHANY 3 (3,1) #21
wire n13059_0;
wire n13060; //CHANY 4 (3,1) #22
wire n13060_0;
wire n13060_1;
buffer_wire buffer_13060_1 (.in(n13060_0), .out(n13060_1));
wire n13061; //CHANY 4 (3,1) #23
wire n13061_0;
wire n13061_1;
buffer_wire buffer_13061_1 (.in(n13061_0), .out(n13061_1));
wire n13062; //CHANY 1 (3,1) #24
wire n13062_0;
wire n13063; //CHANY 1 (3,1) #25
wire n13063_0;
wire n13064; //CHANY 2 (3,1) #26
wire n13064_0;
wire n13065; //CHANY 2 (3,1) #27
wire n13065_0;
wire n13066; //CHANY 3 (3,1) #28
wire n13066_0;
wire n13067; //CHANY 3 (3,1) #29
wire n13067_0;
wire n13068; //CHANY 4 (3,1) #30
wire n13068_0;
wire n13068_1;
buffer_wire buffer_13068_1 (.in(n13068_0), .out(n13068_1));
wire n13069; //CHANY 4 (3,1) #31
wire n13069_0;
wire n13069_1;
buffer_wire buffer_13069_1 (.in(n13069_0), .out(n13069_1));
wire n13070; //CHANY 1 (3,1) #32
wire n13070_0;
wire n13071; //CHANY 1 (3,1) #33
wire n13071_0;
wire n13072; //CHANY 2 (3,1) #34
wire n13072_0;
wire n13073; //CHANY 2 (3,1) #35
wire n13073_0;
wire n13074; //CHANY 3 (3,1) #36
wire n13074_0;
wire n13075; //CHANY 3 (3,1) #37
wire n13075_0;
wire n13076; //CHANY 4 (3,1) #38
wire n13076_0;
wire n13076_1;
buffer_wire buffer_13076_1 (.in(n13076_0), .out(n13076_1));
wire n13077; //CHANY 4 (3,1) #39
wire n13077_0;
wire n13077_1;
buffer_wire buffer_13077_1 (.in(n13077_0), .out(n13077_1));
wire n13078; //CHANY 1 (3,1) #40
wire n13078_0;
wire n13079; //CHANY 1 (3,1) #41
wire n13079_0;
wire n13080; //CHANY 2 (3,1) #42
wire n13080_0;
wire n13081; //CHANY 2 (3,1) #43
wire n13081_0;
wire n13082; //CHANY 3 (3,1) #44
wire n13082_0;
wire n13083; //CHANY 3 (3,1) #45
wire n13083_0;
wire n13084; //CHANY 4 (3,1) #46
wire n13084_0;
wire n13084_1;
buffer_wire buffer_13084_1 (.in(n13084_0), .out(n13084_1));
wire n13085; //CHANY 4 (3,1) #47
wire n13085_0;
wire n13085_1;
buffer_wire buffer_13085_1 (.in(n13085_0), .out(n13085_1));
wire n13086; //CHANY 1 (3,1) #48
wire n13086_0;
wire n13087; //CHANY 1 (3,1) #49
wire n13087_0;
wire n13088; //CHANY 2 (3,1) #50
wire n13088_0;
wire n13089; //CHANY 2 (3,1) #51
wire n13089_0;
wire n13090; //CHANY 3 (3,1) #52
wire n13090_0;
wire n13091; //CHANY 3 (3,1) #53
wire n13091_0;
wire n13092; //CHANY 4 (3,1) #54
wire n13092_0;
wire n13092_1;
buffer_wire buffer_13092_1 (.in(n13092_0), .out(n13092_1));
wire n13093; //CHANY 4 (3,1) #55
wire n13093_0;
wire n13093_1;
buffer_wire buffer_13093_1 (.in(n13093_0), .out(n13093_1));
wire n13094; //CHANY 1 (3,1) #56
wire n13094_0;
wire n13095; //CHANY 1 (3,1) #57
wire n13095_0;
wire n13096; //CHANY 2 (3,1) #58
wire n13096_0;
wire n13097; //CHANY 2 (3,1) #59
wire n13097_0;
wire n13098; //CHANY 3 (3,1) #60
wire n13098_0;
wire n13099; //CHANY 3 (3,1) #61
wire n13099_0;
wire n13100; //CHANY 4 (3,1) #62
wire n13100_0;
wire n13100_1;
buffer_wire buffer_13100_1 (.in(n13100_0), .out(n13100_1));
wire n13101; //CHANY 4 (3,1) #63
wire n13101_0;
wire n13101_1;
buffer_wire buffer_13101_1 (.in(n13101_0), .out(n13101_1));
wire n13102; //CHANY 1 (3,1) #64
wire n13102_0;
wire n13103; //CHANY 1 (3,1) #65
wire n13103_0;
wire n13104; //CHANY 2 (3,1) #66
wire n13104_0;
wire n13105; //CHANY 2 (3,1) #67
wire n13105_0;
wire n13106; //CHANY 3 (3,1) #68
wire n13106_0;
wire n13107; //CHANY 3 (3,1) #69
wire n13107_0;
wire n13108; //CHANY 4 (3,1) #70
wire n13108_0;
wire n13108_1;
buffer_wire buffer_13108_1 (.in(n13108_0), .out(n13108_1));
wire n13109; //CHANY 4 (3,1) #71
wire n13109_0;
wire n13109_1;
buffer_wire buffer_13109_1 (.in(n13109_0), .out(n13109_1));
wire n13110; //CHANY 1 (3,1) #72
wire n13110_0;
wire n13111; //CHANY 1 (3,1) #73
wire n13111_0;
wire n13112; //CHANY 2 (3,1) #74
wire n13112_0;
wire n13113; //CHANY 2 (3,1) #75
wire n13113_0;
wire n13114; //CHANY 3 (3,1) #76
wire n13114_0;
wire n13115; //CHANY 3 (3,1) #77
wire n13115_0;
wire n13116; //CHANY 4 (3,1) #78
wire n13116_0;
wire n13116_1;
buffer_wire buffer_13116_1 (.in(n13116_0), .out(n13116_1));
wire n13117; //CHANY 4 (3,1) #79
wire n13117_0;
wire n13117_1;
buffer_wire buffer_13117_1 (.in(n13117_0), .out(n13117_1));
wire n13118; //CHANY 5 (3,1) #80
wire n13118_0;
wire n13118_1;
buffer_wire buffer_13118_1 (.in(n13118_0), .out(n13118_1));
wire n13119; //CHANY 5 (3,1) #81
wire n13119_0;
wire n13119_1;
buffer_wire buffer_13119_1 (.in(n13119_0), .out(n13119_1));
wire n13120; //CHANY 6 (3,1) #82
wire n13120_0;
wire n13120_1;
buffer_wire buffer_13120_1 (.in(n13120_0), .out(n13120_1));
wire n13121; //CHANY 6 (3,1) #83
wire n13121_0;
wire n13121_1;
buffer_wire buffer_13121_1 (.in(n13121_0), .out(n13121_1));
wire n13122; //CHANY 7 (3,1) #84
wire n13122_0;
wire n13122_1;
wire n13122_2;
buffer_wire buffer_13122_2 (.in(n13122_1), .out(n13122_2));
buffer_wire buffer_13122_1 (.in(n13122_0), .out(n13122_1));
wire n13123; //CHANY 7 (3,1) #85
wire n13123_0;
wire n13123_1;
wire n13123_2;
buffer_wire buffer_13123_2 (.in(n13123_1), .out(n13123_2));
buffer_wire buffer_13123_1 (.in(n13123_0), .out(n13123_1));
wire n13124; //CHANY 8 (3,1) #86
wire n13124_0;
wire n13124_1;
wire n13124_2;
buffer_wire buffer_13124_2 (.in(n13124_1), .out(n13124_2));
buffer_wire buffer_13124_1 (.in(n13124_0), .out(n13124_1));
wire n13125; //CHANY 8 (3,1) #87
wire n13125_0;
wire n13125_1;
wire n13125_2;
buffer_wire buffer_13125_2 (.in(n13125_1), .out(n13125_2));
buffer_wire buffer_13125_1 (.in(n13125_0), .out(n13125_1));
wire n13126; //CHANY 9 (3,1) #88
wire n13126_0;
wire n13126_1;
wire n13126_2;
buffer_wire buffer_13126_2 (.in(n13126_1), .out(n13126_2));
buffer_wire buffer_13126_1 (.in(n13126_0), .out(n13126_1));
wire n13127; //CHANY 9 (3,1) #89
wire n13127_0;
wire n13127_1;
wire n13127_2;
buffer_wire buffer_13127_2 (.in(n13127_1), .out(n13127_2));
buffer_wire buffer_13127_1 (.in(n13127_0), .out(n13127_1));
wire n13128; //CHANY 9 (3,1) #90
wire n13128_0;
wire n13128_1;
wire n13128_2;
buffer_wire buffer_13128_2 (.in(n13128_1), .out(n13128_2));
buffer_wire buffer_13128_1 (.in(n13128_0), .out(n13128_1));
wire n13129; //CHANY 9 (3,1) #91
wire n13129_0;
wire n13129_1;
wire n13129_2;
buffer_wire buffer_13129_2 (.in(n13129_1), .out(n13129_2));
buffer_wire buffer_13129_1 (.in(n13129_0), .out(n13129_1));
wire n13130; //CHANY 4 (3,2) #0
wire n13130_0;
wire n13130_1;
buffer_wire buffer_13130_1 (.in(n13130_0), .out(n13130_1));
wire n13131; //CHANY 4 (3,2) #1
wire n13131_0;
wire n13131_1;
buffer_wire buffer_13131_1 (.in(n13131_0), .out(n13131_1));
wire n13132; //CHANY 4 (3,2) #8
wire n13132_0;
wire n13132_1;
buffer_wire buffer_13132_1 (.in(n13132_0), .out(n13132_1));
wire n13133; //CHANY 4 (3,2) #9
wire n13133_0;
wire n13133_1;
buffer_wire buffer_13133_1 (.in(n13133_0), .out(n13133_1));
wire n13134; //CHANY 4 (3,2) #16
wire n13134_0;
wire n13134_1;
buffer_wire buffer_13134_1 (.in(n13134_0), .out(n13134_1));
wire n13135; //CHANY 4 (3,2) #17
wire n13135_0;
wire n13135_1;
buffer_wire buffer_13135_1 (.in(n13135_0), .out(n13135_1));
wire n13136; //CHANY 4 (3,2) #24
wire n13136_0;
wire n13136_1;
buffer_wire buffer_13136_1 (.in(n13136_0), .out(n13136_1));
wire n13137; //CHANY 4 (3,2) #25
wire n13137_0;
wire n13137_1;
buffer_wire buffer_13137_1 (.in(n13137_0), .out(n13137_1));
wire n13138; //CHANY 4 (3,2) #32
wire n13138_0;
wire n13138_1;
buffer_wire buffer_13138_1 (.in(n13138_0), .out(n13138_1));
wire n13139; //CHANY 4 (3,2) #33
wire n13139_0;
wire n13139_1;
buffer_wire buffer_13139_1 (.in(n13139_0), .out(n13139_1));
wire n13140; //CHANY 4 (3,2) #40
wire n13140_0;
wire n13140_1;
buffer_wire buffer_13140_1 (.in(n13140_0), .out(n13140_1));
wire n13141; //CHANY 4 (3,2) #41
wire n13141_0;
wire n13141_1;
buffer_wire buffer_13141_1 (.in(n13141_0), .out(n13141_1));
wire n13142; //CHANY 4 (3,2) #48
wire n13142_0;
wire n13142_1;
buffer_wire buffer_13142_1 (.in(n13142_0), .out(n13142_1));
wire n13143; //CHANY 4 (3,2) #49
wire n13143_0;
wire n13143_1;
buffer_wire buffer_13143_1 (.in(n13143_0), .out(n13143_1));
wire n13144; //CHANY 4 (3,2) #56
wire n13144_0;
wire n13144_1;
buffer_wire buffer_13144_1 (.in(n13144_0), .out(n13144_1));
wire n13145; //CHANY 4 (3,2) #57
wire n13145_0;
wire n13145_1;
buffer_wire buffer_13145_1 (.in(n13145_0), .out(n13145_1));
wire n13146; //CHANY 4 (3,2) #64
wire n13146_0;
wire n13146_1;
buffer_wire buffer_13146_1 (.in(n13146_0), .out(n13146_1));
wire n13147; //CHANY 4 (3,2) #65
wire n13147_0;
wire n13147_1;
buffer_wire buffer_13147_1 (.in(n13147_0), .out(n13147_1));
wire n13148; //CHANY 4 (3,2) #72
wire n13148_0;
wire n13148_1;
buffer_wire buffer_13148_1 (.in(n13148_0), .out(n13148_1));
wire n13149; //CHANY 4 (3,2) #73
wire n13149_0;
wire n13149_1;
buffer_wire buffer_13149_1 (.in(n13149_0), .out(n13149_1));
wire n13150; //CHANY 4 (3,3) #2
wire n13150_0;
wire n13150_1;
buffer_wire buffer_13150_1 (.in(n13150_0), .out(n13150_1));
wire n13151; //CHANY 4 (3,3) #3
wire n13151_0;
wire n13151_1;
buffer_wire buffer_13151_1 (.in(n13151_0), .out(n13151_1));
wire n13152; //CHANY 4 (3,3) #10
wire n13152_0;
wire n13152_1;
buffer_wire buffer_13152_1 (.in(n13152_0), .out(n13152_1));
wire n13153; //CHANY 4 (3,3) #11
wire n13153_0;
wire n13153_1;
buffer_wire buffer_13153_1 (.in(n13153_0), .out(n13153_1));
wire n13154; //CHANY 4 (3,3) #18
wire n13154_0;
wire n13154_1;
buffer_wire buffer_13154_1 (.in(n13154_0), .out(n13154_1));
wire n13155; //CHANY 4 (3,3) #19
wire n13155_0;
wire n13155_1;
buffer_wire buffer_13155_1 (.in(n13155_0), .out(n13155_1));
wire n13156; //CHANY 4 (3,3) #26
wire n13156_0;
wire n13156_1;
buffer_wire buffer_13156_1 (.in(n13156_0), .out(n13156_1));
wire n13157; //CHANY 4 (3,3) #27
wire n13157_0;
wire n13157_1;
buffer_wire buffer_13157_1 (.in(n13157_0), .out(n13157_1));
wire n13158; //CHANY 4 (3,3) #34
wire n13158_0;
wire n13158_1;
buffer_wire buffer_13158_1 (.in(n13158_0), .out(n13158_1));
wire n13159; //CHANY 4 (3,3) #35
wire n13159_0;
wire n13159_1;
buffer_wire buffer_13159_1 (.in(n13159_0), .out(n13159_1));
wire n13160; //CHANY 4 (3,3) #42
wire n13160_0;
wire n13160_1;
buffer_wire buffer_13160_1 (.in(n13160_0), .out(n13160_1));
wire n13161; //CHANY 4 (3,3) #43
wire n13161_0;
wire n13161_1;
buffer_wire buffer_13161_1 (.in(n13161_0), .out(n13161_1));
wire n13162; //CHANY 4 (3,3) #50
wire n13162_0;
wire n13162_1;
buffer_wire buffer_13162_1 (.in(n13162_0), .out(n13162_1));
wire n13163; //CHANY 4 (3,3) #51
wire n13163_0;
wire n13163_1;
buffer_wire buffer_13163_1 (.in(n13163_0), .out(n13163_1));
wire n13164; //CHANY 4 (3,3) #58
wire n13164_0;
wire n13164_1;
buffer_wire buffer_13164_1 (.in(n13164_0), .out(n13164_1));
wire n13165; //CHANY 4 (3,3) #59
wire n13165_0;
wire n13165_1;
buffer_wire buffer_13165_1 (.in(n13165_0), .out(n13165_1));
wire n13166; //CHANY 4 (3,3) #66
wire n13166_0;
wire n13166_1;
buffer_wire buffer_13166_1 (.in(n13166_0), .out(n13166_1));
wire n13167; //CHANY 4 (3,3) #67
wire n13167_0;
wire n13167_1;
buffer_wire buffer_13167_1 (.in(n13167_0), .out(n13167_1));
wire n13168; //CHANY 4 (3,3) #74
wire n13168_0;
wire n13168_1;
buffer_wire buffer_13168_1 (.in(n13168_0), .out(n13168_1));
wire n13169; //CHANY 4 (3,3) #75
wire n13169_0;
wire n13169_1;
buffer_wire buffer_13169_1 (.in(n13169_0), .out(n13169_1));
wire n13170; //CHANY 4 (3,4) #4
wire n13170_0;
wire n13170_1;
buffer_wire buffer_13170_1 (.in(n13170_0), .out(n13170_1));
wire n13171; //CHANY 4 (3,4) #5
wire n13171_0;
wire n13171_1;
buffer_wire buffer_13171_1 (.in(n13171_0), .out(n13171_1));
wire n13172; //CHANY 4 (3,4) #12
wire n13172_0;
wire n13172_1;
buffer_wire buffer_13172_1 (.in(n13172_0), .out(n13172_1));
wire n13173; //CHANY 4 (3,4) #13
wire n13173_0;
wire n13173_1;
buffer_wire buffer_13173_1 (.in(n13173_0), .out(n13173_1));
wire n13174; //CHANY 4 (3,4) #20
wire n13174_0;
wire n13174_1;
buffer_wire buffer_13174_1 (.in(n13174_0), .out(n13174_1));
wire n13175; //CHANY 4 (3,4) #21
wire n13175_0;
wire n13175_1;
buffer_wire buffer_13175_1 (.in(n13175_0), .out(n13175_1));
wire n13176; //CHANY 4 (3,4) #28
wire n13176_0;
wire n13176_1;
buffer_wire buffer_13176_1 (.in(n13176_0), .out(n13176_1));
wire n13177; //CHANY 4 (3,4) #29
wire n13177_0;
wire n13177_1;
buffer_wire buffer_13177_1 (.in(n13177_0), .out(n13177_1));
wire n13178; //CHANY 4 (3,4) #36
wire n13178_0;
wire n13178_1;
buffer_wire buffer_13178_1 (.in(n13178_0), .out(n13178_1));
wire n13179; //CHANY 4 (3,4) #37
wire n13179_0;
wire n13179_1;
buffer_wire buffer_13179_1 (.in(n13179_0), .out(n13179_1));
wire n13180; //CHANY 4 (3,4) #44
wire n13180_0;
wire n13180_1;
buffer_wire buffer_13180_1 (.in(n13180_0), .out(n13180_1));
wire n13181; //CHANY 4 (3,4) #45
wire n13181_0;
wire n13181_1;
buffer_wire buffer_13181_1 (.in(n13181_0), .out(n13181_1));
wire n13182; //CHANY 4 (3,4) #52
wire n13182_0;
wire n13182_1;
buffer_wire buffer_13182_1 (.in(n13182_0), .out(n13182_1));
wire n13183; //CHANY 4 (3,4) #53
wire n13183_0;
wire n13183_1;
buffer_wire buffer_13183_1 (.in(n13183_0), .out(n13183_1));
wire n13184; //CHANY 4 (3,4) #60
wire n13184_0;
wire n13184_1;
buffer_wire buffer_13184_1 (.in(n13184_0), .out(n13184_1));
wire n13185; //CHANY 4 (3,4) #61
wire n13185_0;
wire n13185_1;
buffer_wire buffer_13185_1 (.in(n13185_0), .out(n13185_1));
wire n13186; //CHANY 4 (3,4) #68
wire n13186_0;
wire n13186_1;
buffer_wire buffer_13186_1 (.in(n13186_0), .out(n13186_1));
wire n13187; //CHANY 4 (3,4) #69
wire n13187_0;
wire n13187_1;
buffer_wire buffer_13187_1 (.in(n13187_0), .out(n13187_1));
wire n13188; //CHANY 4 (3,4) #76
wire n13188_0;
wire n13188_1;
buffer_wire buffer_13188_1 (.in(n13188_0), .out(n13188_1));
wire n13189; //CHANY 4 (3,4) #77
wire n13189_0;
wire n13189_1;
buffer_wire buffer_13189_1 (.in(n13189_0), .out(n13189_1));
wire n13190; //CHANY 4 (3,5) #6
wire n13190_0;
wire n13190_1;
buffer_wire buffer_13190_1 (.in(n13190_0), .out(n13190_1));
wire n13191; //CHANY 4 (3,5) #7
wire n13191_0;
wire n13191_1;
buffer_wire buffer_13191_1 (.in(n13191_0), .out(n13191_1));
wire n13192; //CHANY 4 (3,5) #14
wire n13192_0;
wire n13192_1;
buffer_wire buffer_13192_1 (.in(n13192_0), .out(n13192_1));
wire n13193; //CHANY 4 (3,5) #15
wire n13193_0;
wire n13193_1;
buffer_wire buffer_13193_1 (.in(n13193_0), .out(n13193_1));
wire n13194; //CHANY 4 (3,5) #22
wire n13194_0;
wire n13194_1;
buffer_wire buffer_13194_1 (.in(n13194_0), .out(n13194_1));
wire n13195; //CHANY 4 (3,5) #23
wire n13195_0;
wire n13195_1;
buffer_wire buffer_13195_1 (.in(n13195_0), .out(n13195_1));
wire n13196; //CHANY 4 (3,5) #30
wire n13196_0;
wire n13196_1;
buffer_wire buffer_13196_1 (.in(n13196_0), .out(n13196_1));
wire n13197; //CHANY 4 (3,5) #31
wire n13197_0;
wire n13197_1;
buffer_wire buffer_13197_1 (.in(n13197_0), .out(n13197_1));
wire n13198; //CHANY 4 (3,5) #38
wire n13198_0;
wire n13198_1;
buffer_wire buffer_13198_1 (.in(n13198_0), .out(n13198_1));
wire n13199; //CHANY 4 (3,5) #39
wire n13199_0;
wire n13199_1;
buffer_wire buffer_13199_1 (.in(n13199_0), .out(n13199_1));
wire n13200; //CHANY 4 (3,5) #46
wire n13200_0;
wire n13200_1;
buffer_wire buffer_13200_1 (.in(n13200_0), .out(n13200_1));
wire n13201; //CHANY 4 (3,5) #47
wire n13201_0;
wire n13201_1;
buffer_wire buffer_13201_1 (.in(n13201_0), .out(n13201_1));
wire n13202; //CHANY 4 (3,5) #54
wire n13202_0;
wire n13202_1;
buffer_wire buffer_13202_1 (.in(n13202_0), .out(n13202_1));
wire n13203; //CHANY 4 (3,5) #55
wire n13203_0;
wire n13203_1;
buffer_wire buffer_13203_1 (.in(n13203_0), .out(n13203_1));
wire n13204; //CHANY 4 (3,5) #62
wire n13204_0;
wire n13204_1;
buffer_wire buffer_13204_1 (.in(n13204_0), .out(n13204_1));
wire n13205; //CHANY 4 (3,5) #63
wire n13205_0;
wire n13205_1;
buffer_wire buffer_13205_1 (.in(n13205_0), .out(n13205_1));
wire n13206; //CHANY 4 (3,5) #70
wire n13206_0;
wire n13206_1;
buffer_wire buffer_13206_1 (.in(n13206_0), .out(n13206_1));
wire n13207; //CHANY 4 (3,5) #71
wire n13207_0;
wire n13207_1;
buffer_wire buffer_13207_1 (.in(n13207_0), .out(n13207_1));
wire n13208; //CHANY 4 (3,5) #78
wire n13208_0;
wire n13208_1;
buffer_wire buffer_13208_1 (.in(n13208_0), .out(n13208_1));
wire n13209; //CHANY 4 (3,5) #79
wire n13209_0;
wire n13209_1;
buffer_wire buffer_13209_1 (.in(n13209_0), .out(n13209_1));
wire n13210; //CHANY 4 (3,6) #0
wire n13210_0;
wire n13210_1;
buffer_wire buffer_13210_1 (.in(n13210_0), .out(n13210_1));
wire n13211; //CHANY 4 (3,6) #1
wire n13211_0;
wire n13211_1;
buffer_wire buffer_13211_1 (.in(n13211_0), .out(n13211_1));
wire n13212; //CHANY 4 (3,6) #8
wire n13212_0;
wire n13212_1;
buffer_wire buffer_13212_1 (.in(n13212_0), .out(n13212_1));
wire n13213; //CHANY 4 (3,6) #9
wire n13213_0;
wire n13213_1;
buffer_wire buffer_13213_1 (.in(n13213_0), .out(n13213_1));
wire n13214; //CHANY 4 (3,6) #16
wire n13214_0;
wire n13214_1;
buffer_wire buffer_13214_1 (.in(n13214_0), .out(n13214_1));
wire n13215; //CHANY 4 (3,6) #17
wire n13215_0;
wire n13215_1;
buffer_wire buffer_13215_1 (.in(n13215_0), .out(n13215_1));
wire n13216; //CHANY 4 (3,6) #24
wire n13216_0;
wire n13216_1;
buffer_wire buffer_13216_1 (.in(n13216_0), .out(n13216_1));
wire n13217; //CHANY 4 (3,6) #25
wire n13217_0;
wire n13217_1;
buffer_wire buffer_13217_1 (.in(n13217_0), .out(n13217_1));
wire n13218; //CHANY 4 (3,6) #32
wire n13218_0;
wire n13218_1;
buffer_wire buffer_13218_1 (.in(n13218_0), .out(n13218_1));
wire n13219; //CHANY 4 (3,6) #33
wire n13219_0;
wire n13219_1;
buffer_wire buffer_13219_1 (.in(n13219_0), .out(n13219_1));
wire n13220; //CHANY 4 (3,6) #40
wire n13220_0;
wire n13220_1;
buffer_wire buffer_13220_1 (.in(n13220_0), .out(n13220_1));
wire n13221; //CHANY 4 (3,6) #41
wire n13221_0;
wire n13221_1;
buffer_wire buffer_13221_1 (.in(n13221_0), .out(n13221_1));
wire n13222; //CHANY 4 (3,6) #48
wire n13222_0;
wire n13222_1;
buffer_wire buffer_13222_1 (.in(n13222_0), .out(n13222_1));
wire n13223; //CHANY 4 (3,6) #49
wire n13223_0;
wire n13223_1;
buffer_wire buffer_13223_1 (.in(n13223_0), .out(n13223_1));
wire n13224; //CHANY 4 (3,6) #56
wire n13224_0;
wire n13224_1;
buffer_wire buffer_13224_1 (.in(n13224_0), .out(n13224_1));
wire n13225; //CHANY 4 (3,6) #57
wire n13225_0;
wire n13225_1;
buffer_wire buffer_13225_1 (.in(n13225_0), .out(n13225_1));
wire n13226; //CHANY 4 (3,6) #64
wire n13226_0;
wire n13226_1;
buffer_wire buffer_13226_1 (.in(n13226_0), .out(n13226_1));
wire n13227; //CHANY 4 (3,6) #65
wire n13227_0;
wire n13227_1;
buffer_wire buffer_13227_1 (.in(n13227_0), .out(n13227_1));
wire n13228; //CHANY 4 (3,6) #72
wire n13228_0;
wire n13228_1;
buffer_wire buffer_13228_1 (.in(n13228_0), .out(n13228_1));
wire n13229; //CHANY 4 (3,6) #73
wire n13229_0;
wire n13229_1;
buffer_wire buffer_13229_1 (.in(n13229_0), .out(n13229_1));
wire n13230; //CHANY 4 (3,6) #80
wire n13230_0;
wire n13230_1;
buffer_wire buffer_13230_1 (.in(n13230_0), .out(n13230_1));
wire n13231; //CHANY 4 (3,6) #81
wire n13231_0;
wire n13231_1;
buffer_wire buffer_13231_1 (.in(n13231_0), .out(n13231_1));
wire n13232; //CHANY 3 (3,7) #2
wire n13232_0;
wire n13233; //CHANY 3 (3,7) #3
wire n13233_0;
wire n13234; //CHANY 3 (3,7) #10
wire n13234_0;
wire n13235; //CHANY 3 (3,7) #11
wire n13235_0;
wire n13236; //CHANY 3 (3,7) #18
wire n13236_0;
wire n13237; //CHANY 3 (3,7) #19
wire n13237_0;
wire n13238; //CHANY 3 (3,7) #26
wire n13238_0;
wire n13239; //CHANY 3 (3,7) #27
wire n13239_0;
wire n13240; //CHANY 3 (3,7) #34
wire n13240_0;
wire n13241; //CHANY 3 (3,7) #35
wire n13241_0;
wire n13242; //CHANY 3 (3,7) #42
wire n13242_0;
wire n13243; //CHANY 3 (3,7) #43
wire n13243_0;
wire n13244; //CHANY 3 (3,7) #50
wire n13244_0;
wire n13245; //CHANY 3 (3,7) #51
wire n13245_0;
wire n13246; //CHANY 3 (3,7) #58
wire n13246_0;
wire n13247; //CHANY 3 (3,7) #59
wire n13247_0;
wire n13248; //CHANY 3 (3,7) #66
wire n13248_0;
wire n13249; //CHANY 3 (3,7) #67
wire n13249_0;
wire n13250; //CHANY 3 (3,7) #74
wire n13250_0;
wire n13251; //CHANY 3 (3,7) #75
wire n13251_0;
wire n13252; //CHANY 3 (3,7) #82
wire n13252_0;
wire n13253; //CHANY 3 (3,7) #83
wire n13253_0;
wire n13254; //CHANY 2 (3,8) #4
wire n13254_0;
wire n13255; //CHANY 2 (3,8) #5
wire n13255_0;
wire n13256; //CHANY 2 (3,8) #12
wire n13256_0;
wire n13257; //CHANY 2 (3,8) #13
wire n13257_0;
wire n13258; //CHANY 2 (3,8) #20
wire n13258_0;
wire n13259; //CHANY 2 (3,8) #21
wire n13259_0;
wire n13260; //CHANY 2 (3,8) #28
wire n13260_0;
wire n13261; //CHANY 2 (3,8) #29
wire n13261_0;
wire n13262; //CHANY 2 (3,8) #36
wire n13262_0;
wire n13263; //CHANY 2 (3,8) #37
wire n13263_0;
wire n13264; //CHANY 2 (3,8) #44
wire n13264_0;
wire n13265; //CHANY 2 (3,8) #45
wire n13265_0;
wire n13266; //CHANY 2 (3,8) #52
wire n13266_0;
wire n13267; //CHANY 2 (3,8) #53
wire n13267_0;
wire n13268; //CHANY 2 (3,8) #60
wire n13268_0;
wire n13269; //CHANY 2 (3,8) #61
wire n13269_0;
wire n13270; //CHANY 2 (3,8) #68
wire n13270_0;
wire n13271; //CHANY 2 (3,8) #69
wire n13271_0;
wire n13272; //CHANY 2 (3,8) #76
wire n13272_0;
wire n13273; //CHANY 2 (3,8) #77
wire n13273_0;
wire n13274; //CHANY 2 (3,8) #84
wire n13274_0;
wire n13275; //CHANY 2 (3,8) #85
wire n13275_0;
wire n13276; //CHANY 1 (3,9) #6
wire n13276_0;
wire n13277; //CHANY 1 (3,9) #7
wire n13277_0;
wire n13278; //CHANY 1 (3,9) #14
wire n13278_0;
wire n13279; //CHANY 1 (3,9) #15
wire n13279_0;
wire n13280; //CHANY 1 (3,9) #22
wire n13280_0;
wire n13281; //CHANY 1 (3,9) #23
wire n13281_0;
wire n13282; //CHANY 1 (3,9) #30
wire n13282_0;
wire n13283; //CHANY 1 (3,9) #31
wire n13283_0;
wire n13284; //CHANY 1 (3,9) #38
wire n13284_0;
wire n13285; //CHANY 1 (3,9) #39
wire n13285_0;
wire n13286; //CHANY 1 (3,9) #46
wire n13286_0;
wire n13287; //CHANY 1 (3,9) #47
wire n13287_0;
wire n13288; //CHANY 1 (3,9) #54
wire n13288_0;
wire n13289; //CHANY 1 (3,9) #55
wire n13289_0;
wire n13290; //CHANY 1 (3,9) #62
wire n13290_0;
wire n13291; //CHANY 1 (3,9) #63
wire n13291_0;
wire n13292; //CHANY 1 (3,9) #70
wire n13292_0;
wire n13293; //CHANY 1 (3,9) #71
wire n13293_0;
wire n13294; //CHANY 1 (3,9) #78
wire n13294_0;
wire n13295; //CHANY 1 (3,9) #79
wire n13295_0;
wire n13296; //CHANY 1 (3,9) #86
wire n13296_0;
wire n13297; //CHANY 1 (3,9) #87
wire n13297_0;
wire n13298; //CHANY 4 (4,1) #0
wire n13298_0;
wire n13298_1;
buffer_wire buffer_13298_1 (.in(n13298_0), .out(n13298_1));
wire n13299; //CHANY 4 (4,1) #1
wire n13299_0;
wire n13299_1;
buffer_wire buffer_13299_1 (.in(n13299_0), .out(n13299_1));
wire n13300; //CHANY 1 (4,1) #2
wire n13300_0;
wire n13301; //CHANY 1 (4,1) #3
wire n13301_0;
wire n13302; //CHANY 2 (4,1) #4
wire n13302_0;
wire n13303; //CHANY 2 (4,1) #5
wire n13303_0;
wire n13304; //CHANY 3 (4,1) #6
wire n13304_0;
wire n13305; //CHANY 3 (4,1) #7
wire n13305_0;
wire n13306; //CHANY 4 (4,1) #8
wire n13306_0;
wire n13306_1;
buffer_wire buffer_13306_1 (.in(n13306_0), .out(n13306_1));
wire n13307; //CHANY 4 (4,1) #9
wire n13307_0;
wire n13307_1;
buffer_wire buffer_13307_1 (.in(n13307_0), .out(n13307_1));
wire n13308; //CHANY 1 (4,1) #10
wire n13308_0;
wire n13309; //CHANY 1 (4,1) #11
wire n13309_0;
wire n13310; //CHANY 2 (4,1) #12
wire n13310_0;
wire n13311; //CHANY 2 (4,1) #13
wire n13311_0;
wire n13312; //CHANY 3 (4,1) #14
wire n13312_0;
wire n13313; //CHANY 3 (4,1) #15
wire n13313_0;
wire n13314; //CHANY 4 (4,1) #16
wire n13314_0;
wire n13314_1;
buffer_wire buffer_13314_1 (.in(n13314_0), .out(n13314_1));
wire n13315; //CHANY 4 (4,1) #17
wire n13315_0;
wire n13315_1;
buffer_wire buffer_13315_1 (.in(n13315_0), .out(n13315_1));
wire n13316; //CHANY 1 (4,1) #18
wire n13316_0;
wire n13317; //CHANY 1 (4,1) #19
wire n13317_0;
wire n13318; //CHANY 2 (4,1) #20
wire n13318_0;
wire n13319; //CHANY 2 (4,1) #21
wire n13319_0;
wire n13320; //CHANY 3 (4,1) #22
wire n13320_0;
wire n13321; //CHANY 3 (4,1) #23
wire n13321_0;
wire n13322; //CHANY 4 (4,1) #24
wire n13322_0;
wire n13322_1;
buffer_wire buffer_13322_1 (.in(n13322_0), .out(n13322_1));
wire n13323; //CHANY 4 (4,1) #25
wire n13323_0;
wire n13323_1;
buffer_wire buffer_13323_1 (.in(n13323_0), .out(n13323_1));
wire n13324; //CHANY 1 (4,1) #26
wire n13324_0;
wire n13325; //CHANY 1 (4,1) #27
wire n13325_0;
wire n13326; //CHANY 2 (4,1) #28
wire n13326_0;
wire n13327; //CHANY 2 (4,1) #29
wire n13327_0;
wire n13328; //CHANY 3 (4,1) #30
wire n13328_0;
wire n13329; //CHANY 3 (4,1) #31
wire n13329_0;
wire n13330; //CHANY 4 (4,1) #32
wire n13330_0;
wire n13330_1;
buffer_wire buffer_13330_1 (.in(n13330_0), .out(n13330_1));
wire n13331; //CHANY 4 (4,1) #33
wire n13331_0;
wire n13331_1;
buffer_wire buffer_13331_1 (.in(n13331_0), .out(n13331_1));
wire n13332; //CHANY 1 (4,1) #34
wire n13332_0;
wire n13333; //CHANY 1 (4,1) #35
wire n13333_0;
wire n13334; //CHANY 2 (4,1) #36
wire n13334_0;
wire n13335; //CHANY 2 (4,1) #37
wire n13335_0;
wire n13336; //CHANY 3 (4,1) #38
wire n13336_0;
wire n13337; //CHANY 3 (4,1) #39
wire n13337_0;
wire n13338; //CHANY 4 (4,1) #40
wire n13338_0;
wire n13338_1;
buffer_wire buffer_13338_1 (.in(n13338_0), .out(n13338_1));
wire n13339; //CHANY 4 (4,1) #41
wire n13339_0;
wire n13339_1;
buffer_wire buffer_13339_1 (.in(n13339_0), .out(n13339_1));
wire n13340; //CHANY 1 (4,1) #42
wire n13340_0;
wire n13341; //CHANY 1 (4,1) #43
wire n13341_0;
wire n13342; //CHANY 2 (4,1) #44
wire n13342_0;
wire n13343; //CHANY 2 (4,1) #45
wire n13343_0;
wire n13344; //CHANY 3 (4,1) #46
wire n13344_0;
wire n13345; //CHANY 3 (4,1) #47
wire n13345_0;
wire n13346; //CHANY 4 (4,1) #48
wire n13346_0;
wire n13346_1;
buffer_wire buffer_13346_1 (.in(n13346_0), .out(n13346_1));
wire n13347; //CHANY 4 (4,1) #49
wire n13347_0;
wire n13347_1;
buffer_wire buffer_13347_1 (.in(n13347_0), .out(n13347_1));
wire n13348; //CHANY 1 (4,1) #50
wire n13348_0;
wire n13349; //CHANY 1 (4,1) #51
wire n13349_0;
wire n13350; //CHANY 2 (4,1) #52
wire n13350_0;
wire n13351; //CHANY 2 (4,1) #53
wire n13351_0;
wire n13352; //CHANY 3 (4,1) #54
wire n13352_0;
wire n13353; //CHANY 3 (4,1) #55
wire n13353_0;
wire n13354; //CHANY 4 (4,1) #56
wire n13354_0;
wire n13354_1;
buffer_wire buffer_13354_1 (.in(n13354_0), .out(n13354_1));
wire n13355; //CHANY 4 (4,1) #57
wire n13355_0;
wire n13355_1;
buffer_wire buffer_13355_1 (.in(n13355_0), .out(n13355_1));
wire n13356; //CHANY 1 (4,1) #58
wire n13356_0;
wire n13357; //CHANY 1 (4,1) #59
wire n13357_0;
wire n13358; //CHANY 2 (4,1) #60
wire n13358_0;
wire n13359; //CHANY 2 (4,1) #61
wire n13359_0;
wire n13360; //CHANY 3 (4,1) #62
wire n13360_0;
wire n13361; //CHANY 3 (4,1) #63
wire n13361_0;
wire n13362; //CHANY 4 (4,1) #64
wire n13362_0;
wire n13362_1;
buffer_wire buffer_13362_1 (.in(n13362_0), .out(n13362_1));
wire n13363; //CHANY 4 (4,1) #65
wire n13363_0;
wire n13363_1;
buffer_wire buffer_13363_1 (.in(n13363_0), .out(n13363_1));
wire n13364; //CHANY 1 (4,1) #66
wire n13364_0;
wire n13365; //CHANY 1 (4,1) #67
wire n13365_0;
wire n13366; //CHANY 2 (4,1) #68
wire n13366_0;
wire n13367; //CHANY 2 (4,1) #69
wire n13367_0;
wire n13368; //CHANY 3 (4,1) #70
wire n13368_0;
wire n13369; //CHANY 3 (4,1) #71
wire n13369_0;
wire n13370; //CHANY 4 (4,1) #72
wire n13370_0;
wire n13370_1;
buffer_wire buffer_13370_1 (.in(n13370_0), .out(n13370_1));
wire n13371; //CHANY 4 (4,1) #73
wire n13371_0;
wire n13371_1;
buffer_wire buffer_13371_1 (.in(n13371_0), .out(n13371_1));
wire n13372; //CHANY 1 (4,1) #74
wire n13372_0;
wire n13373; //CHANY 1 (4,1) #75
wire n13373_0;
wire n13374; //CHANY 2 (4,1) #76
wire n13374_0;
wire n13375; //CHANY 2 (4,1) #77
wire n13375_0;
wire n13376; //CHANY 3 (4,1) #78
wire n13376_0;
wire n13377; //CHANY 3 (4,1) #79
wire n13377_0;
wire n13378; //CHANY 4 (4,1) #80
wire n13378_0;
wire n13378_1;
buffer_wire buffer_13378_1 (.in(n13378_0), .out(n13378_1));
wire n13379; //CHANY 4 (4,1) #81
wire n13379_0;
wire n13379_1;
buffer_wire buffer_13379_1 (.in(n13379_0), .out(n13379_1));
wire n13380; //CHANY 5 (4,1) #82
wire n13380_0;
wire n13380_1;
buffer_wire buffer_13380_1 (.in(n13380_0), .out(n13380_1));
wire n13381; //CHANY 5 (4,1) #83
wire n13381_0;
wire n13381_1;
buffer_wire buffer_13381_1 (.in(n13381_0), .out(n13381_1));
wire n13382; //CHANY 6 (4,1) #84
wire n13382_0;
wire n13382_1;
buffer_wire buffer_13382_1 (.in(n13382_0), .out(n13382_1));
wire n13383; //CHANY 6 (4,1) #85
wire n13383_0;
wire n13383_1;
buffer_wire buffer_13383_1 (.in(n13383_0), .out(n13383_1));
wire n13384; //CHANY 7 (4,1) #86
wire n13384_0;
wire n13384_1;
wire n13384_2;
buffer_wire buffer_13384_2 (.in(n13384_1), .out(n13384_2));
buffer_wire buffer_13384_1 (.in(n13384_0), .out(n13384_1));
wire n13385; //CHANY 7 (4,1) #87
wire n13385_0;
wire n13385_1;
wire n13385_2;
buffer_wire buffer_13385_2 (.in(n13385_1), .out(n13385_2));
buffer_wire buffer_13385_1 (.in(n13385_0), .out(n13385_1));
wire n13386; //CHANY 8 (4,1) #88
wire n13386_0;
wire n13386_1;
wire n13386_2;
buffer_wire buffer_13386_2 (.in(n13386_1), .out(n13386_2));
buffer_wire buffer_13386_1 (.in(n13386_0), .out(n13386_1));
wire n13387; //CHANY 8 (4,1) #89
wire n13387_0;
wire n13387_1;
wire n13387_2;
buffer_wire buffer_13387_2 (.in(n13387_1), .out(n13387_2));
buffer_wire buffer_13387_1 (.in(n13387_0), .out(n13387_1));
wire n13388; //CHANY 9 (4,1) #90
wire n13388_0;
wire n13388_1;
wire n13388_2;
buffer_wire buffer_13388_2 (.in(n13388_1), .out(n13388_2));
buffer_wire buffer_13388_1 (.in(n13388_0), .out(n13388_1));
wire n13389; //CHANY 9 (4,1) #91
wire n13389_0;
wire n13389_1;
wire n13389_2;
buffer_wire buffer_13389_2 (.in(n13389_1), .out(n13389_2));
buffer_wire buffer_13389_1 (.in(n13389_0), .out(n13389_1));
wire n13390; //CHANY 4 (4,2) #2
wire n13390_0;
wire n13390_1;
buffer_wire buffer_13390_1 (.in(n13390_0), .out(n13390_1));
wire n13391; //CHANY 4 (4,2) #3
wire n13391_0;
wire n13391_1;
buffer_wire buffer_13391_1 (.in(n13391_0), .out(n13391_1));
wire n13392; //CHANY 4 (4,2) #10
wire n13392_0;
wire n13392_1;
buffer_wire buffer_13392_1 (.in(n13392_0), .out(n13392_1));
wire n13393; //CHANY 4 (4,2) #11
wire n13393_0;
wire n13393_1;
buffer_wire buffer_13393_1 (.in(n13393_0), .out(n13393_1));
wire n13394; //CHANY 4 (4,2) #18
wire n13394_0;
wire n13394_1;
buffer_wire buffer_13394_1 (.in(n13394_0), .out(n13394_1));
wire n13395; //CHANY 4 (4,2) #19
wire n13395_0;
wire n13395_1;
buffer_wire buffer_13395_1 (.in(n13395_0), .out(n13395_1));
wire n13396; //CHANY 4 (4,2) #26
wire n13396_0;
wire n13396_1;
buffer_wire buffer_13396_1 (.in(n13396_0), .out(n13396_1));
wire n13397; //CHANY 4 (4,2) #27
wire n13397_0;
wire n13397_1;
buffer_wire buffer_13397_1 (.in(n13397_0), .out(n13397_1));
wire n13398; //CHANY 4 (4,2) #34
wire n13398_0;
wire n13398_1;
buffer_wire buffer_13398_1 (.in(n13398_0), .out(n13398_1));
wire n13399; //CHANY 4 (4,2) #35
wire n13399_0;
wire n13399_1;
buffer_wire buffer_13399_1 (.in(n13399_0), .out(n13399_1));
wire n13400; //CHANY 4 (4,2) #42
wire n13400_0;
wire n13400_1;
buffer_wire buffer_13400_1 (.in(n13400_0), .out(n13400_1));
wire n13401; //CHANY 4 (4,2) #43
wire n13401_0;
wire n13401_1;
buffer_wire buffer_13401_1 (.in(n13401_0), .out(n13401_1));
wire n13402; //CHANY 4 (4,2) #50
wire n13402_0;
wire n13402_1;
buffer_wire buffer_13402_1 (.in(n13402_0), .out(n13402_1));
wire n13403; //CHANY 4 (4,2) #51
wire n13403_0;
wire n13403_1;
buffer_wire buffer_13403_1 (.in(n13403_0), .out(n13403_1));
wire n13404; //CHANY 4 (4,2) #58
wire n13404_0;
wire n13404_1;
buffer_wire buffer_13404_1 (.in(n13404_0), .out(n13404_1));
wire n13405; //CHANY 4 (4,2) #59
wire n13405_0;
wire n13405_1;
buffer_wire buffer_13405_1 (.in(n13405_0), .out(n13405_1));
wire n13406; //CHANY 4 (4,2) #66
wire n13406_0;
wire n13406_1;
buffer_wire buffer_13406_1 (.in(n13406_0), .out(n13406_1));
wire n13407; //CHANY 4 (4,2) #67
wire n13407_0;
wire n13407_1;
buffer_wire buffer_13407_1 (.in(n13407_0), .out(n13407_1));
wire n13408; //CHANY 4 (4,2) #74
wire n13408_0;
wire n13408_1;
buffer_wire buffer_13408_1 (.in(n13408_0), .out(n13408_1));
wire n13409; //CHANY 4 (4,2) #75
wire n13409_0;
wire n13409_1;
buffer_wire buffer_13409_1 (.in(n13409_0), .out(n13409_1));
wire n13410; //CHANY 4 (4,3) #4
wire n13410_0;
wire n13410_1;
buffer_wire buffer_13410_1 (.in(n13410_0), .out(n13410_1));
wire n13411; //CHANY 4 (4,3) #5
wire n13411_0;
wire n13411_1;
buffer_wire buffer_13411_1 (.in(n13411_0), .out(n13411_1));
wire n13412; //CHANY 4 (4,3) #12
wire n13412_0;
wire n13412_1;
buffer_wire buffer_13412_1 (.in(n13412_0), .out(n13412_1));
wire n13413; //CHANY 4 (4,3) #13
wire n13413_0;
wire n13413_1;
buffer_wire buffer_13413_1 (.in(n13413_0), .out(n13413_1));
wire n13414; //CHANY 4 (4,3) #20
wire n13414_0;
wire n13414_1;
buffer_wire buffer_13414_1 (.in(n13414_0), .out(n13414_1));
wire n13415; //CHANY 4 (4,3) #21
wire n13415_0;
wire n13415_1;
buffer_wire buffer_13415_1 (.in(n13415_0), .out(n13415_1));
wire n13416; //CHANY 4 (4,3) #28
wire n13416_0;
wire n13416_1;
buffer_wire buffer_13416_1 (.in(n13416_0), .out(n13416_1));
wire n13417; //CHANY 4 (4,3) #29
wire n13417_0;
wire n13417_1;
buffer_wire buffer_13417_1 (.in(n13417_0), .out(n13417_1));
wire n13418; //CHANY 4 (4,3) #36
wire n13418_0;
wire n13418_1;
buffer_wire buffer_13418_1 (.in(n13418_0), .out(n13418_1));
wire n13419; //CHANY 4 (4,3) #37
wire n13419_0;
wire n13419_1;
buffer_wire buffer_13419_1 (.in(n13419_0), .out(n13419_1));
wire n13420; //CHANY 4 (4,3) #44
wire n13420_0;
wire n13420_1;
buffer_wire buffer_13420_1 (.in(n13420_0), .out(n13420_1));
wire n13421; //CHANY 4 (4,3) #45
wire n13421_0;
wire n13421_1;
buffer_wire buffer_13421_1 (.in(n13421_0), .out(n13421_1));
wire n13422; //CHANY 4 (4,3) #52
wire n13422_0;
wire n13422_1;
buffer_wire buffer_13422_1 (.in(n13422_0), .out(n13422_1));
wire n13423; //CHANY 4 (4,3) #53
wire n13423_0;
wire n13423_1;
buffer_wire buffer_13423_1 (.in(n13423_0), .out(n13423_1));
wire n13424; //CHANY 4 (4,3) #60
wire n13424_0;
wire n13424_1;
buffer_wire buffer_13424_1 (.in(n13424_0), .out(n13424_1));
wire n13425; //CHANY 4 (4,3) #61
wire n13425_0;
wire n13425_1;
buffer_wire buffer_13425_1 (.in(n13425_0), .out(n13425_1));
wire n13426; //CHANY 4 (4,3) #68
wire n13426_0;
wire n13426_1;
buffer_wire buffer_13426_1 (.in(n13426_0), .out(n13426_1));
wire n13427; //CHANY 4 (4,3) #69
wire n13427_0;
wire n13427_1;
buffer_wire buffer_13427_1 (.in(n13427_0), .out(n13427_1));
wire n13428; //CHANY 4 (4,3) #76
wire n13428_0;
wire n13428_1;
buffer_wire buffer_13428_1 (.in(n13428_0), .out(n13428_1));
wire n13429; //CHANY 4 (4,3) #77
wire n13429_0;
wire n13429_1;
buffer_wire buffer_13429_1 (.in(n13429_0), .out(n13429_1));
wire n13430; //CHANY 4 (4,4) #6
wire n13430_0;
wire n13430_1;
buffer_wire buffer_13430_1 (.in(n13430_0), .out(n13430_1));
wire n13431; //CHANY 4 (4,4) #7
wire n13431_0;
wire n13431_1;
buffer_wire buffer_13431_1 (.in(n13431_0), .out(n13431_1));
wire n13432; //CHANY 4 (4,4) #14
wire n13432_0;
wire n13432_1;
buffer_wire buffer_13432_1 (.in(n13432_0), .out(n13432_1));
wire n13433; //CHANY 4 (4,4) #15
wire n13433_0;
wire n13433_1;
buffer_wire buffer_13433_1 (.in(n13433_0), .out(n13433_1));
wire n13434; //CHANY 4 (4,4) #22
wire n13434_0;
wire n13434_1;
buffer_wire buffer_13434_1 (.in(n13434_0), .out(n13434_1));
wire n13435; //CHANY 4 (4,4) #23
wire n13435_0;
wire n13435_1;
buffer_wire buffer_13435_1 (.in(n13435_0), .out(n13435_1));
wire n13436; //CHANY 4 (4,4) #30
wire n13436_0;
wire n13436_1;
buffer_wire buffer_13436_1 (.in(n13436_0), .out(n13436_1));
wire n13437; //CHANY 4 (4,4) #31
wire n13437_0;
wire n13437_1;
buffer_wire buffer_13437_1 (.in(n13437_0), .out(n13437_1));
wire n13438; //CHANY 4 (4,4) #38
wire n13438_0;
wire n13438_1;
buffer_wire buffer_13438_1 (.in(n13438_0), .out(n13438_1));
wire n13439; //CHANY 4 (4,4) #39
wire n13439_0;
wire n13439_1;
buffer_wire buffer_13439_1 (.in(n13439_0), .out(n13439_1));
wire n13440; //CHANY 4 (4,4) #46
wire n13440_0;
wire n13440_1;
buffer_wire buffer_13440_1 (.in(n13440_0), .out(n13440_1));
wire n13441; //CHANY 4 (4,4) #47
wire n13441_0;
wire n13441_1;
buffer_wire buffer_13441_1 (.in(n13441_0), .out(n13441_1));
wire n13442; //CHANY 4 (4,4) #54
wire n13442_0;
wire n13442_1;
buffer_wire buffer_13442_1 (.in(n13442_0), .out(n13442_1));
wire n13443; //CHANY 4 (4,4) #55
wire n13443_0;
wire n13443_1;
buffer_wire buffer_13443_1 (.in(n13443_0), .out(n13443_1));
wire n13444; //CHANY 4 (4,4) #62
wire n13444_0;
wire n13444_1;
buffer_wire buffer_13444_1 (.in(n13444_0), .out(n13444_1));
wire n13445; //CHANY 4 (4,4) #63
wire n13445_0;
wire n13445_1;
buffer_wire buffer_13445_1 (.in(n13445_0), .out(n13445_1));
wire n13446; //CHANY 4 (4,4) #70
wire n13446_0;
wire n13446_1;
buffer_wire buffer_13446_1 (.in(n13446_0), .out(n13446_1));
wire n13447; //CHANY 4 (4,4) #71
wire n13447_0;
wire n13447_1;
buffer_wire buffer_13447_1 (.in(n13447_0), .out(n13447_1));
wire n13448; //CHANY 4 (4,4) #78
wire n13448_0;
wire n13448_1;
buffer_wire buffer_13448_1 (.in(n13448_0), .out(n13448_1));
wire n13449; //CHANY 4 (4,4) #79
wire n13449_0;
wire n13449_1;
buffer_wire buffer_13449_1 (.in(n13449_0), .out(n13449_1));
wire n13450; //CHANY 4 (4,5) #0
wire n13450_0;
wire n13450_1;
buffer_wire buffer_13450_1 (.in(n13450_0), .out(n13450_1));
wire n13451; //CHANY 4 (4,5) #1
wire n13451_0;
wire n13451_1;
buffer_wire buffer_13451_1 (.in(n13451_0), .out(n13451_1));
wire n13452; //CHANY 4 (4,5) #8
wire n13452_0;
wire n13452_1;
buffer_wire buffer_13452_1 (.in(n13452_0), .out(n13452_1));
wire n13453; //CHANY 4 (4,5) #9
wire n13453_0;
wire n13453_1;
buffer_wire buffer_13453_1 (.in(n13453_0), .out(n13453_1));
wire n13454; //CHANY 4 (4,5) #16
wire n13454_0;
wire n13454_1;
buffer_wire buffer_13454_1 (.in(n13454_0), .out(n13454_1));
wire n13455; //CHANY 4 (4,5) #17
wire n13455_0;
wire n13455_1;
buffer_wire buffer_13455_1 (.in(n13455_0), .out(n13455_1));
wire n13456; //CHANY 4 (4,5) #24
wire n13456_0;
wire n13456_1;
buffer_wire buffer_13456_1 (.in(n13456_0), .out(n13456_1));
wire n13457; //CHANY 4 (4,5) #25
wire n13457_0;
wire n13457_1;
buffer_wire buffer_13457_1 (.in(n13457_0), .out(n13457_1));
wire n13458; //CHANY 4 (4,5) #32
wire n13458_0;
wire n13458_1;
buffer_wire buffer_13458_1 (.in(n13458_0), .out(n13458_1));
wire n13459; //CHANY 4 (4,5) #33
wire n13459_0;
wire n13459_1;
buffer_wire buffer_13459_1 (.in(n13459_0), .out(n13459_1));
wire n13460; //CHANY 4 (4,5) #40
wire n13460_0;
wire n13460_1;
buffer_wire buffer_13460_1 (.in(n13460_0), .out(n13460_1));
wire n13461; //CHANY 4 (4,5) #41
wire n13461_0;
wire n13461_1;
buffer_wire buffer_13461_1 (.in(n13461_0), .out(n13461_1));
wire n13462; //CHANY 4 (4,5) #48
wire n13462_0;
wire n13462_1;
buffer_wire buffer_13462_1 (.in(n13462_0), .out(n13462_1));
wire n13463; //CHANY 4 (4,5) #49
wire n13463_0;
wire n13463_1;
buffer_wire buffer_13463_1 (.in(n13463_0), .out(n13463_1));
wire n13464; //CHANY 4 (4,5) #56
wire n13464_0;
wire n13464_1;
buffer_wire buffer_13464_1 (.in(n13464_0), .out(n13464_1));
wire n13465; //CHANY 4 (4,5) #57
wire n13465_0;
wire n13465_1;
buffer_wire buffer_13465_1 (.in(n13465_0), .out(n13465_1));
wire n13466; //CHANY 4 (4,5) #64
wire n13466_0;
wire n13466_1;
buffer_wire buffer_13466_1 (.in(n13466_0), .out(n13466_1));
wire n13467; //CHANY 4 (4,5) #65
wire n13467_0;
wire n13467_1;
buffer_wire buffer_13467_1 (.in(n13467_0), .out(n13467_1));
wire n13468; //CHANY 4 (4,5) #72
wire n13468_0;
wire n13468_1;
buffer_wire buffer_13468_1 (.in(n13468_0), .out(n13468_1));
wire n13469; //CHANY 4 (4,5) #73
wire n13469_0;
wire n13469_1;
buffer_wire buffer_13469_1 (.in(n13469_0), .out(n13469_1));
wire n13470; //CHANY 5 (4,5) #80
wire n13470_0;
wire n13470_1;
buffer_wire buffer_13470_1 (.in(n13470_0), .out(n13470_1));
wire n13471; //CHANY 5 (4,5) #81
wire n13471_0;
wire n13471_1;
buffer_wire buffer_13471_1 (.in(n13471_0), .out(n13471_1));
wire n13472; //CHANY 4 (4,6) #2
wire n13472_0;
wire n13472_1;
buffer_wire buffer_13472_1 (.in(n13472_0), .out(n13472_1));
wire n13473; //CHANY 4 (4,6) #3
wire n13473_0;
wire n13473_1;
buffer_wire buffer_13473_1 (.in(n13473_0), .out(n13473_1));
wire n13474; //CHANY 4 (4,6) #10
wire n13474_0;
wire n13474_1;
buffer_wire buffer_13474_1 (.in(n13474_0), .out(n13474_1));
wire n13475; //CHANY 4 (4,6) #11
wire n13475_0;
wire n13475_1;
buffer_wire buffer_13475_1 (.in(n13475_0), .out(n13475_1));
wire n13476; //CHANY 4 (4,6) #18
wire n13476_0;
wire n13476_1;
buffer_wire buffer_13476_1 (.in(n13476_0), .out(n13476_1));
wire n13477; //CHANY 4 (4,6) #19
wire n13477_0;
wire n13477_1;
buffer_wire buffer_13477_1 (.in(n13477_0), .out(n13477_1));
wire n13478; //CHANY 4 (4,6) #26
wire n13478_0;
wire n13478_1;
buffer_wire buffer_13478_1 (.in(n13478_0), .out(n13478_1));
wire n13479; //CHANY 4 (4,6) #27
wire n13479_0;
wire n13479_1;
buffer_wire buffer_13479_1 (.in(n13479_0), .out(n13479_1));
wire n13480; //CHANY 4 (4,6) #34
wire n13480_0;
wire n13480_1;
buffer_wire buffer_13480_1 (.in(n13480_0), .out(n13480_1));
wire n13481; //CHANY 4 (4,6) #35
wire n13481_0;
wire n13481_1;
buffer_wire buffer_13481_1 (.in(n13481_0), .out(n13481_1));
wire n13482; //CHANY 4 (4,6) #42
wire n13482_0;
wire n13482_1;
buffer_wire buffer_13482_1 (.in(n13482_0), .out(n13482_1));
wire n13483; //CHANY 4 (4,6) #43
wire n13483_0;
wire n13483_1;
buffer_wire buffer_13483_1 (.in(n13483_0), .out(n13483_1));
wire n13484; //CHANY 4 (4,6) #50
wire n13484_0;
wire n13484_1;
buffer_wire buffer_13484_1 (.in(n13484_0), .out(n13484_1));
wire n13485; //CHANY 4 (4,6) #51
wire n13485_0;
wire n13485_1;
buffer_wire buffer_13485_1 (.in(n13485_0), .out(n13485_1));
wire n13486; //CHANY 4 (4,6) #58
wire n13486_0;
wire n13486_1;
buffer_wire buffer_13486_1 (.in(n13486_0), .out(n13486_1));
wire n13487; //CHANY 4 (4,6) #59
wire n13487_0;
wire n13487_1;
buffer_wire buffer_13487_1 (.in(n13487_0), .out(n13487_1));
wire n13488; //CHANY 4 (4,6) #66
wire n13488_0;
wire n13488_1;
buffer_wire buffer_13488_1 (.in(n13488_0), .out(n13488_1));
wire n13489; //CHANY 4 (4,6) #67
wire n13489_0;
wire n13489_1;
buffer_wire buffer_13489_1 (.in(n13489_0), .out(n13489_1));
wire n13490; //CHANY 4 (4,6) #74
wire n13490_0;
wire n13490_1;
buffer_wire buffer_13490_1 (.in(n13490_0), .out(n13490_1));
wire n13491; //CHANY 4 (4,6) #75
wire n13491_0;
wire n13491_1;
buffer_wire buffer_13491_1 (.in(n13491_0), .out(n13491_1));
wire n13492; //CHANY 4 (4,6) #82
wire n13492_0;
wire n13492_1;
buffer_wire buffer_13492_1 (.in(n13492_0), .out(n13492_1));
wire n13493; //CHANY 4 (4,6) #83
wire n13493_0;
wire n13493_1;
buffer_wire buffer_13493_1 (.in(n13493_0), .out(n13493_1));
wire n13494; //CHANY 3 (4,7) #4
wire n13494_0;
wire n13495; //CHANY 3 (4,7) #5
wire n13495_0;
wire n13496; //CHANY 3 (4,7) #12
wire n13496_0;
wire n13497; //CHANY 3 (4,7) #13
wire n13497_0;
wire n13498; //CHANY 3 (4,7) #20
wire n13498_0;
wire n13499; //CHANY 3 (4,7) #21
wire n13499_0;
wire n13500; //CHANY 3 (4,7) #28
wire n13500_0;
wire n13501; //CHANY 3 (4,7) #29
wire n13501_0;
wire n13502; //CHANY 3 (4,7) #36
wire n13502_0;
wire n13503; //CHANY 3 (4,7) #37
wire n13503_0;
wire n13504; //CHANY 3 (4,7) #44
wire n13504_0;
wire n13505; //CHANY 3 (4,7) #45
wire n13505_0;
wire n13506; //CHANY 3 (4,7) #52
wire n13506_0;
wire n13507; //CHANY 3 (4,7) #53
wire n13507_0;
wire n13508; //CHANY 3 (4,7) #60
wire n13508_0;
wire n13509; //CHANY 3 (4,7) #61
wire n13509_0;
wire n13510; //CHANY 3 (4,7) #68
wire n13510_0;
wire n13511; //CHANY 3 (4,7) #69
wire n13511_0;
wire n13512; //CHANY 3 (4,7) #76
wire n13512_0;
wire n13513; //CHANY 3 (4,7) #77
wire n13513_0;
wire n13514; //CHANY 3 (4,7) #84
wire n13514_0;
wire n13515; //CHANY 3 (4,7) #85
wire n13515_0;
wire n13516; //CHANY 2 (4,8) #6
wire n13516_0;
wire n13517; //CHANY 2 (4,8) #7
wire n13517_0;
wire n13518; //CHANY 2 (4,8) #14
wire n13518_0;
wire n13519; //CHANY 2 (4,8) #15
wire n13519_0;
wire n13520; //CHANY 2 (4,8) #22
wire n13520_0;
wire n13521; //CHANY 2 (4,8) #23
wire n13521_0;
wire n13522; //CHANY 2 (4,8) #30
wire n13522_0;
wire n13523; //CHANY 2 (4,8) #31
wire n13523_0;
wire n13524; //CHANY 2 (4,8) #38
wire n13524_0;
wire n13525; //CHANY 2 (4,8) #39
wire n13525_0;
wire n13526; //CHANY 2 (4,8) #46
wire n13526_0;
wire n13527; //CHANY 2 (4,8) #47
wire n13527_0;
wire n13528; //CHANY 2 (4,8) #54
wire n13528_0;
wire n13529; //CHANY 2 (4,8) #55
wire n13529_0;
wire n13530; //CHANY 2 (4,8) #62
wire n13530_0;
wire n13531; //CHANY 2 (4,8) #63
wire n13531_0;
wire n13532; //CHANY 2 (4,8) #70
wire n13532_0;
wire n13533; //CHANY 2 (4,8) #71
wire n13533_0;
wire n13534; //CHANY 2 (4,8) #78
wire n13534_0;
wire n13535; //CHANY 2 (4,8) #79
wire n13535_0;
wire n13536; //CHANY 2 (4,8) #86
wire n13536_0;
wire n13537; //CHANY 2 (4,8) #87
wire n13537_0;
wire n13538; //CHANY 1 (4,9) #0
wire n13538_0;
wire n13539; //CHANY 1 (4,9) #1
wire n13539_0;
wire n13540; //CHANY 1 (4,9) #8
wire n13540_0;
wire n13541; //CHANY 1 (4,9) #9
wire n13541_0;
wire n13542; //CHANY 1 (4,9) #16
wire n13542_0;
wire n13543; //CHANY 1 (4,9) #17
wire n13543_0;
wire n13544; //CHANY 1 (4,9) #24
wire n13544_0;
wire n13545; //CHANY 1 (4,9) #25
wire n13545_0;
wire n13546; //CHANY 1 (4,9) #32
wire n13546_0;
wire n13547; //CHANY 1 (4,9) #33
wire n13547_0;
wire n13548; //CHANY 1 (4,9) #40
wire n13548_0;
wire n13549; //CHANY 1 (4,9) #41
wire n13549_0;
wire n13550; //CHANY 1 (4,9) #48
wire n13550_0;
wire n13551; //CHANY 1 (4,9) #49
wire n13551_0;
wire n13552; //CHANY 1 (4,9) #56
wire n13552_0;
wire n13553; //CHANY 1 (4,9) #57
wire n13553_0;
wire n13554; //CHANY 1 (4,9) #64
wire n13554_0;
wire n13555; //CHANY 1 (4,9) #65
wire n13555_0;
wire n13556; //CHANY 1 (4,9) #72
wire n13556_0;
wire n13557; //CHANY 1 (4,9) #73
wire n13557_0;
wire n13558; //CHANY 1 (4,9) #88
wire n13558_0;
wire n13559; //CHANY 1 (4,9) #89
wire n13559_0;
wire n13560; //CHANY 3 (5,1) #0
wire n13560_0;
wire n13561; //CHANY 3 (5,1) #1
wire n13561_0;
wire n13562; //CHANY 4 (5,1) #2
wire n13562_0;
wire n13562_1;
buffer_wire buffer_13562_1 (.in(n13562_0), .out(n13562_1));
wire n13563; //CHANY 4 (5,1) #3
wire n13563_0;
wire n13563_1;
buffer_wire buffer_13563_1 (.in(n13563_0), .out(n13563_1));
wire n13564; //CHANY 1 (5,1) #4
wire n13564_0;
wire n13565; //CHANY 1 (5,1) #5
wire n13565_0;
wire n13566; //CHANY 2 (5,1) #6
wire n13566_0;
wire n13567; //CHANY 2 (5,1) #7
wire n13567_0;
wire n13568; //CHANY 3 (5,1) #8
wire n13568_0;
wire n13569; //CHANY 3 (5,1) #9
wire n13569_0;
wire n13570; //CHANY 4 (5,1) #10
wire n13570_0;
wire n13570_1;
buffer_wire buffer_13570_1 (.in(n13570_0), .out(n13570_1));
wire n13571; //CHANY 4 (5,1) #11
wire n13571_0;
wire n13571_1;
buffer_wire buffer_13571_1 (.in(n13571_0), .out(n13571_1));
wire n13572; //CHANY 1 (5,1) #12
wire n13572_0;
wire n13573; //CHANY 1 (5,1) #13
wire n13573_0;
wire n13574; //CHANY 2 (5,1) #14
wire n13574_0;
wire n13575; //CHANY 2 (5,1) #15
wire n13575_0;
wire n13576; //CHANY 3 (5,1) #16
wire n13576_0;
wire n13577; //CHANY 3 (5,1) #17
wire n13577_0;
wire n13578; //CHANY 4 (5,1) #18
wire n13578_0;
wire n13578_1;
buffer_wire buffer_13578_1 (.in(n13578_0), .out(n13578_1));
wire n13579; //CHANY 4 (5,1) #19
wire n13579_0;
wire n13579_1;
buffer_wire buffer_13579_1 (.in(n13579_0), .out(n13579_1));
wire n13580; //CHANY 1 (5,1) #20
wire n13580_0;
wire n13581; //CHANY 1 (5,1) #21
wire n13581_0;
wire n13582; //CHANY 2 (5,1) #22
wire n13582_0;
wire n13583; //CHANY 2 (5,1) #23
wire n13583_0;
wire n13584; //CHANY 3 (5,1) #24
wire n13584_0;
wire n13585; //CHANY 3 (5,1) #25
wire n13585_0;
wire n13586; //CHANY 4 (5,1) #26
wire n13586_0;
wire n13586_1;
buffer_wire buffer_13586_1 (.in(n13586_0), .out(n13586_1));
wire n13587; //CHANY 4 (5,1) #27
wire n13587_0;
wire n13587_1;
buffer_wire buffer_13587_1 (.in(n13587_0), .out(n13587_1));
wire n13588; //CHANY 1 (5,1) #28
wire n13588_0;
wire n13589; //CHANY 1 (5,1) #29
wire n13589_0;
wire n13590; //CHANY 2 (5,1) #30
wire n13590_0;
wire n13591; //CHANY 2 (5,1) #31
wire n13591_0;
wire n13592; //CHANY 3 (5,1) #32
wire n13592_0;
wire n13593; //CHANY 3 (5,1) #33
wire n13593_0;
wire n13594; //CHANY 4 (5,1) #34
wire n13594_0;
wire n13594_1;
buffer_wire buffer_13594_1 (.in(n13594_0), .out(n13594_1));
wire n13595; //CHANY 4 (5,1) #35
wire n13595_0;
wire n13595_1;
buffer_wire buffer_13595_1 (.in(n13595_0), .out(n13595_1));
wire n13596; //CHANY 1 (5,1) #36
wire n13596_0;
wire n13597; //CHANY 1 (5,1) #37
wire n13597_0;
wire n13598; //CHANY 2 (5,1) #38
wire n13598_0;
wire n13599; //CHANY 2 (5,1) #39
wire n13599_0;
wire n13600; //CHANY 3 (5,1) #40
wire n13600_0;
wire n13601; //CHANY 3 (5,1) #41
wire n13601_0;
wire n13602; //CHANY 4 (5,1) #42
wire n13602_0;
wire n13602_1;
buffer_wire buffer_13602_1 (.in(n13602_0), .out(n13602_1));
wire n13603; //CHANY 4 (5,1) #43
wire n13603_0;
wire n13603_1;
buffer_wire buffer_13603_1 (.in(n13603_0), .out(n13603_1));
wire n13604; //CHANY 1 (5,1) #44
wire n13604_0;
wire n13605; //CHANY 1 (5,1) #45
wire n13605_0;
wire n13606; //CHANY 2 (5,1) #46
wire n13606_0;
wire n13607; //CHANY 2 (5,1) #47
wire n13607_0;
wire n13608; //CHANY 3 (5,1) #48
wire n13608_0;
wire n13609; //CHANY 3 (5,1) #49
wire n13609_0;
wire n13610; //CHANY 4 (5,1) #50
wire n13610_0;
wire n13610_1;
buffer_wire buffer_13610_1 (.in(n13610_0), .out(n13610_1));
wire n13611; //CHANY 4 (5,1) #51
wire n13611_0;
wire n13611_1;
buffer_wire buffer_13611_1 (.in(n13611_0), .out(n13611_1));
wire n13612; //CHANY 1 (5,1) #52
wire n13612_0;
wire n13613; //CHANY 1 (5,1) #53
wire n13613_0;
wire n13614; //CHANY 2 (5,1) #54
wire n13614_0;
wire n13615; //CHANY 2 (5,1) #55
wire n13615_0;
wire n13616; //CHANY 3 (5,1) #56
wire n13616_0;
wire n13617; //CHANY 3 (5,1) #57
wire n13617_0;
wire n13618; //CHANY 4 (5,1) #58
wire n13618_0;
wire n13618_1;
buffer_wire buffer_13618_1 (.in(n13618_0), .out(n13618_1));
wire n13619; //CHANY 4 (5,1) #59
wire n13619_0;
wire n13619_1;
buffer_wire buffer_13619_1 (.in(n13619_0), .out(n13619_1));
wire n13620; //CHANY 1 (5,1) #60
wire n13620_0;
wire n13621; //CHANY 1 (5,1) #61
wire n13621_0;
wire n13622; //CHANY 2 (5,1) #62
wire n13622_0;
wire n13623; //CHANY 2 (5,1) #63
wire n13623_0;
wire n13624; //CHANY 3 (5,1) #64
wire n13624_0;
wire n13625; //CHANY 3 (5,1) #65
wire n13625_0;
wire n13626; //CHANY 4 (5,1) #66
wire n13626_0;
wire n13626_1;
buffer_wire buffer_13626_1 (.in(n13626_0), .out(n13626_1));
wire n13627; //CHANY 4 (5,1) #67
wire n13627_0;
wire n13627_1;
buffer_wire buffer_13627_1 (.in(n13627_0), .out(n13627_1));
wire n13628; //CHANY 1 (5,1) #68
wire n13628_0;
wire n13629; //CHANY 1 (5,1) #69
wire n13629_0;
wire n13630; //CHANY 2 (5,1) #70
wire n13630_0;
wire n13631; //CHANY 2 (5,1) #71
wire n13631_0;
wire n13632; //CHANY 3 (5,1) #72
wire n13632_0;
wire n13633; //CHANY 3 (5,1) #73
wire n13633_0;
wire n13634; //CHANY 4 (5,1) #74
wire n13634_0;
wire n13634_1;
buffer_wire buffer_13634_1 (.in(n13634_0), .out(n13634_1));
wire n13635; //CHANY 4 (5,1) #75
wire n13635_0;
wire n13635_1;
buffer_wire buffer_13635_1 (.in(n13635_0), .out(n13635_1));
wire n13636; //CHANY 1 (5,1) #76
wire n13636_0;
wire n13637; //CHANY 1 (5,1) #77
wire n13637_0;
wire n13638; //CHANY 2 (5,1) #78
wire n13638_0;
wire n13639; //CHANY 2 (5,1) #79
wire n13639_0;
wire n13640; //CHANY 3 (5,1) #80
wire n13640_0;
wire n13641; //CHANY 3 (5,1) #81
wire n13641_0;
wire n13642; //CHANY 4 (5,1) #82
wire n13642_0;
wire n13642_1;
buffer_wire buffer_13642_1 (.in(n13642_0), .out(n13642_1));
wire n13643; //CHANY 4 (5,1) #83
wire n13643_0;
wire n13643_1;
buffer_wire buffer_13643_1 (.in(n13643_0), .out(n13643_1));
wire n13644; //CHANY 5 (5,1) #84
wire n13644_0;
wire n13644_1;
buffer_wire buffer_13644_1 (.in(n13644_0), .out(n13644_1));
wire n13645; //CHANY 5 (5,1) #85
wire n13645_0;
wire n13645_1;
buffer_wire buffer_13645_1 (.in(n13645_0), .out(n13645_1));
wire n13646; //CHANY 6 (5,1) #86
wire n13646_0;
wire n13646_1;
buffer_wire buffer_13646_1 (.in(n13646_0), .out(n13646_1));
wire n13647; //CHANY 6 (5,1) #87
wire n13647_0;
wire n13647_1;
buffer_wire buffer_13647_1 (.in(n13647_0), .out(n13647_1));
wire n13648; //CHANY 7 (5,1) #88
wire n13648_0;
wire n13648_1;
wire n13648_2;
buffer_wire buffer_13648_2 (.in(n13648_1), .out(n13648_2));
buffer_wire buffer_13648_1 (.in(n13648_0), .out(n13648_1));
wire n13649; //CHANY 7 (5,1) #89
wire n13649_0;
wire n13649_1;
wire n13649_2;
buffer_wire buffer_13649_2 (.in(n13649_1), .out(n13649_2));
buffer_wire buffer_13649_1 (.in(n13649_0), .out(n13649_1));
wire n13650; //CHANY 8 (5,1) #90
wire n13650_0;
wire n13650_1;
wire n13650_2;
buffer_wire buffer_13650_2 (.in(n13650_1), .out(n13650_2));
buffer_wire buffer_13650_1 (.in(n13650_0), .out(n13650_1));
wire n13651; //CHANY 8 (5,1) #91
wire n13651_0;
wire n13651_1;
wire n13651_2;
buffer_wire buffer_13651_2 (.in(n13651_1), .out(n13651_2));
buffer_wire buffer_13651_1 (.in(n13651_0), .out(n13651_1));
wire n13652; //CHANY 4 (5,2) #4
wire n13652_0;
wire n13652_1;
buffer_wire buffer_13652_1 (.in(n13652_0), .out(n13652_1));
wire n13653; //CHANY 4 (5,2) #5
wire n13653_0;
wire n13653_1;
buffer_wire buffer_13653_1 (.in(n13653_0), .out(n13653_1));
wire n13654; //CHANY 4 (5,2) #12
wire n13654_0;
wire n13654_1;
buffer_wire buffer_13654_1 (.in(n13654_0), .out(n13654_1));
wire n13655; //CHANY 4 (5,2) #13
wire n13655_0;
wire n13655_1;
buffer_wire buffer_13655_1 (.in(n13655_0), .out(n13655_1));
wire n13656; //CHANY 4 (5,2) #20
wire n13656_0;
wire n13656_1;
buffer_wire buffer_13656_1 (.in(n13656_0), .out(n13656_1));
wire n13657; //CHANY 4 (5,2) #21
wire n13657_0;
wire n13657_1;
buffer_wire buffer_13657_1 (.in(n13657_0), .out(n13657_1));
wire n13658; //CHANY 4 (5,2) #28
wire n13658_0;
wire n13658_1;
buffer_wire buffer_13658_1 (.in(n13658_0), .out(n13658_1));
wire n13659; //CHANY 4 (5,2) #29
wire n13659_0;
wire n13659_1;
buffer_wire buffer_13659_1 (.in(n13659_0), .out(n13659_1));
wire n13660; //CHANY 4 (5,2) #36
wire n13660_0;
wire n13660_1;
buffer_wire buffer_13660_1 (.in(n13660_0), .out(n13660_1));
wire n13661; //CHANY 4 (5,2) #37
wire n13661_0;
wire n13661_1;
buffer_wire buffer_13661_1 (.in(n13661_0), .out(n13661_1));
wire n13662; //CHANY 4 (5,2) #44
wire n13662_0;
wire n13662_1;
buffer_wire buffer_13662_1 (.in(n13662_0), .out(n13662_1));
wire n13663; //CHANY 4 (5,2) #45
wire n13663_0;
wire n13663_1;
buffer_wire buffer_13663_1 (.in(n13663_0), .out(n13663_1));
wire n13664; //CHANY 4 (5,2) #52
wire n13664_0;
wire n13664_1;
buffer_wire buffer_13664_1 (.in(n13664_0), .out(n13664_1));
wire n13665; //CHANY 4 (5,2) #53
wire n13665_0;
wire n13665_1;
buffer_wire buffer_13665_1 (.in(n13665_0), .out(n13665_1));
wire n13666; //CHANY 4 (5,2) #60
wire n13666_0;
wire n13666_1;
buffer_wire buffer_13666_1 (.in(n13666_0), .out(n13666_1));
wire n13667; //CHANY 4 (5,2) #61
wire n13667_0;
wire n13667_1;
buffer_wire buffer_13667_1 (.in(n13667_0), .out(n13667_1));
wire n13668; //CHANY 4 (5,2) #68
wire n13668_0;
wire n13668_1;
buffer_wire buffer_13668_1 (.in(n13668_0), .out(n13668_1));
wire n13669; //CHANY 4 (5,2) #69
wire n13669_0;
wire n13669_1;
buffer_wire buffer_13669_1 (.in(n13669_0), .out(n13669_1));
wire n13670; //CHANY 4 (5,2) #76
wire n13670_0;
wire n13670_1;
buffer_wire buffer_13670_1 (.in(n13670_0), .out(n13670_1));
wire n13671; //CHANY 4 (5,2) #77
wire n13671_0;
wire n13671_1;
buffer_wire buffer_13671_1 (.in(n13671_0), .out(n13671_1));
wire n13672; //CHANY 4 (5,3) #6
wire n13672_0;
wire n13672_1;
buffer_wire buffer_13672_1 (.in(n13672_0), .out(n13672_1));
wire n13673; //CHANY 4 (5,3) #7
wire n13673_0;
wire n13673_1;
buffer_wire buffer_13673_1 (.in(n13673_0), .out(n13673_1));
wire n13674; //CHANY 4 (5,3) #14
wire n13674_0;
wire n13674_1;
buffer_wire buffer_13674_1 (.in(n13674_0), .out(n13674_1));
wire n13675; //CHANY 4 (5,3) #15
wire n13675_0;
wire n13675_1;
buffer_wire buffer_13675_1 (.in(n13675_0), .out(n13675_1));
wire n13676; //CHANY 4 (5,3) #22
wire n13676_0;
wire n13676_1;
buffer_wire buffer_13676_1 (.in(n13676_0), .out(n13676_1));
wire n13677; //CHANY 4 (5,3) #23
wire n13677_0;
wire n13677_1;
buffer_wire buffer_13677_1 (.in(n13677_0), .out(n13677_1));
wire n13678; //CHANY 4 (5,3) #30
wire n13678_0;
wire n13678_1;
buffer_wire buffer_13678_1 (.in(n13678_0), .out(n13678_1));
wire n13679; //CHANY 4 (5,3) #31
wire n13679_0;
wire n13679_1;
buffer_wire buffer_13679_1 (.in(n13679_0), .out(n13679_1));
wire n13680; //CHANY 4 (5,3) #38
wire n13680_0;
wire n13680_1;
buffer_wire buffer_13680_1 (.in(n13680_0), .out(n13680_1));
wire n13681; //CHANY 4 (5,3) #39
wire n13681_0;
wire n13681_1;
buffer_wire buffer_13681_1 (.in(n13681_0), .out(n13681_1));
wire n13682; //CHANY 4 (5,3) #46
wire n13682_0;
wire n13682_1;
buffer_wire buffer_13682_1 (.in(n13682_0), .out(n13682_1));
wire n13683; //CHANY 4 (5,3) #47
wire n13683_0;
wire n13683_1;
buffer_wire buffer_13683_1 (.in(n13683_0), .out(n13683_1));
wire n13684; //CHANY 4 (5,3) #54
wire n13684_0;
wire n13684_1;
buffer_wire buffer_13684_1 (.in(n13684_0), .out(n13684_1));
wire n13685; //CHANY 4 (5,3) #55
wire n13685_0;
wire n13685_1;
buffer_wire buffer_13685_1 (.in(n13685_0), .out(n13685_1));
wire n13686; //CHANY 4 (5,3) #62
wire n13686_0;
wire n13686_1;
buffer_wire buffer_13686_1 (.in(n13686_0), .out(n13686_1));
wire n13687; //CHANY 4 (5,3) #63
wire n13687_0;
wire n13687_1;
buffer_wire buffer_13687_1 (.in(n13687_0), .out(n13687_1));
wire n13688; //CHANY 4 (5,3) #70
wire n13688_0;
wire n13688_1;
buffer_wire buffer_13688_1 (.in(n13688_0), .out(n13688_1));
wire n13689; //CHANY 4 (5,3) #71
wire n13689_0;
wire n13689_1;
buffer_wire buffer_13689_1 (.in(n13689_0), .out(n13689_1));
wire n13690; //CHANY 4 (5,3) #78
wire n13690_0;
wire n13690_1;
buffer_wire buffer_13690_1 (.in(n13690_0), .out(n13690_1));
wire n13691; //CHANY 4 (5,3) #79
wire n13691_0;
wire n13691_1;
buffer_wire buffer_13691_1 (.in(n13691_0), .out(n13691_1));
wire n13692; //CHANY 4 (5,4) #0
wire n13692_0;
wire n13692_1;
buffer_wire buffer_13692_1 (.in(n13692_0), .out(n13692_1));
wire n13693; //CHANY 4 (5,4) #1
wire n13693_0;
wire n13693_1;
buffer_wire buffer_13693_1 (.in(n13693_0), .out(n13693_1));
wire n13694; //CHANY 4 (5,4) #8
wire n13694_0;
wire n13694_1;
buffer_wire buffer_13694_1 (.in(n13694_0), .out(n13694_1));
wire n13695; //CHANY 4 (5,4) #9
wire n13695_0;
wire n13695_1;
buffer_wire buffer_13695_1 (.in(n13695_0), .out(n13695_1));
wire n13696; //CHANY 4 (5,4) #16
wire n13696_0;
wire n13696_1;
buffer_wire buffer_13696_1 (.in(n13696_0), .out(n13696_1));
wire n13697; //CHANY 4 (5,4) #17
wire n13697_0;
wire n13697_1;
buffer_wire buffer_13697_1 (.in(n13697_0), .out(n13697_1));
wire n13698; //CHANY 4 (5,4) #24
wire n13698_0;
wire n13698_1;
buffer_wire buffer_13698_1 (.in(n13698_0), .out(n13698_1));
wire n13699; //CHANY 4 (5,4) #25
wire n13699_0;
wire n13699_1;
buffer_wire buffer_13699_1 (.in(n13699_0), .out(n13699_1));
wire n13700; //CHANY 4 (5,4) #32
wire n13700_0;
wire n13700_1;
buffer_wire buffer_13700_1 (.in(n13700_0), .out(n13700_1));
wire n13701; //CHANY 4 (5,4) #33
wire n13701_0;
wire n13701_1;
buffer_wire buffer_13701_1 (.in(n13701_0), .out(n13701_1));
wire n13702; //CHANY 4 (5,4) #40
wire n13702_0;
wire n13702_1;
buffer_wire buffer_13702_1 (.in(n13702_0), .out(n13702_1));
wire n13703; //CHANY 4 (5,4) #41
wire n13703_0;
wire n13703_1;
buffer_wire buffer_13703_1 (.in(n13703_0), .out(n13703_1));
wire n13704; //CHANY 4 (5,4) #48
wire n13704_0;
wire n13704_1;
buffer_wire buffer_13704_1 (.in(n13704_0), .out(n13704_1));
wire n13705; //CHANY 4 (5,4) #49
wire n13705_0;
wire n13705_1;
buffer_wire buffer_13705_1 (.in(n13705_0), .out(n13705_1));
wire n13706; //CHANY 4 (5,4) #56
wire n13706_0;
wire n13706_1;
buffer_wire buffer_13706_1 (.in(n13706_0), .out(n13706_1));
wire n13707; //CHANY 4 (5,4) #57
wire n13707_0;
wire n13707_1;
buffer_wire buffer_13707_1 (.in(n13707_0), .out(n13707_1));
wire n13708; //CHANY 4 (5,4) #64
wire n13708_0;
wire n13708_1;
buffer_wire buffer_13708_1 (.in(n13708_0), .out(n13708_1));
wire n13709; //CHANY 4 (5,4) #65
wire n13709_0;
wire n13709_1;
buffer_wire buffer_13709_1 (.in(n13709_0), .out(n13709_1));
wire n13710; //CHANY 4 (5,4) #72
wire n13710_0;
wire n13710_1;
buffer_wire buffer_13710_1 (.in(n13710_0), .out(n13710_1));
wire n13711; //CHANY 4 (5,4) #73
wire n13711_0;
wire n13711_1;
buffer_wire buffer_13711_1 (.in(n13711_0), .out(n13711_1));
wire n13712; //CHANY 6 (5,4) #80
wire n13712_0;
wire n13712_1;
buffer_wire buffer_13712_1 (.in(n13712_0), .out(n13712_1));
wire n13713; //CHANY 6 (5,4) #81
wire n13713_0;
wire n13713_1;
buffer_wire buffer_13713_1 (.in(n13713_0), .out(n13713_1));
wire n13714; //CHANY 4 (5,5) #2
wire n13714_0;
wire n13714_1;
buffer_wire buffer_13714_1 (.in(n13714_0), .out(n13714_1));
wire n13715; //CHANY 4 (5,5) #3
wire n13715_0;
wire n13715_1;
buffer_wire buffer_13715_1 (.in(n13715_0), .out(n13715_1));
wire n13716; //CHANY 4 (5,5) #10
wire n13716_0;
wire n13716_1;
buffer_wire buffer_13716_1 (.in(n13716_0), .out(n13716_1));
wire n13717; //CHANY 4 (5,5) #11
wire n13717_0;
wire n13717_1;
buffer_wire buffer_13717_1 (.in(n13717_0), .out(n13717_1));
wire n13718; //CHANY 4 (5,5) #18
wire n13718_0;
wire n13718_1;
buffer_wire buffer_13718_1 (.in(n13718_0), .out(n13718_1));
wire n13719; //CHANY 4 (5,5) #19
wire n13719_0;
wire n13719_1;
buffer_wire buffer_13719_1 (.in(n13719_0), .out(n13719_1));
wire n13720; //CHANY 4 (5,5) #26
wire n13720_0;
wire n13720_1;
buffer_wire buffer_13720_1 (.in(n13720_0), .out(n13720_1));
wire n13721; //CHANY 4 (5,5) #27
wire n13721_0;
wire n13721_1;
buffer_wire buffer_13721_1 (.in(n13721_0), .out(n13721_1));
wire n13722; //CHANY 4 (5,5) #34
wire n13722_0;
wire n13722_1;
buffer_wire buffer_13722_1 (.in(n13722_0), .out(n13722_1));
wire n13723; //CHANY 4 (5,5) #35
wire n13723_0;
wire n13723_1;
buffer_wire buffer_13723_1 (.in(n13723_0), .out(n13723_1));
wire n13724; //CHANY 4 (5,5) #42
wire n13724_0;
wire n13724_1;
buffer_wire buffer_13724_1 (.in(n13724_0), .out(n13724_1));
wire n13725; //CHANY 4 (5,5) #43
wire n13725_0;
wire n13725_1;
buffer_wire buffer_13725_1 (.in(n13725_0), .out(n13725_1));
wire n13726; //CHANY 4 (5,5) #50
wire n13726_0;
wire n13726_1;
buffer_wire buffer_13726_1 (.in(n13726_0), .out(n13726_1));
wire n13727; //CHANY 4 (5,5) #51
wire n13727_0;
wire n13727_1;
buffer_wire buffer_13727_1 (.in(n13727_0), .out(n13727_1));
wire n13728; //CHANY 4 (5,5) #58
wire n13728_0;
wire n13728_1;
buffer_wire buffer_13728_1 (.in(n13728_0), .out(n13728_1));
wire n13729; //CHANY 4 (5,5) #59
wire n13729_0;
wire n13729_1;
buffer_wire buffer_13729_1 (.in(n13729_0), .out(n13729_1));
wire n13730; //CHANY 4 (5,5) #66
wire n13730_0;
wire n13730_1;
buffer_wire buffer_13730_1 (.in(n13730_0), .out(n13730_1));
wire n13731; //CHANY 4 (5,5) #67
wire n13731_0;
wire n13731_1;
buffer_wire buffer_13731_1 (.in(n13731_0), .out(n13731_1));
wire n13732; //CHANY 4 (5,5) #74
wire n13732_0;
wire n13732_1;
buffer_wire buffer_13732_1 (.in(n13732_0), .out(n13732_1));
wire n13733; //CHANY 4 (5,5) #75
wire n13733_0;
wire n13733_1;
buffer_wire buffer_13733_1 (.in(n13733_0), .out(n13733_1));
wire n13734; //CHANY 5 (5,5) #82
wire n13734_0;
wire n13734_1;
buffer_wire buffer_13734_1 (.in(n13734_0), .out(n13734_1));
wire n13735; //CHANY 5 (5,5) #83
wire n13735_0;
wire n13735_1;
buffer_wire buffer_13735_1 (.in(n13735_0), .out(n13735_1));
wire n13736; //CHANY 4 (5,6) #4
wire n13736_0;
wire n13736_1;
buffer_wire buffer_13736_1 (.in(n13736_0), .out(n13736_1));
wire n13737; //CHANY 4 (5,6) #5
wire n13737_0;
wire n13737_1;
buffer_wire buffer_13737_1 (.in(n13737_0), .out(n13737_1));
wire n13738; //CHANY 4 (5,6) #12
wire n13738_0;
wire n13738_1;
buffer_wire buffer_13738_1 (.in(n13738_0), .out(n13738_1));
wire n13739; //CHANY 4 (5,6) #13
wire n13739_0;
wire n13739_1;
buffer_wire buffer_13739_1 (.in(n13739_0), .out(n13739_1));
wire n13740; //CHANY 4 (5,6) #20
wire n13740_0;
wire n13740_1;
buffer_wire buffer_13740_1 (.in(n13740_0), .out(n13740_1));
wire n13741; //CHANY 4 (5,6) #21
wire n13741_0;
wire n13741_1;
buffer_wire buffer_13741_1 (.in(n13741_0), .out(n13741_1));
wire n13742; //CHANY 4 (5,6) #28
wire n13742_0;
wire n13742_1;
buffer_wire buffer_13742_1 (.in(n13742_0), .out(n13742_1));
wire n13743; //CHANY 4 (5,6) #29
wire n13743_0;
wire n13743_1;
buffer_wire buffer_13743_1 (.in(n13743_0), .out(n13743_1));
wire n13744; //CHANY 4 (5,6) #36
wire n13744_0;
wire n13744_1;
buffer_wire buffer_13744_1 (.in(n13744_0), .out(n13744_1));
wire n13745; //CHANY 4 (5,6) #37
wire n13745_0;
wire n13745_1;
buffer_wire buffer_13745_1 (.in(n13745_0), .out(n13745_1));
wire n13746; //CHANY 4 (5,6) #44
wire n13746_0;
wire n13746_1;
buffer_wire buffer_13746_1 (.in(n13746_0), .out(n13746_1));
wire n13747; //CHANY 4 (5,6) #45
wire n13747_0;
wire n13747_1;
buffer_wire buffer_13747_1 (.in(n13747_0), .out(n13747_1));
wire n13748; //CHANY 4 (5,6) #52
wire n13748_0;
wire n13748_1;
buffer_wire buffer_13748_1 (.in(n13748_0), .out(n13748_1));
wire n13749; //CHANY 4 (5,6) #53
wire n13749_0;
wire n13749_1;
buffer_wire buffer_13749_1 (.in(n13749_0), .out(n13749_1));
wire n13750; //CHANY 4 (5,6) #60
wire n13750_0;
wire n13750_1;
buffer_wire buffer_13750_1 (.in(n13750_0), .out(n13750_1));
wire n13751; //CHANY 4 (5,6) #61
wire n13751_0;
wire n13751_1;
buffer_wire buffer_13751_1 (.in(n13751_0), .out(n13751_1));
wire n13752; //CHANY 4 (5,6) #68
wire n13752_0;
wire n13752_1;
buffer_wire buffer_13752_1 (.in(n13752_0), .out(n13752_1));
wire n13753; //CHANY 4 (5,6) #69
wire n13753_0;
wire n13753_1;
buffer_wire buffer_13753_1 (.in(n13753_0), .out(n13753_1));
wire n13754; //CHANY 4 (5,6) #76
wire n13754_0;
wire n13754_1;
buffer_wire buffer_13754_1 (.in(n13754_0), .out(n13754_1));
wire n13755; //CHANY 4 (5,6) #77
wire n13755_0;
wire n13755_1;
buffer_wire buffer_13755_1 (.in(n13755_0), .out(n13755_1));
wire n13756; //CHANY 4 (5,6) #84
wire n13756_0;
wire n13756_1;
buffer_wire buffer_13756_1 (.in(n13756_0), .out(n13756_1));
wire n13757; //CHANY 4 (5,6) #85
wire n13757_0;
wire n13757_1;
buffer_wire buffer_13757_1 (.in(n13757_0), .out(n13757_1));
wire n13758; //CHANY 3 (5,7) #6
wire n13758_0;
wire n13759; //CHANY 3 (5,7) #7
wire n13759_0;
wire n13760; //CHANY 3 (5,7) #14
wire n13760_0;
wire n13761; //CHANY 3 (5,7) #15
wire n13761_0;
wire n13762; //CHANY 3 (5,7) #22
wire n13762_0;
wire n13763; //CHANY 3 (5,7) #23
wire n13763_0;
wire n13764; //CHANY 3 (5,7) #30
wire n13764_0;
wire n13765; //CHANY 3 (5,7) #31
wire n13765_0;
wire n13766; //CHANY 3 (5,7) #38
wire n13766_0;
wire n13767; //CHANY 3 (5,7) #39
wire n13767_0;
wire n13768; //CHANY 3 (5,7) #46
wire n13768_0;
wire n13769; //CHANY 3 (5,7) #47
wire n13769_0;
wire n13770; //CHANY 3 (5,7) #54
wire n13770_0;
wire n13771; //CHANY 3 (5,7) #55
wire n13771_0;
wire n13772; //CHANY 3 (5,7) #62
wire n13772_0;
wire n13773; //CHANY 3 (5,7) #63
wire n13773_0;
wire n13774; //CHANY 3 (5,7) #70
wire n13774_0;
wire n13775; //CHANY 3 (5,7) #71
wire n13775_0;
wire n13776; //CHANY 3 (5,7) #78
wire n13776_0;
wire n13777; //CHANY 3 (5,7) #79
wire n13777_0;
wire n13778; //CHANY 3 (5,7) #86
wire n13778_0;
wire n13779; //CHANY 3 (5,7) #87
wire n13779_0;
wire n13780; //CHANY 2 (5,8) #0
wire n13780_0;
wire n13781; //CHANY 2 (5,8) #1
wire n13781_0;
wire n13782; //CHANY 2 (5,8) #8
wire n13782_0;
wire n13783; //CHANY 2 (5,8) #9
wire n13783_0;
wire n13784; //CHANY 2 (5,8) #16
wire n13784_0;
wire n13785; //CHANY 2 (5,8) #17
wire n13785_0;
wire n13786; //CHANY 2 (5,8) #24
wire n13786_0;
wire n13787; //CHANY 2 (5,8) #25
wire n13787_0;
wire n13788; //CHANY 2 (5,8) #32
wire n13788_0;
wire n13789; //CHANY 2 (5,8) #33
wire n13789_0;
wire n13790; //CHANY 2 (5,8) #40
wire n13790_0;
wire n13791; //CHANY 2 (5,8) #41
wire n13791_0;
wire n13792; //CHANY 2 (5,8) #48
wire n13792_0;
wire n13793; //CHANY 2 (5,8) #49
wire n13793_0;
wire n13794; //CHANY 2 (5,8) #56
wire n13794_0;
wire n13795; //CHANY 2 (5,8) #57
wire n13795_0;
wire n13796; //CHANY 2 (5,8) #64
wire n13796_0;
wire n13797; //CHANY 2 (5,8) #65
wire n13797_0;
wire n13798; //CHANY 2 (5,8) #72
wire n13798_0;
wire n13799; //CHANY 2 (5,8) #73
wire n13799_0;
wire n13800; //CHANY 2 (5,8) #88
wire n13800_0;
wire n13801; //CHANY 2 (5,8) #89
wire n13801_0;
wire n13802; //CHANY 1 (5,9) #2
wire n13802_0;
wire n13803; //CHANY 1 (5,9) #3
wire n13803_0;
wire n13804; //CHANY 1 (5,9) #10
wire n13804_0;
wire n13805; //CHANY 1 (5,9) #11
wire n13805_0;
wire n13806; //CHANY 1 (5,9) #18
wire n13806_0;
wire n13807; //CHANY 1 (5,9) #19
wire n13807_0;
wire n13808; //CHANY 1 (5,9) #26
wire n13808_0;
wire n13809; //CHANY 1 (5,9) #27
wire n13809_0;
wire n13810; //CHANY 1 (5,9) #34
wire n13810_0;
wire n13811; //CHANY 1 (5,9) #35
wire n13811_0;
wire n13812; //CHANY 1 (5,9) #42
wire n13812_0;
wire n13813; //CHANY 1 (5,9) #43
wire n13813_0;
wire n13814; //CHANY 1 (5,9) #50
wire n13814_0;
wire n13815; //CHANY 1 (5,9) #51
wire n13815_0;
wire n13816; //CHANY 1 (5,9) #58
wire n13816_0;
wire n13817; //CHANY 1 (5,9) #59
wire n13817_0;
wire n13818; //CHANY 1 (5,9) #66
wire n13818_0;
wire n13819; //CHANY 1 (5,9) #67
wire n13819_0;
wire n13820; //CHANY 1 (5,9) #74
wire n13820_0;
wire n13821; //CHANY 1 (5,9) #75
wire n13821_0;
wire n13822; //CHANY 1 (5,9) #90
wire n13822_0;
wire n13823; //CHANY 1 (5,9) #91
wire n13823_0;
wire n13824; //CHANY 2 (6,1) #0
wire n13824_0;
wire n13825; //CHANY 2 (6,1) #1
wire n13825_0;
wire n13826; //CHANY 3 (6,1) #2
wire n13826_0;
wire n13827; //CHANY 3 (6,1) #3
wire n13827_0;
wire n13828; //CHANY 4 (6,1) #4
wire n13828_0;
wire n13828_1;
buffer_wire buffer_13828_1 (.in(n13828_0), .out(n13828_1));
wire n13829; //CHANY 4 (6,1) #5
wire n13829_0;
wire n13829_1;
buffer_wire buffer_13829_1 (.in(n13829_0), .out(n13829_1));
wire n13830; //CHANY 1 (6,1) #6
wire n13830_0;
wire n13831; //CHANY 1 (6,1) #7
wire n13831_0;
wire n13832; //CHANY 2 (6,1) #8
wire n13832_0;
wire n13833; //CHANY 2 (6,1) #9
wire n13833_0;
wire n13834; //CHANY 3 (6,1) #10
wire n13834_0;
wire n13835; //CHANY 3 (6,1) #11
wire n13835_0;
wire n13836; //CHANY 4 (6,1) #12
wire n13836_0;
wire n13836_1;
buffer_wire buffer_13836_1 (.in(n13836_0), .out(n13836_1));
wire n13837; //CHANY 4 (6,1) #13
wire n13837_0;
wire n13837_1;
buffer_wire buffer_13837_1 (.in(n13837_0), .out(n13837_1));
wire n13838; //CHANY 1 (6,1) #14
wire n13838_0;
wire n13839; //CHANY 1 (6,1) #15
wire n13839_0;
wire n13840; //CHANY 2 (6,1) #16
wire n13840_0;
wire n13841; //CHANY 2 (6,1) #17
wire n13841_0;
wire n13842; //CHANY 3 (6,1) #18
wire n13842_0;
wire n13843; //CHANY 3 (6,1) #19
wire n13843_0;
wire n13844; //CHANY 4 (6,1) #20
wire n13844_0;
wire n13844_1;
buffer_wire buffer_13844_1 (.in(n13844_0), .out(n13844_1));
wire n13845; //CHANY 4 (6,1) #21
wire n13845_0;
wire n13845_1;
buffer_wire buffer_13845_1 (.in(n13845_0), .out(n13845_1));
wire n13846; //CHANY 1 (6,1) #22
wire n13846_0;
wire n13847; //CHANY 1 (6,1) #23
wire n13847_0;
wire n13848; //CHANY 2 (6,1) #24
wire n13848_0;
wire n13849; //CHANY 2 (6,1) #25
wire n13849_0;
wire n13850; //CHANY 3 (6,1) #26
wire n13850_0;
wire n13851; //CHANY 3 (6,1) #27
wire n13851_0;
wire n13852; //CHANY 4 (6,1) #28
wire n13852_0;
wire n13852_1;
buffer_wire buffer_13852_1 (.in(n13852_0), .out(n13852_1));
wire n13853; //CHANY 4 (6,1) #29
wire n13853_0;
wire n13853_1;
buffer_wire buffer_13853_1 (.in(n13853_0), .out(n13853_1));
wire n13854; //CHANY 1 (6,1) #30
wire n13854_0;
wire n13855; //CHANY 1 (6,1) #31
wire n13855_0;
wire n13856; //CHANY 2 (6,1) #32
wire n13856_0;
wire n13857; //CHANY 2 (6,1) #33
wire n13857_0;
wire n13858; //CHANY 3 (6,1) #34
wire n13858_0;
wire n13859; //CHANY 3 (6,1) #35
wire n13859_0;
wire n13860; //CHANY 4 (6,1) #36
wire n13860_0;
wire n13860_1;
buffer_wire buffer_13860_1 (.in(n13860_0), .out(n13860_1));
wire n13861; //CHANY 4 (6,1) #37
wire n13861_0;
wire n13861_1;
buffer_wire buffer_13861_1 (.in(n13861_0), .out(n13861_1));
wire n13862; //CHANY 1 (6,1) #38
wire n13862_0;
wire n13863; //CHANY 1 (6,1) #39
wire n13863_0;
wire n13864; //CHANY 2 (6,1) #40
wire n13864_0;
wire n13865; //CHANY 2 (6,1) #41
wire n13865_0;
wire n13866; //CHANY 3 (6,1) #42
wire n13866_0;
wire n13867; //CHANY 3 (6,1) #43
wire n13867_0;
wire n13868; //CHANY 4 (6,1) #44
wire n13868_0;
wire n13868_1;
buffer_wire buffer_13868_1 (.in(n13868_0), .out(n13868_1));
wire n13869; //CHANY 4 (6,1) #45
wire n13869_0;
wire n13869_1;
buffer_wire buffer_13869_1 (.in(n13869_0), .out(n13869_1));
wire n13870; //CHANY 1 (6,1) #46
wire n13870_0;
wire n13871; //CHANY 1 (6,1) #47
wire n13871_0;
wire n13872; //CHANY 2 (6,1) #48
wire n13872_0;
wire n13873; //CHANY 2 (6,1) #49
wire n13873_0;
wire n13874; //CHANY 3 (6,1) #50
wire n13874_0;
wire n13875; //CHANY 3 (6,1) #51
wire n13875_0;
wire n13876; //CHANY 4 (6,1) #52
wire n13876_0;
wire n13876_1;
buffer_wire buffer_13876_1 (.in(n13876_0), .out(n13876_1));
wire n13877; //CHANY 4 (6,1) #53
wire n13877_0;
wire n13877_1;
buffer_wire buffer_13877_1 (.in(n13877_0), .out(n13877_1));
wire n13878; //CHANY 1 (6,1) #54
wire n13878_0;
wire n13879; //CHANY 1 (6,1) #55
wire n13879_0;
wire n13880; //CHANY 2 (6,1) #56
wire n13880_0;
wire n13881; //CHANY 2 (6,1) #57
wire n13881_0;
wire n13882; //CHANY 3 (6,1) #58
wire n13882_0;
wire n13883; //CHANY 3 (6,1) #59
wire n13883_0;
wire n13884; //CHANY 4 (6,1) #60
wire n13884_0;
wire n13884_1;
buffer_wire buffer_13884_1 (.in(n13884_0), .out(n13884_1));
wire n13885; //CHANY 4 (6,1) #61
wire n13885_0;
wire n13885_1;
buffer_wire buffer_13885_1 (.in(n13885_0), .out(n13885_1));
wire n13886; //CHANY 1 (6,1) #62
wire n13886_0;
wire n13887; //CHANY 1 (6,1) #63
wire n13887_0;
wire n13888; //CHANY 2 (6,1) #64
wire n13888_0;
wire n13889; //CHANY 2 (6,1) #65
wire n13889_0;
wire n13890; //CHANY 3 (6,1) #66
wire n13890_0;
wire n13891; //CHANY 3 (6,1) #67
wire n13891_0;
wire n13892; //CHANY 4 (6,1) #68
wire n13892_0;
wire n13892_1;
buffer_wire buffer_13892_1 (.in(n13892_0), .out(n13892_1));
wire n13893; //CHANY 4 (6,1) #69
wire n13893_0;
wire n13893_1;
buffer_wire buffer_13893_1 (.in(n13893_0), .out(n13893_1));
wire n13894; //CHANY 1 (6,1) #70
wire n13894_0;
wire n13895; //CHANY 1 (6,1) #71
wire n13895_0;
wire n13896; //CHANY 2 (6,1) #72
wire n13896_0;
wire n13897; //CHANY 2 (6,1) #73
wire n13897_0;
wire n13898; //CHANY 3 (6,1) #74
wire n13898_0;
wire n13899; //CHANY 3 (6,1) #75
wire n13899_0;
wire n13900; //CHANY 4 (6,1) #76
wire n13900_0;
wire n13900_1;
buffer_wire buffer_13900_1 (.in(n13900_0), .out(n13900_1));
wire n13901; //CHANY 4 (6,1) #77
wire n13901_0;
wire n13901_1;
buffer_wire buffer_13901_1 (.in(n13901_0), .out(n13901_1));
wire n13902; //CHANY 1 (6,1) #78
wire n13902_0;
wire n13903; //CHANY 1 (6,1) #79
wire n13903_0;
wire n13904; //CHANY 2 (6,1) #80
wire n13904_0;
wire n13905; //CHANY 2 (6,1) #81
wire n13905_0;
wire n13906; //CHANY 3 (6,1) #82
wire n13906_0;
wire n13907; //CHANY 3 (6,1) #83
wire n13907_0;
wire n13908; //CHANY 4 (6,1) #84
wire n13908_0;
wire n13908_1;
buffer_wire buffer_13908_1 (.in(n13908_0), .out(n13908_1));
wire n13909; //CHANY 4 (6,1) #85
wire n13909_0;
wire n13909_1;
buffer_wire buffer_13909_1 (.in(n13909_0), .out(n13909_1));
wire n13910; //CHANY 5 (6,1) #86
wire n13910_0;
wire n13910_1;
buffer_wire buffer_13910_1 (.in(n13910_0), .out(n13910_1));
wire n13911; //CHANY 5 (6,1) #87
wire n13911_0;
wire n13911_1;
buffer_wire buffer_13911_1 (.in(n13911_0), .out(n13911_1));
wire n13912; //CHANY 6 (6,1) #88
wire n13912_0;
wire n13912_1;
buffer_wire buffer_13912_1 (.in(n13912_0), .out(n13912_1));
wire n13913; //CHANY 6 (6,1) #89
wire n13913_0;
wire n13913_1;
buffer_wire buffer_13913_1 (.in(n13913_0), .out(n13913_1));
wire n13914; //CHANY 7 (6,1) #90
wire n13914_0;
wire n13914_1;
wire n13914_2;
buffer_wire buffer_13914_2 (.in(n13914_1), .out(n13914_2));
buffer_wire buffer_13914_1 (.in(n13914_0), .out(n13914_1));
wire n13915; //CHANY 7 (6,1) #91
wire n13915_0;
wire n13915_1;
wire n13915_2;
buffer_wire buffer_13915_2 (.in(n13915_1), .out(n13915_2));
buffer_wire buffer_13915_1 (.in(n13915_0), .out(n13915_1));
wire n13916; //CHANY 4 (6,2) #6
wire n13916_0;
wire n13916_1;
buffer_wire buffer_13916_1 (.in(n13916_0), .out(n13916_1));
wire n13917; //CHANY 4 (6,2) #7
wire n13917_0;
wire n13917_1;
buffer_wire buffer_13917_1 (.in(n13917_0), .out(n13917_1));
wire n13918; //CHANY 4 (6,2) #14
wire n13918_0;
wire n13918_1;
buffer_wire buffer_13918_1 (.in(n13918_0), .out(n13918_1));
wire n13919; //CHANY 4 (6,2) #15
wire n13919_0;
wire n13919_1;
buffer_wire buffer_13919_1 (.in(n13919_0), .out(n13919_1));
wire n13920; //CHANY 4 (6,2) #22
wire n13920_0;
wire n13920_1;
buffer_wire buffer_13920_1 (.in(n13920_0), .out(n13920_1));
wire n13921; //CHANY 4 (6,2) #23
wire n13921_0;
wire n13921_1;
buffer_wire buffer_13921_1 (.in(n13921_0), .out(n13921_1));
wire n13922; //CHANY 4 (6,2) #30
wire n13922_0;
wire n13922_1;
buffer_wire buffer_13922_1 (.in(n13922_0), .out(n13922_1));
wire n13923; //CHANY 4 (6,2) #31
wire n13923_0;
wire n13923_1;
buffer_wire buffer_13923_1 (.in(n13923_0), .out(n13923_1));
wire n13924; //CHANY 4 (6,2) #38
wire n13924_0;
wire n13924_1;
buffer_wire buffer_13924_1 (.in(n13924_0), .out(n13924_1));
wire n13925; //CHANY 4 (6,2) #39
wire n13925_0;
wire n13925_1;
buffer_wire buffer_13925_1 (.in(n13925_0), .out(n13925_1));
wire n13926; //CHANY 4 (6,2) #46
wire n13926_0;
wire n13926_1;
buffer_wire buffer_13926_1 (.in(n13926_0), .out(n13926_1));
wire n13927; //CHANY 4 (6,2) #47
wire n13927_0;
wire n13927_1;
buffer_wire buffer_13927_1 (.in(n13927_0), .out(n13927_1));
wire n13928; //CHANY 4 (6,2) #54
wire n13928_0;
wire n13928_1;
buffer_wire buffer_13928_1 (.in(n13928_0), .out(n13928_1));
wire n13929; //CHANY 4 (6,2) #55
wire n13929_0;
wire n13929_1;
buffer_wire buffer_13929_1 (.in(n13929_0), .out(n13929_1));
wire n13930; //CHANY 4 (6,2) #62
wire n13930_0;
wire n13930_1;
buffer_wire buffer_13930_1 (.in(n13930_0), .out(n13930_1));
wire n13931; //CHANY 4 (6,2) #63
wire n13931_0;
wire n13931_1;
buffer_wire buffer_13931_1 (.in(n13931_0), .out(n13931_1));
wire n13932; //CHANY 4 (6,2) #70
wire n13932_0;
wire n13932_1;
buffer_wire buffer_13932_1 (.in(n13932_0), .out(n13932_1));
wire n13933; //CHANY 4 (6,2) #71
wire n13933_0;
wire n13933_1;
buffer_wire buffer_13933_1 (.in(n13933_0), .out(n13933_1));
wire n13934; //CHANY 4 (6,2) #78
wire n13934_0;
wire n13934_1;
buffer_wire buffer_13934_1 (.in(n13934_0), .out(n13934_1));
wire n13935; //CHANY 4 (6,2) #79
wire n13935_0;
wire n13935_1;
buffer_wire buffer_13935_1 (.in(n13935_0), .out(n13935_1));
wire n13936; //CHANY 4 (6,3) #0
wire n13936_0;
wire n13936_1;
buffer_wire buffer_13936_1 (.in(n13936_0), .out(n13936_1));
wire n13937; //CHANY 4 (6,3) #1
wire n13937_0;
wire n13937_1;
buffer_wire buffer_13937_1 (.in(n13937_0), .out(n13937_1));
wire n13938; //CHANY 4 (6,3) #8
wire n13938_0;
wire n13938_1;
buffer_wire buffer_13938_1 (.in(n13938_0), .out(n13938_1));
wire n13939; //CHANY 4 (6,3) #9
wire n13939_0;
wire n13939_1;
buffer_wire buffer_13939_1 (.in(n13939_0), .out(n13939_1));
wire n13940; //CHANY 4 (6,3) #16
wire n13940_0;
wire n13940_1;
buffer_wire buffer_13940_1 (.in(n13940_0), .out(n13940_1));
wire n13941; //CHANY 4 (6,3) #17
wire n13941_0;
wire n13941_1;
buffer_wire buffer_13941_1 (.in(n13941_0), .out(n13941_1));
wire n13942; //CHANY 4 (6,3) #24
wire n13942_0;
wire n13942_1;
buffer_wire buffer_13942_1 (.in(n13942_0), .out(n13942_1));
wire n13943; //CHANY 4 (6,3) #25
wire n13943_0;
wire n13943_1;
buffer_wire buffer_13943_1 (.in(n13943_0), .out(n13943_1));
wire n13944; //CHANY 4 (6,3) #32
wire n13944_0;
wire n13944_1;
buffer_wire buffer_13944_1 (.in(n13944_0), .out(n13944_1));
wire n13945; //CHANY 4 (6,3) #33
wire n13945_0;
wire n13945_1;
buffer_wire buffer_13945_1 (.in(n13945_0), .out(n13945_1));
wire n13946; //CHANY 4 (6,3) #40
wire n13946_0;
wire n13946_1;
buffer_wire buffer_13946_1 (.in(n13946_0), .out(n13946_1));
wire n13947; //CHANY 4 (6,3) #41
wire n13947_0;
wire n13947_1;
buffer_wire buffer_13947_1 (.in(n13947_0), .out(n13947_1));
wire n13948; //CHANY 4 (6,3) #48
wire n13948_0;
wire n13948_1;
buffer_wire buffer_13948_1 (.in(n13948_0), .out(n13948_1));
wire n13949; //CHANY 4 (6,3) #49
wire n13949_0;
wire n13949_1;
buffer_wire buffer_13949_1 (.in(n13949_0), .out(n13949_1));
wire n13950; //CHANY 4 (6,3) #56
wire n13950_0;
wire n13950_1;
buffer_wire buffer_13950_1 (.in(n13950_0), .out(n13950_1));
wire n13951; //CHANY 4 (6,3) #57
wire n13951_0;
wire n13951_1;
buffer_wire buffer_13951_1 (.in(n13951_0), .out(n13951_1));
wire n13952; //CHANY 4 (6,3) #64
wire n13952_0;
wire n13952_1;
buffer_wire buffer_13952_1 (.in(n13952_0), .out(n13952_1));
wire n13953; //CHANY 4 (6,3) #65
wire n13953_0;
wire n13953_1;
buffer_wire buffer_13953_1 (.in(n13953_0), .out(n13953_1));
wire n13954; //CHANY 4 (6,3) #72
wire n13954_0;
wire n13954_1;
buffer_wire buffer_13954_1 (.in(n13954_0), .out(n13954_1));
wire n13955; //CHANY 4 (6,3) #73
wire n13955_0;
wire n13955_1;
buffer_wire buffer_13955_1 (.in(n13955_0), .out(n13955_1));
wire n13956; //CHANY 7 (6,3) #80
wire n13956_0;
wire n13956_1;
wire n13956_2;
buffer_wire buffer_13956_2 (.in(n13956_1), .out(n13956_2));
buffer_wire buffer_13956_1 (.in(n13956_0), .out(n13956_1));
wire n13957; //CHANY 7 (6,3) #81
wire n13957_0;
wire n13957_1;
wire n13957_2;
buffer_wire buffer_13957_2 (.in(n13957_1), .out(n13957_2));
buffer_wire buffer_13957_1 (.in(n13957_0), .out(n13957_1));
wire n13958; //CHANY 4 (6,4) #2
wire n13958_0;
wire n13958_1;
buffer_wire buffer_13958_1 (.in(n13958_0), .out(n13958_1));
wire n13959; //CHANY 4 (6,4) #3
wire n13959_0;
wire n13959_1;
buffer_wire buffer_13959_1 (.in(n13959_0), .out(n13959_1));
wire n13960; //CHANY 4 (6,4) #10
wire n13960_0;
wire n13960_1;
buffer_wire buffer_13960_1 (.in(n13960_0), .out(n13960_1));
wire n13961; //CHANY 4 (6,4) #11
wire n13961_0;
wire n13961_1;
buffer_wire buffer_13961_1 (.in(n13961_0), .out(n13961_1));
wire n13962; //CHANY 4 (6,4) #18
wire n13962_0;
wire n13962_1;
buffer_wire buffer_13962_1 (.in(n13962_0), .out(n13962_1));
wire n13963; //CHANY 4 (6,4) #19
wire n13963_0;
wire n13963_1;
buffer_wire buffer_13963_1 (.in(n13963_0), .out(n13963_1));
wire n13964; //CHANY 4 (6,4) #26
wire n13964_0;
wire n13964_1;
buffer_wire buffer_13964_1 (.in(n13964_0), .out(n13964_1));
wire n13965; //CHANY 4 (6,4) #27
wire n13965_0;
wire n13965_1;
buffer_wire buffer_13965_1 (.in(n13965_0), .out(n13965_1));
wire n13966; //CHANY 4 (6,4) #34
wire n13966_0;
wire n13966_1;
buffer_wire buffer_13966_1 (.in(n13966_0), .out(n13966_1));
wire n13967; //CHANY 4 (6,4) #35
wire n13967_0;
wire n13967_1;
buffer_wire buffer_13967_1 (.in(n13967_0), .out(n13967_1));
wire n13968; //CHANY 4 (6,4) #42
wire n13968_0;
wire n13968_1;
buffer_wire buffer_13968_1 (.in(n13968_0), .out(n13968_1));
wire n13969; //CHANY 4 (6,4) #43
wire n13969_0;
wire n13969_1;
buffer_wire buffer_13969_1 (.in(n13969_0), .out(n13969_1));
wire n13970; //CHANY 4 (6,4) #50
wire n13970_0;
wire n13970_1;
buffer_wire buffer_13970_1 (.in(n13970_0), .out(n13970_1));
wire n13971; //CHANY 4 (6,4) #51
wire n13971_0;
wire n13971_1;
buffer_wire buffer_13971_1 (.in(n13971_0), .out(n13971_1));
wire n13972; //CHANY 4 (6,4) #58
wire n13972_0;
wire n13972_1;
buffer_wire buffer_13972_1 (.in(n13972_0), .out(n13972_1));
wire n13973; //CHANY 4 (6,4) #59
wire n13973_0;
wire n13973_1;
buffer_wire buffer_13973_1 (.in(n13973_0), .out(n13973_1));
wire n13974; //CHANY 4 (6,4) #66
wire n13974_0;
wire n13974_1;
buffer_wire buffer_13974_1 (.in(n13974_0), .out(n13974_1));
wire n13975; //CHANY 4 (6,4) #67
wire n13975_0;
wire n13975_1;
buffer_wire buffer_13975_1 (.in(n13975_0), .out(n13975_1));
wire n13976; //CHANY 4 (6,4) #74
wire n13976_0;
wire n13976_1;
buffer_wire buffer_13976_1 (.in(n13976_0), .out(n13976_1));
wire n13977; //CHANY 4 (6,4) #75
wire n13977_0;
wire n13977_1;
buffer_wire buffer_13977_1 (.in(n13977_0), .out(n13977_1));
wire n13978; //CHANY 6 (6,4) #82
wire n13978_0;
wire n13978_1;
buffer_wire buffer_13978_1 (.in(n13978_0), .out(n13978_1));
wire n13979; //CHANY 6 (6,4) #83
wire n13979_0;
wire n13979_1;
buffer_wire buffer_13979_1 (.in(n13979_0), .out(n13979_1));
wire n13980; //CHANY 4 (6,5) #4
wire n13980_0;
wire n13980_1;
buffer_wire buffer_13980_1 (.in(n13980_0), .out(n13980_1));
wire n13981; //CHANY 4 (6,5) #5
wire n13981_0;
wire n13981_1;
buffer_wire buffer_13981_1 (.in(n13981_0), .out(n13981_1));
wire n13982; //CHANY 4 (6,5) #12
wire n13982_0;
wire n13982_1;
buffer_wire buffer_13982_1 (.in(n13982_0), .out(n13982_1));
wire n13983; //CHANY 4 (6,5) #13
wire n13983_0;
wire n13983_1;
buffer_wire buffer_13983_1 (.in(n13983_0), .out(n13983_1));
wire n13984; //CHANY 4 (6,5) #20
wire n13984_0;
wire n13984_1;
buffer_wire buffer_13984_1 (.in(n13984_0), .out(n13984_1));
wire n13985; //CHANY 4 (6,5) #21
wire n13985_0;
wire n13985_1;
buffer_wire buffer_13985_1 (.in(n13985_0), .out(n13985_1));
wire n13986; //CHANY 4 (6,5) #28
wire n13986_0;
wire n13986_1;
buffer_wire buffer_13986_1 (.in(n13986_0), .out(n13986_1));
wire n13987; //CHANY 4 (6,5) #29
wire n13987_0;
wire n13987_1;
buffer_wire buffer_13987_1 (.in(n13987_0), .out(n13987_1));
wire n13988; //CHANY 4 (6,5) #36
wire n13988_0;
wire n13988_1;
buffer_wire buffer_13988_1 (.in(n13988_0), .out(n13988_1));
wire n13989; //CHANY 4 (6,5) #37
wire n13989_0;
wire n13989_1;
buffer_wire buffer_13989_1 (.in(n13989_0), .out(n13989_1));
wire n13990; //CHANY 4 (6,5) #44
wire n13990_0;
wire n13990_1;
buffer_wire buffer_13990_1 (.in(n13990_0), .out(n13990_1));
wire n13991; //CHANY 4 (6,5) #45
wire n13991_0;
wire n13991_1;
buffer_wire buffer_13991_1 (.in(n13991_0), .out(n13991_1));
wire n13992; //CHANY 4 (6,5) #52
wire n13992_0;
wire n13992_1;
buffer_wire buffer_13992_1 (.in(n13992_0), .out(n13992_1));
wire n13993; //CHANY 4 (6,5) #53
wire n13993_0;
wire n13993_1;
buffer_wire buffer_13993_1 (.in(n13993_0), .out(n13993_1));
wire n13994; //CHANY 4 (6,5) #60
wire n13994_0;
wire n13994_1;
buffer_wire buffer_13994_1 (.in(n13994_0), .out(n13994_1));
wire n13995; //CHANY 4 (6,5) #61
wire n13995_0;
wire n13995_1;
buffer_wire buffer_13995_1 (.in(n13995_0), .out(n13995_1));
wire n13996; //CHANY 4 (6,5) #68
wire n13996_0;
wire n13996_1;
buffer_wire buffer_13996_1 (.in(n13996_0), .out(n13996_1));
wire n13997; //CHANY 4 (6,5) #69
wire n13997_0;
wire n13997_1;
buffer_wire buffer_13997_1 (.in(n13997_0), .out(n13997_1));
wire n13998; //CHANY 4 (6,5) #76
wire n13998_0;
wire n13998_1;
buffer_wire buffer_13998_1 (.in(n13998_0), .out(n13998_1));
wire n13999; //CHANY 4 (6,5) #77
wire n13999_0;
wire n13999_1;
buffer_wire buffer_13999_1 (.in(n13999_0), .out(n13999_1));
wire n14000; //CHANY 5 (6,5) #84
wire n14000_0;
wire n14000_1;
buffer_wire buffer_14000_1 (.in(n14000_0), .out(n14000_1));
wire n14001; //CHANY 5 (6,5) #85
wire n14001_0;
wire n14001_1;
buffer_wire buffer_14001_1 (.in(n14001_0), .out(n14001_1));
wire n14002; //CHANY 4 (6,6) #6
wire n14002_0;
wire n14002_1;
buffer_wire buffer_14002_1 (.in(n14002_0), .out(n14002_1));
wire n14003; //CHANY 4 (6,6) #7
wire n14003_0;
wire n14003_1;
buffer_wire buffer_14003_1 (.in(n14003_0), .out(n14003_1));
wire n14004; //CHANY 4 (6,6) #14
wire n14004_0;
wire n14004_1;
buffer_wire buffer_14004_1 (.in(n14004_0), .out(n14004_1));
wire n14005; //CHANY 4 (6,6) #15
wire n14005_0;
wire n14005_1;
buffer_wire buffer_14005_1 (.in(n14005_0), .out(n14005_1));
wire n14006; //CHANY 4 (6,6) #22
wire n14006_0;
wire n14006_1;
buffer_wire buffer_14006_1 (.in(n14006_0), .out(n14006_1));
wire n14007; //CHANY 4 (6,6) #23
wire n14007_0;
wire n14007_1;
buffer_wire buffer_14007_1 (.in(n14007_0), .out(n14007_1));
wire n14008; //CHANY 4 (6,6) #30
wire n14008_0;
wire n14008_1;
buffer_wire buffer_14008_1 (.in(n14008_0), .out(n14008_1));
wire n14009; //CHANY 4 (6,6) #31
wire n14009_0;
wire n14009_1;
buffer_wire buffer_14009_1 (.in(n14009_0), .out(n14009_1));
wire n14010; //CHANY 4 (6,6) #38
wire n14010_0;
wire n14010_1;
buffer_wire buffer_14010_1 (.in(n14010_0), .out(n14010_1));
wire n14011; //CHANY 4 (6,6) #39
wire n14011_0;
wire n14011_1;
buffer_wire buffer_14011_1 (.in(n14011_0), .out(n14011_1));
wire n14012; //CHANY 4 (6,6) #46
wire n14012_0;
wire n14012_1;
buffer_wire buffer_14012_1 (.in(n14012_0), .out(n14012_1));
wire n14013; //CHANY 4 (6,6) #47
wire n14013_0;
wire n14013_1;
buffer_wire buffer_14013_1 (.in(n14013_0), .out(n14013_1));
wire n14014; //CHANY 4 (6,6) #54
wire n14014_0;
wire n14014_1;
buffer_wire buffer_14014_1 (.in(n14014_0), .out(n14014_1));
wire n14015; //CHANY 4 (6,6) #55
wire n14015_0;
wire n14015_1;
buffer_wire buffer_14015_1 (.in(n14015_0), .out(n14015_1));
wire n14016; //CHANY 4 (6,6) #62
wire n14016_0;
wire n14016_1;
buffer_wire buffer_14016_1 (.in(n14016_0), .out(n14016_1));
wire n14017; //CHANY 4 (6,6) #63
wire n14017_0;
wire n14017_1;
buffer_wire buffer_14017_1 (.in(n14017_0), .out(n14017_1));
wire n14018; //CHANY 4 (6,6) #70
wire n14018_0;
wire n14018_1;
buffer_wire buffer_14018_1 (.in(n14018_0), .out(n14018_1));
wire n14019; //CHANY 4 (6,6) #71
wire n14019_0;
wire n14019_1;
buffer_wire buffer_14019_1 (.in(n14019_0), .out(n14019_1));
wire n14020; //CHANY 4 (6,6) #78
wire n14020_0;
wire n14020_1;
buffer_wire buffer_14020_1 (.in(n14020_0), .out(n14020_1));
wire n14021; //CHANY 4 (6,6) #79
wire n14021_0;
wire n14021_1;
buffer_wire buffer_14021_1 (.in(n14021_0), .out(n14021_1));
wire n14022; //CHANY 4 (6,6) #86
wire n14022_0;
wire n14022_1;
buffer_wire buffer_14022_1 (.in(n14022_0), .out(n14022_1));
wire n14023; //CHANY 4 (6,6) #87
wire n14023_0;
wire n14023_1;
buffer_wire buffer_14023_1 (.in(n14023_0), .out(n14023_1));
wire n14024; //CHANY 3 (6,7) #0
wire n14024_0;
wire n14025; //CHANY 3 (6,7) #1
wire n14025_0;
wire n14026; //CHANY 3 (6,7) #8
wire n14026_0;
wire n14027; //CHANY 3 (6,7) #9
wire n14027_0;
wire n14028; //CHANY 3 (6,7) #16
wire n14028_0;
wire n14029; //CHANY 3 (6,7) #17
wire n14029_0;
wire n14030; //CHANY 3 (6,7) #24
wire n14030_0;
wire n14031; //CHANY 3 (6,7) #25
wire n14031_0;
wire n14032; //CHANY 3 (6,7) #32
wire n14032_0;
wire n14033; //CHANY 3 (6,7) #33
wire n14033_0;
wire n14034; //CHANY 3 (6,7) #40
wire n14034_0;
wire n14035; //CHANY 3 (6,7) #41
wire n14035_0;
wire n14036; //CHANY 3 (6,7) #48
wire n14036_0;
wire n14037; //CHANY 3 (6,7) #49
wire n14037_0;
wire n14038; //CHANY 3 (6,7) #56
wire n14038_0;
wire n14039; //CHANY 3 (6,7) #57
wire n14039_0;
wire n14040; //CHANY 3 (6,7) #64
wire n14040_0;
wire n14041; //CHANY 3 (6,7) #65
wire n14041_0;
wire n14042; //CHANY 3 (6,7) #72
wire n14042_0;
wire n14043; //CHANY 3 (6,7) #73
wire n14043_0;
wire n14044; //CHANY 3 (6,7) #88
wire n14044_0;
wire n14045; //CHANY 3 (6,7) #89
wire n14045_0;
wire n14046; //CHANY 2 (6,8) #2
wire n14046_0;
wire n14047; //CHANY 2 (6,8) #3
wire n14047_0;
wire n14048; //CHANY 2 (6,8) #10
wire n14048_0;
wire n14049; //CHANY 2 (6,8) #11
wire n14049_0;
wire n14050; //CHANY 2 (6,8) #18
wire n14050_0;
wire n14051; //CHANY 2 (6,8) #19
wire n14051_0;
wire n14052; //CHANY 2 (6,8) #26
wire n14052_0;
wire n14053; //CHANY 2 (6,8) #27
wire n14053_0;
wire n14054; //CHANY 2 (6,8) #34
wire n14054_0;
wire n14055; //CHANY 2 (6,8) #35
wire n14055_0;
wire n14056; //CHANY 2 (6,8) #42
wire n14056_0;
wire n14057; //CHANY 2 (6,8) #43
wire n14057_0;
wire n14058; //CHANY 2 (6,8) #50
wire n14058_0;
wire n14059; //CHANY 2 (6,8) #51
wire n14059_0;
wire n14060; //CHANY 2 (6,8) #58
wire n14060_0;
wire n14061; //CHANY 2 (6,8) #59
wire n14061_0;
wire n14062; //CHANY 2 (6,8) #66
wire n14062_0;
wire n14063; //CHANY 2 (6,8) #67
wire n14063_0;
wire n14064; //CHANY 2 (6,8) #74
wire n14064_0;
wire n14065; //CHANY 2 (6,8) #75
wire n14065_0;
wire n14066; //CHANY 2 (6,8) #90
wire n14066_0;
wire n14067; //CHANY 2 (6,8) #91
wire n14067_0;
wire n14068; //CHANY 1 (6,9) #4
wire n14068_0;
wire n14069; //CHANY 1 (6,9) #5
wire n14069_0;
wire n14070; //CHANY 1 (6,9) #12
wire n14070_0;
wire n14071; //CHANY 1 (6,9) #13
wire n14071_0;
wire n14072; //CHANY 1 (6,9) #20
wire n14072_0;
wire n14073; //CHANY 1 (6,9) #21
wire n14073_0;
wire n14074; //CHANY 1 (6,9) #28
wire n14074_0;
wire n14075; //CHANY 1 (6,9) #29
wire n14075_0;
wire n14076; //CHANY 1 (6,9) #36
wire n14076_0;
wire n14077; //CHANY 1 (6,9) #37
wire n14077_0;
wire n14078; //CHANY 1 (6,9) #44
wire n14078_0;
wire n14079; //CHANY 1 (6,9) #45
wire n14079_0;
wire n14080; //CHANY 1 (6,9) #52
wire n14080_0;
wire n14081; //CHANY 1 (6,9) #53
wire n14081_0;
wire n14082; //CHANY 1 (6,9) #60
wire n14082_0;
wire n14083; //CHANY 1 (6,9) #61
wire n14083_0;
wire n14084; //CHANY 1 (6,9) #68
wire n14084_0;
wire n14085; //CHANY 1 (6,9) #69
wire n14085_0;
wire n14086; //CHANY 1 (6,9) #76
wire n14086_0;
wire n14087; //CHANY 1 (6,9) #77
wire n14087_0;
wire n14088; //CHANY 1 (7,1) #0
wire n14088_0;
wire n14089; //CHANY 1 (7,1) #1
wire n14089_0;
wire n14090; //CHANY 2 (7,1) #2
wire n14090_0;
wire n14091; //CHANY 2 (7,1) #3
wire n14091_0;
wire n14092; //CHANY 3 (7,1) #4
wire n14092_0;
wire n14093; //CHANY 3 (7,1) #5
wire n14093_0;
wire n14094; //CHANY 4 (7,1) #6
wire n14094_0;
wire n14094_1;
buffer_wire buffer_14094_1 (.in(n14094_0), .out(n14094_1));
wire n14095; //CHANY 4 (7,1) #7
wire n14095_0;
wire n14095_1;
buffer_wire buffer_14095_1 (.in(n14095_0), .out(n14095_1));
wire n14096; //CHANY 1 (7,1) #8
wire n14096_0;
wire n14097; //CHANY 1 (7,1) #9
wire n14097_0;
wire n14098; //CHANY 2 (7,1) #10
wire n14098_0;
wire n14099; //CHANY 2 (7,1) #11
wire n14099_0;
wire n14100; //CHANY 3 (7,1) #12
wire n14100_0;
wire n14101; //CHANY 3 (7,1) #13
wire n14101_0;
wire n14102; //CHANY 4 (7,1) #14
wire n14102_0;
wire n14102_1;
buffer_wire buffer_14102_1 (.in(n14102_0), .out(n14102_1));
wire n14103; //CHANY 4 (7,1) #15
wire n14103_0;
wire n14103_1;
buffer_wire buffer_14103_1 (.in(n14103_0), .out(n14103_1));
wire n14104; //CHANY 1 (7,1) #16
wire n14104_0;
wire n14105; //CHANY 1 (7,1) #17
wire n14105_0;
wire n14106; //CHANY 2 (7,1) #18
wire n14106_0;
wire n14107; //CHANY 2 (7,1) #19
wire n14107_0;
wire n14108; //CHANY 3 (7,1) #20
wire n14108_0;
wire n14109; //CHANY 3 (7,1) #21
wire n14109_0;
wire n14110; //CHANY 4 (7,1) #22
wire n14110_0;
wire n14110_1;
buffer_wire buffer_14110_1 (.in(n14110_0), .out(n14110_1));
wire n14111; //CHANY 4 (7,1) #23
wire n14111_0;
wire n14111_1;
buffer_wire buffer_14111_1 (.in(n14111_0), .out(n14111_1));
wire n14112; //CHANY 1 (7,1) #24
wire n14112_0;
wire n14113; //CHANY 1 (7,1) #25
wire n14113_0;
wire n14114; //CHANY 2 (7,1) #26
wire n14114_0;
wire n14115; //CHANY 2 (7,1) #27
wire n14115_0;
wire n14116; //CHANY 3 (7,1) #28
wire n14116_0;
wire n14117; //CHANY 3 (7,1) #29
wire n14117_0;
wire n14118; //CHANY 4 (7,1) #30
wire n14118_0;
wire n14118_1;
buffer_wire buffer_14118_1 (.in(n14118_0), .out(n14118_1));
wire n14119; //CHANY 4 (7,1) #31
wire n14119_0;
wire n14119_1;
buffer_wire buffer_14119_1 (.in(n14119_0), .out(n14119_1));
wire n14120; //CHANY 1 (7,1) #32
wire n14120_0;
wire n14121; //CHANY 1 (7,1) #33
wire n14121_0;
wire n14122; //CHANY 2 (7,1) #34
wire n14122_0;
wire n14123; //CHANY 2 (7,1) #35
wire n14123_0;
wire n14124; //CHANY 3 (7,1) #36
wire n14124_0;
wire n14125; //CHANY 3 (7,1) #37
wire n14125_0;
wire n14126; //CHANY 4 (7,1) #38
wire n14126_0;
wire n14126_1;
buffer_wire buffer_14126_1 (.in(n14126_0), .out(n14126_1));
wire n14127; //CHANY 4 (7,1) #39
wire n14127_0;
wire n14127_1;
buffer_wire buffer_14127_1 (.in(n14127_0), .out(n14127_1));
wire n14128; //CHANY 1 (7,1) #40
wire n14128_0;
wire n14129; //CHANY 1 (7,1) #41
wire n14129_0;
wire n14130; //CHANY 2 (7,1) #42
wire n14130_0;
wire n14131; //CHANY 2 (7,1) #43
wire n14131_0;
wire n14132; //CHANY 3 (7,1) #44
wire n14132_0;
wire n14133; //CHANY 3 (7,1) #45
wire n14133_0;
wire n14134; //CHANY 4 (7,1) #46
wire n14134_0;
wire n14134_1;
buffer_wire buffer_14134_1 (.in(n14134_0), .out(n14134_1));
wire n14135; //CHANY 4 (7,1) #47
wire n14135_0;
wire n14135_1;
buffer_wire buffer_14135_1 (.in(n14135_0), .out(n14135_1));
wire n14136; //CHANY 1 (7,1) #48
wire n14136_0;
wire n14137; //CHANY 1 (7,1) #49
wire n14137_0;
wire n14138; //CHANY 2 (7,1) #50
wire n14138_0;
wire n14139; //CHANY 2 (7,1) #51
wire n14139_0;
wire n14140; //CHANY 3 (7,1) #52
wire n14140_0;
wire n14141; //CHANY 3 (7,1) #53
wire n14141_0;
wire n14142; //CHANY 4 (7,1) #54
wire n14142_0;
wire n14142_1;
buffer_wire buffer_14142_1 (.in(n14142_0), .out(n14142_1));
wire n14143; //CHANY 4 (7,1) #55
wire n14143_0;
wire n14143_1;
buffer_wire buffer_14143_1 (.in(n14143_0), .out(n14143_1));
wire n14144; //CHANY 1 (7,1) #56
wire n14144_0;
wire n14145; //CHANY 1 (7,1) #57
wire n14145_0;
wire n14146; //CHANY 2 (7,1) #58
wire n14146_0;
wire n14147; //CHANY 2 (7,1) #59
wire n14147_0;
wire n14148; //CHANY 3 (7,1) #60
wire n14148_0;
wire n14149; //CHANY 3 (7,1) #61
wire n14149_0;
wire n14150; //CHANY 4 (7,1) #62
wire n14150_0;
wire n14150_1;
buffer_wire buffer_14150_1 (.in(n14150_0), .out(n14150_1));
wire n14151; //CHANY 4 (7,1) #63
wire n14151_0;
wire n14151_1;
buffer_wire buffer_14151_1 (.in(n14151_0), .out(n14151_1));
wire n14152; //CHANY 1 (7,1) #64
wire n14152_0;
wire n14153; //CHANY 1 (7,1) #65
wire n14153_0;
wire n14154; //CHANY 2 (7,1) #66
wire n14154_0;
wire n14155; //CHANY 2 (7,1) #67
wire n14155_0;
wire n14156; //CHANY 3 (7,1) #68
wire n14156_0;
wire n14157; //CHANY 3 (7,1) #69
wire n14157_0;
wire n14158; //CHANY 4 (7,1) #70
wire n14158_0;
wire n14158_1;
buffer_wire buffer_14158_1 (.in(n14158_0), .out(n14158_1));
wire n14159; //CHANY 4 (7,1) #71
wire n14159_0;
wire n14159_1;
buffer_wire buffer_14159_1 (.in(n14159_0), .out(n14159_1));
wire n14160; //CHANY 1 (7,1) #72
wire n14160_0;
wire n14161; //CHANY 1 (7,1) #73
wire n14161_0;
wire n14162; //CHANY 2 (7,1) #74
wire n14162_0;
wire n14163; //CHANY 2 (7,1) #75
wire n14163_0;
wire n14164; //CHANY 3 (7,1) #76
wire n14164_0;
wire n14165; //CHANY 3 (7,1) #77
wire n14165_0;
wire n14166; //CHANY 4 (7,1) #78
wire n14166_0;
wire n14166_1;
buffer_wire buffer_14166_1 (.in(n14166_0), .out(n14166_1));
wire n14167; //CHANY 4 (7,1) #79
wire n14167_0;
wire n14167_1;
buffer_wire buffer_14167_1 (.in(n14167_0), .out(n14167_1));
wire n14168; //CHANY 1 (7,1) #80
wire n14168_0;
wire n14169; //CHANY 1 (7,1) #81
wire n14169_0;
wire n14170; //CHANY 2 (7,1) #82
wire n14170_0;
wire n14171; //CHANY 2 (7,1) #83
wire n14171_0;
wire n14172; //CHANY 3 (7,1) #84
wire n14172_0;
wire n14173; //CHANY 3 (7,1) #85
wire n14173_0;
wire n14174; //CHANY 4 (7,1) #86
wire n14174_0;
wire n14174_1;
buffer_wire buffer_14174_1 (.in(n14174_0), .out(n14174_1));
wire n14175; //CHANY 4 (7,1) #87
wire n14175_0;
wire n14175_1;
buffer_wire buffer_14175_1 (.in(n14175_0), .out(n14175_1));
wire n14176; //CHANY 5 (7,1) #88
wire n14176_0;
wire n14176_1;
buffer_wire buffer_14176_1 (.in(n14176_0), .out(n14176_1));
wire n14177; //CHANY 5 (7,1) #89
wire n14177_0;
wire n14177_1;
buffer_wire buffer_14177_1 (.in(n14177_0), .out(n14177_1));
wire n14178; //CHANY 6 (7,1) #90
wire n14178_0;
wire n14178_1;
buffer_wire buffer_14178_1 (.in(n14178_0), .out(n14178_1));
wire n14179; //CHANY 6 (7,1) #91
wire n14179_0;
wire n14179_1;
buffer_wire buffer_14179_1 (.in(n14179_0), .out(n14179_1));
wire n14180; //CHANY 4 (7,2) #0
wire n14180_0;
wire n14180_1;
buffer_wire buffer_14180_1 (.in(n14180_0), .out(n14180_1));
wire n14181; //CHANY 4 (7,2) #1
wire n14181_0;
wire n14181_1;
buffer_wire buffer_14181_1 (.in(n14181_0), .out(n14181_1));
wire n14182; //CHANY 4 (7,2) #8
wire n14182_0;
wire n14182_1;
buffer_wire buffer_14182_1 (.in(n14182_0), .out(n14182_1));
wire n14183; //CHANY 4 (7,2) #9
wire n14183_0;
wire n14183_1;
buffer_wire buffer_14183_1 (.in(n14183_0), .out(n14183_1));
wire n14184; //CHANY 4 (7,2) #16
wire n14184_0;
wire n14184_1;
buffer_wire buffer_14184_1 (.in(n14184_0), .out(n14184_1));
wire n14185; //CHANY 4 (7,2) #17
wire n14185_0;
wire n14185_1;
buffer_wire buffer_14185_1 (.in(n14185_0), .out(n14185_1));
wire n14186; //CHANY 4 (7,2) #24
wire n14186_0;
wire n14186_1;
buffer_wire buffer_14186_1 (.in(n14186_0), .out(n14186_1));
wire n14187; //CHANY 4 (7,2) #25
wire n14187_0;
wire n14187_1;
buffer_wire buffer_14187_1 (.in(n14187_0), .out(n14187_1));
wire n14188; //CHANY 4 (7,2) #32
wire n14188_0;
wire n14188_1;
buffer_wire buffer_14188_1 (.in(n14188_0), .out(n14188_1));
wire n14189; //CHANY 4 (7,2) #33
wire n14189_0;
wire n14189_1;
buffer_wire buffer_14189_1 (.in(n14189_0), .out(n14189_1));
wire n14190; //CHANY 4 (7,2) #40
wire n14190_0;
wire n14190_1;
buffer_wire buffer_14190_1 (.in(n14190_0), .out(n14190_1));
wire n14191; //CHANY 4 (7,2) #41
wire n14191_0;
wire n14191_1;
buffer_wire buffer_14191_1 (.in(n14191_0), .out(n14191_1));
wire n14192; //CHANY 4 (7,2) #48
wire n14192_0;
wire n14192_1;
buffer_wire buffer_14192_1 (.in(n14192_0), .out(n14192_1));
wire n14193; //CHANY 4 (7,2) #49
wire n14193_0;
wire n14193_1;
buffer_wire buffer_14193_1 (.in(n14193_0), .out(n14193_1));
wire n14194; //CHANY 4 (7,2) #56
wire n14194_0;
wire n14194_1;
buffer_wire buffer_14194_1 (.in(n14194_0), .out(n14194_1));
wire n14195; //CHANY 4 (7,2) #57
wire n14195_0;
wire n14195_1;
buffer_wire buffer_14195_1 (.in(n14195_0), .out(n14195_1));
wire n14196; //CHANY 4 (7,2) #64
wire n14196_0;
wire n14196_1;
buffer_wire buffer_14196_1 (.in(n14196_0), .out(n14196_1));
wire n14197; //CHANY 4 (7,2) #65
wire n14197_0;
wire n14197_1;
buffer_wire buffer_14197_1 (.in(n14197_0), .out(n14197_1));
wire n14198; //CHANY 4 (7,2) #72
wire n14198_0;
wire n14198_1;
buffer_wire buffer_14198_1 (.in(n14198_0), .out(n14198_1));
wire n14199; //CHANY 4 (7,2) #73
wire n14199_0;
wire n14199_1;
buffer_wire buffer_14199_1 (.in(n14199_0), .out(n14199_1));
wire n14200; //CHANY 8 (7,2) #80
wire n14200_0;
wire n14200_1;
wire n14200_2;
buffer_wire buffer_14200_2 (.in(n14200_1), .out(n14200_2));
buffer_wire buffer_14200_1 (.in(n14200_0), .out(n14200_1));
wire n14201; //CHANY 8 (7,2) #81
wire n14201_0;
wire n14201_1;
wire n14201_2;
buffer_wire buffer_14201_2 (.in(n14201_1), .out(n14201_2));
buffer_wire buffer_14201_1 (.in(n14201_0), .out(n14201_1));
wire n14202; //CHANY 4 (7,3) #2
wire n14202_0;
wire n14202_1;
buffer_wire buffer_14202_1 (.in(n14202_0), .out(n14202_1));
wire n14203; //CHANY 4 (7,3) #3
wire n14203_0;
wire n14203_1;
buffer_wire buffer_14203_1 (.in(n14203_0), .out(n14203_1));
wire n14204; //CHANY 4 (7,3) #10
wire n14204_0;
wire n14204_1;
buffer_wire buffer_14204_1 (.in(n14204_0), .out(n14204_1));
wire n14205; //CHANY 4 (7,3) #11
wire n14205_0;
wire n14205_1;
buffer_wire buffer_14205_1 (.in(n14205_0), .out(n14205_1));
wire n14206; //CHANY 4 (7,3) #18
wire n14206_0;
wire n14206_1;
buffer_wire buffer_14206_1 (.in(n14206_0), .out(n14206_1));
wire n14207; //CHANY 4 (7,3) #19
wire n14207_0;
wire n14207_1;
buffer_wire buffer_14207_1 (.in(n14207_0), .out(n14207_1));
wire n14208; //CHANY 4 (7,3) #26
wire n14208_0;
wire n14208_1;
buffer_wire buffer_14208_1 (.in(n14208_0), .out(n14208_1));
wire n14209; //CHANY 4 (7,3) #27
wire n14209_0;
wire n14209_1;
buffer_wire buffer_14209_1 (.in(n14209_0), .out(n14209_1));
wire n14210; //CHANY 4 (7,3) #34
wire n14210_0;
wire n14210_1;
buffer_wire buffer_14210_1 (.in(n14210_0), .out(n14210_1));
wire n14211; //CHANY 4 (7,3) #35
wire n14211_0;
wire n14211_1;
buffer_wire buffer_14211_1 (.in(n14211_0), .out(n14211_1));
wire n14212; //CHANY 4 (7,3) #42
wire n14212_0;
wire n14212_1;
buffer_wire buffer_14212_1 (.in(n14212_0), .out(n14212_1));
wire n14213; //CHANY 4 (7,3) #43
wire n14213_0;
wire n14213_1;
buffer_wire buffer_14213_1 (.in(n14213_0), .out(n14213_1));
wire n14214; //CHANY 4 (7,3) #50
wire n14214_0;
wire n14214_1;
buffer_wire buffer_14214_1 (.in(n14214_0), .out(n14214_1));
wire n14215; //CHANY 4 (7,3) #51
wire n14215_0;
wire n14215_1;
buffer_wire buffer_14215_1 (.in(n14215_0), .out(n14215_1));
wire n14216; //CHANY 4 (7,3) #58
wire n14216_0;
wire n14216_1;
buffer_wire buffer_14216_1 (.in(n14216_0), .out(n14216_1));
wire n14217; //CHANY 4 (7,3) #59
wire n14217_0;
wire n14217_1;
buffer_wire buffer_14217_1 (.in(n14217_0), .out(n14217_1));
wire n14218; //CHANY 4 (7,3) #66
wire n14218_0;
wire n14218_1;
buffer_wire buffer_14218_1 (.in(n14218_0), .out(n14218_1));
wire n14219; //CHANY 4 (7,3) #67
wire n14219_0;
wire n14219_1;
buffer_wire buffer_14219_1 (.in(n14219_0), .out(n14219_1));
wire n14220; //CHANY 4 (7,3) #74
wire n14220_0;
wire n14220_1;
buffer_wire buffer_14220_1 (.in(n14220_0), .out(n14220_1));
wire n14221; //CHANY 4 (7,3) #75
wire n14221_0;
wire n14221_1;
buffer_wire buffer_14221_1 (.in(n14221_0), .out(n14221_1));
wire n14222; //CHANY 7 (7,3) #82
wire n14222_0;
wire n14222_1;
wire n14222_2;
buffer_wire buffer_14222_2 (.in(n14222_1), .out(n14222_2));
buffer_wire buffer_14222_1 (.in(n14222_0), .out(n14222_1));
wire n14223; //CHANY 7 (7,3) #83
wire n14223_0;
wire n14223_1;
wire n14223_2;
buffer_wire buffer_14223_2 (.in(n14223_1), .out(n14223_2));
buffer_wire buffer_14223_1 (.in(n14223_0), .out(n14223_1));
wire n14224; //CHANY 4 (7,4) #4
wire n14224_0;
wire n14224_1;
buffer_wire buffer_14224_1 (.in(n14224_0), .out(n14224_1));
wire n14225; //CHANY 4 (7,4) #5
wire n14225_0;
wire n14225_1;
buffer_wire buffer_14225_1 (.in(n14225_0), .out(n14225_1));
wire n14226; //CHANY 4 (7,4) #12
wire n14226_0;
wire n14226_1;
buffer_wire buffer_14226_1 (.in(n14226_0), .out(n14226_1));
wire n14227; //CHANY 4 (7,4) #13
wire n14227_0;
wire n14227_1;
buffer_wire buffer_14227_1 (.in(n14227_0), .out(n14227_1));
wire n14228; //CHANY 4 (7,4) #20
wire n14228_0;
wire n14228_1;
buffer_wire buffer_14228_1 (.in(n14228_0), .out(n14228_1));
wire n14229; //CHANY 4 (7,4) #21
wire n14229_0;
wire n14229_1;
buffer_wire buffer_14229_1 (.in(n14229_0), .out(n14229_1));
wire n14230; //CHANY 4 (7,4) #28
wire n14230_0;
wire n14230_1;
buffer_wire buffer_14230_1 (.in(n14230_0), .out(n14230_1));
wire n14231; //CHANY 4 (7,4) #29
wire n14231_0;
wire n14231_1;
buffer_wire buffer_14231_1 (.in(n14231_0), .out(n14231_1));
wire n14232; //CHANY 4 (7,4) #36
wire n14232_0;
wire n14232_1;
buffer_wire buffer_14232_1 (.in(n14232_0), .out(n14232_1));
wire n14233; //CHANY 4 (7,4) #37
wire n14233_0;
wire n14233_1;
buffer_wire buffer_14233_1 (.in(n14233_0), .out(n14233_1));
wire n14234; //CHANY 4 (7,4) #44
wire n14234_0;
wire n14234_1;
buffer_wire buffer_14234_1 (.in(n14234_0), .out(n14234_1));
wire n14235; //CHANY 4 (7,4) #45
wire n14235_0;
wire n14235_1;
buffer_wire buffer_14235_1 (.in(n14235_0), .out(n14235_1));
wire n14236; //CHANY 4 (7,4) #52
wire n14236_0;
wire n14236_1;
buffer_wire buffer_14236_1 (.in(n14236_0), .out(n14236_1));
wire n14237; //CHANY 4 (7,4) #53
wire n14237_0;
wire n14237_1;
buffer_wire buffer_14237_1 (.in(n14237_0), .out(n14237_1));
wire n14238; //CHANY 4 (7,4) #60
wire n14238_0;
wire n14238_1;
buffer_wire buffer_14238_1 (.in(n14238_0), .out(n14238_1));
wire n14239; //CHANY 4 (7,4) #61
wire n14239_0;
wire n14239_1;
buffer_wire buffer_14239_1 (.in(n14239_0), .out(n14239_1));
wire n14240; //CHANY 4 (7,4) #68
wire n14240_0;
wire n14240_1;
buffer_wire buffer_14240_1 (.in(n14240_0), .out(n14240_1));
wire n14241; //CHANY 4 (7,4) #69
wire n14241_0;
wire n14241_1;
buffer_wire buffer_14241_1 (.in(n14241_0), .out(n14241_1));
wire n14242; //CHANY 4 (7,4) #76
wire n14242_0;
wire n14242_1;
buffer_wire buffer_14242_1 (.in(n14242_0), .out(n14242_1));
wire n14243; //CHANY 4 (7,4) #77
wire n14243_0;
wire n14243_1;
buffer_wire buffer_14243_1 (.in(n14243_0), .out(n14243_1));
wire n14244; //CHANY 6 (7,4) #84
wire n14244_0;
wire n14244_1;
buffer_wire buffer_14244_1 (.in(n14244_0), .out(n14244_1));
wire n14245; //CHANY 6 (7,4) #85
wire n14245_0;
wire n14245_1;
buffer_wire buffer_14245_1 (.in(n14245_0), .out(n14245_1));
wire n14246; //CHANY 4 (7,5) #6
wire n14246_0;
wire n14246_1;
buffer_wire buffer_14246_1 (.in(n14246_0), .out(n14246_1));
wire n14247; //CHANY 4 (7,5) #7
wire n14247_0;
wire n14247_1;
buffer_wire buffer_14247_1 (.in(n14247_0), .out(n14247_1));
wire n14248; //CHANY 4 (7,5) #14
wire n14248_0;
wire n14248_1;
buffer_wire buffer_14248_1 (.in(n14248_0), .out(n14248_1));
wire n14249; //CHANY 4 (7,5) #15
wire n14249_0;
wire n14249_1;
buffer_wire buffer_14249_1 (.in(n14249_0), .out(n14249_1));
wire n14250; //CHANY 4 (7,5) #22
wire n14250_0;
wire n14250_1;
buffer_wire buffer_14250_1 (.in(n14250_0), .out(n14250_1));
wire n14251; //CHANY 4 (7,5) #23
wire n14251_0;
wire n14251_1;
buffer_wire buffer_14251_1 (.in(n14251_0), .out(n14251_1));
wire n14252; //CHANY 4 (7,5) #30
wire n14252_0;
wire n14252_1;
buffer_wire buffer_14252_1 (.in(n14252_0), .out(n14252_1));
wire n14253; //CHANY 4 (7,5) #31
wire n14253_0;
wire n14253_1;
buffer_wire buffer_14253_1 (.in(n14253_0), .out(n14253_1));
wire n14254; //CHANY 4 (7,5) #38
wire n14254_0;
wire n14254_1;
buffer_wire buffer_14254_1 (.in(n14254_0), .out(n14254_1));
wire n14255; //CHANY 4 (7,5) #39
wire n14255_0;
wire n14255_1;
buffer_wire buffer_14255_1 (.in(n14255_0), .out(n14255_1));
wire n14256; //CHANY 4 (7,5) #46
wire n14256_0;
wire n14256_1;
buffer_wire buffer_14256_1 (.in(n14256_0), .out(n14256_1));
wire n14257; //CHANY 4 (7,5) #47
wire n14257_0;
wire n14257_1;
buffer_wire buffer_14257_1 (.in(n14257_0), .out(n14257_1));
wire n14258; //CHANY 4 (7,5) #54
wire n14258_0;
wire n14258_1;
buffer_wire buffer_14258_1 (.in(n14258_0), .out(n14258_1));
wire n14259; //CHANY 4 (7,5) #55
wire n14259_0;
wire n14259_1;
buffer_wire buffer_14259_1 (.in(n14259_0), .out(n14259_1));
wire n14260; //CHANY 4 (7,5) #62
wire n14260_0;
wire n14260_1;
buffer_wire buffer_14260_1 (.in(n14260_0), .out(n14260_1));
wire n14261; //CHANY 4 (7,5) #63
wire n14261_0;
wire n14261_1;
buffer_wire buffer_14261_1 (.in(n14261_0), .out(n14261_1));
wire n14262; //CHANY 4 (7,5) #70
wire n14262_0;
wire n14262_1;
buffer_wire buffer_14262_1 (.in(n14262_0), .out(n14262_1));
wire n14263; //CHANY 4 (7,5) #71
wire n14263_0;
wire n14263_1;
buffer_wire buffer_14263_1 (.in(n14263_0), .out(n14263_1));
wire n14264; //CHANY 4 (7,5) #78
wire n14264_0;
wire n14264_1;
buffer_wire buffer_14264_1 (.in(n14264_0), .out(n14264_1));
wire n14265; //CHANY 4 (7,5) #79
wire n14265_0;
wire n14265_1;
buffer_wire buffer_14265_1 (.in(n14265_0), .out(n14265_1));
wire n14266; //CHANY 5 (7,5) #86
wire n14266_0;
wire n14266_1;
buffer_wire buffer_14266_1 (.in(n14266_0), .out(n14266_1));
wire n14267; //CHANY 5 (7,5) #87
wire n14267_0;
wire n14267_1;
buffer_wire buffer_14267_1 (.in(n14267_0), .out(n14267_1));
wire n14268; //CHANY 4 (7,6) #0
wire n14268_0;
wire n14268_1;
buffer_wire buffer_14268_1 (.in(n14268_0), .out(n14268_1));
wire n14269; //CHANY 4 (7,6) #1
wire n14269_0;
wire n14269_1;
buffer_wire buffer_14269_1 (.in(n14269_0), .out(n14269_1));
wire n14270; //CHANY 4 (7,6) #8
wire n14270_0;
wire n14270_1;
buffer_wire buffer_14270_1 (.in(n14270_0), .out(n14270_1));
wire n14271; //CHANY 4 (7,6) #9
wire n14271_0;
wire n14271_1;
buffer_wire buffer_14271_1 (.in(n14271_0), .out(n14271_1));
wire n14272; //CHANY 4 (7,6) #16
wire n14272_0;
wire n14272_1;
buffer_wire buffer_14272_1 (.in(n14272_0), .out(n14272_1));
wire n14273; //CHANY 4 (7,6) #17
wire n14273_0;
wire n14273_1;
buffer_wire buffer_14273_1 (.in(n14273_0), .out(n14273_1));
wire n14274; //CHANY 4 (7,6) #24
wire n14274_0;
wire n14274_1;
buffer_wire buffer_14274_1 (.in(n14274_0), .out(n14274_1));
wire n14275; //CHANY 4 (7,6) #25
wire n14275_0;
wire n14275_1;
buffer_wire buffer_14275_1 (.in(n14275_0), .out(n14275_1));
wire n14276; //CHANY 4 (7,6) #32
wire n14276_0;
wire n14276_1;
buffer_wire buffer_14276_1 (.in(n14276_0), .out(n14276_1));
wire n14277; //CHANY 4 (7,6) #33
wire n14277_0;
wire n14277_1;
buffer_wire buffer_14277_1 (.in(n14277_0), .out(n14277_1));
wire n14278; //CHANY 4 (7,6) #40
wire n14278_0;
wire n14278_1;
buffer_wire buffer_14278_1 (.in(n14278_0), .out(n14278_1));
wire n14279; //CHANY 4 (7,6) #41
wire n14279_0;
wire n14279_1;
buffer_wire buffer_14279_1 (.in(n14279_0), .out(n14279_1));
wire n14280; //CHANY 4 (7,6) #48
wire n14280_0;
wire n14280_1;
buffer_wire buffer_14280_1 (.in(n14280_0), .out(n14280_1));
wire n14281; //CHANY 4 (7,6) #49
wire n14281_0;
wire n14281_1;
buffer_wire buffer_14281_1 (.in(n14281_0), .out(n14281_1));
wire n14282; //CHANY 4 (7,6) #56
wire n14282_0;
wire n14282_1;
buffer_wire buffer_14282_1 (.in(n14282_0), .out(n14282_1));
wire n14283; //CHANY 4 (7,6) #57
wire n14283_0;
wire n14283_1;
buffer_wire buffer_14283_1 (.in(n14283_0), .out(n14283_1));
wire n14284; //CHANY 4 (7,6) #64
wire n14284_0;
wire n14284_1;
buffer_wire buffer_14284_1 (.in(n14284_0), .out(n14284_1));
wire n14285; //CHANY 4 (7,6) #65
wire n14285_0;
wire n14285_1;
buffer_wire buffer_14285_1 (.in(n14285_0), .out(n14285_1));
wire n14286; //CHANY 4 (7,6) #72
wire n14286_0;
wire n14286_1;
buffer_wire buffer_14286_1 (.in(n14286_0), .out(n14286_1));
wire n14287; //CHANY 4 (7,6) #73
wire n14287_0;
wire n14287_1;
buffer_wire buffer_14287_1 (.in(n14287_0), .out(n14287_1));
wire n14288; //CHANY 4 (7,6) #88
wire n14288_0;
wire n14288_1;
buffer_wire buffer_14288_1 (.in(n14288_0), .out(n14288_1));
wire n14289; //CHANY 4 (7,6) #89
wire n14289_0;
wire n14289_1;
buffer_wire buffer_14289_1 (.in(n14289_0), .out(n14289_1));
wire n14290; //CHANY 3 (7,7) #2
wire n14290_0;
wire n14291; //CHANY 3 (7,7) #3
wire n14291_0;
wire n14292; //CHANY 3 (7,7) #10
wire n14292_0;
wire n14293; //CHANY 3 (7,7) #11
wire n14293_0;
wire n14294; //CHANY 3 (7,7) #18
wire n14294_0;
wire n14295; //CHANY 3 (7,7) #19
wire n14295_0;
wire n14296; //CHANY 3 (7,7) #26
wire n14296_0;
wire n14297; //CHANY 3 (7,7) #27
wire n14297_0;
wire n14298; //CHANY 3 (7,7) #34
wire n14298_0;
wire n14299; //CHANY 3 (7,7) #35
wire n14299_0;
wire n14300; //CHANY 3 (7,7) #42
wire n14300_0;
wire n14301; //CHANY 3 (7,7) #43
wire n14301_0;
wire n14302; //CHANY 3 (7,7) #50
wire n14302_0;
wire n14303; //CHANY 3 (7,7) #51
wire n14303_0;
wire n14304; //CHANY 3 (7,7) #58
wire n14304_0;
wire n14305; //CHANY 3 (7,7) #59
wire n14305_0;
wire n14306; //CHANY 3 (7,7) #66
wire n14306_0;
wire n14307; //CHANY 3 (7,7) #67
wire n14307_0;
wire n14308; //CHANY 3 (7,7) #74
wire n14308_0;
wire n14309; //CHANY 3 (7,7) #75
wire n14309_0;
wire n14310; //CHANY 3 (7,7) #90
wire n14310_0;
wire n14311; //CHANY 3 (7,7) #91
wire n14311_0;
wire n14312; //CHANY 2 (7,8) #4
wire n14312_0;
wire n14313; //CHANY 2 (7,8) #5
wire n14313_0;
wire n14314; //CHANY 2 (7,8) #12
wire n14314_0;
wire n14315; //CHANY 2 (7,8) #13
wire n14315_0;
wire n14316; //CHANY 2 (7,8) #20
wire n14316_0;
wire n14317; //CHANY 2 (7,8) #21
wire n14317_0;
wire n14318; //CHANY 2 (7,8) #28
wire n14318_0;
wire n14319; //CHANY 2 (7,8) #29
wire n14319_0;
wire n14320; //CHANY 2 (7,8) #36
wire n14320_0;
wire n14321; //CHANY 2 (7,8) #37
wire n14321_0;
wire n14322; //CHANY 2 (7,8) #44
wire n14322_0;
wire n14323; //CHANY 2 (7,8) #45
wire n14323_0;
wire n14324; //CHANY 2 (7,8) #52
wire n14324_0;
wire n14325; //CHANY 2 (7,8) #53
wire n14325_0;
wire n14326; //CHANY 2 (7,8) #60
wire n14326_0;
wire n14327; //CHANY 2 (7,8) #61
wire n14327_0;
wire n14328; //CHANY 2 (7,8) #68
wire n14328_0;
wire n14329; //CHANY 2 (7,8) #69
wire n14329_0;
wire n14330; //CHANY 2 (7,8) #76
wire n14330_0;
wire n14331; //CHANY 2 (7,8) #77
wire n14331_0;
wire n14332; //CHANY 1 (7,9) #6
wire n14332_0;
wire n14333; //CHANY 1 (7,9) #7
wire n14333_0;
wire n14334; //CHANY 1 (7,9) #14
wire n14334_0;
wire n14335; //CHANY 1 (7,9) #15
wire n14335_0;
wire n14336; //CHANY 1 (7,9) #22
wire n14336_0;
wire n14337; //CHANY 1 (7,9) #23
wire n14337_0;
wire n14338; //CHANY 1 (7,9) #30
wire n14338_0;
wire n14339; //CHANY 1 (7,9) #31
wire n14339_0;
wire n14340; //CHANY 1 (7,9) #38
wire n14340_0;
wire n14341; //CHANY 1 (7,9) #39
wire n14341_0;
wire n14342; //CHANY 1 (7,9) #46
wire n14342_0;
wire n14343; //CHANY 1 (7,9) #47
wire n14343_0;
wire n14344; //CHANY 1 (7,9) #54
wire n14344_0;
wire n14345; //CHANY 1 (7,9) #55
wire n14345_0;
wire n14346; //CHANY 1 (7,9) #62
wire n14346_0;
wire n14347; //CHANY 1 (7,9) #63
wire n14347_0;
wire n14348; //CHANY 1 (7,9) #70
wire n14348_0;
wire n14349; //CHANY 1 (7,9) #71
wire n14349_0;
wire n14350; //CHANY 1 (7,9) #78
wire n14350_0;
wire n14351; //CHANY 1 (7,9) #79
wire n14351_0;
wire n14352; //CHANY 4 (8,1) #0
wire n14352_0;
wire n14352_1;
buffer_wire buffer_14352_1 (.in(n14352_0), .out(n14352_1));
wire n14353; //CHANY 4 (8,1) #1
wire n14353_0;
wire n14353_1;
buffer_wire buffer_14353_1 (.in(n14353_0), .out(n14353_1));
wire n14354; //CHANY 1 (8,1) #2
wire n14354_0;
wire n14355; //CHANY 1 (8,1) #3
wire n14355_0;
wire n14356; //CHANY 2 (8,1) #4
wire n14356_0;
wire n14357; //CHANY 2 (8,1) #5
wire n14357_0;
wire n14358; //CHANY 3 (8,1) #6
wire n14358_0;
wire n14359; //CHANY 3 (8,1) #7
wire n14359_0;
wire n14360; //CHANY 4 (8,1) #8
wire n14360_0;
wire n14360_1;
buffer_wire buffer_14360_1 (.in(n14360_0), .out(n14360_1));
wire n14361; //CHANY 4 (8,1) #9
wire n14361_0;
wire n14361_1;
buffer_wire buffer_14361_1 (.in(n14361_0), .out(n14361_1));
wire n14362; //CHANY 1 (8,1) #10
wire n14362_0;
wire n14363; //CHANY 1 (8,1) #11
wire n14363_0;
wire n14364; //CHANY 2 (8,1) #12
wire n14364_0;
wire n14365; //CHANY 2 (8,1) #13
wire n14365_0;
wire n14366; //CHANY 3 (8,1) #14
wire n14366_0;
wire n14367; //CHANY 3 (8,1) #15
wire n14367_0;
wire n14368; //CHANY 4 (8,1) #16
wire n14368_0;
wire n14368_1;
buffer_wire buffer_14368_1 (.in(n14368_0), .out(n14368_1));
wire n14369; //CHANY 4 (8,1) #17
wire n14369_0;
wire n14369_1;
buffer_wire buffer_14369_1 (.in(n14369_0), .out(n14369_1));
wire n14370; //CHANY 1 (8,1) #18
wire n14370_0;
wire n14371; //CHANY 1 (8,1) #19
wire n14371_0;
wire n14372; //CHANY 2 (8,1) #20
wire n14372_0;
wire n14373; //CHANY 2 (8,1) #21
wire n14373_0;
wire n14374; //CHANY 3 (8,1) #22
wire n14374_0;
wire n14375; //CHANY 3 (8,1) #23
wire n14375_0;
wire n14376; //CHANY 4 (8,1) #24
wire n14376_0;
wire n14376_1;
buffer_wire buffer_14376_1 (.in(n14376_0), .out(n14376_1));
wire n14377; //CHANY 4 (8,1) #25
wire n14377_0;
wire n14377_1;
buffer_wire buffer_14377_1 (.in(n14377_0), .out(n14377_1));
wire n14378; //CHANY 1 (8,1) #26
wire n14378_0;
wire n14379; //CHANY 1 (8,1) #27
wire n14379_0;
wire n14380; //CHANY 2 (8,1) #28
wire n14380_0;
wire n14381; //CHANY 2 (8,1) #29
wire n14381_0;
wire n14382; //CHANY 3 (8,1) #30
wire n14382_0;
wire n14383; //CHANY 3 (8,1) #31
wire n14383_0;
wire n14384; //CHANY 4 (8,1) #32
wire n14384_0;
wire n14384_1;
buffer_wire buffer_14384_1 (.in(n14384_0), .out(n14384_1));
wire n14385; //CHANY 4 (8,1) #33
wire n14385_0;
wire n14385_1;
buffer_wire buffer_14385_1 (.in(n14385_0), .out(n14385_1));
wire n14386; //CHANY 1 (8,1) #34
wire n14386_0;
wire n14387; //CHANY 1 (8,1) #35
wire n14387_0;
wire n14388; //CHANY 2 (8,1) #36
wire n14388_0;
wire n14389; //CHANY 2 (8,1) #37
wire n14389_0;
wire n14390; //CHANY 3 (8,1) #38
wire n14390_0;
wire n14391; //CHANY 3 (8,1) #39
wire n14391_0;
wire n14392; //CHANY 4 (8,1) #40
wire n14392_0;
wire n14392_1;
buffer_wire buffer_14392_1 (.in(n14392_0), .out(n14392_1));
wire n14393; //CHANY 4 (8,1) #41
wire n14393_0;
wire n14393_1;
buffer_wire buffer_14393_1 (.in(n14393_0), .out(n14393_1));
wire n14394; //CHANY 1 (8,1) #42
wire n14394_0;
wire n14395; //CHANY 1 (8,1) #43
wire n14395_0;
wire n14396; //CHANY 2 (8,1) #44
wire n14396_0;
wire n14397; //CHANY 2 (8,1) #45
wire n14397_0;
wire n14398; //CHANY 3 (8,1) #46
wire n14398_0;
wire n14399; //CHANY 3 (8,1) #47
wire n14399_0;
wire n14400; //CHANY 4 (8,1) #48
wire n14400_0;
wire n14400_1;
buffer_wire buffer_14400_1 (.in(n14400_0), .out(n14400_1));
wire n14401; //CHANY 4 (8,1) #49
wire n14401_0;
wire n14401_1;
buffer_wire buffer_14401_1 (.in(n14401_0), .out(n14401_1));
wire n14402; //CHANY 1 (8,1) #50
wire n14402_0;
wire n14403; //CHANY 1 (8,1) #51
wire n14403_0;
wire n14404; //CHANY 2 (8,1) #52
wire n14404_0;
wire n14405; //CHANY 2 (8,1) #53
wire n14405_0;
wire n14406; //CHANY 3 (8,1) #54
wire n14406_0;
wire n14407; //CHANY 3 (8,1) #55
wire n14407_0;
wire n14408; //CHANY 4 (8,1) #56
wire n14408_0;
wire n14408_1;
buffer_wire buffer_14408_1 (.in(n14408_0), .out(n14408_1));
wire n14409; //CHANY 4 (8,1) #57
wire n14409_0;
wire n14409_1;
buffer_wire buffer_14409_1 (.in(n14409_0), .out(n14409_1));
wire n14410; //CHANY 1 (8,1) #58
wire n14410_0;
wire n14411; //CHANY 1 (8,1) #59
wire n14411_0;
wire n14412; //CHANY 2 (8,1) #60
wire n14412_0;
wire n14413; //CHANY 2 (8,1) #61
wire n14413_0;
wire n14414; //CHANY 3 (8,1) #62
wire n14414_0;
wire n14415; //CHANY 3 (8,1) #63
wire n14415_0;
wire n14416; //CHANY 4 (8,1) #64
wire n14416_0;
wire n14416_1;
buffer_wire buffer_14416_1 (.in(n14416_0), .out(n14416_1));
wire n14417; //CHANY 4 (8,1) #65
wire n14417_0;
wire n14417_1;
buffer_wire buffer_14417_1 (.in(n14417_0), .out(n14417_1));
wire n14418; //CHANY 1 (8,1) #66
wire n14418_0;
wire n14419; //CHANY 1 (8,1) #67
wire n14419_0;
wire n14420; //CHANY 2 (8,1) #68
wire n14420_0;
wire n14421; //CHANY 2 (8,1) #69
wire n14421_0;
wire n14422; //CHANY 3 (8,1) #70
wire n14422_0;
wire n14423; //CHANY 3 (8,1) #71
wire n14423_0;
wire n14424; //CHANY 4 (8,1) #72
wire n14424_0;
wire n14424_1;
buffer_wire buffer_14424_1 (.in(n14424_0), .out(n14424_1));
wire n14425; //CHANY 4 (8,1) #73
wire n14425_0;
wire n14425_1;
buffer_wire buffer_14425_1 (.in(n14425_0), .out(n14425_1));
wire n14426; //CHANY 1 (8,1) #74
wire n14426_0;
wire n14427; //CHANY 1 (8,1) #75
wire n14427_0;
wire n14428; //CHANY 2 (8,1) #76
wire n14428_0;
wire n14429; //CHANY 2 (8,1) #77
wire n14429_0;
wire n14430; //CHANY 3 (8,1) #78
wire n14430_0;
wire n14431; //CHANY 3 (8,1) #79
wire n14431_0;
wire n14432; //CHANY 9 (8,1) #80
wire n14432_0;
wire n14432_1;
wire n14432_2;
buffer_wire buffer_14432_2 (.in(n14432_1), .out(n14432_2));
buffer_wire buffer_14432_1 (.in(n14432_0), .out(n14432_1));
wire n14433; //CHANY 9 (8,1) #81
wire n14433_0;
wire n14433_1;
wire n14433_2;
buffer_wire buffer_14433_2 (.in(n14433_1), .out(n14433_2));
buffer_wire buffer_14433_1 (.in(n14433_0), .out(n14433_1));
wire n14434; //CHANY 1 (8,1) #82
wire n14434_0;
wire n14435; //CHANY 1 (8,1) #83
wire n14435_0;
wire n14436; //CHANY 2 (8,1) #84
wire n14436_0;
wire n14437; //CHANY 2 (8,1) #85
wire n14437_0;
wire n14438; //CHANY 3 (8,1) #86
wire n14438_0;
wire n14439; //CHANY 3 (8,1) #87
wire n14439_0;
wire n14440; //CHANY 4 (8,1) #88
wire n14440_0;
wire n14440_1;
buffer_wire buffer_14440_1 (.in(n14440_0), .out(n14440_1));
wire n14441; //CHANY 4 (8,1) #89
wire n14441_0;
wire n14441_1;
buffer_wire buffer_14441_1 (.in(n14441_0), .out(n14441_1));
wire n14442; //CHANY 5 (8,1) #90
wire n14442_0;
wire n14442_1;
buffer_wire buffer_14442_1 (.in(n14442_0), .out(n14442_1));
wire n14443; //CHANY 5 (8,1) #91
wire n14443_0;
wire n14443_1;
buffer_wire buffer_14443_1 (.in(n14443_0), .out(n14443_1));
wire n14444; //CHANY 4 (8,2) #2
wire n14444_0;
wire n14444_1;
buffer_wire buffer_14444_1 (.in(n14444_0), .out(n14444_1));
wire n14445; //CHANY 4 (8,2) #3
wire n14445_0;
wire n14445_1;
buffer_wire buffer_14445_1 (.in(n14445_0), .out(n14445_1));
wire n14446; //CHANY 4 (8,2) #10
wire n14446_0;
wire n14446_1;
buffer_wire buffer_14446_1 (.in(n14446_0), .out(n14446_1));
wire n14447; //CHANY 4 (8,2) #11
wire n14447_0;
wire n14447_1;
buffer_wire buffer_14447_1 (.in(n14447_0), .out(n14447_1));
wire n14448; //CHANY 4 (8,2) #18
wire n14448_0;
wire n14448_1;
buffer_wire buffer_14448_1 (.in(n14448_0), .out(n14448_1));
wire n14449; //CHANY 4 (8,2) #19
wire n14449_0;
wire n14449_1;
buffer_wire buffer_14449_1 (.in(n14449_0), .out(n14449_1));
wire n14450; //CHANY 4 (8,2) #26
wire n14450_0;
wire n14450_1;
buffer_wire buffer_14450_1 (.in(n14450_0), .out(n14450_1));
wire n14451; //CHANY 4 (8,2) #27
wire n14451_0;
wire n14451_1;
buffer_wire buffer_14451_1 (.in(n14451_0), .out(n14451_1));
wire n14452; //CHANY 4 (8,2) #34
wire n14452_0;
wire n14452_1;
buffer_wire buffer_14452_1 (.in(n14452_0), .out(n14452_1));
wire n14453; //CHANY 4 (8,2) #35
wire n14453_0;
wire n14453_1;
buffer_wire buffer_14453_1 (.in(n14453_0), .out(n14453_1));
wire n14454; //CHANY 4 (8,2) #42
wire n14454_0;
wire n14454_1;
buffer_wire buffer_14454_1 (.in(n14454_0), .out(n14454_1));
wire n14455; //CHANY 4 (8,2) #43
wire n14455_0;
wire n14455_1;
buffer_wire buffer_14455_1 (.in(n14455_0), .out(n14455_1));
wire n14456; //CHANY 4 (8,2) #50
wire n14456_0;
wire n14456_1;
buffer_wire buffer_14456_1 (.in(n14456_0), .out(n14456_1));
wire n14457; //CHANY 4 (8,2) #51
wire n14457_0;
wire n14457_1;
buffer_wire buffer_14457_1 (.in(n14457_0), .out(n14457_1));
wire n14458; //CHANY 4 (8,2) #58
wire n14458_0;
wire n14458_1;
buffer_wire buffer_14458_1 (.in(n14458_0), .out(n14458_1));
wire n14459; //CHANY 4 (8,2) #59
wire n14459_0;
wire n14459_1;
buffer_wire buffer_14459_1 (.in(n14459_0), .out(n14459_1));
wire n14460; //CHANY 4 (8,2) #66
wire n14460_0;
wire n14460_1;
buffer_wire buffer_14460_1 (.in(n14460_0), .out(n14460_1));
wire n14461; //CHANY 4 (8,2) #67
wire n14461_0;
wire n14461_1;
buffer_wire buffer_14461_1 (.in(n14461_0), .out(n14461_1));
wire n14462; //CHANY 4 (8,2) #74
wire n14462_0;
wire n14462_1;
buffer_wire buffer_14462_1 (.in(n14462_0), .out(n14462_1));
wire n14463; //CHANY 4 (8,2) #75
wire n14463_0;
wire n14463_1;
buffer_wire buffer_14463_1 (.in(n14463_0), .out(n14463_1));
wire n14464; //CHANY 8 (8,2) #82
wire n14464_0;
wire n14464_1;
wire n14464_2;
buffer_wire buffer_14464_2 (.in(n14464_1), .out(n14464_2));
buffer_wire buffer_14464_1 (.in(n14464_0), .out(n14464_1));
wire n14465; //CHANY 8 (8,2) #83
wire n14465_0;
wire n14465_1;
wire n14465_2;
buffer_wire buffer_14465_2 (.in(n14465_1), .out(n14465_2));
buffer_wire buffer_14465_1 (.in(n14465_0), .out(n14465_1));
wire n14466; //CHANY 4 (8,3) #4
wire n14466_0;
wire n14466_1;
buffer_wire buffer_14466_1 (.in(n14466_0), .out(n14466_1));
wire n14467; //CHANY 4 (8,3) #5
wire n14467_0;
wire n14467_1;
buffer_wire buffer_14467_1 (.in(n14467_0), .out(n14467_1));
wire n14468; //CHANY 4 (8,3) #12
wire n14468_0;
wire n14468_1;
buffer_wire buffer_14468_1 (.in(n14468_0), .out(n14468_1));
wire n14469; //CHANY 4 (8,3) #13
wire n14469_0;
wire n14469_1;
buffer_wire buffer_14469_1 (.in(n14469_0), .out(n14469_1));
wire n14470; //CHANY 4 (8,3) #20
wire n14470_0;
wire n14470_1;
buffer_wire buffer_14470_1 (.in(n14470_0), .out(n14470_1));
wire n14471; //CHANY 4 (8,3) #21
wire n14471_0;
wire n14471_1;
buffer_wire buffer_14471_1 (.in(n14471_0), .out(n14471_1));
wire n14472; //CHANY 4 (8,3) #28
wire n14472_0;
wire n14472_1;
buffer_wire buffer_14472_1 (.in(n14472_0), .out(n14472_1));
wire n14473; //CHANY 4 (8,3) #29
wire n14473_0;
wire n14473_1;
buffer_wire buffer_14473_1 (.in(n14473_0), .out(n14473_1));
wire n14474; //CHANY 4 (8,3) #36
wire n14474_0;
wire n14474_1;
buffer_wire buffer_14474_1 (.in(n14474_0), .out(n14474_1));
wire n14475; //CHANY 4 (8,3) #37
wire n14475_0;
wire n14475_1;
buffer_wire buffer_14475_1 (.in(n14475_0), .out(n14475_1));
wire n14476; //CHANY 4 (8,3) #44
wire n14476_0;
wire n14476_1;
buffer_wire buffer_14476_1 (.in(n14476_0), .out(n14476_1));
wire n14477; //CHANY 4 (8,3) #45
wire n14477_0;
wire n14477_1;
buffer_wire buffer_14477_1 (.in(n14477_0), .out(n14477_1));
wire n14478; //CHANY 4 (8,3) #52
wire n14478_0;
wire n14478_1;
buffer_wire buffer_14478_1 (.in(n14478_0), .out(n14478_1));
wire n14479; //CHANY 4 (8,3) #53
wire n14479_0;
wire n14479_1;
buffer_wire buffer_14479_1 (.in(n14479_0), .out(n14479_1));
wire n14480; //CHANY 4 (8,3) #60
wire n14480_0;
wire n14480_1;
buffer_wire buffer_14480_1 (.in(n14480_0), .out(n14480_1));
wire n14481; //CHANY 4 (8,3) #61
wire n14481_0;
wire n14481_1;
buffer_wire buffer_14481_1 (.in(n14481_0), .out(n14481_1));
wire n14482; //CHANY 4 (8,3) #68
wire n14482_0;
wire n14482_1;
buffer_wire buffer_14482_1 (.in(n14482_0), .out(n14482_1));
wire n14483; //CHANY 4 (8,3) #69
wire n14483_0;
wire n14483_1;
buffer_wire buffer_14483_1 (.in(n14483_0), .out(n14483_1));
wire n14484; //CHANY 4 (8,3) #76
wire n14484_0;
wire n14484_1;
buffer_wire buffer_14484_1 (.in(n14484_0), .out(n14484_1));
wire n14485; //CHANY 4 (8,3) #77
wire n14485_0;
wire n14485_1;
buffer_wire buffer_14485_1 (.in(n14485_0), .out(n14485_1));
wire n14486; //CHANY 7 (8,3) #84
wire n14486_0;
wire n14486_1;
wire n14486_2;
buffer_wire buffer_14486_2 (.in(n14486_1), .out(n14486_2));
buffer_wire buffer_14486_1 (.in(n14486_0), .out(n14486_1));
wire n14487; //CHANY 7 (8,3) #85
wire n14487_0;
wire n14487_1;
wire n14487_2;
buffer_wire buffer_14487_2 (.in(n14487_1), .out(n14487_2));
buffer_wire buffer_14487_1 (.in(n14487_0), .out(n14487_1));
wire n14488; //CHANY 4 (8,4) #6
wire n14488_0;
wire n14488_1;
buffer_wire buffer_14488_1 (.in(n14488_0), .out(n14488_1));
wire n14489; //CHANY 4 (8,4) #7
wire n14489_0;
wire n14489_1;
buffer_wire buffer_14489_1 (.in(n14489_0), .out(n14489_1));
wire n14490; //CHANY 4 (8,4) #14
wire n14490_0;
wire n14490_1;
buffer_wire buffer_14490_1 (.in(n14490_0), .out(n14490_1));
wire n14491; //CHANY 4 (8,4) #15
wire n14491_0;
wire n14491_1;
buffer_wire buffer_14491_1 (.in(n14491_0), .out(n14491_1));
wire n14492; //CHANY 4 (8,4) #22
wire n14492_0;
wire n14492_1;
buffer_wire buffer_14492_1 (.in(n14492_0), .out(n14492_1));
wire n14493; //CHANY 4 (8,4) #23
wire n14493_0;
wire n14493_1;
buffer_wire buffer_14493_1 (.in(n14493_0), .out(n14493_1));
wire n14494; //CHANY 4 (8,4) #30
wire n14494_0;
wire n14494_1;
buffer_wire buffer_14494_1 (.in(n14494_0), .out(n14494_1));
wire n14495; //CHANY 4 (8,4) #31
wire n14495_0;
wire n14495_1;
buffer_wire buffer_14495_1 (.in(n14495_0), .out(n14495_1));
wire n14496; //CHANY 4 (8,4) #38
wire n14496_0;
wire n14496_1;
buffer_wire buffer_14496_1 (.in(n14496_0), .out(n14496_1));
wire n14497; //CHANY 4 (8,4) #39
wire n14497_0;
wire n14497_1;
buffer_wire buffer_14497_1 (.in(n14497_0), .out(n14497_1));
wire n14498; //CHANY 4 (8,4) #46
wire n14498_0;
wire n14498_1;
buffer_wire buffer_14498_1 (.in(n14498_0), .out(n14498_1));
wire n14499; //CHANY 4 (8,4) #47
wire n14499_0;
wire n14499_1;
buffer_wire buffer_14499_1 (.in(n14499_0), .out(n14499_1));
wire n14500; //CHANY 4 (8,4) #54
wire n14500_0;
wire n14500_1;
buffer_wire buffer_14500_1 (.in(n14500_0), .out(n14500_1));
wire n14501; //CHANY 4 (8,4) #55
wire n14501_0;
wire n14501_1;
buffer_wire buffer_14501_1 (.in(n14501_0), .out(n14501_1));
wire n14502; //CHANY 4 (8,4) #62
wire n14502_0;
wire n14502_1;
buffer_wire buffer_14502_1 (.in(n14502_0), .out(n14502_1));
wire n14503; //CHANY 4 (8,4) #63
wire n14503_0;
wire n14503_1;
buffer_wire buffer_14503_1 (.in(n14503_0), .out(n14503_1));
wire n14504; //CHANY 4 (8,4) #70
wire n14504_0;
wire n14504_1;
buffer_wire buffer_14504_1 (.in(n14504_0), .out(n14504_1));
wire n14505; //CHANY 4 (8,4) #71
wire n14505_0;
wire n14505_1;
buffer_wire buffer_14505_1 (.in(n14505_0), .out(n14505_1));
wire n14506; //CHANY 4 (8,4) #78
wire n14506_0;
wire n14506_1;
buffer_wire buffer_14506_1 (.in(n14506_0), .out(n14506_1));
wire n14507; //CHANY 4 (8,4) #79
wire n14507_0;
wire n14507_1;
buffer_wire buffer_14507_1 (.in(n14507_0), .out(n14507_1));
wire n14508; //CHANY 6 (8,4) #86
wire n14508_0;
wire n14508_1;
buffer_wire buffer_14508_1 (.in(n14508_0), .out(n14508_1));
wire n14509; //CHANY 6 (8,4) #87
wire n14509_0;
wire n14509_1;
buffer_wire buffer_14509_1 (.in(n14509_0), .out(n14509_1));
wire n14510; //CHANY 4 (8,5) #0
wire n14510_0;
wire n14510_1;
buffer_wire buffer_14510_1 (.in(n14510_0), .out(n14510_1));
wire n14511; //CHANY 4 (8,5) #1
wire n14511_0;
wire n14511_1;
buffer_wire buffer_14511_1 (.in(n14511_0), .out(n14511_1));
wire n14512; //CHANY 4 (8,5) #8
wire n14512_0;
wire n14512_1;
buffer_wire buffer_14512_1 (.in(n14512_0), .out(n14512_1));
wire n14513; //CHANY 4 (8,5) #9
wire n14513_0;
wire n14513_1;
buffer_wire buffer_14513_1 (.in(n14513_0), .out(n14513_1));
wire n14514; //CHANY 4 (8,5) #16
wire n14514_0;
wire n14514_1;
buffer_wire buffer_14514_1 (.in(n14514_0), .out(n14514_1));
wire n14515; //CHANY 4 (8,5) #17
wire n14515_0;
wire n14515_1;
buffer_wire buffer_14515_1 (.in(n14515_0), .out(n14515_1));
wire n14516; //CHANY 4 (8,5) #24
wire n14516_0;
wire n14516_1;
buffer_wire buffer_14516_1 (.in(n14516_0), .out(n14516_1));
wire n14517; //CHANY 4 (8,5) #25
wire n14517_0;
wire n14517_1;
buffer_wire buffer_14517_1 (.in(n14517_0), .out(n14517_1));
wire n14518; //CHANY 4 (8,5) #32
wire n14518_0;
wire n14518_1;
buffer_wire buffer_14518_1 (.in(n14518_0), .out(n14518_1));
wire n14519; //CHANY 4 (8,5) #33
wire n14519_0;
wire n14519_1;
buffer_wire buffer_14519_1 (.in(n14519_0), .out(n14519_1));
wire n14520; //CHANY 4 (8,5) #40
wire n14520_0;
wire n14520_1;
buffer_wire buffer_14520_1 (.in(n14520_0), .out(n14520_1));
wire n14521; //CHANY 4 (8,5) #41
wire n14521_0;
wire n14521_1;
buffer_wire buffer_14521_1 (.in(n14521_0), .out(n14521_1));
wire n14522; //CHANY 4 (8,5) #48
wire n14522_0;
wire n14522_1;
buffer_wire buffer_14522_1 (.in(n14522_0), .out(n14522_1));
wire n14523; //CHANY 4 (8,5) #49
wire n14523_0;
wire n14523_1;
buffer_wire buffer_14523_1 (.in(n14523_0), .out(n14523_1));
wire n14524; //CHANY 4 (8,5) #56
wire n14524_0;
wire n14524_1;
buffer_wire buffer_14524_1 (.in(n14524_0), .out(n14524_1));
wire n14525; //CHANY 4 (8,5) #57
wire n14525_0;
wire n14525_1;
buffer_wire buffer_14525_1 (.in(n14525_0), .out(n14525_1));
wire n14526; //CHANY 4 (8,5) #64
wire n14526_0;
wire n14526_1;
buffer_wire buffer_14526_1 (.in(n14526_0), .out(n14526_1));
wire n14527; //CHANY 4 (8,5) #65
wire n14527_0;
wire n14527_1;
buffer_wire buffer_14527_1 (.in(n14527_0), .out(n14527_1));
wire n14528; //CHANY 4 (8,5) #72
wire n14528_0;
wire n14528_1;
buffer_wire buffer_14528_1 (.in(n14528_0), .out(n14528_1));
wire n14529; //CHANY 4 (8,5) #73
wire n14529_0;
wire n14529_1;
buffer_wire buffer_14529_1 (.in(n14529_0), .out(n14529_1));
wire n14530; //CHANY 5 (8,5) #88
wire n14530_0;
wire n14530_1;
buffer_wire buffer_14530_1 (.in(n14530_0), .out(n14530_1));
wire n14531; //CHANY 5 (8,5) #89
wire n14531_0;
wire n14531_1;
buffer_wire buffer_14531_1 (.in(n14531_0), .out(n14531_1));
wire n14532; //CHANY 4 (8,6) #2
wire n14532_0;
wire n14532_1;
buffer_wire buffer_14532_1 (.in(n14532_0), .out(n14532_1));
wire n14533; //CHANY 4 (8,6) #3
wire n14533_0;
wire n14533_1;
buffer_wire buffer_14533_1 (.in(n14533_0), .out(n14533_1));
wire n14534; //CHANY 4 (8,6) #10
wire n14534_0;
wire n14534_1;
buffer_wire buffer_14534_1 (.in(n14534_0), .out(n14534_1));
wire n14535; //CHANY 4 (8,6) #11
wire n14535_0;
wire n14535_1;
buffer_wire buffer_14535_1 (.in(n14535_0), .out(n14535_1));
wire n14536; //CHANY 4 (8,6) #18
wire n14536_0;
wire n14536_1;
buffer_wire buffer_14536_1 (.in(n14536_0), .out(n14536_1));
wire n14537; //CHANY 4 (8,6) #19
wire n14537_0;
wire n14537_1;
buffer_wire buffer_14537_1 (.in(n14537_0), .out(n14537_1));
wire n14538; //CHANY 4 (8,6) #26
wire n14538_0;
wire n14538_1;
buffer_wire buffer_14538_1 (.in(n14538_0), .out(n14538_1));
wire n14539; //CHANY 4 (8,6) #27
wire n14539_0;
wire n14539_1;
buffer_wire buffer_14539_1 (.in(n14539_0), .out(n14539_1));
wire n14540; //CHANY 4 (8,6) #34
wire n14540_0;
wire n14540_1;
buffer_wire buffer_14540_1 (.in(n14540_0), .out(n14540_1));
wire n14541; //CHANY 4 (8,6) #35
wire n14541_0;
wire n14541_1;
buffer_wire buffer_14541_1 (.in(n14541_0), .out(n14541_1));
wire n14542; //CHANY 4 (8,6) #42
wire n14542_0;
wire n14542_1;
buffer_wire buffer_14542_1 (.in(n14542_0), .out(n14542_1));
wire n14543; //CHANY 4 (8,6) #43
wire n14543_0;
wire n14543_1;
buffer_wire buffer_14543_1 (.in(n14543_0), .out(n14543_1));
wire n14544; //CHANY 4 (8,6) #50
wire n14544_0;
wire n14544_1;
buffer_wire buffer_14544_1 (.in(n14544_0), .out(n14544_1));
wire n14545; //CHANY 4 (8,6) #51
wire n14545_0;
wire n14545_1;
buffer_wire buffer_14545_1 (.in(n14545_0), .out(n14545_1));
wire n14546; //CHANY 4 (8,6) #58
wire n14546_0;
wire n14546_1;
buffer_wire buffer_14546_1 (.in(n14546_0), .out(n14546_1));
wire n14547; //CHANY 4 (8,6) #59
wire n14547_0;
wire n14547_1;
buffer_wire buffer_14547_1 (.in(n14547_0), .out(n14547_1));
wire n14548; //CHANY 4 (8,6) #66
wire n14548_0;
wire n14548_1;
buffer_wire buffer_14548_1 (.in(n14548_0), .out(n14548_1));
wire n14549; //CHANY 4 (8,6) #67
wire n14549_0;
wire n14549_1;
buffer_wire buffer_14549_1 (.in(n14549_0), .out(n14549_1));
wire n14550; //CHANY 4 (8,6) #74
wire n14550_0;
wire n14550_1;
buffer_wire buffer_14550_1 (.in(n14550_0), .out(n14550_1));
wire n14551; //CHANY 4 (8,6) #75
wire n14551_0;
wire n14551_1;
buffer_wire buffer_14551_1 (.in(n14551_0), .out(n14551_1));
wire n14552; //CHANY 4 (8,6) #90
wire n14552_0;
wire n14552_1;
buffer_wire buffer_14552_1 (.in(n14552_0), .out(n14552_1));
wire n14553; //CHANY 4 (8,6) #91
wire n14553_0;
wire n14553_1;
buffer_wire buffer_14553_1 (.in(n14553_0), .out(n14553_1));
wire n14554; //CHANY 3 (8,7) #4
wire n14554_0;
wire n14555; //CHANY 3 (8,7) #5
wire n14555_0;
wire n14556; //CHANY 3 (8,7) #12
wire n14556_0;
wire n14557; //CHANY 3 (8,7) #13
wire n14557_0;
wire n14558; //CHANY 3 (8,7) #20
wire n14558_0;
wire n14559; //CHANY 3 (8,7) #21
wire n14559_0;
wire n14560; //CHANY 3 (8,7) #28
wire n14560_0;
wire n14561; //CHANY 3 (8,7) #29
wire n14561_0;
wire n14562; //CHANY 3 (8,7) #36
wire n14562_0;
wire n14563; //CHANY 3 (8,7) #37
wire n14563_0;
wire n14564; //CHANY 3 (8,7) #44
wire n14564_0;
wire n14565; //CHANY 3 (8,7) #45
wire n14565_0;
wire n14566; //CHANY 3 (8,7) #52
wire n14566_0;
wire n14567; //CHANY 3 (8,7) #53
wire n14567_0;
wire n14568; //CHANY 3 (8,7) #60
wire n14568_0;
wire n14569; //CHANY 3 (8,7) #61
wire n14569_0;
wire n14570; //CHANY 3 (8,7) #68
wire n14570_0;
wire n14571; //CHANY 3 (8,7) #69
wire n14571_0;
wire n14572; //CHANY 3 (8,7) #76
wire n14572_0;
wire n14573; //CHANY 3 (8,7) #77
wire n14573_0;
wire n14574; //CHANY 2 (8,8) #6
wire n14574_0;
wire n14575; //CHANY 2 (8,8) #7
wire n14575_0;
wire n14576; //CHANY 2 (8,8) #14
wire n14576_0;
wire n14577; //CHANY 2 (8,8) #15
wire n14577_0;
wire n14578; //CHANY 2 (8,8) #22
wire n14578_0;
wire n14579; //CHANY 2 (8,8) #23
wire n14579_0;
wire n14580; //CHANY 2 (8,8) #30
wire n14580_0;
wire n14581; //CHANY 2 (8,8) #31
wire n14581_0;
wire n14582; //CHANY 2 (8,8) #38
wire n14582_0;
wire n14583; //CHANY 2 (8,8) #39
wire n14583_0;
wire n14584; //CHANY 2 (8,8) #46
wire n14584_0;
wire n14585; //CHANY 2 (8,8) #47
wire n14585_0;
wire n14586; //CHANY 2 (8,8) #54
wire n14586_0;
wire n14587; //CHANY 2 (8,8) #55
wire n14587_0;
wire n14588; //CHANY 2 (8,8) #62
wire n14588_0;
wire n14589; //CHANY 2 (8,8) #63
wire n14589_0;
wire n14590; //CHANY 2 (8,8) #70
wire n14590_0;
wire n14591; //CHANY 2 (8,8) #71
wire n14591_0;
wire n14592; //CHANY 2 (8,8) #78
wire n14592_0;
wire n14593; //CHANY 2 (8,8) #79
wire n14593_0;
wire n14594; //CHANY 1 (8,9) #0
wire n14594_0;
wire n14595; //CHANY 1 (8,9) #1
wire n14595_0;
wire n14596; //CHANY 1 (8,9) #8
wire n14596_0;
wire n14597; //CHANY 1 (8,9) #9
wire n14597_0;
wire n14598; //CHANY 1 (8,9) #16
wire n14598_0;
wire n14599; //CHANY 1 (8,9) #17
wire n14599_0;
wire n14600; //CHANY 1 (8,9) #24
wire n14600_0;
wire n14601; //CHANY 1 (8,9) #25
wire n14601_0;
wire n14602; //CHANY 1 (8,9) #32
wire n14602_0;
wire n14603; //CHANY 1 (8,9) #33
wire n14603_0;
wire n14604; //CHANY 1 (8,9) #40
wire n14604_0;
wire n14605; //CHANY 1 (8,9) #41
wire n14605_0;
wire n14606; //CHANY 1 (8,9) #48
wire n14606_0;
wire n14607; //CHANY 1 (8,9) #49
wire n14607_0;
wire n14608; //CHANY 1 (8,9) #56
wire n14608_0;
wire n14609; //CHANY 1 (8,9) #57
wire n14609_0;
wire n14610; //CHANY 1 (8,9) #64
wire n14610_0;
wire n14611; //CHANY 1 (8,9) #65
wire n14611_0;
wire n14612; //CHANY 1 (8,9) #72
wire n14612_0;
wire n14613; //CHANY 1 (8,9) #73
wire n14613_0;
wire n14614; //CHANY 3 (9,1) #0
wire n14614_0;
wire n14615; //CHANY 3 (9,1) #1
wire n14615_0;
wire n14616; //CHANY 4 (9,1) #2
wire n14616_0;
wire n14616_1;
buffer_wire buffer_14616_1 (.in(n14616_0), .out(n14616_1));
wire n14617; //CHANY 4 (9,1) #3
wire n14617_0;
wire n14617_1;
buffer_wire buffer_14617_1 (.in(n14617_0), .out(n14617_1));
wire n14618; //CHANY 1 (9,1) #4
wire n14618_0;
wire n14619; //CHANY 1 (9,1) #5
wire n14619_0;
wire n14620; //CHANY 2 (9,1) #6
wire n14620_0;
wire n14621; //CHANY 2 (9,1) #7
wire n14621_0;
wire n14622; //CHANY 3 (9,1) #8
wire n14622_0;
wire n14623; //CHANY 3 (9,1) #9
wire n14623_0;
wire n14624; //CHANY 4 (9,1) #10
wire n14624_0;
wire n14624_1;
buffer_wire buffer_14624_1 (.in(n14624_0), .out(n14624_1));
wire n14625; //CHANY 4 (9,1) #11
wire n14625_0;
wire n14625_1;
buffer_wire buffer_14625_1 (.in(n14625_0), .out(n14625_1));
wire n14626; //CHANY 1 (9,1) #12
wire n14626_0;
wire n14627; //CHANY 1 (9,1) #13
wire n14627_0;
wire n14628; //CHANY 2 (9,1) #14
wire n14628_0;
wire n14629; //CHANY 2 (9,1) #15
wire n14629_0;
wire n14630; //CHANY 3 (9,1) #16
wire n14630_0;
wire n14631; //CHANY 3 (9,1) #17
wire n14631_0;
wire n14632; //CHANY 4 (9,1) #18
wire n14632_0;
wire n14632_1;
buffer_wire buffer_14632_1 (.in(n14632_0), .out(n14632_1));
wire n14633; //CHANY 4 (9,1) #19
wire n14633_0;
wire n14633_1;
buffer_wire buffer_14633_1 (.in(n14633_0), .out(n14633_1));
wire n14634; //CHANY 1 (9,1) #20
wire n14634_0;
wire n14635; //CHANY 1 (9,1) #21
wire n14635_0;
wire n14636; //CHANY 2 (9,1) #22
wire n14636_0;
wire n14637; //CHANY 2 (9,1) #23
wire n14637_0;
wire n14638; //CHANY 3 (9,1) #24
wire n14638_0;
wire n14639; //CHANY 3 (9,1) #25
wire n14639_0;
wire n14640; //CHANY 4 (9,1) #26
wire n14640_0;
wire n14640_1;
buffer_wire buffer_14640_1 (.in(n14640_0), .out(n14640_1));
wire n14641; //CHANY 4 (9,1) #27
wire n14641_0;
wire n14641_1;
buffer_wire buffer_14641_1 (.in(n14641_0), .out(n14641_1));
wire n14642; //CHANY 1 (9,1) #28
wire n14642_0;
wire n14643; //CHANY 1 (9,1) #29
wire n14643_0;
wire n14644; //CHANY 2 (9,1) #30
wire n14644_0;
wire n14645; //CHANY 2 (9,1) #31
wire n14645_0;
wire n14646; //CHANY 3 (9,1) #32
wire n14646_0;
wire n14647; //CHANY 3 (9,1) #33
wire n14647_0;
wire n14648; //CHANY 4 (9,1) #34
wire n14648_0;
wire n14648_1;
buffer_wire buffer_14648_1 (.in(n14648_0), .out(n14648_1));
wire n14649; //CHANY 4 (9,1) #35
wire n14649_0;
wire n14649_1;
buffer_wire buffer_14649_1 (.in(n14649_0), .out(n14649_1));
wire n14650; //CHANY 1 (9,1) #36
wire n14650_0;
wire n14651; //CHANY 1 (9,1) #37
wire n14651_0;
wire n14652; //CHANY 2 (9,1) #38
wire n14652_0;
wire n14653; //CHANY 2 (9,1) #39
wire n14653_0;
wire n14654; //CHANY 3 (9,1) #40
wire n14654_0;
wire n14655; //CHANY 3 (9,1) #41
wire n14655_0;
wire n14656; //CHANY 4 (9,1) #42
wire n14656_0;
wire n14656_1;
buffer_wire buffer_14656_1 (.in(n14656_0), .out(n14656_1));
wire n14657; //CHANY 4 (9,1) #43
wire n14657_0;
wire n14657_1;
buffer_wire buffer_14657_1 (.in(n14657_0), .out(n14657_1));
wire n14658; //CHANY 1 (9,1) #44
wire n14658_0;
wire n14659; //CHANY 1 (9,1) #45
wire n14659_0;
wire n14660; //CHANY 2 (9,1) #46
wire n14660_0;
wire n14661; //CHANY 2 (9,1) #47
wire n14661_0;
wire n14662; //CHANY 3 (9,1) #48
wire n14662_0;
wire n14663; //CHANY 3 (9,1) #49
wire n14663_0;
wire n14664; //CHANY 4 (9,1) #50
wire n14664_0;
wire n14664_1;
buffer_wire buffer_14664_1 (.in(n14664_0), .out(n14664_1));
wire n14665; //CHANY 4 (9,1) #51
wire n14665_0;
wire n14665_1;
buffer_wire buffer_14665_1 (.in(n14665_0), .out(n14665_1));
wire n14666; //CHANY 1 (9,1) #52
wire n14666_0;
wire n14667; //CHANY 1 (9,1) #53
wire n14667_0;
wire n14668; //CHANY 2 (9,1) #54
wire n14668_0;
wire n14669; //CHANY 2 (9,1) #55
wire n14669_0;
wire n14670; //CHANY 3 (9,1) #56
wire n14670_0;
wire n14671; //CHANY 3 (9,1) #57
wire n14671_0;
wire n14672; //CHANY 4 (9,1) #58
wire n14672_0;
wire n14672_1;
buffer_wire buffer_14672_1 (.in(n14672_0), .out(n14672_1));
wire n14673; //CHANY 4 (9,1) #59
wire n14673_0;
wire n14673_1;
buffer_wire buffer_14673_1 (.in(n14673_0), .out(n14673_1));
wire n14674; //CHANY 1 (9,1) #60
wire n14674_0;
wire n14675; //CHANY 1 (9,1) #61
wire n14675_0;
wire n14676; //CHANY 2 (9,1) #62
wire n14676_0;
wire n14677; //CHANY 2 (9,1) #63
wire n14677_0;
wire n14678; //CHANY 3 (9,1) #64
wire n14678_0;
wire n14679; //CHANY 3 (9,1) #65
wire n14679_0;
wire n14680; //CHANY 4 (9,1) #66
wire n14680_0;
wire n14680_1;
buffer_wire buffer_14680_1 (.in(n14680_0), .out(n14680_1));
wire n14681; //CHANY 4 (9,1) #67
wire n14681_0;
wire n14681_1;
buffer_wire buffer_14681_1 (.in(n14681_0), .out(n14681_1));
wire n14682; //CHANY 1 (9,1) #68
wire n14682_0;
wire n14683; //CHANY 1 (9,1) #69
wire n14683_0;
wire n14684; //CHANY 2 (9,1) #70
wire n14684_0;
wire n14685; //CHANY 2 (9,1) #71
wire n14685_0;
wire n14686; //CHANY 3 (9,1) #72
wire n14686_0;
wire n14687; //CHANY 3 (9,1) #73
wire n14687_0;
wire n14688; //CHANY 4 (9,1) #74
wire n14688_0;
wire n14688_1;
buffer_wire buffer_14688_1 (.in(n14688_0), .out(n14688_1));
wire n14689; //CHANY 4 (9,1) #75
wire n14689_0;
wire n14689_1;
buffer_wire buffer_14689_1 (.in(n14689_0), .out(n14689_1));
wire n14690; //CHANY 1 (9,1) #76
wire n14690_0;
wire n14691; //CHANY 1 (9,1) #77
wire n14691_0;
wire n14692; //CHANY 2 (9,1) #78
wire n14692_0;
wire n14693; //CHANY 2 (9,1) #79
wire n14693_0;
wire n14694; //CHANY 9 (9,1) #80
wire n14694_0;
wire n14694_1;
wire n14694_2;
buffer_wire buffer_14694_2 (.in(n14694_1), .out(n14694_2));
buffer_wire buffer_14694_1 (.in(n14694_0), .out(n14694_1));
wire n14695; //CHANY 9 (9,1) #81
wire n14695_0;
wire n14695_1;
wire n14695_2;
buffer_wire buffer_14695_2 (.in(n14695_1), .out(n14695_2));
buffer_wire buffer_14695_1 (.in(n14695_0), .out(n14695_1));
wire n14696; //CHANY 9 (9,1) #82
wire n14696_0;
wire n14696_1;
wire n14696_2;
buffer_wire buffer_14696_2 (.in(n14696_1), .out(n14696_2));
buffer_wire buffer_14696_1 (.in(n14696_0), .out(n14696_1));
wire n14697; //CHANY 9 (9,1) #83
wire n14697_0;
wire n14697_1;
wire n14697_2;
buffer_wire buffer_14697_2 (.in(n14697_1), .out(n14697_2));
buffer_wire buffer_14697_1 (.in(n14697_0), .out(n14697_1));
wire n14698; //CHANY 1 (9,1) #84
wire n14698_0;
wire n14699; //CHANY 1 (9,1) #85
wire n14699_0;
wire n14700; //CHANY 2 (9,1) #86
wire n14700_0;
wire n14701; //CHANY 2 (9,1) #87
wire n14701_0;
wire n14702; //CHANY 3 (9,1) #88
wire n14702_0;
wire n14703; //CHANY 3 (9,1) #89
wire n14703_0;
wire n14704; //CHANY 4 (9,1) #90
wire n14704_0;
wire n14704_1;
buffer_wire buffer_14704_1 (.in(n14704_0), .out(n14704_1));
wire n14705; //CHANY 4 (9,1) #91
wire n14705_0;
wire n14705_1;
buffer_wire buffer_14705_1 (.in(n14705_0), .out(n14705_1));
wire n14706; //CHANY 4 (9,2) #4
wire n14706_0;
wire n14706_1;
buffer_wire buffer_14706_1 (.in(n14706_0), .out(n14706_1));
wire n14707; //CHANY 4 (9,2) #5
wire n14707_0;
wire n14707_1;
buffer_wire buffer_14707_1 (.in(n14707_0), .out(n14707_1));
wire n14708; //CHANY 4 (9,2) #12
wire n14708_0;
wire n14708_1;
buffer_wire buffer_14708_1 (.in(n14708_0), .out(n14708_1));
wire n14709; //CHANY 4 (9,2) #13
wire n14709_0;
wire n14709_1;
buffer_wire buffer_14709_1 (.in(n14709_0), .out(n14709_1));
wire n14710; //CHANY 4 (9,2) #20
wire n14710_0;
wire n14710_1;
buffer_wire buffer_14710_1 (.in(n14710_0), .out(n14710_1));
wire n14711; //CHANY 4 (9,2) #21
wire n14711_0;
wire n14711_1;
buffer_wire buffer_14711_1 (.in(n14711_0), .out(n14711_1));
wire n14712; //CHANY 4 (9,2) #28
wire n14712_0;
wire n14712_1;
buffer_wire buffer_14712_1 (.in(n14712_0), .out(n14712_1));
wire n14713; //CHANY 4 (9,2) #29
wire n14713_0;
wire n14713_1;
buffer_wire buffer_14713_1 (.in(n14713_0), .out(n14713_1));
wire n14714; //CHANY 4 (9,2) #36
wire n14714_0;
wire n14714_1;
buffer_wire buffer_14714_1 (.in(n14714_0), .out(n14714_1));
wire n14715; //CHANY 4 (9,2) #37
wire n14715_0;
wire n14715_1;
buffer_wire buffer_14715_1 (.in(n14715_0), .out(n14715_1));
wire n14716; //CHANY 4 (9,2) #44
wire n14716_0;
wire n14716_1;
buffer_wire buffer_14716_1 (.in(n14716_0), .out(n14716_1));
wire n14717; //CHANY 4 (9,2) #45
wire n14717_0;
wire n14717_1;
buffer_wire buffer_14717_1 (.in(n14717_0), .out(n14717_1));
wire n14718; //CHANY 4 (9,2) #52
wire n14718_0;
wire n14718_1;
buffer_wire buffer_14718_1 (.in(n14718_0), .out(n14718_1));
wire n14719; //CHANY 4 (9,2) #53
wire n14719_0;
wire n14719_1;
buffer_wire buffer_14719_1 (.in(n14719_0), .out(n14719_1));
wire n14720; //CHANY 4 (9,2) #60
wire n14720_0;
wire n14720_1;
buffer_wire buffer_14720_1 (.in(n14720_0), .out(n14720_1));
wire n14721; //CHANY 4 (9,2) #61
wire n14721_0;
wire n14721_1;
buffer_wire buffer_14721_1 (.in(n14721_0), .out(n14721_1));
wire n14722; //CHANY 4 (9,2) #68
wire n14722_0;
wire n14722_1;
buffer_wire buffer_14722_1 (.in(n14722_0), .out(n14722_1));
wire n14723; //CHANY 4 (9,2) #69
wire n14723_0;
wire n14723_1;
buffer_wire buffer_14723_1 (.in(n14723_0), .out(n14723_1));
wire n14724; //CHANY 4 (9,2) #76
wire n14724_0;
wire n14724_1;
buffer_wire buffer_14724_1 (.in(n14724_0), .out(n14724_1));
wire n14725; //CHANY 4 (9,2) #77
wire n14725_0;
wire n14725_1;
buffer_wire buffer_14725_1 (.in(n14725_0), .out(n14725_1));
wire n14726; //CHANY 8 (9,2) #84
wire n14726_0;
wire n14726_1;
wire n14726_2;
buffer_wire buffer_14726_2 (.in(n14726_1), .out(n14726_2));
buffer_wire buffer_14726_1 (.in(n14726_0), .out(n14726_1));
wire n14727; //CHANY 8 (9,2) #85
wire n14727_0;
wire n14727_1;
wire n14727_2;
buffer_wire buffer_14727_2 (.in(n14727_1), .out(n14727_2));
buffer_wire buffer_14727_1 (.in(n14727_0), .out(n14727_1));
wire n14728; //CHANY 4 (9,3) #6
wire n14728_0;
wire n14728_1;
buffer_wire buffer_14728_1 (.in(n14728_0), .out(n14728_1));
wire n14729; //CHANY 4 (9,3) #7
wire n14729_0;
wire n14729_1;
buffer_wire buffer_14729_1 (.in(n14729_0), .out(n14729_1));
wire n14730; //CHANY 4 (9,3) #14
wire n14730_0;
wire n14730_1;
buffer_wire buffer_14730_1 (.in(n14730_0), .out(n14730_1));
wire n14731; //CHANY 4 (9,3) #15
wire n14731_0;
wire n14731_1;
buffer_wire buffer_14731_1 (.in(n14731_0), .out(n14731_1));
wire n14732; //CHANY 4 (9,3) #22
wire n14732_0;
wire n14732_1;
buffer_wire buffer_14732_1 (.in(n14732_0), .out(n14732_1));
wire n14733; //CHANY 4 (9,3) #23
wire n14733_0;
wire n14733_1;
buffer_wire buffer_14733_1 (.in(n14733_0), .out(n14733_1));
wire n14734; //CHANY 4 (9,3) #30
wire n14734_0;
wire n14734_1;
buffer_wire buffer_14734_1 (.in(n14734_0), .out(n14734_1));
wire n14735; //CHANY 4 (9,3) #31
wire n14735_0;
wire n14735_1;
buffer_wire buffer_14735_1 (.in(n14735_0), .out(n14735_1));
wire n14736; //CHANY 4 (9,3) #38
wire n14736_0;
wire n14736_1;
buffer_wire buffer_14736_1 (.in(n14736_0), .out(n14736_1));
wire n14737; //CHANY 4 (9,3) #39
wire n14737_0;
wire n14737_1;
buffer_wire buffer_14737_1 (.in(n14737_0), .out(n14737_1));
wire n14738; //CHANY 4 (9,3) #46
wire n14738_0;
wire n14738_1;
buffer_wire buffer_14738_1 (.in(n14738_0), .out(n14738_1));
wire n14739; //CHANY 4 (9,3) #47
wire n14739_0;
wire n14739_1;
buffer_wire buffer_14739_1 (.in(n14739_0), .out(n14739_1));
wire n14740; //CHANY 4 (9,3) #54
wire n14740_0;
wire n14740_1;
buffer_wire buffer_14740_1 (.in(n14740_0), .out(n14740_1));
wire n14741; //CHANY 4 (9,3) #55
wire n14741_0;
wire n14741_1;
buffer_wire buffer_14741_1 (.in(n14741_0), .out(n14741_1));
wire n14742; //CHANY 4 (9,3) #62
wire n14742_0;
wire n14742_1;
buffer_wire buffer_14742_1 (.in(n14742_0), .out(n14742_1));
wire n14743; //CHANY 4 (9,3) #63
wire n14743_0;
wire n14743_1;
buffer_wire buffer_14743_1 (.in(n14743_0), .out(n14743_1));
wire n14744; //CHANY 4 (9,3) #70
wire n14744_0;
wire n14744_1;
buffer_wire buffer_14744_1 (.in(n14744_0), .out(n14744_1));
wire n14745; //CHANY 4 (9,3) #71
wire n14745_0;
wire n14745_1;
buffer_wire buffer_14745_1 (.in(n14745_0), .out(n14745_1));
wire n14746; //CHANY 4 (9,3) #78
wire n14746_0;
wire n14746_1;
buffer_wire buffer_14746_1 (.in(n14746_0), .out(n14746_1));
wire n14747; //CHANY 4 (9,3) #79
wire n14747_0;
wire n14747_1;
buffer_wire buffer_14747_1 (.in(n14747_0), .out(n14747_1));
wire n14748; //CHANY 7 (9,3) #86
wire n14748_0;
wire n14748_1;
wire n14748_2;
buffer_wire buffer_14748_2 (.in(n14748_1), .out(n14748_2));
buffer_wire buffer_14748_1 (.in(n14748_0), .out(n14748_1));
wire n14749; //CHANY 7 (9,3) #87
wire n14749_0;
wire n14749_1;
wire n14749_2;
buffer_wire buffer_14749_2 (.in(n14749_1), .out(n14749_2));
buffer_wire buffer_14749_1 (.in(n14749_0), .out(n14749_1));
wire n14750; //CHANY 4 (9,4) #0
wire n14750_0;
wire n14750_1;
buffer_wire buffer_14750_1 (.in(n14750_0), .out(n14750_1));
wire n14751; //CHANY 4 (9,4) #1
wire n14751_0;
wire n14751_1;
buffer_wire buffer_14751_1 (.in(n14751_0), .out(n14751_1));
wire n14752; //CHANY 4 (9,4) #8
wire n14752_0;
wire n14752_1;
buffer_wire buffer_14752_1 (.in(n14752_0), .out(n14752_1));
wire n14753; //CHANY 4 (9,4) #9
wire n14753_0;
wire n14753_1;
buffer_wire buffer_14753_1 (.in(n14753_0), .out(n14753_1));
wire n14754; //CHANY 4 (9,4) #16
wire n14754_0;
wire n14754_1;
buffer_wire buffer_14754_1 (.in(n14754_0), .out(n14754_1));
wire n14755; //CHANY 4 (9,4) #17
wire n14755_0;
wire n14755_1;
buffer_wire buffer_14755_1 (.in(n14755_0), .out(n14755_1));
wire n14756; //CHANY 4 (9,4) #24
wire n14756_0;
wire n14756_1;
buffer_wire buffer_14756_1 (.in(n14756_0), .out(n14756_1));
wire n14757; //CHANY 4 (9,4) #25
wire n14757_0;
wire n14757_1;
buffer_wire buffer_14757_1 (.in(n14757_0), .out(n14757_1));
wire n14758; //CHANY 4 (9,4) #32
wire n14758_0;
wire n14758_1;
buffer_wire buffer_14758_1 (.in(n14758_0), .out(n14758_1));
wire n14759; //CHANY 4 (9,4) #33
wire n14759_0;
wire n14759_1;
buffer_wire buffer_14759_1 (.in(n14759_0), .out(n14759_1));
wire n14760; //CHANY 4 (9,4) #40
wire n14760_0;
wire n14760_1;
buffer_wire buffer_14760_1 (.in(n14760_0), .out(n14760_1));
wire n14761; //CHANY 4 (9,4) #41
wire n14761_0;
wire n14761_1;
buffer_wire buffer_14761_1 (.in(n14761_0), .out(n14761_1));
wire n14762; //CHANY 4 (9,4) #48
wire n14762_0;
wire n14762_1;
buffer_wire buffer_14762_1 (.in(n14762_0), .out(n14762_1));
wire n14763; //CHANY 4 (9,4) #49
wire n14763_0;
wire n14763_1;
buffer_wire buffer_14763_1 (.in(n14763_0), .out(n14763_1));
wire n14764; //CHANY 4 (9,4) #56
wire n14764_0;
wire n14764_1;
buffer_wire buffer_14764_1 (.in(n14764_0), .out(n14764_1));
wire n14765; //CHANY 4 (9,4) #57
wire n14765_0;
wire n14765_1;
buffer_wire buffer_14765_1 (.in(n14765_0), .out(n14765_1));
wire n14766; //CHANY 4 (9,4) #64
wire n14766_0;
wire n14766_1;
buffer_wire buffer_14766_1 (.in(n14766_0), .out(n14766_1));
wire n14767; //CHANY 4 (9,4) #65
wire n14767_0;
wire n14767_1;
buffer_wire buffer_14767_1 (.in(n14767_0), .out(n14767_1));
wire n14768; //CHANY 4 (9,4) #72
wire n14768_0;
wire n14768_1;
buffer_wire buffer_14768_1 (.in(n14768_0), .out(n14768_1));
wire n14769; //CHANY 4 (9,4) #73
wire n14769_0;
wire n14769_1;
buffer_wire buffer_14769_1 (.in(n14769_0), .out(n14769_1));
wire n14770; //CHANY 6 (9,4) #88
wire n14770_0;
wire n14770_1;
buffer_wire buffer_14770_1 (.in(n14770_0), .out(n14770_1));
wire n14771; //CHANY 6 (9,4) #89
wire n14771_0;
wire n14771_1;
buffer_wire buffer_14771_1 (.in(n14771_0), .out(n14771_1));
wire n14772; //CHANY 4 (9,5) #2
wire n14772_0;
wire n14772_1;
buffer_wire buffer_14772_1 (.in(n14772_0), .out(n14772_1));
wire n14773; //CHANY 4 (9,5) #3
wire n14773_0;
wire n14773_1;
buffer_wire buffer_14773_1 (.in(n14773_0), .out(n14773_1));
wire n14774; //CHANY 4 (9,5) #10
wire n14774_0;
wire n14774_1;
buffer_wire buffer_14774_1 (.in(n14774_0), .out(n14774_1));
wire n14775; //CHANY 4 (9,5) #11
wire n14775_0;
wire n14775_1;
buffer_wire buffer_14775_1 (.in(n14775_0), .out(n14775_1));
wire n14776; //CHANY 4 (9,5) #18
wire n14776_0;
wire n14776_1;
buffer_wire buffer_14776_1 (.in(n14776_0), .out(n14776_1));
wire n14777; //CHANY 4 (9,5) #19
wire n14777_0;
wire n14777_1;
buffer_wire buffer_14777_1 (.in(n14777_0), .out(n14777_1));
wire n14778; //CHANY 4 (9,5) #26
wire n14778_0;
wire n14778_1;
buffer_wire buffer_14778_1 (.in(n14778_0), .out(n14778_1));
wire n14779; //CHANY 4 (9,5) #27
wire n14779_0;
wire n14779_1;
buffer_wire buffer_14779_1 (.in(n14779_0), .out(n14779_1));
wire n14780; //CHANY 4 (9,5) #34
wire n14780_0;
wire n14780_1;
buffer_wire buffer_14780_1 (.in(n14780_0), .out(n14780_1));
wire n14781; //CHANY 4 (9,5) #35
wire n14781_0;
wire n14781_1;
buffer_wire buffer_14781_1 (.in(n14781_0), .out(n14781_1));
wire n14782; //CHANY 4 (9,5) #42
wire n14782_0;
wire n14782_1;
buffer_wire buffer_14782_1 (.in(n14782_0), .out(n14782_1));
wire n14783; //CHANY 4 (9,5) #43
wire n14783_0;
wire n14783_1;
buffer_wire buffer_14783_1 (.in(n14783_0), .out(n14783_1));
wire n14784; //CHANY 4 (9,5) #50
wire n14784_0;
wire n14784_1;
buffer_wire buffer_14784_1 (.in(n14784_0), .out(n14784_1));
wire n14785; //CHANY 4 (9,5) #51
wire n14785_0;
wire n14785_1;
buffer_wire buffer_14785_1 (.in(n14785_0), .out(n14785_1));
wire n14786; //CHANY 4 (9,5) #58
wire n14786_0;
wire n14786_1;
buffer_wire buffer_14786_1 (.in(n14786_0), .out(n14786_1));
wire n14787; //CHANY 4 (9,5) #59
wire n14787_0;
wire n14787_1;
buffer_wire buffer_14787_1 (.in(n14787_0), .out(n14787_1));
wire n14788; //CHANY 4 (9,5) #66
wire n14788_0;
wire n14788_1;
buffer_wire buffer_14788_1 (.in(n14788_0), .out(n14788_1));
wire n14789; //CHANY 4 (9,5) #67
wire n14789_0;
wire n14789_1;
buffer_wire buffer_14789_1 (.in(n14789_0), .out(n14789_1));
wire n14790; //CHANY 4 (9,5) #74
wire n14790_0;
wire n14790_1;
buffer_wire buffer_14790_1 (.in(n14790_0), .out(n14790_1));
wire n14791; //CHANY 4 (9,5) #75
wire n14791_0;
wire n14791_1;
buffer_wire buffer_14791_1 (.in(n14791_0), .out(n14791_1));
wire n14792; //CHANY 5 (9,5) #90
wire n14792_0;
wire n14792_1;
buffer_wire buffer_14792_1 (.in(n14792_0), .out(n14792_1));
wire n14793; //CHANY 5 (9,5) #91
wire n14793_0;
wire n14793_1;
buffer_wire buffer_14793_1 (.in(n14793_0), .out(n14793_1));
wire n14794; //CHANY 4 (9,6) #4
wire n14794_0;
wire n14794_1;
buffer_wire buffer_14794_1 (.in(n14794_0), .out(n14794_1));
wire n14795; //CHANY 4 (9,6) #5
wire n14795_0;
wire n14795_1;
buffer_wire buffer_14795_1 (.in(n14795_0), .out(n14795_1));
wire n14796; //CHANY 4 (9,6) #12
wire n14796_0;
wire n14796_1;
buffer_wire buffer_14796_1 (.in(n14796_0), .out(n14796_1));
wire n14797; //CHANY 4 (9,6) #13
wire n14797_0;
wire n14797_1;
buffer_wire buffer_14797_1 (.in(n14797_0), .out(n14797_1));
wire n14798; //CHANY 4 (9,6) #20
wire n14798_0;
wire n14798_1;
buffer_wire buffer_14798_1 (.in(n14798_0), .out(n14798_1));
wire n14799; //CHANY 4 (9,6) #21
wire n14799_0;
wire n14799_1;
buffer_wire buffer_14799_1 (.in(n14799_0), .out(n14799_1));
wire n14800; //CHANY 4 (9,6) #28
wire n14800_0;
wire n14800_1;
buffer_wire buffer_14800_1 (.in(n14800_0), .out(n14800_1));
wire n14801; //CHANY 4 (9,6) #29
wire n14801_0;
wire n14801_1;
buffer_wire buffer_14801_1 (.in(n14801_0), .out(n14801_1));
wire n14802; //CHANY 4 (9,6) #36
wire n14802_0;
wire n14802_1;
buffer_wire buffer_14802_1 (.in(n14802_0), .out(n14802_1));
wire n14803; //CHANY 4 (9,6) #37
wire n14803_0;
wire n14803_1;
buffer_wire buffer_14803_1 (.in(n14803_0), .out(n14803_1));
wire n14804; //CHANY 4 (9,6) #44
wire n14804_0;
wire n14804_1;
buffer_wire buffer_14804_1 (.in(n14804_0), .out(n14804_1));
wire n14805; //CHANY 4 (9,6) #45
wire n14805_0;
wire n14805_1;
buffer_wire buffer_14805_1 (.in(n14805_0), .out(n14805_1));
wire n14806; //CHANY 4 (9,6) #52
wire n14806_0;
wire n14806_1;
buffer_wire buffer_14806_1 (.in(n14806_0), .out(n14806_1));
wire n14807; //CHANY 4 (9,6) #53
wire n14807_0;
wire n14807_1;
buffer_wire buffer_14807_1 (.in(n14807_0), .out(n14807_1));
wire n14808; //CHANY 4 (9,6) #60
wire n14808_0;
wire n14808_1;
buffer_wire buffer_14808_1 (.in(n14808_0), .out(n14808_1));
wire n14809; //CHANY 4 (9,6) #61
wire n14809_0;
wire n14809_1;
buffer_wire buffer_14809_1 (.in(n14809_0), .out(n14809_1));
wire n14810; //CHANY 4 (9,6) #68
wire n14810_0;
wire n14810_1;
buffer_wire buffer_14810_1 (.in(n14810_0), .out(n14810_1));
wire n14811; //CHANY 4 (9,6) #69
wire n14811_0;
wire n14811_1;
buffer_wire buffer_14811_1 (.in(n14811_0), .out(n14811_1));
wire n14812; //CHANY 4 (9,6) #76
wire n14812_0;
wire n14812_1;
buffer_wire buffer_14812_1 (.in(n14812_0), .out(n14812_1));
wire n14813; //CHANY 4 (9,6) #77
wire n14813_0;
wire n14813_1;
buffer_wire buffer_14813_1 (.in(n14813_0), .out(n14813_1));
wire n14814; //CHANY 3 (9,7) #6
wire n14814_0;
wire n14815; //CHANY 3 (9,7) #7
wire n14815_0;
wire n14816; //CHANY 3 (9,7) #14
wire n14816_0;
wire n14817; //CHANY 3 (9,7) #15
wire n14817_0;
wire n14818; //CHANY 3 (9,7) #22
wire n14818_0;
wire n14819; //CHANY 3 (9,7) #23
wire n14819_0;
wire n14820; //CHANY 3 (9,7) #30
wire n14820_0;
wire n14821; //CHANY 3 (9,7) #31
wire n14821_0;
wire n14822; //CHANY 3 (9,7) #38
wire n14822_0;
wire n14823; //CHANY 3 (9,7) #39
wire n14823_0;
wire n14824; //CHANY 3 (9,7) #46
wire n14824_0;
wire n14825; //CHANY 3 (9,7) #47
wire n14825_0;
wire n14826; //CHANY 3 (9,7) #54
wire n14826_0;
wire n14827; //CHANY 3 (9,7) #55
wire n14827_0;
wire n14828; //CHANY 3 (9,7) #62
wire n14828_0;
wire n14829; //CHANY 3 (9,7) #63
wire n14829_0;
wire n14830; //CHANY 3 (9,7) #70
wire n14830_0;
wire n14831; //CHANY 3 (9,7) #71
wire n14831_0;
wire n14832; //CHANY 3 (9,7) #78
wire n14832_0;
wire n14833; //CHANY 3 (9,7) #79
wire n14833_0;
wire n14834; //CHANY 2 (9,8) #0
wire n14834_0;
wire n14835; //CHANY 2 (9,8) #1
wire n14835_0;
wire n14836; //CHANY 2 (9,8) #8
wire n14836_0;
wire n14837; //CHANY 2 (9,8) #9
wire n14837_0;
wire n14838; //CHANY 2 (9,8) #16
wire n14838_0;
wire n14839; //CHANY 2 (9,8) #17
wire n14839_0;
wire n14840; //CHANY 2 (9,8) #24
wire n14840_0;
wire n14841; //CHANY 2 (9,8) #25
wire n14841_0;
wire n14842; //CHANY 2 (9,8) #32
wire n14842_0;
wire n14843; //CHANY 2 (9,8) #33
wire n14843_0;
wire n14844; //CHANY 2 (9,8) #40
wire n14844_0;
wire n14845; //CHANY 2 (9,8) #41
wire n14845_0;
wire n14846; //CHANY 2 (9,8) #48
wire n14846_0;
wire n14847; //CHANY 2 (9,8) #49
wire n14847_0;
wire n14848; //CHANY 2 (9,8) #56
wire n14848_0;
wire n14849; //CHANY 2 (9,8) #57
wire n14849_0;
wire n14850; //CHANY 2 (9,8) #64
wire n14850_0;
wire n14851; //CHANY 2 (9,8) #65
wire n14851_0;
wire n14852; //CHANY 2 (9,8) #72
wire n14852_0;
wire n14853; //CHANY 2 (9,8) #73
wire n14853_0;
wire n14854; //CHANY 1 (9,9) #2
wire n14854_0;
wire n14855; //CHANY 1 (9,9) #3
wire n14855_0;
wire n14856; //CHANY 1 (9,9) #10
wire n14856_0;
wire n14857; //CHANY 1 (9,9) #11
wire n14857_0;
wire n14858; //CHANY 1 (9,9) #18
wire n14858_0;
wire n14859; //CHANY 1 (9,9) #19
wire n14859_0;
wire n14860; //CHANY 1 (9,9) #26
wire n14860_0;
wire n14861; //CHANY 1 (9,9) #27
wire n14861_0;
wire n14862; //CHANY 1 (9,9) #34
wire n14862_0;
wire n14863; //CHANY 1 (9,9) #35
wire n14863_0;
wire n14864; //CHANY 1 (9,9) #42
wire n14864_0;
wire n14865; //CHANY 1 (9,9) #43
wire n14865_0;
wire n14866; //CHANY 1 (9,9) #50
wire n14866_0;
wire n14867; //CHANY 1 (9,9) #51
wire n14867_0;
wire n14868; //CHANY 1 (9,9) #58
wire n14868_0;
wire n14869; //CHANY 1 (9,9) #59
wire n14869_0;
wire n14870; //CHANY 1 (9,9) #66
wire n14870_0;
wire n14871; //CHANY 1 (9,9) #67
wire n14871_0;
wire n14872; //CHANY 1 (9,9) #74
wire n14872_0;
wire n14873; //CHANY 1 (9,9) #75
wire n14873_0;
wire [`CONFIG_SIZE-1:0] config_chain;

mux6 mux_0 (.in({n12333_0, n12332_0, n12301_0, n12300_0, n12271_1, n12270_0}), .out(n24), .config_in(config_chain[2:0]), .config_rst(config_rst)); 
mux6 mux_1 (.in({n12337_0, n12336_0, n12305_0, n12304_0, n12275_0, n12274_0}), .out(n27), .config_in(config_chain[5:3]), .config_rst(config_rst)); 
mux6 mux_2 (.in({n12339_0, n12338_0, n12309_0, n12308_0, n12279_1, n12278_0}), .out(n30), .config_in(config_chain[8:6]), .config_rst(config_rst)); 
mux6 mux_3 (.in({n12343_1, n12342_0, n12313_0, n12312_0, n12283_0, n12282_0}), .out(n33), .config_in(config_chain[11:9]), .config_rst(config_rst)); 
mux6 mux_4 (.in({n12347_0, n12346_0, n12317_0, n12316_0, n12287_1, n12286_0}), .out(n36), .config_in(config_chain[14:12]), .config_rst(config_rst)); 
mux6 mux_5 (.in({n12351_2, n12350_0, n12321_0, n12320_0, n12291_0, n12290_0}), .out(n39), .config_in(config_chain[17:15]), .config_rst(config_rst)); 
mux6 mux_6 (.in({n12355_2, n12354_0, n12325_0, n12324_0, n12293_0, n12292_0}), .out(n42), .config_in(config_chain[20:18]), .config_rst(config_rst)); 
mux6 mux_7 (.in({n12359_2, n12358_0, n12329_0, n12328_0, n12297_0, n12296_0}), .out(n45), .config_in(config_chain[23:21]), .config_rst(config_rst)); 
mux6 mux_8 (.in({n12331_0, n12330_0, n12299_0, n12298_0, n12277_0, n12276_0}), .out(n72), .config_in(config_chain[26:24]), .config_rst(config_rst)); 
mux6 mux_9 (.in({n12363_1, n12362_0, n12335_0, n12334_0, n12303_0, n12302_0}), .out(n75), .config_in(config_chain[29:27]), .config_rst(config_rst)); 
mux6 mux_10 (.in({n12379_1, n12378_0, n12307_0, n12306_0, n12285_0, n12284_0}), .out(n78), .config_in(config_chain[32:30]), .config_rst(config_rst)); 
mux6 mux_11 (.in({n12365_1, n12364_0, n12349_0, n12348_0, n12311_0, n12310_0}), .out(n81), .config_in(config_chain[35:33]), .config_rst(config_rst)); 
mux6 mux_12 (.in({n12381_1, n12380_0, n12315_0, n12314_0, n12293_0, n12292_0}), .out(n84), .config_in(config_chain[38:36]), .config_rst(config_rst)); 
mux6 mux_13 (.in({n12367_1, n12366_0, n12361_2, n12360_0, n12319_0, n12318_0}), .out(n87), .config_in(config_chain[41:39]), .config_rst(config_rst)); 
mux6 mux_14 (.in({n12353_2, n12352_0, n12323_0, n12322_0, n12291_0, n12290_0}), .out(n90), .config_in(config_chain[44:42]), .config_rst(config_rst)); 
mux6 mux_15 (.in({n12357_2, n12356_0, n12327_0, n12326_0, n12295_0, n12294_0}), .out(n93), .config_in(config_chain[47:45]), .config_rst(config_rst)); 
mux6 mux_16 (.in({n12383_1, n12382_0, n12377_0, n12376_0, n12369_0, n12368_0}), .out(n120), .config_in(config_chain[50:48]), .config_rst(config_rst)); 
mux6 mux_17 (.in({n12341_0, n12340_0, n12309_0, n12308_0, n12271_0, n12270_0}), .out(n123), .config_in(config_chain[53:51]), .config_rst(config_rst)); 
mux6 mux_18 (.in({n12385_1, n12384_0, n12371_0, n12370_0, n12335_0, n12334_0}), .out(n126), .config_in(config_chain[56:54]), .config_rst(config_rst)); 
mux6 mux_19 (.in({n12401_1, n12400_0, n12317_0, n12316_0, n12279_0, n12278_0}), .out(n129), .config_in(config_chain[59:57]), .config_rst(config_rst)); 
mux6 mux_20 (.in({n12387_1, n12386_0, n12373_0, n12372_0, n12343_0, n12342_0}), .out(n132), .config_in(config_chain[62:60]), .config_rst(config_rst)); 
mux6 mux_21 (.in({n12359_2, n12358_0, n12325_0, n12324_0, n12287_0, n12286_0}), .out(n135), .config_in(config_chain[65:63]), .config_rst(config_rst)); 
mux6 mux_22 (.in({n12375_0, n12374_0, n12367_0, n12366_0, n12351_1, n12350_0}), .out(n138), .config_in(config_chain[68:66]), .config_rst(config_rst)); 
mux6 mux_23 (.in({n12355_2, n12354_0, n12333_0, n12332_0, n12301_0, n12300_0}), .out(n141), .config_in(config_chain[71:69]), .config_rst(config_rst)); 
mux6 mux_24 (.in({n12363_0, n12362_0, n12327_0, n12326_1, n12295_0, n12294_1}), .out(n168), .config_in(config_chain[74:72]), .config_rst(config_rst)); 
mux6 mux_25 (.in({n12403_1, n12402_0, n12399_0, n12398_0, n12391_0, n12390_0}), .out(n171), .config_in(config_chain[77:75]), .config_rst(config_rst)); 
mux6 mux_26 (.in({n12419_1, n12418_0, n12365_0, n12364_0, n12303_0, n12302_1}), .out(n174), .config_in(config_chain[80:78]), .config_rst(config_rst)); 
mux6 mux_27 (.in({n12405_1, n12404_0, n12393_0, n12392_0, n12381_0, n12380_0}), .out(n177), .config_in(config_chain[83:81]), .config_rst(config_rst)); 
mux6 mux_28 (.in({n12421_1, n12420_0, n12367_0, n12366_0, n12311_0, n12310_1}), .out(n180), .config_in(config_chain[86:84]), .config_rst(config_rst)); 
mux6 mux_29 (.in({n12407_1, n12406_0, n12395_0, n12394_0, n12357_1, n12356_1}), .out(n183), .config_in(config_chain[89:87]), .config_rst(config_rst)); 
mux6 mux_30 (.in({n12361_1, n12360_1, n12319_0, n12318_1, n12287_0, n12286_1}), .out(n186), .config_in(config_chain[92:90]), .config_rst(config_rst)); 
mux6 mux_31 (.in({n12397_0, n12396_0, n12389_0, n12388_0, n12353_1, n12352_1}), .out(n189), .config_in(config_chain[95:93]), .config_rst(config_rst)); 
mux6 mux_32 (.in({n12423_1/**/, n12422_0, n12417_0, n12416_0, n12409_0, n12408_0}), .out(n216), .config_in(config_chain[98:96]), .config_rst(config_rst)); 
mux6 mux_33 (.in({n12383_0, n12382_0, n12379_0, n12378_1, n12371_0, n12370_1}), .out(n219), .config_in(config_chain[101:99]), .config_rst(config_rst)); 
mux6 mux_34 (.in({n12425_1, n12424_0, n12411_0, n12410_0, n12399_0, n12398_0}), .out(n222), .config_in(config_chain[104:102]), .config_rst(config_rst)); 
mux6 mux_35 (.in({n12441_1, n12440_0, n12385_0, n12384_0, n12373_0, n12372_1}), .out(n225), .config_in(config_chain[107:105]), .config_rst(config_rst)); 
mux6 mux_36 (.in({n12427_1, n12426_0, n12413_0, n12412_0, n12401_0, n12400_0}), .out(n228), .config_in(config_chain[110:108]), .config_rst(config_rst)); 
mux6 mux_37 (.in({n12387_0, n12386_0, n12375_0, n12374_1, n12355_1, n12354_1}), .out(n231), .config_in(config_chain[113:111]), .config_rst(config_rst)); 
mux6 mux_38 (.in({n12415_0, n12414_0, n12407_0, n12406_0, n12359_1, n12358_1}), .out(n234), .config_in(config_chain[116:114]), .config_rst(config_rst)); 
mux6 mux_39 (.in({n12377_0, n12376_1, n12369_0, n12368_1, n12351_1, n12350_1}), .out(n237), .config_in(config_chain[119:117]), .config_rst(config_rst)); 
mux6 mux_40 (.in({n12403_0, n12402_0, n12397_0, n12396_1, n12389_0, n12388_1}), .out(n264), .config_in(config_chain[122:120]), .config_rst(config_rst)); 
mux6 mux_41 (.in({n12443_1, n12442_0, n12439_0, n12438_0, n12431_0, n12430_0}), .out(n267), .config_in(config_chain[125:123]), .config_rst(config_rst)); 
mux6 mux_42 (.in({n12459_1, n12458_0, n12405_0, n12404_0, n12391_0, n12390_1}), .out(n270), .config_in(config_chain[128:126]), .config_rst(config_rst)); 
mux6 mux_43 (.in({n12445_1, n12444_0, n12433_0, n12432_0, n12421_0, n12420_0}), .out(n273), .config_in(config_chain[131:129]), .config_rst(config_rst)); 
mux6 mux_44 (.in({n12461_1, n12460_0, n12407_0, n12406_0, n12393_0, n12392_1}), .out(n276), .config_in(config_chain[134:132]), .config_rst(config_rst)); 
mux6 mux_45 (.in({n12447_1, n12446_0, n12435_0, n12434_0, n12353_1, n12352_1}), .out(n279), .config_in(config_chain[137:135]), .config_rst(config_rst)); 
mux6 mux_46 (.in({n12395_0, n12394_1, n12387_0, n12386_1, n12357_1, n12356_1}), .out(n282), .config_in(config_chain[140:138]), .config_rst(config_rst)); 
mux6 mux_47 (.in({n12437_0, n12436_0, n12429_0, n12428_0, n12361_1, n12360_1}), .out(n285), .config_in(config_chain[143:141]), .config_rst(config_rst)); 
mux6 mux_48 (.in({n12463_0, n12462_0, n12457_0, n12456_0, n12449_0, n12448_0}), .out(n312), .config_in(config_chain[146:144]), .config_rst(config_rst)); 
mux6 mux_49 (.in({n12423_0, n12422_0, n12419_0, n12418_1, n12411_0, n12410_1}), .out(n315), .config_in(config_chain[149:147]), .config_rst(config_rst)); 
mux6 mux_50 (.in({n12465_0, n12464_0, n12451_0, n12450_0, n12439_0, n12438_0}), .out(n318), .config_in(config_chain[152:150]), .config_rst(config_rst)); 
mux6 mux_51 (.in({n12481_0, n12480_0, n12425_0, n12424_0, n12413_0, n12412_1}), .out(n321), .config_in(config_chain[155:153]), .config_rst(config_rst)); 
mux6 mux_52 (.in({n12467_0, n12466_0, n12453_0, n12452_0, n12441_0, n12440_0}), .out(n324), .config_in(config_chain[158:156]), .config_rst(config_rst)); 
mux6 mux_53 (.in({n12427_0, n12426_0, n12415_0, n12414_1, n12351_0, n12350_2}), .out(n327), .config_in(config_chain[161:159]), .config_rst(config_rst)); 
mux6 mux_54 (.in({n12455_0, n12454_0, n12447_0, n12446_0, n12355_0, n12354_2}), .out(n330), .config_in(config_chain[164:162]), .config_rst(config_rst)); 
mux6 mux_55 (.in({n12417_0, n12416_1, n12409_0, n12408_1, n12359_0, n12358_2}), .out(n333), .config_in(config_chain[167:165]), .config_rst(config_rst)); 
mux6 mux_56 (.in({n12443_0, n12442_0, n12437_0, n12436_1, n12429_0, n12428_1}), .out(n360), .config_in(config_chain[170:168]), .config_rst(config_rst)); 
mux6 mux_57 (.in({n12483_0, n12482_0, n12479_0, n12478_0, n12471_0, n12470_0}), .out(n363), .config_in(config_chain[173:171]), .config_rst(config_rst)); 
mux6 mux_58 (.in({n12499_0, n12498_0, n12445_0, n12444_0, n12431_0, n12430_1}), .out(n366), .config_in(config_chain[176:174]), .config_rst(config_rst)); 
mux6 mux_59 (.in({n12485_0, n12484_0, n12473_0, n12472_0, n12461_0, n12460_0}), .out(n369), .config_in(config_chain[179:177]), .config_rst(config_rst)); 
mux6 mux_60 (.in({n12501_0, n12500_0, n12447_0, n12446_0, n12433_0, n12432_1}), .out(n372), .config_in(config_chain[182:180]), .config_rst(config_rst)); 
mux6 mux_61 (.in({n12487_0, n12486_0, n12475_0, n12474_0, n12361_0, n12360_2}), .out(n375), .config_in(config_chain[185:183]), .config_rst(config_rst)); 
mux6 mux_62 (.in({n12435_0, n12434_1, n12427_0, n12426_1, n12353_0, n12352_2}), .out(n378), .config_in(config_chain[188:186]), .config_rst(config_rst)); 
mux6 mux_63 (.in({n12477_0, n12476_0, n12469_0, n12468_0, n12357_0, n12356_2}), .out(n381), .config_in(config_chain[191:189]), .config_rst(config_rst)); 
mux6 mux_64 (.in({n12503_0, n12502_0, n12497_0, n12496_0, n12489_0, n12488_0}), .out(n408), .config_in(config_chain[194:192]), .config_rst(config_rst)); 
mux6 mux_65 (.in({n12463_0, n12462_0, n12459_0, n12458_1, n12451_0, n12450_1}), .out(n411), .config_in(config_chain[197:195]), .config_rst(config_rst)); 
mux6 mux_66 (.in({n12505_0, n12504_0, n12491_0, n12490_0, n12479_0, n12478_0}), .out(n414), .config_in(config_chain[200:198]), .config_rst(config_rst)); 
mux6 mux_67 (.in({n12521_0, n12520_0, n12465_0, n12464_0, n12453_0, n12452_1}), .out(n417), .config_in(config_chain[203:201]), .config_rst(config_rst)); 
mux6 mux_68 (.in({n12507_0, n12506_0, n12493_0, n12492_0, n12481_0, n12480_0}), .out(n420), .config_in(config_chain[206:204]), .config_rst(config_rst)); 
mux6 mux_69 (.in({n12467_0, n12466_0, n12455_0, n12454_1, n12359_0, n12358_2}), .out(n423), .config_in(config_chain[209:207]), .config_rst(config_rst)); 
mux6 mux_70 (.in({n12523_0, n12522_0, n12495_0, n12494_0, n12487_0, n12486_0}), .out(n426), .config_in(config_chain[212:210]), .config_rst(config_rst)); 
mux6 mux_71 (.in({n12457_0, n12456_1, n12449_0, n12448_1, n12355_0, n12354_2}), .out(n429), .config_in(config_chain[215:213]), .config_rst(config_rst)); 
mux6 mux_72 (.in({n9727_0, n9726_0, n9697_0, n9696_0, n9667_1, n9666_0}), .out(n456), .config_in(config_chain[218:216]), .config_rst(config_rst)); 
mux6 mux_73 (.in({n9731_1, n9730_0, n9701_0, n9700_0, n9669_0, n9668_0}), .out(n459), .config_in(config_chain[221:219]), .config_rst(config_rst)); 
mux6 mux_74 (.in({n9735_0, n9734_0, n9705_0, n9704_0, n9673_0, n9672_0}), .out(n462), .config_in(config_chain[224:222]), .config_rst(config_rst)); 
mux6 mux_75 (.in({n9739_1, n9738_0, n9709_0, n9708_0, n9677_0, n9676_0}), .out(n465), .config_in(config_chain[227:225]), .config_rst(config_rst)); 
mux6 mux_76 (.in({n9743_0, n9742_0, n9713_0, n9712_0, n9681_0, n9680_0}), .out(n468), .config_in(config_chain[230:228]), .config_rst(config_rst)); 
mux6 mux_77 (.in({n9747_2, n9746_0, n9715_1, n9714_0, n9685_0, n9684_0}), .out(n471), .config_in(config_chain[233:231]), .config_rst(config_rst)); 
mux6 mux_78 (.in({n9751_2, n9750_0, n9719_0, n9718_0, n9689_0, n9688_0}), .out(n474), .config_in(config_chain[236:234]), .config_rst(config_rst)); 
mux6 mux_79 (.in({n9755_2, n9754_0, n9723_1, n9722_0, n9693_0, n9692_0}), .out(n477), .config_in(config_chain[239:237]), .config_rst(config_rst)); 
mux6 mux_80 (.in({n9979_1, n9978_0, n9949_0, n9948_0, n9927_0, n9926_0}), .out(n505), .config_in(config_chain[242:240]), .config_rst(config_rst)); 
mux6 mux_81 (.in({n12583_1, n12582_0, n12553_0, n12552_0, n12531_0, n12530_0}), .out(n506), .config_in(config_chain[245:243]), .config_rst(config_rst)); 
mux6 mux_82 (.in({n9729_0, n9728_0, n9697_0, n9696_0, n9667_1, n9666_0}), .out(n507), .config_in(config_chain[248:246]), .config_rst(config_rst)); 
mux6 mux_83 (.in({n12333_0, n12332_0, n12303_1, n12302_0, n12271_1, n12270_0}), .out(n508), .config_in(config_chain[251:249]), .config_rst(config_rst)); 
mux6 mux_84 (.in({n9981_0, n9980_0, n9959_0, n9958_0, n9921_0, n9920_0}), .out(n509), .config_in(config_chain[254:252]), .config_rst(config_rst)); 
mux6 mux_85 (.in({n12595_0, n12594_0, n12563_0, n12562_0, n12525_0, n12524_0}), .out(n510), .config_in(config_chain[257:255]), .config_rst(config_rst)); 
mux6 mux_86 (.in({n9731_1, n9730_0, n9701_0, n9700_0, n9669_0, n9668_0}), .out(n511), .config_in(config_chain[260:258]), .config_rst(config_rst)); 
mux6 mux_87 (.in({n12335_1, n12334_0, n12305_0, n12304_0, n12275_0, n12274_0}), .out(n512), .config_in(config_chain[263:261]), .config_rst(config_rst)); 
mux6 mux_88 (.in({n9985_0, n9984_0, n9953_0, n9952_0, n9923_1, n9922_0}), .out(n513), .config_in(config_chain[266:264]), .config_rst(config_rst)); 
mux6 mux_89 (.in({n12589_0, n12588_0, n12557_0, n12556_0, n12527_1, n12526_0}), .out(n514), .config_in(config_chain[269:267]), .config_rst(config_rst)); 
mux6 mux_90 (.in({n9733_0, n9732_0, n9703_0, n9702_0, n9671_0, n9670_0}), .out(n515), .config_in(config_chain[272:270]), .config_rst(config_rst)); 
mux6 mux_91 (.in({n12337_0, n12336_0, n12307_0, n12306_0, n12277_0, n12276_0}), .out(n516), .config_in(config_chain[275:273]), .config_rst(config_rst)); 
mux6 mux_92 (.in({n9987_1, n9986_0, n9955_1, n9954_0, n9925_0, n9924_0}), .out(n517), .config_in(config_chain[278:276]), .config_rst(config_rst)); 
mux6 mux_93 (.in({n12591_1, n12590_0, n12561_0, n12560_0, n12529_0, n12528_0}), .out(n518), .config_in(config_chain[281:279]), .config_rst(config_rst)); 
mux6 mux_94 (.in({n9735_0, n9734_0, n9705_0, n9704_0, n9675_1, n9674_0}), .out(n519), .config_in(config_chain[284:282]), .config_rst(config_rst)); 
mux6 mux_95 (.in({n12341_0, n12340_0, n12309_0, n12308_0, n12279_1, n12278_0}), .out(n520), .config_in(config_chain[287:285]), .config_rst(config_rst)); 
mux6 mux_96 (.in({n9989_0, n9988_0, n9967_0, n9966_0, n9935_0, n9934_0}), .out(n521), .config_in(config_chain[290:288]), .config_rst(config_rst)); 
mux6 mux_97 (.in({n12593_0, n12592_0, n12571_0, n12570_0, n12533_0, n12532_0}), .out(n522), .config_in(config_chain[293:291]), .config_rst(config_rst)); 
mux6 mux_98 (.in({n9737_0, n9736_0, n9707_1, n9706_0, n9677_0, n9676_0}), .out(n523), .config_in(config_chain[296:294]), .config_rst(config_rst)); 
mux6 mux_99 (.in({n12343_1, n12342_0, n12311_1, n12310_0, n12281_0, n12280_0}), .out(n524), .config_in(config_chain[299:297]), .config_rst(config_rst)); 
mux6 mux_100 (.in({n9999_0, n9998_0, n9961_0, n9960_0, n9929_0, n9928_0}), .out(n525), .config_in(config_chain[302:300]), .config_rst(config_rst)); 
mux6 mux_101 (.in({n12603_0, n12602_0, n12565_0, n12564_0, n12535_1, n12534_0}), .out(n526), .config_in(config_chain[305:303]), .config_rst(config_rst)); 
mux6 mux_102 (.in({n9741_0, n9740_0, n9709_0, n9708_0, n9679_0, n9678_0}), .out(n527), .config_in(config_chain[308:306]), .config_rst(config_rst)); 
mux6 mux_103 (.in({n12345_0, n12344_0, n12315_0, n12314_0, n12283_0, n12282_0}), .out(n528), .config_in(config_chain[311:309]), .config_rst(config_rst)); 
mux6 mux_104 (.in({n9993_0, n9992_0, n9963_1, n9962_0, n9933_0, n9932_0}), .out(n529), .config_in(config_chain[314:312]), .config_rst(config_rst)); 
mux6 mux_105 (.in({n12599_1, n12598_0, n12567_1, n12566_0, n12537_0, n12536_0}), .out(n530), .config_in(config_chain[317:315]), .config_rst(config_rst)); 
mux6 mux_106 (.in({n9743_0, n9742_0, n9713_0, n9712_0, n9681_0, n9680_0}), .out(n531), .config_in(config_chain[320:318]), .config_rst(config_rst)); 
mux6 mux_107 (.in({n12347_0, n12346_0, n12317_0, n12316_0, n12285_0, n12284_0}), .out(n532), .config_in(config_chain[323:321]), .config_rst(config_rst)); 
mux6 mux_108 (.in({n9995_1, n9994_0, n9965_0, n9964_0, n9943_0, n9942_0}), .out(n533), .config_in(config_chain[326:324]), .config_rst(config_rst)); 
mux6 mux_109 (.in({n12601_0, n12600_0, n12569_0, n12568_0, n12547_0, n12546_0}), .out(n534), .config_in(config_chain[329:327]), .config_rst(config_rst)); 
mux6 mux_110 (.in({n9745_0, n9744_0, n9715_1, n9714_0, n9683_1, n9682_0}), .out(n535), .config_in(config_chain[332:330]), .config_rst(config_rst)); 
mux6 mux_111 (.in({n12349_0, n12348_0, n12319_1, n12318_0, n12289_0, n12288_0}), .out(n536), .config_in(config_chain[335:333]), .config_rst(config_rst)); 
mux6 mux_112 (.in({n10011_2, n10010_0, n9975_0, n9974_0, n9937_0, n9936_0}), .out(n537), .config_in(config_chain[338:336]), .config_rst(config_rst)); 
mux6 mux_113 (.in({n12615_2, n12614_0, n12573_0, n12572_0, n12541_0, n12540_0}), .out(n538), .config_in(config_chain[341:339]), .config_rst(config_rst)); 
mux6 mux_114 (.in({n9747_2, n9746_0, n9717_0, n9716_0, n9687_0, n9686_0}), .out(n539), .config_in(config_chain[344:342]), .config_rst(config_rst)); 
mux6 mux_115 (.in({n12351_2, n12350_0, n12321_0, n12320_0, n12291_0, n12290_0}), .out(n540), .config_in(config_chain[347:345]), .config_rst(config_rst)); 
mux6 mux_116 (.in({n10001_2, n10000_0, n9969_0, n9968_0, n9939_1, n9938_0}), .out(n541), .config_in(config_chain[350:348]), .config_rst(config_rst)); 
mux6 mux_117 (.in({n12605_2, n12604_0, n12575_1, n12574_0, n12543_1, n12542_0}), .out(n542), .config_in(config_chain[353:351]), .config_rst(config_rst)); 
mux6 mux_118 (.in({n9749_2, n9748_0, n9719_0, n9718_0, n9689_0, n9688_0}), .out(n543), .config_in(config_chain[356:354]), .config_rst(config_rst)); 
mux6 mux_119 (.in({n12355_2, n12354_0, n12323_0, n12322_0, n12293_0, n12292_0}), .out(n544), .config_in(config_chain[359:357]), .config_rst(config_rst)); 
mux6 mux_120 (.in({n10003_2, n10002_0, n9973_0, n9972_0, n9941_0, n9940_0}), .out(n545), .config_in(config_chain[362:360]), .config_rst(config_rst)); 
mux6 mux_121 (.in({n12607_2, n12606_0, n12577_0, n12576_0, n12555_0, n12554_0}), .out(n546), .config_in(config_chain[365:363]), .config_rst(config_rst)); 
mux6 mux_122 (.in({n9753_2, n9752_0, n9721_0, n9720_0, n9691_1, n9690_0}), .out(n547), .config_in(config_chain[368:366]), .config_rst(config_rst)); 
mux6 mux_123 (.in({n12357_2, n12356_0, n12327_1, n12326_0, n12295_1, n12294_0}), .out(n548), .config_in(config_chain[371:369]), .config_rst(config_rst)); 
mux6 mux_124 (.in({n10005_2, n10004_0, n9983_0, n9982_0, n9951_0, n9950_0}), .out(n549), .config_in(config_chain[374:372]), .config_rst(config_rst)); 
mux6 mux_125 (.in({n12609_2, n12608_0, n12587_0, n12586_0, n12549_0, n12548_0}), .out(n550), .config_in(config_chain[377:375]), .config_rst(config_rst)); 
mux6 mux_126 (.in({n9755_2, n9754_0, n9723_1, n9722_0, n9693_0, n9692_0}), .out(n551), .config_in(config_chain[380:378]), .config_rst(config_rst)); 
mux6 mux_127 (.in({n12359_2, n12358_0, n12329_0, n12328_0, n12297_0, n12296_0}), .out(n552), .config_in(config_chain[383:381]), .config_rst(config_rst)); 
mux6 mux_128 (.in({n10007_2, n10006_0, n9977_0, n9976_0, n9947_1, n9946_0}), .out(n553), .config_in(config_chain[386:384]), .config_rst(config_rst)); 
mux6 mux_129 (.in({n12613_2, n12612_0, n12581_0, n12580_0, n12551_1, n12550_0}), .out(n554), .config_in(config_chain[389:387]), .config_rst(config_rst)); 
mux6 mux_130 (.in({n9757_2, n9756_0, n9727_0, n9726_0, n9695_0, n9694_0}), .out(n555), .config_in(config_chain[392:390]), .config_rst(config_rst)); 
mux6 mux_131 (.in({n12361_2, n12360_0, n12331_0, n12330_0, n12301_0, n12300_0}), .out(n556), .config_in(config_chain[395:393]), .config_rst(config_rst)); 
mux6 mux_132 (.in({n10233_0, n10232_0, n10203_0, n10202_0, n10181_1, n10180_0}), .out(n603), .config_in(config_chain[398:396]), .config_rst(config_rst)); 
mux6 mux_133 (.in({n12617_1, n12616_0, n12581_0, n12580_0, n12551_0, n12550_0}), .out(n604), .config_in(config_chain[401:399]), .config_rst(config_rst)); 
mux6 mux_134 (.in({n9981_0, n9980_0, n9949_0, n9948_0, n9927_0, n9926_0}), .out(n605), .config_in(config_chain[404:402]), .config_rst(config_rst)); 
mux6 mux_135 (.in({n12331_0, n12330_0, n12309_0, n12308_0, n12277_0, n12276_0}), .out(n606), .config_in(config_chain[407:405]), .config_rst(config_rst)); 
mux6 mux_136 (.in({n10235_0, n10234_0, n10213_1, n10212_0, n10183_0, n10182_0}), .out(n607), .config_in(config_chain[410:408]), .config_rst(config_rst)); 
mux6 mux_137 (.in({n12633_1, n12632_0, n12625_1, n12624_0, n12531_0, n12530_0}), .out(n608), .config_in(config_chain[413:411]), .config_rst(config_rst)); 
mux6 mux_138 (.in({n9991_0, n9990_0, n9953_0, n9952_0, n9921_0, n9920_0}), .out(n609), .config_in(config_chain[416:414]), .config_rst(config_rst)); 
mux6 mux_139 (.in({n12363_1, n12362_0, n12341_0, n12340_0, n12303_0, n12302_0}), .out(n610), .config_in(config_chain[419:417]), .config_rst(config_rst)); 
mux6 mux_140 (.in({n10247_0, n10246_0, n10215_0, n10214_0, n10177_0, n10176_0}), .out(n611), .config_in(config_chain[422:420]), .config_rst(config_rst)); 
mux6 mux_141 (.in({n12595_0, n12594_0, n12563_0, n12562_0, n12525_0, n12524_0}), .out(n612), .config_in(config_chain[425:423]), .config_rst(config_rst)); 
mux6 mux_142 (.in({n9985_0, n9984_0, n9955_1, n9954_0, n9923_1, n9922_0}), .out(n613), .config_in(config_chain[428:426]), .config_rst(config_rst)); 
mux6 mux_143 (.in({n12371_1, n12370_0, n12335_0, n12334_0, n12275_0, n12274_0}), .out(n614), .config_in(config_chain[431:429]), .config_rst(config_rst)); 
mux6 mux_144 (.in({n10241_0, n10240_0, n10209_0, n10208_0, n10179_0, n10178_0}), .out(n615), .config_in(config_chain[434:432]), .config_rst(config_rst)); 
mux6 mux_145 (.in({n12589_0, n12588_0, n12559_0, n12558_0, n12527_0, n12526_0}), .out(n616), .config_in(config_chain[437:435]), .config_rst(config_rst)); 
mux6 mux_146 (.in({n9987_1, n9986_0, n9957_0, n9956_0, n9935_0, n9934_0}), .out(n617), .config_in(config_chain[440:438]), .config_rst(config_rst)); 
mux6 mux_147 (.in({n12339_0, n12338_0, n12307_0, n12306_0, n12285_0, n12284_0}), .out(n618), .config_in(config_chain[443:441]), .config_rst(config_rst)); 
mux6 mux_148 (.in({n10243_0, n10242_0, n10221_1, n10220_0, n10189_1, n10188_0}), .out(n619), .config_in(config_chain[446:444]), .config_rst(config_rst)); 
mux6 mux_149 (.in({n12627_1, n12626_0, n12591_0, n12590_0, n12539_0, n12538_0}), .out(n620), .config_in(config_chain[449:447]), .config_rst(config_rst)); 
mux6 mux_150 (.in({n9989_0, n9988_0, n9967_0, n9966_0, n9929_0, n9928_0}), .out(n621), .config_in(config_chain[452:450]), .config_rst(config_rst)); 
mux6 mux_151 (.in({n12349_0, n12348_0, n12317_0, n12316_0, n12279_0, n12278_0}), .out(n622), .config_in(config_chain[455:453]), .config_rst(config_rst)); 
mux6 mux_152 (.in({n10253_1, n10252_0, n10223_0, n10222_0, n10191_0, n10190_0}), .out(n623), .config_in(config_chain[458:456]), .config_rst(config_rst)); 
mux6 mux_153 (.in({n12635_1, n12634_0, n12571_0, n12570_0, n12533_0, n12532_0}), .out(n624), .config_in(config_chain[461:459]), .config_rst(config_rst)); 
mux6 mux_154 (.in({n9993_0, n9992_0, n9961_0, n9960_0, n9931_1, n9930_0}), .out(n625), .config_in(config_chain[464:462]), .config_rst(config_rst)); 
mux6 mux_155 (.in({n12373_1, n12372_0, n12365_1, n12364_0, n12343_0, n12342_0}), .out(n626), .config_in(config_chain[467:465]), .config_rst(config_rst)); 
mux6 mux_156 (.in({n10255_0, n10254_0, n10217_0, n10216_0, n10187_0, n10186_0}), .out(n627), .config_in(config_chain[470:468]), .config_rst(config_rst)); 
mux6 mux_157 (.in({n12597_0, n12596_0, n12565_0, n12564_0, n12535_0, n12534_0}), .out(n628), .config_in(config_chain[473:471]), .config_rst(config_rst)); 
mux6 mux_158 (.in({n9995_1, n9994_0, n9965_0, n9964_0, n9933_0, n9932_0}), .out(n629), .config_in(config_chain[476:474]), .config_rst(config_rst)); 
mux6 mux_159 (.in({n12381_1, n12380_0, n12315_0, n12314_0, n12283_0, n12282_0}), .out(n630), .config_in(config_chain[479:477]), .config_rst(config_rst)); 
mux6 mux_160 (.in({n10249_0, n10248_0, n10219_0, n10218_0, n10197_1, n10196_0}), .out(n631), .config_in(config_chain[482:480]), .config_rst(config_rst)); 
mux6 mux_161 (.in({n12621_1, n12620_0, n12599_0, n12598_0, n12567_0, n12566_0}), .out(n632), .config_in(config_chain[485:483]), .config_rst(config_rst)); 
mux6 mux_162 (.in({n9997_0, n9996_0, n9975_0, n9974_0, n9943_0, n9942_0}), .out(n633), .config_in(config_chain[488:486]), .config_rst(config_rst)); 
mux6 mux_163 (.in({n12347_0, n12346_0, n12325_0, n12324_0, n12287_0, n12286_0}), .out(n634), .config_in(config_chain[491:489]), .config_rst(config_rst)); 
mux6 mux_164 (.in({n10265_2, n10264_0, n10229_1, n10228_0, n10199_0, n10198_0}), .out(n635), .config_in(config_chain[494:492]), .config_rst(config_rst)); 
mux6 mux_165 (.in({n12613_2, n12612_0, n12579_0, n12578_0, n12547_0, n12546_0}), .out(n636), .config_in(config_chain[497:495]), .config_rst(config_rst)); 
mux6 mux_166 (.in({n10011_2, n10010_0, n9969_0, n9968_0, n9939_1, n9938_0}), .out(n637), .config_in(config_chain[500:498]), .config_rst(config_rst)); 
mux6 mux_167 (.in({n12367_1, n12366_0, n12361_2, n12360_0, n12319_0, n12318_0}), .out(n638), .config_in(config_chain[503:501]), .config_rst(config_rst)); 
mux6 mux_168 (.in({n10267_2, n10266_0, n10231_0, n10230_0, n10193_0, n10192_0}), .out(n639), .config_in(config_chain[506:504]), .config_rst(config_rst)); 
mux6 mux_169 (.in({n12615_2, n12614_0, n12573_0, n12572_0, n12541_0, n12540_0}), .out(n640), .config_in(config_chain[509:507]), .config_rst(config_rst)); 
mux6 mux_170 (.in({n10001_2, n10000_0, n9971_1, n9970_0, n9941_0, n9940_0}), .out(n641), .config_in(config_chain[512:510]), .config_rst(config_rst)); 
mux6 mux_171 (.in({n12375_1, n12374_0, n12353_2, n12352_0, n12291_0, n12290_0}), .out(n642), .config_in(config_chain[515:513]), .config_rst(config_rst)); 
mux6 mux_172 (.in({n10257_1, n10256_0, n10227_0, n10226_0, n10195_0, n10194_0}), .out(n643), .config_in(config_chain[518:516]), .config_rst(config_rst)); 
mux6 mux_173 (.in({n12623_1, n12622_0, n12605_1, n12604_0, n12575_0, n12574_0}), .out(n644), .config_in(config_chain[521:519]), .config_rst(config_rst)); 
mux6 mux_174 (.in({n10005_2, n10004_0, n9973_0, n9972_0, n9951_0, n9950_0}), .out(n645), .config_in(config_chain[524:522]), .config_rst(config_rst)); 
mux6 mux_175 (.in({n12355_2, n12354_0, n12333_0, n12332_0, n12301_0, n12300_0}), .out(n646), .config_in(config_chain[527:525]), .config_rst(config_rst)); 
mux6 mux_176 (.in({n10259_2, n10258_0, n10237_1, n10236_0, n10205_1, n10204_0}), .out(n647), .config_in(config_chain[530:528]), .config_rst(config_rst)); 
mux6 mux_177 (.in({n12631_1, n12630_0, n12607_2, n12606_0, n12555_0, n12554_0}), .out(n648), .config_in(config_chain[533:531]), .config_rst(config_rst)); 
mux6 mux_178 (.in({n10007_2, n10006_0, n9983_0, n9982_0, n9945_0, n9944_0}), .out(n649), .config_in(config_chain[536:534]), .config_rst(config_rst)); 
mux6 mux_179 (.in({n12357_2, n12356_0, n12327_0, n12326_0, n12295_0, n12294_0}), .out(n650), .config_in(config_chain[539:537]), .config_rst(config_rst)); 
mux6 mux_180 (.in({n10261_2, n10260_0, n10239_0, n10238_0, n10201_0, n10200_0}), .out(n651), .config_in(config_chain[542:540]), .config_rst(config_rst)); 
mux6 mux_181 (.in({n12611_2, n12610_0, n12587_0, n12586_0, n12549_0, n12548_0}), .out(n652), .config_in(config_chain[545:543]), .config_rst(config_rst)); 
mux6 mux_182 (.in({n10009_2, n10008_0, n9979_1, n9978_0, n9947_1, n9946_0}), .out(n653), .config_in(config_chain[548:546]), .config_rst(config_rst)); 
mux6 mux_183 (.in({n12377_1, n12376_0, n12359_2, n12358_0, n12299_0, n12298_0}), .out(n654), .config_in(config_chain[551:549]), .config_rst(config_rst)); 
mux6 mux_184 (.in({n10497_1, n10496_0, n10459_0, n10458_0, n10437_0, n10436_0}), .out(n701), .config_in(config_chain[554:552]), .config_rst(config_rst)); 
mux6 mux_185 (.in({n12651_1, n12650_0, n12549_0, n12548_0, n12527_0, n12526_0}), .out(n702), .config_in(config_chain[557:555]), .config_rst(config_rst)); 
mux6 mux_186 (.in({n10235_0, n10234_0, n10203_0, n10202_0/**/, n10181_1, n10180_0}), .out(n703), .config_in(config_chain[560:558]), .config_rst(config_rst)); 
mux6 mux_187 (.in({n12391_1, n12390_0, n12383_1, n12382_0, n12377_0, n12376_0}), .out(n704), .config_in(config_chain[563:561]), .config_rst(config_rst)); 
mux6 mux_188 (.in({n10491_0, n10490_0/**/, n10469_0, n10468_0, n10439_0, n10438_0}), .out(n705), .config_in(config_chain[566:564]), .config_rst(config_rst)); 
mux6 mux_189 (.in({n12617_0, n12616_0/**/, n12591_0, n12590_0, n12559_0, n12558_0}), .out(n706), .config_in(config_chain[569:567]), .config_rst(config_rst)); 
mux6 mux_190 (.in({n10245_1, n10244_0, n10215_0, n10214_0, n10183_0, n10182_0}), .out(n707), .config_in(config_chain[572:570]), .config_rst(config_rst)); 
mux6 mux_191 (.in({n12399_1, n12398_0, n12309_0, n12308_0, n12271_0, n12270_0}), .out(n708), .config_in(config_chain[575:573]), .config_rst(config_rst)); 
mux6 mux_192 (.in({n10503_0, n10502_0, n10471_0, n10470_0, n10441_1, n10440_0}), .out(n709), .config_in(config_chain[578:576]), .config_rst(config_rst)); 
mux6 mux_193 (.in({n12637_1, n12636_0, n12633_0, n12632_0, n12625_0, n12624_0}), .out(n710), .config_in(config_chain[581:579]), .config_rst(config_rst)); 
mux6 mux_194 (.in({n10247_0/**/, n10246_0, n10209_0, n10208_0, n10177_0, n10176_0}), .out(n711), .config_in(config_chain[584:582]), .config_rst(config_rst)); 
mux6 mux_195 (.in({n12363_0, n12362_0, n12341_0, n12340_0, n12303_0, n12302_0}), .out(n712), .config_in(config_chain[587:585]), .config_rst(config_rst)); 
mux6 mux_196 (.in({n10505_1, n10504_0, n10473_1, n10472_0, n10435_0, n10434_0}), .out(n713), .config_in(config_chain[590:588]), .config_rst(config_rst)); 
mux6 mux_197 (.in({n12653_1, n12652_0, n12557_0, n12556_0, n12525_0, n12524_0}), .out(n714), .config_in(config_chain[593:591]), .config_rst(config_rst)); 
mux6 mux_198 (.in({n10241_0/**/, n10240_0, n10211_0, n10210_0, n10189_1, n10188_0}), .out(n715), .config_in(config_chain[596:594]), .config_rst(config_rst)); 
mux6 mux_199 (.in({n12385_1, n12384_0, n12379_0, n12378_0, n12371_0, n12370_0}), .out(n716), .config_in(config_chain[599:597]), .config_rst(config_rst)); 
mux6 mux_200 (.in({n10499_0, n10498_0, n10477_0, n10476_0, n10445_0, n10444_0/**/}), .out(n717), .config_in(config_chain[602:600]), .config_rst(config_rst)); 
mux6 mux_201 (.in({n12619_0, n12618_0, n12589_0, n12588_0/**/, n12567_0, n12566_0}), .out(n718), .config_in(config_chain[605:603]), .config_rst(config_rst)); 
mux6 mux_202 (.in({n10243_0, n10242_0, n10221_1, n10220_0, n10191_0, n10190_0}), .out(n719), .config_in(config_chain[608:606]), .config_rst(config_rst)); 
mux6 mux_203 (.in({n12401_1, n12400_0, n12393_1, n12392_0/**/, n12285_0, n12284_0}), .out(n720), .config_in(config_chain[611:609]), .config_rst(config_rst)); 
mux6 mux_204 (.in({n10509_0, n10508_0, n10479_0, n10478_0, n10447_0, n10446_0}), .out(n721), .config_in(config_chain[614:612]), .config_rst(config_rst)); 
mux6 mux_205 (.in({n12639_1, n12638_0, n12627_0, n12626_0, n12599_0, n12598_0}), .out(n722), .config_in(config_chain[617:615]), .config_rst(config_rst)); 
mux6 mux_206 (.in({n10255_0, n10254_0, n10223_0/**/, n10222_0, n10185_0, n10184_0}), .out(n723), .config_in(config_chain[620:618]), .config_rst(config_rst)); 
mux6 mux_207 (.in({n12349_0, n12348_0, n12311_0, n12310_0, n12279_0, n12278_0}), .out(n724), .config_in(config_chain[623:621]), .config_rst(config_rst)); 
mux6 mux_208 (.in({n10511_0, n10510_0, n10481_1, n10480_0, n10443_0, n10442_0}), .out(n725), .config_in(config_chain[626:624]), .config_rst(config_rst)); 
mux6 mux_209 (.in({n12655_1, n12654_0, n12647_1, n12646_0, n12533_0, n12532_0}), .out(n726), .config_in(config_chain[629:627]), .config_rst(config_rst)); 
mux6 mux_210 (.in({n10249_0, n10248_0, n10219_0, n10218_0, n10187_0, n10186_0}), .out(n727), .config_in(config_chain[632:630]), .config_rst(config_rst)); 
mux6 mux_211 (.in({n12373_0/**/, n12372_0, n12365_0, n12364_0, n12343_0, n12342_0}), .out(n728), .config_in(config_chain[635:633]), .config_rst(config_rst)); 
mux6 mux_212 (.in({n10513_1, n10512_0, n10475_0, n10474_0, n10453_0/**/, n10452_0}), .out(n729), .config_in(config_chain[638:636]), .config_rst(config_rst)); 
mux6 mux_213 (.in({n12597_0, n12596_0, n12565_0, n12564_0, n12543_0, n12542_0}), .out(n730), .config_in(config_chain[641:639]), .config_rst(config_rst)); 
mux6 mux_214 (.in({n10251_0, n10250_0, n10229_1, n10228_0, n10197_1, n10196_0}), .out(n731), .config_in(config_chain[644:642]), .config_rst(config_rst)); 
mux6 mux_215 (.in({n12395_1, n12394_0, n12381_0, n12380_0/**/, n12293_0, n12292_0}), .out(n732), .config_in(config_chain[647:645]), .config_rst(config_rst)); 
mux6 mux_216 (.in({n10521_2, n10520_0, n10485_0, n10484_0/**/, n10455_0, n10454_0}), .out(n733), .config_in(config_chain[650:648]), .config_rst(config_rst)); 
mux6 mux_217 (.in({n12629_0/**/, n12628_0, n12621_0, n12620_0, n12611_2, n12610_0}), .out(n734), .config_in(config_chain[653:651]), .config_rst(config_rst)); 
mux6 mux_218 (.in({n10265_2, n10264_0, n10231_0/**/, n10230_0, n10193_0, n10192_0}), .out(n735), .config_in(config_chain[656:654]), .config_rst(config_rst)); 
mux6 mux_219 (.in({n12359_2/**/, n12358_0, n12325_0, n12324_0, n12287_0, n12286_0}), .out(n736), .config_in(config_chain[659:657]), .config_rst(config_rst)); 
mux6 mux_220 (.in({n10523_2, n10522_0, n10487_0, n10486_0, n10457_1, n10456_0}), .out(n737), .config_in(config_chain[662:660]), .config_rst(config_rst)); 
mux6 mux_221 (.in({n12649_1/**/, n12648_0, n12641_1, n12640_0, n12613_2, n12612_0}), .out(n738), .config_in(config_chain[665:663]), .config_rst(config_rst)); 
mux6 mux_222 (.in({n10267_2, n10266_0, n10225_0, n10224_0, n10195_0, n10194_0}), .out(n739), .config_in(config_chain[668:666]), .config_rst(config_rst)); 
mux6 mux_223 (.in({n12367_0, n12366_0, n12351_1, n12350_0, n12319_0, n12318_0}), .out(n740), .config_in(config_chain[671:669]), .config_rst(config_rst)); 
mux6 mux_224 (.in({n10525_2, n10524_0, n10483_0, n10482_0, n10451_0/**/, n10450_0}), .out(n741), .config_in(config_chain[674:672]), .config_rst(config_rst)); 
mux6 mux_225 (.in({n12615_2, n12614_0, n12573_0, n12572_0, n12551_0, n12550_0}), .out(n742), .config_in(config_chain[677:675]), .config_rst(config_rst)); 
mux6 mux_226 (.in({n10259_2, n10258_0, n10227_0, n10226_0, n10205_1/**/, n10204_0}), .out(n743), .config_in(config_chain[680:678]), .config_rst(config_rst)); 
mux6 mux_227 (.in({n12397_1, n12396_0, n12389_1, n12388_0, n12353_2, n12352_0}), .out(n744), .config_in(config_chain[683:681]), .config_rst(config_rst)); 
mux6 mux_228 (.in({n10515_1/**/, n10514_0, n10493_0, n10492_0, n10461_0, n10460_0}), .out(n745), .config_in(config_chain[686:684]), .config_rst(config_rst)); 
mux6 mux_229 (.in({n12623_0, n12622_0, n12605_1, n12604_0, n12583_0, n12582_0}), .out(n746), .config_in(config_chain[689:687]), .config_rst(config_rst)); 
mux6 mux_230 (.in({n10261_2, n10260_0, n10237_1, n10236_0, n10207_0, n10206_0}), .out(n747), .config_in(config_chain[692:690]), .config_rst(config_rst)); 
mux6 mux_231 (.in({n12355_2, n12354_0, n12333_0, n12332_0, n12301_0, n12300_0}), .out(n748), .config_in(config_chain[695:693]), .config_rst(config_rst)); 
mux6 mux_232 (.in({n10517_1, n10516_0, n10495_0, n10494_0, n10465_1, n10464_0}), .out(n749), .config_in(config_chain[698:696]), .config_rst(config_rst)); 
mux6 mux_233 (.in({n12643_1, n12642_0, n12631_0, n12630_0, n12609_2, n12608_0}), .out(n750), .config_in(config_chain[701:699]), .config_rst(config_rst)); 
mux6 mux_234 (.in({n10263_2, n10262_0, n10233_0/**/, n10232_0, n10201_0, n10200_0}), .out(n751), .config_in(config_chain[704:702]), .config_rst(config_rst)); 
mux6 mux_235 (.in({n12369_0/**/, n12368_0, n12357_2, n12356_0, n12327_0, n12326_0}), .out(n752), .config_in(config_chain[707:705]), .config_rst(config_rst)); 
mux6 mux_236 (.in({n10755_0/**/, n10754_0, n10725_0, n10724_0, n10695_1, n10694_0}), .out(n799), .config_in(config_chain[710:708]), .config_rst(config_rst)); 
mux6 mux_237 (.in({n12657_1, n12656_0, n12643_0, n12642_0, n12631_0, n12630_0}), .out(n800), .config_in(config_chain[713:711]), .config_rst(config_rst)); 
mux6 mux_238 (.in({n10491_0, n10490_0, n10459_0, n10458_0, n10437_0, n10436_0}), .out(n801), .config_in(config_chain[716:714]), .config_rst(config_rst)); 
mux6 mux_239 (.in({n12371_0/**/, n12370_0, n12363_0, n12362_0, n12327_0, n12326_1}), .out(n802), .config_in(config_chain[719:717]), .config_rst(config_rst)); 
mux6 mux_240 (.in({n10757_0, n10756_0, n10727_1, n10726_0, n10697_0, n10696_0}), .out(n803), .config_in(config_chain[722:720]), .config_rst(config_rst)); 
mux6 mux_241 (.in({n12673_1, n12672_0, n12665_1, n12664_0, n12527_0, n12526_1}), .out(n804), .config_in(config_chain[725:723]), .config_rst(config_rst)); 
mux6 mux_242 (.in({n10501_0, n10500_0, n10471_0, n10470_0, n10439_0, n10438_0}), .out(n805), .config_in(config_chain[728:726]), .config_rst(config_rst)); 
mux6 mux_243 (.in({n12403_1, n12402_0, n12391_0, n12390_0, n12379_0, n12378_0}), .out(n806), .config_in(config_chain[731:729]), .config_rst(config_rst)); 
mux6 mux_244 (.in({n10761_0, n10760_0, n10729_0, n10728_0, n10699_0, n10698_0}), .out(n807), .config_in(config_chain[734:732]), .config_rst(config_rst)); 
mux6 mux_245 (.in({n12617_0, n12616_0, n12591_0, n12590_1, n12559_0, n12558_1/**/}), .out(n808), .config_in(config_chain[737:735]), .config_rst(config_rst)); 
mux6 mux_246 (.in({n10503_0, n10502_0, n10473_1, n10472_0, n10441_1, n10440_0}), .out(n809), .config_in(config_chain[740:738]), .config_rst(config_rst)); 
mux6 mux_247 (.in({n12411_1, n12410_0, n12399_0, n12398_0, n12271_0, n12270_1}), .out(n810), .config_in(config_chain[743:741]), .config_rst(config_rst)); 
mux6 mux_248 (.in({n10763_0, n10762_0, n10731_0, n10730_0, n10701_0, n10700_0}), .out(n811), .config_in(config_chain[746:744]), .config_rst(config_rst)); 
mux6 mux_249 (.in({n12645_0, n12644_0, n12637_0, n12636_0, n12633_0, n12632_0}), .out(n812), .config_in(config_chain[749:747]), .config_rst(config_rst)); 
mux6 mux_250 (.in({n10505_1, n10504_0, n10467_0, n10466_0/**/, n10445_0, n10444_0}), .out(n813), .config_in(config_chain[752:750]), .config_rst(config_rst)); 
mux6 mux_251 (.in({n12365_0/**/, n12364_0, n12335_0, n12334_1, n12303_0, n12302_1}), .out(n814), .config_in(config_chain[755:753]), .config_rst(config_rst)); 
mux6 mux_252 (.in({n10765_0, n10764_0/**/, n10735_1, n10734_0, n10703_1, n10702_0}), .out(n815), .config_in(config_chain[758:756]), .config_rst(config_rst)); 
mux6 mux_253 (.in({n12667_1, n12666_0, n12653_0, n12652_0, n12535_0, n12534_1}), .out(n816), .config_in(config_chain[761:759]), .config_rst(config_rst)); 
mux6 mux_254 (.in({n10499_0, n10498_0, n10477_0, n10476_0, n10447_0/**/, n10446_0}), .out(n817), .config_in(config_chain[764:762]), .config_rst(config_rst)); 
mux6 mux_255 (.in({n12385_0, n12384_0, n12381_0, n12380_0, n12373_0/**/, n12372_0}), .out(n818), .config_in(config_chain[767:765]), .config_rst(config_rst)); 
mux6 mux_256 (.in({n10767_1, n10766_0, n10737_0, n10736_0, n10705_0/**/, n10704_0}), .out(n819), .config_in(config_chain[770:768]), .config_rst(config_rst)); 
mux6 mux_257 (.in({n12675_1, n12674_0, n12619_0, n12618_0/**/, n12567_0, n12566_1}), .out(n820), .config_in(config_chain[773:771]), .config_rst(config_rst)); 
mux6 mux_258 (.in({n10511_0, n10510_0, n10479_0, n10478_0, n10449_1, n10448_0}), .out(n821), .config_in(config_chain[776:774]), .config_rst(config_rst)); 
mux6 mux_259 (.in({n12413_1, n12412_0, n12405_1, n12404_0/**/, n12401_0, n12400_0}), .out(n822), .config_in(config_chain[779:777]), .config_rst(config_rst)); 
mux6 mux_260 (.in({n10769_0, n10768_0, n10739_0, n10738_0/**/, n10709_0, n10708_0}), .out(n823), .config_in(config_chain[782:780]), .config_rst(config_rst)); 
mux6 mux_261 (.in({n12639_0, n12638_0, n12635_0, n12634_0, n12627_0, n12626_0/**/}), .out(n824), .config_in(config_chain[785:783]), .config_rst(config_rst)); 
mux6 mux_262 (.in({n10513_1, n10512_0, n10475_0, n10474_0, n10443_0, n10442_0}), .out(n825), .config_in(config_chain[788:786]), .config_rst(config_rst)); 
mux6 mux_263 (.in({n12421_1, n12420_0, n12311_0, n12310_1, n12279_0/**/, n12278_1}), .out(n826), .config_in(config_chain[791:789]), .config_rst(config_rst)); 
mux6 mux_264 (.in({n10771_0, n10770_0, n10741_0, n10740_0, n10711_1, n10710_0}), .out(n827), .config_in(config_chain[794:792]), .config_rst(config_rst)); 
mux6 mux_265 (.in({n12661_1, n12660_0, n12655_0, n12654_0, n12647_0, n12646_0}), .out(n828), .config_in(config_chain[797:795]), .config_rst(config_rst)); 
mux6 mux_266 (.in({n10507_0, n10506_0, n10485_0, n10484_0, n10453_0, n10452_0}), .out(n829), .config_in(config_chain[800:798]), .config_rst(config_rst)); 
mux6 mux_267 (.in({n12387_0, n12386_0, n12375_0/**/, n12374_0, n12343_0, n12342_1}), .out(n830), .config_in(config_chain[803:801]), .config_rst(config_rst)); 
mux6 mux_268 (.in({n10779_1, n10778_0, n10743_1, n10742_0, n10713_0, n10712_0}), .out(n831), .config_in(config_chain[806:804]), .config_rst(config_rst)); 
mux6 mux_269 (.in({n12609_1, n12608_1, n12575_0, n12574_1, n12543_0, n12542_1/**/}), .out(n832), .config_in(config_chain[809:807]), .config_rst(config_rst)); 
mux6 mux_270 (.in({n10521_2, n10520_0, n10487_0, n10486_0, n10457_1, n10456_0}), .out(n833), .config_in(config_chain[812:810]), .config_rst(config_rst)); 
mux6 mux_271 (.in({n12407_1, n12406_0, n12395_0/**/, n12394_0, n12357_1, n12356_1}), .out(n834), .config_in(config_chain[815:813]), .config_rst(config_rst)); 
mux6 mux_272 (.in({n10781_2, n10780_0, n10745_0, n10744_0, n10715_0, n10714_0}), .out(n835), .config_in(config_chain[818:816]), .config_rst(config_rst)); 
mux6 mux_273 (.in({n12629_0, n12628_0, n12621_0, n12620_0/**/, n12611_1, n12610_1}), .out(n836), .config_in(config_chain[821:819]), .config_rst(config_rst)); 
mux6 mux_274 (.in({n10523_2, n10522_0, n10489_1, n10488_0, n10451_0/**/, n10450_0}), .out(n837), .config_in(config_chain[824:822]), .config_rst(config_rst)); 
mux6 mux_275 (.in({n12415_1, n12414_0/**/, n12361_1, n12360_1, n12287_0, n12286_1}), .out(n838), .config_in(config_chain[827:825]), .config_rst(config_rst)); 
mux6 mux_276 (.in({n10783_2, n10782_0, n10749_0/**/, n10748_0, n10717_0, n10716_0}), .out(n839), .config_in(config_chain[830:828]), .config_rst(config_rst)); 
mux6 mux_277 (.in({n12663_1, n12662_0/**/, n12649_0, n12648_0, n12613_1, n12612_1}), .out(n840), .config_in(config_chain[833:831]), .config_rst(config_rst)); 
mux6 mux_278 (.in({n10515_1, n10514_0, n10483_0/**/, n10482_0, n10461_0, n10460_0}), .out(n841), .config_in(config_chain[836:834]), .config_rst(config_rst)); 
mux6 mux_279 (.in({n12377_0, n12376_0, n12369_0, n12368_0, n12351_1/**/, n12350_1}), .out(n842), .config_in(config_chain[839:837]), .config_rst(config_rst)); 
mux6 mux_280 (.in({n10785_2, n10784_0, n10751_1, n10750_0, n10719_1, n10718_0}), .out(n843), .config_in(config_chain[842:840]), .config_rst(config_rst)); 
mux6 mux_281 (.in({n12671_1, n12670_0/**/, n12615_1, n12614_1, n12551_0, n12550_1}), .out(n844), .config_in(config_chain[845:843]), .config_rst(config_rst)); 
mux6 mux_282 (.in({n10517_1, n10516_0, n10493_0, n10492_0, n10463_0, n10462_0}), .out(n845), .config_in(config_chain[848:846]), .config_rst(config_rst)); 
mux6 mux_283 (.in({n12397_0, n12396_0, n12389_0, n12388_0, n12353_1, n12352_1}), .out(n846), .config_in(config_chain[851:849]), .config_rst(config_rst)); 
mux6 mux_284 (.in({n10775_1, n10774_0, n10753_0, n10752_0, n10723_0/**/, n10722_0}), .out(n847), .config_in(config_chain[854:852]), .config_rst(config_rst)); 
mux6 mux_285 (.in({n12623_0/**/, n12622_0, n12607_1, n12606_1, n12583_0, n12582_1}), .out(n848), .config_in(config_chain[857:855]), .config_rst(config_rst)); 
mux6 mux_286 (.in({n10519_2, n10518_0, n10497_1, n10496_0, n10465_1, n10464_0}), .out(n849), .config_in(config_chain[860:858]), .config_rst(config_rst)); 
mux6 mux_287 (.in({n12417_1, n12416_0/**/, n12355_1, n12354_1, n12295_0, n12294_1}), .out(n850), .config_in(config_chain[863:861]), .config_rst(config_rst)); 
mux6 mux_288 (.in({n11015_1, n11014_0, n10985_0, n10984_0, n10963_0, n10962_0}), .out(n897), .config_in(config_chain[866:864]), .config_rst(config_rst)); 
mux6 mux_289 (.in({n12691_1, n12690_0, n12637_0, n12636_0, n12623_0, n12622_1}), .out(n898), .config_in(config_chain[869:867]), .config_rst(config_rst)); 
mux6 mux_290 (.in({n10757_0, n10756_0, n10725_0, n10724_0, n10695_1, n10694_0}), .out(n899), .config_in(config_chain[872:870]), .config_rst(config_rst)); 
mux6 mux_291 (.in({n12431_1, n12430_0, n12423_1, n12422_0, n12417_0/**/, n12416_0}), .out(n900), .config_in(config_chain[875:873]), .config_rst(config_rst)); 
mux6 mux_292 (.in({n11017_0/**/, n11016_0, n10995_0, n10994_0, n10957_0, n10956_0}), .out(n901), .config_in(config_chain[878:876]), .config_rst(config_rst)); 
mux6 mux_293 (.in({n12657_0, n12656_0, n12653_0, n12652_0, n12645_0, n12644_0}), .out(n902), .config_in(config_chain[881:879]), .config_rst(config_rst)); 
mux6 mux_294 (.in({n10759_1, n10758_0, n10729_0, n10728_0, n10697_0, n10696_0}), .out(n903), .config_in(config_chain[884:882]), .config_rst(config_rst)); 
mux6 mux_295 (.in({n12439_1, n12438_0, n12383_0, n12382_0, n12371_0/**/, n12370_1}), .out(n904), .config_in(config_chain[887:885]), .config_rst(config_rst)); 
mux6 mux_296 (.in({n11021_0, n11020_0, n10989_0, n10988_0, n10959_1, n10958_0}), .out(n905), .config_in(config_chain[890:888]), .config_rst(config_rst)); 
mux6 mux_297 (.in({n12677_1, n12676_0, n12673_0, n12672_0, n12665_0, n12664_0}), .out(n906), .config_in(config_chain[893:891]), .config_rst(config_rst)); 
mux6 mux_298 (.in({n10761_0, n10760_0, n10731_0, n10730_0, n10699_0, n10698_0}), .out(n907), .config_in(config_chain[896:894]), .config_rst(config_rst)); 
mux6 mux_299 (.in({n12403_0, n12402_0/**/, n12391_0, n12390_0, n12379_0, n12378_1}), .out(n908), .config_in(config_chain[899:897]), .config_rst(config_rst)); 
mux6 mux_300 (.in({n11023_1, n11022_0, n10991_1, n10990_0, n10961_0, n10960_0}), .out(n909), .config_in(config_chain[902:900]), .config_rst(config_rst)); 
mux6 mux_301 (.in({n12693_1, n12692_0, n12625_0, n12624_1/**/, n12617_0, n12616_1}), .out(n910), .config_in(config_chain[905:903]), .config_rst(config_rst)); 
mux6 mux_302 (.in({n10763_0/**/, n10762_0, n10733_0, n10732_0, n10703_1, n10702_0}), .out(n911), .config_in(config_chain[908:906]), .config_rst(config_rst)); 
mux6 mux_303 (.in({n12425_1, n12424_0, n12419_0, n12418_0, n12411_0/**/, n12410_0}), .out(n912), .config_in(config_chain[911:909]), .config_rst(config_rst)); 
mux6 mux_304 (.in({n11025_0, n11024_0/**/, n11003_0, n11002_0, n10971_0, n10970_0}), .out(n913), .config_in(config_chain[914:912]), .config_rst(config_rst)); 
mux6 mux_305 (.in({n12659_0, n12658_0, n12647_0, n12646_0, n12633_0, n12632_1}), .out(n914), .config_in(config_chain[917:915]), .config_rst(config_rst)); 
mux6 mux_306 (.in({n10765_0, n10764_0, n10735_1, n10734_0, n10705_0, n10704_0/**/}), .out(n915), .config_in(config_chain[920:918]), .config_rst(config_rst)); 
mux6 mux_307 (.in({n12441_1, n12440_0/**/, n12433_1, n12432_0, n12365_0, n12364_1}), .out(n916), .config_in(config_chain[923:921]), .config_rst(config_rst)); 
mux6 mux_308 (.in({n11035_0, n11034_0, n10997_0, n10996_0, n10965_0/**/, n10964_0}), .out(n917), .config_in(config_chain[926:924]), .config_rst(config_rst)); 
mux6 mux_309 (.in({n12679_1, n12678_0, n12667_0, n12666_0, n12655_0, n12654_0}), .out(n918), .config_in(config_chain[929:927]), .config_rst(config_rst)); 
mux6 mux_310 (.in({n10769_0, n10768_0, n10737_0, n10736_0, n10707_0, n10706_0}), .out(n919), .config_in(config_chain[932:930]), .config_rst(config_rst)); 
mux6 mux_311 (.in({n12393_0, n12392_0, n12385_0/**/, n12384_0, n12381_0, n12380_1}), .out(n920), .config_in(config_chain[935:933]), .config_rst(config_rst)); 
mux6 mux_312 (.in({n11029_0, n11028_0, n10999_1, n10998_0, n10969_0, n10968_0}), .out(n921), .config_in(config_chain[938:936]), .config_rst(config_rst)); 
mux6 mux_313 (.in({n12695_1, n12694_0, n12687_1, n12686_0, n12619_0, n12618_1}), .out(n922), .config_in(config_chain[941:939]), .config_rst(config_rst)); 
mux6 mux_314 (.in({n10771_0, n10770_0, n10741_0, n10740_0, n10709_0, n10708_0}), .out(n923), .config_in(config_chain[944:942]), .config_rst(config_rst)); 
mux6 mux_315 (.in({n12413_0, n12412_0/**/, n12405_0, n12404_0, n12401_0, n12400_0}), .out(n924), .config_in(config_chain[947:945]), .config_rst(config_rst)); 
mux6 mux_316 (.in({n11031_1, n11030_0, n11001_0/**/, n11000_0, n10979_0, n10978_0}), .out(n925), .config_in(config_chain[950:948]), .config_rst(config_rst)); 
mux6 mux_317 (.in({n12641_0, n12640_0, n12635_0, n12634_1/**/, n12627_0, n12626_1}), .out(n926), .config_in(config_chain[953:951]), .config_rst(config_rst)); 
mux6 mux_318 (.in({n10773_0, n10772_0, n10743_1, n10742_0, n10711_1, n10710_0}), .out(n927), .config_in(config_chain[956:954]), .config_rst(config_rst)); 
mux6 mux_319 (.in({n12435_1, n12434_0/**/, n12421_0, n12420_0, n12367_0, n12366_1}), .out(n928), .config_in(config_chain[959:957]), .config_rst(config_rst)); 
mux6 mux_320 (.in({n11039_1, n11038_0, n11011_0, n11010_0/**/, n10973_0, n10972_0}), .out(n929), .config_in(config_chain[962:960]), .config_rst(config_rst)); 
mux6 mux_321 (.in({n12669_0, n12668_0, n12661_0/**/, n12660_0, n12607_1, n12606_1}), .out(n930), .config_in(config_chain[965:963]), .config_rst(config_rst)); 
mux6 mux_322 (.in({n10779_1, n10778_0, n10745_0/**/, n10744_0, n10715_0, n10714_0}), .out(n931), .config_in(config_chain[968:966]), .config_rst(config_rst)); 
mux6 mux_323 (.in({n12387_0, n12386_0, n12375_0, n12374_1, n12355_1, n12354_1}), .out(n932), .config_in(config_chain[971:969]), .config_rst(config_rst)); 
mux6 mux_324 (.in({n11041_1, n11040_0, n11005_0, n11004_0, n10975_1, n10974_0}), .out(n933), .config_in(config_chain[974:972]), .config_rst(config_rst)); 
mux6 mux_325 (.in({n12689_1/**/, n12688_0, n12681_1, n12680_0, n12609_1, n12608_1}), .out(n934), .config_in(config_chain[977:975]), .config_rst(config_rst)); 
mux6 mux_326 (.in({n10781_2, n10780_0, n10747_0, n10746_0, n10717_0, n10716_0}), .out(n935), .config_in(config_chain[980:978]), .config_rst(config_rst)); 
mux6 mux_327 (.in({n12407_0/**/, n12406_0, n12395_0, n12394_0, n12359_1, n12358_1}), .out(n936), .config_in(config_chain[983:981]), .config_rst(config_rst)); 
mux6 mux_328 (.in({n11043_1, n11042_0, n11009_0, n11008_0, n10977_0/**/, n10976_0}), .out(n937), .config_in(config_chain[986:984]), .config_rst(config_rst)); 
mux6 mux_329 (.in({n12643_0, n12642_0, n12629_0, n12628_1, n12611_1, n12610_1}), .out(n938), .config_in(config_chain[989:987]), .config_rst(config_rst)); 
mux6 mux_330 (.in({n10785_2, n10784_0, n10749_0, n10748_0, n10719_1, n10718_0}), .out(n939), .config_in(config_chain[992:990]), .config_rst(config_rst)); 
mux6 mux_331 (.in({n12437_1, n12436_0, n12429_1, n12428_0, n12361_1, n12360_1}), .out(n940), .config_in(config_chain[995:993]), .config_rst(config_rst)); 
mux6 mux_332 (.in({n11045_2, n11044_0, n11019_0, n11018_0, n10987_0, n10986_0}), .out(n941), .config_in(config_chain[998:996]), .config_rst(config_rst)); 
mux6 mux_333 (.in({n12663_0, n12662_0, n12651_0, n12650_0, n12613_1, n12612_1}), .out(n942), .config_in(config_chain[1001:999]), .config_rst(config_rst)); 
mux6 mux_334 (.in({n10775_1, n10774_0, n10751_1, n10750_0, n10721_0/**/, n10720_0}), .out(n943), .config_in(config_chain[1004:1002]), .config_rst(config_rst)); 
mux6 mux_335 (.in({n12377_0/**/, n12376_1, n12369_0, n12368_1, n12351_1, n12350_1}), .out(n944), .config_in(config_chain[1007:1005]), .config_rst(config_rst)); 
mux6 mux_336 (.in({n11047_2, n11046_0, n11013_0, n11012_0, n10983_1, n10982_0}), .out(n945), .config_in(config_chain[1010:1008]), .config_rst(config_rst)); 
mux6 mux_337 (.in({n12683_1, n12682_0/**/, n12671_0, n12670_0, n12605_0, n12604_1}), .out(n946), .config_in(config_chain[1013:1011]), .config_rst(config_rst)); 
mux6 mux_338 (.in({n10777_1, n10776_0, n10755_0, n10754_0, n10723_0, n10722_0/**/}), .out(n947), .config_in(config_chain[1016:1014]), .config_rst(config_rst)); 
mux6 mux_339 (.in({n12409_0, n12408_0, n12397_0, n12396_0/**/, n12353_1, n12352_1}), .out(n948), .config_in(config_chain[1019:1017]), .config_rst(config_rst)); 
mux6 mux_340 (.in({n11277_0, n11276_0, n11247_0, n11246_0, n11225_1, n11224_0}), .out(n995), .config_in(config_chain[1022:1020]), .config_rst(config_rst)); 
mux6 mux_341 (.in({n12697_1, n12696_0, n12683_0, n12682_0, n12671_0, n12670_0}), .out(n996), .config_in(config_chain[1025:1023]), .config_rst(config_rst)); 
mux6 mux_342 (.in({n11017_0, n11016_0, n10985_0, n10984_0, n10963_0, n10962_0}), .out(n997), .config_in(config_chain[1028:1026]), .config_rst(config_rst)); 
mux6 mux_343 (.in({n12411_0, n12410_0, n12403_0, n12402_0, n12397_0, n12396_1}), .out(n998), .config_in(config_chain[1031:1029]), .config_rst(config_rst)); 
mux6 mux_344 (.in({n11279_0, n11278_0, n11257_1, n11256_0, n11227_0, n11226_0}), .out(n999), .config_in(config_chain[1034:1032]), .config_rst(config_rst)); 
mux6 mux_345 (.in({n12713_1, n12712_0, n12705_1, n12704_0, n12637_0, n12636_1}), .out(n1000), .config_in(config_chain[1037:1035]), .config_rst(config_rst)); 
mux6 mux_346 (.in({n11027_0, n11026_0, n10989_0, n10988_0, n10957_0, n10956_0}), .out(n1001), .config_in(config_chain[1040:1038]), .config_rst(config_rst)); 
mux6 mux_347 (.in({n12443_1, n12442_0, n12431_0, n12430_0, n12419_0, n12418_0/**/}), .out(n1002), .config_in(config_chain[1043:1041]), .config_rst(config_rst)); 
mux6 mux_348 (.in({n11291_0, n11290_0, n11259_0, n11258_0, n11221_0, n11220_0}), .out(n1003), .config_in(config_chain[1046:1044]), .config_rst(config_rst)); 
mux6 mux_349 (.in({n12657_0, n12656_0, n12653_0, n12652_1/**/, n12645_0, n12644_1}), .out(n1004), .config_in(config_chain[1049:1047]), .config_rst(config_rst)); 
mux6 mux_350 (.in({n11021_0, n11020_0, n10991_1, n10990_0, n10959_1, n10958_0}), .out(n1005), .config_in(config_chain[1052:1050]), .config_rst(config_rst)); 
mux6 mux_351 (.in({n12451_1, n12450_0, n12439_0, n12438_0, n12383_0, n12382_1}), .out(n1006), .config_in(config_chain[1055:1053]), .config_rst(config_rst)); 
mux6 mux_352 (.in({n11285_0/**/, n11284_0, n11253_0, n11252_0, n11223_0, n11222_0}), .out(n1007), .config_in(config_chain[1058:1056]), .config_rst(config_rst)); 
mux6 mux_353 (.in({n12685_0, n12684_0, n12677_0/**/, n12676_0, n12673_0, n12672_0}), .out(n1008), .config_in(config_chain[1061:1059]), .config_rst(config_rst)); 
mux6 mux_354 (.in({n11023_1, n11022_0, n10993_0, n10992_0, n10971_0, n10970_0}), .out(n1009), .config_in(config_chain[1064:1062]), .config_rst(config_rst)); 
mux6 mux_355 (.in({n12405_0, n12404_0, n12399_0, n12398_1, n12391_0, n12390_1}), .out(n1010), .config_in(config_chain[1067:1065]), .config_rst(config_rst)); 
mux6 mux_356 (.in({n11287_0, n11286_0, n11265_1, n11264_0, n11233_1, n11232_0}), .out(n1011), .config_in(config_chain[1070:1068]), .config_rst(config_rst)); 
mux6 mux_357 (.in({n12707_1, n12706_0, n12693_0, n12692_0, n12639_0, n12638_1/**/}), .out(n1012), .config_in(config_chain[1073:1071]), .config_rst(config_rst)); 
mux6 mux_358 (.in({n11025_0, n11024_0, n11003_0, n11002_0, n10965_0, n10964_0}), .out(n1013), .config_in(config_chain[1076:1074]), .config_rst(config_rst)); 
mux6 mux_359 (.in({n12425_0, n12424_0, n12421_0/**/, n12420_0, n12413_0, n12412_0}), .out(n1014), .config_in(config_chain[1079:1077]), .config_rst(config_rst)); 
mux6 mux_360 (.in({n11297_1/**/, n11296_0, n11267_0, n11266_0, n11235_0, n11234_0}), .out(n1015), .config_in(config_chain[1082:1080]), .config_rst(config_rst)); 
mux6 mux_361 (.in({n12715_1/**/, n12714_0, n12659_0, n12658_0, n12647_0, n12646_1}), .out(n1016), .config_in(config_chain[1085:1083]), .config_rst(config_rst)); 
mux6 mux_362 (.in({n11029_0, n11028_0, n10997_0/**/, n10996_0, n10967_1, n10966_0}), .out(n1017), .config_in(config_chain[1088:1086]), .config_rst(config_rst)); 
mux6 mux_363 (.in({n12453_1, n12452_0/**/, n12445_1, n12444_0, n12441_0, n12440_0}), .out(n1018), .config_in(config_chain[1091:1089]), .config_rst(config_rst)); 
mux6 mux_364 (.in({n11299_0, n11298_0, n11261_0, n11260_0/**/, n11231_0, n11230_0}), .out(n1019), .config_in(config_chain[1094:1092]), .config_rst(config_rst)); 
mux6 mux_365 (.in({n12679_0, n12678_0, n12675_0, n12674_0, n12667_0, n12666_0}), .out(n1020), .config_in(config_chain[1097:1095]), .config_rst(config_rst)); 
mux6 mux_366 (.in({n11031_1, n11030_0, n11001_0, n11000_0, n10969_0/**/, n10968_0}), .out(n1021), .config_in(config_chain[1100:1098]), .config_rst(config_rst)); 
mux6 mux_367 (.in({n12461_1, n12460_0/**/, n12393_0, n12392_1, n12385_0, n12384_1}), .out(n1022), .config_in(config_chain[1103:1101]), .config_rst(config_rst)); 
mux6 mux_368 (.in({n11293_0, n11292_0/**/, n11263_0, n11262_0, n11241_1, n11240_0}), .out(n1023), .config_in(config_chain[1106:1104]), .config_rst(config_rst)); 
mux6 mux_369 (.in({n12701_1, n12700_0, n12695_0/**/, n12694_0, n12687_0, n12686_0}), .out(n1024), .config_in(config_chain[1109:1107]), .config_rst(config_rst)); 
mux6 mux_370 (.in({n11033_0, n11032_0, n11011_0, n11010_0, n10979_0, n10978_0}), .out(n1025), .config_in(config_chain[1112:1110]), .config_rst(config_rst)); 
mux6 mux_371 (.in({n12427_0/**/, n12426_0, n12415_0, n12414_0, n12401_0, n12400_1}), .out(n1026), .config_in(config_chain[1115:1113]), .config_rst(config_rst)); 
mux6 mux_372 (.in({n11301_0, n11300_0, n11273_1, n11272_0, n11243_0/**/, n11242_0}), .out(n1027), .config_in(config_chain[1118:1116]), .config_rst(config_rst)); 
mux6 mux_373 (.in({n12649_0, n12648_1, n12641_0, n12640_1, n12605_0, n12604_1}), .out(n1028), .config_in(config_chain[1121:1119]), .config_rst(config_rst)); 
mux6 mux_374 (.in({n11039_1, n11038_0, n11005_0, n11004_0, n10975_1, n10974_0}), .out(n1029), .config_in(config_chain[1124:1122]), .config_rst(config_rst)); 
mux6 mux_375 (.in({n12447_1, n12446_0, n12435_0, n12434_0, n12353_1, n12352_1}), .out(n1030), .config_in(config_chain[1127:1125]), .config_rst(config_rst)); 
mux6 mux_376 (.in({n11303_0, n11302_0, n11275_0/**/, n11274_0, n11237_0, n11236_0}), .out(n1031), .config_in(config_chain[1130:1128]), .config_rst(config_rst)); 
mux6 mux_377 (.in({n12669_0, n12668_0, n12661_0, n12660_0, n12607_0/**/, n12606_1}), .out(n1032), .config_in(config_chain[1133:1131]), .config_rst(config_rst)); 
mux6 mux_378 (.in({n11041_1, n11040_0, n11007_1/**/, n11006_0, n10977_0, n10976_0}), .out(n1033), .config_in(config_chain[1136:1134]), .config_rst(config_rst)); 
mux6 mux_379 (.in({n12455_1, n12454_0, n12387_0, n12386_1, n12357_1, n12356_1}), .out(n1034), .config_in(config_chain[1139:1137]), .config_rst(config_rst)); 
mux6 mux_380 (.in({n11305_1, n11304_0, n11271_0, n11270_0, n11239_0, n11238_0/**/}), .out(n1035), .config_in(config_chain[1142:1140]), .config_rst(config_rst)); 
mux6 mux_381 (.in({n12703_1, n12702_0, n12689_0, n12688_0, n12609_1, n12608_1}), .out(n1036), .config_in(config_chain[1145:1143]), .config_rst(config_rst)); 
mux6 mux_382 (.in({n11045_2, n11044_0, n11009_0, n11008_0, n10987_0, n10986_0}), .out(n1037), .config_in(config_chain[1148:1146]), .config_rst(config_rst)); 
mux6 mux_383 (.in({n12417_0, n12416_0, n12409_0, n12408_0, n12359_1, n12358_1}), .out(n1038), .config_in(config_chain[1151:1149]), .config_rst(config_rst)); 
mux6 mux_384 (.in({n11307_1, n11306_0, n11281_1, n11280_0, n11249_1, n11248_0/**/}), .out(n1039), .config_in(config_chain[1154:1152]), .config_rst(config_rst)); 
mux6 mux_385 (.in({n12711_1, n12710_0, n12643_0/**/, n12642_1, n12611_1, n12610_1}), .out(n1040), .config_in(config_chain[1157:1155]), .config_rst(config_rst)); 
mux6 mux_386 (.in({n11047_2, n11046_0, n11019_0, n11018_0/**/, n10981_0, n10980_0}), .out(n1041), .config_in(config_chain[1160:1158]), .config_rst(config_rst)); 
mux6 mux_387 (.in({n12437_0/**/, n12436_0, n12429_0, n12428_0, n12361_1, n12360_1}), .out(n1042), .config_in(config_chain[1163:1161]), .config_rst(config_rst)); 
mux6 mux_388 (.in({n11309_1, n11308_0, n11283_0/**/, n11282_0, n11245_0, n11244_0}), .out(n1043), .config_in(config_chain[1166:1164]), .config_rst(config_rst)); 
mux6 mux_389 (.in({n12663_0, n12662_0, n12651_0, n12650_1, n12615_1, n12614_1}), .out(n1044), .config_in(config_chain[1169:1167]), .config_rst(config_rst)); 
mux6 mux_390 (.in({n11037_0, n11036_0, n11015_1, n11014_0, n10983_1, n10982_0}), .out(n1045), .config_in(config_chain[1172:1170]), .config_rst(config_rst)); 
mux6 mux_391 (.in({n12457_1, n12456_0/**/, n12389_0, n12388_1, n12351_0, n12350_1}), .out(n1046), .config_in(config_chain[1175:1173]), .config_rst(config_rst)); 
mux6 mux_392 (.in({n11547_1, n11546_0, n11509_0, n11508_0, n11487_0, n11486_0}), .out(n1093), .config_in(config_chain[1178:1176]), .config_rst(config_rst)); 
mux6 mux_393 (.in({n12731_0, n12730_0, n12677_0, n12676_0, n12663_0, n12662_1}), .out(n1094), .config_in(config_chain[1181:1179]), .config_rst(config_rst)); 
mux6 mux_394 (.in({n11279_0, n11278_0, n11247_0, n11246_0, n11225_1, n11224_0}), .out(n1095), .config_in(config_chain[1184:1182]), .config_rst(config_rst)); 
mux6 mux_395 (.in({n12471_0, n12470_0, n12463_0, n12462_0, n12457_0, n12456_0}), .out(n1096), .config_in(config_chain[1187:1185]), .config_rst(config_rst)); 
mux6 mux_396 (.in({n11541_0, n11540_0, n11519_0, n11518_0, n11489_0, n11488_0}), .out(n1097), .config_in(config_chain[1190:1188]), .config_rst(config_rst)); 
mux6 mux_397 (.in({n12697_0, n12696_0, n12693_0, n12692_0, n12685_0, n12684_0}), .out(n1098), .config_in(config_chain[1193:1191]), .config_rst(config_rst)); 
mux6 mux_398 (.in({n11289_1, n11288_0, n11259_0/**/, n11258_0, n11227_0, n11226_0}), .out(n1099), .config_in(config_chain[1196:1194]), .config_rst(config_rst)); 
mux6 mux_399 (.in({n12479_0, n12478_0, n12423_0, n12422_0, n12411_0, n12410_1/**/}), .out(n1100), .config_in(config_chain[1199:1197]), .config_rst(config_rst)); 
mux6 mux_400 (.in({n11553_0, n11552_0, n11521_0, n11520_0, n11491_1, n11490_0}), .out(n1101), .config_in(config_chain[1202:1200]), .config_rst(config_rst)); 
mux6 mux_401 (.in({n12717_0, n12716_0, n12713_0, n12712_0, n12705_0, n12704_0}), .out(n1102), .config_in(config_chain[1205:1203]), .config_rst(config_rst)); 
mux6 mux_402 (.in({n11291_0, n11290_0, n11253_0, n11252_0, n11221_0, n11220_0}), .out(n1103), .config_in(config_chain[1208:1206]), .config_rst(config_rst)); 
mux6 mux_403 (.in({n12443_0, n12442_0, n12431_0, n12430_0, n12419_0, n12418_1}), .out(n1104), .config_in(config_chain[1211:1209]), .config_rst(config_rst)); 
mux6 mux_404 (.in({n11555_1, n11554_0, n11523_1, n11522_0, n11485_0, n11484_0}), .out(n1105), .config_in(config_chain[1214:1212]), .config_rst(config_rst)); 
mux6 mux_405 (.in({n12733_0, n12732_0, n12665_0, n12664_1, n12657_0, n12656_1/**/}), .out(n1106), .config_in(config_chain[1217:1215]), .config_rst(config_rst)); 
mux6 mux_406 (.in({n11285_0, n11284_0, n11255_0, n11254_0, n11233_1, n11232_0}), .out(n1107), .config_in(config_chain[1220:1218]), .config_rst(config_rst)); 
mux6 mux_407 (.in({n12465_0, n12464_0, n12459_0, n12458_0, n12451_0, n12450_0}), .out(n1108), .config_in(config_chain[1223:1221]), .config_rst(config_rst)); 
mux6 mux_408 (.in({n11549_0/**/, n11548_0, n11527_0, n11526_0, n11495_0, n11494_0}), .out(n1109), .config_in(config_chain[1226:1224]), .config_rst(config_rst)); 
mux6 mux_409 (.in({n12699_0, n12698_0, n12687_0/**/, n12686_0, n12673_0, n12672_1}), .out(n1110), .config_in(config_chain[1229:1227]), .config_rst(config_rst)); 
mux6 mux_410 (.in({n11287_0, n11286_0, n11265_1, n11264_0, n11235_0/**/, n11234_0}), .out(n1111), .config_in(config_chain[1232:1230]), .config_rst(config_rst)); 
mux6 mux_411 (.in({n12481_0, n12480_0, n12473_0, n12472_0, n12405_0, n12404_1}), .out(n1112), .config_in(config_chain[1235:1233]), .config_rst(config_rst)); 
mux6 mux_412 (.in({n11559_0, n11558_0, n11529_0, n11528_0, n11497_0, n11496_0}), .out(n1113), .config_in(config_chain[1238:1236]), .config_rst(config_rst)); 
mux6 mux_413 (.in({n12719_0, n12718_0, n12707_0, n12706_0, n12695_0, n12694_0}), .out(n1114), .config_in(config_chain[1241:1239]), .config_rst(config_rst)); 
mux6 mux_414 (.in({n11299_0, n11298_0, n11267_0, n11266_0, n11229_0, n11228_0}), .out(n1115), .config_in(config_chain[1244:1242]), .config_rst(config_rst)); 
mux6 mux_415 (.in({n12433_0, n12432_0, n12425_0, n12424_0, n12421_0, n12420_1}), .out(n1116), .config_in(config_chain[1247:1245]), .config_rst(config_rst)); 
mux6 mux_416 (.in({n11561_0, n11560_0, n11531_1, n11530_0, n11493_0, n11492_0}), .out(n1117), .config_in(config_chain[1250:1248]), .config_rst(config_rst)); 
mux6 mux_417 (.in({n12735_0, n12734_0, n12727_0, n12726_0, n12659_0, n12658_1/**/}), .out(n1118), .config_in(config_chain[1253:1251]), .config_rst(config_rst)); 
mux6 mux_418 (.in({n11293_0/**/, n11292_0, n11263_0, n11262_0, n11231_0, n11230_0}), .out(n1119), .config_in(config_chain[1256:1254]), .config_rst(config_rst)); 
mux6 mux_419 (.in({n12453_0, n12452_0, n12445_0, n12444_0, n12441_0/**/, n12440_0}), .out(n1120), .config_in(config_chain[1259:1257]), .config_rst(config_rst)); 
mux6 mux_420 (.in({n11563_1/**/, n11562_0, n11525_0, n11524_0, n11503_0, n11502_0}), .out(n1121), .config_in(config_chain[1262:1260]), .config_rst(config_rst)); 
mux6 mux_421 (.in({n12681_0, n12680_0, n12675_0, n12674_1, n12667_0, n12666_1}), .out(n1122), .config_in(config_chain[1265:1263]), .config_rst(config_rst)); 
mux6 mux_422 (.in({n11295_0, n11294_0, n11273_1, n11272_0, n11241_1/**/, n11240_0}), .out(n1123), .config_in(config_chain[1268:1266]), .config_rst(config_rst)); 
mux6 mux_423 (.in({n12475_0, n12474_0, n12461_0, n12460_0, n12407_0, n12406_1}), .out(n1124), .config_in(config_chain[1271:1269]), .config_rst(config_rst)); 
mux6 mux_424 (.in({n11575_1, n11574_0, n11535_0, n11534_0, n11505_0, n11504_0/**/}), .out(n1125), .config_in(config_chain[1274:1272]), .config_rst(config_rst)); 
mux6 mux_425 (.in({n12709_0, n12708_0, n12701_0, n12700_0, n12615_0, n12614_2}), .out(n1126), .config_in(config_chain[1277:1275]), .config_rst(config_rst)); 
mux6 mux_426 (.in({n11301_0, n11300_0, n11275_0, n11274_0, n11237_0, n11236_0}), .out(n1127), .config_in(config_chain[1280:1278]), .config_rst(config_rst)); 
mux6 mux_427 (.in({n12427_0, n12426_0, n12415_0, n12414_1, n12351_0, n12350_2}), .out(n1128), .config_in(config_chain[1283:1281]), .config_rst(config_rst)); 
mux6 mux_428 (.in({n11565_0, n11564_0, n11537_0, n11536_0, n11507_1/**/, n11506_0}), .out(n1129), .config_in(config_chain[1286:1284]), .config_rst(config_rst)); 
mux6 mux_429 (.in({n12729_0, n12728_0, n12721_0, n12720_0, n12605_0, n12604_2}), .out(n1130), .config_in(config_chain[1289:1287]), .config_rst(config_rst)); 
mux6 mux_430 (.in({n11303_0/**/, n11302_0, n11269_0, n11268_0, n11239_0, n11238_0}), .out(n1131), .config_in(config_chain[1292:1290]), .config_rst(config_rst)); 
mux6 mux_431 (.in({n12447_0, n12446_0, n12435_0/**/, n12434_0, n12355_0, n12354_2}), .out(n1132), .config_in(config_chain[1295:1293]), .config_rst(config_rst)); 
mux6 mux_432 (.in({n11567_0, n11566_0, n11533_0, n11532_0, n11501_0/**/, n11500_0}), .out(n1133), .config_in(config_chain[1298:1296]), .config_rst(config_rst)); 
mux6 mux_433 (.in({n12683_0, n12682_0, n12669_0, n12668_1/**/, n12607_0, n12606_2}), .out(n1134), .config_in(config_chain[1301:1299]), .config_rst(config_rst)); 
mux6 mux_434 (.in({n11307_1, n11306_0, n11271_0, n11270_0, n11249_1, n11248_0}), .out(n1135), .config_in(config_chain[1304:1302]), .config_rst(config_rst)); 
mux6 mux_435 (.in({n12477_0, n12476_0, n12469_0, n12468_0/**/, n12357_0, n12356_2}), .out(n1136), .config_in(config_chain[1307:1305]), .config_rst(config_rst)); 
mux6 mux_436 (.in({n11569_0, n11568_0, n11543_0, n11542_0, n11511_0/**/, n11510_0}), .out(n1137), .config_in(config_chain[1310:1308]), .config_rst(config_rst)); 
mux6 mux_437 (.in({n12703_0, n12702_0, n12691_0, n12690_0, n12609_0, n12608_2}), .out(n1138), .config_in(config_chain[1313:1311]), .config_rst(config_rst)); 
mux6 mux_438 (.in({n11309_1, n11308_0, n11281_1, n11280_0, n11251_0, n11250_0}), .out(n1139), .config_in(config_chain[1316:1314]), .config_rst(config_rst)); 
mux6 mux_439 (.in({n12417_0/**/, n12416_1, n12409_0, n12408_1, n12359_0, n12358_2}), .out(n1140), .config_in(config_chain[1319:1317]), .config_rst(config_rst)); 
mux6 mux_440 (.in({n11571_1, n11570_0, n11545_0, n11544_0, n11515_1, n11514_0}), .out(n1141), .config_in(config_chain[1322:1320]), .config_rst(config_rst)); 
mux6 mux_441 (.in({n12723_0, n12722_0, n12711_0, n12710_0, n12613_0, n12612_2}), .out(n1142), .config_in(config_chain[1325:1323]), .config_rst(config_rst)); 
mux6 mux_442 (.in({n11311_2, n11310_0, n11277_0, n11276_0, n11245_0, n11244_0}), .out(n1143), .config_in(config_chain[1328:1326]), .config_rst(config_rst)); 
mux6 mux_443 (.in({n12449_0, n12448_0, n12437_0, n12436_0, n12361_0, n12360_2}), .out(n1144), .config_in(config_chain[1331:1329]), .config_rst(config_rst)); 
mux6 mux_444 (.in({n11809_0, n11808_0, n11779_0, n11778_0, n11749_1, n11748_0}), .out(n1191), .config_in(config_chain[1334:1332]), .config_rst(config_rst)); 
mux6 mux_445 (.in({n12737_0, n12736_0, n12723_0, n12722_0, n12711_0, n12710_0}), .out(n1192), .config_in(config_chain[1337:1335]), .config_rst(config_rst)); 
mux6 mux_446 (.in({n11541_0, n11540_0, n11509_0, n11508_0, n11487_0, n11486_0}), .out(n1193), .config_in(config_chain[1340:1338]), .config_rst(config_rst)); 
mux6 mux_447 (.in({n12451_0, n12450_0, n12443_0, n12442_0, n12437_0, n12436_1}), .out(n1194), .config_in(config_chain[1343:1341]), .config_rst(config_rst)); 
mux6 mux_448 (.in({n11811_0, n11810_0, n11781_1, n11780_0, n11751_0, n11750_0}), .out(n1195), .config_in(config_chain[1346:1344]), .config_rst(config_rst)); 
mux6 mux_449 (.in({n12753_0, n12752_0, n12745_0/**/, n12744_0, n12677_0, n12676_1}), .out(n1196), .config_in(config_chain[1349:1347]), .config_rst(config_rst)); 
mux6 mux_450 (.in({n11551_0, n11550_0, n11521_0, n11520_0, n11489_0, n11488_0}), .out(n1197), .config_in(config_chain[1352:1350]), .config_rst(config_rst)); 
mux6 mux_451 (.in({n12483_0, n12482_0, n12471_0, n12470_0, n12459_0, n12458_0}), .out(n1198), .config_in(config_chain[1355:1353]), .config_rst(config_rst)); 
mux6 mux_452 (.in({n11815_0, n11814_0, n11783_0, n11782_0, n11753_0, n11752_0}), .out(n1199), .config_in(config_chain[1358:1356]), .config_rst(config_rst)); 
mux6 mux_453 (.in({n12697_0, n12696_0, n12693_0, n12692_1, n12685_0, n12684_1/**/}), .out(n1200), .config_in(config_chain[1361:1359]), .config_rst(config_rst)); 
mux6 mux_454 (.in({n11553_0, n11552_0, n11523_1, n11522_0, n11491_1, n11490_0}), .out(n1201), .config_in(config_chain[1364:1362]), .config_rst(config_rst)); 
mux6 mux_455 (.in({n12491_0, n12490_0, n12479_0, n12478_0, n12423_0, n12422_1}), .out(n1202), .config_in(config_chain[1367:1365]), .config_rst(config_rst)); 
mux6 mux_456 (.in({n11817_0, n11816_0, n11785_0, n11784_0, n11755_0, n11754_0}), .out(n1203), .config_in(config_chain[1370:1368]), .config_rst(config_rst)); 
mux6 mux_457 (.in({n12725_0, n12724_0, n12717_0, n12716_0/**/, n12713_0, n12712_0}), .out(n1204), .config_in(config_chain[1373:1371]), .config_rst(config_rst)); 
mux6 mux_458 (.in({n11555_1, n11554_0/**/, n11517_0, n11516_0, n11495_0, n11494_0}), .out(n1205), .config_in(config_chain[1376:1374]), .config_rst(config_rst)); 
mux6 mux_459 (.in({n12445_0, n12444_0, n12439_0, n12438_1, n12431_0, n12430_1}), .out(n1206), .config_in(config_chain[1379:1377]), .config_rst(config_rst)); 
mux6 mux_460 (.in({n11819_0, n11818_0, n11789_1, n11788_0, n11757_1, n11756_0}), .out(n1207), .config_in(config_chain[1382:1380]), .config_rst(config_rst)); 
mux6 mux_461 (.in({n12747_0, n12746_0/**/, n12733_0, n12732_0, n12679_0, n12678_1}), .out(n1208), .config_in(config_chain[1385:1383]), .config_rst(config_rst)); 
mux6 mux_462 (.in({n11549_0/**/, n11548_0, n11527_0, n11526_0, n11497_0, n11496_0}), .out(n1209), .config_in(config_chain[1388:1386]), .config_rst(config_rst)); 
mux6 mux_463 (.in({n12465_0, n12464_0, n12461_0, n12460_0, n12453_0, n12452_0}), .out(n1210), .config_in(config_chain[1391:1389]), .config_rst(config_rst)); 
mux6 mux_464 (.in({n11821_1, n11820_0, n11791_0, n11790_0, n11759_0, n11758_0}), .out(n1211), .config_in(config_chain[1394:1392]), .config_rst(config_rst)); 
mux6 mux_465 (.in({n12755_0, n12754_0, n12699_0, n12698_0, n12687_0, n12686_1}), .out(n1212), .config_in(config_chain[1397:1395]), .config_rst(config_rst)); 
mux6 mux_466 (.in({n11561_0, n11560_0, n11529_0, n11528_0, n11499_1, n11498_0}), .out(n1213), .config_in(config_chain[1400:1398]), .config_rst(config_rst)); 
mux6 mux_467 (.in({n12493_0, n12492_0, n12485_0, n12484_0, n12481_0, n12480_0}), .out(n1214), .config_in(config_chain[1403:1401]), .config_rst(config_rst)); 
mux6 mux_468 (.in({n11823_0/**/, n11822_0, n11793_0, n11792_0, n11763_0, n11762_0}), .out(n1215), .config_in(config_chain[1406:1404]), .config_rst(config_rst)); 
mux6 mux_469 (.in({n12719_0, n12718_0, n12715_0/**/, n12714_0, n12707_0, n12706_0}), .out(n1216), .config_in(config_chain[1409:1407]), .config_rst(config_rst)); 
mux6 mux_470 (.in({n11563_1, n11562_0, n11525_0/**/, n11524_0, n11493_0, n11492_0}), .out(n1217), .config_in(config_chain[1412:1410]), .config_rst(config_rst)); 
mux6 mux_471 (.in({n12501_0, n12500_0, n12433_0, n12432_1, n12425_0, n12424_1/**/}), .out(n1218), .config_in(config_chain[1415:1413]), .config_rst(config_rst)); 
mux6 mux_472 (.in({n11825_0, n11824_0, n11795_0/**/, n11794_0, n11765_1, n11764_0}), .out(n1219), .config_in(config_chain[1418:1416]), .config_rst(config_rst)); 
mux6 mux_473 (.in({n12741_0, n12740_0, n12735_0, n12734_0, n12727_0, n12726_0}), .out(n1220), .config_in(config_chain[1421:1419]), .config_rst(config_rst)); 
mux6 mux_474 (.in({n11557_0, n11556_0, n11535_0/**/, n11534_0, n11503_0, n11502_0}), .out(n1221), .config_in(config_chain[1424:1422]), .config_rst(config_rst)); 
mux6 mux_475 (.in({n12467_0, n12466_0, n12455_0, n12454_0, n12441_0, n12440_1/**/}), .out(n1222), .config_in(config_chain[1427:1425]), .config_rst(config_rst)); 
mux6 mux_476 (.in({n11837_1, n11836_0, n11797_1, n11796_0, n11767_0, n11766_0}), .out(n1223), .config_in(config_chain[1430:1428]), .config_rst(config_rst)); 
mux6 mux_477 (.in({n12689_0, n12688_1, n12681_0, n12680_1/**/, n12613_0, n12612_2}), .out(n1224), .config_in(config_chain[1433:1431]), .config_rst(config_rst)); 
mux6 mux_478 (.in({n11575_1, n11574_0, n11537_0, n11536_0, n11507_1, n11506_0}), .out(n1225), .config_in(config_chain[1436:1434]), .config_rst(config_rst)); 
mux6 mux_479 (.in({n12487_0, n12486_0, n12475_0, n12474_0/**/, n12361_0, n12360_2}), .out(n1226), .config_in(config_chain[1439:1437]), .config_rst(config_rst)); 
mux6 mux_480 (.in({n11839_1, n11838_0, n11799_0, n11798_0, n11769_0, n11768_0}), .out(n1227), .config_in(config_chain[1442:1440]), .config_rst(config_rst)); 
mux6 mux_481 (.in({n12709_0, n12708_0/**/, n12701_0, n12700_0, n12615_0, n12614_2}), .out(n1228), .config_in(config_chain[1445:1443]), .config_rst(config_rst)); 
mux6 mux_482 (.in({n11565_0, n11564_0, n11539_1, n11538_0, n11501_0, n11500_0}), .out(n1229), .config_in(config_chain[1448:1446]), .config_rst(config_rst)); 
mux6 mux_483 (.in({n12495_0, n12494_0/**/, n12427_0, n12426_1, n12353_0, n12352_2}), .out(n1230), .config_in(config_chain[1451:1449]), .config_rst(config_rst)); 
mux6 mux_484 (.in({n11829_2, n11828_0, n11803_0, n11802_0, n11771_0, n11770_0}), .out(n1231), .config_in(config_chain[1454:1452]), .config_rst(config_rst)); 
mux6 mux_485 (.in({n12757_0, n12756_0, n12743_0, n12742_0/**/, n12729_0, n12728_0}), .out(n1232), .config_in(config_chain[1457:1455]), .config_rst(config_rst)); 
mux6 mux_486 (.in({n11569_0, n11568_0, n11533_0, n11532_0, n11511_0, n11510_0}), .out(n1233), .config_in(config_chain[1460:1458]), .config_rst(config_rst)); 
mux6 mux_487 (.in({n12457_0, n12456_0, n12449_0, n12448_0, n12355_0, n12354_2}), .out(n1234), .config_in(config_chain[1463:1461]), .config_rst(config_rst)); 
mux6 mux_488 (.in({n11831_0, n11830_0, n11805_1, n11804_0, n11773_1/**/, n11772_0}), .out(n1235), .config_in(config_chain[1466:1464]), .config_rst(config_rst)); 
mux6 mux_489 (.in({n12751_0, n12750_0, n12683_0, n12682_1, n12607_0, n12606_2}), .out(n1236), .config_in(config_chain[1469:1467]), .config_rst(config_rst)); 
mux6 mux_490 (.in({n11571_1, n11570_0, n11543_0, n11542_0, n11513_0, n11512_0}), .out(n1237), .config_in(config_chain[1472:1470]), .config_rst(config_rst)); 
mux6 mux_491 (.in({n12477_0, n12476_0, n12469_0, n12468_0, n12357_0, n12356_2}), .out(n1238), .config_in(config_chain[1475:1473]), .config_rst(config_rst)); 
mux6 mux_492 (.in({n11833_0, n11832_0, n11807_0, n11806_0, n11777_0/**/, n11776_0}), .out(n1239), .config_in(config_chain[1478:1476]), .config_rst(config_rst)); 
mux6 mux_493 (.in({n12703_0, n12702_0, n12691_0/**/, n12690_1, n12611_0, n12610_2}), .out(n1240), .config_in(config_chain[1481:1479]), .config_rst(config_rst)); 
mux6 mux_494 (.in({n11573_1, n11572_0, n11547_1, n11546_0, n11515_1, n11514_0}), .out(n1241), .config_in(config_chain[1484:1482]), .config_rst(config_rst)); 
mux6 mux_495 (.in({n12497_0, n12496_0, n12429_0, n12428_1/**/, n12359_0, n12358_2}), .out(n1242), .config_in(config_chain[1487:1485]), .config_rst(config_rst)); 
mux6 mux_496 (.in({n12069_1, n12068_0, n12039_0, n12038_0, n12017_0, n12016_0}), .out(n1289), .config_in(config_chain[1490:1488]), .config_rst(config_rst)); 
mux6 mux_497 (.in({n12773_0, n12772_0, n12717_0, n12716_0, n12703_0, n12702_1}), .out(n1290), .config_in(config_chain[1493:1491]), .config_rst(config_rst)); 
mux6 mux_498 (.in({n11811_0, n11810_0, n11779_0, n11778_0, n11749_1, n11748_0}), .out(n1291), .config_in(config_chain[1496:1494]), .config_rst(config_rst)); 
mux6 mux_499 (.in({n12511_0, n12510_0, n12503_0, n12502_0, n12497_0, n12496_0}), .out(n1292), .config_in(config_chain[1499:1497]), .config_rst(config_rst)); 
mux6 mux_500 (.in({n12071_0, n12070_0, n12049_0, n12048_0, n12011_0, n12010_0}), .out(n1293), .config_in(config_chain[1502:1500]), .config_rst(config_rst)); 
mux6 mux_501 (.in({n12737_0, n12736_0, n12733_0, n12732_0, n12725_0, n12724_0}), .out(n1294), .config_in(config_chain[1505:1503]), .config_rst(config_rst)); 
mux6 mux_502 (.in({n11813_1, n11812_0, n11783_0, n11782_0, n11751_0, n11750_0}), .out(n1295), .config_in(config_chain[1508:1506]), .config_rst(config_rst)); 
mux6 mux_503 (.in({n12519_0, n12518_0, n12463_0, n12462_0, n12451_0, n12450_1}), .out(n1296), .config_in(config_chain[1511:1509]), .config_rst(config_rst)); 
mux6 mux_504 (.in({n12075_0, n12074_0, n12043_0, n12042_0, n12013_1, n12012_0}), .out(n1297), .config_in(config_chain[1514:1512]), .config_rst(config_rst)); 
mux6 mux_505 (.in({n12759_0, n12758_0, n12753_0, n12752_0, n12745_0, n12744_0}), .out(n1298), .config_in(config_chain[1517:1515]), .config_rst(config_rst)); 
mux6 mux_506 (.in({n11815_0, n11814_0, n11785_0, n11784_0, n11753_0, n11752_0}), .out(n1299), .config_in(config_chain[1520:1518]), .config_rst(config_rst)); 
mux6 mux_507 (.in({n12483_0, n12482_0, n12471_0, n12470_0, n12459_0, n12458_1}), .out(n1300), .config_in(config_chain[1523:1521]), .config_rst(config_rst)); 
mux6 mux_508 (.in({n12077_1, n12076_0, n12045_1, n12044_0, n12015_0, n12014_0}), .out(n1301), .config_in(config_chain[1526:1524]), .config_rst(config_rst)); 
mux6 mux_509 (.in({n12775_0, n12774_0, n12705_0, n12704_1, n12697_0, n12696_1}), .out(n1302), .config_in(config_chain[1529:1527]), .config_rst(config_rst)); 
mux6 mux_510 (.in({n11817_0, n11816_0, n11787_0, n11786_0, n11757_1, n11756_0}), .out(n1303), .config_in(config_chain[1532:1530]), .config_rst(config_rst)); 
mux6 mux_511 (.in({n12505_0, n12504_0, n12499_0, n12498_0, n12491_0, n12490_0}), .out(n1304), .config_in(config_chain[1535:1533]), .config_rst(config_rst)); 
mux6 mux_512 (.in({n12079_0, n12078_0, n12057_0, n12056_0, n12025_0, n12024_0}), .out(n1305), .config_in(config_chain[1538:1536]), .config_rst(config_rst)); 
mux6 mux_513 (.in({n12739_0, n12738_0, n12727_0, n12726_0, n12713_0, n12712_1}), .out(n1306), .config_in(config_chain[1541:1539]), .config_rst(config_rst)); 
mux6 mux_514 (.in({n11819_0, n11818_0, n11789_1, n11788_0, n11759_0, n11758_0}), .out(n1307), .config_in(config_chain[1544:1542]), .config_rst(config_rst)); 
mux6 mux_515 (.in({n12521_0, n12520_0, n12513_0, n12512_0, n12445_0, n12444_1}), .out(n1308), .config_in(config_chain[1547:1545]), .config_rst(config_rst)); 
mux6 mux_516 (.in({n12089_0, n12088_0, n12051_0, n12050_0, n12019_0, n12018_0}), .out(n1309), .config_in(config_chain[1550:1548]), .config_rst(config_rst)); 
mux6 mux_517 (.in({n12761_0, n12760_0, n12747_0, n12746_0, n12735_0, n12734_0}), .out(n1310), .config_in(config_chain[1553:1551]), .config_rst(config_rst)); 
mux6 mux_518 (.in({n11823_0, n11822_0, n11791_0, n11790_0, n11761_0, n11760_0}), .out(n1311), .config_in(config_chain[1556:1554]), .config_rst(config_rst)); 
mux6 mux_519 (.in({n12473_0, n12472_0, n12465_0, n12464_0, n12461_0, n12460_1}), .out(n1312), .config_in(config_chain[1559:1557]), .config_rst(config_rst)); 
mux6 mux_520 (.in({n12083_0, n12082_0, n12053_1, n12052_0, n12023_0, n12022_0}), .out(n1313), .config_in(config_chain[1562:1560]), .config_rst(config_rst)); 
mux6 mux_521 (.in({n12777_0, n12776_0, n12769_0, n12768_0, n12699_0, n12698_1}), .out(n1314), .config_in(config_chain[1565:1563]), .config_rst(config_rst)); 
mux6 mux_522 (.in({n11825_0, n11824_0, n11795_0, n11794_0, n11763_0, n11762_0}), .out(n1315), .config_in(config_chain[1568:1566]), .config_rst(config_rst)); 
mux6 mux_523 (.in({n12493_0, n12492_0, n12485_0, n12484_0, n12481_0, n12480_0}), .out(n1316), .config_in(config_chain[1571:1569]), .config_rst(config_rst)); 
mux6 mux_524 (.in({n12085_1, n12084_0, n12055_0, n12054_0, n12033_0, n12032_0}), .out(n1317), .config_in(config_chain[1574:1572]), .config_rst(config_rst)); 
mux6 mux_525 (.in({n12721_0, n12720_0, n12715_0, n12714_1, n12707_0, n12706_1}), .out(n1318), .config_in(config_chain[1577:1575]), .config_rst(config_rst)); 
mux6 mux_526 (.in({n11827_0, n11826_0, n11797_1, n11796_0, n11765_1, n11764_0}), .out(n1319), .config_in(config_chain[1580:1578]), .config_rst(config_rst)); 
mux6 mux_527 (.in({n12515_0, n12514_0, n12501_0, n12500_0, n12447_0, n12446_1}), .out(n1320), .config_in(config_chain[1583:1581]), .config_rst(config_rst)); 
mux6 mux_528 (.in({n12097_0, n12096_0, n12065_0, n12064_0, n12027_0, n12026_0}), .out(n1321), .config_in(config_chain[1586:1584]), .config_rst(config_rst)); 
mux6 mux_529 (.in({n12749_0, n12748_0, n12741_0, n12740_0, n12611_0, n12610_2}), .out(n1322), .config_in(config_chain[1589:1587]), .config_rst(config_rst)); 
mux6 mux_530 (.in({n11837_1, n11836_0, n11799_0, n11798_0, n11769_0, n11768_0}), .out(n1323), .config_in(config_chain[1592:1590]), .config_rst(config_rst)); 
mux6 mux_531 (.in({n12467_0, n12466_0, n12455_0, n12454_1, n12359_0, n12358_2}), .out(n1324), .config_in(config_chain[1595:1593]), .config_rst(config_rst)); 
mux6 mux_532 (.in({n12099_0, n12098_0, n12059_0, n12058_0, n12029_1, n12028_0}), .out(n1325), .config_in(config_chain[1598:1596]), .config_rst(config_rst)); 
mux6 mux_533 (.in({n12771_0, n12770_0, n12763_0, n12762_0, n12613_0, n12612_2}), .out(n1326), .config_in(config_chain[1601:1599]), .config_rst(config_rst)); 
mux6 mux_534 (.in({n11839_1, n11838_0, n11801_0, n11800_0, n11771_0, n11770_0}), .out(n1327), .config_in(config_chain[1604:1602]), .config_rst(config_rst)); 
mux6 mux_535 (.in({n12523_0, n12522_0, n12487_0, n12486_0, n12475_0, n12474_0}), .out(n1328), .config_in(config_chain[1607:1605]), .config_rst(config_rst)); 
mux6 mux_536 (.in({n12101_1, n12100_0, n12063_0, n12062_0, n12031_0, n12030_0}), .out(n1329), .config_in(config_chain[1610:1608]), .config_rst(config_rst)); 
mux6 mux_537 (.in({n12723_0, n12722_0, n12709_0, n12708_1, n12615_0, n12614_2}), .out(n1330), .config_in(config_chain[1613:1611]), .config_rst(config_rst)); 
mux6 mux_538 (.in({n11831_0, n11830_0, n11803_0, n11802_0, n11773_1, n11772_0}), .out(n1331), .config_in(config_chain[1616:1614]), .config_rst(config_rst)); 
mux6 mux_539 (.in({n12517_0, n12516_0, n12509_0, n12508_0, n12353_0, n12352_2}), .out(n1332), .config_in(config_chain[1619:1617]), .config_rst(config_rst)); 
mux6 mux_540 (.in({n12091_2, n12090_0, n12073_0, n12072_0, n12041_0, n12040_0}), .out(n1333), .config_in(config_chain[1622:1620]), .config_rst(config_rst)); 
mux6 mux_541 (.in({n12757_0, n12756_0, n12743_0, n12742_0, n12731_0, n12730_0}), .out(n1334), .config_in(config_chain[1625:1623]), .config_rst(config_rst)); 
mux6 mux_542 (.in({n11833_0, n11832_0, n11805_1, n11804_0, n11775_0, n11774_0}), .out(n1335), .config_in(config_chain[1628:1626]), .config_rst(config_rst)); 
mux6 mux_543 (.in({n12457_0, n12456_1, n12449_0, n12448_1, n12355_0, n12354_2}), .out(n1336), .config_in(config_chain[1631:1629]), .config_rst(config_rst)); 
mux6 mux_544 (.in({n12093_2, n12092_0, n12067_0, n12066_0, n12037_1, n12036_0}), .out(n1337), .config_in(config_chain[1634:1632]), .config_rst(config_rst)); 
mux6 mux_545 (.in({n12765_0, n12764_0, n12751_0, n12750_0, n12609_0, n12608_2}), .out(n1338), .config_in(config_chain[1637:1635]), .config_rst(config_rst)); 
mux6 mux_546 (.in({n11835_0, n11834_0, n11809_0, n11808_0, n11777_0, n11776_0}), .out(n1339), .config_in(config_chain[1640:1638]), .config_rst(config_rst)); 
mux6 mux_547 (.in({n12489_0, n12488_0, n12477_0, n12476_0, n12357_0, n12356_2}), .out(n1340), .config_in(config_chain[1643:1641]), .config_rst(config_rst)); 
mux6 mux_548 (.in({n12071_0, n12070_0, n12049_0, n12048_0, n12017_0, n12016_0}), .out(n1386), .config_in(config_chain[1646:1644]), .config_rst(config_rst)); 
mux6 mux_549 (.in({n12075_0, n12074_0, n12045_1, n12044_0, n12013_1, n12012_0}), .out(n1389), .config_in(config_chain[1649:1647]), .config_rst(config_rst)); 
mux6 mux_550 (.in({n12079_0, n12078_0, n12057_0, n12056_0, n12025_0, n12024_0}), .out(n1392), .config_in(config_chain[1652:1650]), .config_rst(config_rst)); 
mux6 mux_551 (.in({n12083_0, n12082_0, n12053_1, n12052_0, n12021_1, n12020_0}), .out(n1395), .config_in(config_chain[1655:1653]), .config_rst(config_rst)); 
mux6 mux_552 (.in({n12087_0, n12086_0, n12055_0, n12054_0, n12033_0, n12032_0}), .out(n1398), .config_in(config_chain[1658:1656]), .config_rst(config_rst)); 
mux6 mux_553 (.in({n12099_0, n12098_0, n12059_0, n12058_0, n12029_1, n12028_0}), .out(n1401), .config_in(config_chain[1661:1659]), .config_rst(config_rst)); 
mux6 mux_554 (.in({n12091_2, n12090_0, n12063_0, n12062_0, n12041_0, n12040_0}), .out(n1404), .config_in(config_chain[1664:1662]), .config_rst(config_rst)); 
mux6 mux_555 (.in({n12095_0, n12094_0, n12067_0, n12066_0, n12037_1, n12036_0}), .out(n1407), .config_in(config_chain[1667:1665]), .config_rst(config_rst)); 
mux6 mux_556 (.in({n9773_1, n9772_0, n9695_0, n9694_0, n9673_0, n9672_0}), .out(n1434), .config_in(config_chain[1670:1668]), .config_rst(config_rst)); 
mux6 mux_557 (.in({n9737_0, n9736_0, n9699_0, n9698_0, n9667_0, n9666_0}), .out(n1437), .config_in(config_chain[1673:1671]), .config_rst(config_rst)); 
mux6 mux_558 (.in({n9775_1, n9774_0, n9703_0, n9702_0, n9671_0, n9670_0}), .out(n1440), .config_in(config_chain[1676:1674]), .config_rst(config_rst)); 
mux6 mux_559 (.in({n9745_0, n9744_0, n9707_0, n9706_0, n9675_0, n9674_0}), .out(n1443), .config_in(config_chain[1679:1677]), .config_rst(config_rst)); 
mux6 mux_560 (.in({n9777_1, n9776_0, n9711_0, n9710_0, n9679_0, n9678_0}), .out(n1446), .config_in(config_chain[1682:1680]), .config_rst(config_rst)); 
mux6 mux_561 (.in({n9757_2, n9756_0, n9721_0, n9720_0, n9683_0, n9682_0}), .out(n1449), .config_in(config_chain[1685:1683]), .config_rst(config_rst)); 
mux6 mux_562 (.in({n9771_1, n9770_0, n9749_2, n9748_0, n9687_0, n9686_0}), .out(n1452), .config_in(config_chain[1688:1686]), .config_rst(config_rst)); 
mux6 mux_563 (.in({n9753_2, n9752_0, n9729_0, n9728_0, n9691_0, n9690_0}), .out(n1455), .config_in(config_chain[1691:1689]), .config_rst(config_rst)); 
mux6 mux_564 (.in({n10013_1, n10012_0, n9977_0, n9976_0, n9947_0, n9946_0}), .out(n1483), .config_in(config_chain[1694:1692]), .config_rst(config_rst)); 
mux6 mux_565 (.in({n12837_0, n12836_0, n12807_0, n12806_0, n12785_1, n12784_0}), .out(n1484), .config_in(config_chain[1697:1695]), .config_rst(config_rst)); 
mux6 mux_566 (.in({n9727_0, n9726_0, n9695_0, n9694_0, n9673_0, n9672_0}), .out(n1485), .config_in(config_chain[1700:1698]), .config_rst(config_rst)); 
mux6 mux_567 (.in({n12585_0, n12584_0, n12563_0, n12562_0, n12531_0, n12530_0}), .out(n1486), .config_in(config_chain[1703:1701]), .config_rst(config_rst)); 
mux6 mux_568 (.in({n10021_1, n10020_0, n9979_0, n9978_0, n9927_0, n9926_0}), .out(n1487), .config_in(config_chain[1706:1704]), .config_rst(config_rst)); 
mux6 mux_569 (.in({n12849_1, n12848_0, n12817_1, n12816_0, n12787_0, n12786_0}), .out(n1488), .config_in(config_chain[1709:1707]), .config_rst(config_rst)); 
mux6 mux_570 (.in({n9737_0, n9736_0, n9699_0, n9698_0, n9667_0, n9666_0}), .out(n1489), .config_in(config_chain[1712:1710]), .config_rst(config_rst)); 
mux6 mux_571 (.in({n12595_0, n12594_0, n12557_0, n12556_0, n12527_1, n12526_0}), .out(n1490), .config_in(config_chain[1715:1713]), .config_rst(config_rst)); 
mux6 mux_572 (.in({n9991_0, n9990_0, n9959_0, n9958_0, n9921_0, n9920_0}), .out(n1491), .config_in(config_chain[1718:1716]), .config_rst(config_rst)); 
mux6 mux_573 (.in({n12851_0, n12850_0, n12819_0, n12818_0, n12781_0, n12780_0}), .out(n1492), .config_in(config_chain[1721:1719]), .config_rst(config_rst)); 
mux6 mux_574 (.in({n9767_1, n9766_0, n9759_1, n9758_0, n9731_0, n9730_0}), .out(n1493), .config_in(config_chain[1724:1722]), .config_rst(config_rst)); 
mux6 mux_575 (.in({n12589_0, n12588_0, n12559_1, n12558_0, n12529_0, n12528_0}), .out(n1494), .config_in(config_chain[1727:1725]), .config_rst(config_rst)); 
mux6 mux_576 (.in({n9985_0, n9984_0, n9953_0, n9952_0, n9923_0, n9922_0}), .out(n1495), .config_in(config_chain[1730:1728]), .config_rst(config_rst)); 
mux6 mux_577 (.in({n12845_0, n12844_0, n12815_0, n12814_0, n12783_0, n12782_0}), .out(n1496), .config_in(config_chain[1733:1731]), .config_rst(config_rst)); 
mux6 mux_578 (.in({n9775_1, n9774_0, n9703_0, n9702_0, n9681_0, n9680_0}), .out(n1497), .config_in(config_chain[1736:1734]), .config_rst(config_rst)); 
mux6 mux_579 (.in({n12593_0, n12592_0, n12561_0, n12560_0, n12539_0, n12538_0}), .out(n1498), .config_in(config_chain[1739:1737]), .config_rst(config_rst)); 
mux6 mux_580 (.in({n10023_1, n10022_0, n10015_1, n10014_0, n9987_0, n9986_0}), .out(n1499), .config_in(config_chain[1742:1740]), .config_rst(config_rst)); 
mux6 mux_581 (.in({n12847_0, n12846_0, n12825_1, n12824_0, n12795_0, n12794_0}), .out(n1500), .config_in(config_chain[1745:1743]), .config_rst(config_rst)); 
mux6 mux_582 (.in({n9735_0, n9734_0, n9713_0, n9712_0, n9675_0, n9674_0}), .out(n1501), .config_in(config_chain[1748:1746]), .config_rst(config_rst)); 
mux6 mux_583 (.in({n12603_0, n12602_0, n12571_0, n12570_0, n12533_0, n12532_0}), .out(n1502), .config_in(config_chain[1751:1749]), .config_rst(config_rst)); 
mux6 mux_584 (.in({n10031_1, n10030_0, n9967_0, n9966_0, n9935_0, n9934_0}), .out(n1503), .config_in(config_chain[1754:1752]), .config_rst(config_rst)); 
mux6 mux_585 (.in({n12857_1, n12856_0, n12827_0, n12826_0, n12789_0, n12788_0}), .out(n1504), .config_in(config_chain[1757:1755]), .config_rst(config_rst)); 
mux6 mux_586 (.in({n9761_1, n9760_0, n9739_0, n9738_0, n9707_0, n9706_0}), .out(n1505), .config_in(config_chain[1760:1758]), .config_rst(config_rst)); 
mux6 mux_587 (.in({n12597_0, n12596_0, n12567_1, n12566_0, n12535_1, n12534_0}), .out(n1506), .config_in(config_chain[1763:1761]), .config_rst(config_rst)); 
mux6 mux_588 (.in({n9999_0, n9998_0, n9961_0, n9960_0, n9931_0, n9930_0}), .out(n1507), .config_in(config_chain[1766:1764]), .config_rst(config_rst)); 
mux6 mux_589 (.in({n12853_0, n12852_0, n12821_0, n12820_0, n12791_0, n12790_0}), .out(n1508), .config_in(config_chain[1769:1767]), .config_rst(config_rst)); 
mux6 mux_590 (.in({n9777_1, n9776_0, n9711_0, n9710_0, n9679_0, n9678_0}), .out(n1509), .config_in(config_chain[1772:1770]), .config_rst(config_rst)); 
mux6 mux_591 (.in({n12599_1, n12598_0, n12569_0, n12568_0, n12537_0, n12536_0}), .out(n1510), .config_in(config_chain[1775:1773]), .config_rst(config_rst)); 
mux6 mux_592 (.in({n10017_1, n10016_0, n9993_0, n9992_0, n9963_0, n9962_0}), .out(n1511), .config_in(config_chain[1778:1776]), .config_rst(config_rst)); 
mux6 mux_593 (.in({n12855_0, n12854_0, n12823_0, n12822_0, n12801_1, n12800_0}), .out(n1512), .config_in(config_chain[1781:1779]), .config_rst(config_rst)); 
mux6 mux_594 (.in({n9743_0, n9742_0, n9721_0, n9720_0, n9689_0, n9688_0}), .out(n1513), .config_in(config_chain[1784:1782]), .config_rst(config_rst)); 
mux6 mux_595 (.in({n12601_0, n12600_0, n12579_0, n12578_0, n12541_0, n12540_0}), .out(n1514), .config_in(config_chain[1787:1785]), .config_rst(config_rst)); 
mux6 mux_596 (.in({n10025_1, n10024_0, n10009_2, n10008_0, n9943_0, n9942_0}), .out(n1515), .config_in(config_chain[1790:1788]), .config_rst(config_rst)); 
mux6 mux_597 (.in({n12869_2, n12868_0, n12835_0, n12834_0, n12803_0, n12802_0}), .out(n1516), .config_in(config_chain[1793:1791]), .config_rst(config_rst)); 
mux6 mux_598 (.in({n9763_1, n9762_0, n9757_2, n9756_0, n9715_0, n9714_0}), .out(n1517), .config_in(config_chain[1796:1794]), .config_rst(config_rst)); 
mux6 mux_599 (.in({n12615_2, n12614_0, n12573_0, n12572_0, n12543_1, n12542_0}), .out(n1518), .config_in(config_chain[1799:1797]), .config_rst(config_rst)); 
mux6 mux_600 (.in({n10011_2, n10010_0, n9975_0, n9974_0, n9937_0, n9936_0}), .out(n1519), .config_in(config_chain[1802:1800]), .config_rst(config_rst)); 
mux6 mux_601 (.in({n12871_2, n12870_0, n12829_0, n12828_0, n12797_0, n12796_0}), .out(n1520), .config_in(config_chain[1805:1803]), .config_rst(config_rst)); 
mux6 mux_602 (.in({n9771_1, n9770_0, n9747_2, n9746_0, n9687_0, n9686_0}), .out(n1521), .config_in(config_chain[1808:1806]), .config_rst(config_rst)); 
mux6 mux_603 (.in({n12607_2, n12606_0, n12575_1, n12574_0, n12545_0, n12544_0}), .out(n1522), .config_in(config_chain[1811:1809]), .config_rst(config_rst)); 
mux6 mux_604 (.in({n10001_1, n10000_0, n9971_0, n9970_0, n9939_0, n9938_0}), .out(n1523), .config_in(config_chain[1814:1812]), .config_rst(config_rst)); 
mux6 mux_605 (.in({n12861_1, n12860_0, n12831_0, n12830_0, n12809_1, n12808_0}), .out(n1524), .config_in(config_chain[1817:1815]), .config_rst(config_rst)); 
mux6 mux_606 (.in({n9751_2, n9750_0, n9719_0, n9718_0, n9697_0, n9696_0}), .out(n1525), .config_in(config_chain[1820:1818]), .config_rst(config_rst)); 
mux6 mux_607 (.in({n12609_2, n12608_0, n12587_0, n12586_0, n12555_0, n12554_0}), .out(n1526), .config_in(config_chain[1823:1821]), .config_rst(config_rst)); 
mux6 mux_608 (.in({n10027_1, n10026_0, n10019_1, n10018_0, n10003_2, n10002_0}), .out(n1527), .config_in(config_chain[1826:1824]), .config_rst(config_rst)); 
mux6 mux_609 (.in({n12863_2, n12862_0, n12841_1, n12840_0, n12811_0, n12810_0}), .out(n1528), .config_in(config_chain[1829:1827]), .config_rst(config_rst)); 
mux6 mux_610 (.in({n9753_2, n9752_0, n9729_0, n9728_0, n9691_0, n9690_0}), .out(n1529), .config_in(config_chain[1832:1830]), .config_rst(config_rst)); 
mux6 mux_611 (.in({n12611_2, n12610_0, n12581_0, n12580_0, n12549_0, n12548_0}), .out(n1530), .config_in(config_chain[1835:1833]), .config_rst(config_rst)); 
mux6 mux_612 (.in({n10005_2, n10004_0, n9983_0, n9982_0, n9945_0, n9944_0}), .out(n1531), .config_in(config_chain[1838:1836]), .config_rst(config_rst)); 
mux6 mux_613 (.in({n12867_2, n12866_0, n12843_0, n12842_0, n12805_0, n12804_0}), .out(n1532), .config_in(config_chain[1841:1839]), .config_rst(config_rst)); 
mux6 mux_614 (.in({n9773_1, n9772_0, n9765_1, n9764_0, n9755_2, n9754_0}), .out(n1533), .config_in(config_chain[1844:1842]), .config_rst(config_rst)); 
mux6 mux_615 (.in({n12613_2, n12612_0, n12583_1, n12582_0, n12553_0, n12552_0}), .out(n1534), .config_in(config_chain[1847:1845]), .config_rst(config_rst)); 
mux6 mux_616 (.in({n10283_1, n10282_0, n10201_0, n10200_0, n10179_0, n10178_0}), .out(n1581), .config_in(config_chain[1850:1848]), .config_rst(config_rst)); 
mux6 mux_617 (.in({n12887_1, n12886_0, n12805_0, n12804_0, n12783_0, n12782_0}), .out(n1582), .config_in(config_chain[1853:1851]), .config_rst(config_rst)); 
mux6 mux_618 (.in({n10013_1, n10012_0, n9979_0, n9978_0, n9947_0/**/, n9946_0}), .out(n1583), .config_in(config_chain[1856:1854]), .config_rst(config_rst)); 
mux6 mux_619 (.in({n12625_1, n12624_0, n12617_1, n12616_0, n12583_0, n12582_0}), .out(n1584), .config_in(config_chain[1859:1857]), .config_rst(config_rst)); 
mux6 mux_620 (.in({n10233_0, n10232_0/**/, n10211_0, n10210_0, n10181_0, n10180_0}), .out(n1585), .config_in(config_chain[1862:1860]), .config_rst(config_rst)); 
mux6 mux_621 (.in({n12847_0, n12846_0/**/, n12815_0, n12814_0, n12785_0, n12784_0}), .out(n1586), .config_in(config_chain[1865:1863]), .config_rst(config_rst)); 
mux6 mux_622 (.in({n10029_1, n10028_0, n9959_0, n9958_0, n9927_0, n9926_0}), .out(n1587), .config_in(config_chain[1868:1866]), .config_rst(config_rst)); 
mux6 mux_623 (.in({n12633_1, n12632_0, n12563_0, n12562_0, n12525_0, n12524_0}), .out(n1588), .config_in(config_chain[1871:1869]), .config_rst(config_rst)); 
mux6 mux_624 (.in({n10269_1, n10268_0, n10245_0, n10244_0, n10213_0, n10212_0}), .out(n1589), .config_in(config_chain[1874:1872]), .config_rst(config_rst)); 
mux6 mux_625 (.in({n12873_1, n12872_0, n12849_0, n12848_0, n12817_0, n12816_0}), .out(n1590), .config_in(config_chain[1877:1875]), .config_rst(config_rst)); 
mux6 mux_626 (.in({n9991_0, n9990_0, n9953_0, n9952_0, n9921_0, n9920_0}), .out(n1591), .config_in(config_chain[1880:1878]), .config_rst(config_rst)); 
mux6 mux_627 (.in({n12595_0, n12594_0, n12557_0, n12556_0, n12527_0, n12526_0}), .out(n1592), .config_in(config_chain[1883:1881]), .config_rst(config_rst)); 
mux6 mux_628 (.in({n10285_1, n10284_0, n10277_1, n10276_0, n10177_0, n10176_0}), .out(n1593), .config_in(config_chain[1886:1884]), .config_rst(config_rst)); 
mux6 mux_629 (.in({n12889_1, n12888_0, n12813_0, n12812_0, n12781_0, n12780_0}), .out(n1594), .config_in(config_chain[1889:1887]), .config_rst(config_rst)); 
mux6 mux_630 (.in({n10015_1, n10014_0, n9985_0, n9984_0, n9955_0, n9954_0}), .out(n1595), .config_in(config_chain[1892:1890]), .config_rst(config_rst)); 
mux6 mux_631 (.in({n12619_1, n12618_0, n12591_0, n12590_0/**/, n12559_0, n12558_0}), .out(n1596), .config_in(config_chain[1895:1893]), .config_rst(config_rst)); 
mux6 mux_632 (.in({n10241_0, n10240_0, n10219_0/**/, n10218_0, n10187_0, n10186_0}), .out(n1597), .config_in(config_chain[1898:1896]), .config_rst(config_rst)); 
mux6 mux_633 (.in({n12845_0, n12844_0, n12823_0, n12822_0/**/, n12793_0, n12792_0}), .out(n1598), .config_in(config_chain[1901:1899]), .config_rst(config_rst)); 
mux6 mux_634 (.in({n10023_1, n10022_0, n9987_0, n9986_0/**/, n9935_0, n9934_0}), .out(n1599), .config_in(config_chain[1904:1902]), .config_rst(config_rst)); 
mux6 mux_635 (.in({n12635_1/**/, n12634_0, n12627_1, n12626_0, n12539_0, n12538_0}), .out(n1600), .config_in(config_chain[1907:1905]), .config_rst(config_rst)); 
mux6 mux_636 (.in({n10251_0, n10250_0, n10221_0/**/, n10220_0, n10189_0, n10188_0}), .out(n1601), .config_in(config_chain[1910:1908]), .config_rst(config_rst)); 
mux6 mux_637 (.in({n12875_1, n12874_0, n12855_0, n12854_0/**/, n12825_0, n12824_0}), .out(n1602), .config_in(config_chain[1913:1911]), .config_rst(config_rst)); 
mux6 mux_638 (.in({n9999_0/**/, n9998_0, n9967_0, n9966_0, n9929_0, n9928_0}), .out(n1603), .config_in(config_chain[1916:1914]), .config_rst(config_rst)); 
mux6 mux_639 (.in({n12603_0, n12602_0, n12565_0, n12564_0, n12533_0, n12532_0}), .out(n1604), .config_in(config_chain[1919:1917]), .config_rst(config_rst)); 
mux6 mux_640 (.in({n10279_1, n10278_0, n10253_0, n10252_0, n10185_0, n10184_0}), .out(n1605), .config_in(config_chain[1922:1920]), .config_rst(config_rst)); 
mux6 mux_641 (.in({n12891_1, n12890_0, n12883_1, n12882_0, n12789_0, n12788_0}), .out(n1606), .config_in(config_chain[1925:1923]), .config_rst(config_rst)); 
mux6 mux_642 (.in({n9993_0, n9992_0, n9963_0, n9962_0, n9931_0/**/, n9930_0}), .out(n1607), .config_in(config_chain[1928:1926]), .config_rst(config_rst)); 
mux6 mux_643 (.in({n12597_0, n12596_0, n12567_0, n12566_0, n12535_0, n12534_0}), .out(n1608), .config_in(config_chain[1931:1929]), .config_rst(config_rst)); 
mux6 mux_644 (.in({n10287_1, n10286_0, n10217_0, n10216_0/**/, n10195_0, n10194_0}), .out(n1609), .config_in(config_chain[1934:1932]), .config_rst(config_rst)); 
mux6 mux_645 (.in({n12853_0, n12852_0, n12821_0, n12820_0, n12799_0, n12798_0}), .out(n1610), .config_in(config_chain[1937:1935]), .config_rst(config_rst)); 
mux6 mux_646 (.in({n10025_1, n10024_0, n10017_1, n10016_0, n9995_0, n9994_0/**/}), .out(n1611), .config_in(config_chain[1940:1938]), .config_rst(config_rst)); 
mux6 mux_647 (.in({n12629_1, n12628_0, n12599_0, n12598_0, n12547_0/**/, n12546_0}), .out(n1612), .config_in(config_chain[1943:1941]), .config_rst(config_rst)); 
mux6 mux_648 (.in({n10263_2, n10262_0, n10227_0, n10226_0, n10197_0/**/, n10196_0}), .out(n1613), .config_in(config_chain[1946:1944]), .config_rst(config_rst)); 
mux6 mux_649 (.in({n12867_2, n12866_0, n12833_0, n12832_0/**/, n12801_0, n12800_0}), .out(n1614), .config_in(config_chain[1949:1947]), .config_rst(config_rst)); 
mux6 mux_650 (.in({n10009_2, n10008_0, n9975_0/**/, n9974_0, n9937_0, n9936_0}), .out(n1615), .config_in(config_chain[1952:1950]), .config_rst(config_rst)); 
mux6 mux_651 (.in({n12613_2, n12612_0, n12579_0, n12578_0, n12541_0, n12540_0}), .out(n1616), .config_in(config_chain[1955:1953]), .config_rst(config_rst)); 
mux6 mux_652 (.in({n10273_1, n10272_0, n10265_2, n10264_0, n10229_0, n10228_0}), .out(n1617), .config_in(config_chain[1958:1956]), .config_rst(config_rst)); 
mux6 mux_653 (.in({n12885_1, n12884_0, n12877_1, n12876_0/**/, n12869_2, n12868_0}), .out(n1618), .config_in(config_chain[1961:1959]), .config_rst(config_rst)); 
mux6 mux_654 (.in({n10011_2, n10010_0, n9969_0, n9968_0, n9939_0, n9938_0/**/}), .out(n1619), .config_in(config_chain[1964:1962]), .config_rst(config_rst)); 
mux6 mux_655 (.in({n12605_1/**/, n12604_0, n12573_0, n12572_0, n12543_0, n12542_0}), .out(n1620), .config_in(config_chain[1967:1965]), .config_rst(config_rst)); 
mux6 mux_656 (.in({n10267_2, n10266_0, n10225_0, n10224_0, n10193_0, n10192_0}), .out(n1621), .config_in(config_chain[1970:1968]), .config_rst(config_rst)); 
mux6 mux_657 (.in({n12871_2/**/, n12870_0, n12829_0, n12828_0, n12807_0, n12806_0}), .out(n1622), .config_in(config_chain[1973:1971]), .config_rst(config_rst)); 
mux6 mux_658 (.in({n10019_1, n10018_0, n10003_2, n10002_0, n9971_0, n9970_0/**/}), .out(n1623), .config_in(config_chain[1976:1974]), .config_rst(config_rst)); 
mux6 mux_659 (.in({n12631_1, n12630_0, n12623_1, n12622_0, n12607_2, n12606_0}), .out(n1624), .config_in(config_chain[1979:1977]), .config_rst(config_rst)); 
mux6 mux_660 (.in({n10257_1, n10256_0, n10235_0/**/, n10234_0, n10203_0, n10202_0}), .out(n1625), .config_in(config_chain[1982:1980]), .config_rst(config_rst)); 
mux6 mux_661 (.in({n12861_1, n12860_0, n12839_0, n12838_0, n12809_0, n12808_0}), .out(n1626), .config_in(config_chain[1985:1983]), .config_rst(config_rst)); 
mux6 mux_662 (.in({n10027_1/**/, n10026_0, n10005_2, n10004_0, n9951_0, n9950_0}), .out(n1627), .config_in(config_chain[1988:1986]), .config_rst(config_rst)); 
mux6 mux_663 (.in({n12609_2, n12608_0, n12587_0/**/, n12586_0, n12555_0, n12554_0}), .out(n1628), .config_in(config_chain[1991:1989]), .config_rst(config_rst)); 
mux6 mux_664 (.in({n10275_1, n10274_0, n10259_1, n10258_0, n10237_0, n10236_0}), .out(n1629), .config_in(config_chain[1994:1992]), .config_rst(config_rst)); 
mux6 mux_665 (.in({n12879_1, n12878_0, n12865_2/**/, n12864_0, n12841_0, n12840_0}), .out(n1630), .config_in(config_chain[1997:1995]), .config_rst(config_rst)); 
mux6 mux_666 (.in({n10007_2, n10006_0, n9977_0/**/, n9976_0, n9945_0, n9944_0}), .out(n1631), .config_in(config_chain[2000:1998]), .config_rst(config_rst)); 
mux6 mux_667 (.in({n12611_2, n12610_0, n12581_0, n12580_0, n12551_0, n12550_0}), .out(n1632), .config_in(config_chain[2003:2001]), .config_rst(config_rst)); 
mux6 mux_668 (.in({n10527_1, n10526_0, n10495_0, n10494_0, n10465_0, n10464_0}), .out(n1679), .config_in(config_chain[2006:2004]), .config_rst(config_rst)); 
mux6 mux_669 (.in({n12893_1, n12892_0, n12879_0, n12878_0, n12841_0, n12840_0}), .out(n1680), .config_in(config_chain[2009:2007]), .config_rst(config_rst)); 
mux6 mux_670 (.in({n10233_0, n10232_0, n10201_0, n10200_0, n10179_0, n10178_0}), .out(n1681), .config_in(config_chain[2012:2010]), .config_rst(config_rst)); 
mux6 mux_671 (.in({n12581_0, n12580_0, n12559_0, n12558_0, n12527_0, n12526_0}), .out(n1682), .config_in(config_chain[2015:2013]), .config_rst(config_rst)); 
mux6 mux_672 (.in({n10535_1, n10534_0, n10497_0/**/, n10496_0, n10437_0, n10436_0}), .out(n1683), .config_in(config_chain[2018:2016]), .config_rst(config_rst)); 
mux6 mux_673 (.in({n12909_1, n12908_0, n12901_1, n12900_0, n12783_0, n12782_0}), .out(n1684), .config_in(config_chain[2021:2019]), .config_rst(config_rst)); 
mux6 mux_674 (.in({n10243_0, n10242_0, n10213_0, n10212_0, n10181_0, n10180_0}), .out(n1685), .config_in(config_chain[2024:2022]), .config_rst(config_rst)); 
mux6 mux_675 (.in({n12637_1, n12636_0, n12625_0, n12624_0, n12591_0, n12590_0}), .out(n1686), .config_in(config_chain[2027:2025]), .config_rst(config_rst)); 
mux6 mux_676 (.in({n10501_0/**/, n10500_0, n10469_0, n10468_0, n10439_0, n10438_0}), .out(n1687), .config_in(config_chain[2030:2028]), .config_rst(config_rst)); 
mux6 mux_677 (.in({n12847_0, n12846_0, n12815_0, n12814_0, n12785_0, n12784_0}), .out(n1688), .config_in(config_chain[2033:2031]), .config_rst(config_rst)); 
mux6 mux_678 (.in({n10277_1, n10276_0, n10269_1, n10268_0, n10245_0, n10244_0}), .out(n1689), .config_in(config_chain[2036:2034]), .config_rst(config_rst)); 
mux6 mux_679 (.in({n12645_1, n12644_0, n12633_0, n12632_0, n12525_0, n12524_0}), .out(n1690), .config_in(config_chain[2039:2037]), .config_rst(config_rst)); 
mux6 mux_680 (.in({n10503_0, n10502_0, n10471_0/**/, n10470_0, n10441_0, n10440_0}), .out(n1691), .config_in(config_chain[2042:2040]), .config_rst(config_rst)); 
mux6 mux_681 (.in({n12881_0, n12880_0, n12873_0/**/, n12872_0, n12849_0, n12848_0}), .out(n1692), .config_in(config_chain[2045:2043]), .config_rst(config_rst)); 
mux6 mux_682 (.in({n10285_1, n10284_0, n10209_0, n10208_0, n10187_0/**/, n10186_0}), .out(n1693), .config_in(config_chain[2048:2046]), .config_rst(config_rst)); 
mux6 mux_683 (.in({n12589_0, n12588_0, n12557_0, n12556_0, n12535_0/**/, n12534_0}), .out(n1694), .config_in(config_chain[2051:2049]), .config_rst(config_rst)); 
mux6 mux_684 (.in({n10537_1, n10536_0, n10529_1, n10528_0, n10505_0, n10504_0/**/}), .out(n1695), .config_in(config_chain[2054:2052]), .config_rst(config_rst)); 
mux6 mux_685 (.in({n12903_1, n12902_0, n12889_0, n12888_0, n12791_0, n12790_0}), .out(n1696), .config_in(config_chain[2057:2055]), .config_rst(config_rst)); 
mux6 mux_686 (.in({n10241_0/**/, n10240_0, n10219_0, n10218_0, n10189_0, n10188_0}), .out(n1697), .config_in(config_chain[2060:2058]), .config_rst(config_rst)); 
mux6 mux_687 (.in({n12619_0, n12618_0, n12599_0, n12598_0/**/, n12567_0, n12566_0}), .out(n1698), .config_in(config_chain[2063:2061]), .config_rst(config_rst)); 
mux6 mux_688 (.in({n10545_1, n10544_0, n10477_0, n10476_0, n10445_0/**/, n10444_0}), .out(n1699), .config_in(config_chain[2066:2064]), .config_rst(config_rst)); 
mux6 mux_689 (.in({n12911_1, n12910_0, n12823_0, n12822_0, n12793_0, n12792_0}), .out(n1700), .config_in(config_chain[2069:2067]), .config_rst(config_rst)); 
mux6 mux_690 (.in({n10271_1, n10270_0, n10253_0, n10252_0/**/, n10221_0, n10220_0}), .out(n1701), .config_in(config_chain[2072:2070]), .config_rst(config_rst)); 
mux6 mux_691 (.in({n12647_1, n12646_0, n12639_1, n12638_0, n12635_0, n12634_0}), .out(n1702), .config_in(config_chain[2075:2073]), .config_rst(config_rst)); 
mux6 mux_692 (.in({n10509_0, n10508_0, n10479_0, n10478_0, n10449_0/**/, n10448_0}), .out(n1703), .config_in(config_chain[2078:2076]), .config_rst(config_rst)); 
mux6 mux_693 (.in({n12875_0, n12874_0, n12857_0, n12856_0, n12825_0, n12824_0}), .out(n1704), .config_in(config_chain[2081:2079]), .config_rst(config_rst)); 
mux6 mux_694 (.in({n10287_1, n10286_0, n10217_0, n10216_0, n10185_0/**/, n10184_0}), .out(n1705), .config_in(config_chain[2084:2082]), .config_rst(config_rst)); 
mux6 mux_695 (.in({n12655_1, n12654_0, n12565_0, n12564_0, n12533_0, n12532_0/**/}), .out(n1706), .config_in(config_chain[2087:2085]), .config_rst(config_rst)); 
mux6 mux_696 (.in({n10531_1, n10530_0, n10511_0, n10510_0, n10481_0, n10480_0}), .out(n1707), .config_in(config_chain[2090:2088]), .config_rst(config_rst)); 
mux6 mux_697 (.in({n12897_1, n12896_0, n12891_0/**/, n12890_0, n12883_0, n12882_0}), .out(n1708), .config_in(config_chain[2093:2091]), .config_rst(config_rst)); 
mux6 mux_698 (.in({n10249_0, n10248_0, n10227_0, n10226_0/**/, n10195_0, n10194_0}), .out(n1709), .config_in(config_chain[2096:2094]), .config_rst(config_rst)); 
mux6 mux_699 (.in({n12621_0, n12620_0, n12597_0, n12596_0, n12575_0/**/, n12574_0}), .out(n1710), .config_in(config_chain[2099:2097]), .config_rst(config_rst)); 
mux6 mux_700 (.in({n10539_1, n10538_0, n10519_1, n10518_0, n10453_0, n10452_0}), .out(n1711), .config_in(config_chain[2102:2100]), .config_rst(config_rst)); 
mux6 mux_701 (.in({n12865_1, n12864_0, n12831_0, n12830_0, n12799_0/**/, n12798_0}), .out(n1712), .config_in(config_chain[2105:2103]), .config_rst(config_rst)); 
mux6 mux_702 (.in({n10273_1, n10272_0/**/, n10263_2, n10262_0, n10229_0, n10228_0}), .out(n1713), .config_in(config_chain[2108:2106]), .config_rst(config_rst)); 
mux6 mux_703 (.in({n12641_1/**/, n12640_0, n12629_0, n12628_0, n12611_2, n12610_0}), .out(n1714), .config_in(config_chain[2111:2109]), .config_rst(config_rst)); 
mux6 mux_704 (.in({n10521_2, n10520_0, n10485_0, n10484_0, n10455_0, n10454_0/**/}), .out(n1715), .config_in(config_chain[2114:2112]), .config_rst(config_rst)); 
mux6 mux_705 (.in({n12867_2, n12866_0, n12833_0/**/, n12832_0, n12801_0, n12800_0}), .out(n1716), .config_in(config_chain[2117:2115]), .config_rst(config_rst)); 
mux6 mux_706 (.in({n10281_1, n10280_0, n10265_2, n10264_0, n10193_0, n10192_0}), .out(n1717), .config_in(config_chain[2120:2118]), .config_rst(config_rst)); 
mux6 mux_707 (.in({n12649_1, n12648_0, n12615_2, n12614_0, n12541_0/**/, n12540_0}), .out(n1718), .config_in(config_chain[2123:2121]), .config_rst(config_rst)); 
mux6 mux_708 (.in({n10523_2, n10522_0, n10489_0, n10488_0, n10457_0/**/, n10456_0}), .out(n1719), .config_in(config_chain[2126:2124]), .config_rst(config_rst)); 
mux6 mux_709 (.in({n12899_1/**/, n12898_0, n12885_0, n12884_0, n12869_2, n12868_0}), .out(n1720), .config_in(config_chain[2129:2127]), .config_rst(config_rst)); 
mux6 mux_710 (.in({n10257_1, n10256_0, n10225_0/**/, n10224_0, n10203_0, n10202_0}), .out(n1721), .config_in(config_chain[2132:2130]), .config_rst(config_rst)); 
mux6 mux_711 (.in({n12605_1, n12604_0, n12583_0, n12582_0, n12551_0/**/, n12550_0}), .out(n1722), .config_in(config_chain[2135:2133]), .config_rst(config_rst)); 
mux6 mux_712 (.in({n10541_1, n10540_0, n10533_1, n10532_0, n10525_2, n10524_0}), .out(n1723), .config_in(config_chain[2138:2136]), .config_rst(config_rst)); 
mux6 mux_713 (.in({n12907_1, n12906_0, n12871_2, n12870_0, n12807_0, n12806_0}), .out(n1724), .config_in(config_chain[2141:2139]), .config_rst(config_rst)); 
mux6 mux_714 (.in({n10259_1, n10258_0, n10235_0, n10234_0, n10205_0, n10204_0}), .out(n1725), .config_in(config_chain[2144:2142]), .config_rst(config_rst)); 
mux6 mux_715 (.in({n12631_0, n12630_0, n12623_0, n12622_0, n12607_1, n12606_0}), .out(n1726), .config_in(config_chain[2147:2145]), .config_rst(config_rst)); 
mux6 mux_716 (.in({n10515_1, n10514_0, n10493_0/**/, n10492_0, n10463_0, n10462_0}), .out(n1727), .config_in(config_chain[2150:2148]), .config_rst(config_rst)); 
mux6 mux_717 (.in({n12863_1, n12862_0, n12839_0/**/, n12838_0, n12809_0, n12808_0}), .out(n1728), .config_in(config_chain[2153:2151]), .config_rst(config_rst)); 
mux6 mux_718 (.in({n10283_1, n10282_0/**/, n10275_1, n10274_0, n10261_2, n10260_0}), .out(n1729), .config_in(config_chain[2156:2154]), .config_rst(config_rst)); 
mux6 mux_719 (.in({n12651_1/**/, n12650_0, n12609_2, n12608_0, n12549_0, n12548_0}), .out(n1730), .config_in(config_chain[2159:2157]), .config_rst(config_rst)); 
mux6 mux_720 (.in({n10801_1, n10800_0, n10723_0/**/, n10722_0, n10701_0, n10700_0}), .out(n1777), .config_in(config_chain[2162:2160]), .config_rst(config_rst)); 
mux6 mux_721 (.in({n12927_1, n12926_0, n12873_0, n12872_0, n12809_0, n12808_1}), .out(n1778), .config_in(config_chain[2165:2163]), .config_rst(config_rst)); 
mux6 mux_722 (.in({n10527_1, n10526_0, n10497_0, n10496_0, n10465_0, n10464_0}), .out(n1779), .config_in(config_chain[2168:2166]), .config_rst(config_rst)); 
mux6 mux_723 (.in({n12665_1, n12664_0, n12657_1, n12656_0, n12651_0, n12650_0}), .out(n1780), .config_in(config_chain[2171:2169]), .config_rst(config_rst)); 
mux6 mux_724 (.in({n10755_0, n10754_0, n10733_0, n10732_0, n10695_0, n10694_0}), .out(n1781), .config_in(config_chain[2174:2172]), .config_rst(config_rst)); 
mux6 mux_725 (.in({n12893_0, n12892_0, n12889_0, n12888_0, n12881_0, n12880_0}), .out(n1782), .config_in(config_chain[2177:2175]), .config_rst(config_rst)); 
mux6 mux_726 (.in({n10543_1, n10542_0, n10469_0, n10468_0, n10437_0, n10436_0}), .out(n1783), .config_in(config_chain[2180:2178]), .config_rst(config_rst)); 
mux6 mux_727 (.in({n12673_1, n12672_0, n12617_0, n12616_0, n12559_0, n12558_1}), .out(n1784), .config_in(config_chain[2183:2181]), .config_rst(config_rst)); 
mux6 mux_728 (.in({n10787_1, n10786_0, n10759_0, n10758_0, n10727_0, n10726_0}), .out(n1785), .config_in(config_chain[2186:2184]), .config_rst(config_rst)); 
mux6 mux_729 (.in({n12913_1, n12912_0, n12909_0, n12908_0, n12901_0, n12900_0}), .out(n1786), .config_in(config_chain[2189:2187]), .config_rst(config_rst)); 
mux6 mux_730 (.in({n10501_0, n10500_0, n10471_0, n10470_0, n10439_0, n10438_0}), .out(n1787), .config_in(config_chain[2192:2190]), .config_rst(config_rst)); 
mux6 mux_731 (.in({n12637_0, n12636_0, n12625_0, n12624_0, n12591_0, n12590_1}), .out(n1788), .config_in(config_chain[2195:2193]), .config_rst(config_rst)); 
mux6 mux_732 (.in({n10803_1, n10802_0, n10795_1, n10794_0, n10699_0, n10698_0}), .out(n1789), .config_in(config_chain[2198:2196]), .config_rst(config_rst)); 
mux6 mux_733 (.in({n12929_1, n12928_0, n12817_0, n12816_1, n12785_0, n12784_1}), .out(n1790), .config_in(config_chain[2201:2199]), .config_rst(config_rst)); 
mux6 mux_734 (.in({n10529_1, n10528_0/**/, n10503_0, n10502_0, n10473_0, n10472_0}), .out(n1791), .config_in(config_chain[2204:2202]), .config_rst(config_rst)); 
mux6 mux_735 (.in({n12659_1, n12658_0, n12653_0, n12652_0, n12645_0, n12644_0}), .out(n1792), .config_in(config_chain[2207:2205]), .config_rst(config_rst)); 
mux6 mux_736 (.in({n10763_0, n10762_0, n10741_0/**/, n10740_0, n10709_0, n10708_0}), .out(n1793), .config_in(config_chain[2210:2208]), .config_rst(config_rst)); 
mux6 mux_737 (.in({n12895_0, n12894_0, n12883_0, n12882_0, n12849_0, n12848_1}), .out(n1794), .config_in(config_chain[2213:2211]), .config_rst(config_rst)); 
mux6 mux_738 (.in({n10537_1, n10536_0, n10505_0, n10504_0, n10445_0/**/, n10444_0}), .out(n1795), .config_in(config_chain[2216:2214]), .config_rst(config_rst)); 
mux6 mux_739 (.in({n12675_1, n12674_0, n12667_1, n12666_0/**/, n12535_0, n12534_1}), .out(n1796), .config_in(config_chain[2219:2217]), .config_rst(config_rst)); 
mux6 mux_740 (.in({n10773_0, n10772_0, n10735_0/**/, n10734_0, n10703_0, n10702_0}), .out(n1797), .config_in(config_chain[2222:2220]), .config_rst(config_rst)); 
mux6 mux_741 (.in({n12915_1, n12914_0, n12903_0, n12902_0, n12891_0, n12890_0}), .out(n1798), .config_in(config_chain[2225:2223]), .config_rst(config_rst)); 
mux6 mux_742 (.in({n10509_0/**/, n10508_0, n10477_0, n10476_0, n10447_0, n10446_0}), .out(n1799), .config_in(config_chain[2228:2226]), .config_rst(config_rst)); 
mux6 mux_743 (.in({n12627_0, n12626_0, n12619_0, n12618_0, n12599_0, n12598_1/**/}), .out(n1800), .config_in(config_chain[2231:2229]), .config_rst(config_rst)); 
mux6 mux_744 (.in({n10797_1, n10796_0/**/, n10767_0, n10766_0, n10707_0, n10706_0}), .out(n1801), .config_in(config_chain[2234:2232]), .config_rst(config_rst)); 
mux6 mux_745 (.in({n12931_1/**/, n12930_0, n12923_1, n12922_0, n12793_0, n12792_1}), .out(n1802), .config_in(config_chain[2237:2235]), .config_rst(config_rst)); 
mux6 mux_746 (.in({n10511_0/**/, n10510_0, n10481_0, n10480_0, n10449_0, n10448_0}), .out(n1803), .config_in(config_chain[2240:2238]), .config_rst(config_rst)); 
mux6 mux_747 (.in({n12647_0/**/, n12646_0, n12639_0, n12638_0, n12635_0, n12634_0}), .out(n1804), .config_in(config_chain[2243:2241]), .config_rst(config_rst)); 
mux6 mux_748 (.in({n10805_1, n10804_0, n10739_0, n10738_0, n10717_0, n10716_0}), .out(n1805), .config_in(config_chain[2246:2244]), .config_rst(config_rst)); 
mux6 mux_749 (.in({n12877_0, n12876_0, n12857_0, n12856_1/**/, n12825_0, n12824_1}), .out(n1806), .config_in(config_chain[2249:2247]), .config_rst(config_rst)); 
mux6 mux_750 (.in({n10539_1, n10538_0, n10531_1, n10530_0, n10513_0, n10512_0}), .out(n1807), .config_in(config_chain[2252:2250]), .config_rst(config_rst)); 
mux6 mux_751 (.in({n12669_1, n12668_0, n12655_0, n12654_0/**/, n12543_0, n12542_1}), .out(n1808), .config_in(config_chain[2255:2253]), .config_rst(config_rst)); 
mux6 mux_752 (.in({n10777_1, n10776_0, n10749_0/**/, n10748_0, n10711_0, n10710_0}), .out(n1809), .config_in(config_chain[2258:2256]), .config_rst(config_rst)); 
mux6 mux_753 (.in({n12905_0, n12904_0/**/, n12897_0, n12896_0, n12863_1, n12862_1}), .out(n1810), .config_in(config_chain[2261:2259]), .config_rst(config_rst)); 
mux6 mux_754 (.in({n10519_1, n10518_0, n10485_0, n10484_0/**/, n10455_0, n10454_0}), .out(n1811), .config_in(config_chain[2264:2262]), .config_rst(config_rst)); 
mux6 mux_755 (.in({n12621_0/**/, n12620_0, n12609_1, n12608_1, n12575_0, n12574_1}), .out(n1812), .config_in(config_chain[2267:2265]), .config_rst(config_rst)); 
mux6 mux_756 (.in({n10791_1, n10790_0, n10779_1, n10778_0, n10743_0, n10742_0/**/}), .out(n1813), .config_in(config_chain[2270:2268]), .config_rst(config_rst)); 
mux6 mux_757 (.in({n12925_1, n12924_0, n12917_1, n12916_0, n12865_1/**/, n12864_1}), .out(n1814), .config_in(config_chain[2273:2271]), .config_rst(config_rst)); 
mux6 mux_758 (.in({n10521_2, n10520_0, n10487_0, n10486_0, n10457_0, n10456_0}), .out(n1815), .config_in(config_chain[2276:2274]), .config_rst(config_rst)); 
mux6 mux_759 (.in({n12641_0, n12640_0, n12629_0, n12628_0, n12613_1, n12612_1}), .out(n1816), .config_in(config_chain[2279:2277]), .config_rst(config_rst)); 
mux6 mux_760 (.in({n10781_1, n10780_0, n10747_0, n10746_0/**/, n10715_0, n10714_0}), .out(n1817), .config_in(config_chain[2282:2280]), .config_rst(config_rst)); 
mux6 mux_761 (.in({n12879_0, n12878_0, n12867_1, n12866_1, n12833_0/**/, n12832_1}), .out(n1818), .config_in(config_chain[2285:2283]), .config_rst(config_rst)); 
mux6 mux_762 (.in({n10533_1, n10532_0, n10525_2, n10524_0, n10489_0, n10488_0}), .out(n1819), .config_in(config_chain[2288:2286]), .config_rst(config_rst)); 
mux6 mux_763 (.in({n12671_1, n12670_0, n12663_1, n12662_0, n12615_1, n12614_1}), .out(n1820), .config_in(config_chain[2291:2289]), .config_rst(config_rst)); 
mux6 mux_764 (.in({n10783_2, n10782_0, n10757_0/**/, n10756_0, n10725_0, n10724_0}), .out(n1821), .config_in(config_chain[2294:2292]), .config_rst(config_rst)); 
mux6 mux_765 (.in({n12899_0, n12898_0, n12887_0, n12886_0, n12869_1, n12868_1}), .out(n1822), .config_in(config_chain[2297:2295]), .config_rst(config_rst)); 
mux6 mux_766 (.in({n10541_1, n10540_0, n10515_1, n10514_0, n10461_0, n10460_0}), .out(n1823), .config_in(config_chain[2300:2298]), .config_rst(config_rst)); 
mux6 mux_767 (.in({n12605_1, n12604_1, n12583_0, n12582_1, n12551_0, n12550_1}), .out(n1824), .config_in(config_chain[2303:2301]), .config_rst(config_rst)); 
mux6 mux_768 (.in({n10793_1, n10792_0, n10785_2, n10784_0, n10751_0/**/, n10750_0}), .out(n1825), .config_in(config_chain[2306:2304]), .config_rst(config_rst)); 
mux6 mux_769 (.in({n12919_1, n12918_0, n12907_0, n12906_0, n12861_0, n12860_1}), .out(n1826), .config_in(config_chain[2309:2307]), .config_rst(config_rst)); 
mux6 mux_770 (.in({n10517_1, n10516_0, n10495_0, n10494_0, n10463_0/**/, n10462_0}), .out(n1827), .config_in(config_chain[2312:2310]), .config_rst(config_rst)); 
mux6 mux_771 (.in({n12643_0, n12642_0, n12631_0, n12630_0, n12607_1, n12606_1}), .out(n1828), .config_in(config_chain[2315:2313]), .config_rst(config_rst)); 
mux6 mux_772 (.in({n11049_1, n11048_0, n11013_0, n11012_0, n10983_0, n10982_0}), .out(n1875), .config_in(config_chain[2318:2316]), .config_rst(config_rst)); 
mux6 mux_773 (.in({n12933_1, n12932_0, n12919_0, n12918_0, n12907_0, n12906_0}), .out(n1876), .config_in(config_chain[2321:2319]), .config_rst(config_rst)); 
mux6 mux_774 (.in({n10755_0, n10754_0, n10723_0, n10722_0, n10701_0, n10700_0}), .out(n1877), .config_in(config_chain[2324:2322]), .config_rst(config_rst)); 
mux6 mux_775 (.in({n12645_0, n12644_0, n12637_0, n12636_0/**/, n12631_0, n12630_1}), .out(n1878), .config_in(config_chain[2327:2325]), .config_rst(config_rst)); 
mux6 mux_776 (.in({n11057_1, n11056_0, n11015_0, n11014_0, n10963_0, n10962_0}), .out(n1879), .config_in(config_chain[2330:2328]), .config_rst(config_rst)); 
mux6 mux_777 (.in({n12949_1, n12948_0, n12941_1, n12940_0, n12873_0, n12872_1}), .out(n1880), .config_in(config_chain[2333:2331]), .config_rst(config_rst)); 
mux6 mux_778 (.in({n10765_0, n10764_0, n10727_0, n10726_0, n10695_0, n10694_0}), .out(n1881), .config_in(config_chain[2336:2334]), .config_rst(config_rst)); 
mux6 mux_779 (.in({n12677_1, n12676_0, n12665_0/**/, n12664_0, n12653_0, n12652_0}), .out(n1882), .config_in(config_chain[2339:2337]), .config_rst(config_rst)); 
mux6 mux_780 (.in({n11027_0, n11026_0, n10995_0/**/, n10994_0, n10957_0, n10956_0}), .out(n1883), .config_in(config_chain[2342:2340]), .config_rst(config_rst)); 
mux6 mux_781 (.in({n12893_0, n12892_0, n12889_0, n12888_1, n12881_0, n12880_1}), .out(n1884), .config_in(config_chain[2345:2343]), .config_rst(config_rst)); 
mux6 mux_782 (.in({n10795_1, n10794_0, n10787_1, n10786_0, n10759_0, n10758_0}), .out(n1885), .config_in(config_chain[2348:2346]), .config_rst(config_rst)); 
mux6 mux_783 (.in({n12685_1, n12684_0, n12673_0, n12672_0, n12617_0, n12616_1}), .out(n1886), .config_in(config_chain[2351:2349]), .config_rst(config_rst)); 
mux6 mux_784 (.in({n11021_0, n11020_0/**/, n10989_0, n10988_0, n10959_0, n10958_0}), .out(n1887), .config_in(config_chain[2354:2352]), .config_rst(config_rst)); 
mux6 mux_785 (.in({n12921_0, n12920_0, n12913_0, n12912_0, n12909_0, n12908_0}), .out(n1888), .config_in(config_chain[2357:2355]), .config_rst(config_rst)); 
mux6 mux_786 (.in({n10803_1, n10802_0, n10731_0/**/, n10730_0, n10709_0, n10708_0}), .out(n1889), .config_in(config_chain[2360:2358]), .config_rst(config_rst)); 
mux6 mux_787 (.in({n12639_0, n12638_0, n12633_0, n12632_1, n12625_0, n12624_1}), .out(n1890), .config_in(config_chain[2363:2361]), .config_rst(config_rst)); 
mux6 mux_788 (.in({n11059_1, n11058_0, n11051_1, n11050_0, n11023_0, n11022_0/**/}), .out(n1891), .config_in(config_chain[2366:2364]), .config_rst(config_rst)); 
mux6 mux_789 (.in({n12943_1, n12942_0, n12929_0, n12928_0/**/, n12875_0, n12874_1}), .out(n1892), .config_in(config_chain[2369:2367]), .config_rst(config_rst)); 
mux6 mux_790 (.in({n10763_0, n10762_0, n10741_0, n10740_0, n10703_0, n10702_0}), .out(n1893), .config_in(config_chain[2372:2370]), .config_rst(config_rst)); 
mux6 mux_791 (.in({n12659_0, n12658_0, n12655_0, n12654_0/**/, n12647_0, n12646_0}), .out(n1894), .config_in(config_chain[2375:2373]), .config_rst(config_rst)); 
mux6 mux_792 (.in({n11067_1, n11066_0, n11003_0, n11002_0, n10971_0/**/, n10970_0}), .out(n1895), .config_in(config_chain[2378:2376]), .config_rst(config_rst)); 
mux6 mux_793 (.in({n12951_1/**/, n12950_0, n12895_0, n12894_0, n12883_0, n12882_1}), .out(n1896), .config_in(config_chain[2381:2379]), .config_rst(config_rst)); 
mux6 mux_794 (.in({n10789_1, n10788_0, n10767_0, n10766_0, n10735_0, n10734_0}), .out(n1897), .config_in(config_chain[2384:2382]), .config_rst(config_rst)); 
mux6 mux_795 (.in({n12687_1, n12686_0, n12679_1, n12678_0, n12675_0, n12674_0}), .out(n1898), .config_in(config_chain[2387:2385]), .config_rst(config_rst)); 
mux6 mux_796 (.in({n11035_0, n11034_0, n10997_0, n10996_0, n10967_0, n10966_0}), .out(n1899), .config_in(config_chain[2390:2388]), .config_rst(config_rst)); 
mux6 mux_797 (.in({n12915_0, n12914_0, n12911_0/**/, n12910_0, n12903_0, n12902_0}), .out(n1900), .config_in(config_chain[2393:2391]), .config_rst(config_rst)); 
mux6 mux_798 (.in({n10805_1, n10804_0, n10739_0/**/, n10738_0, n10707_0, n10706_0}), .out(n1901), .config_in(config_chain[2396:2394]), .config_rst(config_rst)); 
mux6 mux_799 (.in({n12695_1, n12694_0, n12627_0, n12626_1, n12619_0/**/, n12618_1}), .out(n1902), .config_in(config_chain[2399:2397]), .config_rst(config_rst)); 
mux6 mux_800 (.in({n11053_1/**/, n11052_0, n11029_0, n11028_0, n10999_0, n10998_0}), .out(n1903), .config_in(config_chain[2402:2400]), .config_rst(config_rst)); 
mux6 mux_801 (.in({n12937_1, n12936_0, n12931_0, n12930_0, n12923_0, n12922_0}), .out(n1904), .config_in(config_chain[2405:2403]), .config_rst(config_rst)); 
mux6 mux_802 (.in({n10771_0, n10770_0, n10749_0, n10748_0, n10717_0, n10716_0}), .out(n1905), .config_in(config_chain[2408:2406]), .config_rst(config_rst)); 
mux6 mux_803 (.in({n12661_0/**/, n12660_0, n12649_0, n12648_0, n12635_0, n12634_1}), .out(n1906), .config_in(config_chain[2411:2409]), .config_rst(config_rst)); 
mux6 mux_804 (.in({n11061_1, n11060_0, n11037_0, n11036_0, n10979_0, n10978_0}), .out(n1907), .config_in(config_chain[2414:2412]), .config_rst(config_rst)); 
mux6 mux_805 (.in({n12885_0, n12884_1, n12877_0, n12876_1, n12861_0, n12860_1}), .out(n1908), .config_in(config_chain[2417:2415]), .config_rst(config_rst)); 
mux6 mux_806 (.in({n10791_1, n10790_0, n10777_1, n10776_0, n10743_0, n10742_0}), .out(n1909), .config_in(config_chain[2420:2418]), .config_rst(config_rst)); 
mux6 mux_807 (.in({n12681_1/**/, n12680_0, n12669_0, n12668_0, n12607_1, n12606_1}), .out(n1910), .config_in(config_chain[2423:2421]), .config_rst(config_rst)); 
mux6 mux_808 (.in({n11039_0, n11038_0, n11011_0, n11010_0, n10973_0, n10972_0/**/}), .out(n1911), .config_in(config_chain[2426:2424]), .config_rst(config_rst)); 
mux6 mux_809 (.in({n12905_0, n12904_0, n12897_0, n12896_0/**/, n12863_0, n12862_1}), .out(n1912), .config_in(config_chain[2429:2427]), .config_rst(config_rst)); 
mux6 mux_810 (.in({n10799_1, n10798_0, n10779_1, n10778_0, n10715_0, n10714_0/**/}), .out(n1913), .config_in(config_chain[2432:2430]), .config_rst(config_rst)); 
mux6 mux_811 (.in({n12689_1, n12688_0, n12621_0, n12620_1, n12611_1, n12610_1}), .out(n1914), .config_in(config_chain[2435:2433]), .config_rst(config_rst)); 
mux6 mux_812 (.in({n11041_1, n11040_0, n11007_0, n11006_0, n10975_0, n10974_0}), .out(n1915), .config_in(config_chain[2438:2436]), .config_rst(config_rst)); 
mux6 mux_813 (.in({n12939_1, n12938_0, n12925_0, n12924_0, n12865_1, n12864_1}), .out(n1916), .config_in(config_chain[2441:2439]), .config_rst(config_rst)); 
mux6 mux_814 (.in({n10783_2, n10782_0, n10747_0/**/, n10746_0, n10725_0, n10724_0}), .out(n1917), .config_in(config_chain[2444:2442]), .config_rst(config_rst)); 
mux6 mux_815 (.in({n12651_0, n12650_0/**/, n12643_0, n12642_0, n12613_1, n12612_1}), .out(n1918), .config_in(config_chain[2447:2445]), .config_rst(config_rst)); 
mux6 mux_816 (.in({n11063_1, n11062_0, n11055_1, n11054_0, n11043_1, n11042_0}), .out(n1919), .config_in(config_chain[2450:2448]), .config_rst(config_rst)); 
mux6 mux_817 (.in({n12947_1, n12946_0, n12879_0/**/, n12878_1, n12867_1, n12866_1}), .out(n1920), .config_in(config_chain[2453:2451]), .config_rst(config_rst)); 
mux6 mux_818 (.in({n10785_2, n10784_0, n10757_0/**/, n10756_0, n10719_0, n10718_0}), .out(n1921), .config_in(config_chain[2456:2454]), .config_rst(config_rst)); 
mux6 mux_819 (.in({n12671_0, n12670_0, n12663_0, n12662_0/**/, n12615_1, n12614_1}), .out(n1922), .config_in(config_chain[2459:2457]), .config_rst(config_rst)); 
mux6 mux_820 (.in({n11045_1, n11044_0, n11019_0/**/, n11018_0, n10981_0, n10980_0}), .out(n1923), .config_in(config_chain[2462:2460]), .config_rst(config_rst)); 
mux6 mux_821 (.in({n12899_0, n12898_0, n12887_0/**/, n12886_1, n12871_1, n12870_1}), .out(n1924), .config_in(config_chain[2465:2463]), .config_rst(config_rst)); 
mux6 mux_822 (.in({n10801_1, n10800_0, n10793_1, n10792_0/**/, n10775_0, n10774_0}), .out(n1925), .config_in(config_chain[2468:2466]), .config_rst(config_rst)); 
mux6 mux_823 (.in({n12691_1, n12690_0, n12623_0, n12622_1/**/, n12605_0, n12604_1}), .out(n1926), .config_in(config_chain[2471:2469]), .config_rst(config_rst)); 
mux6 mux_824 (.in({n11327_1, n11326_0, n11245_0, n11244_0, n11223_0, n11222_0}), .out(n1973), .config_in(config_chain[2474:2472]), .config_rst(config_rst)); 
mux6 mux_825 (.in({n12967_1, n12966_0, n12913_0, n12912_0, n12899_0, n12898_1}), .out(n1974), .config_in(config_chain[2477:2475]), .config_rst(config_rst)); 
mux6 mux_826 (.in({n11049_1, n11048_0, n11015_0, n11014_0, n10983_0, n10982_0}), .out(n1975), .config_in(config_chain[2480:2478]), .config_rst(config_rst)); 
mux6 mux_827 (.in({n12705_1, n12704_0, n12697_1, n12696_0, n12691_0, n12690_0}), .out(n1976), .config_in(config_chain[2483:2481]), .config_rst(config_rst)); 
mux6 mux_828 (.in({n11277_0, n11276_0, n11255_0, n11254_0, n11225_0, n11224_0}), .out(n1977), .config_in(config_chain[2486:2484]), .config_rst(config_rst)); 
mux6 mux_829 (.in({n12933_0, n12932_0, n12929_0, n12928_0, n12921_0, n12920_0}), .out(n1978), .config_in(config_chain[2489:2487]), .config_rst(config_rst)); 
mux6 mux_830 (.in({n11065_1, n11064_0, n10995_0, n10994_0, n10963_0, n10962_0}), .out(n1979), .config_in(config_chain[2492:2490]), .config_rst(config_rst)); 
mux6 mux_831 (.in({n12713_1, n12712_0, n12657_0, n12656_0, n12645_0, n12644_1}), .out(n1980), .config_in(config_chain[2495:2493]), .config_rst(config_rst)); 
mux6 mux_832 (.in({n11313_1, n11312_0, n11289_0, n11288_0, n11257_0, n11256_0}), .out(n1981), .config_in(config_chain[2498:2496]), .config_rst(config_rst)); 
mux6 mux_833 (.in({n12953_1, n12952_0, n12949_0, n12948_0, n12941_0/**/, n12940_0}), .out(n1982), .config_in(config_chain[2501:2499]), .config_rst(config_rst)); 
mux6 mux_834 (.in({n11027_0, n11026_0/**/, n10989_0, n10988_0, n10957_0, n10956_0}), .out(n1983), .config_in(config_chain[2504:2502]), .config_rst(config_rst)); 
mux6 mux_835 (.in({n12677_0, n12676_0, n12665_0, n12664_0, n12653_0, n12652_1}), .out(n1984), .config_in(config_chain[2507:2505]), .config_rst(config_rst)); 
mux6 mux_836 (.in({n11329_1, n11328_0, n11321_1, n11320_0, n11221_0, n11220_0}), .out(n1985), .config_in(config_chain[2510:2508]), .config_rst(config_rst)); 
mux6 mux_837 (.in({n12969_1, n12968_0, n12901_0, n12900_1, n12893_0, n12892_1}), .out(n1986), .config_in(config_chain[2513:2511]), .config_rst(config_rst)); 
mux6 mux_838 (.in({n11051_1, n11050_0, n11021_0, n11020_0, n10991_0/**/, n10990_0}), .out(n1987), .config_in(config_chain[2516:2514]), .config_rst(config_rst)); 
mux6 mux_839 (.in({n12699_1, n12698_0, n12693_0, n12692_0/**/, n12685_0, n12684_0}), .out(n1988), .config_in(config_chain[2519:2517]), .config_rst(config_rst)); 
mux6 mux_840 (.in({n11285_0, n11284_0, n11263_0, n11262_0, n11231_0/**/, n11230_0}), .out(n1989), .config_in(config_chain[2522:2520]), .config_rst(config_rst)); 
mux6 mux_841 (.in({n12935_0, n12934_0, n12923_0, n12922_0, n12909_0, n12908_1}), .out(n1990), .config_in(config_chain[2525:2523]), .config_rst(config_rst)); 
mux6 mux_842 (.in({n11059_1, n11058_0, n11023_0, n11022_0, n10971_0, n10970_0/**/}), .out(n1991), .config_in(config_chain[2528:2526]), .config_rst(config_rst)); 
mux6 mux_843 (.in({n12715_1, n12714_0, n12707_1, n12706_0/**/, n12639_0, n12638_1}), .out(n1992), .config_in(config_chain[2531:2529]), .config_rst(config_rst)); 
mux6 mux_844 (.in({n11295_0/**/, n11294_0, n11265_0, n11264_0, n11233_0, n11232_0}), .out(n1993), .config_in(config_chain[2534:2532]), .config_rst(config_rst)); 
mux6 mux_845 (.in({n12955_1, n12954_0, n12943_0, n12942_0, n12931_0/**/, n12930_0}), .out(n1994), .config_in(config_chain[2537:2535]), .config_rst(config_rst)); 
mux6 mux_846 (.in({n11035_0, n11034_0, n11003_0, n11002_0, n10965_0, n10964_0}), .out(n1995), .config_in(config_chain[2540:2538]), .config_rst(config_rst)); 
mux6 mux_847 (.in({n12667_0, n12666_0, n12659_0, n12658_0, n12655_0, n12654_1}), .out(n1996), .config_in(config_chain[2543:2541]), .config_rst(config_rst)); 
mux6 mux_848 (.in({n11323_1, n11322_0, n11297_0, n11296_0, n11229_0, n11228_0}), .out(n1997), .config_in(config_chain[2546:2544]), .config_rst(config_rst)); 
mux6 mux_849 (.in({n12971_1, n12970_0, n12963_1, n12962_0, n12895_0, n12894_1}), .out(n1998), .config_in(config_chain[2549:2547]), .config_rst(config_rst)); 
mux6 mux_850 (.in({n11029_0, n11028_0, n10999_0, n10998_0, n10967_0, n10966_0/**/}), .out(n1999), .config_in(config_chain[2552:2550]), .config_rst(config_rst)); 
mux6 mux_851 (.in({n12687_0, n12686_0, n12679_0, n12678_0/**/, n12675_0, n12674_0}), .out(n2000), .config_in(config_chain[2555:2553]), .config_rst(config_rst)); 
mux6 mux_852 (.in({n11331_1, n11330_0, n11261_0, n11260_0/**/, n11239_0, n11238_0}), .out(n2001), .config_in(config_chain[2558:2556]), .config_rst(config_rst)); 
mux6 mux_853 (.in({n12917_0, n12916_0, n12911_0, n12910_1/**/, n12903_0, n12902_1}), .out(n2002), .config_in(config_chain[2561:2559]), .config_rst(config_rst)); 
mux6 mux_854 (.in({n11061_1, n11060_0, n11053_1, n11052_0, n11031_0, n11030_0}), .out(n2003), .config_in(config_chain[2564:2562]), .config_rst(config_rst)); 
mux6 mux_855 (.in({n12709_1, n12708_0, n12695_0, n12694_0/**/, n12641_0, n12640_1}), .out(n2004), .config_in(config_chain[2567:2565]), .config_rst(config_rst)); 
mux6 mux_856 (.in({n11311_1, n11310_0, n11271_0, n11270_0, n11241_0, n11240_0}), .out(n2005), .config_in(config_chain[2570:2568]), .config_rst(config_rst)); 
mux6 mux_857 (.in({n12945_0, n12944_0, n12937_0/**/, n12936_0, n12871_1, n12870_1}), .out(n2006), .config_in(config_chain[2573:2571]), .config_rst(config_rst)); 
mux6 mux_858 (.in({n11037_0, n11036_0, n11011_0, n11010_0, n10973_0, n10972_0}), .out(n2007), .config_in(config_chain[2576:2574]), .config_rst(config_rst)); 
mux6 mux_859 (.in({n12661_0, n12660_0, n12649_0, n12648_1/**/, n12605_0, n12604_1}), .out(n2008), .config_in(config_chain[2579:2577]), .config_rst(config_rst)); 
mux6 mux_860 (.in({n11317_1, n11316_0, n11301_0, n11300_0, n11273_0/**/, n11272_0}), .out(n2009), .config_in(config_chain[2582:2580]), .config_rst(config_rst)); 
mux6 mux_861 (.in({n12965_1, n12964_0, n12957_1, n12956_0, n12861_0, n12860_1}), .out(n2010), .config_in(config_chain[2585:2583]), .config_rst(config_rst)); 
mux6 mux_862 (.in({n11039_0, n11038_0, n11005_0, n11004_0, n10975_0, n10974_0}), .out(n2011), .config_in(config_chain[2588:2586]), .config_rst(config_rst)); 
mux6 mux_863 (.in({n12681_0, n12680_0, n12669_0, n12668_0, n12609_1, n12608_1}), .out(n2012), .config_in(config_chain[2591:2589]), .config_rst(config_rst)); 
mux6 mux_864 (.in({n11303_0, n11302_0, n11269_0/**/, n11268_0, n11237_0, n11236_0}), .out(n2013), .config_in(config_chain[2594:2592]), .config_rst(config_rst)); 
mux6 mux_865 (.in({n12919_0, n12918_0, n12905_0, n12904_1, n12863_0, n12862_1}), .out(n2014), .config_in(config_chain[2597:2595]), .config_rst(config_rst)); 
mux6 mux_866 (.in({n11055_1, n11054_0, n11043_1, n11042_0, n11007_0, n11006_0}), .out(n2015), .config_in(config_chain[2600:2598]), .config_rst(config_rst)); 
mux6 mux_867 (.in({n12711_1, n12710_0, n12703_1/**/, n12702_0, n12611_1, n12610_1}), .out(n2016), .config_in(config_chain[2603:2601]), .config_rst(config_rst)); 
mux6 mux_868 (.in({n11305_0, n11304_0, n11279_0, n11278_0, n11247_0/**/, n11246_0}), .out(n2017), .config_in(config_chain[2606:2604]), .config_rst(config_rst)); 
mux6 mux_869 (.in({n12939_0, n12938_0, n12927_0, n12926_0, n12865_0/**/, n12864_1}), .out(n2018), .config_in(config_chain[2609:2607]), .config_rst(config_rst)); 
mux6 mux_870 (.in({n11063_1, n11062_0, n11045_1, n11044_0, n10987_0, n10986_0/**/}), .out(n2019), .config_in(config_chain[2612:2610]), .config_rst(config_rst)); 
mux6 mux_871 (.in({n12651_0, n12650_1, n12643_0, n12642_1, n12613_1, n12612_1}), .out(n2020), .config_in(config_chain[2615:2613]), .config_rst(config_rst)); 
mux6 mux_872 (.in({n11319_1, n11318_0, n11307_1, n11306_0, n11281_0, n11280_0}), .out(n2021), .config_in(config_chain[2618:2616]), .config_rst(config_rst)); 
mux6 mux_873 (.in({n12959_1, n12958_0, n12947_0, n12946_0, n12869_1, n12868_1}), .out(n2022), .config_in(config_chain[2621:2619]), .config_rst(config_rst)); 
mux6 mux_874 (.in({n11047_2, n11046_0, n11013_0/**/, n11012_0, n10981_0, n10980_0}), .out(n2023), .config_in(config_chain[2624:2622]), .config_rst(config_rst)); 
mux6 mux_875 (.in({n12683_0, n12682_0, n12671_0/**/, n12670_0, n12615_1, n12614_1}), .out(n2024), .config_in(config_chain[2627:2625]), .config_rst(config_rst)); 
mux6 mux_876 (.in({n11577_1, n11576_0, n11545_0, n11544_0, n11515_0, n11514_0}), .out(n2071), .config_in(config_chain[2630:2628]), .config_rst(config_rst)); 
mux6 mux_877 (.in({n12973_0, n12972_0, n12959_0, n12958_0, n12947_0, n12946_0}), .out(n2072), .config_in(config_chain[2633:2631]), .config_rst(config_rst)); 
mux6 mux_878 (.in({n11277_0, n11276_0, n11245_0, n11244_0, n11223_0, n11222_0}), .out(n2073), .config_in(config_chain[2636:2634]), .config_rst(config_rst)); 
mux6 mux_879 (.in({n12685_0, n12684_0, n12677_0, n12676_0, n12671_0, n12670_1}), .out(n2074), .config_in(config_chain[2639:2637]), .config_rst(config_rst)); 
mux6 mux_880 (.in({n11585_1, n11584_0, n11547_0, n11546_0, n11487_0, n11486_0}), .out(n2075), .config_in(config_chain[2642:2640]), .config_rst(config_rst)); 
mux6 mux_881 (.in({n12989_0, n12988_0, n12981_0/**/, n12980_0, n12913_0, n12912_1}), .out(n2076), .config_in(config_chain[2645:2643]), .config_rst(config_rst)); 
mux6 mux_882 (.in({n11287_0, n11286_0, n11257_0/**/, n11256_0, n11225_0, n11224_0}), .out(n2077), .config_in(config_chain[2648:2646]), .config_rst(config_rst)); 
mux6 mux_883 (.in({n12717_0, n12716_0, n12705_0, n12704_0, n12693_0, n12692_0}), .out(n2078), .config_in(config_chain[2651:2649]), .config_rst(config_rst)); 
mux6 mux_884 (.in({n11551_0, n11550_0, n11519_0, n11518_0, n11489_0, n11488_0}), .out(n2079), .config_in(config_chain[2654:2652]), .config_rst(config_rst)); 
mux6 mux_885 (.in({n12933_0, n12932_0, n12929_0, n12928_1/**/, n12921_0, n12920_1}), .out(n2080), .config_in(config_chain[2657:2655]), .config_rst(config_rst)); 
mux6 mux_886 (.in({n11321_1, n11320_0, n11313_1, n11312_0, n11289_0, n11288_0}), .out(n2081), .config_in(config_chain[2660:2658]), .config_rst(config_rst)); 
mux6 mux_887 (.in({n12725_0, n12724_0, n12713_0/**/, n12712_0, n12657_0, n12656_1}), .out(n2082), .config_in(config_chain[2663:2661]), .config_rst(config_rst)); 
mux6 mux_888 (.in({n11553_0, n11552_0, n11521_0, n11520_0, n11491_0, n11490_0}), .out(n2083), .config_in(config_chain[2666:2664]), .config_rst(config_rst)); 
mux6 mux_889 (.in({n12961_0/**/, n12960_0, n12953_0, n12952_0, n12949_0, n12948_0}), .out(n2084), .config_in(config_chain[2669:2667]), .config_rst(config_rst)); 
mux6 mux_890 (.in({n11329_1, n11328_0, n11253_0, n11252_0, n11231_0, n11230_0}), .out(n2085), .config_in(config_chain[2672:2670]), .config_rst(config_rst)); 
mux6 mux_891 (.in({n12679_0, n12678_0, n12673_0/**/, n12672_1, n12665_0, n12664_1}), .out(n2086), .config_in(config_chain[2675:2673]), .config_rst(config_rst)); 
mux6 mux_892 (.in({n11587_1, n11586_0, n11579_1, n11578_0, n11555_0, n11554_0}), .out(n2087), .config_in(config_chain[2678:2676]), .config_rst(config_rst)); 
mux6 mux_893 (.in({n12983_0, n12982_0, n12969_0/**/, n12968_0, n12915_0, n12914_1}), .out(n2088), .config_in(config_chain[2681:2679]), .config_rst(config_rst)); 
mux6 mux_894 (.in({n11285_0, n11284_0/**/, n11263_0, n11262_0, n11233_0, n11232_0}), .out(n2089), .config_in(config_chain[2684:2682]), .config_rst(config_rst)); 
mux6 mux_895 (.in({n12699_0, n12698_0, n12695_0, n12694_0/**/, n12687_0, n12686_0}), .out(n2090), .config_in(config_chain[2687:2685]), .config_rst(config_rst)); 
mux6 mux_896 (.in({n11595_1, n11594_0, n11527_0/**/, n11526_0, n11495_0, n11494_0}), .out(n2091), .config_in(config_chain[2690:2688]), .config_rst(config_rst)); 
mux6 mux_897 (.in({n12991_0/**/, n12990_0, n12935_0, n12934_0, n12923_0, n12922_1}), .out(n2092), .config_in(config_chain[2693:2691]), .config_rst(config_rst)); 
mux6 mux_898 (.in({n11315_1, n11314_0, n11297_0, n11296_0, n11265_0, n11264_0}), .out(n2093), .config_in(config_chain[2696:2694]), .config_rst(config_rst)); 
mux6 mux_899 (.in({n12727_0, n12726_0/**/, n12719_0, n12718_0, n12715_0, n12714_0}), .out(n2094), .config_in(config_chain[2699:2697]), .config_rst(config_rst)); 
mux6 mux_900 (.in({n11559_0, n11558_0, n11529_0, n11528_0, n11499_0, n11498_0}), .out(n2095), .config_in(config_chain[2702:2700]), .config_rst(config_rst)); 
mux6 mux_901 (.in({n12955_0, n12954_0, n12951_0, n12950_0, n12943_0, n12942_0}), .out(n2096), .config_in(config_chain[2705:2703]), .config_rst(config_rst)); 
mux6 mux_902 (.in({n11331_1, n11330_0, n11261_0, n11260_0, n11229_0, n11228_0}), .out(n2097), .config_in(config_chain[2708:2706]), .config_rst(config_rst)); 
mux6 mux_903 (.in({n12735_0, n12734_0, n12667_0, n12666_1, n12659_0/**/, n12658_1}), .out(n2098), .config_in(config_chain[2711:2709]), .config_rst(config_rst)); 
mux6 mux_904 (.in({n11581_1, n11580_0, n11561_0, n11560_0/**/, n11531_0, n11530_0}), .out(n2099), .config_in(config_chain[2714:2712]), .config_rst(config_rst)); 
mux6 mux_905 (.in({n12977_0, n12976_0, n12971_0, n12970_0, n12963_0, n12962_0}), .out(n2100), .config_in(config_chain[2717:2715]), .config_rst(config_rst)); 
mux6 mux_906 (.in({n11293_0, n11292_0, n11271_0, n11270_0, n11239_0/**/, n11238_0}), .out(n2101), .config_in(config_chain[2720:2718]), .config_rst(config_rst)); 
mux6 mux_907 (.in({n12701_0, n12700_0, n12689_0, n12688_0, n12675_0, n12674_1}), .out(n2102), .config_in(config_chain[2723:2721]), .config_rst(config_rst)); 
mux6 mux_908 (.in({n11589_1, n11588_0, n11573_1, n11572_0, n11503_0/**/, n11502_0}), .out(n2103), .config_in(config_chain[2726:2724]), .config_rst(config_rst)); 
mux6 mux_909 (.in({n12925_0, n12924_1, n12917_0, n12916_1, n12869_0/**/, n12868_2}), .out(n2104), .config_in(config_chain[2729:2727]), .config_rst(config_rst)); 
mux6 mux_910 (.in({n11317_1, n11316_0, n11311_1, n11310_0, n11273_0, n11272_0}), .out(n2105), .config_in(config_chain[2732:2730]), .config_rst(config_rst)); 
mux6 mux_911 (.in({n12721_0, n12720_0/**/, n12709_0, n12708_0, n12615_0, n12614_2}), .out(n2106), .config_in(config_chain[2735:2733]), .config_rst(config_rst)); 
mux6 mux_912 (.in({n11575_1, n11574_0, n11535_0/**/, n11534_0, n11505_0, n11504_0}), .out(n2107), .config_in(config_chain[2738:2736]), .config_rst(config_rst)); 
mux6 mux_913 (.in({n12945_0, n12944_0, n12937_0, n12936_0, n12871_0, n12870_2}), .out(n2108), .config_in(config_chain[2741:2739]), .config_rst(config_rst)); 
mux6 mux_914 (.in({n11325_1, n11324_0, n11301_0, n11300_0, n11237_0/**/, n11236_0}), .out(n2109), .config_in(config_chain[2744:2742]), .config_rst(config_rst)); 
mux6 mux_915 (.in({n12729_0, n12728_0, n12661_0, n12660_1/**/, n12607_0, n12606_2}), .out(n2110), .config_in(config_chain[2747:2745]), .config_rst(config_rst)); 
mux6 mux_916 (.in({n11597_2, n11596_0, n11539_0, n11538_0, n11507_0, n11506_0/**/}), .out(n2111), .config_in(config_chain[2750:2748]), .config_rst(config_rst)); 
mux6 mux_917 (.in({n12993_0, n12992_0, n12979_0/**/, n12978_0, n12965_0, n12964_0}), .out(n2112), .config_in(config_chain[2753:2751]), .config_rst(config_rst)); 
mux6 mux_918 (.in({n11305_0, n11304_0, n11269_0, n11268_0/**/, n11247_0, n11246_0}), .out(n2113), .config_in(config_chain[2756:2754]), .config_rst(config_rst)); 
mux6 mux_919 (.in({n12691_0, n12690_0, n12683_0, n12682_0, n12609_0, n12608_2}), .out(n2114), .config_in(config_chain[2759:2757]), .config_rst(config_rst)); 
mux6 mux_920 (.in({n11591_1, n11590_0, n11583_1, n11582_0, n11567_0, n11566_0}), .out(n2115), .config_in(config_chain[2762:2760]), .config_rst(config_rst)); 
mux6 mux_921 (.in({n12987_0, n12986_0, n12919_0, n12918_1, n12863_0/**/, n12862_2}), .out(n2116), .config_in(config_chain[2765:2763]), .config_rst(config_rst)); 
mux6 mux_922 (.in({n11307_1, n11306_0, n11279_0, n11278_0, n11249_0, n11248_0}), .out(n2117), .config_in(config_chain[2768:2766]), .config_rst(config_rst)); 
mux6 mux_923 (.in({n12711_0, n12710_0, n12703_0, n12702_0/**/, n12611_0, n12610_2}), .out(n2118), .config_in(config_chain[2771:2769]), .config_rst(config_rst)); 
mux6 mux_924 (.in({n11569_0, n11568_0, n11543_0, n11542_0, n11513_0, n11512_0}), .out(n2119), .config_in(config_chain[2774:2772]), .config_rst(config_rst)); 
mux6 mux_925 (.in({n12939_0, n12938_0, n12927_0/**/, n12926_1, n12867_0, n12866_2}), .out(n2120), .config_in(config_chain[2777:2775]), .config_rst(config_rst)); 
mux6 mux_926 (.in({n11327_1, n11326_0, n11319_1, n11318_0, n11309_1, n11308_0}), .out(n2121), .config_in(config_chain[2780:2778]), .config_rst(config_rst)); 
mux6 mux_927 (.in({n12731_0, n12730_0, n12663_0/**/, n12662_1, n12613_0, n12612_2}), .out(n2122), .config_in(config_chain[2783:2781]), .config_rst(config_rst)); 
mux6 mux_928 (.in({n11855_1, n11854_0, n11777_0, n11776_0, n11755_0, n11754_0}), .out(n2169), .config_in(config_chain[2786:2784]), .config_rst(config_rst)); 
mux6 mux_929 (.in({n13009_0, n13008_0, n12953_0, n12952_0, n12939_0, n12938_1}), .out(n2170), .config_in(config_chain[2789:2787]), .config_rst(config_rst)); 
mux6 mux_930 (.in({n11577_1, n11576_0, n11547_0, n11546_0, n11515_0, n11514_0}), .out(n2171), .config_in(config_chain[2792:2790]), .config_rst(config_rst)); 
mux6 mux_931 (.in({n12745_0, n12744_0, n12737_0, n12736_0, n12731_0, n12730_0}), .out(n2172), .config_in(config_chain[2795:2793]), .config_rst(config_rst)); 
mux6 mux_932 (.in({n11809_0, n11808_0, n11787_0, n11786_0, n11749_0, n11748_0/**/}), .out(n2173), .config_in(config_chain[2798:2796]), .config_rst(config_rst)); 
mux6 mux_933 (.in({n12973_0, n12972_0, n12969_0, n12968_0, n12961_0, n12960_0}), .out(n2174), .config_in(config_chain[2801:2799]), .config_rst(config_rst)); 
mux6 mux_934 (.in({n11593_1, n11592_0, n11519_0, n11518_0, n11487_0, n11486_0}), .out(n2175), .config_in(config_chain[2804:2802]), .config_rst(config_rst)); 
mux6 mux_935 (.in({n12753_0, n12752_0/**/, n12697_0, n12696_0, n12685_0, n12684_1}), .out(n2176), .config_in(config_chain[2807:2805]), .config_rst(config_rst)); 
mux6 mux_936 (.in({n11841_1, n11840_0, n11813_0, n11812_0/**/, n11781_0, n11780_0}), .out(n2177), .config_in(config_chain[2810:2808]), .config_rst(config_rst)); 
mux6 mux_937 (.in({n12995_0/**/, n12994_0, n12989_0, n12988_0, n12981_0, n12980_0}), .out(n2178), .config_in(config_chain[2813:2811]), .config_rst(config_rst)); 
mux6 mux_938 (.in({n11551_0, n11550_0, n11521_0, n11520_0, n11489_0, n11488_0}), .out(n2179), .config_in(config_chain[2816:2814]), .config_rst(config_rst)); 
mux6 mux_939 (.in({n12717_0, n12716_0, n12705_0, n12704_0, n12693_0, n12692_1}), .out(n2180), .config_in(config_chain[2819:2817]), .config_rst(config_rst)); 
mux6 mux_940 (.in({n11857_1, n11856_0, n11849_1, n11848_0, n11753_0, n11752_0}), .out(n2181), .config_in(config_chain[2822:2820]), .config_rst(config_rst)); 
mux6 mux_941 (.in({n13011_0, n13010_0, n12941_0, n12940_1, n12933_0, n12932_1}), .out(n2182), .config_in(config_chain[2825:2823]), .config_rst(config_rst)); 
mux6 mux_942 (.in({n11579_1, n11578_0, n11553_0, n11552_0, n11523_0, n11522_0}), .out(n2183), .config_in(config_chain[2828:2826]), .config_rst(config_rst)); 
mux6 mux_943 (.in({n12739_0, n12738_0, n12733_0, n12732_0, n12725_0, n12724_0/**/}), .out(n2184), .config_in(config_chain[2831:2829]), .config_rst(config_rst)); 
mux6 mux_944 (.in({n11817_0, n11816_0, n11795_0, n11794_0, n11763_0/**/, n11762_0}), .out(n2185), .config_in(config_chain[2834:2832]), .config_rst(config_rst)); 
mux6 mux_945 (.in({n12975_0, n12974_0/**/, n12963_0, n12962_0, n12949_0, n12948_1}), .out(n2186), .config_in(config_chain[2837:2835]), .config_rst(config_rst)); 
mux6 mux_946 (.in({n11587_1, n11586_0, n11555_0, n11554_0, n11495_0, n11494_0}), .out(n2187), .config_in(config_chain[2840:2838]), .config_rst(config_rst)); 
mux6 mux_947 (.in({n12755_0, n12754_0, n12747_0, n12746_0, n12679_0/**/, n12678_1}), .out(n2188), .config_in(config_chain[2843:2841]), .config_rst(config_rst)); 
mux6 mux_948 (.in({n11827_0, n11826_0, n11789_0, n11788_0, n11757_0, n11756_0}), .out(n2189), .config_in(config_chain[2846:2844]), .config_rst(config_rst)); 
mux6 mux_949 (.in({n12997_0, n12996_0, n12983_0, n12982_0, n12971_0, n12970_0}), .out(n2190), .config_in(config_chain[2849:2847]), .config_rst(config_rst)); 
mux6 mux_950 (.in({n11559_0, n11558_0/**/, n11527_0, n11526_0, n11497_0, n11496_0}), .out(n2191), .config_in(config_chain[2852:2850]), .config_rst(config_rst)); 
mux6 mux_951 (.in({n12707_0, n12706_0, n12699_0, n12698_0, n12695_0, n12694_1/**/}), .out(n2192), .config_in(config_chain[2855:2853]), .config_rst(config_rst)); 
mux6 mux_952 (.in({n11851_1, n11850_0, n11821_0, n11820_0, n11761_0, n11760_0}), .out(n2193), .config_in(config_chain[2858:2856]), .config_rst(config_rst)); 
mux6 mux_953 (.in({n13013_0/**/, n13012_0, n13005_0, n13004_0, n12935_0, n12934_1}), .out(n2194), .config_in(config_chain[2861:2859]), .config_rst(config_rst)); 
mux6 mux_954 (.in({n11561_0/**/, n11560_0, n11531_0, n11530_0, n11499_0, n11498_0}), .out(n2195), .config_in(config_chain[2864:2862]), .config_rst(config_rst)); 
mux6 mux_955 (.in({n12727_0, n12726_0, n12719_0, n12718_0, n12715_0, n12714_0}), .out(n2196), .config_in(config_chain[2867:2865]), .config_rst(config_rst)); 
mux6 mux_956 (.in({n11859_1, n11858_0, n11793_0, n11792_0, n11771_0, n11770_0}), .out(n2197), .config_in(config_chain[2870:2868]), .config_rst(config_rst)); 
mux6 mux_957 (.in({n12957_0, n12956_0, n12951_0, n12950_1/**/, n12943_0, n12942_1}), .out(n2198), .config_in(config_chain[2873:2871]), .config_rst(config_rst)); 
mux6 mux_958 (.in({n11589_1, n11588_0, n11581_1, n11580_0, n11563_0, n11562_0}), .out(n2199), .config_in(config_chain[2876:2874]), .config_rst(config_rst)); 
mux6 mux_959 (.in({n12749_0, n12748_0, n12735_0, n12734_0/**/, n12681_0, n12680_1}), .out(n2200), .config_in(config_chain[2879:2877]), .config_rst(config_rst)); 
mux6 mux_960 (.in({n11835_0, n11834_0, n11803_0, n11802_0, n11765_0, n11764_0}), .out(n2201), .config_in(config_chain[2882:2880]), .config_rst(config_rst)); 
mux6 mux_961 (.in({n12985_0, n12984_0, n12977_0/**/, n12976_0, n12867_0, n12866_2}), .out(n2202), .config_in(config_chain[2885:2883]), .config_rst(config_rst)); 
mux6 mux_962 (.in({n11573_1/**/, n11572_0, n11535_0, n11534_0, n11505_0, n11504_0}), .out(n2203), .config_in(config_chain[2888:2886]), .config_rst(config_rst)); 
mux6 mux_963 (.in({n12701_0, n12700_0, n12689_0, n12688_1, n12613_0, n12612_2}), .out(n2204), .config_in(config_chain[2891:2889]), .config_rst(config_rst)); 
mux6 mux_964 (.in({n11845_1, n11844_0/**/, n11837_0, n11836_0, n11797_0, n11796_0}), .out(n2205), .config_in(config_chain[2894:2892]), .config_rst(config_rst)); 
mux6 mux_965 (.in({n13007_0, n13006_0, n12999_0, n12998_0, n12869_0, n12868_2}), .out(n2206), .config_in(config_chain[2897:2895]), .config_rst(config_rst)); 
mux6 mux_966 (.in({n11575_1, n11574_0, n11537_0, n11536_0, n11507_0, n11506_0}), .out(n2207), .config_in(config_chain[2900:2898]), .config_rst(config_rst)); 
mux6 mux_967 (.in({n12757_0, n12756_0, n12721_0/**/, n12720_0, n12709_0, n12708_0}), .out(n2208), .config_in(config_chain[2903:2901]), .config_rst(config_rst)); 
mux6 mux_968 (.in({n11839_1, n11838_0, n11801_0, n11800_0, n11769_0/**/, n11768_0}), .out(n2209), .config_in(config_chain[2906:2904]), .config_rst(config_rst)); 
mux6 mux_969 (.in({n12959_0, n12958_0, n12945_0, n12944_1, n12871_0, n12870_2}), .out(n2210), .config_in(config_chain[2909:2907]), .config_rst(config_rst)); 
mux6 mux_970 (.in({n11583_1, n11582_0, n11567_0, n11566_0, n11539_0, n11538_0/**/}), .out(n2211), .config_in(config_chain[2912:2910]), .config_rst(config_rst)); 
mux6 mux_971 (.in({n12751_0, n12750_0, n12743_0, n12742_0, n12607_0, n12606_2}), .out(n2212), .config_in(config_chain[2915:2913]), .config_rst(config_rst)); 
mux6 mux_972 (.in({n11829_2, n11828_0, n11811_0, n11810_0, n11779_0, n11778_0}), .out(n2213), .config_in(config_chain[2918:2916]), .config_rst(config_rst)); 
mux6 mux_973 (.in({n12993_0, n12992_0, n12979_0/**/, n12978_0, n12967_0, n12966_0}), .out(n2214), .config_in(config_chain[2921:2919]), .config_rst(config_rst)); 
mux6 mux_974 (.in({n11591_1, n11590_0, n11569_0/**/, n11568_0, n11511_0, n11510_0}), .out(n2215), .config_in(config_chain[2924:2922]), .config_rst(config_rst)); 
mux6 mux_975 (.in({n12691_0, n12690_1, n12683_0, n12682_1, n12609_0, n12608_2}), .out(n2216), .config_in(config_chain[2927:2925]), .config_rst(config_rst)); 
mux6 mux_976 (.in({n11861_2, n11860_0, n11847_1, n11846_0, n11805_0, n11804_0}), .out(n2217), .config_in(config_chain[2930:2928]), .config_rst(config_rst)); 
mux6 mux_977 (.in({n13001_0, n13000_0/**/, n12987_0, n12986_0, n12865_0, n12864_2}), .out(n2218), .config_in(config_chain[2933:2931]), .config_rst(config_rst)); 
mux6 mux_978 (.in({n11571_0, n11570_0, n11545_0, n11544_0, n11513_0, n11512_0}), .out(n2219), .config_in(config_chain[2936:2934]), .config_rst(config_rst)); 
mux6 mux_979 (.in({n12723_0, n12722_0, n12711_0, n12710_0, n12611_0, n12610_2}), .out(n2220), .config_in(config_chain[2939:2937]), .config_rst(config_rst)); 
mux6 mux_980 (.in({n12103_1, n12102_0, n12067_0, n12066_0, n12037_0, n12036_0}), .out(n2267), .config_in(config_chain[2942:2940]), .config_rst(config_rst)); 
mux6 mux_981 (.in({n13017_0, n13016_0, n13001_0, n13000_0, n12987_0, n12986_0}), .out(n2268), .config_in(config_chain[2945:2943]), .config_rst(config_rst)); 
mux6 mux_982 (.in({n11809_0, n11808_0, n11777_0, n11776_0, n11755_0, n11754_0}), .out(n2269), .config_in(config_chain[2948:2946]), .config_rst(config_rst)); 
mux6 mux_983 (.in({n12725_0, n12724_0/**/, n12717_0, n12716_0, n12711_0, n12710_1}), .out(n2270), .config_in(config_chain[2951:2949]), .config_rst(config_rst)); 
mux6 mux_984 (.in({n12111_1, n12110_0, n12069_0, n12068_0, n12017_0, n12016_0}), .out(n2271), .config_in(config_chain[2954:2952]), .config_rst(config_rst)); 
mux6 mux_985 (.in({n13033_0, n13032_0, n13025_0, n13024_0, n12953_0, n12952_1}), .out(n2272), .config_in(config_chain[2957:2955]), .config_rst(config_rst)); 
mux6 mux_986 (.in({n11819_0, n11818_0, n11781_0, n11780_0, n11749_0, n11748_0}), .out(n2273), .config_in(config_chain[2960:2958]), .config_rst(config_rst)); 
mux6 mux_987 (.in({n12759_0, n12758_0, n12745_0, n12744_0, n12733_0, n12732_0}), .out(n2274), .config_in(config_chain[2963:2961]), .config_rst(config_rst)); 
mux6 mux_988 (.in({n12081_0, n12080_0, n12049_0, n12048_0, n12011_0, n12010_0}), .out(n2275), .config_in(config_chain[2966:2964]), .config_rst(config_rst)); 
mux6 mux_989 (.in({n12973_0, n12972_0, n12969_0, n12968_1, n12961_0, n12960_1}), .out(n2276), .config_in(config_chain[2969:2967]), .config_rst(config_rst)); 
mux6 mux_990 (.in({n11849_1, n11848_0, n11841_1, n11840_0, n11813_0, n11812_0}), .out(n2277), .config_in(config_chain[2972:2970]), .config_rst(config_rst)); 
mux6 mux_991 (.in({n12767_0, n12766_0, n12753_0, n12752_0, n12697_0, n12696_1}), .out(n2278), .config_in(config_chain[2975:2973]), .config_rst(config_rst)); 
mux6 mux_992 (.in({n12075_0, n12074_0, n12043_0, n12042_0/**/, n12013_0, n12012_0}), .out(n2279), .config_in(config_chain[2978:2976]), .config_rst(config_rst)); 
mux6 mux_993 (.in({n13003_0, n13002_0, n12995_0, n12994_0, n12989_0, n12988_0}), .out(n2280), .config_in(config_chain[2981:2979]), .config_rst(config_rst)); 
mux6 mux_994 (.in({n11857_1, n11856_0, n11785_0, n11784_0, n11763_0, n11762_0}), .out(n2281), .config_in(config_chain[2984:2982]), .config_rst(config_rst)); 
mux6 mux_995 (.in({n12719_0, n12718_0, n12713_0, n12712_1/**/, n12705_0, n12704_1}), .out(n2282), .config_in(config_chain[2987:2985]), .config_rst(config_rst)); 
mux6 mux_996 (.in({n12113_1, n12112_0, n12105_1, n12104_0/**/, n12077_0, n12076_0}), .out(n2283), .config_in(config_chain[2990:2988]), .config_rst(config_rst)); 
mux6 mux_997 (.in({n13027_0, n13026_0, n13011_0, n13010_0, n12955_0, n12954_1}), .out(n2284), .config_in(config_chain[2993:2991]), .config_rst(config_rst)); 
mux6 mux_998 (.in({n11817_0/**/, n11816_0, n11795_0, n11794_0, n11757_0, n11756_0}), .out(n2285), .config_in(config_chain[2996:2994]), .config_rst(config_rst)); 
mux6 mux_999 (.in({n12739_0/**/, n12738_0, n12735_0, n12734_0, n12727_0, n12726_0}), .out(n2286), .config_in(config_chain[2999:2997]), .config_rst(config_rst)); 
mux6 mux_1000 (.in({n12121_1, n12120_0, n12057_0, n12056_0, n12025_0/**/, n12024_0}), .out(n2287), .config_in(config_chain[3002:3000]), .config_rst(config_rst)); 
mux6 mux_1001 (.in({n13035_0, n13034_0, n12975_0, n12974_0, n12963_0, n12962_1}), .out(n2288), .config_in(config_chain[3005:3003]), .config_rst(config_rst)); 
mux6 mux_1002 (.in({n11843_1, n11842_0, n11821_0, n11820_0, n11789_0, n11788_0/**/}), .out(n2289), .config_in(config_chain[3008:3006]), .config_rst(config_rst)); 
mux6 mux_1003 (.in({n12769_0, n12768_0, n12761_0, n12760_0, n12755_0, n12754_0}), .out(n2290), .config_in(config_chain[3011:3009]), .config_rst(config_rst)); 
mux6 mux_1004 (.in({n12089_0, n12088_0, n12051_0, n12050_0, n12021_0, n12020_0}), .out(n2291), .config_in(config_chain[3014:3012]), .config_rst(config_rst)); 
mux6 mux_1005 (.in({n12997_0, n12996_0, n12991_0, n12990_0, n12983_0, n12982_0}), .out(n2292), .config_in(config_chain[3017:3015]), .config_rst(config_rst)); 
mux6 mux_1006 (.in({n11859_1/**/, n11858_0, n11793_0, n11792_0, n11761_0, n11760_0}), .out(n2293), .config_in(config_chain[3020:3018]), .config_rst(config_rst)); 
mux6 mux_1007 (.in({n12777_0, n12776_0, n12707_0, n12706_1/**/, n12699_0, n12698_1}), .out(n2294), .config_in(config_chain[3023:3021]), .config_rst(config_rst)); 
mux6 mux_1008 (.in({n12107_1, n12106_0, n12083_0/**/, n12082_0, n12053_0, n12052_0}), .out(n2295), .config_in(config_chain[3026:3024]), .config_rst(config_rst)); 
mux6 mux_1009 (.in({n13021_0, n13020_0/**/, n13013_0, n13012_0, n13005_0, n13004_0}), .out(n2296), .config_in(config_chain[3029:3027]), .config_rst(config_rst)); 
mux6 mux_1010 (.in({n11825_0, n11824_0/**/, n11803_0, n11802_0, n11771_0, n11770_0}), .out(n2297), .config_in(config_chain[3032:3030]), .config_rst(config_rst)); 
mux6 mux_1011 (.in({n12741_0, n12740_0, n12729_0, n12728_0, n12715_0, n12714_1}), .out(n2298), .config_in(config_chain[3035:3033]), .config_rst(config_rst)); 
mux6 mux_1012 (.in({n12123_2, n12122_0, n12115_1, n12114_0, n12033_0, n12032_0}), .out(n2299), .config_in(config_chain[3038:3036]), .config_rst(config_rst)); 
mux6 mux_1013 (.in({n13037_0, n13036_0, n12965_0, n12964_1, n12957_0, n12956_1/**/}), .out(n2300), .config_in(config_chain[3041:3039]), .config_rst(config_rst)); 
mux6 mux_1014 (.in({n11845_1, n11844_0, n11835_0, n11834_0, n11797_0/**/, n11796_0}), .out(n2301), .config_in(config_chain[3044:3042]), .config_rst(config_rst)); 
mux6 mux_1015 (.in({n12763_0, n12762_0, n12749_0, n12748_0, n12611_0, n12610_2}), .out(n2302), .config_in(config_chain[3047:3045]), .config_rst(config_rst)); 
mux6 mux_1016 (.in({n12097_0, n12096_0, n12065_0, n12064_0, n12027_0/**/, n12026_0}), .out(n2303), .config_in(config_chain[3050:3048]), .config_rst(config_rst)); 
mux6 mux_1017 (.in({n12985_0, n12984_0, n12977_0, n12976_0/**/, n12867_0, n12866_2}), .out(n2304), .config_in(config_chain[3053:3051]), .config_rst(config_rst)); 
mux6 mux_1018 (.in({n11853_1, n11852_0, n11837_0, n11836_0, n11769_0, n11768_0}), .out(n2305), .config_in(config_chain[3056:3054]), .config_rst(config_rst)); 
mux6 mux_1019 (.in({n12771_0, n12770_0, n12701_0, n12700_1, n12615_0, n12614_2}), .out(n2306), .config_in(config_chain[3059:3057]), .config_rst(config_rst)); 
mux6 mux_1020 (.in({n12099_0, n12098_0, n12061_0, n12060_0, n12029_0, n12028_0}), .out(n2307), .config_in(config_chain[3062:3060]), .config_rst(config_rst)); 
mux6 mux_1021 (.in({n13023_0, n13022_0, n13007_0, n13006_0, n12869_0, n12868_2}), .out(n2308), .config_in(config_chain[3065:3063]), .config_rst(config_rst)); 
mux6 mux_1022 (.in({n11829_2, n11828_0, n11801_0, n11800_0, n11779_0/**/, n11778_0}), .out(n2309), .config_in(config_chain[3068:3066]), .config_rst(config_rst)); 
mux6 mux_1023 (.in({n12757_0, n12756_0, n12731_0, n12730_0, n12723_0, n12722_0/**/}), .out(n2310), .config_in(config_chain[3071:3069]), .config_rst(config_rst)); 
mux6 mux_1024 (.in({n12117_1, n12116_0, n12109_1, n12108_0, n12101_0, n12100_0}), .out(n2311), .config_in(config_chain[3074:3072]), .config_rst(config_rst)); 
mux6 mux_1025 (.in({n13031_0, n13030_0/**/, n12959_0, n12958_1, n12871_0, n12870_2}), .out(n2312), .config_in(config_chain[3077:3075]), .config_rst(config_rst)); 
mux6 mux_1026 (.in({n11861_2, n11860_0, n11811_0, n11810_0, n11773_0, n11772_0}), .out(n2313), .config_in(config_chain[3080:3078]), .config_rst(config_rst)); 
mux6 mux_1027 (.in({n12779_0, n12778_0, n12751_0, n12750_0, n12743_0, n12742_0}), .out(n2314), .config_in(config_chain[3083:3081]), .config_rst(config_rst)); 
mux6 mux_1028 (.in({n12091_2, n12090_0, n12073_0, n12072_0, n12035_0, n12034_0}), .out(n2315), .config_in(config_chain[3086:3084]), .config_rst(config_rst)); 
mux6 mux_1029 (.in({n13015_0, n13014_0, n12979_0, n12978_0/**/, n12967_0, n12966_1}), .out(n2316), .config_in(config_chain[3089:3087]), .config_rst(config_rst)); 
mux6 mux_1030 (.in({n11855_1, n11854_0/**/, n11847_1, n11846_0, n11833_0, n11832_0}), .out(n2317), .config_in(config_chain[3092:3090]), .config_rst(config_rst)); 
mux6 mux_1031 (.in({n12773_0, n12772_0/**/, n12703_0, n12702_1, n12609_0, n12608_2}), .out(n2318), .config_in(config_chain[3095:3093]), .config_rst(config_rst)); 
mux6 mux_1032 (.in({n12111_1, n12110_0, n12103_1, n12102_0, n12069_0, n12068_0}), .out(n2364), .config_in(config_chain[3098:3096]), .config_rst(config_rst)); 
mux6 mux_1033 (.in({n12081_0, n12080_0, n12043_0, n12042_0, n12011_0, n12010_0}), .out(n2367), .config_in(config_chain[3101:3099]), .config_rst(config_rst)); 
mux6 mux_1034 (.in({n12113_1, n12112_0, n12105_1, n12104_0, n12077_0, n12076_0}), .out(n2370), .config_in(config_chain[3104:3102]), .config_rst(config_rst)); 
mux6 mux_1035 (.in({n12089_0, n12088_0, n12051_0, n12050_0, n12019_0, n12018_0}), .out(n2373), .config_in(config_chain[3107:3105]), .config_rst(config_rst)); 
mux6 mux_1036 (.in({n12107_1, n12106_0, n12085_0, n12084_0, n12053_0, n12052_0}), .out(n2376), .config_in(config_chain[3110:3108]), .config_rst(config_rst)); 
mux6 mux_1037 (.in({n12097_0, n12096_0, n12065_0, n12064_0, n12027_0, n12026_0}), .out(n2379), .config_in(config_chain[3113:3111]), .config_rst(config_rst)); 
mux6 mux_1038 (.in({n12109_1, n12108_0, n12101_0, n12100_0, n12061_0, n12060_0}), .out(n2382), .config_in(config_chain[3116:3114]), .config_rst(config_rst)); 
mux6 mux_1039 (.in({n12093_2, n12092_0, n12073_0, n12072_0, n12035_0, n12034_0}), .out(n2385), .config_in(config_chain[3119:3117]), .config_rst(config_rst)); 
mux6 mux_1040 (.in({n9779_1, n9778_0, n9765_0, n9764_0, n9723_0, n9722_0}), .out(n2412), .config_in(config_chain[3122:3120]), .config_rst(config_rst)); 
mux6 mux_1041 (.in({n9795_1, n9794_0, n9705_0, n9704_0, n9673_0, n9672_0}), .out(n2415), .config_in(config_chain[3125:3123]), .config_rst(config_rst)); 
mux6 mux_1042 (.in({n9767_0, n9766_0, n9759_0, n9758_0, n9731_0, n9730_0}), .out(n2418), .config_in(config_chain[3128:3126]), .config_rst(config_rst)); 
mux6 mux_1043 (.in({n9797_1, n9796_0, n9713_0, n9712_0, n9681_0, n9680_0}), .out(n2421), .config_in(config_chain[3131:3129]), .config_rst(config_rst)); 
mux6 mux_1044 (.in({n9769_0, n9768_0, n9761_0, n9760_0, n9739_0, n9738_0}), .out(n2424), .config_in(config_chain[3134:3132]), .config_rst(config_rst)); 
mux6 mux_1045 (.in({n9791_1, n9790_0, n9755_2, n9754_0, n9689_0, n9688_0}), .out(n2427), .config_in(config_chain[3137:3135]), .config_rst(config_rst)); 
mux6 mux_1046 (.in({n9763_0, n9762_0, n9747_1, n9746_0, n9715_0, n9714_0}), .out(n2430), .config_in(config_chain[3140:3138]), .config_rst(config_rst)); 
mux6 mux_1047 (.in({n9793_1, n9792_0, n9751_2, n9750_0, n9697_0, n9696_0}), .out(n2433), .config_in(config_chain[3143:3141]), .config_rst(config_rst)); 
mux6 mux_1048 (.in({n10047_1, n10046_0, n9945_0, n9944_0, n9923_0, n9922_0}), .out(n2461), .config_in(config_chain[3146:3144]), .config_rst(config_rst)); 
mux6 mux_1049 (.in({n13101_1, n13100_0, n13063_0, n13062_0, n13041_0, n13040_0}), .out(n2462), .config_in(config_chain[3149:3147]), .config_rst(config_rst)); 
mux6 mux_1050 (.in({n9779_1, n9778_0, n9773_0/**/, n9772_0, n9765_0, n9764_0}), .out(n2463), .config_in(config_chain[3152:3150]), .config_rst(config_rst)); 
mux6 mux_1051 (.in({n12839_0, n12838_0, n12817_1, n12816_0, n12785_1, n12784_0}), .out(n2464), .config_in(config_chain[3155:3153]), .config_rst(config_rst)); 
mux6 mux_1052 (.in({n10013_0, n10012_0, n9977_0, n9976_0, n9955_0, n9954_0/**/}), .out(n2465), .config_in(config_chain[3158:3156]), .config_rst(config_rst)); 
mux6 mux_1053 (.in({n13105_0, n13104_0, n13073_0, n13072_0/**/, n13043_0, n13042_0}), .out(n2466), .config_in(config_chain[3161:3159]), .config_rst(config_rst)); 
mux6 mux_1054 (.in({n9795_1, n9794_0, n9705_0, n9704_0, n9673_0, n9672_0}), .out(n2467), .config_in(config_chain[3164:3162]), .config_rst(config_rst)); 
mux6 mux_1055 (.in({n12849_1, n12848_0, n12819_0, n12818_0, n12781_0, n12780_0}), .out(n2468), .config_in(config_chain[3167:3165]), .config_rst(config_rst)); 
mux6 mux_1056 (.in({n10033_1, n10032_0, n10029_0, n10028_0, n10021_0, n10020_0}), .out(n2469), .config_in(config_chain[3170:3168]), .config_rst(config_rst)); 
mux6 mux_1057 (.in({n13107_0, n13106_0, n13075_0, n13074_0, n13045_1, n13044_0}), .out(n2470), .config_in(config_chain[3173:3171]), .config_rst(config_rst)); 
mux6 mux_1058 (.in({n9737_0, n9736_0, n9699_0, n9698_0, n9667_0, n9666_0}), .out(n2471), .config_in(config_chain[3176:3174]), .config_rst(config_rst)); 
mux6 mux_1059 (.in({n12851_0, n12850_0, n12813_0, n12812_0, n12783_0, n12782_0}), .out(n2472), .config_in(config_chain[3179:3177]), .config_rst(config_rst)); 
mux6 mux_1060 (.in({n10049_1, n10048_0, n10041_1, n10040_0, n9921_0, n9920_0}), .out(n2473), .config_in(config_chain[3182:3180]), .config_rst(config_rst)); 
mux6 mux_1061 (.in({n13109_1/**/, n13108_0, n13071_0, n13070_0, n13039_0, n13038_0}), .out(n2474), .config_in(config_chain[3185:3183]), .config_rst(config_rst)); 
mux6 mux_1062 (.in({n9781_1, n9780_0, n9767_0, n9766_0, n9731_0, n9730_0}), .out(n2475), .config_in(config_chain[3188:3186]), .config_rst(config_rst)); 
mux6 mux_1063 (.in({n12847_0, n12846_0, n12815_0, n12814_0, n12793_1, n12792_0}), .out(n2476), .config_in(config_chain[3191:3189]), .config_rst(config_rst)); 
mux6 mux_1064 (.in({n9985_0, n9984_0, n9963_0, n9962_0, n9931_0, n9930_0}), .out(n2477), .config_in(config_chain[3194:3192]), .config_rst(config_rst)); 
mux6 mux_1065 (.in({n13103_0, n13102_0, n13081_0, n13080_0, n13051_0, n13050_0}), .out(n2478), .config_in(config_chain[3197:3195]), .config_rst(config_rst)); 
mux6 mux_1066 (.in({n9789_1, n9788_0, n9775_0/**/, n9774_0, n9681_0, n9680_0}), .out(n2479), .config_in(config_chain[3200:3198]), .config_rst(config_rst)); 
mux6 mux_1067 (.in({n12857_1, n12856_0, n12825_1, n12824_0, n12795_0, n12794_0}), .out(n2480), .config_in(config_chain[3203:3201]), .config_rst(config_rst)); 
mux6 mux_1068 (.in({n10023_0, n10022_0, n10015_0/**/, n10014_0, n9995_0, n9994_0}), .out(n2481), .config_in(config_chain[3206:3204]), .config_rst(config_rst)); 
mux6 mux_1069 (.in({n13113_0, n13112_0/**/, n13083_0, n13082_0, n13053_1, n13052_0}), .out(n2482), .config_in(config_chain[3209:3207]), .config_rst(config_rst)); 
mux6 mux_1070 (.in({n9745_0/**/, n9744_0, n9713_0, n9712_0, n9675_0, n9674_0}), .out(n2483), .config_in(config_chain[3212:3210]), .config_rst(config_rst)); 
mux6 mux_1071 (.in({n12859_0, n12858_0, n12821_0, n12820_0, n12789_0, n12788_0}), .out(n2484), .config_in(config_chain[3215:3213]), .config_rst(config_rst)); 
mux6 mux_1072 (.in({n10043_1, n10042_0, n10031_0/**/, n10030_0, n9929_0, n9928_0}), .out(n2485), .config_in(config_chain[3218:3216]), .config_rst(config_rst)); 
mux6 mux_1073 (.in({n13117_1, n13116_0, n13085_1, n13084_0/**/, n13047_0, n13046_0}), .out(n2486), .config_in(config_chain[3221:3219]), .config_rst(config_rst)); 
mux6 mux_1074 (.in({n9769_0/**/, n9768_0, n9761_0, n9760_0, n9739_0, n9738_0}), .out(n2487), .config_in(config_chain[3224:3222]), .config_rst(config_rst)); 
mux6 mux_1075 (.in({n12853_0, n12852_0, n12823_0, n12822_0, n12791_0, n12790_0/**/}), .out(n2488), .config_in(config_chain[3227:3225]), .config_rst(config_rst)); 
mux6 mux_1076 (.in({n10051_1, n10050_0, n9961_0, n9960_0, n9939_0, n9938_0}), .out(n2489), .config_in(config_chain[3230:3228]), .config_rst(config_rst)); 
mux6 mux_1077 (.in({n13111_0, n13110_0, n13079_0, n13078_0, n13057_0/**/, n13056_0}), .out(n2490), .config_in(config_chain[3233:3231]), .config_rst(config_rst)); 
mux6 mux_1078 (.in({n9791_1, n9790_0/**/, n9783_1, n9782_0, n9777_0, n9776_0}), .out(n2491), .config_in(config_chain[3236:3234]), .config_rst(config_rst)); 
mux6 mux_1079 (.in({n12855_0, n12854_0, n12833_1, n12832_0, n12803_0, n12802_0}), .out(n2492), .config_in(config_chain[3239:3237]), .config_rst(config_rst)); 
mux6 mux_1080 (.in({n10017_0, n10016_0, n10007_2, n10006_0, n9971_0/**/, n9970_0}), .out(n2493), .config_in(config_chain[3242:3240]), .config_rst(config_rst)); 
mux6 mux_1081 (.in({n13125_2, n13124_0, n13091_0, n13090_0, n13059_0, n13058_0}), .out(n2494), .config_in(config_chain[3245:3243]), .config_rst(config_rst)); 
mux6 mux_1082 (.in({n9755_2, n9754_0, n9721_0, n9720_0, n9683_0/**/, n9682_0}), .out(n2495), .config_in(config_chain[3248:3246]), .config_rst(config_rst)); 
mux6 mux_1083 (.in({n12869_2, n12868_0, n12835_0, n12834_0/**/, n12797_0, n12796_0}), .out(n2496), .config_in(config_chain[3251:3249]), .config_rst(config_rst)); 
mux6 mux_1084 (.in({n10037_1, n10036_0, n10025_0, n10024_0, n10009_2, n10008_0}), .out(n2497), .config_in(config_chain[3254:3252]), .config_rst(config_rst)); 
mux6 mux_1085 (.in({n13127_2, n13126_0, n13093_1, n13092_0, n13061_1, n13060_0}), .out(n2498), .config_in(config_chain[3257:3255]), .config_rst(config_rst)); 
mux6 mux_1086 (.in({n9763_0/**/, n9762_0, n9757_2, n9756_0, n9715_0, n9714_0}), .out(n2499), .config_in(config_chain[3260:3258]), .config_rst(config_rst)); 
mux6 mux_1087 (.in({n12861_1, n12860_0, n12829_0/**/, n12828_0, n12799_0, n12798_0}), .out(n2500), .config_in(config_chain[3263:3261]), .config_rst(config_rst)); 
mux6 mux_1088 (.in({n10011_2, n10010_0, n9969_0, n9968_0/**/, n9937_0, n9936_0}), .out(n2501), .config_in(config_chain[3266:3264]), .config_rst(config_rst)); 
mux6 mux_1089 (.in({n13129_2, n13128_0, n13087_0/**/, n13086_0, n13065_0, n13064_0}), .out(n2502), .config_in(config_chain[3269:3267]), .config_rst(config_rst)); 
mux6 mux_1090 (.in({n9785_1/**/, n9784_0, n9771_0, n9770_0, n9749_2, n9748_0}), .out(n2503), .config_in(config_chain[3272:3270]), .config_rst(config_rst)); 
mux6 mux_1091 (.in({n12863_2, n12862_0, n12841_1, n12840_0, n12809_1, n12808_0}), .out(n2504), .config_in(config_chain[3275:3273]), .config_rst(config_rst)); 
mux6 mux_1092 (.in({n10001_1, n10000_0, n9979_0, n9978_0/**/, n9947_0, n9946_0}), .out(n2505), .config_in(config_chain[3278:3276]), .config_rst(config_rst)); 
mux6 mux_1093 (.in({n13119_1, n13118_0, n13097_0, n13096_0, n13067_0, n13066_0}), .out(n2506), .config_in(config_chain[3281:3279]), .config_rst(config_rst)); 
mux6 mux_1094 (.in({n9793_1, n9792_0, n9751_2, n9750_0, n9697_0/**/, n9696_0}), .out(n2507), .config_in(config_chain[3284:3282]), .config_rst(config_rst)); 
mux6 mux_1095 (.in({n12865_2/**/, n12864_0, n12843_0, n12842_0, n12811_0, n12810_0}), .out(n2508), .config_in(config_chain[3287:3285]), .config_rst(config_rst)); 
mux6 mux_1096 (.in({n10039_1, n10038_0, n10027_0, n10026_0, n10003_1, n10002_0}), .out(n2509), .config_in(config_chain[3290:3288]), .config_rst(config_rst)); 
mux6 mux_1097 (.in({n13123_2, n13122_0, n13099_0/**/, n13098_0, n13069_1, n13068_0}), .out(n2510), .config_in(config_chain[3293:3291]), .config_rst(config_rst)); 
mux6 mux_1098 (.in({n9753_2, n9752_0, n9723_0, n9722_0, n9691_0, n9690_0}), .out(n2511), .config_in(config_chain[3296:3294]), .config_rst(config_rst)); 
mux6 mux_1099 (.in({n12867_2, n12866_0, n12837_0/**/, n12836_0, n12807_0, n12806_0}), .out(n2512), .config_in(config_chain[3299:3297]), .config_rst(config_rst)); 
mux6 mux_1100 (.in({n10289_1, n10288_0, n10275_0, n10274_0, n10237_0, n10236_0}), .out(n2559), .config_in(config_chain[3302:3300]), .config_rst(config_rst)); 
mux6 mux_1101 (.in({n13131_1/**/, n13130_0, n13099_0, n13098_0, n13069_0, n13068_0}), .out(n2560), .config_in(config_chain[3305:3303]), .config_rst(config_rst)); 
mux6 mux_1102 (.in({n9977_0, n9976_0/**/, n9945_0, n9944_0, n9923_0, n9922_0}), .out(n2561), .config_in(config_chain[3308:3306]), .config_rst(config_rst)); 
mux6 mux_1103 (.in({n12837_0, n12836_0, n12815_0, n12814_0, n12783_0, n12782_0}), .out(n2562), .config_in(config_chain[3311:3309]), .config_rst(config_rst)); 
mux6 mux_1104 (.in({n10297_1, n10296_0, n10283_0, n10282_0, n10179_0, n10178_0}), .out(n2563), .config_in(config_chain[3314:3312]), .config_rst(config_rst)); 
mux6 mux_1105 (.in({n13147_1, n13146_0, n13139_1, n13138_0, n13041_0, n13040_0}), .out(n2564), .config_in(config_chain[3317:3315]), .config_rst(config_rst)); 
mux6 mux_1106 (.in({n10021_0, n10020_0, n10013_0, n10012_0, n9987_0, n9986_0}), .out(n2565), .config_in(config_chain[3320:3318]), .config_rst(config_rst)); 
mux6 mux_1107 (.in({n12873_1, n12872_0, n12847_0, n12846_0, n12817_0, n12816_0}), .out(n2566), .config_in(config_chain[3323:3321]), .config_rst(config_rst)); 
mux6 mux_1108 (.in({n10243_0, n10242_0, n10211_0, n10210_0, n10181_0, n10180_0}), .out(n2567), .config_in(config_chain[3326:3324]), .config_rst(config_rst)); 
mux6 mux_1109 (.in({n13105_0, n13104_0, n13073_0, n13072_0, n13043_0, n13042_0}), .out(n2568), .config_in(config_chain[3329:3327]), .config_rst(config_rst)); 
mux6 mux_1110 (.in({n10041_1, n10040_0, n10033_1, n10032_0, n10029_0, n10028_0}), .out(n2569), .config_in(config_chain[3332:3330]), .config_rst(config_rst)); 
mux6 mux_1111 (.in({n12881_1, n12880_0, n12849_0, n12848_0, n12781_0, n12780_0}), .out(n2570), .config_in(config_chain[3335:3333]), .config_rst(config_rst)); 
mux6 mux_1112 (.in({n10269_0, n10268_0, n10245_0, n10244_0, n10213_0, n10212_0}), .out(n2571), .config_in(config_chain[3338:3336]), .config_rst(config_rst)); 
mux6 mux_1113 (.in({n13107_0, n13106_0, n13077_0, n13076_0, n13045_0, n13044_0}), .out(n2572), .config_in(config_chain[3341:3339]), .config_rst(config_rst)); 
mux6 mux_1114 (.in({n10049_1, n10048_0, n9953_0, n9952_0, n9931_0, n9930_0}), .out(n2573), .config_in(config_chain[3344:3342]), .config_rst(config_rst)); 
mux6 mux_1115 (.in({n12845_0, n12844_0, n12813_0/**/, n12812_0, n12791_0, n12790_0}), .out(n2574), .config_in(config_chain[3347:3345]), .config_rst(config_rst)); 
mux6 mux_1116 (.in({n10299_1, n10298_0, n10291_1, n10290_0, n10285_0, n10284_0/**/}), .out(n2575), .config_in(config_chain[3350:3348]), .config_rst(config_rst)); 
mux6 mux_1117 (.in({n13141_1, n13140_0, n13109_0, n13108_0, n13049_0/**/, n13048_0}), .out(n2576), .config_in(config_chain[3353:3351]), .config_rst(config_rst)); 
mux6 mux_1118 (.in({n10015_0, n10014_0, n9985_0/**/, n9984_0, n9963_0, n9962_0}), .out(n2577), .config_in(config_chain[3356:3354]), .config_rst(config_rst)); 
mux6 mux_1119 (.in({n12855_0, n12854_0/**/, n12823_0, n12822_0, n12793_0, n12792_0}), .out(n2578), .config_in(config_chain[3359:3357]), .config_rst(config_rst)); 
mux6 mux_1120 (.in({n10307_1, n10306_0/**/, n10219_0, n10218_0, n10187_0, n10186_0}), .out(n2579), .config_in(config_chain[3362:3360]), .config_rst(config_rst)); 
mux6 mux_1121 (.in({n13149_1, n13148_0, n13081_0, n13080_0, n13051_0, n13050_0}), .out(n2580), .config_in(config_chain[3365:3363]), .config_rst(config_rst)); 
mux6 mux_1122 (.in({n10035_1, n10034_0, n10031_0, n10030_0, n10023_0, n10022_0/**/}), .out(n2581), .config_in(config_chain[3368:3366]), .config_rst(config_rst)); 
mux6 mux_1123 (.in({n12883_1, n12882_0, n12875_1, n12874_0, n12857_0, n12856_0}), .out(n2582), .config_in(config_chain[3371:3369]), .config_rst(config_rst)); 
mux6 mux_1124 (.in({n10271_0, n10270_0, n10251_0, n10250_0/**/, n10221_0, n10220_0}), .out(n2583), .config_in(config_chain[3374:3372]), .config_rst(config_rst)); 
mux6 mux_1125 (.in({n13115_0, n13114_0, n13083_0/**/, n13082_0, n13053_0, n13052_0}), .out(n2584), .config_in(config_chain[3377:3375]), .config_rst(config_rst)); 
mux6 mux_1126 (.in({n10051_1, n10050_0, n9961_0, n9960_0, n9929_0, n9928_0}), .out(n2585), .config_in(config_chain[3380:3378]), .config_rst(config_rst)); 
mux6 mux_1127 (.in({n12891_1, n12890_0, n12821_0, n12820_0, n12789_0, n12788_0/**/}), .out(n2586), .config_in(config_chain[3383:3381]), .config_rst(config_rst)); 
mux6 mux_1128 (.in({n10293_1, n10292_0, n10279_0, n10278_0, n10253_0/**/, n10252_0}), .out(n2587), .config_in(config_chain[3386:3384]), .config_rst(config_rst)); 
mux6 mux_1129 (.in({n13135_1, n13134_0, n13117_0, n13116_0, n13085_0, n13084_0}), .out(n2588), .config_in(config_chain[3389:3387]), .config_rst(config_rst)); 
mux6 mux_1130 (.in({n9993_0, n9992_0, n9971_0, n9970_0, n9939_0, n9938_0/**/}), .out(n2589), .config_in(config_chain[3392:3390]), .config_rst(config_rst)); 
mux6 mux_1131 (.in({n12853_0, n12852_0, n12831_0, n12830_0, n12801_0, n12800_0}), .out(n2590), .config_in(config_chain[3395:3393]), .config_rst(config_rst)); 
mux6 mux_1132 (.in({n10301_1/**/, n10300_0, n10261_1, n10260_0, n10195_0, n10194_0}), .out(n2591), .config_in(config_chain[3398:3396]), .config_rst(config_rst)); 
mux6 mux_1133 (.in({n13123_1, n13122_0, n13089_0, n13088_0/**/, n13057_0, n13056_0}), .out(n2592), .config_in(config_chain[3401:3399]), .config_rst(config_rst)); 
mux6 mux_1134 (.in({n10037_1, n10036_0/**/, n10025_0, n10024_0, n10007_2, n10006_0}), .out(n2593), .config_in(config_chain[3404:3402]), .config_rst(config_rst)); 
mux6 mux_1135 (.in({n12877_1/**/, n12876_0, n12867_2, n12866_0, n12833_0, n12832_0}), .out(n2594), .config_in(config_chain[3407:3405]), .config_rst(config_rst)); 
mux6 mux_1136 (.in({n10263_2, n10262_0, n10227_0, n10226_0, n10197_0, n10196_0}), .out(n2595), .config_in(config_chain[3410:3408]), .config_rst(config_rst)); 
mux6 mux_1137 (.in({n13125_2, n13124_0, n13091_0, n13090_0, n13059_0/**/, n13058_0}), .out(n2596), .config_in(config_chain[3413:3411]), .config_rst(config_rst)); 
mux6 mux_1138 (.in({n10045_1, n10044_0, n10009_2, n10008_0, n9937_0, n9936_0}), .out(n2597), .config_in(config_chain[3416:3414]), .config_rst(config_rst)); 
mux6 mux_1139 (.in({n12885_1, n12884_0, n12871_2, n12870_0, n12797_0, n12796_0}), .out(n2598), .config_in(config_chain[3419:3417]), .config_rst(config_rst)); 
mux6 mux_1140 (.in({n10281_0, n10280_0, n10273_0, n10272_0, n10265_2, n10264_0}), .out(n2599), .config_in(config_chain[3422:3420]), .config_rst(config_rst)); 
mux6 mux_1141 (.in({n13137_1, n13136_0, n13127_2, n13126_0, n13093_0, n13092_0}), .out(n2600), .config_in(config_chain[3425:3423]), .config_rst(config_rst)); 
mux6 mux_1142 (.in({n10001_1, n10000_0, n9969_0, n9968_0/**/, n9947_0, n9946_0}), .out(n2601), .config_in(config_chain[3428:3426]), .config_rst(config_rst)); 
mux6 mux_1143 (.in({n12861_1, n12860_0, n12839_0, n12838_0, n12807_0/**/, n12806_0}), .out(n2602), .config_in(config_chain[3431:3429]), .config_rst(config_rst)); 
mux6 mux_1144 (.in({n10303_1, n10302_0/**/, n10295_1, n10294_0, n10267_2, n10266_0}), .out(n2603), .config_in(config_chain[3434:3432]), .config_rst(config_rst)); 
mux6 mux_1145 (.in({n13145_1, n13144_0, n13129_2, n13128_0, n13065_0, n13064_0}), .out(n2604), .config_in(config_chain[3437:3435]), .config_rst(config_rst)); 
mux6 mux_1146 (.in({n10019_0, n10018_0/**/, n10003_1, n10002_0, n9979_0, n9978_0}), .out(n2605), .config_in(config_chain[3440:3438]), .config_rst(config_rst)); 
mux6 mux_1147 (.in({n12863_1, n12862_0, n12841_0, n12840_0, n12809_0, n12808_0}), .out(n2606), .config_in(config_chain[3443:3441]), .config_rst(config_rst)); 
mux6 mux_1148 (.in({n10257_1, n10256_0, n10235_0, n10234_0, n10205_0, n10204_0}), .out(n2607), .config_in(config_chain[3446:3444]), .config_rst(config_rst)); 
mux6 mux_1149 (.in({n13121_1/**/, n13120_0, n13097_0, n13096_0, n13067_0, n13066_0}), .out(n2608), .config_in(config_chain[3449:3447]), .config_rst(config_rst)); 
mux6 mux_1150 (.in({n10047_1, n10046_0, n10039_1, n10038_0/**/, n10005_2, n10004_0}), .out(n2609), .config_in(config_chain[3452:3450]), .config_rst(config_rst)); 
mux6 mux_1151 (.in({n12887_1, n12886_0, n12865_2, n12864_0, n12805_0, n12804_0}), .out(n2610), .config_in(config_chain[3455:3453]), .config_rst(config_rst)); 
mux6 mux_1152 (.in({n10561_1/**/, n10560_0, n10463_0, n10462_0, n10441_0, n10440_0}), .out(n2657), .config_in(config_chain[3458:3456]), .config_rst(config_rst)); 
mux6 mux_1153 (.in({n13165_1, n13164_0, n13067_0, n13066_0, n13045_0, n13044_0}), .out(n2658), .config_in(config_chain[3461:3459]), .config_rst(config_rst)); 
mux6 mux_1154 (.in({n10289_1, n10288_0, n10283_0, n10282_0, n10275_0, n10274_0}), .out(n2659), .config_in(config_chain[3464:3462]), .config_rst(config_rst)); 
mux6 mux_1155 (.in({n12901_1, n12900_0/**/, n12893_1, n12892_0, n12887_0, n12886_0}), .out(n2660), .config_in(config_chain[3467:3465]), .config_rst(config_rst)); 
mux6 mux_1156 (.in({n10527_0, n10526_0, n10495_0, n10494_0, n10473_0, n10472_0}), .out(n2661), .config_in(config_chain[3470:3468]), .config_rst(config_rst)); 
mux6 mux_1157 (.in({n13131_0, n13130_0, n13109_0, n13108_0, n13077_0, n13076_0}), .out(n2662), .config_in(config_chain[3473:3471]), .config_rst(config_rst)); 
mux6 mux_1158 (.in({n10305_1, n10304_0, n10211_0, n10210_0, n10179_0, n10178_0}), .out(n2663), .config_in(config_chain[3476:3474]), .config_rst(config_rst)); 
mux6 mux_1159 (.in({n12909_1, n12908_0, n12815_0, n12814_0, n12785_0, n12784_0}), .out(n2664), .config_in(config_chain[3479:3477]), .config_rst(config_rst)); 
mux6 mux_1160 (.in({n10547_1, n10546_0, n10543_0, n10542_0, n10535_0, n10534_0}), .out(n2665), .config_in(config_chain[3482:3480]), .config_rst(config_rst)); 
mux6 mux_1161 (.in({n13151_1, n13150_0, n13147_0, n13146_0, n13139_0, n13138_0}), .out(n2666), .config_in(config_chain[3485:3483]), .config_rst(config_rst)); 
mux6 mux_1162 (.in({n10243_0, n10242_0/**/, n10213_0, n10212_0, n10181_0, n10180_0}), .out(n2667), .config_in(config_chain[3488:3486]), .config_rst(config_rst)); 
mux6 mux_1163 (.in({n12873_0, n12872_0, n12847_0, n12846_0, n12817_0, n12816_0}), .out(n2668), .config_in(config_chain[3491:3489]), .config_rst(config_rst)); 
mux6 mux_1164 (.in({n10563_1, n10562_0, n10555_1, n10554_0, n10439_0, n10438_0/**/}), .out(n2669), .config_in(config_chain[3494:3492]), .config_rst(config_rst)); 
mux6 mux_1165 (.in({n13167_1, n13166_0, n13075_0, n13074_0, n13043_0, n13042_0}), .out(n2670), .config_in(config_chain[3497:3495]), .config_rst(config_rst)); 
mux6 mux_1166 (.in({n10291_1, n10290_0, n10277_0, n10276_0, n10245_0/**/, n10244_0}), .out(n2671), .config_in(config_chain[3500:3498]), .config_rst(config_rst)); 
mux6 mux_1167 (.in({n12895_1, n12894_0, n12889_0, n12888_0/**/, n12881_0, n12880_0}), .out(n2672), .config_in(config_chain[3503:3501]), .config_rst(config_rst)); 
mux6 mux_1168 (.in({n10503_0, n10502_0/**/, n10481_0, n10480_0, n10449_0, n10448_0}), .out(n2673), .config_in(config_chain[3506:3504]), .config_rst(config_rst)); 
mux6 mux_1169 (.in({n13133_0/**/, n13132_0, n13107_0, n13106_0, n13085_0, n13084_0}), .out(n2674), .config_in(config_chain[3509:3507]), .config_rst(config_rst)); 
mux6 mux_1170 (.in({n10299_1, n10298_0/**/, n10285_0, n10284_0, n10187_0, n10186_0}), .out(n2675), .config_in(config_chain[3512:3510]), .config_rst(config_rst)); 
mux6 mux_1171 (.in({n12911_1, n12910_0, n12903_1, n12902_0, n12791_0/**/, n12790_0}), .out(n2676), .config_in(config_chain[3515:3513]), .config_rst(config_rst)); 
mux6 mux_1172 (.in({n10537_0/**/, n10536_0, n10529_0, n10528_0, n10513_0, n10512_0}), .out(n2677), .config_in(config_chain[3518:3516]), .config_rst(config_rst)); 
mux6 mux_1173 (.in({n13153_1, n13152_0, n13141_0/**/, n13140_0, n13117_0, n13116_0}), .out(n2678), .config_in(config_chain[3521:3519]), .config_rst(config_rst)); 
mux6 mux_1174 (.in({n10251_0/**/, n10250_0, n10219_0, n10218_0, n10189_0, n10188_0}), .out(n2679), .config_in(config_chain[3524:3522]), .config_rst(config_rst)); 
mux6 mux_1175 (.in({n12855_0, n12854_0, n12825_0, n12824_0, n12793_0, n12792_0}), .out(n2680), .config_in(config_chain[3527:3525]), .config_rst(config_rst)); 
mux6 mux_1176 (.in({n10557_1/**/, n10556_0, n10545_0, n10544_0, n10447_0, n10446_0}), .out(n2681), .config_in(config_chain[3530:3528]), .config_rst(config_rst)); 
mux6 mux_1177 (.in({n13169_1, n13168_0, n13161_1, n13160_0/**/, n13051_0, n13050_0}), .out(n2682), .config_in(config_chain[3533:3531]), .config_rst(config_rst)); 
mux6 mux_1178 (.in({n10279_0, n10278_0, n10271_0, n10270_0/**/, n10253_0, n10252_0}), .out(n2683), .config_in(config_chain[3536:3534]), .config_rst(config_rst)); 
mux6 mux_1179 (.in({n12883_0, n12882_0, n12875_0, n12874_0, n12857_0, n12856_0}), .out(n2684), .config_in(config_chain[3539:3537]), .config_rst(config_rst)); 
mux6 mux_1180 (.in({n10565_1, n10564_0, n10479_0, n10478_0, n10457_0, n10456_0}), .out(n2685), .config_in(config_chain[3542:3540]), .config_rst(config_rst)); 
mux6 mux_1181 (.in({n13115_0, n13114_0, n13083_0, n13082_0/**/, n13061_0, n13060_0}), .out(n2686), .config_in(config_chain[3545:3543]), .config_rst(config_rst)); 
mux6 mux_1182 (.in({n10301_1/**/, n10300_0, n10293_1, n10292_0, n10287_0, n10286_0}), .out(n2687), .config_in(config_chain[3548:3546]), .config_rst(config_rst)); 
mux6 mux_1183 (.in({n12905_1/**/, n12904_0, n12891_0, n12890_0, n12799_0, n12798_0}), .out(n2688), .config_in(config_chain[3551:3549]), .config_rst(config_rst)); 
mux6 mux_1184 (.in({n10531_0, n10530_0, n10517_1, n10516_0, n10489_0, n10488_0/**/}), .out(n2689), .config_in(config_chain[3554:3552]), .config_rst(config_rst)); 
mux6 mux_1185 (.in({n13143_0, n13142_0, n13135_0, n13134_0, n13121_1, n13120_0}), .out(n2690), .config_in(config_chain[3557:3555]), .config_rst(config_rst)); 
mux6 mux_1186 (.in({n10261_1, n10260_0, n10227_0, n10226_0, n10197_0/**/, n10196_0}), .out(n2691), .config_in(config_chain[3560:3558]), .config_rst(config_rst)); 
mux6 mux_1187 (.in({n12865_1, n12864_0, n12831_0/**/, n12830_0, n12801_0, n12800_0}), .out(n2692), .config_in(config_chain[3563:3561]), .config_rst(config_rst)); 
mux6 mux_1188 (.in({n10551_1, n10550_0, n10539_0, n10538_0, n10519_1, n10518_0}), .out(n2693), .config_in(config_chain[3566:3564]), .config_rst(config_rst)); 
mux6 mux_1189 (.in({n13163_1, n13162_0, n13155_1, n13154_0, n13123_1, n13122_0}), .out(n2694), .config_in(config_chain[3569:3567]), .config_rst(config_rst)); 
mux6 mux_1190 (.in({n10273_0, n10272_0/**/, n10263_2, n10262_0, n10229_0, n10228_0}), .out(n2695), .config_in(config_chain[3572:3570]), .config_rst(config_rst)); 
mux6 mux_1191 (.in({n12877_0, n12876_0, n12869_2, n12868_0, n12833_0, n12832_0}), .out(n2696), .config_in(config_chain[3575:3573]), .config_rst(config_rst)); 
mux6 mux_1192 (.in({n10521_1, n10520_0, n10487_0/**/, n10486_0, n10455_0, n10454_0}), .out(n2697), .config_in(config_chain[3578:3576]), .config_rst(config_rst)); 
mux6 mux_1193 (.in({n13125_1, n13124_0, n13091_0, n13090_0, n13069_0/**/, n13068_0}), .out(n2698), .config_in(config_chain[3581:3579]), .config_rst(config_rst)); 
mux6 mux_1194 (.in({n10295_1, n10294_0, n10281_0, n10280_0, n10267_2, n10266_0}), .out(n2699), .config_in(config_chain[3584:3582]), .config_rst(config_rst)); 
mux6 mux_1195 (.in({n12907_1/**/, n12906_0, n12899_1, n12898_0, n12871_2, n12870_0}), .out(n2700), .config_in(config_chain[3587:3585]), .config_rst(config_rst)); 
mux6 mux_1196 (.in({n10523_2, n10522_0, n10497_0, n10496_0, n10465_0, n10464_0}), .out(n2701), .config_in(config_chain[3590:3588]), .config_rst(config_rst)); 
mux6 mux_1197 (.in({n13137_0, n13136_0/**/, n13127_2, n13126_0, n13101_0, n13100_0}), .out(n2702), .config_in(config_chain[3593:3591]), .config_rst(config_rst)); 
mux6 mux_1198 (.in({n10303_1, n10302_0, n10257_1, n10256_0, n10203_0/**/, n10202_0}), .out(n2703), .config_in(config_chain[3596:3594]), .config_rst(config_rst)); 
mux6 mux_1199 (.in({n12861_1, n12860_0, n12839_0, n12838_0, n12807_0, n12806_0/**/}), .out(n2704), .config_in(config_chain[3599:3597]), .config_rst(config_rst)); 
mux6 mux_1200 (.in({n10553_1, n10552_0, n10541_0/**/, n10540_0, n10525_2, n10524_0}), .out(n2705), .config_in(config_chain[3602:3600]), .config_rst(config_rst)); 
mux6 mux_1201 (.in({n13157_1, n13156_0, n13145_0, n13144_0, n13119_0/**/, n13118_0}), .out(n2706), .config_in(config_chain[3605:3603]), .config_rst(config_rst)); 
mux6 mux_1202 (.in({n10259_1, n10258_0, n10237_0, n10236_0, n10205_0, n10204_0}), .out(n2707), .config_in(config_chain[3608:3606]), .config_rst(config_rst)); 
mux6 mux_1203 (.in({n12879_0, n12878_0/**/, n12863_1, n12862_0, n12841_0, n12840_0}), .out(n2708), .config_in(config_chain[3611:3609]), .config_rst(config_rst)); 
mux6 mux_1204 (.in({n10807_1, n10806_0, n10793_0, n10792_0, n10751_0, n10750_0}), .out(n2755), .config_in(config_chain[3614:3612]), .config_rst(config_rst)); 
mux6 mux_1205 (.in({n13171_1, n13170_0, n13157_0, n13156_0, n13145_0, n13144_0}), .out(n2756), .config_in(config_chain[3617:3615]), .config_rst(config_rst)); 
mux6 mux_1206 (.in({n10495_0, n10494_0, n10463_0, n10462_0, n10441_0, n10440_0}), .out(n2757), .config_in(config_chain[3620:3618]), .config_rst(config_rst)); 
mux6 mux_1207 (.in({n12881_0, n12880_0, n12873_0, n12872_0, n12841_0, n12840_1}), .out(n2758), .config_in(config_chain[3623:3621]), .config_rst(config_rst)); 
mux6 mux_1208 (.in({n10815_1, n10814_0, n10801_0, n10800_0, n10701_0, n10700_0}), .out(n2759), .config_in(config_chain[3626:3624]), .config_rst(config_rst)); 
mux6 mux_1209 (.in({n13187_1, n13186_0, n13179_1, n13178_0, n13045_0, n13044_1}), .out(n2760), .config_in(config_chain[3629:3627]), .config_rst(config_rst)); 
mux6 mux_1210 (.in({n10535_0, n10534_0, n10527_0, n10526_0, n10505_0, n10504_0}), .out(n2761), .config_in(config_chain[3632:3630]), .config_rst(config_rst)); 
mux6 mux_1211 (.in({n12913_1, n12912_0, n12901_0, n12900_0, n12889_0, n12888_0}), .out(n2762), .config_in(config_chain[3635:3633]), .config_rst(config_rst)); 
mux6 mux_1212 (.in({n10765_0, n10764_0, n10733_0, n10732_0, n10695_0, n10694_0}), .out(n2763), .config_in(config_chain[3638:3636]), .config_rst(config_rst)); 
mux6 mux_1213 (.in({n13131_0, n13130_0/**/, n13109_0, n13108_1, n13077_0, n13076_1}), .out(n2764), .config_in(config_chain[3641:3639]), .config_rst(config_rst)); 
mux6 mux_1214 (.in({n10555_1, n10554_0/**/, n10547_1, n10546_0, n10543_0, n10542_0}), .out(n2765), .config_in(config_chain[3644:3642]), .config_rst(config_rst)); 
mux6 mux_1215 (.in({n12921_1, n12920_0, n12909_0, n12908_0/**/, n12785_0, n12784_1}), .out(n2766), .config_in(config_chain[3647:3645]), .config_rst(config_rst)); 
mux6 mux_1216 (.in({n10787_0, n10786_0, n10759_0, n10758_0, n10727_0, n10726_0}), .out(n2767), .config_in(config_chain[3650:3648]), .config_rst(config_rst)); 
mux6 mux_1217 (.in({n13159_0, n13158_0/**/, n13151_0, n13150_0, n13147_0, n13146_0}), .out(n2768), .config_in(config_chain[3653:3651]), .config_rst(config_rst)); 
mux6 mux_1218 (.in({n10563_1, n10562_0, n10471_0, n10470_0, n10449_0, n10448_0}), .out(n2769), .config_in(config_chain[3656:3654]), .config_rst(config_rst)); 
mux6 mux_1219 (.in({n12875_0/**/, n12874_0, n12849_0, n12848_1, n12817_0, n12816_1}), .out(n2770), .config_in(config_chain[3659:3657]), .config_rst(config_rst)); 
mux6 mux_1220 (.in({n10817_1, n10816_0, n10809_1/**/, n10808_0, n10803_0, n10802_0}), .out(n2771), .config_in(config_chain[3662:3660]), .config_rst(config_rst)); 
mux6 mux_1221 (.in({n13181_1, n13180_0, n13167_0, n13166_0, n13053_0, n13052_1}), .out(n2772), .config_in(config_chain[3665:3663]), .config_rst(config_rst)); 
mux6 mux_1222 (.in({n10529_0, n10528_0, n10503_0/**/, n10502_0, n10481_0, n10480_0}), .out(n2773), .config_in(config_chain[3668:3666]), .config_rst(config_rst)); 
mux6 mux_1223 (.in({n12895_0, n12894_0/**/, n12891_0, n12890_0, n12883_0, n12882_0}), .out(n2774), .config_in(config_chain[3671:3669]), .config_rst(config_rst)); 
mux6 mux_1224 (.in({n10825_1/**/, n10824_0, n10741_0, n10740_0, n10709_0, n10708_0}), .out(n2775), .config_in(config_chain[3674:3672]), .config_rst(config_rst)); 
mux6 mux_1225 (.in({n13189_1/**/, n13188_0, n13133_0, n13132_0, n13085_0, n13084_1}), .out(n2776), .config_in(config_chain[3677:3675]), .config_rst(config_rst)); 
mux6 mux_1226 (.in({n10549_1, n10548_0, n10545_0/**/, n10544_0, n10537_0, n10536_0}), .out(n2777), .config_in(config_chain[3680:3678]), .config_rst(config_rst)); 
mux6 mux_1227 (.in({n12923_1, n12922_0, n12915_1, n12914_0, n12911_0, n12910_0/**/}), .out(n2778), .config_in(config_chain[3683:3681]), .config_rst(config_rst)); 
mux6 mux_1228 (.in({n10789_0, n10788_0, n10773_0, n10772_0, n10735_0, n10734_0}), .out(n2779), .config_in(config_chain[3686:3684]), .config_rst(config_rst)); 
mux6 mux_1229 (.in({n13153_0, n13152_0, n13149_0, n13148_0, n13141_0, n13140_0}), .out(n2780), .config_in(config_chain[3689:3687]), .config_rst(config_rst)); 
mux6 mux_1230 (.in({n10565_1, n10564_0/**/, n10479_0, n10478_0, n10447_0, n10446_0}), .out(n2781), .config_in(config_chain[3692:3690]), .config_rst(config_rst)); 
mux6 mux_1231 (.in({n12931_1, n12930_0, n12825_0, n12824_1/**/, n12793_0, n12792_1}), .out(n2782), .config_in(config_chain[3695:3693]), .config_rst(config_rst)); 
mux6 mux_1232 (.in({n10811_1, n10810_0, n10797_0, n10796_0, n10767_0, n10766_0}), .out(n2783), .config_in(config_chain[3698:3696]), .config_rst(config_rst)); 
mux6 mux_1233 (.in({n13175_1, n13174_0, n13169_0, n13168_0, n13161_0, n13160_0/**/}), .out(n2784), .config_in(config_chain[3701:3699]), .config_rst(config_rst)); 
mux6 mux_1234 (.in({n10511_0, n10510_0, n10489_0/**/, n10488_0, n10457_0, n10456_0}), .out(n2785), .config_in(config_chain[3704:3702]), .config_rst(config_rst)); 
mux6 mux_1235 (.in({n12897_0, n12896_0, n12885_0, n12884_0, n12857_0/**/, n12856_1}), .out(n2786), .config_in(config_chain[3707:3705]), .config_rst(config_rst)); 
mux6 mux_1236 (.in({n10819_1, n10818_0, n10775_0, n10774_0, n10717_0, n10716_0}), .out(n2787), .config_in(config_chain[3710:3708]), .config_rst(config_rst)); 
mux6 mux_1237 (.in({n13119_0, n13118_1, n13093_0, n13092_1, n13061_0, n13060_1}), .out(n2788), .config_in(config_chain[3713:3711]), .config_rst(config_rst)); 
mux6 mux_1238 (.in({n10551_1, n10550_0, n10539_0/**/, n10538_0, n10517_1, n10516_0}), .out(n2789), .config_in(config_chain[3716:3714]), .config_rst(config_rst)); 
mux6 mux_1239 (.in({n12917_1, n12916_0, n12905_0, n12904_0, n12863_1, n12862_1}), .out(n2790), .config_in(config_chain[3719:3717]), .config_rst(config_rst)); 
mux6 mux_1240 (.in({n10777_0, n10776_0, n10749_0, n10748_0, n10711_0/**/, n10710_0}), .out(n2791), .config_in(config_chain[3722:3720]), .config_rst(config_rst)); 
mux6 mux_1241 (.in({n13143_0, n13142_0, n13135_0/**/, n13134_0, n13121_0, n13120_1}), .out(n2792), .config_in(config_chain[3725:3723]), .config_rst(config_rst)); 
mux6 mux_1242 (.in({n10559_1, n10558_0, n10519_1/**/, n10518_0, n10455_0, n10454_0}), .out(n2793), .config_in(config_chain[3728:3726]), .config_rst(config_rst)); 
mux6 mux_1243 (.in({n12925_1, n12924_0, n12867_1, n12866_1, n12801_0, n12800_1/**/}), .out(n2794), .config_in(config_chain[3731:3729]), .config_rst(config_rst)); 
mux6 mux_1244 (.in({n10799_0, n10798_0, n10791_0, n10790_0, n10779_1, n10778_0}), .out(n2795), .config_in(config_chain[3734:3732]), .config_rst(config_rst)); 
mux6 mux_1245 (.in({n13177_1, n13176_0, n13163_0, n13162_0/**/, n13123_1, n13122_1}), .out(n2796), .config_in(config_chain[3737:3735]), .config_rst(config_rst)); 
mux6 mux_1246 (.in({n10523_2, n10522_0, n10487_0, n10486_0, n10465_0, n10464_0}), .out(n2797), .config_in(config_chain[3740:3738]), .config_rst(config_rst)); 
mux6 mux_1247 (.in({n12887_0/**/, n12886_0, n12879_0, n12878_0, n12869_1, n12868_1}), .out(n2798), .config_in(config_chain[3743:3741]), .config_rst(config_rst)); 
mux6 mux_1248 (.in({n10821_1, n10820_0, n10813_1, n10812_0, n10781_1, n10780_0}), .out(n2799), .config_in(config_chain[3746:3744]), .config_rst(config_rst)); 
mux6 mux_1249 (.in({n13185_1, n13184_0/**/, n13125_1, n13124_1, n13069_0, n13068_1}), .out(n2800), .config_in(config_chain[3749:3747]), .config_rst(config_rst)); 
mux6 mux_1250 (.in({n10533_0, n10532_0, n10525_2, n10524_0, n10497_0, n10496_0}), .out(n2801), .config_in(config_chain[3752:3750]), .config_rst(config_rst)); 
mux6 mux_1251 (.in({n12907_0, n12906_0, n12899_0, n12898_0/**/, n12871_1, n12870_1}), .out(n2802), .config_in(config_chain[3755:3753]), .config_rst(config_rst)); 
mux6 mux_1252 (.in({n10783_1, n10782_0, n10757_0, n10756_0, n10719_0/**/, n10718_0}), .out(n2803), .config_in(config_chain[3758:3756]), .config_rst(config_rst)); 
mux6 mux_1253 (.in({n13137_0, n13136_0, n13129_1, n13128_1, n13101_0, n13100_1}), .out(n2804), .config_in(config_chain[3761:3759]), .config_rst(config_rst)); 
mux6 mux_1254 (.in({n10561_1, n10560_0, n10553_1, n10552_0, n10515_0/**/, n10514_0}), .out(n2805), .config_in(config_chain[3764:3762]), .config_rst(config_rst)); 
mux6 mux_1255 (.in({n12927_1, n12926_0, n12861_0, n12860_1, n12809_0, n12808_1}), .out(n2806), .config_in(config_chain[3767:3765]), .config_rst(config_rst)); 
mux6 mux_1256 (.in({n11083_1, n11082_0, n10981_0, n10980_0, n10959_0, n10958_0}), .out(n2853), .config_in(config_chain[3770:3768]), .config_rst(config_rst)); 
mux6 mux_1257 (.in({n13205_1, n13204_0, n13151_0, n13150_0, n13137_0, n13136_1}), .out(n2854), .config_in(config_chain[3773:3771]), .config_rst(config_rst)); 
mux6 mux_1258 (.in({n10807_1, n10806_0, n10801_0, n10800_0, n10793_0, n10792_0}), .out(n2855), .config_in(config_chain[3776:3774]), .config_rst(config_rst)); 
mux6 mux_1259 (.in({n12941_1, n12940_0, n12933_1, n12932_0, n12927_0, n12926_0}), .out(n2856), .config_in(config_chain[3779:3777]), .config_rst(config_rst)); 
mux6 mux_1260 (.in({n11049_0, n11048_0, n11013_0, n11012_0, n10991_0, n10990_0}), .out(n2857), .config_in(config_chain[3782:3780]), .config_rst(config_rst)); 
mux6 mux_1261 (.in({n13171_0, n13170_0, n13167_0, n13166_0, n13159_0, n13158_0}), .out(n2858), .config_in(config_chain[3785:3783]), .config_rst(config_rst)); 
mux6 mux_1262 (.in({n10823_1, n10822_0, n10733_0, n10732_0, n10701_0, n10700_0}), .out(n2859), .config_in(config_chain[3788:3786]), .config_rst(config_rst)); 
mux6 mux_1263 (.in({n12949_1, n12948_0, n12893_0, n12892_0, n12881_0, n12880_1}), .out(n2860), .config_in(config_chain[3791:3789]), .config_rst(config_rst)); 
mux6 mux_1264 (.in({n11069_1/**/, n11068_0, n11065_0, n11064_0, n11057_0, n11056_0}), .out(n2861), .config_in(config_chain[3794:3792]), .config_rst(config_rst)); 
mux6 mux_1265 (.in({n13191_1, n13190_0, n13187_0, n13186_0, n13179_0, n13178_0/**/}), .out(n2862), .config_in(config_chain[3797:3795]), .config_rst(config_rst)); 
mux6 mux_1266 (.in({n10765_0, n10764_0, n10727_0, n10726_0, n10695_0, n10694_0}), .out(n2863), .config_in(config_chain[3800:3798]), .config_rst(config_rst)); 
mux6 mux_1267 (.in({n12913_0, n12912_0, n12901_0/**/, n12900_0, n12889_0, n12888_1}), .out(n2864), .config_in(config_chain[3803:3801]), .config_rst(config_rst)); 
mux6 mux_1268 (.in({n11085_1, n11084_0, n11077_1, n11076_0, n10957_0, n10956_0}), .out(n2865), .config_in(config_chain[3806:3804]), .config_rst(config_rst)); 
mux6 mux_1269 (.in({n13207_1, n13206_0, n13139_0, n13138_1, n13131_0, n13130_1}), .out(n2866), .config_in(config_chain[3809:3807]), .config_rst(config_rst)); 
mux6 mux_1270 (.in({n10809_1, n10808_0, n10795_0, n10794_0/**/, n10759_0, n10758_0}), .out(n2867), .config_in(config_chain[3812:3810]), .config_rst(config_rst)); 
mux6 mux_1271 (.in({n12935_1, n12934_0/**/, n12929_0, n12928_0, n12921_0, n12920_0}), .out(n2868), .config_in(config_chain[3815:3813]), .config_rst(config_rst)); 
mux6 mux_1272 (.in({n11021_0, n11020_0/**/, n10999_0, n10998_0, n10967_0, n10966_0}), .out(n2869), .config_in(config_chain[3818:3816]), .config_rst(config_rst)); 
mux6 mux_1273 (.in({n13173_0, n13172_0, n13161_0, n13160_0, n13147_0, n13146_1}), .out(n2870), .config_in(config_chain[3821:3819]), .config_rst(config_rst)); 
mux6 mux_1274 (.in({n10817_1, n10816_0, n10803_0, n10802_0, n10709_0, n10708_0/**/}), .out(n2871), .config_in(config_chain[3824:3822]), .config_rst(config_rst)); 
mux6 mux_1275 (.in({n12951_1, n12950_0, n12943_1/**/, n12942_0, n12875_0, n12874_1}), .out(n2872), .config_in(config_chain[3827:3825]), .config_rst(config_rst)); 
mux6 mux_1276 (.in({n11059_0, n11058_0, n11051_0, n11050_0, n11031_0, n11030_0}), .out(n2873), .config_in(config_chain[3830:3828]), .config_rst(config_rst)); 
mux6 mux_1277 (.in({n13193_1, n13192_0, n13181_0, n13180_0, n13169_0, n13168_0/**/}), .out(n2874), .config_in(config_chain[3833:3831]), .config_rst(config_rst)); 
mux6 mux_1278 (.in({n10773_0, n10772_0, n10741_0, n10740_0/**/, n10703_0, n10702_0}), .out(n2875), .config_in(config_chain[3836:3834]), .config_rst(config_rst)); 
mux6 mux_1279 (.in({n12903_0, n12902_0, n12895_0/**/, n12894_0, n12891_0, n12890_1}), .out(n2876), .config_in(config_chain[3839:3837]), .config_rst(config_rst)); 
mux6 mux_1280 (.in({n11079_1, n11078_0, n11067_0, n11066_0, n10965_0, n10964_0/**/}), .out(n2877), .config_in(config_chain[3842:3840]), .config_rst(config_rst)); 
mux6 mux_1281 (.in({n13209_1, n13208_0, n13201_1, n13200_0, n13133_0, n13132_1}), .out(n2878), .config_in(config_chain[3845:3843]), .config_rst(config_rst)); 
mux6 mux_1282 (.in({n10797_0, n10796_0, n10789_0, n10788_0, n10767_0, n10766_0}), .out(n2879), .config_in(config_chain[3848:3846]), .config_rst(config_rst)); 
mux6 mux_1283 (.in({n12923_0, n12922_0, n12915_0, n12914_0, n12911_0, n12910_0}), .out(n2880), .config_in(config_chain[3851:3849]), .config_rst(config_rst)); 
mux6 mux_1284 (.in({n11087_1, n11086_0, n10997_0, n10996_0/**/, n10975_0, n10974_0}), .out(n2881), .config_in(config_chain[3854:3852]), .config_rst(config_rst)); 
mux6 mux_1285 (.in({n13155_0, n13154_0, n13149_0, n13148_1, n13141_0, n13140_1/**/}), .out(n2882), .config_in(config_chain[3857:3855]), .config_rst(config_rst)); 
mux6 mux_1286 (.in({n10819_1, n10818_0, n10811_1, n10810_0, n10805_0, n10804_0}), .out(n2883), .config_in(config_chain[3860:3858]), .config_rst(config_rst)); 
mux6 mux_1287 (.in({n12945_1, n12944_0, n12931_0, n12930_0/**/, n12877_0, n12876_1}), .out(n2884), .config_in(config_chain[3863:3861]), .config_rst(config_rst)); 
mux6 mux_1288 (.in({n11053_0/**/, n11052_0, n11047_1, n11046_0, n11007_0, n11006_0}), .out(n2885), .config_in(config_chain[3866:3864]), .config_rst(config_rst)); 
mux6 mux_1289 (.in({n13183_0, n13182_0, n13175_0, n13174_0, n13129_1, n13128_1}), .out(n2886), .config_in(config_chain[3869:3867]), .config_rst(config_rst)); 
mux6 mux_1290 (.in({n10775_0, n10774_0, n10749_0, n10748_0, n10711_0, n10710_0}), .out(n2887), .config_in(config_chain[3872:3870]), .config_rst(config_rst)); 
mux6 mux_1291 (.in({n12897_0, n12896_0, n12885_0, n12884_1/**/, n12861_0, n12860_1}), .out(n2888), .config_in(config_chain[3875:3873]), .config_rst(config_rst)); 
mux6 mux_1292 (.in({n11073_1, n11072_0, n11061_0, n11060_0, n11037_0, n11036_0}), .out(n2889), .config_in(config_chain[3878:3876]), .config_rst(config_rst)); 
mux6 mux_1293 (.in({n13203_1, n13202_0, n13195_1, n13194_0, n13119_0, n13118_1}), .out(n2890), .config_in(config_chain[3881:3879]), .config_rst(config_rst)); 
mux6 mux_1294 (.in({n10791_0, n10790_0, n10777_0, n10776_0, n10743_0/**/, n10742_0}), .out(n2891), .config_in(config_chain[3884:3882]), .config_rst(config_rst)); 
mux6 mux_1295 (.in({n12917_0, n12916_0, n12905_0, n12904_0, n12865_1, n12864_1}), .out(n2892), .config_in(config_chain[3887:3885]), .config_rst(config_rst)); 
mux6 mux_1296 (.in({n11039_0, n11038_0, n11005_0/**/, n11004_0, n10973_0, n10972_0}), .out(n2893), .config_in(config_chain[3890:3888]), .config_rst(config_rst)); 
mux6 mux_1297 (.in({n13157_0, n13156_0/**/, n13143_0, n13142_1, n13121_0, n13120_1}), .out(n2894), .config_in(config_chain[3893:3891]), .config_rst(config_rst)); 
mux6 mux_1298 (.in({n10813_1, n10812_0, n10799_0, n10798_0, n10781_1, n10780_0}), .out(n2895), .config_in(config_chain[3896:3894]), .config_rst(config_rst)); 
mux6 mux_1299 (.in({n12947_1, n12946_0, n12939_1, n12938_0, n12867_1, n12866_1}), .out(n2896), .config_in(config_chain[3899:3897]), .config_rst(config_rst)); 
mux6 mux_1300 (.in({n11041_0, n11040_0, n11015_0, n11014_0, n10983_0, n10982_0}), .out(n2897), .config_in(config_chain[3902:3900]), .config_rst(config_rst)); 
mux6 mux_1301 (.in({n13177_0, n13176_0, n13165_0, n13164_0, n13123_0, n13122_1}), .out(n2898), .config_in(config_chain[3905:3903]), .config_rst(config_rst)); 
mux6 mux_1302 (.in({n10821_1, n10820_0, n10783_1, n10782_0, n10725_0, n10724_0}), .out(n2899), .config_in(config_chain[3908:3906]), .config_rst(config_rst)); 
mux6 mux_1303 (.in({n12887_0, n12886_1/**/, n12879_0, n12878_1, n12869_1, n12868_1}), .out(n2900), .config_in(config_chain[3911:3909]), .config_rst(config_rst)); 
mux6 mux_1304 (.in({n11075_1/**/, n11074_0, n11063_0, n11062_0, n11043_1, n11042_0}), .out(n2901), .config_in(config_chain[3914:3912]), .config_rst(config_rst)); 
mux6 mux_1305 (.in({n13197_1, n13196_0, n13185_0, n13184_0, n13127_1, n13126_1}), .out(n2902), .config_in(config_chain[3917:3915]), .config_rst(config_rst)); 
mux6 mux_1306 (.in({n10785_2, n10784_0, n10751_0, n10750_0, n10719_0, n10718_0}), .out(n2903), .config_in(config_chain[3920:3918]), .config_rst(config_rst)); 
mux6 mux_1307 (.in({n12919_0, n12918_0, n12907_0, n12906_0, n12871_1, n12870_1}), .out(n2904), .config_in(config_chain[3923:3921]), .config_rst(config_rst)); 
mux6 mux_1308 (.in({n11333_1, n11332_0, n11319_0, n11318_0, n11281_0, n11280_0}), .out(n2951), .config_in(config_chain[3926:3924]), .config_rst(config_rst)); 
mux6 mux_1309 (.in({n13211_1, n13210_0, n13197_0, n13196_0, n13185_0, n13184_0}), .out(n2952), .config_in(config_chain[3929:3927]), .config_rst(config_rst)); 
mux6 mux_1310 (.in({n11013_0, n11012_0, n10981_0, n10980_0, n10959_0, n10958_0}), .out(n2953), .config_in(config_chain[3932:3930]), .config_rst(config_rst)); 
mux6 mux_1311 (.in({n12921_0, n12920_0, n12913_0, n12912_0, n12907_0, n12906_1}), .out(n2954), .config_in(config_chain[3935:3933]), .config_rst(config_rst)); 
mux6 mux_1312 (.in({n11341_1, n11340_0/**/, n11327_0, n11326_0, n11223_0, n11222_0}), .out(n2955), .config_in(config_chain[3938:3936]), .config_rst(config_rst)); 
mux6 mux_1313 (.in({n13227_1, n13226_0, n13219_1, n13218_0, n13151_0, n13150_1/**/}), .out(n2956), .config_in(config_chain[3941:3939]), .config_rst(config_rst)); 
mux6 mux_1314 (.in({n11057_0, n11056_0/**/, n11049_0, n11048_0, n11023_0, n11022_0}), .out(n2957), .config_in(config_chain[3944:3942]), .config_rst(config_rst)); 
mux6 mux_1315 (.in({n12953_1, n12952_0, n12941_0, n12940_0, n12929_0, n12928_0}), .out(n2958), .config_in(config_chain[3947:3945]), .config_rst(config_rst)); 
mux6 mux_1316 (.in({n11287_0, n11286_0, n11255_0, n11254_0, n11225_0, n11224_0}), .out(n2959), .config_in(config_chain[3950:3948]), .config_rst(config_rst)); 
mux6 mux_1317 (.in({n13171_0, n13170_0, n13167_0, n13166_1, n13159_0, n13158_1}), .out(n2960), .config_in(config_chain[3953:3951]), .config_rst(config_rst)); 
mux6 mux_1318 (.in({n11077_1, n11076_0, n11069_1, n11068_0, n11065_0, n11064_0}), .out(n2961), .config_in(config_chain[3956:3954]), .config_rst(config_rst)); 
mux6 mux_1319 (.in({n12961_1, n12960_0, n12949_0, n12948_0, n12893_0, n12892_1}), .out(n2962), .config_in(config_chain[3959:3957]), .config_rst(config_rst)); 
mux6 mux_1320 (.in({n11313_0, n11312_0, n11289_0, n11288_0, n11257_0, n11256_0}), .out(n2963), .config_in(config_chain[3962:3960]), .config_rst(config_rst)); 
mux6 mux_1321 (.in({n13199_0, n13198_0/**/, n13191_0, n13190_0, n13187_0, n13186_0}), .out(n2964), .config_in(config_chain[3965:3963]), .config_rst(config_rst)); 
mux6 mux_1322 (.in({n11085_1, n11084_0, n10989_0, n10988_0/**/, n10967_0, n10966_0}), .out(n2965), .config_in(config_chain[3968:3966]), .config_rst(config_rst)); 
mux6 mux_1323 (.in({n12915_0, n12914_0/**/, n12909_0, n12908_1, n12901_0, n12900_1}), .out(n2966), .config_in(config_chain[3971:3969]), .config_rst(config_rst)); 
mux6 mux_1324 (.in({n11343_1, n11342_0, n11335_1, n11334_0/**/, n11329_0, n11328_0}), .out(n2967), .config_in(config_chain[3974:3972]), .config_rst(config_rst)); 
mux6 mux_1325 (.in({n13221_1, n13220_0, n13207_0, n13206_0, n13153_0, n13152_1}), .out(n2968), .config_in(config_chain[3977:3975]), .config_rst(config_rst)); 
mux6 mux_1326 (.in({n11051_0, n11050_0, n11021_0, n11020_0, n10999_0, n10998_0/**/}), .out(n2969), .config_in(config_chain[3980:3978]), .config_rst(config_rst)); 
mux6 mux_1327 (.in({n12935_0, n12934_0, n12931_0, n12930_0, n12923_0, n12922_0}), .out(n2970), .config_in(config_chain[3983:3981]), .config_rst(config_rst)); 
mux6 mux_1328 (.in({n11351_1, n11350_0, n11263_0, n11262_0, n11231_0, n11230_0}), .out(n2971), .config_in(config_chain[3986:3984]), .config_rst(config_rst)); 
mux6 mux_1329 (.in({n13229_1, n13228_0, n13173_0, n13172_0, n13161_0/**/, n13160_1}), .out(n2972), .config_in(config_chain[3989:3987]), .config_rst(config_rst)); 
mux6 mux_1330 (.in({n11071_1, n11070_0, n11067_0/**/, n11066_0, n11059_0, n11058_0}), .out(n2973), .config_in(config_chain[3992:3990]), .config_rst(config_rst)); 
mux6 mux_1331 (.in({n12963_1, n12962_0, n12955_1, n12954_0, n12951_0/**/, n12950_0}), .out(n2974), .config_in(config_chain[3995:3993]), .config_rst(config_rst)); 
mux6 mux_1332 (.in({n11315_0, n11314_0/**/, n11295_0, n11294_0, n11265_0, n11264_0}), .out(n2975), .config_in(config_chain[3998:3996]), .config_rst(config_rst)); 
mux6 mux_1333 (.in({n13193_0, n13192_0, n13189_0, n13188_0, n13181_0, n13180_0}), .out(n2976), .config_in(config_chain[4001:3999]), .config_rst(config_rst)); 
mux6 mux_1334 (.in({n11087_1, n11086_0, n10997_0, n10996_0, n10965_0, n10964_0}), .out(n2977), .config_in(config_chain[4004:4002]), .config_rst(config_rst)); 
mux6 mux_1335 (.in({n12971_1, n12970_0, n12903_0, n12902_1, n12895_0, n12894_1}), .out(n2978), .config_in(config_chain[4007:4005]), .config_rst(config_rst)); 
mux6 mux_1336 (.in({n11337_1, n11336_0, n11323_0, n11322_0, n11297_0, n11296_0}), .out(n2979), .config_in(config_chain[4010:4008]), .config_rst(config_rst)); 
mux6 mux_1337 (.in({n13215_1, n13214_0, n13209_0, n13208_0, n13201_0, n13200_0}), .out(n2980), .config_in(config_chain[4013:4011]), .config_rst(config_rst)); 
mux6 mux_1338 (.in({n11029_0, n11028_0, n11007_0, n11006_0, n10975_0/**/, n10974_0}), .out(n2981), .config_in(config_chain[4016:4014]), .config_rst(config_rst)); 
mux6 mux_1339 (.in({n12937_0, n12936_0/**/, n12925_0, n12924_0, n12911_0, n12910_1}), .out(n2982), .config_in(config_chain[4019:4017]), .config_rst(config_rst)); 
mux6 mux_1340 (.in({n11345_1/**/, n11344_0, n11309_1, n11308_0, n11239_0, n11238_0}), .out(n2983), .config_in(config_chain[4022:4020]), .config_rst(config_rst)); 
mux6 mux_1341 (.in({n13163_0, n13162_1, n13155_0, n13154_1, n13127_1, n13126_1}), .out(n2984), .config_in(config_chain[4025:4023]), .config_rst(config_rst)); 
mux6 mux_1342 (.in({n11073_1, n11072_0, n11061_0, n11060_0, n11047_1/**/, n11046_0}), .out(n2985), .config_in(config_chain[4028:4026]), .config_rst(config_rst)); 
mux6 mux_1343 (.in({n12957_1, n12956_0, n12945_0, n12944_0/**/, n12871_1, n12870_1}), .out(n2986), .config_in(config_chain[4031:4029]), .config_rst(config_rst)); 
mux6 mux_1344 (.in({n11311_1, n11310_0, n11271_0/**/, n11270_0, n11241_0, n11240_0}), .out(n2987), .config_in(config_chain[4034:4032]), .config_rst(config_rst)); 
mux6 mux_1345 (.in({n13183_0, n13182_0, n13175_0, n13174_0, n13129_1, n13128_1}), .out(n2988), .config_in(config_chain[4037:4035]), .config_rst(config_rst)); 
mux6 mux_1346 (.in({n11081_1, n11080_0, n11037_0, n11036_0, n10973_0, n10972_0/**/}), .out(n2989), .config_in(config_chain[4040:4038]), .config_rst(config_rst)); 
mux6 mux_1347 (.in({n12965_1, n12964_0, n12897_0, n12896_1, n12863_0, n12862_1}), .out(n2990), .config_in(config_chain[4043:4041]), .config_rst(config_rst)); 
mux6 mux_1348 (.in({n11353_2, n11352_0, n11325_0, n11324_0, n11317_0, n11316_0}), .out(n2991), .config_in(config_chain[4046:4044]), .config_rst(config_rst)); 
mux6 mux_1349 (.in({n13231_1, n13230_0, n13217_1, n13216_0, n13203_0, n13202_0}), .out(n2992), .config_in(config_chain[4049:4047]), .config_rst(config_rst)); 
mux6 mux_1350 (.in({n11041_0, n11040_0, n11005_0, n11004_0, n10983_0/**/, n10982_0}), .out(n2993), .config_in(config_chain[4052:4050]), .config_rst(config_rst)); 
mux6 mux_1351 (.in({n12927_0, n12926_0, n12919_0, n12918_0, n12865_0, n12864_1}), .out(n2994), .config_in(config_chain[4055:4053]), .config_rst(config_rst)); 
mux6 mux_1352 (.in({n11347_1/**/, n11346_0, n11339_1, n11338_0, n11303_0, n11302_0}), .out(n2995), .config_in(config_chain[4058:4056]), .config_rst(config_rst)); 
mux6 mux_1353 (.in({n13225_1, n13224_0, n13157_0, n13156_1, n13121_0, n13120_1}), .out(n2996), .config_in(config_chain[4061:4059]), .config_rst(config_rst)); 
mux6 mux_1354 (.in({n11055_0, n11054_0, n11043_1, n11042_0, n11015_0, n11014_0}), .out(n2997), .config_in(config_chain[4064:4062]), .config_rst(config_rst)); 
mux6 mux_1355 (.in({n12947_0, n12946_0, n12939_0, n12938_0, n12867_1, n12866_1}), .out(n2998), .config_in(config_chain[4067:4065]), .config_rst(config_rst)); 
mux6 mux_1356 (.in({n11305_0, n11304_0, n11279_0, n11278_0, n11249_0, n11248_0}), .out(n2999), .config_in(config_chain[4070:4068]), .config_rst(config_rst)); 
mux6 mux_1357 (.in({n13177_0, n13176_0, n13165_0, n13164_1/**/, n13125_0, n13124_1}), .out(n3000), .config_in(config_chain[4073:4071]), .config_rst(config_rst)); 
mux6 mux_1358 (.in({n11083_1, n11082_0, n11075_1, n11074_0, n11045_1, n11044_0}), .out(n3001), .config_in(config_chain[4076:4074]), .config_rst(config_rst)); 
mux6 mux_1359 (.in({n12967_1, n12966_0, n12899_0, n12898_1, n12869_1, n12868_1}), .out(n3002), .config_in(config_chain[4079:4077]), .config_rst(config_rst)); 
mux6 mux_1360 (.in({n11613_1, n11612_0, n11513_0, n11512_0, n11491_0, n11490_0}), .out(n3049), .config_in(config_chain[4082:4080]), .config_rst(config_rst)); 
mux6 mux_1361 (.in({n13247_0, n13246_0, n13191_0, n13190_0, n13177_0, n13176_1}), .out(n3050), .config_in(config_chain[4085:4083]), .config_rst(config_rst)); 
mux6 mux_1362 (.in({n11333_1, n11332_0, n11327_0, n11326_0, n11319_0, n11318_0}), .out(n3051), .config_in(config_chain[4088:4086]), .config_rst(config_rst)); 
mux6 mux_1363 (.in({n12981_0, n12980_0, n12973_0, n12972_0, n12967_0, n12966_0}), .out(n3052), .config_in(config_chain[4091:4089]), .config_rst(config_rst)); 
mux6 mux_1364 (.in({n11577_0, n11576_0, n11545_0, n11544_0, n11523_0, n11522_0}), .out(n3053), .config_in(config_chain[4094:4092]), .config_rst(config_rst)); 
mux6 mux_1365 (.in({n13211_0, n13210_0, n13207_0, n13206_0, n13199_0, n13198_0}), .out(n3054), .config_in(config_chain[4097:4095]), .config_rst(config_rst)); 
mux6 mux_1366 (.in({n11349_1, n11348_0/**/, n11255_0, n11254_0, n11223_0, n11222_0}), .out(n3055), .config_in(config_chain[4100:4098]), .config_rst(config_rst)); 
mux6 mux_1367 (.in({n12989_0, n12988_0, n12933_0, n12932_0, n12921_0, n12920_1/**/}), .out(n3056), .config_in(config_chain[4103:4101]), .config_rst(config_rst)); 
mux6 mux_1368 (.in({n11599_1, n11598_0, n11593_0, n11592_0, n11585_0, n11584_0}), .out(n3057), .config_in(config_chain[4106:4104]), .config_rst(config_rst)); 
mux6 mux_1369 (.in({n13233_0, n13232_0, n13227_0, n13226_0/**/, n13219_0, n13218_0}), .out(n3058), .config_in(config_chain[4109:4107]), .config_rst(config_rst)); 
mux6 mux_1370 (.in({n11287_0, n11286_0, n11257_0, n11256_0, n11225_0, n11224_0}), .out(n3059), .config_in(config_chain[4112:4110]), .config_rst(config_rst)); 
mux6 mux_1371 (.in({n12953_0, n12952_0, n12941_0, n12940_0, n12929_0, n12928_1/**/}), .out(n3060), .config_in(config_chain[4115:4113]), .config_rst(config_rst)); 
mux6 mux_1372 (.in({n11615_1, n11614_0, n11607_1, n11606_0, n11489_0, n11488_0}), .out(n3061), .config_in(config_chain[4118:4116]), .config_rst(config_rst)); 
mux6 mux_1373 (.in({n13249_0, n13248_0, n13179_0/**/, n13178_1, n13171_0, n13170_1}), .out(n3062), .config_in(config_chain[4121:4119]), .config_rst(config_rst)); 
mux6 mux_1374 (.in({n11335_1, n11334_0, n11321_0, n11320_0, n11289_0, n11288_0}), .out(n3063), .config_in(config_chain[4124:4122]), .config_rst(config_rst)); 
mux6 mux_1375 (.in({n12975_0, n12974_0, n12969_0, n12968_0, n12961_0, n12960_0}), .out(n3064), .config_in(config_chain[4127:4125]), .config_rst(config_rst)); 
mux6 mux_1376 (.in({n11553_0, n11552_0, n11531_0, n11530_0/**/, n11499_0, n11498_0}), .out(n3065), .config_in(config_chain[4130:4128]), .config_rst(config_rst)); 
mux6 mux_1377 (.in({n13213_0, n13212_0, n13201_0, n13200_0, n13187_0, n13186_1}), .out(n3066), .config_in(config_chain[4133:4131]), .config_rst(config_rst)); 
mux6 mux_1378 (.in({n11343_1, n11342_0, n11329_0, n11328_0, n11231_0/**/, n11230_0}), .out(n3067), .config_in(config_chain[4136:4134]), .config_rst(config_rst)); 
mux6 mux_1379 (.in({n12991_0, n12990_0, n12983_0, n12982_0/**/, n12915_0, n12914_1}), .out(n3068), .config_in(config_chain[4139:4137]), .config_rst(config_rst)); 
mux6 mux_1380 (.in({n11587_0, n11586_0, n11579_0, n11578_0, n11563_0, n11562_0}), .out(n3069), .config_in(config_chain[4142:4140]), .config_rst(config_rst)); 
mux6 mux_1381 (.in({n13235_0, n13234_0, n13221_0, n13220_0, n13209_0, n13208_0}), .out(n3070), .config_in(config_chain[4145:4143]), .config_rst(config_rst)); 
mux6 mux_1382 (.in({n11295_0, n11294_0, n11263_0, n11262_0, n11233_0, n11232_0}), .out(n3071), .config_in(config_chain[4148:4146]), .config_rst(config_rst)); 
mux6 mux_1383 (.in({n12943_0/**/, n12942_0, n12935_0, n12934_0, n12931_0, n12930_1}), .out(n3072), .config_in(config_chain[4151:4149]), .config_rst(config_rst)); 
mux6 mux_1384 (.in({n11609_1, n11608_0, n11595_0, n11594_0, n11497_0, n11496_0}), .out(n3073), .config_in(config_chain[4154:4152]), .config_rst(config_rst)); 
mux6 mux_1385 (.in({n13251_0, n13250_0/**/, n13243_0, n13242_0, n13173_0, n13172_1}), .out(n3074), .config_in(config_chain[4157:4155]), .config_rst(config_rst)); 
mux6 mux_1386 (.in({n11323_0, n11322_0, n11315_0, n11314_0, n11297_0, n11296_0}), .out(n3075), .config_in(config_chain[4160:4158]), .config_rst(config_rst)); 
mux6 mux_1387 (.in({n12963_0, n12962_0, n12955_0/**/, n12954_0, n12951_0, n12950_0}), .out(n3076), .config_in(config_chain[4163:4161]), .config_rst(config_rst)); 
mux6 mux_1388 (.in({n11617_1/**/, n11616_0, n11529_0, n11528_0, n11507_0, n11506_0}), .out(n3077), .config_in(config_chain[4166:4164]), .config_rst(config_rst)); 
mux6 mux_1389 (.in({n13195_0/**/, n13194_0, n13189_0, n13188_1, n13181_0, n13180_1}), .out(n3078), .config_in(config_chain[4169:4167]), .config_rst(config_rst)); 
mux6 mux_1390 (.in({n11345_1, n11344_0, n11337_1, n11336_0, n11331_0, n11330_0}), .out(n3079), .config_in(config_chain[4172:4170]), .config_rst(config_rst)); 
mux6 mux_1391 (.in({n12985_0, n12984_0, n12971_0, n12970_0/**/, n12917_0, n12916_1}), .out(n3080), .config_in(config_chain[4175:4173]), .config_rst(config_rst)); 
mux6 mux_1392 (.in({n11581_0, n11580_0, n11571_0, n11570_0, n11539_0, n11538_0}), .out(n3081), .config_in(config_chain[4178:4176]), .config_rst(config_rst)); 
mux6 mux_1393 (.in({n13223_0, n13222_0, n13215_0/**/, n13214_0, n13125_0, n13124_2}), .out(n3082), .config_in(config_chain[4181:4179]), .config_rst(config_rst)); 
mux6 mux_1394 (.in({n11309_1, n11308_0, n11271_0, n11270_0, n11241_0, n11240_0}), .out(n3083), .config_in(config_chain[4184:4182]), .config_rst(config_rst)); 
mux6 mux_1395 (.in({n12937_0/**/, n12936_0, n12925_0, n12924_1, n12869_0, n12868_2}), .out(n3084), .config_in(config_chain[4187:4185]), .config_rst(config_rst)); 
mux6 mux_1396 (.in({n11603_1, n11602_0, n11589_0, n11588_0/**/, n11573_0, n11572_0}), .out(n3085), .config_in(config_chain[4190:4188]), .config_rst(config_rst)); 
mux6 mux_1397 (.in({n13245_0/**/, n13244_0, n13237_0, n13236_0, n13127_0, n13126_2}), .out(n3086), .config_in(config_chain[4193:4191]), .config_rst(config_rst)); 
mux6 mux_1398 (.in({n11317_0, n11316_0, n11311_1, n11310_0, n11273_0, n11272_0}), .out(n3087), .config_in(config_chain[4196:4194]), .config_rst(config_rst)); 
mux6 mux_1399 (.in({n12993_0, n12992_0, n12957_0, n12956_0, n12945_0, n12944_0}), .out(n3088), .config_in(config_chain[4199:4197]), .config_rst(config_rst)); 
mux6 mux_1400 (.in({n11575_1, n11574_0, n11537_0, n11536_0, n11505_0/**/, n11504_0}), .out(n3089), .config_in(config_chain[4202:4200]), .config_rst(config_rst)); 
mux6 mux_1401 (.in({n13197_0, n13196_0, n13183_0, n13182_1, n13129_0, n13128_2}), .out(n3090), .config_in(config_chain[4205:4203]), .config_rst(config_rst)); 
mux6 mux_1402 (.in({n11339_1/**/, n11338_0, n11325_0, n11324_0, n11303_0, n11302_0}), .out(n3091), .config_in(config_chain[4208:4206]), .config_rst(config_rst)); 
mux6 mux_1403 (.in({n12987_0, n12986_0/**/, n12979_0, n12978_0, n12863_0, n12862_2}), .out(n3092), .config_in(config_chain[4211:4209]), .config_rst(config_rst)); 
mux6 mux_1404 (.in({n11597_2, n11596_0, n11547_0, n11546_0, n11515_0, n11514_0}), .out(n3093), .config_in(config_chain[4214:4212]), .config_rst(config_rst)); 
mux6 mux_1405 (.in({n13231_0, n13230_0, n13217_0, n13216_0/**/, n13205_0, n13204_0}), .out(n3094), .config_in(config_chain[4217:4215]), .config_rst(config_rst)); 
mux6 mux_1406 (.in({n11347_1, n11346_0, n11305_0, n11304_0, n11247_0, n11246_0/**/}), .out(n3095), .config_in(config_chain[4220:4218]), .config_rst(config_rst)); 
mux6 mux_1407 (.in({n12927_0, n12926_1/**/, n12919_0, n12918_1, n12865_0, n12864_2}), .out(n3096), .config_in(config_chain[4223:4221]), .config_rst(config_rst)); 
mux6 mux_1408 (.in({n11619_2, n11618_0, n11605_1, n11604_0, n11591_0, n11590_0/**/}), .out(n3097), .config_in(config_chain[4226:4224]), .config_rst(config_rst)); 
mux6 mux_1409 (.in({n13239_0, n13238_0, n13225_0, n13224_0, n13123_0, n13122_2}), .out(n3098), .config_in(config_chain[4229:4227]), .config_rst(config_rst)); 
mux6 mux_1410 (.in({n11307_0, n11306_0, n11281_0, n11280_0, n11249_0, n11248_0}), .out(n3099), .config_in(config_chain[4232:4230]), .config_rst(config_rst)); 
mux6 mux_1411 (.in({n12959_0, n12958_0/**/, n12947_0, n12946_0, n12867_0, n12866_2}), .out(n3100), .config_in(config_chain[4235:4233]), .config_rst(config_rst)); 
mux6 mux_1412 (.in({n11863_1, n11862_0, n11847_0, n11846_0, n11805_0, n11804_0}), .out(n3147), .config_in(config_chain[4238:4236]), .config_rst(config_rst)); 
mux6 mux_1413 (.in({n13255_0, n13254_0, n13239_0, n13238_0, n13225_0, n13224_0}), .out(n3148), .config_in(config_chain[4241:4239]), .config_rst(config_rst)); 
mux6 mux_1414 (.in({n11545_0, n11544_0, n11513_0, n11512_0, n11491_0, n11490_0}), .out(n3149), .config_in(config_chain[4244:4242]), .config_rst(config_rst)); 
mux6 mux_1415 (.in({n12961_0, n12960_0, n12953_0, n12952_0, n12947_0, n12946_1}), .out(n3150), .config_in(config_chain[4247:4245]), .config_rst(config_rst)); 
mux6 mux_1416 (.in({n11871_1, n11870_0, n11855_0, n11854_0, n11755_0, n11754_0}), .out(n3151), .config_in(config_chain[4250:4248]), .config_rst(config_rst)); 
mux6 mux_1417 (.in({n13271_0, n13270_0, n13263_0, n13262_0, n13191_0, n13190_1}), .out(n3152), .config_in(config_chain[4253:4251]), .config_rst(config_rst)); 
mux6 mux_1418 (.in({n11585_0, n11584_0, n11577_0, n11576_0, n11555_0, n11554_0}), .out(n3153), .config_in(config_chain[4256:4254]), .config_rst(config_rst)); 
mux6 mux_1419 (.in({n12995_0, n12994_0, n12981_0, n12980_0, n12969_0, n12968_0}), .out(n3154), .config_in(config_chain[4259:4257]), .config_rst(config_rst)); 
mux6 mux_1420 (.in({n11819_0, n11818_0, n11787_0, n11786_0, n11749_0, n11748_0}), .out(n3155), .config_in(config_chain[4262:4260]), .config_rst(config_rst)); 
mux6 mux_1421 (.in({n13211_0, n13210_0, n13207_0, n13206_1, n13199_0, n13198_1}), .out(n3156), .config_in(config_chain[4265:4263]), .config_rst(config_rst)); 
mux6 mux_1422 (.in({n11607_1, n11606_0, n11599_1, n11598_0, n11593_0, n11592_0}), .out(n3157), .config_in(config_chain[4268:4266]), .config_rst(config_rst)); 
mux6 mux_1423 (.in({n13003_0, n13002_0, n12989_0, n12988_0/**/, n12933_0, n12932_1}), .out(n3158), .config_in(config_chain[4271:4269]), .config_rst(config_rst)); 
mux6 mux_1424 (.in({n11841_0, n11840_0, n11813_0, n11812_0, n11781_0, n11780_0}), .out(n3159), .config_in(config_chain[4274:4272]), .config_rst(config_rst)); 
mux6 mux_1425 (.in({n13241_0, n13240_0, n13233_0, n13232_0/**/, n13227_0, n13226_0}), .out(n3160), .config_in(config_chain[4277:4275]), .config_rst(config_rst)); 
mux6 mux_1426 (.in({n11615_1, n11614_0/**/, n11521_0, n11520_0, n11499_0, n11498_0}), .out(n3161), .config_in(config_chain[4280:4278]), .config_rst(config_rst)); 
mux6 mux_1427 (.in({n12955_0, n12954_0/**/, n12949_0, n12948_1, n12941_0, n12940_1}), .out(n3162), .config_in(config_chain[4283:4281]), .config_rst(config_rst)); 
mux6 mux_1428 (.in({n11873_1, n11872_0, n11865_1, n11864_0, n11857_0/**/, n11856_0}), .out(n3163), .config_in(config_chain[4286:4284]), .config_rst(config_rst)); 
mux6 mux_1429 (.in({n13265_0/**/, n13264_0, n13249_0, n13248_0, n13193_0, n13192_1}), .out(n3164), .config_in(config_chain[4289:4287]), .config_rst(config_rst)); 
mux6 mux_1430 (.in({n11579_0, n11578_0, n11553_0, n11552_0, n11531_0, n11530_0/**/}), .out(n3165), .config_in(config_chain[4292:4290]), .config_rst(config_rst)); 
mux6 mux_1431 (.in({n12975_0, n12974_0, n12971_0, n12970_0, n12963_0, n12962_0}), .out(n3166), .config_in(config_chain[4295:4293]), .config_rst(config_rst)); 
mux6 mux_1432 (.in({n11881_1, n11880_0, n11795_0, n11794_0, n11763_0, n11762_0}), .out(n3167), .config_in(config_chain[4298:4296]), .config_rst(config_rst)); 
mux6 mux_1433 (.in({n13273_0, n13272_0, n13213_0, n13212_0, n13201_0, n13200_1/**/}), .out(n3168), .config_in(config_chain[4301:4299]), .config_rst(config_rst)); 
mux6 mux_1434 (.in({n11601_1, n11600_0/**/, n11595_0, n11594_0, n11587_0, n11586_0}), .out(n3169), .config_in(config_chain[4304:4302]), .config_rst(config_rst)); 
mux6 mux_1435 (.in({n13005_0, n13004_0/**/, n12997_0, n12996_0, n12991_0, n12990_0}), .out(n3170), .config_in(config_chain[4307:4305]), .config_rst(config_rst)); 
mux6 mux_1436 (.in({n11843_0, n11842_0, n11827_0/**/, n11826_0, n11789_0, n11788_0}), .out(n3171), .config_in(config_chain[4310:4308]), .config_rst(config_rst)); 
mux6 mux_1437 (.in({n13235_0, n13234_0, n13229_0, n13228_0, n13221_0, n13220_0}), .out(n3172), .config_in(config_chain[4313:4311]), .config_rst(config_rst)); 
mux6 mux_1438 (.in({n11617_1, n11616_0, n11529_0, n11528_0, n11497_0/**/, n11496_0}), .out(n3173), .config_in(config_chain[4316:4314]), .config_rst(config_rst)); 
mux6 mux_1439 (.in({n13013_0, n13012_0/**/, n12943_0, n12942_1, n12935_0, n12934_1}), .out(n3174), .config_in(config_chain[4319:4317]), .config_rst(config_rst)); 
mux6 mux_1440 (.in({n11867_1, n11866_0, n11851_0, n11850_0, n11821_0, n11820_0}), .out(n3175), .config_in(config_chain[4322:4320]), .config_rst(config_rst)); 
mux6 mux_1441 (.in({n13259_0, n13258_0, n13251_0, n13250_0, n13243_0, n13242_0}), .out(n3176), .config_in(config_chain[4325:4323]), .config_rst(config_rst)); 
mux6 mux_1442 (.in({n11561_0, n11560_0, n11539_0/**/, n11538_0, n11507_0, n11506_0}), .out(n3177), .config_in(config_chain[4328:4326]), .config_rst(config_rst)); 
mux6 mux_1443 (.in({n12977_0, n12976_0, n12965_0, n12964_0/**/, n12951_0, n12950_1}), .out(n3178), .config_in(config_chain[4331:4329]), .config_rst(config_rst)); 
mux6 mux_1444 (.in({n11883_2, n11882_0, n11875_1, n11874_0, n11771_0/**/, n11770_0}), .out(n3179), .config_in(config_chain[4334:4332]), .config_rst(config_rst)); 
mux6 mux_1445 (.in({n13275_0, n13274_0, n13203_0, n13202_1, n13195_0, n13194_1}), .out(n3180), .config_in(config_chain[4337:4335]), .config_rst(config_rst)); 
mux6 mux_1446 (.in({n11603_1, n11602_0, n11589_0/**/, n11588_0, n11571_0, n11570_0}), .out(n3181), .config_in(config_chain[4340:4338]), .config_rst(config_rst)); 
mux6 mux_1447 (.in({n12999_0, n12998_0, n12985_0, n12984_0, n12867_0, n12866_2}), .out(n3182), .config_in(config_chain[4343:4341]), .config_rst(config_rst)); 
mux6 mux_1448 (.in({n11835_0, n11834_0, n11803_0, n11802_0, n11765_0/**/, n11764_0}), .out(n3183), .config_in(config_chain[4346:4344]), .config_rst(config_rst)); 
mux6 mux_1449 (.in({n13223_0, n13222_0/**/, n13215_0, n13214_0, n13125_0, n13124_2}), .out(n3184), .config_in(config_chain[4349:4347]), .config_rst(config_rst)); 
mux6 mux_1450 (.in({n11611_1, n11610_0, n11573_0, n11572_0, n11505_0, n11504_0}), .out(n3185), .config_in(config_chain[4352:4350]), .config_rst(config_rst)); 
mux6 mux_1451 (.in({n13007_0, n13006_0, n12937_0, n12936_1, n12871_0, n12870_2}), .out(n3186), .config_in(config_chain[4355:4353]), .config_rst(config_rst)); 
mux6 mux_1452 (.in({n11853_0, n11852_0, n11845_0, n11844_0, n11837_0, n11836_0}), .out(n3187), .config_in(config_chain[4358:4356]), .config_rst(config_rst)); 
mux6 mux_1453 (.in({n13261_0, n13260_0, n13245_0, n13244_0, n13127_0, n13126_2}), .out(n3188), .config_in(config_chain[4361:4359]), .config_rst(config_rst)); 
mux6 mux_1454 (.in({n11597_2, n11596_0, n11537_0, n11536_0, n11515_0, n11514_0}), .out(n3189), .config_in(config_chain[4364:4362]), .config_rst(config_rst)); 
mux6 mux_1455 (.in({n12993_0, n12992_0, n12967_0, n12966_0/**/, n12959_0, n12958_0}), .out(n3190), .config_in(config_chain[4367:4365]), .config_rst(config_rst)); 
mux6 mux_1456 (.in({n11877_1, n11876_0, n11869_1, n11868_0, n11839_0/**/, n11838_0}), .out(n3191), .config_in(config_chain[4370:4368]), .config_rst(config_rst)); 
mux6 mux_1457 (.in({n13269_0/**/, n13268_0, n13197_0, n13196_1, n13129_0, n13128_2}), .out(n3192), .config_in(config_chain[4373:4371]), .config_rst(config_rst)); 
mux6 mux_1458 (.in({n11619_2, n11618_0, n11583_0, n11582_0, n11547_0, n11546_0}), .out(n3193), .config_in(config_chain[4376:4374]), .config_rst(config_rst)); 
mux6 mux_1459 (.in({n13015_0, n13014_0, n12987_0, n12986_0, n12979_0, n12978_0}), .out(n3194), .config_in(config_chain[4379:4377]), .config_rst(config_rst)); 
mux6 mux_1460 (.in({n11829_2, n11828_0, n11811_0/**/, n11810_0, n11773_0, n11772_0}), .out(n3195), .config_in(config_chain[4382:4380]), .config_rst(config_rst)); 
mux6 mux_1461 (.in({n13253_0, n13252_0, n13217_0, n13216_0, n13205_0/**/, n13204_1}), .out(n3196), .config_in(config_chain[4385:4383]), .config_rst(config_rst)); 
mux6 mux_1462 (.in({n11613_1, n11612_0, n11605_1, n11604_0, n11569_0, n11568_0}), .out(n3197), .config_in(config_chain[4388:4386]), .config_rst(config_rst)); 
mux6 mux_1463 (.in({n13009_0, n13008_0, n12939_0, n12938_1/**/, n12865_0, n12864_2}), .out(n3198), .config_in(config_chain[4391:4389]), .config_rst(config_rst)); 
mux6 mux_1464 (.in({n12139_1, n12138_0, n12035_0, n12034_0, n12013_0, n12012_0}), .out(n3245), .config_in(config_chain[4394:4392]), .config_rst(config_rst)); 
mux6 mux_1465 (.in({n13291_0, n13290_0, n13233_0, n13232_0, n13217_0, n13216_1}), .out(n3246), .config_in(config_chain[4397:4395]), .config_rst(config_rst)); 
mux6 mux_1466 (.in({n11863_1, n11862_0, n11855_0, n11854_0, n11847_0, n11846_0}), .out(n3247), .config_in(config_chain[4400:4398]), .config_rst(config_rst)); 
mux6 mux_1467 (.in({n13025_0, n13024_0, n13017_0, n13016_0/**/, n13009_0, n13008_0}), .out(n3248), .config_in(config_chain[4403:4401]), .config_rst(config_rst)); 
mux6 mux_1468 (.in({n12103_0, n12102_0, n12067_0, n12066_0, n12045_0, n12044_0}), .out(n3249), .config_in(config_chain[4406:4404]), .config_rst(config_rst)); 
mux6 mux_1469 (.in({n13255_0, n13254_0, n13249_0, n13248_0, n13241_0, n13240_0}), .out(n3250), .config_in(config_chain[4409:4407]), .config_rst(config_rst)); 
mux6 mux_1470 (.in({n11879_1, n11878_0, n11787_0, n11786_0, n11755_0, n11754_0}), .out(n3251), .config_in(config_chain[4412:4410]), .config_rst(config_rst)); 
mux6 mux_1471 (.in({n13033_0, n13032_0, n12973_0, n12972_0, n12961_0, n12960_1}), .out(n3252), .config_in(config_chain[4415:4413]), .config_rst(config_rst)); 
mux6 mux_1472 (.in({n12125_1, n12124_0, n12119_0, n12118_0, n12111_0, n12110_0}), .out(n3253), .config_in(config_chain[4418:4416]), .config_rst(config_rst)); 
mux6 mux_1473 (.in({n13277_0, n13276_0/**/, n13271_0, n13270_0, n13263_0, n13262_0}), .out(n3254), .config_in(config_chain[4421:4419]), .config_rst(config_rst)); 
mux6 mux_1474 (.in({n11819_0, n11818_0, n11781_0, n11780_0, n11749_0, n11748_0}), .out(n3255), .config_in(config_chain[4424:4422]), .config_rst(config_rst)); 
mux6 mux_1475 (.in({n12995_0, n12994_0, n12981_0, n12980_0, n12969_0, n12968_1}), .out(n3256), .config_in(config_chain[4427:4425]), .config_rst(config_rst)); 
mux6 mux_1476 (.in({n12141_1, n12140_0, n12133_1, n12132_0, n12011_0, n12010_0}), .out(n3257), .config_in(config_chain[4430:4428]), .config_rst(config_rst)); 
mux6 mux_1477 (.in({n13293_0, n13292_0, n13219_0, n13218_1, n13211_0, n13210_1}), .out(n3258), .config_in(config_chain[4433:4431]), .config_rst(config_rst)); 
mux6 mux_1478 (.in({n11865_1, n11864_0, n11849_0, n11848_0, n11813_0/**/, n11812_0}), .out(n3259), .config_in(config_chain[4436:4434]), .config_rst(config_rst)); 
mux6 mux_1479 (.in({n13019_0, n13018_0, n13011_0, n13010_0/**/, n13003_0, n13002_0}), .out(n3260), .config_in(config_chain[4439:4437]), .config_rst(config_rst)); 
mux6 mux_1480 (.in({n12075_0, n12074_0, n12053_0, n12052_0, n12021_0, n12020_0}), .out(n3261), .config_in(config_chain[4442:4440]), .config_rst(config_rst)); 
mux6 mux_1481 (.in({n13257_0, n13256_0, n13243_0, n13242_0/**/, n13227_0, n13226_1}), .out(n3262), .config_in(config_chain[4445:4443]), .config_rst(config_rst)); 
mux6 mux_1482 (.in({n11873_1, n11872_0/**/, n11857_0, n11856_0, n11763_0, n11762_0}), .out(n3263), .config_in(config_chain[4448:4446]), .config_rst(config_rst)); 
mux6 mux_1483 (.in({n13035_0, n13034_0, n13027_0, n13026_0, n12955_0, n12954_1}), .out(n3264), .config_in(config_chain[4451:4449]), .config_rst(config_rst)); 
mux6 mux_1484 (.in({n12113_0, n12112_0/**/, n12105_0, n12104_0, n12085_0, n12084_0}), .out(n3265), .config_in(config_chain[4454:4452]), .config_rst(config_rst)); 
mux6 mux_1485 (.in({n13279_0, n13278_0/**/, n13265_0, n13264_0, n13251_0, n13250_0}), .out(n3266), .config_in(config_chain[4457:4455]), .config_rst(config_rst)); 
mux6 mux_1486 (.in({n11827_0, n11826_0, n11795_0, n11794_0/**/, n11757_0, n11756_0}), .out(n3267), .config_in(config_chain[4460:4458]), .config_rst(config_rst)); 
mux6 mux_1487 (.in({n12983_0, n12982_0, n12975_0, n12974_0, n12971_0, n12970_1}), .out(n3268), .config_in(config_chain[4463:4461]), .config_rst(config_rst)); 
mux6 mux_1488 (.in({n12135_1, n12134_0, n12121_0/**/, n12120_0, n12019_0, n12018_0}), .out(n3269), .config_in(config_chain[4466:4464]), .config_rst(config_rst)); 
mux6 mux_1489 (.in({n13295_0, n13294_0/**/, n13287_0, n13286_0, n13213_0, n13212_1}), .out(n3270), .config_in(config_chain[4469:4467]), .config_rst(config_rst)); 
mux6 mux_1490 (.in({n11851_0, n11850_0, n11843_0, n11842_0, n11821_0, n11820_0/**/}), .out(n3271), .config_in(config_chain[4472:4470]), .config_rst(config_rst)); 
mux6 mux_1491 (.in({n13005_0, n13004_0, n12997_0, n12996_0, n12991_0, n12990_0/**/}), .out(n3272), .config_in(config_chain[4475:4473]), .config_rst(config_rst)); 
mux6 mux_1492 (.in({n12143_1, n12142_0, n12051_0/**/, n12050_0, n12029_0, n12028_0}), .out(n3273), .config_in(config_chain[4478:4476]), .config_rst(config_rst)); 
mux6 mux_1493 (.in({n13237_0, n13236_0, n13229_0, n13228_1, n13221_0, n13220_1}), .out(n3274), .config_in(config_chain[4481:4479]), .config_rst(config_rst)); 
mux6 mux_1494 (.in({n11875_1, n11874_0, n11867_1, n11866_0/**/, n11859_0, n11858_0}), .out(n3275), .config_in(config_chain[4484:4482]), .config_rst(config_rst)); 
mux6 mux_1495 (.in({n13029_0, n13028_0, n13013_0, n13012_0/**/, n12957_0, n12956_1}), .out(n3276), .config_in(config_chain[4487:4485]), .config_rst(config_rst)); 
mux6 mux_1496 (.in({n12107_0, n12106_0, n12093_2, n12092_0, n12061_0, n12060_0}), .out(n3277), .config_in(config_chain[4490:4488]), .config_rst(config_rst)); 
mux6 mux_1497 (.in({n13267_0, n13266_0, n13259_0, n13258_0, n13253_0, n13252_0}), .out(n3278), .config_in(config_chain[4493:4491]), .config_rst(config_rst)); 
mux6 mux_1498 (.in({n11883_2, n11882_0, n11803_0, n11802_0, n11765_0, n11764_0/**/}), .out(n3279), .config_in(config_chain[4496:4494]), .config_rst(config_rst)); 
mux6 mux_1499 (.in({n13037_0, n13036_0/**/, n12977_0, n12976_0, n12965_0, n12964_1}), .out(n3280), .config_in(config_chain[4499:4497]), .config_rst(config_rst)); 
mux6 mux_1500 (.in({n12129_1, n12128_0/**/, n12123_2, n12122_0, n12115_0, n12114_0}), .out(n3281), .config_in(config_chain[4502:4500]), .config_rst(config_rst)); 
mux6 mux_1501 (.in({n13289_0, n13288_0/**/, n13281_0, n13280_0, n13275_0, n13274_0}), .out(n3282), .config_in(config_chain[4505:4503]), .config_rst(config_rst)); 
mux6 mux_1502 (.in({n11845_0, n11844_0, n11835_0, n11834_0, n11797_0, n11796_0}), .out(n3283), .config_in(config_chain[4508:4506]), .config_rst(config_rst)); 
mux6 mux_1503 (.in({n12999_0, n12998_0, n12985_0, n12984_0, n12869_0, n12868_2}), .out(n3284), .config_in(config_chain[4511:4509]), .config_rst(config_rst)); 
mux6 mux_1504 (.in({n12145_2, n12144_0, n12059_0, n12058_0/**/, n12027_0, n12026_0}), .out(n3285), .config_in(config_chain[4514:4512]), .config_rst(config_rst)); 
mux6 mux_1505 (.in({n13297_0, n13296_0, n13239_0, n13238_0, n13223_0, n13222_1}), .out(n3286), .config_in(config_chain[4517:4515]), .config_rst(config_rst)); 
mux6 mux_1506 (.in({n11869_1/**/, n11868_0, n11853_0, n11852_0, n11839_0, n11838_0}), .out(n3287), .config_in(config_chain[4520:4518]), .config_rst(config_rst)); 
mux6 mux_1507 (.in({n13031_0, n13030_0, n13023_0, n13022_0/**/, n12871_0, n12870_2}), .out(n3288), .config_in(config_chain[4523:4521]), .config_rst(config_rst)); 
mux6 mux_1508 (.in({n12099_0, n12098_0, n12069_0/**/, n12068_0, n12037_0, n12036_0}), .out(n3289), .config_in(config_chain[4526:4524]), .config_rst(config_rst)); 
mux6 mux_1509 (.in({n13261_0, n13260_0/**/, n13247_0, n13246_0, n13127_0, n13126_2}), .out(n3290), .config_in(config_chain[4529:4527]), .config_rst(config_rst)); 
mux6 mux_1510 (.in({n11877_1, n11876_0, n11829_2, n11828_0, n11779_0, n11778_0}), .out(n3291), .config_in(config_chain[4532:4530]), .config_rst(config_rst)); 
mux6 mux_1511 (.in({n12993_0, n12992_0, n12967_0, n12966_1, n12959_0, n12958_1}), .out(n3292), .config_in(config_chain[4535:4533]), .config_rst(config_rst)); 
mux6 mux_1512 (.in({n12131_1/**/, n12130_0, n12117_0, n12116_0, n12101_0, n12100_0}), .out(n3293), .config_in(config_chain[4538:4536]), .config_rst(config_rst)); 
mux6 mux_1513 (.in({n13283_0, n13282_0, n13269_0, n13268_0, n13231_0, n13230_1}), .out(n3294), .config_in(config_chain[4541:4539]), .config_rst(config_rst)); 
mux6 mux_1514 (.in({n11861_2, n11860_0, n11805_0, n11804_0, n11773_0, n11772_0}), .out(n3295), .config_in(config_chain[4544:4542]), .config_rst(config_rst)); 
mux6 mux_1515 (.in({n13015_0, n13014_0, n13001_0, n13000_0, n12987_0, n12986_0}), .out(n3296), .config_in(config_chain[4547:4545]), .config_rst(config_rst)); 
mux6 mux_1516 (.in({n12067_0, n12066_0, n12045_0, n12044_0, n12013_0, n12012_0}), .out(n3342), .config_in(config_chain[4550:4548]), .config_rst(config_rst)); 
mux6 mux_1517 (.in({n12133_1, n12132_0, n12125_1, n12124_0, n12119_0, n12118_0}), .out(n3345), .config_in(config_chain[4553:4551]), .config_rst(config_rst)); 
mux6 mux_1518 (.in({n12075_0, n12074_0, n12053_0, n12052_0, n12021_0, n12020_0}), .out(n3348), .config_in(config_chain[4556:4554]), .config_rst(config_rst)); 
mux6 mux_1519 (.in({n12135_1, n12134_0, n12127_1, n12126_0, n12121_0, n12120_0}), .out(n3351), .config_in(config_chain[4559:4557]), .config_rst(config_rst)); 
mux6 mux_1520 (.in({n12083_0, n12082_0, n12051_0, n12050_0, n12029_0, n12028_0}), .out(n3354), .config_in(config_chain[4562:4560]), .config_rst(config_rst)); 
mux6 mux_1521 (.in({n12129_1, n12128_0, n12123_2, n12122_0, n12115_0, n12114_0}), .out(n3357), .config_in(config_chain[4565:4563]), .config_rst(config_rst)); 
mux6 mux_1522 (.in({n12099_0, n12098_0, n12059_0, n12058_0, n12037_0, n12036_0}), .out(n3360), .config_in(config_chain[4568:4566]), .config_rst(config_rst)); 
mux6 mux_1523 (.in({n12131_1, n12130_0, n12117_0, n12116_0, n12091_2, n12090_0}), .out(n3363), .config_in(config_chain[4571:4569]), .config_rst(config_rst)); 
mux6 mux_1524 (.in({n9813_1, n9812_0, n9759_0, n9758_0, n9691_0, n9690_1}), .out(n3390), .config_in(config_chain[4574:4572]), .config_rst(config_rst)); 
mux6 mux_1525 (.in({n9787_0, n9786_0, n9779_0, n9778_0, n9775_0, n9774_0}), .out(n3393), .config_in(config_chain[4577:4575]), .config_rst(config_rst)); 
mux6 mux_1526 (.in({n9815_1, n9814_0, n9699_0, n9698_1, n9667_0, n9666_1}), .out(n3396), .config_in(config_chain[4580:4578]), .config_rst(config_rst)); 
mux6 mux_1527 (.in({n9789_0, n9788_0, n9781_0, n9780_0, n9777_0, n9776_0}), .out(n3399), .config_in(config_chain[4583:4581]), .config_rst(config_rst)); 
mux6 mux_1528 (.in({n9817_1, n9816_0, n9707_0, n9706_1, n9675_0, n9674_1}), .out(n3402), .config_in(config_chain[4586:4584]), .config_rst(config_rst)); 
mux6 mux_1529 (.in({n9783_0, n9782_0, n9771_0, n9770_0, n9753_1, n9752_1}), .out(n3405), .config_in(config_chain[4589:4587]), .config_rst(config_rst)); 
mux6 mux_1530 (.in({n9811_1, n9810_0, n9757_1, n9756_1, n9683_0, n9682_1}), .out(n3408), .config_in(config_chain[4592:4590]), .config_rst(config_rst)); 
mux6 mux_1531 (.in({n9785_0, n9784_0, n9773_0, n9772_0, n9749_1, n9748_1}), .out(n3411), .config_in(config_chain[4595:4593]), .config_rst(config_rst)); 
mux6 mux_1532 (.in({n10053_1, n10052_0, n10039_0, n10038_0, n10027_0, n10026_0}), .out(n3439), .config_in(config_chain[4598:4596]), .config_rst(config_rst)); 
mux6 mux_1533 (.in({n13359_0, n13358_0, n13329_0, n13328_0, n13299_1, n13298_0}), .out(n3440), .config_in(config_chain[4601:4599]), .config_rst(config_rst)); 
mux6 mux_1534 (.in({n9759_0, n9758_0, n9723_0, n9722_1, n9691_0, n9690_1}), .out(n3441), .config_in(config_chain[4604:4602]), .config_rst(config_rst)); 
mux6 mux_1535 (.in({n13095_0, n13094_0, n13073_0, n13072_0, n13041_0, n13040_0}), .out(n3442), .config_in(config_chain[4607:4605]), .config_rst(config_rst)); 
mux6 mux_1536 (.in({n10061_1, n10060_0, n10047_0, n10046_0, n9923_0/**/, n9922_1}), .out(n3443), .config_in(config_chain[4610:4608]), .config_rst(config_rst)); 
mux6 mux_1537 (.in({n13363_1, n13362_0, n13331_1, n13330_0, n13301_0/**/, n13300_0}), .out(n3444), .config_in(config_chain[4613:4611]), .config_rst(config_rst)); 
mux6 mux_1538 (.in({n9787_0, n9786_0, n9779_0, n9778_0, n9775_0, n9774_0}), .out(n3445), .config_in(config_chain[4616:4614]), .config_rst(config_rst)); 
mux6 mux_1539 (.in({n13105_0, n13104_0, n13075_0, n13074_0, n13045_1, n13044_0}), .out(n3446), .config_in(config_chain[4619:4617]), .config_rst(config_rst)); 
mux6 mux_1540 (.in({n10013_0, n10012_0, n9987_0, n9986_1, n9955_0, n9954_1/**/}), .out(n3447), .config_in(config_chain[4622:4620]), .config_rst(config_rst)); 
mux6 mux_1541 (.in({n13365_0, n13364_0, n13333_0, n13332_0, n13303_0, n13302_0}), .out(n3448), .config_in(config_chain[4625:4623]), .config_rst(config_rst)); 
mux6 mux_1542 (.in({n9807_1, n9806_0, n9799_1, n9798_0, n9795_0, n9794_0}), .out(n3449), .config_in(config_chain[4628:4626]), .config_rst(config_rst)); 
mux6 mux_1543 (.in({n13107_0, n13106_0, n13077_1, n13076_0, n13039_0, n13038_0}), .out(n3450), .config_in(config_chain[4631:4629]), .config_rst(config_rst)); 
mux6 mux_1544 (.in({n10033_0, n10032_0, n10029_0, n10028_0, n10021_0, n10020_0}), .out(n3451), .config_in(config_chain[4634:4632]), .config_rst(config_rst)); 
mux6 mux_1545 (.in({n13367_0, n13366_0/**/, n13337_0, n13336_0, n13305_0, n13304_0}), .out(n3452), .config_in(config_chain[4637:4635]), .config_rst(config_rst)); 
mux6 mux_1546 (.in({n9815_1, n9814_0, n9761_0, n9760_0, n9699_0, n9698_1}), .out(n3453), .config_in(config_chain[4640:4638]), .config_rst(config_rst)); 
mux6 mux_1547 (.in({n13103_0/**/, n13102_0, n13071_0, n13070_0, n13049_0, n13048_0}), .out(n3454), .config_in(config_chain[4643:4641]), .config_rst(config_rst)); 
mux6 mux_1548 (.in({n10063_1, n10062_0, n10055_1, n10054_0, n10049_0, n10048_0}), .out(n3455), .config_in(config_chain[4646:4644]), .config_rst(config_rst)); 
mux6 mux_1549 (.in({n13369_0, n13368_0, n13339_1/**/, n13338_0, n13309_0, n13308_0}), .out(n3456), .config_in(config_chain[4649:4647]), .config_rst(config_rst)); 
mux6 mux_1550 (.in({n9781_0, n9780_0, n9769_0/**/, n9768_0, n9731_0, n9730_1}), .out(n3457), .config_in(config_chain[4652:4650]), .config_rst(config_rst)); 
mux6 mux_1551 (.in({n13113_0, n13112_0, n13081_0, n13080_0, n13051_0, n13050_0}), .out(n3458), .config_in(config_chain[4655:4653]), .config_rst(config_rst)); 
mux6 mux_1552 (.in({n10071_1/**/, n10070_0, n9963_0, n9962_1, n9931_0, n9930_1}), .out(n3459), .config_in(config_chain[4658:4656]), .config_rst(config_rst)); 
mux6 mux_1553 (.in({n13371_1/**/, n13370_0, n13341_0, n13340_0, n13311_0, n13310_0}), .out(n3460), .config_in(config_chain[4661:4659]), .config_rst(config_rst)); 
mux6 mux_1554 (.in({n9801_1, n9800_0, n9797_0, n9796_0, n9789_0, n9788_0}), .out(n3461), .config_in(config_chain[4664:4662]), .config_rst(config_rst)); 
mux6 mux_1555 (.in({n13115_0, n13114_0, n13085_1, n13084_0, n13053_1, n13052_0}), .out(n3462), .config_in(config_chain[4667:4665]), .config_rst(config_rst)); 
mux6 mux_1556 (.in({n10035_0, n10034_0, n10023_0/**/, n10022_0, n9995_0, n9994_1}), .out(n3463), .config_in(config_chain[4670:4668]), .config_rst(config_rst)); 
mux6 mux_1557 (.in({n13375_0, n13374_0, n13343_0, n13342_0, n13313_0, n13312_0}), .out(n3464), .config_in(config_chain[4673:4671]), .config_rst(config_rst)); 
mux6 mux_1558 (.in({n9817_1, n9816_0, n9707_0, n9706_1, n9675_0, n9674_1}), .out(n3465), .config_in(config_chain[4676:4674]), .config_rst(config_rst)); 
mux6 mux_1559 (.in({n13117_1, n13116_0, n13079_0/**/, n13078_0, n13047_0, n13046_0}), .out(n3466), .config_in(config_chain[4679:4677]), .config_rst(config_rst)); 
mux6 mux_1560 (.in({n10057_1, n10056_0, n10043_0, n10042_0, n10031_0, n10030_0}), .out(n3467), .config_in(config_chain[4682:4680]), .config_rst(config_rst)); 
mux6 mux_1561 (.in({n13377_0, n13376_0, n13345_0, n13344_0/**/, n13315_1, n13314_0}), .out(n3468), .config_in(config_chain[4685:4683]), .config_rst(config_rst)); 
mux6 mux_1562 (.in({n9771_0, n9770_0, n9763_0, n9762_0, n9739_0, n9738_1/**/}), .out(n3469), .config_in(config_chain[4688:4686]), .config_rst(config_rst)); 
mux6 mux_1563 (.in({n13111_0, n13110_0, n13089_0, n13088_0, n13059_0, n13058_0}), .out(n3470), .config_in(config_chain[4691:4689]), .config_rst(config_rst)); 
mux6 mux_1564 (.in({n10065_1, n10064_0, n10005_1, n10004_1, n9939_0, n9938_1/**/}), .out(n3471), .config_in(config_chain[4694:4692]), .config_rst(config_rst)); 
mux6 mux_1565 (.in({n13383_1, n13382_0, n13349_0, n13348_0, n13317_0/**/, n13316_0}), .out(n3472), .config_in(config_chain[4697:4695]), .config_rst(config_rst)); 
mux6 mux_1566 (.in({n9803_1, n9802_0, n9791_0, n9790_0, n9753_1, n9752_1}), .out(n3473), .config_in(config_chain[4700:4698]), .config_rst(config_rst)); 
mux6 mux_1567 (.in({n13125_2, n13124_0, n13091_0, n13090_0, n13061_1/**/, n13060_0}), .out(n3474), .config_in(config_chain[4703:4701]), .config_rst(config_rst)); 
mux6 mux_1568 (.in({n10017_0/**/, n10016_0, n10007_1, n10006_1, n9971_0, n9970_1}), .out(n3475), .config_in(config_chain[4706:4704]), .config_rst(config_rst)); 
mux6 mux_1569 (.in({n13385_2, n13384_0, n13351_0/**/, n13350_0, n13319_0, n13318_0}), .out(n3476), .config_in(config_chain[4709:4707]), .config_rst(config_rst)); 
mux6 mux_1570 (.in({n9811_1/**/, n9810_0, n9755_1, n9754_1, n9683_0, n9682_1}), .out(n3477), .config_in(config_chain[4712:4710]), .config_rst(config_rst)); 
mux6 mux_1571 (.in({n13129_2, n13128_0, n13093_1, n13092_0, n13055_0, n13054_0/**/}), .out(n3478), .config_in(config_chain[4715:4713]), .config_rst(config_rst)); 
mux6 mux_1572 (.in({n10045_0, n10044_0, n10037_0, n10036_0/**/, n10009_1, n10008_1}), .out(n3479), .config_in(config_chain[4718:4716]), .config_rst(config_rst)); 
mux6 mux_1573 (.in({n13387_2, n13386_0, n13353_0, n13352_0, n13323_1/**/, n13322_0}), .out(n3480), .config_in(config_chain[4721:4719]), .config_rst(config_rst)); 
mux6 mux_1574 (.in({n9765_0/**/, n9764_0, n9747_1, n9746_1, n9715_0, n9714_1}), .out(n3481), .config_in(config_chain[4724:4722]), .config_rst(config_rst)); 
mux6 mux_1575 (.in({n13119_1, n13118_0, n13097_0, n13096_0, n13065_0/**/, n13064_0}), .out(n3482), .config_in(config_chain[4727:4725]), .config_rst(config_rst)); 
mux6 mux_1576 (.in({n10067_1, n10066_0, n10059_1, n10058_0, n10011_1, n10010_1}), .out(n3483), .config_in(config_chain[4730:4728]), .config_rst(config_rst)); 
mux6 mux_1577 (.in({n13389_2, n13388_0, n13355_1, n13354_0, n13325_0, n13324_0}), .out(n3484), .config_in(config_chain[4733:4731]), .config_rst(config_rst)); 
mux6 mux_1578 (.in({n9785_0, n9784_0, n9773_0, n9772_0, n9749_1, n9748_1}), .out(n3485), .config_in(config_chain[4736:4734]), .config_rst(config_rst)); 
mux6 mux_1579 (.in({n13121_1, n13120_0, n13099_0, n13098_0, n13067_0, n13066_0}), .out(n3486), .config_in(config_chain[4739:4737]), .config_rst(config_rst)); 
mux6 mux_1580 (.in({n10019_0, n10018_0, n10001_1, n10000_1, n9979_0, n9978_1/**/}), .out(n3487), .config_in(config_chain[4742:4740]), .config_rst(config_rst)); 
mux6 mux_1581 (.in({n13381_1, n13380_0, n13357_0/**/, n13356_0, n13327_0, n13326_0}), .out(n3488), .config_in(config_chain[4745:4743]), .config_rst(config_rst)); 
mux6 mux_1582 (.in({n9813_1/**/, n9812_0, n9805_1, n9804_0, n9751_1, n9750_1}), .out(n3489), .config_in(config_chain[4748:4746]), .config_rst(config_rst)); 
mux6 mux_1583 (.in({n13123_2, n13122_0, n13101_1, n13100_0, n13063_0, n13062_0}), .out(n3490), .config_in(config_chain[4751:4749]), .config_rst(config_rst)); 
mux6 mux_1584 (.in({n10323_1, n10322_0, n10269_0, n10268_0, n10205_0, n10204_1}), .out(n3537), .config_in(config_chain[4754:4752]), .config_rst(config_rst)); 
mux6 mux_1585 (.in({n13405_1, n13404_0, n13327_0, n13326_0, n13305_0, n13304_0}), .out(n3538), .config_in(config_chain[4757:4755]), .config_rst(config_rst)); 
mux6 mux_1586 (.in({n10053_1, n10052_0, n10047_0, n10046_0, n10039_0, n10038_0}), .out(n3539), .config_in(config_chain[4760:4758]), .config_rst(config_rst)); 
mux6 mux_1587 (.in({n13139_1, n13138_0/**/, n13131_1, n13130_0, n13101_0, n13100_0}), .out(n3540), .config_in(config_chain[4763:4761]), .config_rst(config_rst)); 
mux6 mux_1588 (.in({n10289_0, n10288_0, n10277_0, n10276_0, n10237_0, n10236_1}), .out(n3541), .config_in(config_chain[4766:4764]), .config_rst(config_rst)); 
mux6 mux_1589 (.in({n13369_0, n13368_0, n13337_0, n13336_0, n13299_0, n13298_0}), .out(n3542), .config_in(config_chain[4769:4767]), .config_rst(config_rst)); 
mux6 mux_1590 (.in({n10069_1, n10068_0, n9955_0, n9954_1, n9923_0, n9922_1}), .out(n3543), .config_in(config_chain[4772:4770]), .config_rst(config_rst)); 
mux6 mux_1591 (.in({n13147_1, n13146_0, n13073_0, n13072_0, n13043_0, n13042_0}), .out(n3544), .config_in(config_chain[4775:4773]), .config_rst(config_rst)); 
mux6 mux_1592 (.in({n10309_1, n10308_0, n10305_0, n10304_0, n10297_0, n10296_0}), .out(n3545), .config_in(config_chain[4778:4776]), .config_rst(config_rst)); 
mux6 mux_1593 (.in({n13391_1, n13390_0/**/, n13363_0, n13362_0, n13331_0, n13330_0}), .out(n3546), .config_in(config_chain[4781:4779]), .config_rst(config_rst)); 
mux6 mux_1594 (.in({n10021_0, n10020_0, n10013_0, n10012_0, n9987_0, n9986_1}), .out(n3547), .config_in(config_chain[4784:4782]), .config_rst(config_rst)); 
mux6 mux_1595 (.in({n13105_0, n13104_0, n13075_0, n13074_0, n13045_0, n13044_0}), .out(n3548), .config_in(config_chain[4787:4785]), .config_rst(config_rst)); 
mux6 mux_1596 (.in({n10325_1, n10324_0, n10317_1, n10316_0, n10181_0, n10180_1}), .out(n3549), .config_in(config_chain[4790:4788]), .config_rst(config_rst)); 
mux6 mux_1597 (.in({n13407_1, n13406_0, n13335_0/**/, n13334_0, n13303_0, n13302_0}), .out(n3550), .config_in(config_chain[4793:4791]), .config_rst(config_rst)); 
mux6 mux_1598 (.in({n10055_1, n10054_0, n10041_0, n10040_0, n10029_0, n10028_0}), .out(n3551), .config_in(config_chain[4796:4794]), .config_rst(config_rst)); 
mux6 mux_1599 (.in({n13133_1, n13132_0, n13109_0, n13108_0, n13077_0, n13076_0}), .out(n3552), .config_in(config_chain[4799:4797]), .config_rst(config_rst)); 
mux6 mux_1600 (.in({n10279_0/**/, n10278_0, n10271_0, n10270_0, n10245_0, n10244_1}), .out(n3553), .config_in(config_chain[4802:4800]), .config_rst(config_rst)); 
mux6 mux_1601 (.in({n13367_0, n13366_0, n13345_0, n13344_0, n13307_0, n13306_0}), .out(n3554), .config_in(config_chain[4805:4803]), .config_rst(config_rst)); 
mux6 mux_1602 (.in({n10063_1, n10062_0, n10049_0, n10048_0, n9931_0, n9930_1/**/}), .out(n3555), .config_in(config_chain[4808:4806]), .config_rst(config_rst)); 
mux6 mux_1603 (.in({n13149_1, n13148_0, n13141_1, n13140_0, n13049_0, n13048_0}), .out(n3556), .config_in(config_chain[4811:4809]), .config_rst(config_rst)); 
mux6 mux_1604 (.in({n10299_0/**/, n10298_0, n10291_0, n10290_0, n10287_0, n10286_0}), .out(n3557), .config_in(config_chain[4814:4812]), .config_rst(config_rst)); 
mux6 mux_1605 (.in({n13393_1, n13392_0, n13377_0/**/, n13376_0, n13339_0, n13338_0}), .out(n3558), .config_in(config_chain[4817:4815]), .config_rst(config_rst)); 
mux6 mux_1606 (.in({n10015_0, n10014_0, n9995_0, n9994_1/**/, n9963_0, n9962_1}), .out(n3559), .config_in(config_chain[4820:4818]), .config_rst(config_rst)); 
mux6 mux_1607 (.in({n13113_0, n13112_0/**/, n13083_0, n13082_0, n13051_0, n13050_0}), .out(n3560), .config_in(config_chain[4823:4821]), .config_rst(config_rst)); 
mux6 mux_1608 (.in({n10319_1, n10318_0, n10307_0, n10306_0, n10189_0, n10188_1/**/}), .out(n3561), .config_in(config_chain[4826:4824]), .config_rst(config_rst)); 
mux6 mux_1609 (.in({n13409_1/**/, n13408_0, n13401_1, n13400_0, n13311_0, n13310_0}), .out(n3562), .config_in(config_chain[4829:4827]), .config_rst(config_rst)); 
mux6 mux_1610 (.in({n10043_0/**/, n10042_0, n10035_0, n10034_0, n10031_0, n10030_0}), .out(n3563), .config_in(config_chain[4832:4830]), .config_rst(config_rst)); 
mux6 mux_1611 (.in({n13115_0/**/, n13114_0, n13085_0, n13084_0, n13053_0, n13052_0}), .out(n3564), .config_in(config_chain[4835:4833]), .config_rst(config_rst)); 
mux6 mux_1612 (.in({n10327_1/**/, n10326_0, n10273_0, n10272_0, n10221_0, n10220_1}), .out(n3565), .config_in(config_chain[4838:4836]), .config_rst(config_rst)); 
mux6 mux_1613 (.in({n13375_0, n13374_0, n13343_0, n13342_0, n13321_0, n13320_0}), .out(n3566), .config_in(config_chain[4841:4839]), .config_rst(config_rst)); 
mux6 mux_1614 (.in({n10065_1, n10064_0, n10057_1, n10056_0, n10051_0, n10050_0}), .out(n3567), .config_in(config_chain[4844:4842]), .config_rst(config_rst)); 
mux6 mux_1615 (.in({n13143_1, n13142_0, n13117_0, n13116_0, n13057_0, n13056_0/**/}), .out(n3568), .config_in(config_chain[4847:4845]), .config_rst(config_rst)); 
mux6 mux_1616 (.in({n10293_0, n10292_0, n10281_0, n10280_0, n10259_1, n10258_1}), .out(n3569), .config_in(config_chain[4850:4848]), .config_rst(config_rst)); 
mux6 mux_1617 (.in({n13381_1, n13380_0, n13347_0/**/, n13346_0, n13315_0, n13314_0}), .out(n3570), .config_in(config_chain[4853:4851]), .config_rst(config_rst)); 
mux6 mux_1618 (.in({n10017_0, n10016_0, n10005_1, n10004_1, n9971_0, n9970_1}), .out(n3571), .config_in(config_chain[4856:4854]), .config_rst(config_rst)); 
mux6 mux_1619 (.in({n13123_1, n13122_0, n13089_0, n13088_0/**/, n13059_0, n13058_0}), .out(n3572), .config_in(config_chain[4859:4857]), .config_rst(config_rst)); 
mux6 mux_1620 (.in({n10313_1, n10312_0, n10301_0, n10300_0, n10261_1, n10260_1}), .out(n3573), .config_in(config_chain[4862:4860]), .config_rst(config_rst)); 
mux6 mux_1621 (.in({n13403_1, n13402_0, n13395_1, n13394_0/**/, n13383_1, n13382_0}), .out(n3574), .config_in(config_chain[4865:4863]), .config_rst(config_rst)); 
mux6 mux_1622 (.in({n10037_0, n10036_0, n10025_0, n10024_0, n10007_1, n10006_1}), .out(n3575), .config_in(config_chain[4868:4866]), .config_rst(config_rst)); 
mux6 mux_1623 (.in({n13127_2, n13126_0, n13091_0, n13090_0, n13061_0, n13060_0/**/}), .out(n3576), .config_in(config_chain[4871:4869]), .config_rst(config_rst)); 
mux6 mux_1624 (.in({n10263_1, n10262_1, n10229_0, n10228_1, n10197_0/**/, n10196_1}), .out(n3577), .config_in(config_chain[4874:4872]), .config_rst(config_rst)); 
mux6 mux_1625 (.in({n13385_1, n13384_0, n13351_0, n13350_0, n13329_0, n13328_0}), .out(n3578), .config_in(config_chain[4877:4875]), .config_rst(config_rst)); 
mux6 mux_1626 (.in({n10059_1, n10058_0, n10045_0, n10044_0/**/, n10011_1, n10010_1}), .out(n3579), .config_in(config_chain[4880:4878]), .config_rst(config_rst)); 
mux6 mux_1627 (.in({n13145_1, n13144_0, n13137_1, n13136_0/**/, n13129_2, n13128_0}), .out(n3580), .config_in(config_chain[4883:4881]), .config_rst(config_rst)); 
mux6 mux_1628 (.in({n10283_0, n10282_0, n10275_0, n10274_0, n10265_1, n10264_1}), .out(n3581), .config_in(config_chain[4886:4884]), .config_rst(config_rst)); 
mux6 mux_1629 (.in({n13387_2, n13386_0, n13361_0, n13360_0, n13323_0, n13322_0}), .out(n3582), .config_in(config_chain[4889:4887]), .config_rst(config_rst)); 
mux6 mux_1630 (.in({n10067_1, n10066_0, n10001_1, n10000_1, n9947_0, n9946_1/**/}), .out(n3583), .config_in(config_chain[4892:4890]), .config_rst(config_rst)); 
mux6 mux_1631 (.in({n13119_1, n13118_0, n13097_0/**/, n13096_0, n13065_0, n13064_0}), .out(n3584), .config_in(config_chain[4895:4893]), .config_rst(config_rst)); 
mux6 mux_1632 (.in({n10315_1, n10314_0, n10303_0, n10302_0, n10267_1, n10266_1}), .out(n3585), .config_in(config_chain[4898:4896]), .config_rst(config_rst)); 
mux6 mux_1633 (.in({n13397_1, n13396_0, n13379_0, n13378_0, n13355_0, n13354_0}), .out(n3586), .config_in(config_chain[4901:4899]), .config_rst(config_rst)); 
mux6 mux_1634 (.in({n10027_0, n10026_0, n10019_0, n10018_0, n10003_1, n10002_1}), .out(n3587), .config_in(config_chain[4904:4902]), .config_rst(config_rst)); 
mux6 mux_1635 (.in({n13121_1, n13120_0, n13099_0, n13098_0, n13069_0, n13068_0}), .out(n3588), .config_in(config_chain[4907:4905]), .config_rst(config_rst)); 
mux6 mux_1636 (.in({n10567_1, n10566_0, n10553_0, n10552_0, n10541_0, n10540_0}), .out(n3635), .config_in(config_chain[4910:4908]), .config_rst(config_rst)); 
mux6 mux_1637 (.in({n13411_1, n13410_0, n13397_0, n13396_0, n13355_0, n13354_0}), .out(n3636), .config_in(config_chain[4913:4911]), .config_rst(config_rst)); 
mux6 mux_1638 (.in({n10269_0, n10268_0, n10237_0, n10236_1, n10205_0, n10204_1}), .out(n3637), .config_in(config_chain[4916:4914]), .config_rst(config_rst)); 
mux6 mux_1639 (.in({n13099_0, n13098_0, n13077_0/**/, n13076_0, n13045_0, n13044_0}), .out(n3638), .config_in(config_chain[4919:4917]), .config_rst(config_rst)); 
mux6 mux_1640 (.in({n10575_1, n10574_0, n10561_0, n10560_0, n10441_0, n10440_1}), .out(n3639), .config_in(config_chain[4922:4920]), .config_rst(config_rst)); 
mux6 mux_1641 (.in({n13427_1, n13426_0, n13419_1, n13418_0, n13305_0, n13304_0}), .out(n3640), .config_in(config_chain[4925:4923]), .config_rst(config_rst)); 
mux6 mux_1642 (.in({n10297_0, n10296_0, n10289_0, n10288_0, n10285_0, n10284_0}), .out(n3641), .config_in(config_chain[4928:4926]), .config_rst(config_rst)); 
mux6 mux_1643 (.in({n13151_1, n13150_0/**/, n13139_0, n13138_0, n13109_0, n13108_0}), .out(n3642), .config_in(config_chain[4931:4929]), .config_rst(config_rst)); 
mux6 mux_1644 (.in({n10527_0, n10526_0, n10505_0, n10504_1, n10473_0, n10472_1}), .out(n3643), .config_in(config_chain[4934:4932]), .config_rst(config_rst)); 
mux6 mux_1645 (.in({n13369_0, n13368_0, n13337_0, n13336_0, n13299_0, n13298_0}), .out(n3644), .config_in(config_chain[4937:4935]), .config_rst(config_rst)); 
mux6 mux_1646 (.in({n10317_1, n10316_0, n10309_1, n10308_0, n10305_0, n10304_0/**/}), .out(n3645), .config_in(config_chain[4940:4938]), .config_rst(config_rst)); 
mux6 mux_1647 (.in({n13159_1, n13158_0, n13147_0/**/, n13146_0, n13043_0, n13042_0}), .out(n3646), .config_in(config_chain[4943:4941]), .config_rst(config_rst)); 
mux6 mux_1648 (.in({n10547_0, n10546_0, n10543_0, n10542_0, n10535_0, n10534_0/**/}), .out(n3647), .config_in(config_chain[4946:4944]), .config_rst(config_rst)); 
mux6 mux_1649 (.in({n13399_0, n13398_0, n13391_0, n13390_0, n13363_0, n13362_0/**/}), .out(n3648), .config_in(config_chain[4949:4947]), .config_rst(config_rst)); 
mux6 mux_1650 (.in({n10325_1, n10324_0, n10271_0, n10270_0, n10213_0, n10212_1}), .out(n3649), .config_in(config_chain[4952:4950]), .config_rst(config_rst)); 
mux6 mux_1651 (.in({n13107_0, n13106_0, n13075_0, n13074_0, n13053_0/**/, n13052_0}), .out(n3650), .config_in(config_chain[4955:4953]), .config_rst(config_rst)); 
mux6 mux_1652 (.in({n10577_1, n10576_0, n10569_1, n10568_0/**/, n10563_0, n10562_0}), .out(n3651), .config_in(config_chain[4958:4956]), .config_rst(config_rst)); 
mux6 mux_1653 (.in({n13421_1, n13420_0, n13407_0, n13406_0, n13313_0/**/, n13312_0}), .out(n3652), .config_in(config_chain[4961:4959]), .config_rst(config_rst)); 
mux6 mux_1654 (.in({n10291_0/**/, n10290_0, n10279_0, n10278_0, n10245_0, n10244_1}), .out(n3653), .config_in(config_chain[4964:4962]), .config_rst(config_rst)); 
mux6 mux_1655 (.in({n13133_0, n13132_0/**/, n13117_0, n13116_0, n13085_0, n13084_0}), .out(n3654), .config_in(config_chain[4967:4965]), .config_rst(config_rst)); 
mux6 mux_1656 (.in({n10585_1, n10584_0, n10481_0, n10480_1, n10449_0, n10448_1}), .out(n3655), .config_in(config_chain[4970:4968]), .config_rst(config_rst)); 
mux6 mux_1657 (.in({n13429_1, n13428_0, n13345_0, n13344_0, n13307_0/**/, n13306_0}), .out(n3656), .config_in(config_chain[4973:4971]), .config_rst(config_rst)); 
mux6 mux_1658 (.in({n10311_1, n10310_0, n10307_0, n10306_0, n10299_0, n10298_0}), .out(n3657), .config_in(config_chain[4976:4974]), .config_rst(config_rst)); 
mux6 mux_1659 (.in({n13161_1, n13160_0, n13153_1, n13152_0/**/, n13149_0, n13148_0}), .out(n3658), .config_in(config_chain[4979:4977]), .config_rst(config_rst)); 
mux6 mux_1660 (.in({n10549_0/**/, n10548_0, n10537_0, n10536_0, n10513_0, n10512_1}), .out(n3659), .config_in(config_chain[4982:4980]), .config_rst(config_rst)); 
mux6 mux_1661 (.in({n13393_0/**/, n13392_0, n13371_0, n13370_0, n13339_0, n13338_0}), .out(n3660), .config_in(config_chain[4985:4983]), .config_rst(config_rst)); 
mux6 mux_1662 (.in({n10327_1, n10326_0, n10221_0, n10220_1, n10189_0/**/, n10188_1}), .out(n3661), .config_in(config_chain[4988:4986]), .config_rst(config_rst)); 
mux6 mux_1663 (.in({n13169_1, n13168_0, n13083_0, n13082_0, n13051_0, n13050_0}), .out(n3662), .config_in(config_chain[4991:4989]), .config_rst(config_rst)); 
mux6 mux_1664 (.in({n10571_1, n10570_0, n10557_0/**/, n10556_0, n10545_0, n10544_0}), .out(n3663), .config_in(config_chain[4994:4992]), .config_rst(config_rst)); 
mux6 mux_1665 (.in({n13415_1, n13414_0, n13409_0, n13408_0, n13401_0, n13400_0/**/}), .out(n3664), .config_in(config_chain[4997:4995]), .config_rst(config_rst)); 
mux6 mux_1666 (.in({n10281_0, n10280_0, n10273_0, n10272_0, n10253_0, n10252_1}), .out(n3665), .config_in(config_chain[5000:4998]), .config_rst(config_rst)); 
mux6 mux_1667 (.in({n13135_0, n13134_0, n13115_0, n13114_0/**/, n13093_0, n13092_0}), .out(n3666), .config_in(config_chain[5003:5001]), .config_rst(config_rst)); 
mux6 mux_1668 (.in({n10579_1, n10578_0, n10515_0, n10514_1, n10457_0, n10456_1}), .out(n3667), .config_in(config_chain[5006:5004]), .config_rst(config_rst)); 
mux6 mux_1669 (.in({n13379_0, n13378_0, n13353_0, n13352_0/**/, n13321_0, n13320_0}), .out(n3668), .config_in(config_chain[5009:5007]), .config_rst(config_rst)); 
mux6 mux_1670 (.in({n10313_1, n10312_0/**/, n10301_0, n10300_0, n10259_1, n10258_1}), .out(n3669), .config_in(config_chain[5012:5010]), .config_rst(config_rst)); 
mux6 mux_1671 (.in({n13155_1, n13154_0, n13143_0, n13142_0, n13121_1, n13120_0}), .out(n3670), .config_in(config_chain[5015:5013]), .config_rst(config_rst)); 
mux6 mux_1672 (.in({n10531_0, n10530_0, n10517_0, n10516_1, n10489_0, n10488_1}), .out(n3671), .config_in(config_chain[5018:5016]), .config_rst(config_rst)); 
mux6 mux_1673 (.in({n13381_0, n13380_0, n13347_0, n13346_0, n13315_0/**/, n13314_0}), .out(n3672), .config_in(config_chain[5021:5019]), .config_rst(config_rst)); 
mux6 mux_1674 (.in({n10321_1, n10320_0/**/, n10261_1, n10260_1, n10197_0, n10196_1}), .out(n3673), .config_in(config_chain[5024:5022]), .config_rst(config_rst)); 
mux6 mux_1675 (.in({n13163_1, n13162_0, n13125_1, n13124_0, n13059_0, n13058_0/**/}), .out(n3674), .config_in(config_chain[5027:5025]), .config_rst(config_rst)); 
mux6 mux_1676 (.in({n10559_0, n10558_0, n10551_0, n10550_0, n10519_1, n10518_1}), .out(n3675), .config_in(config_chain[5030:5028]), .config_rst(config_rst)); 
mux6 mux_1677 (.in({n13417_1, n13416_0, n13403_0, n13402_0/**/, n13383_1, n13382_0}), .out(n3676), .config_in(config_chain[5033:5031]), .config_rst(config_rst)); 
mux6 mux_1678 (.in({n10275_0, n10274_0, n10265_1, n10264_1, n10229_0, n10228_1}), .out(n3677), .config_in(config_chain[5036:5034]), .config_rst(config_rst)); 
mux6 mux_1679 (.in({n13127_2, n13126_0, n13101_0/**/, n13100_0, n13069_0, n13068_0}), .out(n3678), .config_in(config_chain[5039:5037]), .config_rst(config_rst)); 
mux6 mux_1680 (.in({n10581_1, n10580_0, n10573_1, n10572_0, n10521_1, n10520_1}), .out(n3679), .config_in(config_chain[5042:5040]), .config_rst(config_rst)); 
mux6 mux_1681 (.in({n13425_1/**/, n13424_0, n13385_1, n13384_0, n13329_0, n13328_0}), .out(n3680), .config_in(config_chain[5045:5043]), .config_rst(config_rst)); 
mux6 mux_1682 (.in({n10295_0, n10294_0, n10283_0, n10282_0, n10267_1, n10266_1}), .out(n3681), .config_in(config_chain[5048:5046]), .config_rst(config_rst)); 
mux6 mux_1683 (.in({n13145_0, n13144_0, n13137_0, n13136_0/**/, n13129_2, n13128_0}), .out(n3682), .config_in(config_chain[5051:5049]), .config_rst(config_rst)); 
mux6 mux_1684 (.in({n10533_0/**/, n10532_0, n10523_1, n10522_1, n10497_0, n10496_1}), .out(n3683), .config_in(config_chain[5054:5052]), .config_rst(config_rst)); 
mux6 mux_1685 (.in({n13389_2, n13388_0, n13361_0, n13360_0, n13323_0, n13322_0/**/}), .out(n3684), .config_in(config_chain[5057:5055]), .config_rst(config_rst)); 
mux6 mux_1686 (.in({n10323_1, n10322_0, n10315_1, n10314_0, n10257_0, n10256_1}), .out(n3685), .config_in(config_chain[5060:5058]), .config_rst(config_rst)); 
mux6 mux_1687 (.in({n13165_1/**/, n13164_0, n13119_0, n13118_0, n13067_0, n13066_0}), .out(n3686), .config_in(config_chain[5063:5061]), .config_rst(config_rst)); 
mux6 mux_1688 (.in({n10841_1, n10840_0, n10787_0, n10786_0, n10719_0, n10718_1}), .out(n3733), .config_in(config_chain[5066:5064]), .config_rst(config_rst)); 
mux6 mux_1689 (.in({n13445_1, n13444_0, n13391_0, n13390_0, n13323_0, n13322_1}), .out(n3734), .config_in(config_chain[5069:5067]), .config_rst(config_rst)); 
mux6 mux_1690 (.in({n10567_1, n10566_0, n10561_0, n10560_0, n10553_0, n10552_0}), .out(n3735), .config_in(config_chain[5072:5070]), .config_rst(config_rst)); 
mux6 mux_1691 (.in({n13179_1, n13178_0, n13171_1, n13170_0, n13165_0, n13164_0}), .out(n3736), .config_in(config_chain[5075:5073]), .config_rst(config_rst)); 
mux6 mux_1692 (.in({n10807_0, n10806_0, n10795_0, n10794_0, n10751_0, n10750_1}), .out(n3737), .config_in(config_chain[5078:5076]), .config_rst(config_rst)); 
mux6 mux_1693 (.in({n13411_0, n13410_0, n13407_0, n13406_0, n13399_0, n13398_0}), .out(n3738), .config_in(config_chain[5081:5079]), .config_rst(config_rst)); 
mux6 mux_1694 (.in({n10583_1, n10582_0, n10473_0, n10472_1, n10441_0, n10440_1}), .out(n3739), .config_in(config_chain[5084:5082]), .config_rst(config_rst)); 
mux6 mux_1695 (.in({n13187_1, n13186_0, n13131_0, n13130_0, n13077_0, n13076_1}), .out(n3740), .config_in(config_chain[5087:5085]), .config_rst(config_rst)); 
mux6 mux_1696 (.in({n10827_1, n10826_0, n10823_0, n10822_0, n10815_0, n10814_0}), .out(n3741), .config_in(config_chain[5090:5088]), .config_rst(config_rst)); 
mux6 mux_1697 (.in({n13431_1, n13430_0, n13427_0, n13426_0, n13419_0, n13418_0}), .out(n3742), .config_in(config_chain[5093:5091]), .config_rst(config_rst)); 
mux6 mux_1698 (.in({n10535_0, n10534_0, n10527_0, n10526_0, n10505_0, n10504_1}), .out(n3743), .config_in(config_chain[5096:5094]), .config_rst(config_rst)); 
mux6 mux_1699 (.in({n13151_0, n13150_0, n13139_0, n13138_0/**/, n13109_0, n13108_1}), .out(n3744), .config_in(config_chain[5099:5097]), .config_rst(config_rst)); 
mux6 mux_1700 (.in({n10843_1, n10842_0, n10835_1, n10834_0, n10695_0, n10694_1}), .out(n3745), .config_in(config_chain[5102:5100]), .config_rst(config_rst)); 
mux6 mux_1701 (.in({n13447_1/**/, n13446_0, n13331_0, n13330_1, n13299_0, n13298_1}), .out(n3746), .config_in(config_chain[5105:5103]), .config_rst(config_rst)); 
mux6 mux_1702 (.in({n10569_1, n10568_0, n10555_0, n10554_0, n10543_0/**/, n10542_0}), .out(n3747), .config_in(config_chain[5108:5106]), .config_rst(config_rst)); 
mux6 mux_1703 (.in({n13173_1, n13172_0, n13167_0, n13166_0, n13159_0, n13158_0}), .out(n3748), .config_in(config_chain[5111:5109]), .config_rst(config_rst)); 
mux6 mux_1704 (.in({n10797_0, n10796_0, n10789_0, n10788_0, n10759_0, n10758_1/**/}), .out(n3749), .config_in(config_chain[5114:5112]), .config_rst(config_rst)); 
mux6 mux_1705 (.in({n13413_0, n13412_0/**/, n13401_0, n13400_0, n13363_0, n13362_1}), .out(n3750), .config_in(config_chain[5117:5115]), .config_rst(config_rst)); 
mux6 mux_1706 (.in({n10577_1, n10576_0, n10563_0, n10562_0, n10449_0, n10448_1}), .out(n3751), .config_in(config_chain[5120:5118]), .config_rst(config_rst)); 
mux6 mux_1707 (.in({n13189_1/**/, n13188_0, n13181_1, n13180_0, n13053_0, n13052_1}), .out(n3752), .config_in(config_chain[5123:5121]), .config_rst(config_rst)); 
mux6 mux_1708 (.in({n10817_0, n10816_0, n10809_0, n10808_0, n10805_0/**/, n10804_0}), .out(n3753), .config_in(config_chain[5126:5124]), .config_rst(config_rst)); 
mux6 mux_1709 (.in({n13433_1, n13432_0/**/, n13421_0, n13420_0, n13409_0, n13408_0}), .out(n3754), .config_in(config_chain[5129:5127]), .config_rst(config_rst)); 
mux6 mux_1710 (.in({n10529_0, n10528_0, n10513_0/**/, n10512_1, n10481_0, n10480_1}), .out(n3755), .config_in(config_chain[5132:5130]), .config_rst(config_rst)); 
mux6 mux_1711 (.in({n13141_0, n13140_0, n13133_0, n13132_0, n13117_0, n13116_1}), .out(n3756), .config_in(config_chain[5135:5133]), .config_rst(config_rst)); 
mux6 mux_1712 (.in({n10837_1, n10836_0, n10825_0, n10824_0, n10703_0, n10702_1}), .out(n3757), .config_in(config_chain[5138:5136]), .config_rst(config_rst)); 
mux6 mux_1713 (.in({n13449_1, n13448_0, n13441_1, n13440_0, n13307_0, n13306_1}), .out(n3758), .config_in(config_chain[5141:5139]), .config_rst(config_rst)); 
mux6 mux_1714 (.in({n10557_0, n10556_0/**/, n10549_0, n10548_0, n10545_0, n10544_0}), .out(n3759), .config_in(config_chain[5144:5142]), .config_rst(config_rst)); 
mux6 mux_1715 (.in({n13161_0, n13160_0, n13153_0/**/, n13152_0, n13149_0, n13148_0}), .out(n3760), .config_in(config_chain[5147:5145]), .config_rst(config_rst)); 
mux6 mux_1716 (.in({n10845_1, n10844_0, n10791_0, n10790_0, n10735_0, n10734_1/**/}), .out(n3761), .config_in(config_chain[5150:5148]), .config_rst(config_rst)); 
mux6 mux_1717 (.in({n13395_0, n13394_0, n13371_0, n13370_1, n13339_0, n13338_1}), .out(n3762), .config_in(config_chain[5153:5151]), .config_rst(config_rst)); 
mux6 mux_1718 (.in({n10579_1, n10578_0, n10571_1, n10570_0, n10565_0, n10564_0/**/}), .out(n3763), .config_in(config_chain[5156:5154]), .config_rst(config_rst)); 
mux6 mux_1719 (.in({n13183_1/**/, n13182_0, n13169_0, n13168_0, n13061_0, n13060_1}), .out(n3764), .config_in(config_chain[5159:5157]), .config_rst(config_rst)); 
mux6 mux_1720 (.in({n10811_0/**/, n10810_0, n10799_0, n10798_0, n10785_1, n10784_1}), .out(n3765), .config_in(config_chain[5162:5160]), .config_rst(config_rst)); 
mux6 mux_1721 (.in({n13423_0, n13422_0, n13415_0, n13414_0/**/, n13389_1, n13388_1}), .out(n3766), .config_in(config_chain[5165:5163]), .config_rst(config_rst)); 
mux6 mux_1722 (.in({n10531_0, n10530_0, n10515_0, n10514_1, n10489_0, n10488_1}), .out(n3767), .config_in(config_chain[5168:5166]), .config_rst(config_rst)); 
mux6 mux_1723 (.in({n13135_0/**/, n13134_0, n13119_0, n13118_1, n13093_0, n13092_1}), .out(n3768), .config_in(config_chain[5171:5169]), .config_rst(config_rst)); 
mux6 mux_1724 (.in({n10831_1, n10830_0/**/, n10819_0, n10818_0, n10775_0, n10774_1}), .out(n3769), .config_in(config_chain[5174:5172]), .config_rst(config_rst)); 
mux6 mux_1725 (.in({n13443_1, n13442_0, n13435_1/**/, n13434_0, n13379_0, n13378_1}), .out(n3770), .config_in(config_chain[5177:5175]), .config_rst(config_rst)); 
mux6 mux_1726 (.in({n10551_0, n10550_0, n10539_0/**/, n10538_0, n10517_0, n10516_1}), .out(n3771), .config_in(config_chain[5180:5178]), .config_rst(config_rst)); 
mux6 mux_1727 (.in({n13155_0, n13154_0, n13143_0, n13142_0/**/, n13123_1, n13122_1}), .out(n3772), .config_in(config_chain[5183:5181]), .config_rst(config_rst)); 
mux6 mux_1728 (.in({n10777_0, n10776_1, n10743_0, n10742_1, n10711_0, n10710_1/**/}), .out(n3773), .config_in(config_chain[5186:5184]), .config_rst(config_rst)); 
mux6 mux_1729 (.in({n13397_0, n13396_0, n13381_0, n13380_1, n13347_0, n13346_1}), .out(n3774), .config_in(config_chain[5189:5187]), .config_rst(config_rst)); 
mux6 mux_1730 (.in({n10573_1, n10572_0, n10559_0, n10558_0, n10521_1, n10520_1}), .out(n3775), .config_in(config_chain[5192:5190]), .config_rst(config_rst)); 
mux6 mux_1731 (.in({n13185_1/**/, n13184_0, n13177_1, n13176_0, n13125_1, n13124_1}), .out(n3776), .config_in(config_chain[5195:5193]), .config_rst(config_rst)); 
mux6 mux_1732 (.in({n10801_0/**/, n10800_0, n10793_0, n10792_0, n10779_0, n10778_1}), .out(n3777), .config_in(config_chain[5198:5196]), .config_rst(config_rst)); 
mux6 mux_1733 (.in({n13417_0, n13416_0, n13405_0, n13404_0, n13383_0, n13382_1}), .out(n3778), .config_in(config_chain[5201:5199]), .config_rst(config_rst)); 
mux6 mux_1734 (.in({n10581_1, n10580_0, n10523_1, n10522_1, n10465_0, n10464_1}), .out(n3779), .config_in(config_chain[5204:5202]), .config_rst(config_rst)); 
mux6 mux_1735 (.in({n13127_1, n13126_1, n13101_0, n13100_1, n13069_0, n13068_1}), .out(n3780), .config_in(config_chain[5207:5205]), .config_rst(config_rst)); 
mux6 mux_1736 (.in({n10833_1, n10832_0, n10821_0, n10820_0/**/, n10781_1, n10780_1}), .out(n3781), .config_in(config_chain[5210:5208]), .config_rst(config_rst)); 
mux6 mux_1737 (.in({n13437_1, n13436_0, n13425_0, n13424_0, n13387_1, n13386_1}), .out(n3782), .config_in(config_chain[5213:5211]), .config_rst(config_rst)); 
mux6 mux_1738 (.in({n10541_0, n10540_0, n10533_0, n10532_0, n10525_1, n10524_1}), .out(n3783), .config_in(config_chain[5216:5214]), .config_rst(config_rst)); 
mux6 mux_1739 (.in({n13157_0, n13156_0, n13145_0, n13144_0, n13129_1, n13128_1}), .out(n3784), .config_in(config_chain[5219:5217]), .config_rst(config_rst)); 
mux6 mux_1740 (.in({n11089_1, n11088_0, n11075_0, n11074_0, n11063_0, n11062_0}), .out(n3831), .config_in(config_chain[5222:5220]), .config_rst(config_rst)); 
mux6 mux_1741 (.in({n13451_1, n13450_0, n13437_0, n13436_0, n13425_0, n13424_0}), .out(n3832), .config_in(config_chain[5225:5223]), .config_rst(config_rst)); 
mux6 mux_1742 (.in({n10787_0, n10786_0, n10751_0, n10750_1, n10719_0, n10718_1}), .out(n3833), .config_in(config_chain[5228:5226]), .config_rst(config_rst)); 
mux6 mux_1743 (.in({n13159_0/**/, n13158_0, n13151_0, n13150_0, n13145_0, n13144_1}), .out(n3834), .config_in(config_chain[5231:5229]), .config_rst(config_rst)); 
mux6 mux_1744 (.in({n11097_1, n11096_0, n11083_0, n11082_0, n10959_0, n10958_1}), .out(n3835), .config_in(config_chain[5234:5232]), .config_rst(config_rst)); 
mux6 mux_1745 (.in({n13467_1, n13466_0, n13459_1, n13458_0, n13391_0, n13390_1/**/}), .out(n3836), .config_in(config_chain[5237:5235]), .config_rst(config_rst)); 
mux6 mux_1746 (.in({n10815_0, n10814_0, n10807_0, n10806_0, n10803_0, n10802_0}), .out(n3837), .config_in(config_chain[5240:5238]), .config_rst(config_rst)); 
mux6 mux_1747 (.in({n13191_1, n13190_0, n13179_0, n13178_0, n13167_0, n13166_0}), .out(n3838), .config_in(config_chain[5243:5241]), .config_rst(config_rst)); 
mux6 mux_1748 (.in({n11049_0, n11048_0, n11023_0, n11022_1, n10991_0, n10990_1}), .out(n3839), .config_in(config_chain[5246:5244]), .config_rst(config_rst)); 
mux6 mux_1749 (.in({n13411_0, n13410_0, n13407_0, n13406_1/**/, n13399_0, n13398_1}), .out(n3840), .config_in(config_chain[5249:5247]), .config_rst(config_rst)); 
mux6 mux_1750 (.in({n10835_1, n10834_0/**/, n10827_1, n10826_0, n10823_0, n10822_0}), .out(n3841), .config_in(config_chain[5252:5250]), .config_rst(config_rst)); 
mux6 mux_1751 (.in({n13199_1/**/, n13198_0, n13187_0, n13186_0, n13131_0, n13130_1}), .out(n3842), .config_in(config_chain[5255:5253]), .config_rst(config_rst)); 
mux6 mux_1752 (.in({n11069_0, n11068_0, n11065_0, n11064_0, n11057_0, n11056_0}), .out(n3843), .config_in(config_chain[5258:5256]), .config_rst(config_rst)); 
mux6 mux_1753 (.in({n13439_0, n13438_0, n13431_0, n13430_0, n13427_0, n13426_0}), .out(n3844), .config_in(config_chain[5261:5259]), .config_rst(config_rst)); 
mux6 mux_1754 (.in({n10843_1, n10842_0, n10789_0, n10788_0/**/, n10727_0, n10726_1}), .out(n3845), .config_in(config_chain[5264:5262]), .config_rst(config_rst)); 
mux6 mux_1755 (.in({n13153_0, n13152_0, n13147_0, n13146_1, n13139_0, n13138_1}), .out(n3846), .config_in(config_chain[5267:5265]), .config_rst(config_rst)); 
mux6 mux_1756 (.in({n11099_1, n11098_0, n11091_1, n11090_0, n11085_0, n11084_0/**/}), .out(n3847), .config_in(config_chain[5270:5268]), .config_rst(config_rst)); 
mux6 mux_1757 (.in({n13461_1, n13460_0, n13447_0, n13446_0/**/, n13393_0, n13392_1}), .out(n3848), .config_in(config_chain[5273:5271]), .config_rst(config_rst)); 
mux6 mux_1758 (.in({n10809_0, n10808_0, n10797_0/**/, n10796_0, n10759_0, n10758_1}), .out(n3849), .config_in(config_chain[5276:5274]), .config_rst(config_rst)); 
mux6 mux_1759 (.in({n13173_0, n13172_0, n13169_0, n13168_0, n13161_0, n13160_0}), .out(n3850), .config_in(config_chain[5279:5277]), .config_rst(config_rst)); 
mux6 mux_1760 (.in({n11107_1, n11106_0, n10999_0, n10998_1, n10967_0, n10966_1/**/}), .out(n3851), .config_in(config_chain[5282:5280]), .config_rst(config_rst)); 
mux6 mux_1761 (.in({n13469_1, n13468_0, n13413_0, n13412_0, n13401_0/**/, n13400_1}), .out(n3852), .config_in(config_chain[5285:5283]), .config_rst(config_rst)); 
mux6 mux_1762 (.in({n10829_1, n10828_0, n10825_0, n10824_0, n10817_0, n10816_0/**/}), .out(n3853), .config_in(config_chain[5288:5286]), .config_rst(config_rst)); 
mux6 mux_1763 (.in({n13201_1, n13200_0, n13193_1/**/, n13192_0, n13189_0, n13188_0}), .out(n3854), .config_in(config_chain[5291:5289]), .config_rst(config_rst)); 
mux6 mux_1764 (.in({n11071_0, n11070_0, n11059_0, n11058_0, n11031_0/**/, n11030_1}), .out(n3855), .config_in(config_chain[5294:5292]), .config_rst(config_rst)); 
mux6 mux_1765 (.in({n13433_0, n13432_0, n13429_0, n13428_0, n13421_0, n13420_0}), .out(n3856), .config_in(config_chain[5297:5295]), .config_rst(config_rst)); 
mux6 mux_1766 (.in({n10845_1, n10844_0, n10735_0, n10734_1, n10703_0, n10702_1/**/}), .out(n3857), .config_in(config_chain[5300:5298]), .config_rst(config_rst)); 
mux6 mux_1767 (.in({n13209_1, n13208_0, n13141_0, n13140_1, n13133_0, n13132_1}), .out(n3858), .config_in(config_chain[5303:5301]), .config_rst(config_rst)); 
mux6 mux_1768 (.in({n11093_1, n11092_0, n11079_0, n11078_0, n11067_0, n11066_0}), .out(n3859), .config_in(config_chain[5306:5304]), .config_rst(config_rst)); 
mux6 mux_1769 (.in({n13455_1, n13454_0, n13449_0, n13448_0, n13441_0, n13440_0}), .out(n3860), .config_in(config_chain[5309:5307]), .config_rst(config_rst)); 
mux6 mux_1770 (.in({n10799_0, n10798_0, n10791_0, n10790_0, n10767_0/**/, n10766_1}), .out(n3861), .config_in(config_chain[5312:5310]), .config_rst(config_rst)); 
mux6 mux_1771 (.in({n13175_0, n13174_0, n13163_0, n13162_0/**/, n13149_0, n13148_1}), .out(n3862), .config_in(config_chain[5315:5313]), .config_rst(config_rst)); 
mux6 mux_1772 (.in({n11101_1, n11100_0, n11045_1, n11044_1, n10975_0, n10974_1/**/}), .out(n3863), .config_in(config_chain[5318:5316]), .config_rst(config_rst)); 
mux6 mux_1773 (.in({n13403_0, n13402_1, n13395_0, n13394_1, n13387_1, n13386_1}), .out(n3864), .config_in(config_chain[5321:5319]), .config_rst(config_rst)); 
mux6 mux_1774 (.in({n10831_1, n10830_0, n10819_0, n10818_0, n10785_1, n10784_1}), .out(n3865), .config_in(config_chain[5324:5322]), .config_rst(config_rst)); 
mux6 mux_1775 (.in({n13195_1/**/, n13194_0, n13183_0, n13182_0, n13129_1, n13128_1}), .out(n3866), .config_in(config_chain[5327:5325]), .config_rst(config_rst)); 
mux6 mux_1776 (.in({n11053_0, n11052_0, n11047_1, n11046_1, n11007_0, n11006_1}), .out(n3867), .config_in(config_chain[5330:5328]), .config_rst(config_rst)); 
mux6 mux_1777 (.in({n13423_0/**/, n13422_0, n13415_0, n13414_0, n13389_1, n13388_1}), .out(n3868), .config_in(config_chain[5333:5331]), .config_rst(config_rst)); 
mux6 mux_1778 (.in({n10839_1/**/, n10838_0, n10775_0, n10774_1, n10711_0, n10710_1}), .out(n3869), .config_in(config_chain[5336:5334]), .config_rst(config_rst)); 
mux6 mux_1779 (.in({n13203_1, n13202_0, n13135_0, n13134_1/**/, n13121_0, n13120_1}), .out(n3870), .config_in(config_chain[5339:5337]), .config_rst(config_rst)); 
mux6 mux_1780 (.in({n11109_1, n11108_0, n11081_0, n11080_0, n11073_0, n11072_0/**/}), .out(n3871), .config_in(config_chain[5342:5340]), .config_rst(config_rst)); 
mux6 mux_1781 (.in({n13471_1, n13470_0, n13457_1, n13456_0, n13443_0, n13442_0}), .out(n3872), .config_in(config_chain[5345:5343]), .config_rst(config_rst)); 
mux6 mux_1782 (.in({n10793_0/**/, n10792_0, n10779_0, n10778_1, n10743_0, n10742_1}), .out(n3873), .config_in(config_chain[5348:5346]), .config_rst(config_rst)); 
mux6 mux_1783 (.in({n13165_0, n13164_0/**/, n13157_0, n13156_0, n13123_0, n13122_1}), .out(n3874), .config_in(config_chain[5351:5349]), .config_rst(config_rst)); 
mux6 mux_1784 (.in({n11103_1, n11102_0, n11095_1, n11094_0, n11039_0, n11038_1/**/}), .out(n3875), .config_in(config_chain[5354:5352]), .config_rst(config_rst)); 
mux6 mux_1785 (.in({n13465_1, n13464_0, n13397_0, n13396_1, n13381_0, n13380_1}), .out(n3876), .config_in(config_chain[5357:5355]), .config_rst(config_rst)); 
mux6 mux_1786 (.in({n10813_0, n10812_0, n10801_0, n10800_0, n10781_1, n10780_1}), .out(n3877), .config_in(config_chain[5360:5358]), .config_rst(config_rst)); 
mux6 mux_1787 (.in({n13185_0, n13184_0, n13177_0/**/, n13176_0, n13125_1, n13124_1}), .out(n3878), .config_in(config_chain[5363:5361]), .config_rst(config_rst)); 
mux6 mux_1788 (.in({n11055_0, n11054_0, n11041_0, n11040_1, n11015_0, n11014_1/**/}), .out(n3879), .config_in(config_chain[5366:5364]), .config_rst(config_rst)); 
mux6 mux_1789 (.in({n13417_0, n13416_0, n13405_0, n13404_1, n13385_0, n13384_1}), .out(n3880), .config_in(config_chain[5369:5367]), .config_rst(config_rst)); 
mux6 mux_1790 (.in({n10841_1, n10840_0, n10833_1, n10832_0, n10783_1, n10782_1}), .out(n3881), .config_in(config_chain[5372:5370]), .config_rst(config_rst)); 
mux6 mux_1791 (.in({n13205_1/**/, n13204_0, n13137_0, n13136_1, n13127_1, n13126_1}), .out(n3882), .config_in(config_chain[5375:5373]), .config_rst(config_rst)); 
mux6 mux_1792 (.in({n11369_1/**/, n11368_0, n11313_0, n11312_0, n11249_0, n11248_1}), .out(n3929), .config_in(config_chain[5378:5376]), .config_rst(config_rst)); 
mux6 mux_1793 (.in({n13487_1, n13486_0, n13431_0, n13430_0, n13417_0, n13416_1}), .out(n3930), .config_in(config_chain[5381:5379]), .config_rst(config_rst)); 
mux6 mux_1794 (.in({n11089_1, n11088_0/**/, n11083_0, n11082_0, n11075_0, n11074_0}), .out(n3931), .config_in(config_chain[5384:5382]), .config_rst(config_rst)); 
mux6 mux_1795 (.in({n13219_1, n13218_0, n13211_1, n13210_0/**/, n13205_0, n13204_0}), .out(n3932), .config_in(config_chain[5387:5385]), .config_rst(config_rst)); 
mux6 mux_1796 (.in({n11333_0, n11332_0, n11321_0, n11320_0, n11281_0, n11280_1}), .out(n3933), .config_in(config_chain[5390:5388]), .config_rst(config_rst)); 
mux6 mux_1797 (.in({n13451_0, n13450_0, n13447_0, n13446_0, n13439_0, n13438_0}), .out(n3934), .config_in(config_chain[5393:5391]), .config_rst(config_rst)); 
mux6 mux_1798 (.in({n11105_1, n11104_0, n10991_0, n10990_1, n10959_0, n10958_1}), .out(n3935), .config_in(config_chain[5396:5394]), .config_rst(config_rst)); 
mux6 mux_1799 (.in({n13227_1, n13226_0, n13171_0, n13170_0, n13159_0, n13158_1}), .out(n3936), .config_in(config_chain[5399:5397]), .config_rst(config_rst)); 
mux6 mux_1800 (.in({n11355_1, n11354_0, n11349_0, n11348_0, n11341_0, n11340_0}), .out(n3937), .config_in(config_chain[5402:5400]), .config_rst(config_rst)); 
mux6 mux_1801 (.in({n13473_1, n13472_0, n13467_0, n13466_0, n13459_0, n13458_0}), .out(n3938), .config_in(config_chain[5405:5403]), .config_rst(config_rst)); 
mux6 mux_1802 (.in({n11057_0, n11056_0, n11049_0, n11048_0, n11023_0, n11022_1}), .out(n3939), .config_in(config_chain[5408:5406]), .config_rst(config_rst)); 
mux6 mux_1803 (.in({n13191_0, n13190_0, n13179_0, n13178_0, n13167_0, n13166_1}), .out(n3940), .config_in(config_chain[5411:5409]), .config_rst(config_rst)); 
mux6 mux_1804 (.in({n11371_1, n11370_0, n11363_1, n11362_0, n11225_0, n11224_1}), .out(n3941), .config_in(config_chain[5414:5412]), .config_rst(config_rst)); 
mux6 mux_1805 (.in({n13489_1, n13488_0, n13419_0, n13418_1, n13411_0, n13410_1}), .out(n3942), .config_in(config_chain[5417:5415]), .config_rst(config_rst)); 
mux6 mux_1806 (.in({n11091_1, n11090_0, n11077_0, n11076_0, n11065_0, n11064_0}), .out(n3943), .config_in(config_chain[5420:5418]), .config_rst(config_rst)); 
mux6 mux_1807 (.in({n13213_1, n13212_0, n13207_0/**/, n13206_0, n13199_0, n13198_0}), .out(n3944), .config_in(config_chain[5423:5421]), .config_rst(config_rst)); 
mux6 mux_1808 (.in({n11323_0, n11322_0, n11315_0, n11314_0, n11289_0, n11288_1/**/}), .out(n3945), .config_in(config_chain[5426:5424]), .config_rst(config_rst)); 
mux6 mux_1809 (.in({n13453_0, n13452_0, n13441_0, n13440_0, n13427_0, n13426_1/**/}), .out(n3946), .config_in(config_chain[5429:5427]), .config_rst(config_rst)); 
mux6 mux_1810 (.in({n11099_1, n11098_0, n11085_0, n11084_0/**/, n10967_0, n10966_1}), .out(n3947), .config_in(config_chain[5432:5430]), .config_rst(config_rst)); 
mux6 mux_1811 (.in({n13229_1/**/, n13228_0, n13221_1, n13220_0, n13153_0, n13152_1}), .out(n3948), .config_in(config_chain[5435:5433]), .config_rst(config_rst)); 
mux6 mux_1812 (.in({n11343_0, n11342_0, n11335_0, n11334_0/**/, n11331_0, n11330_0}), .out(n3949), .config_in(config_chain[5438:5436]), .config_rst(config_rst)); 
mux6 mux_1813 (.in({n13475_1, n13474_0, n13461_0/**/, n13460_0, n13449_0, n13448_0}), .out(n3950), .config_in(config_chain[5441:5439]), .config_rst(config_rst)); 
mux6 mux_1814 (.in({n11051_0, n11050_0, n11031_0, n11030_1, n10999_0, n10998_1}), .out(n3951), .config_in(config_chain[5444:5442]), .config_rst(config_rst)); 
mux6 mux_1815 (.in({n13181_0, n13180_0, n13173_0, n13172_0, n13169_0, n13168_1}), .out(n3952), .config_in(config_chain[5447:5445]), .config_rst(config_rst)); 
mux6 mux_1816 (.in({n11365_1, n11364_0, n11351_0, n11350_0/**/, n11233_0, n11232_1}), .out(n3953), .config_in(config_chain[5450:5448]), .config_rst(config_rst)); 
mux6 mux_1817 (.in({n13491_1, n13490_0, n13483_1, n13482_0, n13413_0, n13412_1}), .out(n3954), .config_in(config_chain[5453:5451]), .config_rst(config_rst)); 
mux6 mux_1818 (.in({n11079_0, n11078_0, n11071_0, n11070_0/**/, n11067_0, n11066_0}), .out(n3955), .config_in(config_chain[5456:5454]), .config_rst(config_rst)); 
mux6 mux_1819 (.in({n13201_0, n13200_0/**/, n13193_0, n13192_0, n13189_0, n13188_0}), .out(n3956), .config_in(config_chain[5459:5457]), .config_rst(config_rst)); 
mux6 mux_1820 (.in({n11373_1, n11372_0, n11317_0, n11316_0, n11265_0, n11264_1}), .out(n3957), .config_in(config_chain[5462:5460]), .config_rst(config_rst)); 
mux6 mux_1821 (.in({n13435_0, n13434_0, n13429_0, n13428_1, n13421_0, n13420_1}), .out(n3958), .config_in(config_chain[5465:5463]), .config_rst(config_rst)); 
mux6 mux_1822 (.in({n11101_1, n11100_0, n11093_1, n11092_0, n11087_0, n11086_0}), .out(n3959), .config_in(config_chain[5468:5466]), .config_rst(config_rst)); 
mux6 mux_1823 (.in({n13223_1, n13222_0, n13209_0, n13208_0, n13155_0, n13154_1}), .out(n3960), .config_in(config_chain[5471:5469]), .config_rst(config_rst)); 
mux6 mux_1824 (.in({n11337_0, n11336_0/**/, n11325_0, n11324_0, n11307_0, n11306_1}), .out(n3961), .config_in(config_chain[5474:5472]), .config_rst(config_rst)); 
mux6 mux_1825 (.in({n13463_0, n13462_0, n13455_0, n13454_0, n13385_0, n13384_1/**/}), .out(n3962), .config_in(config_chain[5477:5475]), .config_rst(config_rst)); 
mux6 mux_1826 (.in({n11053_0, n11052_0, n11045_1, n11044_1, n11007_0, n11006_1/**/}), .out(n3963), .config_in(config_chain[5480:5478]), .config_rst(config_rst)); 
mux6 mux_1827 (.in({n13175_0, n13174_0/**/, n13163_0, n13162_1, n13127_1, n13126_1}), .out(n3964), .config_in(config_chain[5483:5481]), .config_rst(config_rst)); 
mux6 mux_1828 (.in({n11359_1, n11358_0, n11345_0, n11344_0, n11309_0/**/, n11308_1}), .out(n3965), .config_in(config_chain[5486:5484]), .config_rst(config_rst)); 
mux6 mux_1829 (.in({n13485_1/**/, n13484_0, n13477_1, n13476_0, n13387_0, n13386_1}), .out(n3966), .config_in(config_chain[5489:5487]), .config_rst(config_rst)); 
mux6 mux_1830 (.in({n11073_0, n11072_0, n11061_0, n11060_0, n11047_1, n11046_1}), .out(n3967), .config_in(config_chain[5492:5490]), .config_rst(config_rst)); 
mux6 mux_1831 (.in({n13231_1, n13230_0, n13195_0/**/, n13194_0, n13183_0, n13182_0}), .out(n3968), .config_in(config_chain[5495:5493]), .config_rst(config_rst)); 
mux6 mux_1832 (.in({n11311_1/**/, n11310_1, n11273_0, n11272_1, n11241_0, n11240_1}), .out(n3969), .config_in(config_chain[5498:5496]), .config_rst(config_rst)); 
mux6 mux_1833 (.in({n13437_0, n13436_0, n13423_0, n13422_1, n13389_1, n13388_1}), .out(n3970), .config_in(config_chain[5501:5499]), .config_rst(config_rst)); 
mux6 mux_1834 (.in({n11095_1, n11094_0, n11081_0, n11080_0, n11039_0, n11038_1}), .out(n3971), .config_in(config_chain[5504:5502]), .config_rst(config_rst)); 
mux6 mux_1835 (.in({n13225_1, n13224_0, n13217_1, n13216_0, n13121_0, n13120_1}), .out(n3972), .config_in(config_chain[5507:5505]), .config_rst(config_rst)); 
mux6 mux_1836 (.in({n11353_1, n11352_0, n11327_0, n11326_0/**/, n11319_0, n11318_0}), .out(n3973), .config_in(config_chain[5510:5508]), .config_rst(config_rst)); 
mux6 mux_1837 (.in({n13471_1, n13470_0, n13457_0, n13456_0, n13445_0, n13444_0}), .out(n3974), .config_in(config_chain[5513:5511]), .config_rst(config_rst)); 
mux6 mux_1838 (.in({n11103_1, n11102_0, n11041_0, n11040_1, n10983_0, n10982_1}), .out(n3975), .config_in(config_chain[5516:5514]), .config_rst(config_rst)); 
mux6 mux_1839 (.in({n13165_0, n13164_1/**/, n13157_0, n13156_1, n13123_0, n13122_1}), .out(n3976), .config_in(config_chain[5519:5517]), .config_rst(config_rst)); 
mux6 mux_1840 (.in({n11375_1, n11374_0, n11361_1, n11360_0, n11347_0, n11346_0/**/}), .out(n3977), .config_in(config_chain[5522:5520]), .config_rst(config_rst)); 
mux6 mux_1841 (.in({n13479_1, n13478_0, n13465_0, n13464_0/**/, n13383_0, n13382_1}), .out(n3978), .config_in(config_chain[5525:5523]), .config_rst(config_rst)); 
mux6 mux_1842 (.in({n11063_0, n11062_0, n11055_0, n11054_0/**/, n11043_0, n11042_1}), .out(n3979), .config_in(config_chain[5528:5526]), .config_rst(config_rst)); 
mux6 mux_1843 (.in({n13197_0/**/, n13196_0, n13185_0, n13184_0, n13125_0, n13124_1}), .out(n3980), .config_in(config_chain[5531:5529]), .config_rst(config_rst)); 
mux6 mux_1844 (.in({n11621_1, n11620_0, n11605_0, n11604_0, n11591_0, n11590_0}), .out(n4027), .config_in(config_chain[5534:5532]), .config_rst(config_rst)); 
mux6 mux_1845 (.in({n13495_0, n13494_0, n13479_0, n13478_0, n13465_0/**/, n13464_0}), .out(n4028), .config_in(config_chain[5537:5535]), .config_rst(config_rst)); 
mux6 mux_1846 (.in({n11313_0, n11312_0, n11281_0, n11280_1, n11249_0, n11248_1}), .out(n4029), .config_in(config_chain[5540:5538]), .config_rst(config_rst)); 
mux6 mux_1847 (.in({n13199_0, n13198_0, n13191_0, n13190_0, n13185_0, n13184_1}), .out(n4030), .config_in(config_chain[5543:5541]), .config_rst(config_rst)); 
mux6 mux_1848 (.in({n11629_1, n11628_0, n11613_0, n11612_0, n11491_0, n11490_1}), .out(n4031), .config_in(config_chain[5546:5544]), .config_rst(config_rst)); 
mux6 mux_1849 (.in({n13511_0, n13510_0, n13503_0, n13502_0, n13431_0, n13430_1}), .out(n4032), .config_in(config_chain[5549:5547]), .config_rst(config_rst)); 
mux6 mux_1850 (.in({n11341_0, n11340_0, n11333_0, n11332_0, n11329_0, n11328_0}), .out(n4033), .config_in(config_chain[5552:5550]), .config_rst(config_rst)); 
mux6 mux_1851 (.in({n13233_0, n13232_0, n13219_0, n13218_0, n13207_0, n13206_0}), .out(n4034), .config_in(config_chain[5555:5553]), .config_rst(config_rst)); 
mux6 mux_1852 (.in({n11577_0, n11576_0, n11555_0, n11554_1, n11523_0, n11522_1}), .out(n4035), .config_in(config_chain[5558:5556]), .config_rst(config_rst)); 
mux6 mux_1853 (.in({n13451_0, n13450_0, n13447_0, n13446_1, n13439_0, n13438_1}), .out(n4036), .config_in(config_chain[5561:5559]), .config_rst(config_rst)); 
mux6 mux_1854 (.in({n11363_1/**/, n11362_0, n11355_1, n11354_0, n11349_0, n11348_0}), .out(n4037), .config_in(config_chain[5564:5562]), .config_rst(config_rst)); 
mux6 mux_1855 (.in({n13241_0, n13240_0, n13227_0, n13226_0/**/, n13171_0, n13170_1}), .out(n4038), .config_in(config_chain[5567:5565]), .config_rst(config_rst)); 
mux6 mux_1856 (.in({n11599_0, n11598_0/**/, n11593_0, n11592_0, n11585_0, n11584_0}), .out(n4039), .config_in(config_chain[5570:5568]), .config_rst(config_rst)); 
mux6 mux_1857 (.in({n13481_0/**/, n13480_0, n13473_0, n13472_0, n13467_0, n13466_0}), .out(n4040), .config_in(config_chain[5573:5571]), .config_rst(config_rst)); 
mux6 mux_1858 (.in({n11371_1, n11370_0, n11315_0, n11314_0, n11257_0, n11256_1}), .out(n4041), .config_in(config_chain[5576:5574]), .config_rst(config_rst)); 
mux6 mux_1859 (.in({n13193_0, n13192_0, n13187_0/**/, n13186_1, n13179_0, n13178_1}), .out(n4042), .config_in(config_chain[5579:5577]), .config_rst(config_rst)); 
mux6 mux_1860 (.in({n11631_1, n11630_0, n11623_1, n11622_0, n11615_0, n11614_0}), .out(n4043), .config_in(config_chain[5582:5580]), .config_rst(config_rst)); 
mux6 mux_1861 (.in({n13505_0, n13504_0/**/, n13489_0, n13488_0, n13433_0, n13432_1}), .out(n4044), .config_in(config_chain[5585:5583]), .config_rst(config_rst)); 
mux6 mux_1862 (.in({n11335_0, n11334_0/**/, n11323_0, n11322_0, n11289_0, n11288_1}), .out(n4045), .config_in(config_chain[5588:5586]), .config_rst(config_rst)); 
mux6 mux_1863 (.in({n13213_0, n13212_0/**/, n13209_0, n13208_0, n13201_0, n13200_0}), .out(n4046), .config_in(config_chain[5591:5589]), .config_rst(config_rst)); 
mux6 mux_1864 (.in({n11639_1, n11638_0, n11531_0, n11530_1, n11499_0/**/, n11498_1}), .out(n4047), .config_in(config_chain[5594:5592]), .config_rst(config_rst)); 
mux6 mux_1865 (.in({n13513_0, n13512_0, n13453_0, n13452_0, n13441_0, n13440_1}), .out(n4048), .config_in(config_chain[5597:5595]), .config_rst(config_rst)); 
mux6 mux_1866 (.in({n11357_1, n11356_0, n11351_0, n11350_0, n11343_0, n11342_0/**/}), .out(n4049), .config_in(config_chain[5600:5598]), .config_rst(config_rst)); 
mux6 mux_1867 (.in({n13243_0/**/, n13242_0, n13235_0, n13234_0, n13229_0, n13228_0}), .out(n4050), .config_in(config_chain[5603:5601]), .config_rst(config_rst)); 
mux6 mux_1868 (.in({n11601_0, n11600_0, n11587_0/**/, n11586_0, n11563_0, n11562_1}), .out(n4051), .config_in(config_chain[5606:5604]), .config_rst(config_rst)); 
mux6 mux_1869 (.in({n13475_0, n13474_0, n13469_0/**/, n13468_0, n13461_0, n13460_0}), .out(n4052), .config_in(config_chain[5609:5607]), .config_rst(config_rst)); 
mux6 mux_1870 (.in({n11373_1, n11372_0/**/, n11265_0, n11264_1, n11233_0, n11232_1}), .out(n4053), .config_in(config_chain[5612:5610]), .config_rst(config_rst)); 
mux6 mux_1871 (.in({n13251_0, n13250_0, n13181_0, n13180_1, n13173_0, n13172_1}), .out(n4054), .config_in(config_chain[5615:5613]), .config_rst(config_rst)); 
mux6 mux_1872 (.in({n11625_1, n11624_0, n11609_0, n11608_0, n11595_0, n11594_0}), .out(n4055), .config_in(config_chain[5618:5616]), .config_rst(config_rst)); 
mux6 mux_1873 (.in({n13499_0, n13498_0, n13491_0, n13490_0, n13483_0, n13482_0}), .out(n4056), .config_in(config_chain[5621:5619]), .config_rst(config_rst)); 
mux6 mux_1874 (.in({n11325_0, n11324_0, n11317_0/**/, n11316_0, n11297_0, n11296_1}), .out(n4057), .config_in(config_chain[5624:5622]), .config_rst(config_rst)); 
mux6 mux_1875 (.in({n13215_0, n13214_0, n13203_0, n13202_0, n13189_0, n13188_1/**/}), .out(n4058), .config_in(config_chain[5627:5625]), .config_rst(config_rst)); 
mux6 mux_1876 (.in({n11641_1, n11640_0, n11633_1/**/, n11632_0, n11507_0, n11506_1}), .out(n4059), .config_in(config_chain[5630:5628]), .config_rst(config_rst)); 
mux6 mux_1877 (.in({n13515_0, n13514_0, n13443_0, n13442_1, n13435_0, n13434_1}), .out(n4060), .config_in(config_chain[5633:5631]), .config_rst(config_rst)); 
mux6 mux_1878 (.in({n11359_1, n11358_0, n11345_0, n11344_0, n11307_0, n11306_1}), .out(n4061), .config_in(config_chain[5636:5634]), .config_rst(config_rst)); 
mux6 mux_1879 (.in({n13237_0, n13236_0, n13223_0, n13222_0, n13125_0, n13124_2}), .out(n4062), .config_in(config_chain[5639:5637]), .config_rst(config_rst)); 
mux6 mux_1880 (.in({n11581_0, n11580_0, n11571_0/**/, n11570_1, n11539_0, n11538_1}), .out(n4063), .config_in(config_chain[5642:5640]), .config_rst(config_rst)); 
mux6 mux_1881 (.in({n13463_0, n13462_0/**/, n13455_0, n13454_0, n13385_0, n13384_2}), .out(n4064), .config_in(config_chain[5645:5643]), .config_rst(config_rst)); 
mux6 mux_1882 (.in({n11367_1, n11366_0, n11309_0, n11308_1, n11241_0, n11240_1}), .out(n4065), .config_in(config_chain[5648:5646]), .config_rst(config_rst)); 
mux6 mux_1883 (.in({n13245_0, n13244_0/**/, n13175_0, n13174_1, n13129_0, n13128_2}), .out(n4066), .config_in(config_chain[5651:5649]), .config_rst(config_rst)); 
mux6 mux_1884 (.in({n11611_0, n11610_0, n11603_0/**/, n11602_0, n11573_0, n11572_1}), .out(n4067), .config_in(config_chain[5654:5652]), .config_rst(config_rst)); 
mux6 mux_1885 (.in({n13501_0, n13500_0, n13485_0, n13484_0/**/, n13387_0, n13386_2}), .out(n4068), .config_in(config_chain[5657:5655]), .config_rst(config_rst)); 
mux6 mux_1886 (.in({n11353_1, n11352_0, n11319_0/**/, n11318_0, n11273_0, n11272_1}), .out(n4069), .config_in(config_chain[5660:5658]), .config_rst(config_rst)); 
mux6 mux_1887 (.in({n13231_0, n13230_0, n13205_0/**/, n13204_0, n13197_0, n13196_0}), .out(n4070), .config_in(config_chain[5663:5661]), .config_rst(config_rst)); 
mux6 mux_1888 (.in({n11635_1, n11634_0, n11627_1, n11626_0, n11575_0/**/, n11574_1}), .out(n4071), .config_in(config_chain[5666:5664]), .config_rst(config_rst)); 
mux6 mux_1889 (.in({n13509_0/**/, n13508_0, n13437_0, n13436_1, n13389_0, n13388_2}), .out(n4072), .config_in(config_chain[5669:5667]), .config_rst(config_rst)); 
mux6 mux_1890 (.in({n11375_1, n11374_0, n11339_0, n11338_0, n11327_0, n11326_0}), .out(n4073), .config_in(config_chain[5672:5670]), .config_rst(config_rst)); 
mux6 mux_1891 (.in({n13253_0, n13252_0, n13225_0, n13224_0, n13217_0, n13216_0/**/}), .out(n4074), .config_in(config_chain[5675:5673]), .config_rst(config_rst)); 
mux6 mux_1892 (.in({n11597_1, n11596_0, n11583_0, n11582_0, n11547_0, n11546_1}), .out(n4075), .config_in(config_chain[5678:5676]), .config_rst(config_rst)); 
mux6 mux_1893 (.in({n13493_0, n13492_0, n13457_0, n13456_0, n13445_0, n13444_1}), .out(n4076), .config_in(config_chain[5681:5679]), .config_rst(config_rst)); 
mux6 mux_1894 (.in({n11369_1, n11368_0, n11361_1, n11360_0, n11305_0, n11304_1}), .out(n4077), .config_in(config_chain[5684:5682]), .config_rst(config_rst)); 
mux6 mux_1895 (.in({n13247_0, n13246_0/**/, n13177_0, n13176_1, n13123_0, n13122_2}), .out(n4078), .config_in(config_chain[5687:5685]), .config_rst(config_rst)); 
mux6 mux_1896 (.in({n11899_1, n11898_0, n11841_0, n11840_0, n11773_0, n11772_1}), .out(n4125), .config_in(config_chain[5690:5688]), .config_rst(config_rst)); 
mux6 mux_1897 (.in({n13531_0, n13530_0, n13473_0, n13472_0, n13457_0, n13456_1}), .out(n4126), .config_in(config_chain[5693:5691]), .config_rst(config_rst)); 
mux6 mux_1898 (.in({n11621_1, n11620_0, n11613_0, n11612_0/**/, n11605_0, n11604_0}), .out(n4127), .config_in(config_chain[5696:5694]), .config_rst(config_rst)); 
mux6 mux_1899 (.in({n13263_0, n13262_0, n13255_0, n13254_0, n13247_0, n13246_0}), .out(n4128), .config_in(config_chain[5699:5697]), .config_rst(config_rst)); 
mux6 mux_1900 (.in({n11863_0, n11862_0/**/, n11849_0, n11848_0, n11805_0, n11804_1}), .out(n4129), .config_in(config_chain[5702:5700]), .config_rst(config_rst)); 
mux6 mux_1901 (.in({n13495_0, n13494_0, n13489_0, n13488_0, n13481_0, n13480_0}), .out(n4130), .config_in(config_chain[5705:5703]), .config_rst(config_rst)); 
mux6 mux_1902 (.in({n11637_1/**/, n11636_0, n11523_0, n11522_1, n11491_0, n11490_1}), .out(n4131), .config_in(config_chain[5708:5706]), .config_rst(config_rst)); 
mux6 mux_1903 (.in({n13271_0/**/, n13270_0, n13211_0, n13210_0, n13199_0, n13198_1}), .out(n4132), .config_in(config_chain[5711:5709]), .config_rst(config_rst)); 
mux6 mux_1904 (.in({n11885_1, n11884_0, n11879_0, n11878_0, n11871_0, n11870_0}), .out(n4133), .config_in(config_chain[5714:5712]), .config_rst(config_rst)); 
mux6 mux_1905 (.in({n13517_0, n13516_0, n13511_0, n13510_0, n13503_0, n13502_0}), .out(n4134), .config_in(config_chain[5717:5715]), .config_rst(config_rst)); 
mux6 mux_1906 (.in({n11585_0, n11584_0, n11577_0, n11576_0, n11555_0, n11554_1}), .out(n4135), .config_in(config_chain[5720:5718]), .config_rst(config_rst)); 
mux6 mux_1907 (.in({n13233_0, n13232_0, n13219_0, n13218_0, n13207_0, n13206_1}), .out(n4136), .config_in(config_chain[5723:5721]), .config_rst(config_rst)); 
mux6 mux_1908 (.in({n11901_1, n11900_0, n11893_1, n11892_0, n11749_0, n11748_1/**/}), .out(n4137), .config_in(config_chain[5726:5724]), .config_rst(config_rst)); 
mux6 mux_1909 (.in({n13533_0, n13532_0, n13459_0, n13458_1, n13451_0/**/, n13450_1}), .out(n4138), .config_in(config_chain[5729:5727]), .config_rst(config_rst)); 
mux6 mux_1910 (.in({n11623_1, n11622_0, n11607_0, n11606_0/**/, n11593_0, n11592_0}), .out(n4139), .config_in(config_chain[5732:5730]), .config_rst(config_rst)); 
mux6 mux_1911 (.in({n13257_0, n13256_0/**/, n13249_0, n13248_0, n13241_0, n13240_0}), .out(n4140), .config_in(config_chain[5735:5733]), .config_rst(config_rst)); 
mux6 mux_1912 (.in({n11851_0, n11850_0, n11843_0, n11842_0, n11813_0, n11812_1/**/}), .out(n4141), .config_in(config_chain[5738:5736]), .config_rst(config_rst)); 
mux6 mux_1913 (.in({n13497_0, n13496_0, n13483_0, n13482_0, n13467_0, n13466_1}), .out(n4142), .config_in(config_chain[5741:5739]), .config_rst(config_rst)); 
mux6 mux_1914 (.in({n11631_1, n11630_0, n11615_0/**/, n11614_0, n11499_0, n11498_1}), .out(n4143), .config_in(config_chain[5744:5742]), .config_rst(config_rst)); 
mux6 mux_1915 (.in({n13273_0, n13272_0/**/, n13265_0, n13264_0, n13193_0, n13192_1}), .out(n4144), .config_in(config_chain[5747:5745]), .config_rst(config_rst)); 
mux6 mux_1916 (.in({n11873_0, n11872_0, n11865_0, n11864_0, n11859_0, n11858_0}), .out(n4145), .config_in(config_chain[5750:5748]), .config_rst(config_rst)); 
mux6 mux_1917 (.in({n13519_0, n13518_0, n13505_0, n13504_0, n13491_0, n13490_0}), .out(n4146), .config_in(config_chain[5753:5751]), .config_rst(config_rst)); 
mux6 mux_1918 (.in({n11579_0, n11578_0, n11563_0, n11562_1, n11531_0, n11530_1/**/}), .out(n4147), .config_in(config_chain[5756:5754]), .config_rst(config_rst)); 
mux6 mux_1919 (.in({n13221_0, n13220_0, n13213_0, n13212_0, n13209_0/**/, n13208_1}), .out(n4148), .config_in(config_chain[5759:5757]), .config_rst(config_rst)); 
mux6 mux_1920 (.in({n11895_1, n11894_0, n11881_0, n11880_0, n11757_0, n11756_1}), .out(n4149), .config_in(config_chain[5762:5760]), .config_rst(config_rst)); 
mux6 mux_1921 (.in({n13535_0, n13534_0/**/, n13527_0, n13526_0, n13453_0, n13452_1}), .out(n4150), .config_in(config_chain[5765:5763]), .config_rst(config_rst)); 
mux6 mux_1922 (.in({n11609_0, n11608_0, n11601_0, n11600_0, n11595_0, n11594_0}), .out(n4151), .config_in(config_chain[5768:5766]), .config_rst(config_rst)); 
mux6 mux_1923 (.in({n13243_0, n13242_0, n13235_0, n13234_0, n13229_0, n13228_0}), .out(n4152), .config_in(config_chain[5771:5769]), .config_rst(config_rst)); 
mux6 mux_1924 (.in({n11903_1, n11902_0, n11845_0, n11844_0, n11789_0, n11788_1}), .out(n4153), .config_in(config_chain[5774:5772]), .config_rst(config_rst)); 
mux6 mux_1925 (.in({n13477_0, n13476_0, n13469_0, n13468_1, n13461_0, n13460_1}), .out(n4154), .config_in(config_chain[5777:5775]), .config_rst(config_rst)); 
mux6 mux_1926 (.in({n11633_1, n11632_0, n11625_1, n11624_0/**/, n11617_0, n11616_0}), .out(n4155), .config_in(config_chain[5780:5778]), .config_rst(config_rst)); 
mux6 mux_1927 (.in({n13267_0, n13266_0, n13251_0, n13250_0, n13195_0, n13194_1/**/}), .out(n4156), .config_in(config_chain[5783:5781]), .config_rst(config_rst)); 
mux6 mux_1928 (.in({n11867_0, n11866_0, n11861_1, n11860_0, n11853_0, n11852_0}), .out(n4157), .config_in(config_chain[5786:5784]), .config_rst(config_rst)); 
mux6 mux_1929 (.in({n13507_0, n13506_0/**/, n13499_0, n13498_0, n13493_0, n13492_0}), .out(n4158), .config_in(config_chain[5789:5787]), .config_rst(config_rst)); 
mux6 mux_1930 (.in({n11641_1, n11640_0, n11581_0, n11580_0, n11539_0, n11538_1}), .out(n4159), .config_in(config_chain[5792:5790]), .config_rst(config_rst)); 
mux6 mux_1931 (.in({n13275_0, n13274_0, n13215_0, n13214_0, n13203_0/**/, n13202_1}), .out(n4160), .config_in(config_chain[5795:5793]), .config_rst(config_rst)); 
mux6 mux_1932 (.in({n11889_1, n11888_0, n11883_1, n11882_0, n11875_0, n11874_0/**/}), .out(n4161), .config_in(config_chain[5798:5796]), .config_rst(config_rst)); 
mux6 mux_1933 (.in({n13529_0, n13528_0, n13521_0/**/, n13520_0, n13515_0, n13514_0}), .out(n4162), .config_in(config_chain[5801:5799]), .config_rst(config_rst)); 
mux6 mux_1934 (.in({n11603_0, n11602_0, n11589_0/**/, n11588_0, n11571_0, n11570_1}), .out(n4163), .config_in(config_chain[5804:5802]), .config_rst(config_rst)); 
mux6 mux_1935 (.in({n13237_0, n13236_0, n13223_0, n13222_0, n13127_0/**/, n13126_2}), .out(n4164), .config_in(config_chain[5807:5805]), .config_rst(config_rst)); 
mux6 mux_1936 (.in({n11905_1, n11904_0/**/, n11797_0, n11796_1, n11765_0, n11764_1}), .out(n4165), .config_in(config_chain[5810:5808]), .config_rst(config_rst)); 
mux6 mux_1937 (.in({n13537_0, n13536_0, n13479_0, n13478_0, n13463_0, n13462_1}), .out(n4166), .config_in(config_chain[5813:5811]), .config_rst(config_rst)); 
mux6 mux_1938 (.in({n11627_1, n11626_0, n11611_0, n11610_0, n11575_0/**/, n11574_1}), .out(n4167), .config_in(config_chain[5816:5814]), .config_rst(config_rst)); 
mux6 mux_1939 (.in({n13269_0, n13268_0/**/, n13261_0, n13260_0, n13129_0, n13128_2}), .out(n4168), .config_in(config_chain[5819:5817]), .config_rst(config_rst)); 
mux6 mux_1940 (.in({n11855_0, n11854_0, n11847_0, n11846_0/**/, n11837_0, n11836_1}), .out(n4169), .config_in(config_chain[5822:5820]), .config_rst(config_rst)); 
mux6 mux_1941 (.in({n13501_0, n13500_0, n13487_0, n13486_0/**/, n13387_0, n13386_2}), .out(n4170), .config_in(config_chain[5825:5823]), .config_rst(config_rst)); 
mux6 mux_1942 (.in({n11635_1/**/, n11634_0, n11597_1, n11596_0, n11515_0, n11514_1}), .out(n4171), .config_in(config_chain[5828:5826]), .config_rst(config_rst)); 
mux6 mux_1943 (.in({n13231_0, n13230_0, n13205_0, n13204_1, n13197_0, n13196_1}), .out(n4172), .config_in(config_chain[5831:5829]), .config_rst(config_rst)); 
mux6 mux_1944 (.in({n11891_1, n11890_0, n11877_0, n11876_0, n11839_0, n11838_1}), .out(n4173), .config_in(config_chain[5834:5832]), .config_rst(config_rst)); 
mux6 mux_1945 (.in({n13523_0, n13522_0, n13509_0, n13508_0, n13471_0, n13470_1}), .out(n4174), .config_in(config_chain[5837:5835]), .config_rst(config_rst)); 
mux6 mux_1946 (.in({n11619_1, n11618_0, n11591_0, n11590_0, n11583_0, n11582_0}), .out(n4175), .config_in(config_chain[5840:5838]), .config_rst(config_rst)); 
mux6 mux_1947 (.in({n13253_0, n13252_0, n13239_0, n13238_0, n13225_0, n13224_0/**/}), .out(n4176), .config_in(config_chain[5843:5841]), .config_rst(config_rst)); 
mux6 mux_1948 (.in({n12147_1, n12146_0, n12131_0, n12130_0, n12117_0, n12116_0}), .out(n4223), .config_in(config_chain[5846:5844]), .config_rst(config_rst)); 
mux6 mux_1949 (.in({n13539_0, n13538_0, n13523_0, n13522_0, n13509_0, n13508_0}), .out(n4224), .config_in(config_chain[5849:5847]), .config_rst(config_rst)); 
mux6 mux_1950 (.in({n11841_0, n11840_0, n11805_0, n11804_1, n11773_0, n11772_1/**/}), .out(n4225), .config_in(config_chain[5852:5850]), .config_rst(config_rst)); 
mux6 mux_1951 (.in({n13241_0, n13240_0, n13233_0, n13232_0, n13225_0, n13224_1}), .out(n4226), .config_in(config_chain[5855:5853]), .config_rst(config_rst)); 
mux6 mux_1952 (.in({n12155_1, n12154_0, n12139_0, n12138_0, n12013_0, n12012_1}), .out(n4227), .config_in(config_chain[5858:5856]), .config_rst(config_rst)); 
mux6 mux_1953 (.in({n13555_0, n13554_0, n13547_0, n13546_0, n13473_0, n13472_1}), .out(n4228), .config_in(config_chain[5861:5859]), .config_rst(config_rst)); 
mux6 mux_1954 (.in({n11871_0, n11870_0, n11863_0, n11862_0, n11857_0, n11856_0}), .out(n4229), .config_in(config_chain[5864:5862]), .config_rst(config_rst)); 
mux6 mux_1955 (.in({n13277_0, n13276_0, n13263_0, n13262_0, n13249_0, n13248_0}), .out(n4230), .config_in(config_chain[5867:5865]), .config_rst(config_rst)); 
mux6 mux_1956 (.in({n12103_0, n12102_0, n12077_0/**/, n12076_1, n12045_0, n12044_1}), .out(n4231), .config_in(config_chain[5870:5868]), .config_rst(config_rst)); 
mux6 mux_1957 (.in({n13495_0, n13494_0, n13489_0, n13488_1, n13481_0, n13480_1}), .out(n4232), .config_in(config_chain[5873:5871]), .config_rst(config_rst)); 
mux6 mux_1958 (.in({n11893_1/**/, n11892_0, n11885_1, n11884_0, n11879_0, n11878_0}), .out(n4233), .config_in(config_chain[5876:5874]), .config_rst(config_rst)); 
mux6 mux_1959 (.in({n13285_0, n13284_0, n13271_0, n13270_0, n13211_0, n13210_1}), .out(n4234), .config_in(config_chain[5879:5877]), .config_rst(config_rst)); 
mux6 mux_1960 (.in({n12125_0, n12124_0, n12119_0, n12118_0, n12111_0, n12110_0}), .out(n4235), .config_in(config_chain[5882:5880]), .config_rst(config_rst)); 
mux6 mux_1961 (.in({n13525_0/**/, n13524_0, n13517_0, n13516_0, n13511_0, n13510_0}), .out(n4236), .config_in(config_chain[5885:5883]), .config_rst(config_rst)); 
mux6 mux_1962 (.in({n11901_1, n11900_0, n11843_0, n11842_0/**/, n11781_0, n11780_1}), .out(n4237), .config_in(config_chain[5888:5886]), .config_rst(config_rst)); 
mux6 mux_1963 (.in({n13235_0, n13234_0/**/, n13227_0, n13226_1, n13219_0, n13218_1}), .out(n4238), .config_in(config_chain[5891:5889]), .config_rst(config_rst)); 
mux6 mux_1964 (.in({n12157_1, n12156_0, n12149_1, n12148_0, n12141_0, n12140_0}), .out(n4239), .config_in(config_chain[5894:5892]), .config_rst(config_rst)); 
mux6 mux_1965 (.in({n13549_0, n13548_0/**/, n13533_0, n13532_0, n13475_0, n13474_1}), .out(n4240), .config_in(config_chain[5897:5895]), .config_rst(config_rst)); 
mux6 mux_1966 (.in({n11865_0, n11864_0, n11851_0, n11850_0, n11813_0, n11812_1}), .out(n4241), .config_in(config_chain[5900:5898]), .config_rst(config_rst)); 
mux6 mux_1967 (.in({n13257_0, n13256_0, n13251_0, n13250_0, n13243_0, n13242_0}), .out(n4242), .config_in(config_chain[5903:5901]), .config_rst(config_rst)); 
mux6 mux_1968 (.in({n12165_1, n12164_0, n12053_0, n12052_1, n12021_0, n12020_1}), .out(n4243), .config_in(config_chain[5906:5904]), .config_rst(config_rst)); 
mux6 mux_1969 (.in({n13557_0, n13556_0, n13497_0, n13496_0, n13483_0, n13482_1}), .out(n4244), .config_in(config_chain[5909:5907]), .config_rst(config_rst)); 
mux6 mux_1970 (.in({n11887_1, n11886_0, n11881_0, n11880_0/**/, n11873_0, n11872_0}), .out(n4245), .config_in(config_chain[5912:5910]), .config_rst(config_rst)); 
mux6 mux_1971 (.in({n13287_0, n13286_0, n13279_0/**/, n13278_0, n13273_0, n13272_0}), .out(n4246), .config_in(config_chain[5915:5913]), .config_rst(config_rst)); 
mux6 mux_1972 (.in({n12127_0, n12126_0, n12113_0/**/, n12112_0, n12085_0, n12084_1}), .out(n4247), .config_in(config_chain[5918:5916]), .config_rst(config_rst)); 
mux6 mux_1973 (.in({n13519_0, n13518_0/**/, n13513_0, n13512_0, n13505_0, n13504_0}), .out(n4248), .config_in(config_chain[5921:5919]), .config_rst(config_rst)); 
mux6 mux_1974 (.in({n11903_1, n11902_0, n11789_0/**/, n11788_1, n11757_0, n11756_1}), .out(n4249), .config_in(config_chain[5924:5922]), .config_rst(config_rst)); 
mux6 mux_1975 (.in({n13295_0, n13294_0, n13221_0, n13220_1, n13213_0/**/, n13212_1}), .out(n4250), .config_in(config_chain[5927:5925]), .config_rst(config_rst)); 
mux6 mux_1976 (.in({n12151_1, n12150_0, n12135_0, n12134_0, n12121_0, n12120_0}), .out(n4251), .config_in(config_chain[5930:5928]), .config_rst(config_rst)); 
mux6 mux_1977 (.in({n13543_0, n13542_0, n13535_0, n13534_0, n13527_0, n13526_0/**/}), .out(n4252), .config_in(config_chain[5933:5931]), .config_rst(config_rst)); 
mux6 mux_1978 (.in({n11853_0, n11852_0, n11845_0, n11844_0, n11821_0/**/, n11820_1}), .out(n4253), .config_in(config_chain[5936:5934]), .config_rst(config_rst)); 
mux6 mux_1979 (.in({n13259_0, n13258_0, n13245_0, n13244_0, n13229_0, n13228_1}), .out(n4254), .config_in(config_chain[5939:5937]), .config_rst(config_rst)); 
mux6 mux_1980 (.in({n12159_1, n12158_0, n12091_1, n12090_1, n12029_0/**/, n12028_1}), .out(n4255), .config_in(config_chain[5942:5940]), .config_rst(config_rst)); 
mux6 mux_1981 (.in({n13485_0, n13484_1, n13477_0, n13476_1, n13471_0, n13470_1}), .out(n4256), .config_in(config_chain[5945:5943]), .config_rst(config_rst)); 
mux6 mux_1982 (.in({n11889_1, n11888_0, n11875_0, n11874_0, n11861_1, n11860_0}), .out(n4257), .config_in(config_chain[5948:5946]), .config_rst(config_rst)); 
mux6 mux_1983 (.in({n13281_0, n13280_0/**/, n13267_0, n13266_0, n13253_0, n13252_0}), .out(n4258), .config_in(config_chain[5951:5949]), .config_rst(config_rst)); 
mux6 mux_1984 (.in({n12107_0, n12106_0, n12093_1, n12092_1, n12061_0/**/, n12060_1}), .out(n4259), .config_in(config_chain[5954:5952]), .config_rst(config_rst)); 
mux6 mux_1985 (.in({n13507_0, n13506_0, n13499_0, n13498_0, n13493_0, n13492_1/**/}), .out(n4260), .config_in(config_chain[5957:5955]), .config_rst(config_rst)); 
mux6 mux_1986 (.in({n11897_1/**/, n11896_0, n11883_1, n11882_0, n11765_0, n11764_1}), .out(n4261), .config_in(config_chain[5960:5958]), .config_rst(config_rst)); 
mux6 mux_1987 (.in({n13297_0, n13296_0/**/, n13289_0, n13288_0, n13215_0, n13214_1}), .out(n4262), .config_in(config_chain[5963:5961]), .config_rst(config_rst)); 
mux6 mux_1988 (.in({n12137_0, n12136_0, n12129_0, n12128_0, n12123_1, n12122_0}), .out(n4263), .config_in(config_chain[5966:5964]), .config_rst(config_rst)); 
mux6 mux_1989 (.in({n13545_0, n13544_0, n13529_0, n13528_0/**/, n13515_0, n13514_0}), .out(n4264), .config_in(config_chain[5969:5967]), .config_rst(config_rst)); 
mux6 mux_1990 (.in({n11847_0, n11846_0, n11837_0, n11836_1, n11797_0, n11796_1/**/}), .out(n4265), .config_in(config_chain[5972:5970]), .config_rst(config_rst)); 
mux6 mux_1991 (.in({n13247_0, n13246_0, n13239_0, n13238_0, n13127_0, n13126_2}), .out(n4266), .config_in(config_chain[5975:5973]), .config_rst(config_rst)); 
mux6 mux_1992 (.in({n12161_1, n12160_0, n12153_1, n12152_0, n12145_1, n12144_0}), .out(n4267), .config_in(config_chain[5978:5976]), .config_rst(config_rst)); 
mux6 mux_1993 (.in({n13553_0, n13552_0, n13537_0, n13536_0, n13479_0, n13478_1}), .out(n4268), .config_in(config_chain[5981:5979]), .config_rst(config_rst)); 
mux6 mux_1994 (.in({n11869_0, n11868_0, n11855_0, n11854_0, n11839_0, n11838_1}), .out(n4269), .config_in(config_chain[5984:5982]), .config_rst(config_rst)); 
mux6 mux_1995 (.in({n13269_0, n13268_0, n13261_0, n13260_0/**/, n13129_0, n13128_2}), .out(n4270), .config_in(config_chain[5987:5985]), .config_rst(config_rst)); 
mux6 mux_1996 (.in({n12167_1, n12166_0, n12109_0, n12108_0, n12069_0, n12068_1}), .out(n4271), .config_in(config_chain[5990:5988]), .config_rst(config_rst)); 
mux6 mux_1997 (.in({n13501_0, n13500_0, n13487_0, n13486_1, n13389_0, n13388_2}), .out(n4272), .config_in(config_chain[5993:5991]), .config_rst(config_rst)); 
mux6 mux_1998 (.in({n11899_1, n11898_0, n11891_1, n11890_0, n11829_1, n11828_1}), .out(n4273), .config_in(config_chain[5996:5994]), .config_rst(config_rst)); 
mux6 mux_1999 (.in({n13291_0, n13290_0, n13231_0, n13230_1, n13217_0, n13216_1/**/}), .out(n4274), .config_in(config_chain[5999:5997]), .config_rst(config_rst)); 
mux6 mux_2000 (.in({n12155_1, n12154_0, n12147_1, n12146_0, n12139_0, n12138_0}), .out(n4320), .config_in(config_chain[6002:6000]), .config_rst(config_rst)); 
mux6 mux_2001 (.in({n12111_0, n12110_0, n12103_0, n12102_0, n12077_0, n12076_1}), .out(n4323), .config_in(config_chain[6005:6003]), .config_rst(config_rst)); 
mux6 mux_2002 (.in({n12157_1, n12156_0, n12149_1, n12148_0, n12141_0, n12140_0}), .out(n4326), .config_in(config_chain[6008:6006]), .config_rst(config_rst)); 
mux6 mux_2003 (.in({n12113_0, n12112_0, n12105_0, n12104_0, n12085_0, n12084_1}), .out(n4329), .config_in(config_chain[6011:6009]), .config_rst(config_rst)); 
mux6 mux_2004 (.in({n12151_1, n12150_0, n12143_0, n12142_0, n12135_0, n12134_0}), .out(n4332), .config_in(config_chain[6014:6012]), .config_rst(config_rst)); 
mux6 mux_2005 (.in({n12107_0, n12106_0, n12093_1, n12092_1, n12061_0, n12060_1}), .out(n4335), .config_in(config_chain[6017:6015]), .config_rst(config_rst)); 
mux6 mux_2006 (.in({n12153_1, n12152_0, n12145_1, n12144_0, n12137_0, n12136_0}), .out(n4338), .config_in(config_chain[6020:6018]), .config_rst(config_rst)); 
mux6 mux_2007 (.in({n12109_0, n12108_0, n12101_0, n12100_1, n12069_0, n12068_1}), .out(n4341), .config_in(config_chain[6023:6021]), .config_rst(config_rst)); 
mux6 mux_2008 (.in({n9819_1, n9818_0, n9805_0, n9804_0, n9793_0, n9792_0}), .out(n4368), .config_in(config_chain[6026:6024]), .config_rst(config_rst)); 
mux6 mux_2009 (.in({n9835_1, n9834_0, n9767_0, n9766_1, n9759_0, n9758_1}), .out(n4371), .config_in(config_chain[6029:6027]), .config_rst(config_rst)); 
mux6 mux_2010 (.in({n9807_0, n9806_0, n9799_0, n9798_0, n9795_0, n9794_0}), .out(n4374), .config_in(config_chain[6032:6030]), .config_rst(config_rst)); 
mux6 mux_2011 (.in({n9837_1, n9836_0, n9769_0, n9768_1, n9761_0, n9760_1}), .out(n4377), .config_in(config_chain[6035:6033]), .config_rst(config_rst)); 
mux6 mux_2012 (.in({n9809_0, n9808_0, n9801_0, n9800_0, n9797_0, n9796_0}), .out(n4380), .config_in(config_chain[6038:6036]), .config_rst(config_rst)); 
mux6 mux_2013 (.in({n9831_1, n9830_0, n9763_0, n9762_1, n9751_1, n9750_1}), .out(n4383), .config_in(config_chain[6041:6039]), .config_rst(config_rst)); 
mux6 mux_2014 (.in({n9803_0, n9802_0, n9791_0, n9790_0, n9755_1, n9754_1}), .out(n4386), .config_in(config_chain[6044:6042]), .config_rst(config_rst)); 
mux6 mux_2015 (.in({n9833_1, n9832_0, n9765_0, n9764_1, n9747_1, n9746_1}), .out(n4389), .config_in(config_chain[6047:6045]), .config_rst(config_rst)); 
mux6 mux_2016 (.in({n10087_1, n10086_0, n10033_0, n10032_0, n10019_0, n10018_1}), .out(n4417), .config_in(config_chain[6050:6048]), .config_rst(config_rst)); 
mux6 mux_2017 (.in({n13619_1, n13618_0, n13589_0, n13588_0, n13567_0, n13566_0}), .out(n4418), .config_in(config_chain[6053:6051]), .config_rst(config_rst)); 
mux6 mux_2018 (.in({n9819_1, n9818_0, n9813_0, n9812_0, n9805_0, n9804_0}), .out(n4419), .config_in(config_chain[6056:6054]), .config_rst(config_rst)); 
mux6 mux_2019 (.in({n13361_0, n13360_0, n13331_1, n13330_0, n13299_1, n13298_0}), .out(n4420), .config_in(config_chain[6059:6057]), .config_rst(config_rst)); 
mux6 mux_2020 (.in({n10053_0, n10052_0, n10041_0, n10040_0, n10027_0, n10026_1}), .out(n4421), .config_in(config_chain[6062:6060]), .config_rst(config_rst)); 
mux6 mux_2021 (.in({n13631_0, n13630_0, n13599_0, n13598_0, n13561_0, n13560_0}), .out(n4422), .config_in(config_chain[6065:6063]), .config_rst(config_rst)); 
mux6 mux_2022 (.in({n9835_1, n9834_0, n9767_0, n9766_1, n9759_0, n9758_1}), .out(n4423), .config_in(config_chain[6068:6066]), .config_rst(config_rst)); 
mux6 mux_2023 (.in({n13363_1, n13362_0, n13333_0, n13332_0, n13303_0, n13302_0}), .out(n4424), .config_in(config_chain[6071:6069]), .config_rst(config_rst)); 
mux6 mux_2024 (.in({n10073_1, n10072_0, n10069_0, n10068_0, n10061_0, n10060_0}), .out(n4425), .config_in(config_chain[6074:6072]), .config_rst(config_rst)); 
mux6 mux_2025 (.in({n13625_0, n13624_0, n13593_0, n13592_0, n13563_1, n13562_0}), .out(n4426), .config_in(config_chain[6077:6075]), .config_rst(config_rst)); 
mux6 mux_2026 (.in({n9787_0, n9786_0, n9779_0, n9778_0, n9775_0, n9774_1}), .out(n4427), .config_in(config_chain[6080:6078]), .config_rst(config_rst)); 
mux6 mux_2027 (.in({n13365_0, n13364_0, n13335_0, n13334_0, n13305_0, n13304_0}), .out(n4428), .config_in(config_chain[6083:6081]), .config_rst(config_rst)); 
mux6 mux_2028 (.in({n10089_1, n10088_0, n10081_1, n10080_0, n10013_0/**/, n10012_1}), .out(n4429), .config_in(config_chain[6086:6084]), .config_rst(config_rst)); 
mux6 mux_2029 (.in({n13627_1, n13626_0, n13597_0/**/, n13596_0, n13565_0, n13564_0}), .out(n4430), .config_in(config_chain[6089:6087]), .config_rst(config_rst)); 
mux6 mux_2030 (.in({n9821_1, n9820_0, n9807_0, n9806_0, n9795_0, n9794_0}), .out(n4431), .config_in(config_chain[6092:6090]), .config_rst(config_rst)); 
mux6 mux_2031 (.in({n13369_0, n13368_0, n13337_0, n13336_0, n13307_1, n13306_0}), .out(n4432), .config_in(config_chain[6095:6093]), .config_rst(config_rst)); 
mux6 mux_2032 (.in({n10043_0/**/, n10042_0, n10035_0, n10034_0, n10029_0, n10028_1}), .out(n4433), .config_in(config_chain[6098:6096]), .config_rst(config_rst)); 
mux6 mux_2033 (.in({n13629_0, n13628_0, n13607_0, n13606_0, n13569_0, n13568_0}), .out(n4434), .config_in(config_chain[6101:6099]), .config_rst(config_rst)); 
mux6 mux_2034 (.in({n9829_1, n9828_0, n9815_0, n9814_0, n9761_0, n9760_1}), .out(n4435), .config_in(config_chain[6104:6102]), .config_rst(config_rst)); 
mux6 mux_2035 (.in({n13371_1, n13370_0, n13339_1, n13338_0, n13309_0/**/, n13308_0}), .out(n4436), .config_in(config_chain[6107:6105]), .config_rst(config_rst)); 
mux6 mux_2036 (.in({n10063_0, n10062_0, n10055_0, n10054_0/**/, n10051_0, n10050_0}), .out(n4437), .config_in(config_chain[6110:6108]), .config_rst(config_rst)); 
mux6 mux_2037 (.in({n13639_0, n13638_0, n13601_0, n13600_0, n13571_1, n13570_0}), .out(n4438), .config_in(config_chain[6113:6111]), .config_rst(config_rst)); 
mux6 mux_2038 (.in({n9781_0, n9780_0, n9777_0/**/, n9776_1, n9769_0, n9768_1}), .out(n4439), .config_in(config_chain[6116:6114]), .config_rst(config_rst)); 
mux6 mux_2039 (.in({n13373_0, n13372_0, n13343_0, n13342_0, n13311_0, n13310_0}), .out(n4440), .config_in(config_chain[6119:6117]), .config_rst(config_rst)); 
mux6 mux_2040 (.in({n10083_1, n10082_0, n10071_0, n10070_0/**/, n10015_0, n10014_1}), .out(n4441), .config_in(config_chain[6122:6120]), .config_rst(config_rst)); 
mux6 mux_2041 (.in({n13635_1, n13634_0, n13603_1, n13602_0, n13573_0, n13572_0/**/}), .out(n4442), .config_in(config_chain[6125:6123]), .config_rst(config_rst)); 
mux6 mux_2042 (.in({n9809_0, n9808_0, n9801_0, n9800_0, n9797_0, n9796_0/**/}), .out(n4443), .config_in(config_chain[6128:6126]), .config_rst(config_rst)); 
mux6 mux_2043 (.in({n13375_0, n13374_0, n13345_0, n13344_0, n13313_0, n13312_0}), .out(n4444), .config_in(config_chain[6131:6129]), .config_rst(config_rst)); 
mux6 mux_2044 (.in({n10091_1, n10090_0/**/, n10037_0, n10036_0, n10023_0, n10022_1}), .out(n4445), .config_in(config_chain[6134:6132]), .config_rst(config_rst)); 
mux6 mux_2045 (.in({n13637_0, n13636_0, n13605_0, n13604_0/**/, n13583_0, n13582_0}), .out(n4446), .config_in(config_chain[6137:6135]), .config_rst(config_rst)); 
mux6 mux_2046 (.in({n9831_1/**/, n9830_0, n9823_1, n9822_0, n9817_0, n9816_0}), .out(n4447), .config_in(config_chain[6140:6138]), .config_rst(config_rst)); 
mux6 mux_2047 (.in({n13377_0, n13376_0, n13347_1, n13346_0, n13317_0, n13316_0/**/}), .out(n4448), .config_in(config_chain[6143:6141]), .config_rst(config_rst)); 
mux6 mux_2048 (.in({n10057_0, n10056_0, n10045_0, n10044_0, n10003_1, n10002_1}), .out(n4449), .config_in(config_chain[6146:6144]), .config_rst(config_rst)); 
mux6 mux_2049 (.in({n13643_1, n13642_0, n13609_0, n13608_0, n13577_0, n13576_0}), .out(n4450), .config_in(config_chain[6149:6147]), .config_rst(config_rst)); 
mux6 mux_2050 (.in({n9783_0, n9782_0, n9771_0/**/, n9770_1, n9751_1, n9750_1}), .out(n4451), .config_in(config_chain[6152:6150]), .config_rst(config_rst)); 
mux6 mux_2051 (.in({n13383_1, n13382_0, n13349_0, n13348_0, n13319_0, n13318_0}), .out(n4452), .config_in(config_chain[6155:6153]), .config_rst(config_rst)); 
mux6 mux_2052 (.in({n10077_1, n10076_0, n10065_0, n10064_0, n10005_1, n10004_1}), .out(n4453), .config_in(config_chain[6158:6156]), .config_rst(config_rst)); 
mux6 mux_2053 (.in({n13645_1, n13644_0, n13611_1, n13610_0, n13579_1, n13578_0}), .out(n4454), .config_in(config_chain[6161:6159]), .config_rst(config_rst)); 
mux6 mux_2054 (.in({n9803_0, n9802_0, n9791_0, n9790_0, n9753_1, n9752_1}), .out(n4455), .config_in(config_chain[6164:6162]), .config_rst(config_rst)); 
mux6 mux_2055 (.in({n13387_2, n13386_0, n13351_0, n13350_0, n13321_0, n13320_0}), .out(n4456), .config_in(config_chain[6167:6165]), .config_rst(config_rst)); 
mux6 mux_2056 (.in({n10025_0, n10024_1, n10017_0, n10016_1/**/, n10007_1, n10006_1}), .out(n4457), .config_in(config_chain[6170:6168]), .config_rst(config_rst)); 
mux6 mux_2057 (.in({n13647_1, n13646_0, n13613_0, n13612_0, n13591_0, n13590_0}), .out(n4458), .config_in(config_chain[6173:6171]), .config_rst(config_rst)); 
mux6 mux_2058 (.in({n9825_1, n9824_0, n9811_0, n9810_0, n9757_1, n9756_1}), .out(n4459), .config_in(config_chain[6176:6174]), .config_rst(config_rst)); 
mux6 mux_2059 (.in({n13389_2, n13388_0, n13355_1, n13354_0, n13323_1/**/, n13322_0}), .out(n4460), .config_in(config_chain[6179:6177]), .config_rst(config_rst)); 
mux6 mux_2060 (.in({n10047_0, n10046_0, n10039_0/**/, n10038_0, n10009_1, n10008_1}), .out(n4461), .config_in(config_chain[6182:6180]), .config_rst(config_rst)); 
mux6 mux_2061 (.in({n13649_2, n13648_0, n13623_0, n13622_0, n13585_0, n13584_0}), .out(n4462), .config_in(config_chain[6185:6183]), .config_rst(config_rst)); 
mux6 mux_2062 (.in({n9833_1, n9832_0, n9765_0, n9764_1, n9747_1, n9746_1}), .out(n4463), .config_in(config_chain[6188:6186]), .config_rst(config_rst)); 
mux6 mux_2063 (.in({n13379_1, n13378_0, n13357_0/**/, n13356_0, n13325_0, n13324_0}), .out(n4464), .config_in(config_chain[6191:6189]), .config_rst(config_rst)); 
mux6 mux_2064 (.in({n10079_1/**/, n10078_0, n10067_0, n10066_0, n10011_1, n10010_1}), .out(n4465), .config_in(config_chain[6194:6192]), .config_rst(config_rst)); 
mux6 mux_2065 (.in({n13641_0, n13640_0, n13617_0, n13616_0, n13587_1, n13586_0}), .out(n4466), .config_in(config_chain[6197:6195]), .config_rst(config_rst)); 
mux6 mux_2066 (.in({n9793_0, n9792_0/**/, n9785_0, n9784_0, n9749_1, n9748_1}), .out(n4467), .config_in(config_chain[6200:6198]), .config_rst(config_rst)); 
mux6 mux_2067 (.in({n13381_1, n13380_0, n13359_0, n13358_0, n13329_0, n13328_0}), .out(n4468), .config_in(config_chain[6203:6201]), .config_rst(config_rst)); 
mux6 mux_2068 (.in({n10329_1, n10328_0, n10315_0, n10314_0, n10303_0, n10302_0}), .out(n4515), .config_in(config_chain[6206:6204]), .config_rst(config_rst)); 
mux6 mux_2069 (.in({n13653_1, n13652_0, n13617_0, n13616_0, n13587_0, n13586_0}), .out(n4516), .config_in(config_chain[6209:6207]), .config_rst(config_rst)); 
mux6 mux_2070 (.in({n10033_0, n10032_0, n10027_0, n10026_1/**/, n10019_0, n10018_1}), .out(n4517), .config_in(config_chain[6212:6210]), .config_rst(config_rst)); 
mux6 mux_2071 (.in({n13359_0, n13358_0, n13337_0, n13336_0, n13305_0, n13304_0}), .out(n4518), .config_in(config_chain[6215:6213]), .config_rst(config_rst)); 
mux6 mux_2072 (.in({n10337_1, n10336_0, n10323_0, n10322_0, n10269_0, n10268_1}), .out(n4519), .config_in(config_chain[6218:6216]), .config_rst(config_rst)); 
mux6 mux_2073 (.in({n13669_1, n13668_0, n13661_1, n13660_0, n13567_0, n13566_0}), .out(n4520), .config_in(config_chain[6221:6219]), .config_rst(config_rst)); 
mux6 mux_2074 (.in({n10061_0, n10060_0, n10053_0, n10052_0, n10049_0, n10048_0}), .out(n4521), .config_in(config_chain[6224:6222]), .config_rst(config_rst)); 
mux6 mux_2075 (.in({n13391_1, n13390_0, n13369_0, n13368_0, n13331_0, n13330_0}), .out(n4522), .config_in(config_chain[6227:6225]), .config_rst(config_rst)); 
mux6 mux_2076 (.in({n10289_0, n10288_0, n10285_0, n10284_1, n10277_0, n10276_1}), .out(n4523), .config_in(config_chain[6230:6228]), .config_rst(config_rst)); 
mux6 mux_2077 (.in({n13631_0, n13630_0, n13599_0, n13598_0, n13561_0, n13560_0}), .out(n4524), .config_in(config_chain[6233:6231]), .config_rst(config_rst)); 
mux6 mux_2078 (.in({n10081_1, n10080_0, n10073_1, n10072_0, n10069_0, n10068_0}), .out(n4525), .config_in(config_chain[6236:6234]), .config_rst(config_rst)); 
mux6 mux_2079 (.in({n13399_1, n13398_0, n13363_0, n13362_0, n13303_0, n13302_0}), .out(n4526), .config_in(config_chain[6239:6237]), .config_rst(config_rst)); 
mux6 mux_2080 (.in({n10309_0, n10308_0, n10305_0, n10304_0/**/, n10297_0, n10296_0}), .out(n4527), .config_in(config_chain[6242:6240]), .config_rst(config_rst)); 
mux6 mux_2081 (.in({n13625_0, n13624_0, n13595_0, n13594_0, n13563_0, n13562_0/**/}), .out(n4528), .config_in(config_chain[6245:6243]), .config_rst(config_rst)); 
mux6 mux_2082 (.in({n10089_1, n10088_0/**/, n10035_0, n10034_0, n10021_0, n10020_1}), .out(n4529), .config_in(config_chain[6248:6246]), .config_rst(config_rst)); 
mux6 mux_2083 (.in({n13367_0, n13366_0, n13335_0, n13334_0, n13313_0/**/, n13312_0}), .out(n4530), .config_in(config_chain[6251:6249]), .config_rst(config_rst)); 
mux6 mux_2084 (.in({n10339_1, n10338_0, n10331_1, n10330_0, n10325_0/**/, n10324_0}), .out(n4531), .config_in(config_chain[6254:6252]), .config_rst(config_rst)); 
mux6 mux_2085 (.in({n13663_1, n13662_0, n13627_0, n13626_0, n13575_0, n13574_0}), .out(n4532), .config_in(config_chain[6257:6255]), .config_rst(config_rst)); 
mux6 mux_2086 (.in({n10055_0, n10054_0, n10043_0, n10042_0, n10029_0, n10028_1/**/}), .out(n4533), .config_in(config_chain[6260:6258]), .config_rst(config_rst)); 
mux6 mux_2087 (.in({n13377_0, n13376_0, n13345_0/**/, n13344_0, n13307_0, n13306_0}), .out(n4534), .config_in(config_chain[6263:6261]), .config_rst(config_rst)); 
mux6 mux_2088 (.in({n10347_1, n10346_0, n10279_0, n10278_1, n10271_0/**/, n10270_1}), .out(n4535), .config_in(config_chain[6266:6264]), .config_rst(config_rst)); 
mux6 mux_2089 (.in({n13671_1, n13670_0, n13607_0, n13606_0, n13569_0, n13568_0}), .out(n4536), .config_in(config_chain[6269:6267]), .config_rst(config_rst)); 
mux6 mux_2090 (.in({n10075_1, n10074_0, n10071_0, n10070_0, n10063_0, n10062_0}), .out(n4537), .config_in(config_chain[6272:6270]), .config_rst(config_rst)); 
mux6 mux_2091 (.in({n13401_1, n13400_0, n13393_1, n13392_0, n13371_0, n13370_0}), .out(n4538), .config_in(config_chain[6275:6273]), .config_rst(config_rst)); 
mux6 mux_2092 (.in({n10311_0, n10310_0, n10299_0, n10298_0, n10287_0, n10286_1}), .out(n4539), .config_in(config_chain[6278:6276]), .config_rst(config_rst)); 
mux6 mux_2093 (.in({n13633_0, n13632_0, n13601_0/**/, n13600_0, n13571_0, n13570_0}), .out(n4540), .config_in(config_chain[6281:6279]), .config_rst(config_rst)); 
mux6 mux_2094 (.in({n10091_1, n10090_0/**/, n10023_0, n10022_1, n10015_0, n10014_1}), .out(n4541), .config_in(config_chain[6284:6282]), .config_rst(config_rst)); 
mux6 mux_2095 (.in({n13409_1, n13408_0, n13343_0, n13342_0, n13311_0, n13310_0}), .out(n4542), .config_in(config_chain[6287:6285]), .config_rst(config_rst)); 
mux6 mux_2096 (.in({n10333_1, n10332_0, n10319_0, n10318_0, n10307_0, n10306_0}), .out(n4543), .config_in(config_chain[6290:6288]), .config_rst(config_rst)); 
mux6 mux_2097 (.in({n13657_1, n13656_0, n13635_0, n13634_0, n13603_0, n13602_0}), .out(n4544), .config_in(config_chain[6293:6291]), .config_rst(config_rst)); 
mux6 mux_2098 (.in({n10045_0, n10044_0, n10037_0, n10036_0/**/, n10031_0, n10030_1}), .out(n4545), .config_in(config_chain[6296:6294]), .config_rst(config_rst)); 
mux6 mux_2099 (.in({n13375_0/**/, n13374_0, n13353_0, n13352_0, n13315_0, n13314_0}), .out(n4546), .config_in(config_chain[6299:6297]), .config_rst(config_rst)); 
mux6 mux_2100 (.in({n10341_1, n10340_0, n10273_0, n10272_1/**/, n10257_0, n10256_1}), .out(n4547), .config_in(config_chain[6302:6300]), .config_rst(config_rst)); 
mux6 mux_2101 (.in({n13641_0, n13640_0, n13615_0, n13614_0, n13583_0/**/, n13582_0}), .out(n4548), .config_in(config_chain[6305:6303]), .config_rst(config_rst)); 
mux6 mux_2102 (.in({n10077_1, n10076_0, n10065_0, n10064_0, n10003_1, n10002_1}), .out(n4549), .config_in(config_chain[6308:6306]), .config_rst(config_rst)); 
mux6 mux_2103 (.in({n13395_1/**/, n13394_0, n13381_1, n13380_0, n13347_0, n13346_0}), .out(n4550), .config_in(config_chain[6311:6309]), .config_rst(config_rst)); 
mux6 mux_2104 (.in({n10293_0, n10292_0, n10281_0, n10280_1/**/, n10259_0, n10258_1}), .out(n4551), .config_in(config_chain[6314:6312]), .config_rst(config_rst)); 
mux6 mux_2105 (.in({n13643_0, n13642_0, n13609_0, n13608_0/**/, n13577_0, n13576_0}), .out(n4552), .config_in(config_chain[6317:6315]), .config_rst(config_rst)); 
mux6 mux_2106 (.in({n10085_1, n10084_0, n10017_0, n10016_1, n10005_1, n10004_1}), .out(n4553), .config_in(config_chain[6320:6318]), .config_rst(config_rst)); 
mux6 mux_2107 (.in({n13403_1/**/, n13402_0, n13385_1, n13384_0, n13319_0, n13318_0}), .out(n4554), .config_in(config_chain[6323:6321]), .config_rst(config_rst)); 
mux6 mux_2108 (.in({n10321_0, n10320_0, n10313_0, n10312_0, n10261_1/**/, n10260_1}), .out(n4555), .config_in(config_chain[6326:6324]), .config_rst(config_rst)); 
mux6 mux_2109 (.in({n13659_1, n13658_0, n13645_1, n13644_0, n13611_0, n13610_0}), .out(n4556), .config_in(config_chain[6329:6327]), .config_rst(config_rst)); 
mux6 mux_2110 (.in({n10039_0, n10038_0, n10025_0, n10024_1/**/, n10009_1, n10008_1}), .out(n4557), .config_in(config_chain[6332:6330]), .config_rst(config_rst)); 
mux6 mux_2111 (.in({n13387_2, n13386_0, n13361_0/**/, n13360_0, n13329_0, n13328_0}), .out(n4558), .config_in(config_chain[6335:6333]), .config_rst(config_rst)); 
mux6 mux_2112 (.in({n10343_1, n10342_0, n10335_1/**/, n10334_0, n10263_1, n10262_1}), .out(n4559), .config_in(config_chain[6338:6336]), .config_rst(config_rst)); 
mux6 mux_2113 (.in({n13667_1, n13666_0, n13647_1, n13646_0, n13591_0/**/, n13590_0}), .out(n4560), .config_in(config_chain[6341:6339]), .config_rst(config_rst)); 
mux6 mux_2114 (.in({n10059_0, n10058_0, n10047_0/**/, n10046_0, n10011_1, n10010_1}), .out(n4561), .config_in(config_chain[6344:6342]), .config_rst(config_rst)); 
mux6 mux_2115 (.in({n13389_2, n13388_0, n13355_0, n13354_0, n13323_0/**/, n13322_0}), .out(n4562), .config_in(config_chain[6347:6345]), .config_rst(config_rst)); 
mux6 mux_2116 (.in({n10295_0/**/, n10294_0, n10283_0, n10282_1, n10265_1, n10264_1}), .out(n4563), .config_in(config_chain[6350:6348]), .config_rst(config_rst)); 
mux6 mux_2117 (.in({n13651_2, n13650_0, n13623_0, n13622_0, n13585_0, n13584_0}), .out(n4564), .config_in(config_chain[6353:6351]), .config_rst(config_rst)); 
mux6 mux_2118 (.in({n10087_1, n10086_0, n10079_1, n10078_0/**/, n10001_0, n10000_1}), .out(n4565), .config_in(config_chain[6356:6354]), .config_rst(config_rst)); 
mux6 mux_2119 (.in({n13405_1, n13404_0/**/, n13379_0, n13378_0, n13327_0, n13326_0}), .out(n4566), .config_in(config_chain[6359:6357]), .config_rst(config_rst)); 
mux6 mux_2120 (.in({n10601_1, n10600_0, n10547_0, n10546_0, n10533_0, n10532_1}), .out(n4613), .config_in(config_chain[6362:6360]), .config_rst(config_rst)); 
mux6 mux_2121 (.in({n13687_1, n13686_0, n13585_0, n13584_0, n13563_0/**/, n13562_0}), .out(n4614), .config_in(config_chain[6365:6363]), .config_rst(config_rst)); 
mux6 mux_2122 (.in({n10329_1, n10328_0, n10323_0, n10322_0, n10315_0, n10314_0}), .out(n4615), .config_in(config_chain[6368:6366]), .config_rst(config_rst)); 
mux6 mux_2123 (.in({n13419_1, n13418_0, n13411_1, n13410_0, n13405_0, n13404_0}), .out(n4616), .config_in(config_chain[6371:6369]), .config_rst(config_rst)); 
mux6 mux_2124 (.in({n10567_0, n10566_0, n10555_0, n10554_0, n10541_0, n10540_1/**/}), .out(n4617), .config_in(config_chain[6374:6372]), .config_rst(config_rst)); 
mux6 mux_2125 (.in({n13653_0, n13652_0, n13627_0/**/, n13626_0, n13595_0, n13594_0}), .out(n4618), .config_in(config_chain[6377:6375]), .config_rst(config_rst)); 
mux6 mux_2126 (.in({n10345_1, n10344_0, n10277_0, n10276_1, n10269_0, n10268_1}), .out(n4619), .config_in(config_chain[6380:6378]), .config_rst(config_rst)); 
mux6 mux_2127 (.in({n13427_1, n13426_0, n13337_0, n13336_0, n13299_0, n13298_0}), .out(n4620), .config_in(config_chain[6383:6381]), .config_rst(config_rst)); 
mux6 mux_2128 (.in({n10587_1, n10586_0, n10583_0, n10582_0, n10575_0, n10574_0}), .out(n4621), .config_in(config_chain[6386:6384]), .config_rst(config_rst)); 
mux6 mux_2129 (.in({n13673_1, n13672_0, n13669_0, n13668_0, n13661_0, n13660_0}), .out(n4622), .config_in(config_chain[6389:6387]), .config_rst(config_rst)); 
mux6 mux_2130 (.in({n10297_0, n10296_0, n10289_0, n10288_0, n10285_0, n10284_1}), .out(n4623), .config_in(config_chain[6392:6390]), .config_rst(config_rst)); 
mux6 mux_2131 (.in({n13391_0, n13390_0, n13369_0, n13368_0, n13331_0, n13330_0}), .out(n4624), .config_in(config_chain[6395:6393]), .config_rst(config_rst)); 
mux6 mux_2132 (.in({n10603_1, n10602_0, n10595_1, n10594_0, n10527_0, n10526_1/**/}), .out(n4625), .config_in(config_chain[6398:6396]), .config_rst(config_rst)); 
mux6 mux_2133 (.in({n13689_1, n13688_0, n13593_0, n13592_0, n13561_0/**/, n13560_0}), .out(n4626), .config_in(config_chain[6401:6399]), .config_rst(config_rst)); 
mux6 mux_2134 (.in({n10331_1, n10330_0, n10317_0, n10316_0, n10305_0, n10304_0/**/}), .out(n4627), .config_in(config_chain[6404:6402]), .config_rst(config_rst)); 
mux6 mux_2135 (.in({n13413_1, n13412_0, n13407_0, n13406_0, n13399_0/**/, n13398_0}), .out(n4628), .config_in(config_chain[6407:6405]), .config_rst(config_rst)); 
mux6 mux_2136 (.in({n10557_0, n10556_0, n10549_0, n10548_0, n10543_0/**/, n10542_1}), .out(n4629), .config_in(config_chain[6410:6408]), .config_rst(config_rst)); 
mux6 mux_2137 (.in({n13655_0, n13654_0, n13625_0, n13624_0, n13603_0, n13602_0}), .out(n4630), .config_in(config_chain[6413:6411]), .config_rst(config_rst)); 
mux6 mux_2138 (.in({n10339_1, n10338_0, n10325_0, n10324_0, n10271_0, n10270_1/**/}), .out(n4631), .config_in(config_chain[6416:6414]), .config_rst(config_rst)); 
mux6 mux_2139 (.in({n13429_1, n13428_0, n13421_1, n13420_0, n13313_0, n13312_0}), .out(n4632), .config_in(config_chain[6419:6417]), .config_rst(config_rst)); 
mux6 mux_2140 (.in({n10577_0, n10576_0, n10569_0, n10568_0, n10565_0, n10564_0}), .out(n4633), .config_in(config_chain[6422:6420]), .config_rst(config_rst)); 
mux6 mux_2141 (.in({n13675_1, n13674_0, n13663_0, n13662_0, n13635_0, n13634_0}), .out(n4634), .config_in(config_chain[6425:6423]), .config_rst(config_rst)); 
mux6 mux_2142 (.in({n10291_0, n10290_0, n10287_0, n10286_1, n10279_0, n10278_1/**/}), .out(n4635), .config_in(config_chain[6428:6426]), .config_rst(config_rst)); 
mux6 mux_2143 (.in({n13377_0, n13376_0, n13339_0, n13338_0, n13307_0, n13306_0}), .out(n4636), .config_in(config_chain[6431:6429]), .config_rst(config_rst)); 
mux6 mux_2144 (.in({n10597_1, n10596_0, n10585_0, n10584_0, n10529_0, n10528_1}), .out(n4637), .config_in(config_chain[6434:6432]), .config_rst(config_rst)); 
mux6 mux_2145 (.in({n13691_1, n13690_0, n13683_1, n13682_0, n13569_0, n13568_0/**/}), .out(n4638), .config_in(config_chain[6437:6435]), .config_rst(config_rst)); 
mux6 mux_2146 (.in({n10319_0, n10318_0, n10311_0/**/, n10310_0, n10307_0, n10306_0}), .out(n4639), .config_in(config_chain[6440:6438]), .config_rst(config_rst)); 
mux6 mux_2147 (.in({n13401_0, n13400_0, n13393_0, n13392_0/**/, n13371_0, n13370_0}), .out(n4640), .config_in(config_chain[6443:6441]), .config_rst(config_rst)); 
mux6 mux_2148 (.in({n10605_1/**/, n10604_0, n10551_0, n10550_0, n10537_0, n10536_1}), .out(n4641), .config_in(config_chain[6446:6444]), .config_rst(config_rst)); 
mux6 mux_2149 (.in({n13633_0, n13632_0, n13601_0, n13600_0/**/, n13579_0, n13578_0}), .out(n4642), .config_in(config_chain[6449:6447]), .config_rst(config_rst)); 
mux6 mux_2150 (.in({n10341_1/**/, n10340_0, n10333_1, n10332_0, n10327_0, n10326_0}), .out(n4643), .config_in(config_chain[6452:6450]), .config_rst(config_rst)); 
mux6 mux_2151 (.in({n13423_1, n13422_0, n13409_0, n13408_0, n13321_0, n13320_0/**/}), .out(n4644), .config_in(config_chain[6455:6453]), .config_rst(config_rst)); 
mux6 mux_2152 (.in({n10571_0, n10570_0, n10559_0, n10558_0, n10525_1, n10524_1}), .out(n4645), .config_in(config_chain[6458:6456]), .config_rst(config_rst)); 
mux6 mux_2153 (.in({n13665_0/**/, n13664_0, n13657_0, n13656_0, n13651_1, n13650_0}), .out(n4646), .config_in(config_chain[6461:6459]), .config_rst(config_rst)); 
mux6 mux_2154 (.in({n10293_0, n10292_0, n10281_0/**/, n10280_1, n10257_0, n10256_1}), .out(n4647), .config_in(config_chain[6464:6462]), .config_rst(config_rst)); 
mux6 mux_2155 (.in({n13379_0, n13378_0, n13353_0, n13352_0, n13315_0/**/, n13314_0}), .out(n4648), .config_in(config_chain[6467:6465]), .config_rst(config_rst)); 
mux6 mux_2156 (.in({n10591_1, n10590_0, n10579_0, n10578_0, n10515_0, n10514_1}), .out(n4649), .config_in(config_chain[6470:6468]), .config_rst(config_rst)); 
mux6 mux_2157 (.in({n13685_1, n13684_0, n13677_1, n13676_0, n13641_0, n13640_0}), .out(n4650), .config_in(config_chain[6473:6471]), .config_rst(config_rst)); 
mux6 mux_2158 (.in({n10313_0, n10312_0, n10301_0, n10300_0, n10259_0, n10258_1}), .out(n4651), .config_in(config_chain[6476:6474]), .config_rst(config_rst)); 
mux6 mux_2159 (.in({n13395_0, n13394_0, n13383_1, n13382_0, n13347_0, n13346_0}), .out(n4652), .config_in(config_chain[6479:6477]), .config_rst(config_rst)); 
mux6 mux_2160 (.in({n10539_0, n10538_1/**/, n10531_0, n10530_1, n10517_0, n10516_1}), .out(n4653), .config_in(config_chain[6482:6480]), .config_rst(config_rst)); 
mux6 mux_2161 (.in({n13643_0, n13642_0, n13609_0, n13608_0, n13587_0, n13586_0}), .out(n4654), .config_in(config_chain[6485:6483]), .config_rst(config_rst)); 
mux6 mux_2162 (.in({n10335_1, n10334_0/**/, n10321_0, n10320_0, n10263_1, n10262_1}), .out(n4655), .config_in(config_chain[6488:6486]), .config_rst(config_rst)); 
mux6 mux_2163 (.in({n13425_1, n13424_0, n13417_1/**/, n13416_0, n13385_1, n13384_0}), .out(n4656), .config_in(config_chain[6491:6489]), .config_rst(config_rst)); 
mux6 mux_2164 (.in({n10561_0, n10560_0, n10553_0, n10552_0/**/, n10519_0, n10518_1}), .out(n4657), .config_in(config_chain[6494:6492]), .config_rst(config_rst)); 
mux6 mux_2165 (.in({n13659_0, n13658_0, n13645_0, n13644_0, n13619_0, n13618_0}), .out(n4658), .config_in(config_chain[6497:6495]), .config_rst(config_rst)); 
mux6 mux_2166 (.in({n10343_1, n10342_0, n10275_0, n10274_1/**/, n10265_1, n10264_1}), .out(n4659), .config_in(config_chain[6500:6498]), .config_rst(config_rst)); 
mux6 mux_2167 (.in({n13387_1, n13386_0, n13361_0, n13360_0, n13329_0/**/, n13328_0}), .out(n4660), .config_in(config_chain[6503:6501]), .config_rst(config_rst)); 
mux6 mux_2168 (.in({n10593_1, n10592_0, n10581_0, n10580_0/**/, n10521_1, n10520_1}), .out(n4661), .config_in(config_chain[6506:6504]), .config_rst(config_rst)); 
mux6 mux_2169 (.in({n13679_1, n13678_0, n13667_0/**/, n13666_0, n13649_1, n13648_0}), .out(n4662), .config_in(config_chain[6509:6507]), .config_rst(config_rst)); 
mux6 mux_2170 (.in({n10303_0, n10302_0, n10295_0/**/, n10294_0, n10267_1, n10266_1}), .out(n4663), .config_in(config_chain[6512:6510]), .config_rst(config_rst)); 
mux6 mux_2171 (.in({n13397_0, n13396_0, n13389_2, n13388_0, n13355_0/**/, n13354_0}), .out(n4664), .config_in(config_chain[6515:6513]), .config_rst(config_rst)); 
mux6 mux_2172 (.in({n10847_1, n10846_0, n10833_0, n10832_0, n10821_0, n10820_0}), .out(n4711), .config_in(config_chain[6518:6516]), .config_rst(config_rst)); 
mux6 mux_2173 (.in({n13693_1, n13692_0, n13679_0, n13678_0/**/, n13667_0, n13666_0}), .out(n4712), .config_in(config_chain[6521:6519]), .config_rst(config_rst)); 
mux6 mux_2174 (.in({n10547_0, n10546_0, n10541_0, n10540_1, n10533_0, n10532_1}), .out(n4713), .config_in(config_chain[6524:6522]), .config_rst(config_rst)); 
mux6 mux_2175 (.in({n13399_0, n13398_0, n13391_0, n13390_0, n13355_0, n13354_1}), .out(n4714), .config_in(config_chain[6527:6525]), .config_rst(config_rst)); 
mux6 mux_2176 (.in({n10855_1, n10854_0, n10841_0, n10840_0, n10787_0, n10786_1}), .out(n4715), .config_in(config_chain[6530:6528]), .config_rst(config_rst)); 
mux6 mux_2177 (.in({n13709_1, n13708_0, n13701_1, n13700_0, n13563_0, n13562_1}), .out(n4716), .config_in(config_chain[6533:6531]), .config_rst(config_rst)); 
mux6 mux_2178 (.in({n10575_0, n10574_0, n10567_0, n10566_0, n10563_0, n10562_0}), .out(n4717), .config_in(config_chain[6536:6534]), .config_rst(config_rst)); 
mux6 mux_2179 (.in({n13431_1, n13430_0, n13419_0, n13418_0, n13407_0, n13406_0/**/}), .out(n4718), .config_in(config_chain[6539:6537]), .config_rst(config_rst)); 
mux6 mux_2180 (.in({n10807_0, n10806_0, n10803_0, n10802_1, n10795_0, n10794_1}), .out(n4719), .config_in(config_chain[6542:6540]), .config_rst(config_rst)); 
mux6 mux_2181 (.in({n13653_0, n13652_0, n13627_0, n13626_1, n13595_0, n13594_1}), .out(n4720), .config_in(config_chain[6545:6543]), .config_rst(config_rst)); 
mux6 mux_2182 (.in({n10595_1, n10594_0, n10587_1, n10586_0, n10583_0, n10582_0}), .out(n4721), .config_in(config_chain[6548:6546]), .config_rst(config_rst)); 
mux6 mux_2183 (.in({n13439_1, n13438_0, n13427_0, n13426_0, n13299_0, n13298_1}), .out(n4722), .config_in(config_chain[6551:6549]), .config_rst(config_rst)); 
mux6 mux_2184 (.in({n10827_0, n10826_0, n10823_0, n10822_0, n10815_0, n10814_0}), .out(n4723), .config_in(config_chain[6554:6552]), .config_rst(config_rst)); 
mux6 mux_2185 (.in({n13681_0, n13680_0, n13673_0, n13672_0, n13669_0, n13668_0}), .out(n4724), .config_in(config_chain[6557:6555]), .config_rst(config_rst)); 
mux6 mux_2186 (.in({n10603_1/**/, n10602_0, n10549_0, n10548_0, n10535_0, n10534_1}), .out(n4725), .config_in(config_chain[6560:6558]), .config_rst(config_rst)); 
mux6 mux_2187 (.in({n13393_0, n13392_0, n13363_0, n13362_1, n13331_0/**/, n13330_1}), .out(n4726), .config_in(config_chain[6563:6561]), .config_rst(config_rst)); 
mux6 mux_2188 (.in({n10857_1, n10856_0, n10849_1, n10848_0, n10843_0, n10842_0/**/}), .out(n4727), .config_in(config_chain[6566:6564]), .config_rst(config_rst)); 
mux6 mux_2189 (.in({n13703_1, n13702_0, n13689_0, n13688_0, n13571_0, n13570_1}), .out(n4728), .config_in(config_chain[6569:6567]), .config_rst(config_rst)); 
mux6 mux_2190 (.in({n10569_0, n10568_0, n10557_0, n10556_0, n10543_0, n10542_1}), .out(n4729), .config_in(config_chain[6572:6570]), .config_rst(config_rst)); 
mux6 mux_2191 (.in({n13413_0, n13412_0, n13409_0, n13408_0, n13401_0, n13400_0}), .out(n4730), .config_in(config_chain[6575:6573]), .config_rst(config_rst)); 
mux6 mux_2192 (.in({n10865_1, n10864_0, n10797_0, n10796_1, n10789_0, n10788_1/**/}), .out(n4731), .config_in(config_chain[6578:6576]), .config_rst(config_rst)); 
mux6 mux_2193 (.in({n13711_1, n13710_0, n13655_0, n13654_0, n13603_0/**/, n13602_1}), .out(n4732), .config_in(config_chain[6581:6579]), .config_rst(config_rst)); 
mux6 mux_2194 (.in({n10589_1, n10588_0, n10585_0, n10584_0/**/, n10577_0, n10576_0}), .out(n4733), .config_in(config_chain[6584:6582]), .config_rst(config_rst)); 
mux6 mux_2195 (.in({n13441_1, n13440_0, n13433_1, n13432_0/**/, n13429_0, n13428_0}), .out(n4734), .config_in(config_chain[6587:6585]), .config_rst(config_rst)); 
mux6 mux_2196 (.in({n10829_0/**/, n10828_0, n10817_0, n10816_0, n10805_0, n10804_1}), .out(n4735), .config_in(config_chain[6590:6588]), .config_rst(config_rst)); 
mux6 mux_2197 (.in({n13675_0, n13674_0, n13671_0, n13670_0/**/, n13663_0, n13662_0}), .out(n4736), .config_in(config_chain[6593:6591]), .config_rst(config_rst)); 
mux6 mux_2198 (.in({n10605_1, n10604_0, n10537_0, n10536_1, n10529_0, n10528_1}), .out(n4737), .config_in(config_chain[6596:6594]), .config_rst(config_rst)); 
mux6 mux_2199 (.in({n13449_1, n13448_0, n13339_0, n13338_1, n13307_0, n13306_1/**/}), .out(n4738), .config_in(config_chain[6599:6597]), .config_rst(config_rst)); 
mux6 mux_2200 (.in({n10851_1, n10850_0, n10837_0, n10836_0, n10825_0, n10824_0/**/}), .out(n4739), .config_in(config_chain[6602:6600]), .config_rst(config_rst)); 
mux6 mux_2201 (.in({n13697_1, n13696_0, n13691_0/**/, n13690_0, n13683_0, n13682_0}), .out(n4740), .config_in(config_chain[6605:6603]), .config_rst(config_rst)); 
mux6 mux_2202 (.in({n10559_0, n10558_0, n10551_0, n10550_0, n10545_0, n10544_1}), .out(n4741), .config_in(config_chain[6608:6606]), .config_rst(config_rst)); 
mux6 mux_2203 (.in({n13415_0, n13414_0, n13403_0, n13402_0, n13371_0, n13370_1}), .out(n4742), .config_in(config_chain[6611:6609]), .config_rst(config_rst)); 
mux6 mux_2204 (.in({n10859_1, n10858_0, n10791_0, n10790_1/**/, n10783_1, n10782_1}), .out(n4743), .config_in(config_chain[6614:6612]), .config_rst(config_rst)); 
mux6 mux_2205 (.in({n13649_1, n13648_1, n13611_0/**/, n13610_1, n13579_0, n13578_1}), .out(n4744), .config_in(config_chain[6617:6615]), .config_rst(config_rst)); 
mux6 mux_2206 (.in({n10591_1, n10590_0, n10579_0, n10578_0/**/, n10525_1, n10524_1}), .out(n4745), .config_in(config_chain[6620:6618]), .config_rst(config_rst)); 
mux6 mux_2207 (.in({n13435_1, n13434_0/**/, n13423_0, n13422_0, n13389_1, n13388_1}), .out(n4746), .config_in(config_chain[6623:6621]), .config_rst(config_rst)); 
mux6 mux_2208 (.in({n10811_0, n10810_0, n10799_0, n10798_1, n10785_1/**/, n10784_1}), .out(n4747), .config_in(config_chain[6626:6624]), .config_rst(config_rst)); 
mux6 mux_2209 (.in({n13665_0, n13664_0, n13657_0, n13656_0, n13651_1, n13650_1}), .out(n4748), .config_in(config_chain[6629:6627]), .config_rst(config_rst)); 
mux6 mux_2210 (.in({n10599_1, n10598_0, n10531_0, n10530_1/**/, n10515_0, n10514_1}), .out(n4749), .config_in(config_chain[6632:6630]), .config_rst(config_rst)); 
mux6 mux_2211 (.in({n13443_1, n13442_0, n13381_0, n13380_1, n13315_0, n13314_1}), .out(n4750), .config_in(config_chain[6635:6633]), .config_rst(config_rst)); 
mux6 mux_2212 (.in({n10867_1, n10866_0, n10839_0, n10838_0/**/, n10831_0, n10830_0}), .out(n4751), .config_in(config_chain[6638:6636]), .config_rst(config_rst)); 
mux6 mux_2213 (.in({n13713_1, n13712_0, n13699_1, n13698_0, n13685_0, n13684_0}), .out(n4752), .config_in(config_chain[6641:6639]), .config_rst(config_rst)); 
mux6 mux_2214 (.in({n10553_0, n10552_0, n10539_0, n10538_1, n10519_0, n10518_1}), .out(n4753), .config_in(config_chain[6644:6642]), .config_rst(config_rst)); 
mux6 mux_2215 (.in({n13405_0, n13404_0, n13397_0, n13396_0, n13383_0, n13382_1}), .out(n4754), .config_in(config_chain[6647:6645]), .config_rst(config_rst)); 
mux6 mux_2216 (.in({n10861_1, n10860_0, n10853_1, n10852_0, n10777_0/**/, n10776_1}), .out(n4755), .config_in(config_chain[6650:6648]), .config_rst(config_rst)); 
mux6 mux_2217 (.in({n13707_1/**/, n13706_0, n13643_0, n13642_1, n13587_0, n13586_1}), .out(n4756), .config_in(config_chain[6653:6651]), .config_rst(config_rst)); 
mux6 mux_2218 (.in({n10573_0/**/, n10572_0, n10561_0, n10560_0, n10521_1, n10520_1}), .out(n4757), .config_in(config_chain[6656:6654]), .config_rst(config_rst)); 
mux6 mux_2219 (.in({n13425_0/**/, n13424_0, n13417_0, n13416_0, n13385_1, n13384_1}), .out(n4758), .config_in(config_chain[6659:6657]), .config_rst(config_rst)); 
mux6 mux_2220 (.in({n10813_0, n10812_0, n10801_0, n10800_1, n10779_0, n10778_1}), .out(n4759), .config_in(config_chain[6662:6660]), .config_rst(config_rst)); 
mux6 mux_2221 (.in({n13659_0/**/, n13658_0, n13647_0, n13646_1, n13619_0, n13618_1}), .out(n4760), .config_in(config_chain[6665:6663]), .config_rst(config_rst)); 
mux6 mux_2222 (.in({n10601_1, n10600_0, n10593_1, n10592_0, n10523_1, n10522_1}), .out(n4761), .config_in(config_chain[6668:6666]), .config_rst(config_rst)); 
mux6 mux_2223 (.in({n13445_1, n13444_0, n13387_1, n13386_1, n13323_0, n13322_1}), .out(n4762), .config_in(config_chain[6671:6669]), .config_rst(config_rst)); 
mux6 mux_2224 (.in({n11125_1, n11124_0, n11069_0/**/, n11068_0, n11055_0, n11054_1}), .out(n4809), .config_in(config_chain[6674:6672]), .config_rst(config_rst)); 
mux6 mux_2225 (.in({n13729_1, n13728_0, n13673_0, n13672_0, n13659_0, n13658_1}), .out(n4810), .config_in(config_chain[6677:6675]), .config_rst(config_rst)); 
mux6 mux_2226 (.in({n10847_1, n10846_0, n10841_0, n10840_0, n10833_0, n10832_0}), .out(n4811), .config_in(config_chain[6680:6678]), .config_rst(config_rst)); 
mux6 mux_2227 (.in({n13459_1, n13458_0, n13451_1, n13450_0, n13445_0, n13444_0/**/}), .out(n4812), .config_in(config_chain[6683:6681]), .config_rst(config_rst)); 
mux6 mux_2228 (.in({n11089_0, n11088_0, n11077_0, n11076_0/**/, n11063_0, n11062_1}), .out(n4813), .config_in(config_chain[6686:6684]), .config_rst(config_rst)); 
mux6 mux_2229 (.in({n13693_0, n13692_0, n13689_0, n13688_0, n13681_0, n13680_0}), .out(n4814), .config_in(config_chain[6689:6687]), .config_rst(config_rst)); 
mux6 mux_2230 (.in({n10863_1/**/, n10862_0, n10795_0, n10794_1, n10787_0, n10786_1}), .out(n4815), .config_in(config_chain[6692:6690]), .config_rst(config_rst)); 
mux6 mux_2231 (.in({n13467_1, n13466_0, n13411_0, n13410_0, n13399_0, n13398_1/**/}), .out(n4816), .config_in(config_chain[6695:6693]), .config_rst(config_rst)); 
mux6 mux_2232 (.in({n11111_1, n11110_0/**/, n11105_0, n11104_0, n11097_0, n11096_0}), .out(n4817), .config_in(config_chain[6698:6696]), .config_rst(config_rst)); 
mux6 mux_2233 (.in({n13715_1, n13714_0, n13709_0, n13708_0, n13701_0, n13700_0}), .out(n4818), .config_in(config_chain[6701:6699]), .config_rst(config_rst)); 
mux6 mux_2234 (.in({n10815_0, n10814_0, n10807_0, n10806_0, n10803_0, n10802_1}), .out(n4819), .config_in(config_chain[6704:6702]), .config_rst(config_rst)); 
mux6 mux_2235 (.in({n13431_0/**/, n13430_0, n13419_0, n13418_0, n13407_0, n13406_1}), .out(n4820), .config_in(config_chain[6707:6705]), .config_rst(config_rst)); 
mux6 mux_2236 (.in({n11127_1/**/, n11126_0, n11119_1, n11118_0, n11049_0, n11048_1}), .out(n4821), .config_in(config_chain[6710:6708]), .config_rst(config_rst)); 
mux6 mux_2237 (.in({n13731_1, n13730_0, n13661_0, n13660_1, n13653_0/**/, n13652_1}), .out(n4822), .config_in(config_chain[6713:6711]), .config_rst(config_rst)); 
mux6 mux_2238 (.in({n10849_1, n10848_0, n10835_0, n10834_0, n10823_0, n10822_0}), .out(n4823), .config_in(config_chain[6716:6714]), .config_rst(config_rst)); 
mux6 mux_2239 (.in({n13453_1, n13452_0/**/, n13447_0, n13446_0, n13439_0, n13438_0}), .out(n4824), .config_in(config_chain[6719:6717]), .config_rst(config_rst)); 
mux6 mux_2240 (.in({n11079_0, n11078_0, n11071_0/**/, n11070_0, n11065_0, n11064_1}), .out(n4825), .config_in(config_chain[6722:6720]), .config_rst(config_rst)); 
mux6 mux_2241 (.in({n13695_0, n13694_0, n13683_0, n13682_0, n13669_0, n13668_1}), .out(n4826), .config_in(config_chain[6725:6723]), .config_rst(config_rst)); 
mux6 mux_2242 (.in({n10857_1, n10856_0/**/, n10843_0, n10842_0, n10789_0, n10788_1}), .out(n4827), .config_in(config_chain[6728:6726]), .config_rst(config_rst)); 
mux6 mux_2243 (.in({n13469_1, n13468_0, n13461_1, n13460_0/**/, n13393_0, n13392_1}), .out(n4828), .config_in(config_chain[6731:6729]), .config_rst(config_rst)); 
mux6 mux_2244 (.in({n11099_0, n11098_0, n11091_0, n11090_0/**/, n11087_0, n11086_0}), .out(n4829), .config_in(config_chain[6734:6732]), .config_rst(config_rst)); 
mux6 mux_2245 (.in({n13717_1, n13716_0, n13703_0, n13702_0, n13691_0, n13690_0}), .out(n4830), .config_in(config_chain[6737:6735]), .config_rst(config_rst)); 
mux6 mux_2246 (.in({n10809_0, n10808_0, n10805_0, n10804_1/**/, n10797_0, n10796_1}), .out(n4831), .config_in(config_chain[6740:6738]), .config_rst(config_rst)); 
mux6 mux_2247 (.in({n13421_0/**/, n13420_0, n13413_0, n13412_0, n13409_0, n13408_1}), .out(n4832), .config_in(config_chain[6743:6741]), .config_rst(config_rst)); 
mux6 mux_2248 (.in({n11121_1, n11120_0, n11107_0, n11106_0, n11051_0, n11050_1/**/}), .out(n4833), .config_in(config_chain[6746:6744]), .config_rst(config_rst)); 
mux6 mux_2249 (.in({n13733_1, n13732_0/**/, n13725_1, n13724_0, n13655_0, n13654_1}), .out(n4834), .config_in(config_chain[6749:6747]), .config_rst(config_rst)); 
mux6 mux_2250 (.in({n10837_0, n10836_0/**/, n10829_0, n10828_0, n10825_0, n10824_0}), .out(n4835), .config_in(config_chain[6752:6750]), .config_rst(config_rst)); 
mux6 mux_2251 (.in({n13441_0, n13440_0, n13433_0, n13432_0, n13429_0/**/, n13428_0}), .out(n4836), .config_in(config_chain[6755:6753]), .config_rst(config_rst)); 
mux6 mux_2252 (.in({n11129_1, n11128_0/**/, n11073_0, n11072_0, n11059_0, n11058_1}), .out(n4837), .config_in(config_chain[6758:6756]), .config_rst(config_rst)); 
mux6 mux_2253 (.in({n13677_0, n13676_0/**/, n13671_0, n13670_1, n13663_0, n13662_1}), .out(n4838), .config_in(config_chain[6761:6759]), .config_rst(config_rst)); 
mux6 mux_2254 (.in({n10859_1, n10858_0, n10851_1, n10850_0, n10845_0, n10844_0/**/}), .out(n4839), .config_in(config_chain[6764:6762]), .config_rst(config_rst)); 
mux6 mux_2255 (.in({n13463_1, n13462_0, n13449_0, n13448_0, n13395_0, n13394_1}), .out(n4840), .config_in(config_chain[6767:6765]), .config_rst(config_rst)); 
mux6 mux_2256 (.in({n11093_0, n11092_0, n11081_0/**/, n11080_0, n11043_0, n11042_1}), .out(n4841), .config_in(config_chain[6770:6768]), .config_rst(config_rst)); 
mux6 mux_2257 (.in({n13705_0, n13704_0, n13697_0, n13696_0, n13647_0, n13646_1}), .out(n4842), .config_in(config_chain[6773:6771]), .config_rst(config_rst)); 
mux6 mux_2258 (.in({n10811_0, n10810_0, n10799_0, n10798_1, n10783_1, n10782_1}), .out(n4843), .config_in(config_chain[6776:6774]), .config_rst(config_rst)); 
mux6 mux_2259 (.in({n13415_0, n13414_0, n13403_0, n13402_1/**/, n13387_1, n13386_1}), .out(n4844), .config_in(config_chain[6779:6777]), .config_rst(config_rst)); 
mux6 mux_2260 (.in({n11115_1, n11114_0, n11101_0, n11100_0, n11045_0/**/, n11044_1}), .out(n4845), .config_in(config_chain[6782:6780]), .config_rst(config_rst)); 
mux6 mux_2261 (.in({n13727_1, n13726_0, n13719_1, n13718_0/**/, n13649_0, n13648_1}), .out(n4846), .config_in(config_chain[6785:6783]), .config_rst(config_rst)); 
mux6 mux_2262 (.in({n10831_0, n10830_0, n10819_0, n10818_0, n10785_1, n10784_1}), .out(n4847), .config_in(config_chain[6788:6786]), .config_rst(config_rst)); 
mux6 mux_2263 (.in({n13471_1/**/, n13470_0, n13435_0, n13434_0, n13423_0, n13422_0}), .out(n4848), .config_in(config_chain[6791:6789]), .config_rst(config_rst)); 
mux6 mux_2264 (.in({n11061_0/**/, n11060_1, n11053_0, n11052_1, n11047_1, n11046_1}), .out(n4849), .config_in(config_chain[6794:6792]), .config_rst(config_rst)); 
mux6 mux_2265 (.in({n13679_0, n13678_0, n13665_0, n13664_1/**/, n13651_1, n13650_1}), .out(n4850), .config_in(config_chain[6797:6795]), .config_rst(config_rst)); 
mux6 mux_2266 (.in({n10853_1, n10852_0, n10839_0, n10838_0, n10777_0, n10776_1}), .out(n4851), .config_in(config_chain[6800:6798]), .config_rst(config_rst)); 
mux6 mux_2267 (.in({n13465_1, n13464_0, n13457_1/**/, n13456_0, n13381_0, n13380_1}), .out(n4852), .config_in(config_chain[6803:6801]), .config_rst(config_rst)); 
mux6 mux_2268 (.in({n11109_1, n11108_0, n11083_0, n11082_0, n11075_0, n11074_0}), .out(n4853), .config_in(config_chain[6806:6804]), .config_rst(config_rst)); 
mux6 mux_2269 (.in({n13713_1, n13712_0, n13699_0, n13698_0/**/, n13687_0, n13686_0}), .out(n4854), .config_in(config_chain[6809:6807]), .config_rst(config_rst)); 
mux6 mux_2270 (.in({n10861_1, n10860_0, n10793_0, n10792_1, n10779_0/**/, n10778_1}), .out(n4855), .config_in(config_chain[6812:6810]), .config_rst(config_rst)); 
mux6 mux_2271 (.in({n13405_0, n13404_1/**/, n13397_0, n13396_1, n13383_0, n13382_1}), .out(n4856), .config_in(config_chain[6815:6813]), .config_rst(config_rst)); 
mux6 mux_2272 (.in({n11131_1, n11130_0, n11117_1, n11116_0, n11103_0, n11102_0/**/}), .out(n4857), .config_in(config_chain[6818:6816]), .config_rst(config_rst)); 
mux6 mux_2273 (.in({n13721_1, n13720_0, n13707_0, n13706_0, n13645_0, n13644_1}), .out(n4858), .config_in(config_chain[6821:6819]), .config_rst(config_rst)); 
mux6 mux_2274 (.in({n10821_0, n10820_0, n10813_0, n10812_0/**/, n10781_0, n10780_1}), .out(n4859), .config_in(config_chain[6824:6822]), .config_rst(config_rst)); 
mux6 mux_2275 (.in({n13437_0, n13436_0, n13425_0/**/, n13424_0, n13385_0, n13384_1}), .out(n4860), .config_in(config_chain[6827:6825]), .config_rst(config_rst)); 
mux6 mux_2276 (.in({n11377_1, n11376_0, n11361_0, n11360_0, n11347_0, n11346_0}), .out(n4907), .config_in(config_chain[6830:6828]), .config_rst(config_rst)); 
mux6 mux_2277 (.in({n13737_1, n13736_0, n13721_0, n13720_0, n13707_0, n13706_0}), .out(n4908), .config_in(config_chain[6833:6831]), .config_rst(config_rst)); 
mux6 mux_2278 (.in({n11069_0, n11068_0, n11063_0, n11062_1, n11055_0/**/, n11054_1}), .out(n4909), .config_in(config_chain[6836:6834]), .config_rst(config_rst)); 
mux6 mux_2279 (.in({n13439_0, n13438_0, n13431_0, n13430_0, n13425_0, n13424_1}), .out(n4910), .config_in(config_chain[6839:6837]), .config_rst(config_rst)); 
mux6 mux_2280 (.in({n11385_1, n11384_0, n11369_0, n11368_0, n11313_0, n11312_1/**/}), .out(n4911), .config_in(config_chain[6842:6840]), .config_rst(config_rst)); 
mux6 mux_2281 (.in({n13753_1, n13752_0, n13745_1/**/, n13744_0, n13673_0, n13672_1}), .out(n4912), .config_in(config_chain[6845:6843]), .config_rst(config_rst)); 
mux6 mux_2282 (.in({n11097_0, n11096_0/**/, n11089_0, n11088_0, n11085_0, n11084_0}), .out(n4913), .config_in(config_chain[6848:6846]), .config_rst(config_rst)); 
mux6 mux_2283 (.in({n13473_1/**/, n13472_0, n13459_0, n13458_0, n13447_0, n13446_0}), .out(n4914), .config_in(config_chain[6851:6849]), .config_rst(config_rst)); 
mux6 mux_2284 (.in({n11333_0, n11332_0, n11329_0, n11328_1/**/, n11321_0, n11320_1}), .out(n4915), .config_in(config_chain[6854:6852]), .config_rst(config_rst)); 
mux6 mux_2285 (.in({n13693_0, n13692_0/**/, n13689_0, n13688_1, n13681_0, n13680_1}), .out(n4916), .config_in(config_chain[6857:6855]), .config_rst(config_rst)); 
mux6 mux_2286 (.in({n11119_1, n11118_0, n11111_1, n11110_0, n11105_0, n11104_0}), .out(n4917), .config_in(config_chain[6860:6858]), .config_rst(config_rst)); 
mux6 mux_2287 (.in({n13481_1, n13480_0, n13467_0, n13466_0, n13411_0, n13410_1}), .out(n4918), .config_in(config_chain[6863:6861]), .config_rst(config_rst)); 
mux6 mux_2288 (.in({n11355_0, n11354_0, n11349_0, n11348_0, n11341_0, n11340_0}), .out(n4919), .config_in(config_chain[6866:6864]), .config_rst(config_rst)); 
mux6 mux_2289 (.in({n13723_0, n13722_0, n13715_0, n13714_0, n13709_0, n13708_0/**/}), .out(n4920), .config_in(config_chain[6869:6867]), .config_rst(config_rst)); 
mux6 mux_2290 (.in({n11127_1, n11126_0, n11071_0, n11070_0, n11057_0, n11056_1}), .out(n4921), .config_in(config_chain[6872:6870]), .config_rst(config_rst)); 
mux6 mux_2291 (.in({n13433_0, n13432_0, n13427_0, n13426_1, n13419_0, n13418_1/**/}), .out(n4922), .config_in(config_chain[6875:6873]), .config_rst(config_rst)); 
mux6 mux_2292 (.in({n11387_1, n11386_0, n11379_1, n11378_0, n11371_0/**/, n11370_0}), .out(n4923), .config_in(config_chain[6878:6876]), .config_rst(config_rst)); 
mux6 mux_2293 (.in({n13747_1, n13746_0, n13731_0, n13730_0, n13675_0, n13674_1}), .out(n4924), .config_in(config_chain[6881:6879]), .config_rst(config_rst)); 
mux6 mux_2294 (.in({n11091_0, n11090_0, n11079_0, n11078_0/**/, n11065_0, n11064_1}), .out(n4925), .config_in(config_chain[6884:6882]), .config_rst(config_rst)); 
mux6 mux_2295 (.in({n13453_0/**/, n13452_0, n13449_0, n13448_0, n13441_0, n13440_0}), .out(n4926), .config_in(config_chain[6887:6885]), .config_rst(config_rst)); 
mux6 mux_2296 (.in({n11395_1, n11394_0, n11323_0, n11322_1, n11315_0, n11314_1}), .out(n4927), .config_in(config_chain[6890:6888]), .config_rst(config_rst)); 
mux6 mux_2297 (.in({n13755_1, n13754_0, n13695_0, n13694_0/**/, n13683_0, n13682_1}), .out(n4928), .config_in(config_chain[6893:6891]), .config_rst(config_rst)); 
mux6 mux_2298 (.in({n11113_1, n11112_0, n11107_0, n11106_0, n11099_0, n11098_0/**/}), .out(n4929), .config_in(config_chain[6896:6894]), .config_rst(config_rst)); 
mux6 mux_2299 (.in({n13483_1, n13482_0, n13475_1, n13474_0, n13469_0, n13468_0/**/}), .out(n4930), .config_in(config_chain[6899:6897]), .config_rst(config_rst)); 
mux6 mux_2300 (.in({n11357_0, n11356_0/**/, n11343_0, n11342_0, n11331_0, n11330_1}), .out(n4931), .config_in(config_chain[6902:6900]), .config_rst(config_rst)); 
mux6 mux_2301 (.in({n13717_0, n13716_0, n13711_0, n13710_0, n13703_0/**/, n13702_0}), .out(n4932), .config_in(config_chain[6905:6903]), .config_rst(config_rst)); 
mux6 mux_2302 (.in({n11129_1, n11128_0, n11059_0, n11058_1, n11051_0, n11050_1}), .out(n4933), .config_in(config_chain[6908:6906]), .config_rst(config_rst)); 
mux6 mux_2303 (.in({n13491_1, n13490_0, n13421_0, n13420_1, n13413_0/**/, n13412_1}), .out(n4934), .config_in(config_chain[6911:6909]), .config_rst(config_rst)); 
mux6 mux_2304 (.in({n11381_1, n11380_0, n11365_0, n11364_0, n11351_0, n11350_0/**/}), .out(n4935), .config_in(config_chain[6914:6912]), .config_rst(config_rst)); 
mux6 mux_2305 (.in({n13741_1, n13740_0, n13733_0, n13732_0, n13725_0/**/, n13724_0}), .out(n4936), .config_in(config_chain[6917:6915]), .config_rst(config_rst)); 
mux6 mux_2306 (.in({n11081_0, n11080_0, n11073_0/**/, n11072_0, n11067_0, n11066_1}), .out(n4937), .config_in(config_chain[6920:6918]), .config_rst(config_rst)); 
mux6 mux_2307 (.in({n13455_0/**/, n13454_0, n13443_0, n13442_0, n13429_0, n13428_1}), .out(n4938), .config_in(config_chain[6923:6921]), .config_rst(config_rst)); 
mux6 mux_2308 (.in({n11397_1, n11396_0, n11389_1, n11388_0, n11317_0, n11316_1/**/}), .out(n4939), .config_in(config_chain[6926:6924]), .config_rst(config_rst)); 
mux6 mux_2309 (.in({n13757_1, n13756_0, n13685_0, n13684_1, n13677_0/**/, n13676_1}), .out(n4940), .config_in(config_chain[6929:6927]), .config_rst(config_rst)); 
mux6 mux_2310 (.in({n11115_1, n11114_0/**/, n11101_0, n11100_0, n11043_0, n11042_1}), .out(n4941), .config_in(config_chain[6932:6930]), .config_rst(config_rst)); 
mux6 mux_2311 (.in({n13477_1, n13476_0, n13463_0, n13462_0, n13385_0/**/, n13384_1}), .out(n4942), .config_in(config_chain[6935:6933]), .config_rst(config_rst)); 
mux6 mux_2312 (.in({n11337_0, n11336_0, n11325_0, n11324_1, n11307_0/**/, n11306_1}), .out(n4943), .config_in(config_chain[6938:6936]), .config_rst(config_rst)); 
mux6 mux_2313 (.in({n13705_0, n13704_0, n13697_0, n13696_0/**/, n13647_0, n13646_1}), .out(n4944), .config_in(config_chain[6941:6939]), .config_rst(config_rst)); 
mux6 mux_2314 (.in({n11123_1, n11122_0/**/, n11053_0, n11052_1, n11045_0, n11044_1}), .out(n4945), .config_in(config_chain[6944:6942]), .config_rst(config_rst)); 
mux6 mux_2315 (.in({n13485_1, n13484_0, n13415_0/**/, n13414_1, n13389_1, n13388_1}), .out(n4946), .config_in(config_chain[6947:6945]), .config_rst(config_rst)); 
mux6 mux_2316 (.in({n11367_0, n11366_0, n11359_0, n11358_0, n11309_0, n11308_1}), .out(n4947), .config_in(config_chain[6950:6948]), .config_rst(config_rst)); 
mux6 mux_2317 (.in({n13743_1, n13742_0, n13727_0, n13726_0, n13649_0/**/, n13648_1}), .out(n4948), .config_in(config_chain[6953:6951]), .config_rst(config_rst)); 
mux6 mux_2318 (.in({n11109_1, n11108_0/**/, n11075_0, n11074_0, n11061_0, n11060_1}), .out(n4949), .config_in(config_chain[6956:6954]), .config_rst(config_rst)); 
mux6 mux_2319 (.in({n13471_1, n13470_0, n13445_0/**/, n13444_0, n13437_0, n13436_0}), .out(n4950), .config_in(config_chain[6959:6957]), .config_rst(config_rst)); 
mux6 mux_2320 (.in({n11391_1, n11390_0, n11383_1, n11382_0, n11311_0, n11310_1}), .out(n4951), .config_in(config_chain[6962:6960]), .config_rst(config_rst)); 
mux6 mux_2321 (.in({n13751_1, n13750_0, n13679_0/**/, n13678_1, n13651_0, n13650_1}), .out(n4952), .config_in(config_chain[6965:6963]), .config_rst(config_rst)); 
mux6 mux_2322 (.in({n11131_1, n11130_0/**/, n11095_0, n11094_0, n11083_0, n11082_0}), .out(n4953), .config_in(config_chain[6968:6966]), .config_rst(config_rst)); 
mux6 mux_2323 (.in({n13493_1, n13492_0, n13465_0, n13464_0, n13457_0, n13456_0/**/}), .out(n4954), .config_in(config_chain[6971:6969]), .config_rst(config_rst)); 
mux6 mux_2324 (.in({n11353_1, n11352_0, n11339_0/**/, n11338_0, n11327_0, n11326_1}), .out(n4955), .config_in(config_chain[6974:6972]), .config_rst(config_rst)); 
mux6 mux_2325 (.in({n13735_1, n13734_0, n13699_0, n13698_0, n13687_0, n13686_1/**/}), .out(n4956), .config_in(config_chain[6977:6975]), .config_rst(config_rst)); 
mux6 mux_2326 (.in({n11125_1, n11124_0/**/, n11117_1, n11116_0, n11041_0, n11040_1}), .out(n4957), .config_in(config_chain[6980:6978]), .config_rst(config_rst)); 
mux6 mux_2327 (.in({n13487_1, n13486_0, n13417_0, n13416_1/**/, n13383_0, n13382_1}), .out(n4958), .config_in(config_chain[6983:6981]), .config_rst(config_rst)); 
mux6 mux_2328 (.in({n11657_1, n11656_0, n11599_0, n11598_0, n11583_0, n11582_1}), .out(n5005), .config_in(config_chain[6986:6984]), .config_rst(config_rst)); 
mux6 mux_2329 (.in({n13773_0, n13772_0/**/, n13715_0, n13714_0, n13699_0, n13698_1}), .out(n5006), .config_in(config_chain[6989:6987]), .config_rst(config_rst)); 
mux6 mux_2330 (.in({n11377_1, n11376_0, n11369_0, n11368_0, n11361_0, n11360_0}), .out(n5007), .config_in(config_chain[6992:6990]), .config_rst(config_rst)); 
mux6 mux_2331 (.in({n13503_0, n13502_0, n13495_0, n13494_0, n13487_0, n13486_0}), .out(n5008), .config_in(config_chain[6995:6993]), .config_rst(config_rst)); 
mux6 mux_2332 (.in({n11621_0, n11620_0, n11607_0, n11606_0, n11591_0, n11590_1}), .out(n5009), .config_in(config_chain[6998:6996]), .config_rst(config_rst)); 
mux6 mux_2333 (.in({n13737_0, n13736_0, n13731_0, n13730_0, n13723_0, n13722_0}), .out(n5010), .config_in(config_chain[7001:6999]), .config_rst(config_rst)); 
mux6 mux_2334 (.in({n11393_1, n11392_0, n11321_0, n11320_1, n11313_0, n11312_1}), .out(n5011), .config_in(config_chain[7004:7002]), .config_rst(config_rst)); 
mux6 mux_2335 (.in({n13511_0, n13510_0, n13451_0, n13450_0, n13439_0, n13438_1}), .out(n5012), .config_in(config_chain[7007:7005]), .config_rst(config_rst)); 
mux6 mux_2336 (.in({n11643_1, n11642_0, n11637_0, n11636_0, n11629_0, n11628_0}), .out(n5013), .config_in(config_chain[7010:7008]), .config_rst(config_rst)); 
mux6 mux_2337 (.in({n13759_0, n13758_0, n13753_0, n13752_0, n13745_0, n13744_0}), .out(n5014), .config_in(config_chain[7013:7011]), .config_rst(config_rst)); 
mux6 mux_2338 (.in({n11341_0, n11340_0, n11333_0, n11332_0, n11329_0, n11328_1}), .out(n5015), .config_in(config_chain[7016:7014]), .config_rst(config_rst)); 
mux6 mux_2339 (.in({n13473_0, n13472_0, n13459_0, n13458_0, n13447_0, n13446_1}), .out(n5016), .config_in(config_chain[7019:7017]), .config_rst(config_rst)); 
mux6 mux_2340 (.in({n11659_1, n11658_0, n11651_1, n11650_0, n11577_0, n11576_1}), .out(n5017), .config_in(config_chain[7022:7020]), .config_rst(config_rst)); 
mux6 mux_2341 (.in({n13775_0, n13774_0, n13701_0, n13700_1/**/, n13693_0, n13692_1}), .out(n5018), .config_in(config_chain[7025:7023]), .config_rst(config_rst)); 
mux6 mux_2342 (.in({n11379_1, n11378_0, n11363_0, n11362_0, n11349_0, n11348_0}), .out(n5019), .config_in(config_chain[7028:7026]), .config_rst(config_rst)); 
mux6 mux_2343 (.in({n13497_0, n13496_0, n13489_0, n13488_0, n13481_0, n13480_0}), .out(n5020), .config_in(config_chain[7031:7029]), .config_rst(config_rst)); 
mux6 mux_2344 (.in({n11609_0, n11608_0, n11601_0, n11600_0, n11593_0, n11592_1/**/}), .out(n5021), .config_in(config_chain[7034:7032]), .config_rst(config_rst)); 
mux6 mux_2345 (.in({n13739_0, n13738_0, n13725_0, n13724_0, n13709_0, n13708_1}), .out(n5022), .config_in(config_chain[7037:7035]), .config_rst(config_rst)); 
mux6 mux_2346 (.in({n11387_1, n11386_0/**/, n11371_0, n11370_0, n11315_0, n11314_1}), .out(n5023), .config_in(config_chain[7040:7038]), .config_rst(config_rst)); 
mux6 mux_2347 (.in({n13513_0, n13512_0, n13505_0, n13504_0, n13433_0/**/, n13432_1}), .out(n5024), .config_in(config_chain[7043:7041]), .config_rst(config_rst)); 
mux6 mux_2348 (.in({n11631_0, n11630_0, n11623_0, n11622_0, n11617_0, n11616_0}), .out(n5025), .config_in(config_chain[7046:7044]), .config_rst(config_rst)); 
mux6 mux_2349 (.in({n13761_0, n13760_0, n13747_0, n13746_0, n13733_0, n13732_0/**/}), .out(n5026), .config_in(config_chain[7049:7047]), .config_rst(config_rst)); 
mux6 mux_2350 (.in({n11335_0/**/, n11334_0, n11331_0, n11330_1, n11323_0, n11322_1}), .out(n5027), .config_in(config_chain[7052:7050]), .config_rst(config_rst)); 
mux6 mux_2351 (.in({n13461_0, n13460_0, n13453_0, n13452_0, n13449_0/**/, n13448_1}), .out(n5028), .config_in(config_chain[7055:7053]), .config_rst(config_rst)); 
mux6 mux_2352 (.in({n11653_1, n11652_0, n11639_0, n11638_0/**/, n11579_0, n11578_1}), .out(n5029), .config_in(config_chain[7058:7056]), .config_rst(config_rst)); 
mux6 mux_2353 (.in({n13777_0, n13776_0, n13769_0, n13768_0, n13695_0, n13694_1}), .out(n5030), .config_in(config_chain[7061:7059]), .config_rst(config_rst)); 
mux6 mux_2354 (.in({n11365_0, n11364_0, n11357_0, n11356_0, n11351_0, n11350_0}), .out(n5031), .config_in(config_chain[7064:7062]), .config_rst(config_rst)); 
mux6 mux_2355 (.in({n13483_0, n13482_0, n13475_0, n13474_0, n13469_0, n13468_0}), .out(n5032), .config_in(config_chain[7067:7065]), .config_rst(config_rst)); 
mux6 mux_2356 (.in({n11661_1, n11660_0, n11603_0, n11602_0, n11587_0/**/, n11586_1}), .out(n5033), .config_in(config_chain[7070:7068]), .config_rst(config_rst)); 
mux6 mux_2357 (.in({n13719_0, n13718_0, n13711_0, n13710_1/**/, n13703_0, n13702_1}), .out(n5034), .config_in(config_chain[7073:7071]), .config_rst(config_rst)); 
mux6 mux_2358 (.in({n11389_1, n11388_0, n11381_1, n11380_0, n11373_0, n11372_0}), .out(n5035), .config_in(config_chain[7076:7074]), .config_rst(config_rst)); 
mux6 mux_2359 (.in({n13507_0/**/, n13506_0, n13491_0, n13490_0, n13435_0, n13434_1}), .out(n5036), .config_in(config_chain[7079:7077]), .config_rst(config_rst)); 
mux6 mux_2360 (.in({n11625_0, n11624_0, n11619_1, n11618_0, n11611_0, n11610_0}), .out(n5037), .config_in(config_chain[7082:7080]), .config_rst(config_rst)); 
mux6 mux_2361 (.in({n13749_0, n13748_0, n13741_0, n13740_0, n13735_0, n13734_0}), .out(n5038), .config_in(config_chain[7085:7083]), .config_rst(config_rst)); 
mux6 mux_2362 (.in({n11397_1, n11396_0, n11337_0, n11336_0, n11325_0, n11324_1/**/}), .out(n5039), .config_in(config_chain[7088:7086]), .config_rst(config_rst)); 
mux6 mux_2363 (.in({n13515_0, n13514_0, n13455_0/**/, n13454_0, n13443_0, n13442_1}), .out(n5040), .config_in(config_chain[7091:7089]), .config_rst(config_rst)); 
mux6 mux_2364 (.in({n11647_1, n11646_0, n11641_1, n11640_0, n11633_0, n11632_0}), .out(n5041), .config_in(config_chain[7094:7092]), .config_rst(config_rst)); 
mux6 mux_2365 (.in({n13771_0, n13770_0, n13763_0, n13762_0, n13757_0, n13756_0}), .out(n5042), .config_in(config_chain[7097:7095]), .config_rst(config_rst)); 
mux6 mux_2366 (.in({n11359_0, n11358_0, n11345_0, n11344_0/**/, n11307_0, n11306_1}), .out(n5043), .config_in(config_chain[7100:7098]), .config_rst(config_rst)); 
mux6 mux_2367 (.in({n13477_0, n13476_0, n13463_0/**/, n13462_0, n13387_0, n13386_2}), .out(n5044), .config_in(config_chain[7103:7101]), .config_rst(config_rst)); 
mux6 mux_2368 (.in({n11663_1, n11662_0, n11589_0, n11588_1, n11581_0, n11580_1}), .out(n5045), .config_in(config_chain[7106:7104]), .config_rst(config_rst)); 
mux6 mux_2369 (.in({n13779_0, n13778_0, n13721_0, n13720_0/**/, n13705_0, n13704_1}), .out(n5046), .config_in(config_chain[7109:7107]), .config_rst(config_rst)); 
mux6 mux_2370 (.in({n11383_1, n11382_0, n11367_0, n11366_0, n11311_0/**/, n11310_1}), .out(n5047), .config_in(config_chain[7112:7110]), .config_rst(config_rst)); 
mux6 mux_2371 (.in({n13509_0, n13508_0, n13501_0/**/, n13500_0, n13389_0, n13388_2}), .out(n5048), .config_in(config_chain[7115:7113]), .config_rst(config_rst)); 
mux6 mux_2372 (.in({n11613_0, n11612_0, n11605_0, n11604_0, n11573_0, n11572_1}), .out(n5049), .config_in(config_chain[7118:7116]), .config_rst(config_rst)); 
mux6 mux_2373 (.in({n13743_0, n13742_0, n13729_0, n13728_0, n13649_0, n13648_2}), .out(n5050), .config_in(config_chain[7121:7119]), .config_rst(config_rst)); 
mux6 mux_2374 (.in({n11391_1, n11390_0, n11353_1, n11352_0, n11319_0, n11318_1}), .out(n5051), .config_in(config_chain[7124:7122]), .config_rst(config_rst)); 
mux6 mux_2375 (.in({n13471_0, n13470_0, n13445_0, n13444_1, n13437_0, n13436_1}), .out(n5052), .config_in(config_chain[7127:7125]), .config_rst(config_rst)); 
mux6 mux_2376 (.in({n11649_1, n11648_0, n11635_0, n11634_0, n11575_0, n11574_1}), .out(n5053), .config_in(config_chain[7130:7128]), .config_rst(config_rst)); 
mux6 mux_2377 (.in({n13765_0, n13764_0, n13751_0, n13750_0/**/, n13713_0, n13712_1}), .out(n5054), .config_in(config_chain[7133:7131]), .config_rst(config_rst)); 
mux6 mux_2378 (.in({n11375_1, n11374_0, n11347_0, n11346_0, n11339_0, n11338_0/**/}), .out(n5055), .config_in(config_chain[7136:7134]), .config_rst(config_rst)); 
mux6 mux_2379 (.in({n13493_0, n13492_0, n13479_0, n13478_0, n13465_0, n13464_0}), .out(n5056), .config_in(config_chain[7139:7137]), .config_rst(config_rst)); 
mux6 mux_2380 (.in({n11907_1, n11906_0, n11891_0, n11890_0, n11877_0, n11876_0}), .out(n5103), .config_in(config_chain[7142:7140]), .config_rst(config_rst)); 
mux6 mux_2381 (.in({n13781_0, n13780_0, n13765_0, n13764_0, n13751_0, n13750_0}), .out(n5104), .config_in(config_chain[7145:7143]), .config_rst(config_rst)); 
mux6 mux_2382 (.in({n11599_0, n11598_0, n11591_0, n11590_1, n11583_0, n11582_1/**/}), .out(n5105), .config_in(config_chain[7148:7146]), .config_rst(config_rst)); 
mux6 mux_2383 (.in({n13481_0, n13480_0, n13473_0, n13472_0, n13465_0, n13464_1}), .out(n5106), .config_in(config_chain[7151:7149]), .config_rst(config_rst)); 
mux6 mux_2384 (.in({n11915_1, n11914_0, n11899_0, n11898_0, n11841_0, n11840_1}), .out(n5107), .config_in(config_chain[7154:7152]), .config_rst(config_rst)); 
mux6 mux_2385 (.in({n13797_0, n13796_0, n13789_0, n13788_0, n13715_0/**/, n13714_1}), .out(n5108), .config_in(config_chain[7157:7155]), .config_rst(config_rst)); 
mux6 mux_2386 (.in({n11629_0, n11628_0, n11621_0, n11620_0, n11615_0, n11614_0}), .out(n5109), .config_in(config_chain[7160:7158]), .config_rst(config_rst)); 
mux6 mux_2387 (.in({n13517_0, n13516_0, n13503_0, n13502_0, n13489_0, n13488_0/**/}), .out(n5110), .config_in(config_chain[7163:7161]), .config_rst(config_rst)); 
mux6 mux_2388 (.in({n11863_0, n11862_0, n11857_0, n11856_1, n11849_0, n11848_1}), .out(n5111), .config_in(config_chain[7166:7164]), .config_rst(config_rst)); 
mux6 mux_2389 (.in({n13737_0, n13736_0, n13731_0, n13730_1, n13723_0, n13722_1}), .out(n5112), .config_in(config_chain[7169:7167]), .config_rst(config_rst)); 
mux6 mux_2390 (.in({n11651_1, n11650_0, n11643_1, n11642_0, n11637_0, n11636_0}), .out(n5113), .config_in(config_chain[7172:7170]), .config_rst(config_rst)); 
mux6 mux_2391 (.in({n13525_0, n13524_0, n13511_0, n13510_0, n13451_0, n13450_1}), .out(n5114), .config_in(config_chain[7175:7173]), .config_rst(config_rst)); 
mux6 mux_2392 (.in({n11885_0, n11884_0, n11879_0, n11878_0, n11871_0, n11870_0}), .out(n5115), .config_in(config_chain[7178:7176]), .config_rst(config_rst)); 
mux6 mux_2393 (.in({n13767_0, n13766_0, n13759_0, n13758_0/**/, n13753_0, n13752_0}), .out(n5116), .config_in(config_chain[7181:7179]), .config_rst(config_rst)); 
mux6 mux_2394 (.in({n11659_1, n11658_0, n11601_0, n11600_0, n11585_0, n11584_1/**/}), .out(n5117), .config_in(config_chain[7184:7182]), .config_rst(config_rst)); 
mux6 mux_2395 (.in({n13475_0, n13474_0, n13467_0, n13466_1, n13459_0/**/, n13458_1}), .out(n5118), .config_in(config_chain[7187:7185]), .config_rst(config_rst)); 
mux6 mux_2396 (.in({n11917_1, n11916_0, n11909_1, n11908_0, n11901_0, n11900_0}), .out(n5119), .config_in(config_chain[7190:7188]), .config_rst(config_rst)); 
mux6 mux_2397 (.in({n13791_0, n13790_0, n13775_0, n13774_0, n13717_0, n13716_1}), .out(n5120), .config_in(config_chain[7193:7191]), .config_rst(config_rst)); 
mux6 mux_2398 (.in({n11623_0, n11622_0/**/, n11609_0, n11608_0, n11593_0, n11592_1}), .out(n5121), .config_in(config_chain[7196:7194]), .config_rst(config_rst)); 
mux6 mux_2399 (.in({n13497_0, n13496_0/**/, n13491_0, n13490_0, n13483_0, n13482_0}), .out(n5122), .config_in(config_chain[7199:7197]), .config_rst(config_rst)); 
mux6 mux_2400 (.in({n11925_1/**/, n11924_0, n11851_0, n11850_1, n11843_0, n11842_1}), .out(n5123), .config_in(config_chain[7202:7200]), .config_rst(config_rst)); 
mux6 mux_2401 (.in({n13799_0, n13798_0, n13739_0, n13738_0/**/, n13725_0, n13724_1}), .out(n5124), .config_in(config_chain[7205:7203]), .config_rst(config_rst)); 
mux6 mux_2402 (.in({n11645_1, n11644_0, n11639_0, n11638_0, n11631_0/**/, n11630_0}), .out(n5125), .config_in(config_chain[7208:7206]), .config_rst(config_rst)); 
mux6 mux_2403 (.in({n13527_0/**/, n13526_0, n13519_0, n13518_0, n13513_0, n13512_0}), .out(n5126), .config_in(config_chain[7211:7209]), .config_rst(config_rst)); 
mux6 mux_2404 (.in({n11887_0/**/, n11886_0, n11873_0, n11872_0, n11859_0, n11858_1}), .out(n5127), .config_in(config_chain[7214:7212]), .config_rst(config_rst)); 
mux6 mux_2405 (.in({n13761_0, n13760_0, n13755_0, n13754_0, n13747_0, n13746_0}), .out(n5128), .config_in(config_chain[7217:7215]), .config_rst(config_rst)); 
mux6 mux_2406 (.in({n11661_1, n11660_0, n11587_0, n11586_1/**/, n11579_0, n11578_1}), .out(n5129), .config_in(config_chain[7220:7218]), .config_rst(config_rst)); 
mux6 mux_2407 (.in({n13535_0, n13534_0, n13461_0, n13460_1, n13453_0, n13452_1}), .out(n5130), .config_in(config_chain[7223:7221]), .config_rst(config_rst)); 
mux6 mux_2408 (.in({n11911_1/**/, n11910_0, n11895_0, n11894_0, n11881_0, n11880_0}), .out(n5131), .config_in(config_chain[7226:7224]), .config_rst(config_rst)); 
mux6 mux_2409 (.in({n13785_0, n13784_0, n13777_0, n13776_0, n13769_0, n13768_0/**/}), .out(n5132), .config_in(config_chain[7229:7227]), .config_rst(config_rst)); 
mux6 mux_2410 (.in({n11611_0, n11610_0, n11603_0, n11602_0, n11595_0, n11594_1/**/}), .out(n5133), .config_in(config_chain[7232:7230]), .config_rst(config_rst)); 
mux6 mux_2411 (.in({n13499_0, n13498_0, n13485_0, n13484_0, n13469_0, n13468_1}), .out(n5134), .config_in(config_chain[7235:7233]), .config_rst(config_rst)); 
mux6 mux_2412 (.in({n11919_1, n11918_0, n11845_0, n11844_1, n11829_1, n11828_1}), .out(n5135), .config_in(config_chain[7238:7236]), .config_rst(config_rst)); 
mux6 mux_2413 (.in({n13727_0, n13726_1/**/, n13719_0, n13718_1, n13713_0, n13712_1}), .out(n5136), .config_in(config_chain[7241:7239]), .config_rst(config_rst)); 
mux6 mux_2414 (.in({n11647_1, n11646_0, n11633_0, n11632_0/**/, n11619_1, n11618_0}), .out(n5137), .config_in(config_chain[7244:7242]), .config_rst(config_rst)); 
mux6 mux_2415 (.in({n13521_0, n13520_0, n13507_0, n13506_0, n13493_0, n13492_0}), .out(n5138), .config_in(config_chain[7247:7245]), .config_rst(config_rst)); 
mux6 mux_2416 (.in({n11867_0/**/, n11866_0, n11861_1, n11860_1, n11853_0, n11852_1}), .out(n5139), .config_in(config_chain[7250:7248]), .config_rst(config_rst)); 
mux6 mux_2417 (.in({n13749_0, n13748_0, n13741_0, n13740_0, n13735_0, n13734_1/**/}), .out(n5140), .config_in(config_chain[7253:7251]), .config_rst(config_rst)); 
mux6 mux_2418 (.in({n11655_1, n11654_0, n11641_1, n11640_0, n11581_0, n11580_1}), .out(n5141), .config_in(config_chain[7256:7254]), .config_rst(config_rst)); 
mux6 mux_2419 (.in({n13537_0, n13536_0, n13529_0, n13528_0, n13455_0, n13454_1}), .out(n5142), .config_in(config_chain[7259:7257]), .config_rst(config_rst)); 
mux6 mux_2420 (.in({n11897_0, n11896_0, n11889_0, n11888_0/**/, n11883_1, n11882_0}), .out(n5143), .config_in(config_chain[7262:7260]), .config_rst(config_rst)); 
mux6 mux_2421 (.in({n13787_0, n13786_0, n13771_0, n13770_0, n13757_0, n13756_0}), .out(n5144), .config_in(config_chain[7265:7263]), .config_rst(config_rst)); 
mux6 mux_2422 (.in({n11605_0, n11604_0, n11589_0, n11588_1, n11573_0, n11572_1}), .out(n5145), .config_in(config_chain[7268:7266]), .config_rst(config_rst)); 
mux6 mux_2423 (.in({n13487_0, n13486_0, n13479_0, n13478_0, n13387_0, n13386_2}), .out(n5146), .config_in(config_chain[7271:7269]), .config_rst(config_rst)); 
mux6 mux_2424 (.in({n11921_1/**/, n11920_0, n11913_1, n11912_0, n11905_1, n11904_0}), .out(n5147), .config_in(config_chain[7274:7272]), .config_rst(config_rst)); 
mux6 mux_2425 (.in({n13795_0, n13794_0, n13779_0, n13778_0, n13721_0, n13720_1}), .out(n5148), .config_in(config_chain[7277:7275]), .config_rst(config_rst)); 
mux6 mux_2426 (.in({n11627_0, n11626_0, n11613_0, n11612_0, n11575_0, n11574_1}), .out(n5149), .config_in(config_chain[7280:7278]), .config_rst(config_rst)); 
mux6 mux_2427 (.in({n13509_0, n13508_0, n13501_0, n13500_0, n13389_0, n13388_2}), .out(n5150), .config_in(config_chain[7283:7281]), .config_rst(config_rst)); 
mux6 mux_2428 (.in({n11927_1, n11926_0, n11869_0, n11868_0, n11855_0/**/, n11854_1}), .out(n5151), .config_in(config_chain[7286:7284]), .config_rst(config_rst)); 
mux6 mux_2429 (.in({n13743_0, n13742_0, n13729_0, n13728_1, n13651_0, n13650_2}), .out(n5152), .config_in(config_chain[7289:7287]), .config_rst(config_rst)); 
mux6 mux_2430 (.in({n11657_1, n11656_0, n11649_1, n11648_0, n11597_1, n11596_1}), .out(n5153), .config_in(config_chain[7292:7290]), .config_rst(config_rst)); 
mux6 mux_2431 (.in({n13531_0, n13530_0/**/, n13471_0, n13470_1, n13457_0, n13456_1}), .out(n5154), .config_in(config_chain[7295:7293]), .config_rst(config_rst)); 
mux6 mux_2432 (.in({n12183_1, n12182_0, n12125_0, n12124_0, n12109_0, n12108_1}), .out(n5201), .config_in(config_chain[7298:7296]), .config_rst(config_rst)); 
mux6 mux_2433 (.in({n13817_0, n13816_0, n13759_0, n13758_0, n13743_0, n13742_1}), .out(n5202), .config_in(config_chain[7301:7299]), .config_rst(config_rst)); 
mux6 mux_2434 (.in({n11907_1, n11906_0, n11899_0, n11898_0, n11891_0, n11890_0}), .out(n5203), .config_in(config_chain[7304:7302]), .config_rst(config_rst)); 
mux6 mux_2435 (.in({n13547_0, n13546_0, n13539_0, n13538_0/**/, n13531_0, n13530_0}), .out(n5204), .config_in(config_chain[7307:7305]), .config_rst(config_rst)); 
mux6 mux_2436 (.in({n12147_0/**/, n12146_0, n12133_0, n12132_0, n12117_0, n12116_1}), .out(n5205), .config_in(config_chain[7310:7308]), .config_rst(config_rst)); 
mux6 mux_2437 (.in({n13781_0, n13780_0, n13775_0, n13774_0, n13767_0, n13766_0}), .out(n5206), .config_in(config_chain[7313:7311]), .config_rst(config_rst)); 
mux6 mux_2438 (.in({n11923_1, n11922_0, n11849_0, n11848_1, n11841_0, n11840_1}), .out(n5207), .config_in(config_chain[7316:7314]), .config_rst(config_rst)); 
mux6 mux_2439 (.in({n13555_0, n13554_0, n13495_0, n13494_0, n13481_0, n13480_1}), .out(n5208), .config_in(config_chain[7319:7317]), .config_rst(config_rst)); 
mux6 mux_2440 (.in({n12169_1, n12168_0, n12163_0, n12162_0, n12155_0, n12154_0}), .out(n5209), .config_in(config_chain[7322:7320]), .config_rst(config_rst)); 
mux6 mux_2441 (.in({n13803_0, n13802_0, n13797_0, n13796_0, n13789_0, n13788_0}), .out(n5210), .config_in(config_chain[7325:7323]), .config_rst(config_rst)); 
mux6 mux_2442 (.in({n11871_0, n11870_0, n11863_0, n11862_0, n11857_0, n11856_1}), .out(n5211), .config_in(config_chain[7328:7326]), .config_rst(config_rst)); 
mux6 mux_2443 (.in({n13517_0, n13516_0, n13503_0, n13502_0, n13489_0, n13488_1}), .out(n5212), .config_in(config_chain[7331:7329]), .config_rst(config_rst)); 
mux6 mux_2444 (.in({n12185_1, n12184_0, n12177_1, n12176_0, n12103_0, n12102_1}), .out(n5213), .config_in(config_chain[7334:7332]), .config_rst(config_rst)); 
mux6 mux_2445 (.in({n13819_0, n13818_0, n13745_0, n13744_1, n13737_0/**/, n13736_1}), .out(n5214), .config_in(config_chain[7337:7335]), .config_rst(config_rst)); 
mux6 mux_2446 (.in({n11909_1, n11908_0, n11893_0, n11892_0, n11879_0, n11878_0}), .out(n5215), .config_in(config_chain[7340:7338]), .config_rst(config_rst)); 
mux6 mux_2447 (.in({n13541_0, n13540_0, n13533_0, n13532_0/**/, n13525_0, n13524_0}), .out(n5216), .config_in(config_chain[7343:7341]), .config_rst(config_rst)); 
mux6 mux_2448 (.in({n12135_0, n12134_0/**/, n12127_0, n12126_0, n12119_0, n12118_1}), .out(n5217), .config_in(config_chain[7346:7344]), .config_rst(config_rst)); 
mux6 mux_2449 (.in({n13783_0, n13782_0, n13769_0, n13768_0, n13753_0, n13752_1}), .out(n5218), .config_in(config_chain[7349:7347]), .config_rst(config_rst)); 
mux6 mux_2450 (.in({n11917_1/**/, n11916_0, n11901_0, n11900_0, n11843_0, n11842_1}), .out(n5219), .config_in(config_chain[7352:7350]), .config_rst(config_rst)); 
mux6 mux_2451 (.in({n13557_0, n13556_0, n13549_0, n13548_0/**/, n13475_0, n13474_1}), .out(n5220), .config_in(config_chain[7355:7353]), .config_rst(config_rst)); 
mux6 mux_2452 (.in({n12157_0, n12156_0, n12149_0, n12148_0, n12143_0, n12142_0}), .out(n5221), .config_in(config_chain[7358:7356]), .config_rst(config_rst)); 
mux6 mux_2453 (.in({n13805_0/**/, n13804_0, n13791_0, n13790_0, n13777_0, n13776_0}), .out(n5222), .config_in(config_chain[7361:7359]), .config_rst(config_rst)); 
mux6 mux_2454 (.in({n11865_0, n11864_0, n11859_0, n11858_1/**/, n11851_0, n11850_1}), .out(n5223), .config_in(config_chain[7364:7362]), .config_rst(config_rst)); 
mux6 mux_2455 (.in({n13505_0, n13504_0, n13497_0, n13496_0, n13491_0, n13490_1}), .out(n5224), .config_in(config_chain[7367:7365]), .config_rst(config_rst)); 
mux6 mux_2456 (.in({n12179_1, n12178_0, n12165_0, n12164_0, n12105_0, n12104_1/**/}), .out(n5225), .config_in(config_chain[7370:7368]), .config_rst(config_rst)); 
mux6 mux_2457 (.in({n13821_0, n13820_0, n13813_0, n13812_0, n13739_0, n13738_1}), .out(n5226), .config_in(config_chain[7373:7371]), .config_rst(config_rst)); 
mux6 mux_2458 (.in({n11895_0/**/, n11894_0, n11887_0, n11886_0, n11881_0, n11880_0}), .out(n5227), .config_in(config_chain[7376:7374]), .config_rst(config_rst)); 
mux6 mux_2459 (.in({n13527_0, n13526_0/**/, n13519_0, n13518_0, n13513_0, n13512_0}), .out(n5228), .config_in(config_chain[7379:7377]), .config_rst(config_rst)); 
mux6 mux_2460 (.in({n12187_1, n12186_0, n12129_0, n12128_0/**/, n12113_0, n12112_1}), .out(n5229), .config_in(config_chain[7382:7380]), .config_rst(config_rst)); 
mux6 mux_2461 (.in({n13763_0, n13762_0/**/, n13755_0, n13754_1, n13747_0, n13746_1}), .out(n5230), .config_in(config_chain[7385:7383]), .config_rst(config_rst)); 
mux6 mux_2462 (.in({n11919_1, n11918_0, n11911_1, n11910_0/**/, n11903_0, n11902_0}), .out(n5231), .config_in(config_chain[7388:7386]), .config_rst(config_rst)); 
mux6 mux_2463 (.in({n13551_0, n13550_0, n13535_0, n13534_0, n13477_0, n13476_1}), .out(n5232), .config_in(config_chain[7391:7389]), .config_rst(config_rst)); 
mux6 mux_2464 (.in({n12189_1, n12188_0, n12151_0, n12150_0/**/, n12137_0, n12136_0}), .out(n5233), .config_in(config_chain[7394:7392]), .config_rst(config_rst)); 
mux6 mux_2465 (.in({n13823_0, n13822_0/**/, n13793_0, n13792_0, n13785_0, n13784_0}), .out(n5234), .config_in(config_chain[7397:7395]), .config_rst(config_rst)); 
mux6 mux_2466 (.in({n11867_0, n11866_0, n11853_0, n11852_1, n11829_1, n11828_1}), .out(n5235), .config_in(config_chain[7400:7398]), .config_rst(config_rst)); 
mux6 mux_2467 (.in({n13499_0, n13498_0/**/, n13485_0, n13484_1, n13471_0, n13470_1}), .out(n5236), .config_in(config_chain[7403:7401]), .config_rst(config_rst)); 
mux6 mux_2468 (.in({n12173_1, n12172_0, n12159_0, n12158_0, n12091_1, n12090_1}), .out(n5237), .config_in(config_chain[7406:7404]), .config_rst(config_rst)); 
mux6 mux_2469 (.in({n13815_0, n13814_0, n13807_0, n13806_0, n13713_0, n13712_1}), .out(n5238), .config_in(config_chain[7409:7407]), .config_rst(config_rst)); 
mux6 mux_2470 (.in({n11889_0, n11888_0, n11875_0, n11874_0, n11861_1, n11860_1}), .out(n5239), .config_in(config_chain[7412:7410]), .config_rst(config_rst)); 
mux6 mux_2471 (.in({n13521_0, n13520_0, n13515_0, n13514_0, n13507_0, n13506_0}), .out(n5240), .config_in(config_chain[7415:7413]), .config_rst(config_rst)); 
mux6 mux_2472 (.in({n12115_0, n12114_1, n12107_0/**/, n12106_1, n12093_1, n12092_1}), .out(n5241), .config_in(config_chain[7418:7416]), .config_rst(config_rst)); 
mux6 mux_2473 (.in({n13765_0, n13764_0, n13749_0, n13748_1, n13735_0, n13734_1}), .out(n5242), .config_in(config_chain[7421:7419]), .config_rst(config_rst)); 
mux6 mux_2474 (.in({n11913_1, n11912_0, n11905_1, n11904_0, n11897_0, n11896_0}), .out(n5243), .config_in(config_chain[7424:7422]), .config_rst(config_rst)); 
mux6 mux_2475 (.in({n13553_0, n13552_0, n13545_0, n13544_0/**/, n13537_0, n13536_0}), .out(n5244), .config_in(config_chain[7427:7425]), .config_rst(config_rst)); 
mux6 mux_2476 (.in({n12139_0, n12138_0, n12131_0, n12130_0, n12123_1, n12122_1}), .out(n5245), .config_in(config_chain[7430:7428]), .config_rst(config_rst)); 
mux6 mux_2477 (.in({n13787_0, n13786_0, n13773_0, n13772_0/**/, n13757_0, n13756_1}), .out(n5246), .config_in(config_chain[7433:7431]), .config_rst(config_rst)); 
mux6 mux_2478 (.in({n11927_1/**/, n11926_0, n11921_1, n11920_0, n11847_0, n11846_1}), .out(n5247), .config_in(config_chain[7436:7434]), .config_rst(config_rst)); 
mux6 mux_2479 (.in({n13559_0, n13558_0, n13487_0, n13486_1, n13479_0, n13478_1}), .out(n5248), .config_in(config_chain[7439:7437]), .config_rst(config_rst)); 
mux6 mux_2480 (.in({n12175_1, n12174_0, n12161_0, n12160_0/**/, n12145_1, n12144_0}), .out(n5249), .config_in(config_chain[7442:7440]), .config_rst(config_rst)); 
mux6 mux_2481 (.in({n13809_0, n13808_0, n13801_0, n13800_0, n13795_0, n13794_0}), .out(n5250), .config_in(config_chain[7445:7443]), .config_rst(config_rst)); 
mux6 mux_2482 (.in({n11877_0, n11876_0/**/, n11869_0, n11868_0, n11839_0, n11838_1}), .out(n5251), .config_in(config_chain[7448:7446]), .config_rst(config_rst)); 
mux6 mux_2483 (.in({n13523_0, n13522_0, n13509_0, n13508_0/**/, n13389_0, n13388_2}), .out(n5252), .config_in(config_chain[7451:7449]), .config_rst(config_rst)); 
mux6 mux_2484 (.in({n12133_0, n12132_0, n12125_0, n12124_0, n12117_0, n12116_1}), .out(n5298), .config_in(config_chain[7454:7452]), .config_rst(config_rst)); 
mux6 mux_2485 (.in({n12177_1, n12176_0, n12169_1, n12168_0, n12163_0, n12162_0}), .out(n5301), .config_in(config_chain[7457:7455]), .config_rst(config_rst)); 
mux6 mux_2486 (.in({n12135_0, n12134_0, n12127_0, n12126_0, n12119_0, n12118_1}), .out(n5304), .config_in(config_chain[7460:7458]), .config_rst(config_rst)); 
mux6 mux_2487 (.in({n12179_1, n12178_0, n12171_1, n12170_0, n12165_0, n12164_0}), .out(n5307), .config_in(config_chain[7463:7461]), .config_rst(config_rst)); 
mux6 mux_2488 (.in({n12129_0, n12128_0, n12121_0, n12120_1, n12113_0, n12112_1}), .out(n5310), .config_in(config_chain[7466:7464]), .config_rst(config_rst)); 
mux6 mux_2489 (.in({n12173_1, n12172_0, n12159_0, n12158_0, n12091_1, n12090_1}), .out(n5313), .config_in(config_chain[7469:7467]), .config_rst(config_rst)); 
mux6 mux_2490 (.in({n12131_0, n12130_0, n12123_1, n12122_1, n12115_0, n12114_1}), .out(n5316), .config_in(config_chain[7472:7470]), .config_rst(config_rst)); 
mux6 mux_2491 (.in({n12175_1, n12174_0/**/, n12167_1, n12166_0, n12161_0, n12160_0}), .out(n5319), .config_in(config_chain[7475:7473]), .config_rst(config_rst)); 
mux6 mux_2492 (.in({n9853_1, n9852_0, n9799_0, n9798_0, n9785_0, n9784_1}), .out(n5346), .config_in(config_chain[7478:7476]), .config_rst(config_rst)); 
mux6 mux_2493 (.in({n9827_0, n9826_0, n9819_0, n9818_0, n9815_0, n9814_0}), .out(n5349), .config_in(config_chain[7481:7479]), .config_rst(config_rst)); 
mux6 mux_2494 (.in({n9855_1, n9854_0, n9787_0, n9786_1, n9779_0, n9778_1}), .out(n5352), .config_in(config_chain[7484:7482]), .config_rst(config_rst)); 
mux6 mux_2495 (.in({n9829_0, n9828_0, n9821_0, n9820_0, n9817_0, n9816_0}), .out(n5355), .config_in(config_chain[7487:7485]), .config_rst(config_rst)); 
mux6 mux_2496 (.in({n9857_1, n9856_0, n9789_0, n9788_1, n9781_0, n9780_1}), .out(n5358), .config_in(config_chain[7490:7488]), .config_rst(config_rst)); 
mux6 mux_2497 (.in({n9823_0, n9822_0, n9811_0, n9810_0, n9749_1, n9748_1}), .out(n5361), .config_in(config_chain[7493:7491]), .config_rst(config_rst)); 
mux6 mux_2498 (.in({n9851_1, n9850_0, n9783_0, n9782_1, n9753_1, n9752_1}), .out(n5364), .config_in(config_chain[7496:7494]), .config_rst(config_rst)); 
mux6 mux_2499 (.in({n9825_0, n9824_0, n9813_0, n9812_0, n9757_1, n9756_1}), .out(n5367), .config_in(config_chain[7499:7497]), .config_rst(config_rst)); 
mux6 mux_2500 (.in({n10093_1, n10092_0, n10079_0, n10078_0, n10067_0, n10066_0}), .out(n5395), .config_in(config_chain[7502:7500]), .config_rst(config_rst)); 
mux6 mux_2501 (.in({n13881_0, n13880_0, n13851_0, n13850_0, n13829_1, n13828_0}), .out(n5396), .config_in(config_chain[7505:7503]), .config_rst(config_rst)); 
mux6 mux_2502 (.in({n9799_0, n9798_0, n9793_0, n9792_1, n9785_0, n9784_1}), .out(n5397), .config_in(config_chain[7508:7506]), .config_rst(config_rst)); 
mux6 mux_2503 (.in({n13621_0, n13620_0, n13599_0, n13598_0, n13567_0, n13566_0}), .out(n5398), .config_in(config_chain[7511:7509]), .config_rst(config_rst)); 
mux6 mux_2504 (.in({n10101_1, n10100_0, n10087_0/**/, n10086_0, n10033_0, n10032_1}), .out(n5399), .config_in(config_chain[7514:7512]), .config_rst(config_rst)); 
mux6 mux_2505 (.in({n13893_1, n13892_0, n13861_1, n13860_0, n13831_0, n13830_0}), .out(n5400), .config_in(config_chain[7517:7515]), .config_rst(config_rst)); 
mux6 mux_2506 (.in({n9827_0, n9826_0, n9819_0, n9818_0, n9815_0, n9814_0}), .out(n5401), .config_in(config_chain[7520:7518]), .config_rst(config_rst)); 
mux6 mux_2507 (.in({n13631_0, n13630_0, n13593_0, n13592_0, n13563_1, n13562_0}), .out(n5402), .config_in(config_chain[7523:7521]), .config_rst(config_rst)); 
mux6 mux_2508 (.in({n10053_0, n10052_0, n10049_0, n10048_1, n10041_0, n10040_1}), .out(n5403), .config_in(config_chain[7526:7524]), .config_rst(config_rst)); 
mux6 mux_2509 (.in({n13895_0, n13894_0, n13863_0/**/, n13862_0, n13825_0, n13824_0}), .out(n5404), .config_in(config_chain[7529:7527]), .config_rst(config_rst)); 
mux6 mux_2510 (.in({n9847_1, n9846_0, n9839_1, n9838_0, n9835_0, n9834_0}), .out(n5405), .config_in(config_chain[7532:7530]), .config_rst(config_rst)); 
mux6 mux_2511 (.in({n13625_0, n13624_0, n13595_1, n13594_0, n13565_0, n13564_0}), .out(n5406), .config_in(config_chain[7535:7533]), .config_rst(config_rst)); 
mux6 mux_2512 (.in({n10073_0, n10072_0, n10069_0, n10068_0, n10061_0/**/, n10060_0}), .out(n5407), .config_in(config_chain[7538:7536]), .config_rst(config_rst)); 
mux6 mux_2513 (.in({n13889_0, n13888_0, n13859_0, n13858_0, n13827_0, n13826_0}), .out(n5408), .config_in(config_chain[7541:7539]), .config_rst(config_rst)); 
mux6 mux_2514 (.in({n9855_1, n9854_0, n9801_0, n9800_0, n9787_0/**/, n9786_1}), .out(n5409), .config_in(config_chain[7544:7542]), .config_rst(config_rst)); 
mux6 mux_2515 (.in({n13629_0/**/, n13628_0, n13597_0, n13596_0, n13575_0, n13574_0}), .out(n5410), .config_in(config_chain[7547:7545]), .config_rst(config_rst)); 
mux6 mux_2516 (.in({n10103_1, n10102_0, n10095_1/**/, n10094_0, n10089_0, n10088_0}), .out(n5411), .config_in(config_chain[7550:7548]), .config_rst(config_rst)); 
mux6 mux_2517 (.in({n13891_0, n13890_0, n13869_1, n13868_0, n13839_0/**/, n13838_0}), .out(n5412), .config_in(config_chain[7553:7551]), .config_rst(config_rst)); 
mux6 mux_2518 (.in({n9821_0, n9820_0/**/, n9809_0, n9808_0, n9795_0, n9794_1}), .out(n5413), .config_in(config_chain[7556:7554]), .config_rst(config_rst)); 
mux6 mux_2519 (.in({n13639_0, n13638_0, n13607_0, n13606_0, n13569_0, n13568_0}), .out(n5414), .config_in(config_chain[7559:7557]), .config_rst(config_rst)); 
mux6 mux_2520 (.in({n10111_1, n10110_0, n10043_0/**/, n10042_1, n10035_0, n10034_1}), .out(n5415), .config_in(config_chain[7562:7560]), .config_rst(config_rst)); 
mux6 mux_2521 (.in({n13901_1, n13900_0, n13871_0, n13870_0, n13833_0, n13832_0}), .out(n5416), .config_in(config_chain[7565:7563]), .config_rst(config_rst)); 
mux6 mux_2522 (.in({n9841_1, n9840_0, n9837_0, n9836_0, n9829_0/**/, n9828_0}), .out(n5417), .config_in(config_chain[7568:7566]), .config_rst(config_rst)); 
mux6 mux_2523 (.in({n13633_0, n13632_0, n13603_1, n13602_0, n13571_1/**/, n13570_0}), .out(n5418), .config_in(config_chain[7571:7569]), .config_rst(config_rst)); 
mux6 mux_2524 (.in({n10075_0, n10074_0, n10063_0, n10062_0, n10051_0, n10050_1}), .out(n5419), .config_in(config_chain[7574:7572]), .config_rst(config_rst)); 
mux6 mux_2525 (.in({n13897_0, n13896_0, n13865_0, n13864_0, n13835_0/**/, n13834_0}), .out(n5420), .config_in(config_chain[7577:7575]), .config_rst(config_rst)); 
mux6 mux_2526 (.in({n9857_1, n9856_0, n9789_0, n9788_1, n9781_0, n9780_1}), .out(n5421), .config_in(config_chain[7580:7578]), .config_rst(config_rst)); 
mux6 mux_2527 (.in({n13635_1, n13634_0, n13605_0/**/, n13604_0, n13573_0, n13572_0}), .out(n5422), .config_in(config_chain[7583:7581]), .config_rst(config_rst)); 
mux6 mux_2528 (.in({n10097_1, n10096_0, n10083_0, n10082_0, n10071_0, n10070_0/**/}), .out(n5423), .config_in(config_chain[7586:7584]), .config_rst(config_rst)); 
mux6 mux_2529 (.in({n13899_0, n13898_0, n13867_0, n13866_0, n13845_1/**/, n13844_0}), .out(n5424), .config_in(config_chain[7589:7587]), .config_rst(config_rst)); 
mux6 mux_2530 (.in({n9811_0, n9810_0, n9803_0, n9802_0, n9797_0, n9796_1}), .out(n5425), .config_in(config_chain[7592:7590]), .config_rst(config_rst)); 
mux6 mux_2531 (.in({n13637_0, n13636_0, n13615_0/**/, n13614_0, n13577_0, n13576_0}), .out(n5426), .config_in(config_chain[7595:7593]), .config_rst(config_rst)); 
mux6 mux_2532 (.in({n10105_1/**/, n10104_0, n10037_0, n10036_1, n10001_0, n10000_1}), .out(n5427), .config_in(config_chain[7598:7596]), .config_rst(config_rst)); 
mux6 mux_2533 (.in({n13905_0, n13904_0, n13879_0, n13878_0, n13847_0, n13846_0}), .out(n5428), .config_in(config_chain[7601:7599]), .config_rst(config_rst)); 
mux6 mux_2534 (.in({n9843_1, n9842_0, n9831_0, n9830_0/**/, n9749_1, n9748_1}), .out(n5429), .config_in(config_chain[7604:7602]), .config_rst(config_rst)); 
mux6 mux_2535 (.in({n13643_1, n13642_0, n13609_0, n13608_0, n13579_1, n13578_0}), .out(n5430), .config_in(config_chain[7607:7605]), .config_rst(config_rst)); 
mux6 mux_2536 (.in({n10057_0, n10056_0, n10045_0/**/, n10044_1, n10003_0, n10002_1}), .out(n5431), .config_in(config_chain[7610:7608]), .config_rst(config_rst)); 
mux6 mux_2537 (.in({n13907_0, n13906_0, n13873_0, n13872_0, n13841_0, n13840_0}), .out(n5432), .config_in(config_chain[7613:7611]), .config_rst(config_rst)); 
mux6 mux_2538 (.in({n9851_1, n9850_0, n9783_0, n9782_1, n9751_1, n9750_1}), .out(n5433), .config_in(config_chain[7616:7614]), .config_rst(config_rst)); 
mux6 mux_2539 (.in({n13647_1, n13646_0, n13611_1, n13610_0, n13581_0, n13580_0}), .out(n5434), .config_in(config_chain[7619:7617]), .config_rst(config_rst)); 
mux6 mux_2540 (.in({n10085_0, n10084_0/**/, n10077_0, n10076_0, n10005_1, n10004_1}), .out(n5435), .config_in(config_chain[7622:7620]), .config_rst(config_rst)); 
mux6 mux_2541 (.in({n13909_1, n13908_0, n13875_0, n13874_0, n13853_1/**/, n13852_0}), .out(n5436), .config_in(config_chain[7625:7623]), .config_rst(config_rst)); 
mux6 mux_2542 (.in({n9805_0, n9804_0, n9791_0/**/, n9790_1, n9755_1, n9754_1}), .out(n5437), .config_in(config_chain[7628:7626]), .config_rst(config_rst)); 
mux6 mux_2543 (.in({n13649_2, n13648_0, n13623_0, n13622_0, n13591_0, n13590_0}), .out(n5438), .config_in(config_chain[7631:7629]), .config_rst(config_rst)); 
mux6 mux_2544 (.in({n10107_1, n10106_0, n10099_1, n10098_0, n10007_1, n10006_1}), .out(n5439), .config_in(config_chain[7634:7632]), .config_rst(config_rst)); 
mux6 mux_2545 (.in({n13911_1, n13910_0, n13885_1, n13884_0/**/, n13855_0, n13854_0}), .out(n5440), .config_in(config_chain[7637:7635]), .config_rst(config_rst)); 
mux6 mux_2546 (.in({n9825_0, n9824_0, n9813_0, n9812_0, n9757_1, n9756_1}), .out(n5441), .config_in(config_chain[7640:7638]), .config_rst(config_rst)); 
mux6 mux_2547 (.in({n13651_2, n13650_0, n13617_0, n13616_0/**/, n13585_0, n13584_0}), .out(n5442), .config_in(config_chain[7643:7641]), .config_rst(config_rst)); 
mux6 mux_2548 (.in({n10059_0, n10058_0, n10047_0/**/, n10046_1, n10009_1, n10008_1}), .out(n5443), .config_in(config_chain[7646:7644]), .config_rst(config_rst)); 
mux6 mux_2549 (.in({n13915_2, n13914_0, n13887_0, n13886_0, n13849_0, n13848_0}), .out(n5444), .config_in(config_chain[7649:7647]), .config_rst(config_rst)); 
mux6 mux_2550 (.in({n9853_1, n9852_0, n9845_1, n9844_0, n9747_0, n9746_1}), .out(n5445), .config_in(config_chain[7652:7650]), .config_rst(config_rst)); 
mux6 mux_2551 (.in({n13641_0, n13640_0, n13619_1, n13618_0, n13589_0, n13588_0/**/}), .out(n5446), .config_in(config_chain[7655:7653]), .config_rst(config_rst)); 
mux6 mux_2552 (.in({n10363_1, n10362_0, n10309_0, n10308_0, n10295_0, n10294_1}), .out(n5493), .config_in(config_chain[7658:7656]), .config_rst(config_rst)); 
mux6 mux_2553 (.in({n13931_1, n13930_0, n13849_0, n13848_0, n13827_0, n13826_0}), .out(n5494), .config_in(config_chain[7661:7659]), .config_rst(config_rst)); 
mux6 mux_2554 (.in({n10093_1, n10092_0, n10087_0, n10086_0, n10079_0, n10078_0}), .out(n5495), .config_in(config_chain[7664:7662]), .config_rst(config_rst)); 
mux6 mux_2555 (.in({n13661_1, n13660_0, n13653_1, n13652_0/**/, n13619_0, n13618_0}), .out(n5496), .config_in(config_chain[7667:7665]), .config_rst(config_rst)); 
mux6 mux_2556 (.in({n10329_0, n10328_0, n10317_0, n10316_0, n10303_0, n10302_1}), .out(n5497), .config_in(config_chain[7670:7668]), .config_rst(config_rst)); 
mux6 mux_2557 (.in({n13891_0, n13890_0, n13859_0, n13858_0, n13829_0, n13828_0}), .out(n5498), .config_in(config_chain[7673:7671]), .config_rst(config_rst)); 
mux6 mux_2558 (.in({n10109_1, n10108_0, n10041_0, n10040_1, n10033_0, n10032_1}), .out(n5499), .config_in(config_chain[7676:7674]), .config_rst(config_rst)); 
mux6 mux_2559 (.in({n13669_1, n13668_0, n13599_0, n13598_0, n13561_0, n13560_0}), .out(n5500), .config_in(config_chain[7679:7677]), .config_rst(config_rst)); 
mux6 mux_2560 (.in({n10349_1, n10348_0, n10345_0, n10344_0, n10337_0, n10336_0}), .out(n5501), .config_in(config_chain[7682:7680]), .config_rst(config_rst)); 
mux6 mux_2561 (.in({n13917_1, n13916_0, n13893_0, n13892_0, n13861_0, n13860_0}), .out(n5502), .config_in(config_chain[7685:7683]), .config_rst(config_rst)); 
mux6 mux_2562 (.in({n10061_0, n10060_0/**/, n10053_0, n10052_0, n10049_0, n10048_1}), .out(n5503), .config_in(config_chain[7688:7686]), .config_rst(config_rst)); 
mux6 mux_2563 (.in({n13631_0, n13630_0, n13593_0/**/, n13592_0, n13563_0, n13562_0}), .out(n5504), .config_in(config_chain[7691:7689]), .config_rst(config_rst)); 
mux6 mux_2564 (.in({n10365_1, n10364_0, n10357_1, n10356_0, n10289_0, n10288_1}), .out(n5505), .config_in(config_chain[7694:7692]), .config_rst(config_rst)); 
mux6 mux_2565 (.in({n13933_1, n13932_0, n13857_0, n13856_0, n13825_0, n13824_0/**/}), .out(n5506), .config_in(config_chain[7697:7695]), .config_rst(config_rst)); 
mux6 mux_2566 (.in({n10095_1/**/, n10094_0, n10081_0, n10080_0, n10069_0, n10068_0}), .out(n5507), .config_in(config_chain[7700:7698]), .config_rst(config_rst)); 
mux6 mux_2567 (.in({n13655_1, n13654_0, n13627_0, n13626_0, n13595_0, n13594_0}), .out(n5508), .config_in(config_chain[7703:7701]), .config_rst(config_rst)); 
mux6 mux_2568 (.in({n10319_0/**/, n10318_0, n10311_0, n10310_0, n10305_0, n10304_1}), .out(n5509), .config_in(config_chain[7706:7704]), .config_rst(config_rst)); 
mux6 mux_2569 (.in({n13889_0, n13888_0, n13867_0/**/, n13866_0, n13837_0, n13836_0}), .out(n5510), .config_in(config_chain[7709:7707]), .config_rst(config_rst)); 
mux6 mux_2570 (.in({n10103_1, n10102_0, n10089_0, n10088_0, n10035_0, n10034_1/**/}), .out(n5511), .config_in(config_chain[7712:7710]), .config_rst(config_rst)); 
mux6 mux_2571 (.in({n13671_1, n13670_0, n13663_1, n13662_0, n13575_0/**/, n13574_0}), .out(n5512), .config_in(config_chain[7715:7713]), .config_rst(config_rst)); 
mux6 mux_2572 (.in({n10339_0, n10338_0, n10331_0, n10330_0, n10327_0/**/, n10326_0}), .out(n5513), .config_in(config_chain[7718:7716]), .config_rst(config_rst)); 
mux6 mux_2573 (.in({n13919_1, n13918_0, n13899_0, n13898_0, n13869_0, n13868_0}), .out(n5514), .config_in(config_chain[7721:7719]), .config_rst(config_rst)); 
mux6 mux_2574 (.in({n10055_0, n10054_0/**/, n10051_0, n10050_1, n10043_0, n10042_1}), .out(n5515), .config_in(config_chain[7724:7722]), .config_rst(config_rst)); 
mux6 mux_2575 (.in({n13639_0/**/, n13638_0, n13601_0, n13600_0, n13569_0, n13568_0}), .out(n5516), .config_in(config_chain[7727:7725]), .config_rst(config_rst)); 
mux6 mux_2576 (.in({n10359_1, n10358_0, n10347_0, n10346_0, n10291_0, n10290_1}), .out(n5517), .config_in(config_chain[7730:7728]), .config_rst(config_rst)); 
mux6 mux_2577 (.in({n13935_1, n13934_0, n13927_1, n13926_0, n13833_0/**/, n13832_0}), .out(n5518), .config_in(config_chain[7733:7731]), .config_rst(config_rst)); 
mux6 mux_2578 (.in({n10083_0, n10082_0/**/, n10075_0, n10074_0, n10071_0, n10070_0}), .out(n5519), .config_in(config_chain[7736:7734]), .config_rst(config_rst)); 
mux6 mux_2579 (.in({n13633_0, n13632_0/**/, n13603_0, n13602_0, n13571_0, n13570_0}), .out(n5520), .config_in(config_chain[7739:7737]), .config_rst(config_rst)); 
mux6 mux_2580 (.in({n10367_1, n10366_0/**/, n10313_0, n10312_0, n10299_0, n10298_1}), .out(n5521), .config_in(config_chain[7742:7740]), .config_rst(config_rst)); 
mux6 mux_2581 (.in({n13897_0, n13896_0, n13865_0, n13864_0, n13843_0, n13842_0}), .out(n5522), .config_in(config_chain[7745:7743]), .config_rst(config_rst)); 
mux6 mux_2582 (.in({n10105_1, n10104_0, n10097_1, n10096_0, n10091_0, n10090_0}), .out(n5523), .config_in(config_chain[7748:7746]), .config_rst(config_rst)); 
mux6 mux_2583 (.in({n13665_1, n13664_0, n13635_0, n13634_0, n13583_0, n13582_0}), .out(n5524), .config_in(config_chain[7751:7749]), .config_rst(config_rst)); 
mux6 mux_2584 (.in({n10333_0, n10332_0/**/, n10321_0, n10320_0, n10267_1, n10266_1}), .out(n5525), .config_in(config_chain[7754:7752]), .config_rst(config_rst)); 
mux6 mux_2585 (.in({n13915_1, n13914_0, n13877_0, n13876_0, n13845_0, n13844_0}), .out(n5526), .config_in(config_chain[7757:7755]), .config_rst(config_rst)); 
mux6 mux_2586 (.in({n10057_0, n10056_0, n10045_0, n10044_1, n10001_0/**/, n10000_1}), .out(n5527), .config_in(config_chain[7760:7758]), .config_rst(config_rst)); 
mux6 mux_2587 (.in({n13641_0, n13640_0, n13615_0, n13614_0, n13577_0, n13576_0/**/}), .out(n5528), .config_in(config_chain[7763:7761]), .config_rst(config_rst)); 
mux6 mux_2588 (.in({n10353_1, n10352_0, n10341_0, n10340_0, n10257_0, n10256_1}), .out(n5529), .config_in(config_chain[7766:7764]), .config_rst(config_rst)); 
mux6 mux_2589 (.in({n13929_1/**/, n13928_0, n13921_1, n13920_0, n13905_0, n13904_0}), .out(n5530), .config_in(config_chain[7769:7767]), .config_rst(config_rst)); 
mux6 mux_2590 (.in({n10077_0, n10076_0, n10065_0, n10064_0/**/, n10003_0, n10002_1}), .out(n5531), .config_in(config_chain[7772:7770]), .config_rst(config_rst)); 
mux6 mux_2591 (.in({n13645_1, n13644_0, n13609_0/**/, n13608_0, n13579_0, n13578_0}), .out(n5532), .config_in(config_chain[7775:7773]), .config_rst(config_rst)); 
mux6 mux_2592 (.in({n10301_0, n10300_1, n10293_0, n10292_1/**/, n10259_0, n10258_1}), .out(n5533), .config_in(config_chain[7778:7776]), .config_rst(config_rst)); 
mux6 mux_2593 (.in({n13907_0, n13906_0, n13873_0, n13872_0, n13851_0, n13850_0}), .out(n5534), .config_in(config_chain[7781:7779]), .config_rst(config_rst)); 
mux6 mux_2594 (.in({n10099_1/**/, n10098_0, n10085_0, n10084_0, n10007_1, n10006_1}), .out(n5535), .config_in(config_chain[7784:7782]), .config_rst(config_rst)); 
mux6 mux_2595 (.in({n13667_1, n13666_0, n13659_1, n13658_0/**/, n13647_1, n13646_0}), .out(n5536), .config_in(config_chain[7787:7785]), .config_rst(config_rst)); 
mux6 mux_2596 (.in({n10323_0, n10322_0, n10315_0, n10314_0, n10261_0, n10260_1}), .out(n5537), .config_in(config_chain[7790:7788]), .config_rst(config_rst)); 
mux6 mux_2597 (.in({n13909_0, n13908_0, n13883_0, n13882_0/**/, n13853_0, n13852_0}), .out(n5538), .config_in(config_chain[7793:7791]), .config_rst(config_rst)); 
mux6 mux_2598 (.in({n10107_1/**/, n10106_0, n10039_0, n10038_1, n10009_1, n10008_1}), .out(n5539), .config_in(config_chain[7796:7794]), .config_rst(config_rst)); 
mux6 mux_2599 (.in({n13649_1, n13648_0, n13623_0/**/, n13622_0, n13591_0, n13590_0}), .out(n5540), .config_in(config_chain[7799:7797]), .config_rst(config_rst)); 
mux6 mux_2600 (.in({n10355_1, n10354_0, n10343_0, n10342_0, n10263_1, n10262_1}), .out(n5541), .config_in(config_chain[7802:7800]), .config_rst(config_rst)); 
mux6 mux_2601 (.in({n13923_1, n13922_0, n13913_1, n13912_0, n13885_0/**/, n13884_0}), .out(n5542), .config_in(config_chain[7805:7803]), .config_rst(config_rst)); 
mux6 mux_2602 (.in({n10067_0, n10066_0, n10059_0/**/, n10058_0, n10011_1, n10010_1}), .out(n5543), .config_in(config_chain[7808:7806]), .config_rst(config_rst)); 
mux6 mux_2603 (.in({n13651_2, n13650_0, n13617_0, n13616_0/**/, n13587_0, n13586_0}), .out(n5544), .config_in(config_chain[7811:7809]), .config_rst(config_rst)); 
mux6 mux_2604 (.in({n10607_1/**/, n10606_0, n10593_0, n10592_0, n10581_0, n10580_0}), .out(n5591), .config_in(config_chain[7814:7812]), .config_rst(config_rst)); 
mux6 mux_2605 (.in({n13937_1, n13936_0, n13923_0, n13922_0, n13885_0, n13884_0}), .out(n5592), .config_in(config_chain[7817:7815]), .config_rst(config_rst)); 
mux6 mux_2606 (.in({n10309_0, n10308_0, n10303_0, n10302_1, n10295_0/**/, n10294_1}), .out(n5593), .config_in(config_chain[7820:7818]), .config_rst(config_rst)); 
mux6 mux_2607 (.in({n13617_0, n13616_0, n13595_0, n13594_0, n13563_0, n13562_0}), .out(n5594), .config_in(config_chain[7823:7821]), .config_rst(config_rst)); 
mux6 mux_2608 (.in({n10615_1, n10614_0, n10601_0, n10600_0, n10547_0, n10546_1}), .out(n5595), .config_in(config_chain[7826:7824]), .config_rst(config_rst)); 
mux6 mux_2609 (.in({n13953_1, n13952_0, n13945_1, n13944_0, n13827_0, n13826_0}), .out(n5596), .config_in(config_chain[7829:7827]), .config_rst(config_rst)); 
mux6 mux_2610 (.in({n10337_0, n10336_0, n10329_0, n10328_0, n10325_0, n10324_0}), .out(n5597), .config_in(config_chain[7832:7830]), .config_rst(config_rst)); 
mux6 mux_2611 (.in({n13673_1, n13672_0, n13661_0, n13660_0, n13627_0, n13626_0}), .out(n5598), .config_in(config_chain[7835:7833]), .config_rst(config_rst)); 
mux6 mux_2612 (.in({n10567_0, n10566_0, n10563_0, n10562_1, n10555_0, n10554_1}), .out(n5599), .config_in(config_chain[7838:7836]), .config_rst(config_rst)); 
mux6 mux_2613 (.in({n13891_0, n13890_0, n13859_0, n13858_0, n13829_0, n13828_0}), .out(n5600), .config_in(config_chain[7841:7839]), .config_rst(config_rst)); 
mux6 mux_2614 (.in({n10357_1, n10356_0/**/, n10349_1, n10348_0, n10345_0, n10344_0}), .out(n5601), .config_in(config_chain[7844:7842]), .config_rst(config_rst)); 
mux6 mux_2615 (.in({n13681_1, n13680_0, n13669_0, n13668_0, n13561_0, n13560_0}), .out(n5602), .config_in(config_chain[7847:7845]), .config_rst(config_rst)); 
mux6 mux_2616 (.in({n10587_0, n10586_0, n10583_0, n10582_0, n10575_0, n10574_0}), .out(n5603), .config_in(config_chain[7850:7848]), .config_rst(config_rst)); 
mux6 mux_2617 (.in({n13925_0/**/, n13924_0, n13917_0, n13916_0, n13893_0, n13892_0}), .out(n5604), .config_in(config_chain[7853:7851]), .config_rst(config_rst)); 
mux6 mux_2618 (.in({n10365_1, n10364_0/**/, n10311_0, n10310_0, n10297_0, n10296_1}), .out(n5605), .config_in(config_chain[7856:7854]), .config_rst(config_rst)); 
mux6 mux_2619 (.in({n13625_0, n13624_0, n13593_0, n13592_0, n13571_0, n13570_0}), .out(n5606), .config_in(config_chain[7859:7857]), .config_rst(config_rst)); 
mux6 mux_2620 (.in({n10617_1, n10616_0, n10609_1, n10608_0, n10603_0, n10602_0}), .out(n5607), .config_in(config_chain[7862:7860]), .config_rst(config_rst)); 
mux6 mux_2621 (.in({n13947_1, n13946_0, n13933_0, n13932_0, n13835_0, n13834_0}), .out(n5608), .config_in(config_chain[7865:7863]), .config_rst(config_rst)); 
mux6 mux_2622 (.in({n10331_0/**/, n10330_0, n10319_0, n10318_0, n10305_0, n10304_1}), .out(n5609), .config_in(config_chain[7868:7866]), .config_rst(config_rst)); 
mux6 mux_2623 (.in({n13655_0, n13654_0/**/, n13635_0, n13634_0, n13603_0, n13602_0}), .out(n5610), .config_in(config_chain[7871:7869]), .config_rst(config_rst)); 
mux6 mux_2624 (.in({n10625_1, n10624_0, n10557_0, n10556_1, n10549_0, n10548_1}), .out(n5611), .config_in(config_chain[7874:7872]), .config_rst(config_rst)); 
mux6 mux_2625 (.in({n13955_1, n13954_0, n13867_0, n13866_0, n13837_0, n13836_0}), .out(n5612), .config_in(config_chain[7877:7875]), .config_rst(config_rst)); 
mux6 mux_2626 (.in({n10351_1, n10350_0, n10347_0, n10346_0/**/, n10339_0, n10338_0}), .out(n5613), .config_in(config_chain[7880:7878]), .config_rst(config_rst)); 
mux6 mux_2627 (.in({n13683_1/**/, n13682_0, n13675_1, n13674_0, n13671_0, n13670_0}), .out(n5614), .config_in(config_chain[7883:7881]), .config_rst(config_rst)); 
mux6 mux_2628 (.in({n10589_0, n10588_0, n10577_0, n10576_0, n10565_0, n10564_1/**/}), .out(n5615), .config_in(config_chain[7886:7884]), .config_rst(config_rst)); 
mux6 mux_2629 (.in({n13919_0, n13918_0, n13901_0/**/, n13900_0, n13869_0, n13868_0}), .out(n5616), .config_in(config_chain[7889:7887]), .config_rst(config_rst)); 
mux6 mux_2630 (.in({n10367_1, n10366_0, n10299_0, n10298_1/**/, n10291_0, n10290_1}), .out(n5617), .config_in(config_chain[7892:7890]), .config_rst(config_rst)); 
mux6 mux_2631 (.in({n13691_1, n13690_0, n13601_0, n13600_0, n13569_0/**/, n13568_0}), .out(n5618), .config_in(config_chain[7895:7893]), .config_rst(config_rst)); 
mux6 mux_2632 (.in({n10611_1/**/, n10610_0, n10597_0, n10596_0, n10585_0, n10584_0}), .out(n5619), .config_in(config_chain[7898:7896]), .config_rst(config_rst)); 
mux6 mux_2633 (.in({n13941_1, n13940_0/**/, n13935_0, n13934_0, n13927_0, n13926_0}), .out(n5620), .config_in(config_chain[7901:7899]), .config_rst(config_rst)); 
mux6 mux_2634 (.in({n10321_0, n10320_0/**/, n10313_0, n10312_0, n10307_0, n10306_1}), .out(n5621), .config_in(config_chain[7904:7902]), .config_rst(config_rst)); 
mux6 mux_2635 (.in({n13657_0, n13656_0, n13633_0/**/, n13632_0, n13611_0, n13610_0}), .out(n5622), .config_in(config_chain[7907:7905]), .config_rst(config_rst)); 
mux6 mux_2636 (.in({n10619_1, n10618_0, n10551_0, n10550_1, n10523_1, n10522_1}), .out(n5623), .config_in(config_chain[7910:7908]), .config_rst(config_rst)); 
mux6 mux_2637 (.in({n13913_1, n13912_0, n13875_0, n13874_0, n13843_0, n13842_0}), .out(n5624), .config_in(config_chain[7913:7911]), .config_rst(config_rst)); 
mux6 mux_2638 (.in({n10353_1, n10352_0, n10341_0, n10340_0, n10267_1, n10266_1}), .out(n5625), .config_in(config_chain[7916:7914]), .config_rst(config_rst)); 
mux6 mux_2639 (.in({n13677_1, n13676_0, n13665_0/**/, n13664_0, n13651_1, n13650_0}), .out(n5626), .config_in(config_chain[7919:7917]), .config_rst(config_rst)); 
mux6 mux_2640 (.in({n10571_0, n10570_0, n10559_0, n10558_1, n10525_1, n10524_1}), .out(n5627), .config_in(config_chain[7922:7920]), .config_rst(config_rst)); 
mux6 mux_2641 (.in({n13915_1, n13914_0, n13877_0, n13876_0, n13845_0, n13844_0}), .out(n5628), .config_in(config_chain[7925:7923]), .config_rst(config_rst)); 
mux6 mux_2642 (.in({n10361_1, n10360_0, n10293_0, n10292_1, n10257_0, n10256_1}), .out(n5629), .config_in(config_chain[7928:7926]), .config_rst(config_rst)); 
mux6 mux_2643 (.in({n13685_1, n13684_0, n13643_0, n13642_0, n13577_0, n13576_0/**/}), .out(n5630), .config_in(config_chain[7931:7929]), .config_rst(config_rst)); 
mux6 mux_2644 (.in({n10627_1, n10626_0, n10599_0/**/, n10598_0, n10591_0, n10590_0}), .out(n5631), .config_in(config_chain[7934:7932]), .config_rst(config_rst)); 
mux6 mux_2645 (.in({n13957_2, n13956_0, n13943_1, n13942_0, n13929_0, n13928_0}), .out(n5632), .config_in(config_chain[7937:7935]), .config_rst(config_rst)); 
mux6 mux_2646 (.in({n10315_0/**/, n10314_0, n10301_0, n10300_1, n10261_0, n10260_1}), .out(n5633), .config_in(config_chain[7940:7938]), .config_rst(config_rst)); 
mux6 mux_2647 (.in({n13645_0, n13644_0, n13619_0/**/, n13618_0, n13587_0, n13586_0}), .out(n5634), .config_in(config_chain[7943:7941]), .config_rst(config_rst)); 
mux6 mux_2648 (.in({n10621_1, n10620_0, n10613_1/**/, n10612_0, n10517_0, n10516_1}), .out(n5635), .config_in(config_chain[7946:7944]), .config_rst(config_rst)); 
mux6 mux_2649 (.in({n13951_1, n13950_0, n13907_0, n13906_0, n13851_0, n13850_0/**/}), .out(n5636), .config_in(config_chain[7949:7947]), .config_rst(config_rst)); 
mux6 mux_2650 (.in({n10335_0, n10334_0/**/, n10323_0, n10322_0, n10263_1, n10262_1}), .out(n5637), .config_in(config_chain[7952:7950]), .config_rst(config_rst)); 
mux6 mux_2651 (.in({n13667_0, n13666_0, n13659_0, n13658_0, n13647_1, n13646_0}), .out(n5638), .config_in(config_chain[7955:7953]), .config_rst(config_rst)); 
mux6 mux_2652 (.in({n10573_0, n10572_0, n10561_0, n10560_1/**/, n10519_0, n10518_1}), .out(n5639), .config_in(config_chain[7958:7956]), .config_rst(config_rst)); 
mux6 mux_2653 (.in({n13911_0, n13910_0/**/, n13883_0, n13882_0, n13853_0, n13852_0}), .out(n5640), .config_in(config_chain[7961:7959]), .config_rst(config_rst)); 
mux6 mux_2654 (.in({n10363_1, n10362_0, n10355_1/**/, n10354_0, n10265_1, n10264_1}), .out(n5641), .config_in(config_chain[7964:7962]), .config_rst(config_rst)); 
mux6 mux_2655 (.in({n13687_1/**/, n13686_0, n13649_1, n13648_0, n13585_0, n13584_0}), .out(n5642), .config_in(config_chain[7967:7965]), .config_rst(config_rst)); 
mux6 mux_2656 (.in({n10883_1, n10882_0, n10827_0, n10826_0/**/, n10813_0, n10812_1}), .out(n5689), .config_in(config_chain[7970:7968]), .config_rst(config_rst)); 
mux6 mux_2657 (.in({n13973_1, n13972_0, n13917_0/**/, n13916_0, n13853_0, n13852_1}), .out(n5690), .config_in(config_chain[7973:7971]), .config_rst(config_rst)); 
mux6 mux_2658 (.in({n10607_1, n10606_0/**/, n10601_0, n10600_0, n10593_0, n10592_0}), .out(n5691), .config_in(config_chain[7976:7974]), .config_rst(config_rst)); 
mux6 mux_2659 (.in({n13701_1, n13700_0, n13693_1/**/, n13692_0, n13687_0, n13686_0}), .out(n5692), .config_in(config_chain[7979:7977]), .config_rst(config_rst)); 
mux6 mux_2660 (.in({n10847_0, n10846_0, n10835_0, n10834_0, n10821_0, n10820_1}), .out(n5693), .config_in(config_chain[7982:7980]), .config_rst(config_rst)); 
mux6 mux_2661 (.in({n13937_0, n13936_0, n13933_0, n13932_0, n13925_0, n13924_0}), .out(n5694), .config_in(config_chain[7985:7983]), .config_rst(config_rst)); 
mux6 mux_2662 (.in({n10623_1, n10622_0, n10555_0, n10554_1, n10547_0, n10546_1}), .out(n5695), .config_in(config_chain[7988:7986]), .config_rst(config_rst)); 
mux6 mux_2663 (.in({n13709_1, n13708_0, n13653_0, n13652_0, n13595_0, n13594_1}), .out(n5696), .config_in(config_chain[7991:7989]), .config_rst(config_rst)); 
mux6 mux_2664 (.in({n10869_1, n10868_0, n10863_0/**/, n10862_0, n10855_0, n10854_0}), .out(n5697), .config_in(config_chain[7994:7992]), .config_rst(config_rst)); 
mux6 mux_2665 (.in({n13959_1, n13958_0, n13953_0, n13952_0, n13945_0, n13944_0}), .out(n5698), .config_in(config_chain[7997:7995]), .config_rst(config_rst)); 
mux6 mux_2666 (.in({n10575_0, n10574_0, n10567_0, n10566_0, n10563_0, n10562_1}), .out(n5699), .config_in(config_chain[8000:7998]), .config_rst(config_rst)); 
mux6 mux_2667 (.in({n13673_0, n13672_0, n13661_0, n13660_0, n13627_0, n13626_1/**/}), .out(n5700), .config_in(config_chain[8003:8001]), .config_rst(config_rst)); 
mux6 mux_2668 (.in({n10885_1, n10884_0, n10877_1, n10876_0, n10807_0, n10806_1}), .out(n5701), .config_in(config_chain[8006:8004]), .config_rst(config_rst)); 
mux6 mux_2669 (.in({n13975_1, n13974_0, n13861_0/**/, n13860_1, n13829_0, n13828_1}), .out(n5702), .config_in(config_chain[8009:8007]), .config_rst(config_rst)); 
mux6 mux_2670 (.in({n10609_1/**/, n10608_0, n10595_0, n10594_0, n10583_0, n10582_0}), .out(n5703), .config_in(config_chain[8012:8010]), .config_rst(config_rst)); 
mux6 mux_2671 (.in({n13695_1, n13694_0, n13689_0/**/, n13688_0, n13681_0, n13680_0}), .out(n5704), .config_in(config_chain[8015:8013]), .config_rst(config_rst)); 
mux6 mux_2672 (.in({n10837_0, n10836_0, n10829_0, n10828_0, n10823_0, n10822_1}), .out(n5705), .config_in(config_chain[8018:8016]), .config_rst(config_rst)); 
mux6 mux_2673 (.in({n13939_0, n13938_0, n13927_0, n13926_0/**/, n13893_0, n13892_1}), .out(n5706), .config_in(config_chain[8021:8019]), .config_rst(config_rst)); 
mux6 mux_2674 (.in({n10617_1, n10616_0, n10603_0, n10602_0/**/, n10549_0, n10548_1}), .out(n5707), .config_in(config_chain[8024:8022]), .config_rst(config_rst)); 
mux6 mux_2675 (.in({n13711_1, n13710_0, n13703_1, n13702_0, n13571_0, n13570_1}), .out(n5708), .config_in(config_chain[8027:8025]), .config_rst(config_rst)); 
mux6 mux_2676 (.in({n10857_0, n10856_0, n10849_0, n10848_0/**/, n10845_0, n10844_0}), .out(n5709), .config_in(config_chain[8030:8028]), .config_rst(config_rst)); 
mux6 mux_2677 (.in({n13961_1, n13960_0, n13947_0/**/, n13946_0, n13935_0, n13934_0}), .out(n5710), .config_in(config_chain[8033:8031]), .config_rst(config_rst)); 
mux6 mux_2678 (.in({n10569_0, n10568_0, n10565_0/**/, n10564_1, n10557_0, n10556_1}), .out(n5711), .config_in(config_chain[8036:8034]), .config_rst(config_rst)); 
mux6 mux_2679 (.in({n13663_0, n13662_0, n13655_0, n13654_0, n13635_0/**/, n13634_1}), .out(n5712), .config_in(config_chain[8039:8037]), .config_rst(config_rst)); 
mux6 mux_2680 (.in({n10879_1/**/, n10878_0, n10865_0, n10864_0, n10809_0, n10808_1}), .out(n5713), .config_in(config_chain[8042:8040]), .config_rst(config_rst)); 
mux6 mux_2681 (.in({n13977_1, n13976_0, n13969_1, n13968_0, n13837_0/**/, n13836_1}), .out(n5714), .config_in(config_chain[8045:8043]), .config_rst(config_rst)); 
mux6 mux_2682 (.in({n10597_0, n10596_0, n10589_0, n10588_0, n10585_0/**/, n10584_0}), .out(n5715), .config_in(config_chain[8048:8046]), .config_rst(config_rst)); 
mux6 mux_2683 (.in({n13683_0, n13682_0, n13675_0/**/, n13674_0, n13671_0, n13670_0}), .out(n5716), .config_in(config_chain[8051:8049]), .config_rst(config_rst)); 
mux6 mux_2684 (.in({n10887_1, n10886_0, n10831_0/**/, n10830_0, n10817_0, n10816_1}), .out(n5717), .config_in(config_chain[8054:8052]), .config_rst(config_rst)); 
mux6 mux_2685 (.in({n13921_0, n13920_0, n13901_0/**/, n13900_1, n13869_0, n13868_1}), .out(n5718), .config_in(config_chain[8057:8055]), .config_rst(config_rst)); 
mux6 mux_2686 (.in({n10619_1/**/, n10618_0, n10611_1, n10610_0, n10605_0, n10604_0}), .out(n5719), .config_in(config_chain[8060:8058]), .config_rst(config_rst)); 
mux6 mux_2687 (.in({n13705_1, n13704_0, n13691_0, n13690_0, n13579_0, n13578_1/**/}), .out(n5720), .config_in(config_chain[8063:8061]), .config_rst(config_rst)); 
mux6 mux_2688 (.in({n10851_0, n10850_0, n10839_0, n10838_0, n10781_0/**/, n10780_1}), .out(n5721), .config_in(config_chain[8066:8064]), .config_rst(config_rst)); 
mux6 mux_2689 (.in({n13949_0, n13948_0, n13941_0, n13940_0, n13911_0, n13910_1}), .out(n5722), .config_in(config_chain[8069:8067]), .config_rst(config_rst)); 
mux6 mux_2690 (.in({n10571_0, n10570_0, n10559_0, n10558_1, n10523_1, n10522_1}), .out(n5723), .config_in(config_chain[8072:8070]), .config_rst(config_rst)); 
mux6 mux_2691 (.in({n13657_0, n13656_0/**/, n13649_1, n13648_1, n13611_0, n13610_1}), .out(n5724), .config_in(config_chain[8075:8073]), .config_rst(config_rst)); 
mux6 mux_2692 (.in({n10873_1, n10872_0, n10859_0, n10858_0, n10783_0, n10782_1/**/}), .out(n5725), .config_in(config_chain[8078:8076]), .config_rst(config_rst)); 
mux6 mux_2693 (.in({n13971_1, n13970_0, n13963_1/**/, n13962_0, n13913_0, n13912_1}), .out(n5726), .config_in(config_chain[8081:8079]), .config_rst(config_rst)); 
mux6 mux_2694 (.in({n10591_0, n10590_0, n10579_0, n10578_0, n10525_1/**/, n10524_1}), .out(n5727), .config_in(config_chain[8084:8082]), .config_rst(config_rst)); 
mux6 mux_2695 (.in({n13713_1, n13712_0, n13677_0, n13676_0/**/, n13665_0, n13664_0}), .out(n5728), .config_in(config_chain[8087:8085]), .config_rst(config_rst)); 
mux6 mux_2696 (.in({n10819_0/**/, n10818_1, n10811_0, n10810_1, n10785_1, n10784_1}), .out(n5729), .config_in(config_chain[8090:8088]), .config_rst(config_rst)); 
mux6 mux_2697 (.in({n13923_0, n13922_0/**/, n13915_1, n13914_1, n13877_0, n13876_1}), .out(n5730), .config_in(config_chain[8093:8091]), .config_rst(config_rst)); 
mux6 mux_2698 (.in({n10613_1, n10612_0, n10599_0/**/, n10598_0, n10517_0, n10516_1}), .out(n5731), .config_in(config_chain[8096:8094]), .config_rst(config_rst)); 
mux6 mux_2699 (.in({n13707_1, n13706_0, n13699_1, n13698_0, n13643_0, n13642_1}), .out(n5732), .config_in(config_chain[8099:8097]), .config_rst(config_rst)); 
mux6 mux_2700 (.in({n10867_1, n10866_0, n10841_0, n10840_0, n10833_0, n10832_0}), .out(n5733), .config_in(config_chain[8102:8100]), .config_rst(config_rst)); 
mux6 mux_2701 (.in({n13957_1, n13956_0, n13943_0, n13942_0, n13931_0, n13930_0/**/}), .out(n5734), .config_in(config_chain[8105:8103]), .config_rst(config_rst)); 
mux6 mux_2702 (.in({n10621_1, n10620_0, n10553_0, n10552_1/**/, n10519_0, n10518_1}), .out(n5735), .config_in(config_chain[8108:8106]), .config_rst(config_rst)); 
mux6 mux_2703 (.in({n13645_0, n13644_1, n13619_0, n13618_1, n13587_0/**/, n13586_1}), .out(n5736), .config_in(config_chain[8111:8109]), .config_rst(config_rst)); 
mux6 mux_2704 (.in({n10889_1, n10888_0/**/, n10875_1, n10874_0, n10861_0, n10860_0}), .out(n5737), .config_in(config_chain[8114:8112]), .config_rst(config_rst)); 
mux6 mux_2705 (.in({n13965_1, n13964_0, n13951_0/**/, n13950_0, n13909_0, n13908_1}), .out(n5738), .config_in(config_chain[8117:8115]), .config_rst(config_rst)); 
mux6 mux_2706 (.in({n10581_0/**/, n10580_0, n10573_0, n10572_0, n10521_0, n10520_1}), .out(n5739), .config_in(config_chain[8120:8118]), .config_rst(config_rst)); 
mux6 mux_2707 (.in({n13679_0, n13678_0, n13667_0, n13666_0, n13647_0, n13646_1}), .out(n5740), .config_in(config_chain[8123:8121]), .config_rst(config_rst)); 
mux6 mux_2708 (.in({n11133_1, n11132_0, n11117_0, n11116_0, n11103_0, n11102_0}), .out(n5787), .config_in(config_chain[8126:8124]), .config_rst(config_rst)); 
mux6 mux_2709 (.in({n13981_1, n13980_0, n13965_0, n13964_0/**/, n13951_0, n13950_0}), .out(n5788), .config_in(config_chain[8129:8127]), .config_rst(config_rst)); 
mux6 mux_2710 (.in({n10827_0, n10826_0, n10821_0, n10820_1, n10813_0, n10812_1}), .out(n5789), .config_in(config_chain[8132:8130]), .config_rst(config_rst)); 
mux6 mux_2711 (.in({n13681_0, n13680_0, n13673_0, n13672_0, n13667_0, n13666_1}), .out(n5790), .config_in(config_chain[8135:8133]), .config_rst(config_rst)); 
mux6 mux_2712 (.in({n11141_1, n11140_0, n11125_0/**/, n11124_0, n11069_0, n11068_1}), .out(n5791), .config_in(config_chain[8138:8136]), .config_rst(config_rst)); 
mux6 mux_2713 (.in({n13997_1, n13996_0, n13989_1, n13988_0, n13917_0, n13916_1}), .out(n5792), .config_in(config_chain[8141:8139]), .config_rst(config_rst)); 
mux6 mux_2714 (.in({n10855_0, n10854_0, n10847_0, n10846_0, n10843_0, n10842_0}), .out(n5793), .config_in(config_chain[8144:8142]), .config_rst(config_rst)); 
mux6 mux_2715 (.in({n13715_1/**/, n13714_0, n13701_0, n13700_0, n13689_0, n13688_0}), .out(n5794), .config_in(config_chain[8147:8145]), .config_rst(config_rst)); 
mux6 mux_2716 (.in({n11089_0, n11088_0, n11085_0, n11084_1, n11077_0, n11076_1}), .out(n5795), .config_in(config_chain[8150:8148]), .config_rst(config_rst)); 
mux6 mux_2717 (.in({n13937_0, n13936_0, n13933_0/**/, n13932_1, n13925_0, n13924_1}), .out(n5796), .config_in(config_chain[8153:8151]), .config_rst(config_rst)); 
mux6 mux_2718 (.in({n10877_1, n10876_0, n10869_1, n10868_0, n10863_0, n10862_0}), .out(n5797), .config_in(config_chain[8156:8154]), .config_rst(config_rst)); 
mux6 mux_2719 (.in({n13723_1, n13722_0, n13709_0/**/, n13708_0, n13653_0, n13652_1}), .out(n5798), .config_in(config_chain[8159:8157]), .config_rst(config_rst)); 
mux6 mux_2720 (.in({n11111_0, n11110_0, n11105_0, n11104_0, n11097_0, n11096_0}), .out(n5799), .config_in(config_chain[8162:8160]), .config_rst(config_rst)); 
mux6 mux_2721 (.in({n13967_0, n13966_0, n13959_0, n13958_0/**/, n13953_0, n13952_0}), .out(n5800), .config_in(config_chain[8165:8163]), .config_rst(config_rst)); 
mux6 mux_2722 (.in({n10885_1, n10884_0, n10829_0, n10828_0, n10815_0/**/, n10814_1}), .out(n5801), .config_in(config_chain[8168:8166]), .config_rst(config_rst)); 
mux6 mux_2723 (.in({n13675_0, n13674_0/**/, n13669_0, n13668_1, n13661_0, n13660_1}), .out(n5802), .config_in(config_chain[8171:8169]), .config_rst(config_rst)); 
mux6 mux_2724 (.in({n11143_1, n11142_0, n11135_1, n11134_0, n11127_0, n11126_0}), .out(n5803), .config_in(config_chain[8174:8172]), .config_rst(config_rst)); 
mux6 mux_2725 (.in({n13991_1, n13990_0, n13975_0, n13974_0, n13919_0, n13918_1/**/}), .out(n5804), .config_in(config_chain[8177:8175]), .config_rst(config_rst)); 
mux6 mux_2726 (.in({n10849_0, n10848_0, n10837_0, n10836_0, n10823_0, n10822_1/**/}), .out(n5805), .config_in(config_chain[8180:8178]), .config_rst(config_rst)); 
mux6 mux_2727 (.in({n13695_0, n13694_0, n13691_0, n13690_0, n13683_0, n13682_0}), .out(n5806), .config_in(config_chain[8183:8181]), .config_rst(config_rst)); 
mux6 mux_2728 (.in({n11151_1, n11150_0, n11079_0, n11078_1/**/, n11071_0, n11070_1}), .out(n5807), .config_in(config_chain[8186:8184]), .config_rst(config_rst)); 
mux6 mux_2729 (.in({n13999_1, n13998_0, n13939_0, n13938_0, n13927_0/**/, n13926_1}), .out(n5808), .config_in(config_chain[8189:8187]), .config_rst(config_rst)); 
mux6 mux_2730 (.in({n10871_1/**/, n10870_0, n10865_0, n10864_0, n10857_0, n10856_0}), .out(n5809), .config_in(config_chain[8192:8190]), .config_rst(config_rst)); 
mux6 mux_2731 (.in({n13725_1, n13724_0, n13717_1, n13716_0, n13711_0, n13710_0}), .out(n5810), .config_in(config_chain[8195:8193]), .config_rst(config_rst)); 
mux6 mux_2732 (.in({n11113_0, n11112_0, n11099_0, n11098_0, n11087_0/**/, n11086_1}), .out(n5811), .config_in(config_chain[8198:8196]), .config_rst(config_rst)); 
mux6 mux_2733 (.in({n13961_0, n13960_0, n13955_0, n13954_0, n13947_0, n13946_0}), .out(n5812), .config_in(config_chain[8201:8199]), .config_rst(config_rst)); 
mux6 mux_2734 (.in({n10887_1, n10886_0, n10817_0, n10816_1, n10809_0, n10808_1}), .out(n5813), .config_in(config_chain[8204:8202]), .config_rst(config_rst)); 
mux6 mux_2735 (.in({n13733_1, n13732_0, n13663_0, n13662_1, n13655_0, n13654_1}), .out(n5814), .config_in(config_chain[8207:8205]), .config_rst(config_rst)); 
mux6 mux_2736 (.in({n11137_1/**/, n11136_0, n11121_0, n11120_0, n11107_0, n11106_0}), .out(n5815), .config_in(config_chain[8210:8208]), .config_rst(config_rst)); 
mux6 mux_2737 (.in({n13985_1, n13984_0, n13977_0, n13976_0, n13969_0/**/, n13968_0}), .out(n5816), .config_in(config_chain[8213:8211]), .config_rst(config_rst)); 
mux6 mux_2738 (.in({n10839_0, n10838_0/**/, n10831_0, n10830_0, n10825_0, n10824_1}), .out(n5817), .config_in(config_chain[8216:8214]), .config_rst(config_rst)); 
mux6 mux_2739 (.in({n13697_0, n13696_0, n13685_0, n13684_0, n13671_0/**/, n13670_1}), .out(n5818), .config_in(config_chain[8219:8217]), .config_rst(config_rst)); 
mux6 mux_2740 (.in({n11153_1, n11152_0, n11145_1, n11144_0, n11073_0, n11072_1}), .out(n5819), .config_in(config_chain[8222:8220]), .config_rst(config_rst)); 
mux6 mux_2741 (.in({n14001_1, n14000_0, n13929_0, n13928_1, n13921_0/**/, n13920_1}), .out(n5820), .config_in(config_chain[8225:8223]), .config_rst(config_rst)); 
mux6 mux_2742 (.in({n10873_1, n10872_0, n10859_0/**/, n10858_0, n10781_0, n10780_1}), .out(n5821), .config_in(config_chain[8228:8226]), .config_rst(config_rst)); 
mux6 mux_2743 (.in({n13719_1, n13718_0, n13705_0, n13704_0/**/, n13647_0, n13646_1}), .out(n5822), .config_in(config_chain[8231:8229]), .config_rst(config_rst)); 
mux6 mux_2744 (.in({n11093_0, n11092_0, n11081_0, n11080_1/**/, n11043_0, n11042_1}), .out(n5823), .config_in(config_chain[8234:8232]), .config_rst(config_rst)); 
mux6 mux_2745 (.in({n13949_0, n13948_0/**/, n13941_0, n13940_0, n13911_0, n13910_1}), .out(n5824), .config_in(config_chain[8237:8235]), .config_rst(config_rst)); 
mux6 mux_2746 (.in({n10881_1, n10880_0, n10811_0, n10810_1/**/, n10783_0, n10782_1}), .out(n5825), .config_in(config_chain[8240:8238]), .config_rst(config_rst)); 
mux6 mux_2747 (.in({n13727_1, n13726_0, n13657_0/**/, n13656_1, n13651_1, n13650_1}), .out(n5826), .config_in(config_chain[8243:8241]), .config_rst(config_rst)); 
mux6 mux_2748 (.in({n11123_0, n11122_0, n11115_0, n11114_0, n11045_0, n11044_1}), .out(n5827), .config_in(config_chain[8246:8244]), .config_rst(config_rst)); 
mux6 mux_2749 (.in({n13987_1/**/, n13986_0, n13971_0, n13970_0, n13913_0, n13912_1}), .out(n5828), .config_in(config_chain[8249:8247]), .config_rst(config_rst)); 
mux6 mux_2750 (.in({n10867_1, n10866_0, n10833_0, n10832_0, n10819_0, n10818_1}), .out(n5829), .config_in(config_chain[8252:8250]), .config_rst(config_rst)); 
mux6 mux_2751 (.in({n13713_1, n13712_0, n13687_0, n13686_0, n13679_0, n13678_0}), .out(n5830), .config_in(config_chain[8255:8253]), .config_rst(config_rst)); 
mux6 mux_2752 (.in({n11147_1, n11146_0, n11139_1, n11138_0, n11047_0, n11046_1}), .out(n5831), .config_in(config_chain[8258:8256]), .config_rst(config_rst)); 
mux6 mux_2753 (.in({n13995_1/**/, n13994_0, n13923_0, n13922_1, n13915_0, n13914_1}), .out(n5832), .config_in(config_chain[8261:8259]), .config_rst(config_rst)); 
mux6 mux_2754 (.in({n10889_1, n10888_0, n10853_0, n10852_0, n10841_0/**/, n10840_0}), .out(n5833), .config_in(config_chain[8264:8262]), .config_rst(config_rst)); 
mux6 mux_2755 (.in({n13735_1, n13734_0, n13707_0, n13706_0/**/, n13699_0, n13698_0}), .out(n5834), .config_in(config_chain[8267:8265]), .config_rst(config_rst)); 
mux6 mux_2756 (.in({n11109_1, n11108_0, n11095_0, n11094_0, n11083_0, n11082_1/**/}), .out(n5835), .config_in(config_chain[8270:8268]), .config_rst(config_rst)); 
mux6 mux_2757 (.in({n13979_1, n13978_0, n13943_0, n13942_0, n13931_0, n13930_1}), .out(n5836), .config_in(config_chain[8273:8271]), .config_rst(config_rst)); 
mux6 mux_2758 (.in({n10883_1, n10882_0, n10875_1, n10874_0/**/, n10779_0, n10778_1}), .out(n5837), .config_in(config_chain[8276:8274]), .config_rst(config_rst)); 
mux6 mux_2759 (.in({n13729_1/**/, n13728_0, n13659_0, n13658_1, n13645_0, n13644_1}), .out(n5838), .config_in(config_chain[8279:8277]), .config_rst(config_rst)); 
mux6 mux_2760 (.in({n11413_1, n11412_0, n11355_0/**/, n11354_0, n11339_0, n11338_1}), .out(n5885), .config_in(config_chain[8282:8280]), .config_rst(config_rst)); 
mux6 mux_2761 (.in({n14017_1, n14016_0, n13959_0, n13958_0, n13943_0, n13942_1}), .out(n5886), .config_in(config_chain[8285:8283]), .config_rst(config_rst)); 
mux6 mux_2762 (.in({n11133_1, n11132_0, n11125_0, n11124_0, n11117_0, n11116_0}), .out(n5887), .config_in(config_chain[8288:8286]), .config_rst(config_rst)); 
mux6 mux_2763 (.in({n13745_1, n13744_0, n13737_1, n13736_0, n13729_0/**/, n13728_0}), .out(n5888), .config_in(config_chain[8291:8289]), .config_rst(config_rst)); 
mux6 mux_2764 (.in({n11377_0, n11376_0, n11363_0, n11362_0, n11347_0, n11346_1}), .out(n5889), .config_in(config_chain[8294:8292]), .config_rst(config_rst)); 
mux6 mux_2765 (.in({n13981_0, n13980_0, n13975_0/**/, n13974_0, n13967_0, n13966_0}), .out(n5890), .config_in(config_chain[8297:8295]), .config_rst(config_rst)); 
mux6 mux_2766 (.in({n11149_1, n11148_0, n11077_0, n11076_1, n11069_0, n11068_1}), .out(n5891), .config_in(config_chain[8300:8298]), .config_rst(config_rst)); 
mux6 mux_2767 (.in({n13753_1, n13752_0, n13693_0, n13692_0, n13681_0, n13680_1}), .out(n5892), .config_in(config_chain[8303:8301]), .config_rst(config_rst)); 
mux6 mux_2768 (.in({n11399_1, n11398_0, n11393_0, n11392_0, n11385_0, n11384_0}), .out(n5893), .config_in(config_chain[8306:8304]), .config_rst(config_rst)); 
mux6 mux_2769 (.in({n14003_1, n14002_0, n13997_0, n13996_0/**/, n13989_0, n13988_0}), .out(n5894), .config_in(config_chain[8309:8307]), .config_rst(config_rst)); 
mux6 mux_2770 (.in({n11097_0, n11096_0, n11089_0, n11088_0, n11085_0, n11084_1}), .out(n5895), .config_in(config_chain[8312:8310]), .config_rst(config_rst)); 
mux6 mux_2771 (.in({n13715_0, n13714_0, n13701_0, n13700_0, n13689_0, n13688_1}), .out(n5896), .config_in(config_chain[8315:8313]), .config_rst(config_rst)); 
mux6 mux_2772 (.in({n11415_1, n11414_0, n11407_1/**/, n11406_0, n11333_0, n11332_1}), .out(n5897), .config_in(config_chain[8318:8316]), .config_rst(config_rst)); 
mux6 mux_2773 (.in({n14019_1, n14018_0, n13945_0, n13944_1, n13937_0, n13936_1}), .out(n5898), .config_in(config_chain[8321:8319]), .config_rst(config_rst)); 
mux6 mux_2774 (.in({n11135_1, n11134_0, n11119_0/**/, n11118_0, n11105_0, n11104_0}), .out(n5899), .config_in(config_chain[8324:8322]), .config_rst(config_rst)); 
mux6 mux_2775 (.in({n13739_1, n13738_0/**/, n13731_0, n13730_0, n13723_0, n13722_0}), .out(n5900), .config_in(config_chain[8327:8325]), .config_rst(config_rst)); 
mux6 mux_2776 (.in({n11365_0, n11364_0, n11357_0, n11356_0, n11349_0, n11348_1/**/}), .out(n5901), .config_in(config_chain[8330:8328]), .config_rst(config_rst)); 
mux6 mux_2777 (.in({n13983_0, n13982_0, n13969_0, n13968_0, n13953_0, n13952_1}), .out(n5902), .config_in(config_chain[8333:8331]), .config_rst(config_rst)); 
mux6 mux_2778 (.in({n11143_1, n11142_0, n11127_0, n11126_0/**/, n11071_0, n11070_1}), .out(n5903), .config_in(config_chain[8336:8334]), .config_rst(config_rst)); 
mux6 mux_2779 (.in({n13755_1, n13754_0, n13747_1, n13746_0, n13675_0, n13674_1}), .out(n5904), .config_in(config_chain[8339:8337]), .config_rst(config_rst)); 
mux6 mux_2780 (.in({n11387_0, n11386_0, n11379_0/**/, n11378_0, n11373_0, n11372_0}), .out(n5905), .config_in(config_chain[8342:8340]), .config_rst(config_rst)); 
mux6 mux_2781 (.in({n14005_1, n14004_0, n13991_0/**/, n13990_0, n13977_0, n13976_0}), .out(n5906), .config_in(config_chain[8345:8343]), .config_rst(config_rst)); 
mux6 mux_2782 (.in({n11091_0, n11090_0, n11087_0, n11086_1/**/, n11079_0, n11078_1}), .out(n5907), .config_in(config_chain[8348:8346]), .config_rst(config_rst)); 
mux6 mux_2783 (.in({n13703_0, n13702_0/**/, n13695_0, n13694_0, n13691_0, n13690_1}), .out(n5908), .config_in(config_chain[8351:8349]), .config_rst(config_rst)); 
mux6 mux_2784 (.in({n11409_1, n11408_0, n11395_0, n11394_0/**/, n11335_0, n11334_1}), .out(n5909), .config_in(config_chain[8354:8352]), .config_rst(config_rst)); 
mux6 mux_2785 (.in({n14021_1, n14020_0, n14013_1, n14012_0, n13939_0, n13938_1}), .out(n5910), .config_in(config_chain[8357:8355]), .config_rst(config_rst)); 
mux6 mux_2786 (.in({n11121_0, n11120_0, n11113_0/**/, n11112_0, n11107_0, n11106_0}), .out(n5911), .config_in(config_chain[8360:8358]), .config_rst(config_rst)); 
mux6 mux_2787 (.in({n13725_0, n13724_0, n13717_0, n13716_0, n13711_0, n13710_0/**/}), .out(n5912), .config_in(config_chain[8363:8361]), .config_rst(config_rst)); 
mux6 mux_2788 (.in({n11417_1, n11416_0, n11359_0/**/, n11358_0, n11343_0, n11342_1}), .out(n5913), .config_in(config_chain[8366:8364]), .config_rst(config_rst)); 
mux6 mux_2789 (.in({n13963_0, n13962_0, n13955_0, n13954_1, n13947_0, n13946_1}), .out(n5914), .config_in(config_chain[8369:8367]), .config_rst(config_rst)); 
mux6 mux_2790 (.in({n11145_1, n11144_0, n11137_1, n11136_0, n11129_0, n11128_0/**/}), .out(n5915), .config_in(config_chain[8372:8370]), .config_rst(config_rst)); 
mux6 mux_2791 (.in({n13749_1, n13748_0/**/, n13733_0, n13732_0, n13677_0, n13676_1}), .out(n5916), .config_in(config_chain[8375:8373]), .config_rst(config_rst)); 
mux6 mux_2792 (.in({n11381_0, n11380_0/**/, n11375_1, n11374_0, n11367_0, n11366_0}), .out(n5917), .config_in(config_chain[8378:8376]), .config_rst(config_rst)); 
mux6 mux_2793 (.in({n13993_0/**/, n13992_0, n13985_0, n13984_0, n13979_1, n13978_0}), .out(n5918), .config_in(config_chain[8381:8379]), .config_rst(config_rst)); 
mux6 mux_2794 (.in({n11153_1, n11152_0, n11093_0, n11092_0, n11081_0, n11080_1}), .out(n5919), .config_in(config_chain[8384:8382]), .config_rst(config_rst)); 
mux6 mux_2795 (.in({n13757_1, n13756_0/**/, n13697_0, n13696_0, n13685_0, n13684_1}), .out(n5920), .config_in(config_chain[8387:8385]), .config_rst(config_rst)); 
mux6 mux_2796 (.in({n11403_1, n11402_0, n11397_1, n11396_0, n11389_0, n11388_0}), .out(n5921), .config_in(config_chain[8390:8388]), .config_rst(config_rst)); 
mux6 mux_2797 (.in({n14015_1, n14014_0, n14007_1, n14006_0/**/, n14001_1, n14000_0}), .out(n5922), .config_in(config_chain[8393:8391]), .config_rst(config_rst)); 
mux6 mux_2798 (.in({n11115_0, n11114_0, n11101_0/**/, n11100_0, n11043_0, n11042_1}), .out(n5923), .config_in(config_chain[8396:8394]), .config_rst(config_rst)); 
mux6 mux_2799 (.in({n13719_0, n13718_0/**/, n13705_0, n13704_0, n13649_0, n13648_1}), .out(n5924), .config_in(config_chain[8399:8397]), .config_rst(config_rst)); 
mux6 mux_2800 (.in({n11419_1, n11418_0, n11345_0, n11344_1, n11337_0, n11336_1}), .out(n5925), .config_in(config_chain[8402:8400]), .config_rst(config_rst)); 
mux6 mux_2801 (.in({n14023_1, n14022_0, n13965_0, n13964_0, n13949_0, n13948_1}), .out(n5926), .config_in(config_chain[8405:8403]), .config_rst(config_rst)); 
mux6 mux_2802 (.in({n11139_1, n11138_0, n11123_0, n11122_0, n11047_0/**/, n11046_1}), .out(n5927), .config_in(config_chain[8408:8406]), .config_rst(config_rst)); 
mux6 mux_2803 (.in({n13751_1, n13750_0, n13743_1, n13742_0, n13651_0/**/, n13650_1}), .out(n5928), .config_in(config_chain[8411:8409]), .config_rst(config_rst)); 
mux6 mux_2804 (.in({n11369_0, n11368_0, n11361_0/**/, n11360_0, n11309_0, n11308_1}), .out(n5929), .config_in(config_chain[8414:8412]), .config_rst(config_rst)); 
mux6 mux_2805 (.in({n13987_0, n13986_0, n13973_0, n13972_0, n13913_0, n13912_1}), .out(n5930), .config_in(config_chain[8417:8415]), .config_rst(config_rst)); 
mux6 mux_2806 (.in({n11147_1, n11146_0/**/, n11109_1, n11108_0, n11075_0, n11074_1}), .out(n5931), .config_in(config_chain[8420:8418]), .config_rst(config_rst)); 
mux6 mux_2807 (.in({n13713_1, n13712_0, n13687_0, n13686_1, n13679_0, n13678_1}), .out(n5932), .config_in(config_chain[8423:8421]), .config_rst(config_rst)); 
mux6 mux_2808 (.in({n11405_1, n11404_0, n11391_0/**/, n11390_0, n11311_0, n11310_1}), .out(n5933), .config_in(config_chain[8426:8424]), .config_rst(config_rst)); 
mux6 mux_2809 (.in({n14009_1, n14008_0, n13995_0/**/, n13994_0, n13957_1, n13956_1}), .out(n5934), .config_in(config_chain[8429:8427]), .config_rst(config_rst)); 
mux6 mux_2810 (.in({n11131_1, n11130_0, n11103_0, n11102_0, n11095_0, n11094_0/**/}), .out(n5935), .config_in(config_chain[8432:8430]), .config_rst(config_rst)); 
mux6 mux_2811 (.in({n13735_1, n13734_0, n13721_0, n13720_0, n13707_0, n13706_0}), .out(n5936), .config_in(config_chain[8435:8433]), .config_rst(config_rst)); 
mux6 mux_2812 (.in({n11665_1, n11664_0, n11649_0, n11648_0, n11635_0, n11634_0}), .out(n5983), .config_in(config_chain[8438:8436]), .config_rst(config_rst)); 
mux6 mux_2813 (.in({n14025_0, n14024_0, n14009_0, n14008_0, n13995_0, n13994_0}), .out(n5984), .config_in(config_chain[8441:8439]), .config_rst(config_rst)); 
mux6 mux_2814 (.in({n11355_0, n11354_0, n11347_0, n11346_1, n11339_0, n11338_1}), .out(n5985), .config_in(config_chain[8444:8442]), .config_rst(config_rst)); 
mux6 mux_2815 (.in({n13723_0, n13722_0, n13715_0, n13714_0, n13707_0, n13706_1}), .out(n5986), .config_in(config_chain[8447:8445]), .config_rst(config_rst)); 
mux6 mux_2816 (.in({n11673_1, n11672_0, n11657_0, n11656_0, n11599_0, n11598_1}), .out(n5987), .config_in(config_chain[8450:8448]), .config_rst(config_rst)); 
mux6 mux_2817 (.in({n14041_0, n14040_0, n14033_0, n14032_0, n13959_0, n13958_1}), .out(n5988), .config_in(config_chain[8453:8451]), .config_rst(config_rst)); 
mux6 mux_2818 (.in({n11385_0, n11384_0, n11377_0, n11376_0, n11371_0, n11370_0}), .out(n5989), .config_in(config_chain[8456:8454]), .config_rst(config_rst)); 
mux6 mux_2819 (.in({n13759_0, n13758_0, n13745_0, n13744_0, n13731_0, n13730_0}), .out(n5990), .config_in(config_chain[8459:8457]), .config_rst(config_rst)); 
mux6 mux_2820 (.in({n11621_0, n11620_0, n11615_0, n11614_1, n11607_0, n11606_1}), .out(n5991), .config_in(config_chain[8462:8460]), .config_rst(config_rst)); 
mux6 mux_2821 (.in({n13981_0, n13980_0, n13975_0, n13974_1, n13967_0, n13966_1}), .out(n5992), .config_in(config_chain[8465:8463]), .config_rst(config_rst)); 
mux6 mux_2822 (.in({n11407_1, n11406_0, n11399_1, n11398_0, n11393_0, n11392_0}), .out(n5993), .config_in(config_chain[8468:8466]), .config_rst(config_rst)); 
mux6 mux_2823 (.in({n13767_0, n13766_0/**/, n13753_0, n13752_0, n13693_0, n13692_1}), .out(n5994), .config_in(config_chain[8471:8469]), .config_rst(config_rst)); 
mux6 mux_2824 (.in({n11643_0, n11642_0, n11637_0, n11636_0/**/, n11629_0, n11628_0}), .out(n5995), .config_in(config_chain[8474:8472]), .config_rst(config_rst)); 
mux6 mux_2825 (.in({n14011_0, n14010_0/**/, n14003_0, n14002_0, n13997_0, n13996_0}), .out(n5996), .config_in(config_chain[8477:8475]), .config_rst(config_rst)); 
mux6 mux_2826 (.in({n11415_1, n11414_0, n11357_0, n11356_0/**/, n11341_0, n11340_1}), .out(n5997), .config_in(config_chain[8480:8478]), .config_rst(config_rst)); 
mux6 mux_2827 (.in({n13717_0, n13716_0, n13709_0, n13708_1, n13701_0, n13700_1/**/}), .out(n5998), .config_in(config_chain[8483:8481]), .config_rst(config_rst)); 
mux6 mux_2828 (.in({n11675_1, n11674_0, n11667_1, n11666_0, n11659_0, n11658_0}), .out(n5999), .config_in(config_chain[8486:8484]), .config_rst(config_rst)); 
mux6 mux_2829 (.in({n14035_0, n14034_0/**/, n14019_0, n14018_0, n13961_0, n13960_1}), .out(n6000), .config_in(config_chain[8489:8487]), .config_rst(config_rst)); 
mux6 mux_2830 (.in({n11379_0, n11378_0, n11365_0, n11364_0, n11349_0, n11348_1/**/}), .out(n6001), .config_in(config_chain[8492:8490]), .config_rst(config_rst)); 
mux6 mux_2831 (.in({n13739_0, n13738_0, n13733_0, n13732_0/**/, n13725_0, n13724_0}), .out(n6002), .config_in(config_chain[8495:8493]), .config_rst(config_rst)); 
mux6 mux_2832 (.in({n11683_1, n11682_0/**/, n11609_0, n11608_1, n11601_0, n11600_1}), .out(n6003), .config_in(config_chain[8498:8496]), .config_rst(config_rst)); 
mux6 mux_2833 (.in({n14043_0, n14042_0, n13983_0, n13982_0, n13969_0, n13968_1}), .out(n6004), .config_in(config_chain[8501:8499]), .config_rst(config_rst)); 
mux6 mux_2834 (.in({n11401_1, n11400_0, n11395_0, n11394_0, n11387_0, n11386_0}), .out(n6005), .config_in(config_chain[8504:8502]), .config_rst(config_rst)); 
mux6 mux_2835 (.in({n13769_0, n13768_0, n13761_0, n13760_0/**/, n13755_0, n13754_0}), .out(n6006), .config_in(config_chain[8507:8505]), .config_rst(config_rst)); 
mux6 mux_2836 (.in({n11645_0, n11644_0, n11631_0, n11630_0, n11617_0/**/, n11616_1}), .out(n6007), .config_in(config_chain[8510:8508]), .config_rst(config_rst)); 
mux6 mux_2837 (.in({n14005_0, n14004_0, n13999_0, n13998_0, n13991_0, n13990_0}), .out(n6008), .config_in(config_chain[8513:8511]), .config_rst(config_rst)); 
mux6 mux_2838 (.in({n11417_1, n11416_0, n11343_0/**/, n11342_1, n11335_0, n11334_1}), .out(n6009), .config_in(config_chain[8516:8514]), .config_rst(config_rst)); 
mux6 mux_2839 (.in({n13777_0, n13776_0/**/, n13703_0, n13702_1, n13695_0, n13694_1}), .out(n6010), .config_in(config_chain[8519:8517]), .config_rst(config_rst)); 
mux6 mux_2840 (.in({n11669_1, n11668_0, n11653_0, n11652_0/**/, n11639_0, n11638_0}), .out(n6011), .config_in(config_chain[8522:8520]), .config_rst(config_rst)); 
mux6 mux_2841 (.in({n14029_0, n14028_0, n14021_0, n14020_0, n14013_0, n14012_0}), .out(n6012), .config_in(config_chain[8525:8523]), .config_rst(config_rst)); 
mux6 mux_2842 (.in({n11367_0, n11366_0, n11359_0, n11358_0/**/, n11351_0, n11350_1}), .out(n6013), .config_in(config_chain[8528:8526]), .config_rst(config_rst)); 
mux6 mux_2843 (.in({n13741_0, n13740_0/**/, n13727_0, n13726_0, n13711_0, n13710_1}), .out(n6014), .config_in(config_chain[8531:8529]), .config_rst(config_rst)); 
mux6 mux_2844 (.in({n11677_1, n11676_0, n11603_0, n11602_1, n11597_1, n11596_1}), .out(n6015), .config_in(config_chain[8534:8532]), .config_rst(config_rst)); 
mux6 mux_2845 (.in({n13971_0, n13970_1, n13963_0, n13962_1/**/, n13957_0, n13956_1}), .out(n6016), .config_in(config_chain[8537:8535]), .config_rst(config_rst)); 
mux6 mux_2846 (.in({n11403_1, n11402_0, n11389_0, n11388_0, n11375_1, n11374_0}), .out(n6017), .config_in(config_chain[8540:8538]), .config_rst(config_rst)); 
mux6 mux_2847 (.in({n13763_0/**/, n13762_0, n13749_0, n13748_0, n13735_0, n13734_0}), .out(n6018), .config_in(config_chain[8543:8541]), .config_rst(config_rst)); 
mux6 mux_2848 (.in({n11625_0/**/, n11624_0, n11619_1, n11618_1, n11611_0, n11610_1}), .out(n6019), .config_in(config_chain[8546:8544]), .config_rst(config_rst)); 
mux6 mux_2849 (.in({n13993_0, n13992_0, n13985_0, n13984_0, n13979_0, n13978_1}), .out(n6020), .config_in(config_chain[8549:8547]), .config_rst(config_rst)); 
mux6 mux_2850 (.in({n11411_1, n11410_0, n11397_1, n11396_0, n11337_0, n11336_1}), .out(n6021), .config_in(config_chain[8552:8550]), .config_rst(config_rst)); 
mux6 mux_2851 (.in({n13779_0, n13778_0, n13771_0, n13770_0/**/, n13697_0, n13696_1}), .out(n6022), .config_in(config_chain[8555:8553]), .config_rst(config_rst)); 
mux6 mux_2852 (.in({n11655_0, n11654_0, n11647_0, n11646_0, n11641_1, n11640_0}), .out(n6023), .config_in(config_chain[8558:8556]), .config_rst(config_rst)); 
mux6 mux_2853 (.in({n14031_0, n14030_0, n14015_0, n14014_0, n14001_0, n14000_0/**/}), .out(n6024), .config_in(config_chain[8561:8559]), .config_rst(config_rst)); 
mux6 mux_2854 (.in({n11361_0, n11360_0/**/, n11345_0, n11344_1, n11309_0, n11308_1}), .out(n6025), .config_in(config_chain[8564:8562]), .config_rst(config_rst)); 
mux6 mux_2855 (.in({n13729_0, n13728_0, n13721_0, n13720_0, n13649_0, n13648_2}), .out(n6026), .config_in(config_chain[8567:8565]), .config_rst(config_rst)); 
mux6 mux_2856 (.in({n11679_1, n11678_0, n11671_1, n11670_0, n11663_1, n11662_0}), .out(n6027), .config_in(config_chain[8570:8568]), .config_rst(config_rst)); 
mux6 mux_2857 (.in({n14039_0, n14038_0/**/, n14023_0, n14022_0, n13965_0, n13964_1}), .out(n6028), .config_in(config_chain[8573:8571]), .config_rst(config_rst)); 
mux6 mux_2858 (.in({n11383_0, n11382_0, n11369_0/**/, n11368_0, n11311_0, n11310_1}), .out(n6029), .config_in(config_chain[8576:8574]), .config_rst(config_rst)); 
mux6 mux_2859 (.in({n13751_0, n13750_0, n13743_0, n13742_0, n13651_0, n13650_2}), .out(n6030), .config_in(config_chain[8579:8577]), .config_rst(config_rst)); 
mux6 mux_2860 (.in({n11685_1, n11684_0, n11627_0, n11626_0, n11613_0, n11612_1}), .out(n6031), .config_in(config_chain[8582:8580]), .config_rst(config_rst)); 
mux6 mux_2861 (.in({n13987_0, n13986_0, n13973_0, n13972_1, n13915_0, n13914_2}), .out(n6032), .config_in(config_chain[8585:8583]), .config_rst(config_rst)); 
mux6 mux_2862 (.in({n11413_1, n11412_0, n11405_1, n11404_0, n11353_1, n11352_1}), .out(n6033), .config_in(config_chain[8588:8586]), .config_rst(config_rst)); 
mux6 mux_2863 (.in({n13773_0/**/, n13772_0, n13713_0, n13712_1, n13699_0, n13698_1}), .out(n6034), .config_in(config_chain[8591:8589]), .config_rst(config_rst)); 
mux6 mux_2864 (.in({n11943_1, n11942_0, n11885_0, n11884_0, n11869_0, n11868_1}), .out(n6081), .config_in(config_chain[8594:8592]), .config_rst(config_rst)); 
mux6 mux_2865 (.in({n14061_0, n14060_0, n14003_0, n14002_0, n13987_0, n13986_1}), .out(n6082), .config_in(config_chain[8597:8595]), .config_rst(config_rst)); 
mux6 mux_2866 (.in({n11665_1, n11664_0, n11657_0, n11656_0, n11649_0, n11648_0}), .out(n6083), .config_in(config_chain[8600:8598]), .config_rst(config_rst)); 
mux6 mux_2867 (.in({n13789_0, n13788_0, n13781_0, n13780_0, n13773_0, n13772_0}), .out(n6084), .config_in(config_chain[8603:8601]), .config_rst(config_rst)); 
mux6 mux_2868 (.in({n11907_0, n11906_0, n11893_0, n11892_0, n11877_0, n11876_1}), .out(n6085), .config_in(config_chain[8606:8604]), .config_rst(config_rst)); 
mux6 mux_2869 (.in({n14025_0, n14024_0, n14019_0, n14018_0, n14011_0, n14010_0}), .out(n6086), .config_in(config_chain[8609:8607]), .config_rst(config_rst)); 
mux6 mux_2870 (.in({n11681_1, n11680_0, n11607_0, n11606_1, n11599_0, n11598_1}), .out(n6087), .config_in(config_chain[8612:8610]), .config_rst(config_rst)); 
mux6 mux_2871 (.in({n13797_0, n13796_0, n13737_0, n13736_0, n13723_0, n13722_1}), .out(n6088), .config_in(config_chain[8615:8613]), .config_rst(config_rst)); 
mux6 mux_2872 (.in({n11929_1, n11928_0, n11923_0, n11922_0/**/, n11915_0, n11914_0}), .out(n6089), .config_in(config_chain[8618:8616]), .config_rst(config_rst)); 
mux6 mux_2873 (.in({n14047_0, n14046_0, n14041_0, n14040_0/**/, n14033_0, n14032_0}), .out(n6090), .config_in(config_chain[8621:8619]), .config_rst(config_rst)); 
mux6 mux_2874 (.in({n11629_0, n11628_0, n11621_0, n11620_0, n11615_0, n11614_1}), .out(n6091), .config_in(config_chain[8624:8622]), .config_rst(config_rst)); 
mux6 mux_2875 (.in({n13759_0, n13758_0, n13745_0, n13744_0, n13731_0, n13730_1}), .out(n6092), .config_in(config_chain[8627:8625]), .config_rst(config_rst)); 
mux6 mux_2876 (.in({n11945_1, n11944_0, n11937_1, n11936_0/**/, n11863_0, n11862_1}), .out(n6093), .config_in(config_chain[8630:8628]), .config_rst(config_rst)); 
mux6 mux_2877 (.in({n14063_0, n14062_0, n13989_0/**/, n13988_1, n13981_0, n13980_1}), .out(n6094), .config_in(config_chain[8633:8631]), .config_rst(config_rst)); 
mux6 mux_2878 (.in({n11667_1, n11666_0/**/, n11651_0, n11650_0, n11637_0, n11636_0}), .out(n6095), .config_in(config_chain[8636:8634]), .config_rst(config_rst)); 
mux6 mux_2879 (.in({n13783_0, n13782_0, n13775_0, n13774_0, n13767_0, n13766_0}), .out(n6096), .config_in(config_chain[8639:8637]), .config_rst(config_rst)); 
mux6 mux_2880 (.in({n11895_0, n11894_0, n11887_0, n11886_0/**/, n11879_0, n11878_1}), .out(n6097), .config_in(config_chain[8642:8640]), .config_rst(config_rst)); 
mux6 mux_2881 (.in({n14027_0, n14026_0/**/, n14013_0, n14012_0, n13997_0, n13996_1}), .out(n6098), .config_in(config_chain[8645:8643]), .config_rst(config_rst)); 
mux6 mux_2882 (.in({n11675_1, n11674_0, n11659_0/**/, n11658_0, n11601_0, n11600_1}), .out(n6099), .config_in(config_chain[8648:8646]), .config_rst(config_rst)); 
mux6 mux_2883 (.in({n13799_0/**/, n13798_0, n13791_0, n13790_0, n13717_0, n13716_1}), .out(n6100), .config_in(config_chain[8651:8649]), .config_rst(config_rst)); 
mux6 mux_2884 (.in({n11917_0, n11916_0, n11909_0, n11908_0, n11903_0, n11902_0}), .out(n6101), .config_in(config_chain[8654:8652]), .config_rst(config_rst)); 
mux6 mux_2885 (.in({n14049_0, n14048_0, n14035_0, n14034_0/**/, n14021_0, n14020_0}), .out(n6102), .config_in(config_chain[8657:8655]), .config_rst(config_rst)); 
mux6 mux_2886 (.in({n11623_0, n11622_0, n11617_0, n11616_1, n11609_0, n11608_1/**/}), .out(n6103), .config_in(config_chain[8660:8658]), .config_rst(config_rst)); 
mux6 mux_2887 (.in({n13747_0, n13746_0, n13739_0, n13738_0, n13733_0, n13732_1}), .out(n6104), .config_in(config_chain[8663:8661]), .config_rst(config_rst)); 
mux6 mux_2888 (.in({n11939_1, n11938_0, n11925_0, n11924_0, n11865_0/**/, n11864_1}), .out(n6105), .config_in(config_chain[8666:8664]), .config_rst(config_rst)); 
mux6 mux_2889 (.in({n14065_0, n14064_0/**/, n14057_0, n14056_0, n13983_0, n13982_1}), .out(n6106), .config_in(config_chain[8669:8667]), .config_rst(config_rst)); 
mux6 mux_2890 (.in({n11653_0, n11652_0, n11645_0, n11644_0, n11639_0/**/, n11638_0}), .out(n6107), .config_in(config_chain[8672:8670]), .config_rst(config_rst)); 
mux6 mux_2891 (.in({n13769_0, n13768_0, n13761_0, n13760_0, n13755_0/**/, n13754_0}), .out(n6108), .config_in(config_chain[8675:8673]), .config_rst(config_rst)); 
mux6 mux_2892 (.in({n11947_1/**/, n11946_0, n11889_0, n11888_0, n11873_0, n11872_1}), .out(n6109), .config_in(config_chain[8678:8676]), .config_rst(config_rst)); 
mux6 mux_2893 (.in({n14007_0, n14006_0, n13999_0, n13998_1, n13991_0, n13990_1}), .out(n6110), .config_in(config_chain[8681:8679]), .config_rst(config_rst)); 
mux6 mux_2894 (.in({n11677_1/**/, n11676_0, n11669_1, n11668_0, n11661_0, n11660_0}), .out(n6111), .config_in(config_chain[8684:8682]), .config_rst(config_rst)); 
mux6 mux_2895 (.in({n13793_0, n13792_0, n13777_0/**/, n13776_0, n13719_0, n13718_1}), .out(n6112), .config_in(config_chain[8687:8685]), .config_rst(config_rst)); 
mux6 mux_2896 (.in({n11949_1, n11948_0, n11911_0, n11910_0/**/, n11897_0, n11896_0}), .out(n6113), .config_in(config_chain[8690:8688]), .config_rst(config_rst)); 
mux6 mux_2897 (.in({n14067_0, n14066_0, n14037_0, n14036_0/**/, n14029_0, n14028_0}), .out(n6114), .config_in(config_chain[8693:8691]), .config_rst(config_rst)); 
mux6 mux_2898 (.in({n11625_0, n11624_0, n11611_0/**/, n11610_1, n11597_1, n11596_1}), .out(n6115), .config_in(config_chain[8696:8694]), .config_rst(config_rst)); 
mux6 mux_2899 (.in({n13741_0, n13740_0, n13727_0, n13726_1, n13713_0, n13712_1}), .out(n6116), .config_in(config_chain[8699:8697]), .config_rst(config_rst)); 
mux6 mux_2900 (.in({n11933_1, n11932_0, n11919_0, n11918_0, n11829_1, n11828_1}), .out(n6117), .config_in(config_chain[8702:8700]), .config_rst(config_rst)); 
mux6 mux_2901 (.in({n14059_0, n14058_0, n14051_0, n14050_0/**/, n13957_0, n13956_1}), .out(n6118), .config_in(config_chain[8705:8703]), .config_rst(config_rst)); 
mux6 mux_2902 (.in({n11647_0, n11646_0, n11633_0, n11632_0, n11619_1, n11618_1}), .out(n6119), .config_in(config_chain[8708:8706]), .config_rst(config_rst)); 
mux6 mux_2903 (.in({n13763_0, n13762_0, n13757_0, n13756_0, n13749_0/**/, n13748_0}), .out(n6120), .config_in(config_chain[8711:8709]), .config_rst(config_rst)); 
mux6 mux_2904 (.in({n11875_0/**/, n11874_1, n11867_0, n11866_1, n11861_1, n11860_1}), .out(n6121), .config_in(config_chain[8714:8712]), .config_rst(config_rst)); 
mux6 mux_2905 (.in({n14009_0, n14008_0, n13993_0, n13992_1, n13979_0, n13978_1}), .out(n6122), .config_in(config_chain[8717:8715]), .config_rst(config_rst)); 
mux6 mux_2906 (.in({n11671_1, n11670_0, n11663_1, n11662_0, n11655_0, n11654_0/**/}), .out(n6123), .config_in(config_chain[8720:8718]), .config_rst(config_rst)); 
mux6 mux_2907 (.in({n13795_0, n13794_0/**/, n13787_0, n13786_0, n13779_0, n13778_0}), .out(n6124), .config_in(config_chain[8723:8721]), .config_rst(config_rst)); 
mux6 mux_2908 (.in({n11899_0, n11898_0, n11891_0, n11890_0, n11883_1, n11882_1}), .out(n6125), .config_in(config_chain[8726:8724]), .config_rst(config_rst)); 
mux6 mux_2909 (.in({n14031_0, n14030_0, n14017_0, n14016_0, n14001_0, n14000_1}), .out(n6126), .config_in(config_chain[8729:8727]), .config_rst(config_rst)); 
mux6 mux_2910 (.in({n11685_1, n11684_0, n11679_1, n11678_0, n11605_0/**/, n11604_1}), .out(n6127), .config_in(config_chain[8732:8730]), .config_rst(config_rst)); 
mux6 mux_2911 (.in({n13801_0, n13800_0, n13729_0, n13728_1/**/, n13721_0, n13720_1}), .out(n6128), .config_in(config_chain[8735:8733]), .config_rst(config_rst)); 
mux6 mux_2912 (.in({n11935_1, n11934_0, n11921_0, n11920_0, n11905_1, n11904_0}), .out(n6129), .config_in(config_chain[8738:8736]), .config_rst(config_rst)); 
mux6 mux_2913 (.in({n14053_0, n14052_0, n14045_0, n14044_0, n14039_0, n14038_0/**/}), .out(n6130), .config_in(config_chain[8741:8739]), .config_rst(config_rst)); 
mux6 mux_2914 (.in({n11635_0, n11634_0/**/, n11627_0, n11626_0, n11575_0, n11574_1}), .out(n6131), .config_in(config_chain[8744:8742]), .config_rst(config_rst)); 
mux6 mux_2915 (.in({n13765_0, n13764_0/**/, n13751_0, n13750_0, n13651_0, n13650_2}), .out(n6132), .config_in(config_chain[8747:8745]), .config_rst(config_rst)); 
mux6 mux_2916 (.in({n12191_1, n12190_0, n12175_0, n12174_0, n12161_0, n12160_0}), .out(n6179), .config_in(config_chain[8750:8748]), .config_rst(config_rst)); 
mux6 mux_2917 (.in({n14069_0, n14068_0, n14053_0, n14052_0, n14039_0, n14038_0}), .out(n6180), .config_in(config_chain[8753:8751]), .config_rst(config_rst)); 
mux6 mux_2918 (.in({n11885_0, n11884_0, n11877_0, n11876_1, n11869_0, n11868_1}), .out(n6181), .config_in(config_chain[8756:8754]), .config_rst(config_rst)); 
mux6 mux_2919 (.in({n13767_0, n13766_0, n13759_0, n13758_0, n13751_0, n13750_1}), .out(n6182), .config_in(config_chain[8759:8757]), .config_rst(config_rst)); 
mux6 mux_2920 (.in({n12199_1, n12198_0, n12183_0, n12182_0, n12125_0, n12124_1}), .out(n6183), .config_in(config_chain[8762:8760]), .config_rst(config_rst)); 
mux6 mux_2921 (.in({n14085_0, n14084_0, n14077_0, n14076_0, n14003_0, n14002_1}), .out(n6184), .config_in(config_chain[8765:8763]), .config_rst(config_rst)); 
mux6 mux_2922 (.in({n11915_0, n11914_0, n11907_0, n11906_0, n11901_0, n11900_0}), .out(n6185), .config_in(config_chain[8768:8766]), .config_rst(config_rst)); 
mux6 mux_2923 (.in({n13803_0, n13802_0, n13789_0, n13788_0, n13775_0, n13774_0/**/}), .out(n6186), .config_in(config_chain[8771:8769]), .config_rst(config_rst)); 
mux6 mux_2924 (.in({n12147_0, n12146_0, n12141_0, n12140_1, n12133_0, n12132_1/**/}), .out(n6187), .config_in(config_chain[8774:8772]), .config_rst(config_rst)); 
mux6 mux_2925 (.in({n14025_0, n14024_0, n14019_0, n14018_1, n14011_0, n14010_1}), .out(n6188), .config_in(config_chain[8777:8775]), .config_rst(config_rst)); 
mux6 mux_2926 (.in({n11937_1, n11936_0, n11929_1, n11928_0, n11923_0, n11922_0}), .out(n6189), .config_in(config_chain[8780:8778]), .config_rst(config_rst)); 
mux6 mux_2927 (.in({n13811_0/**/, n13810_0, n13797_0, n13796_0, n13737_0, n13736_1}), .out(n6190), .config_in(config_chain[8783:8781]), .config_rst(config_rst)); 
mux6 mux_2928 (.in({n12169_0, n12168_0, n12163_0, n12162_0, n12155_0, n12154_0}), .out(n6191), .config_in(config_chain[8786:8784]), .config_rst(config_rst)); 
mux6 mux_2929 (.in({n14055_0, n14054_0, n14047_0, n14046_0/**/, n14041_0, n14040_0}), .out(n6192), .config_in(config_chain[8789:8787]), .config_rst(config_rst)); 
mux6 mux_2930 (.in({n11945_1, n11944_0, n11887_0, n11886_0, n11871_0/**/, n11870_1}), .out(n6193), .config_in(config_chain[8792:8790]), .config_rst(config_rst)); 
mux6 mux_2931 (.in({n13761_0, n13760_0, n13753_0, n13752_1/**/, n13745_0, n13744_1}), .out(n6194), .config_in(config_chain[8795:8793]), .config_rst(config_rst)); 
mux6 mux_2932 (.in({n12201_1, n12200_0, n12193_1, n12192_0, n12185_0/**/, n12184_0}), .out(n6195), .config_in(config_chain[8798:8796]), .config_rst(config_rst)); 
mux6 mux_2933 (.in({n14079_0, n14078_0, n14063_0, n14062_0, n14005_0, n14004_1}), .out(n6196), .config_in(config_chain[8801:8799]), .config_rst(config_rst)); 
mux6 mux_2934 (.in({n11909_0, n11908_0, n11895_0, n11894_0, n11879_0, n11878_1}), .out(n6197), .config_in(config_chain[8804:8802]), .config_rst(config_rst)); 
mux6 mux_2935 (.in({n13783_0, n13782_0/**/, n13777_0, n13776_0, n13769_0, n13768_0}), .out(n6198), .config_in(config_chain[8807:8805]), .config_rst(config_rst)); 
mux6 mux_2936 (.in({n12209_1, n12208_0, n12135_0, n12134_1, n12127_0/**/, n12126_1}), .out(n6199), .config_in(config_chain[8810:8808]), .config_rst(config_rst)); 
mux6 mux_2937 (.in({n14087_0/**/, n14086_0, n14027_0, n14026_0, n14013_0, n14012_1}), .out(n6200), .config_in(config_chain[8813:8811]), .config_rst(config_rst)); 
mux6 mux_2938 (.in({n11931_1, n11930_0, n11925_0, n11924_0, n11917_0, n11916_0}), .out(n6201), .config_in(config_chain[8816:8814]), .config_rst(config_rst)); 
mux6 mux_2939 (.in({n13813_0, n13812_0/**/, n13805_0, n13804_0, n13799_0, n13798_0}), .out(n6202), .config_in(config_chain[8819:8817]), .config_rst(config_rst)); 
mux6 mux_2940 (.in({n12171_0, n12170_0, n12157_0, n12156_0, n12143_0, n12142_1/**/}), .out(n6203), .config_in(config_chain[8822:8820]), .config_rst(config_rst)); 
mux6 mux_2941 (.in({n14049_0, n14048_0/**/, n14043_0, n14042_0, n14035_0, n14034_0}), .out(n6204), .config_in(config_chain[8825:8823]), .config_rst(config_rst)); 
mux6 mux_2942 (.in({n11947_1/**/, n11946_0, n11873_0, n11872_1, n11865_0, n11864_1}), .out(n6205), .config_in(config_chain[8828:8826]), .config_rst(config_rst)); 
mux6 mux_2943 (.in({n13821_0, n13820_0, n13747_0, n13746_1, n13739_0/**/, n13738_1}), .out(n6206), .config_in(config_chain[8831:8829]), .config_rst(config_rst)); 
mux6 mux_2944 (.in({n12195_1, n12194_0, n12179_0, n12178_0, n12165_0, n12164_0/**/}), .out(n6207), .config_in(config_chain[8834:8832]), .config_rst(config_rst)); 
mux6 mux_2945 (.in({n14073_0, n14072_0, n14065_0, n14064_0, n14057_0, n14056_0}), .out(n6208), .config_in(config_chain[8837:8835]), .config_rst(config_rst)); 
mux6 mux_2946 (.in({n11897_0, n11896_0, n11889_0, n11888_0, n11881_0, n11880_1}), .out(n6209), .config_in(config_chain[8840:8838]), .config_rst(config_rst)); 
mux6 mux_2947 (.in({n13785_0, n13784_0, n13771_0, n13770_0, n13755_0, n13754_1/**/}), .out(n6210), .config_in(config_chain[8843:8841]), .config_rst(config_rst)); 
mux6 mux_2948 (.in({n12203_1, n12202_0, n12167_1, n12166_0, n12129_0/**/, n12128_1}), .out(n6211), .config_in(config_chain[8846:8844]), .config_rst(config_rst)); 
mux6 mux_2949 (.in({n14045_0, n14044_0, n14015_0, n14014_1, n14007_0, n14006_1}), .out(n6212), .config_in(config_chain[8849:8847]), .config_rst(config_rst)); 
mux6 mux_2950 (.in({n11949_1, n11948_0, n11933_1, n11932_0, n11919_0, n11918_0}), .out(n6213), .config_in(config_chain[8852:8850]), .config_rst(config_rst)); 
mux6 mux_2951 (.in({n13823_0, n13822_0, n13807_0, n13806_0, n13793_0, n13792_0}), .out(n6214), .config_in(config_chain[8855:8853]), .config_rst(config_rst)); 
mux6 mux_2952 (.in({n12189_1, n12188_0, n12151_0, n12150_0/**/, n12137_0, n12136_1}), .out(n6215), .config_in(config_chain[8858:8856]), .config_rst(config_rst)); 
mux6 mux_2953 (.in({n14067_0, n14066_0, n14037_0, n14036_0, n14029_0, n14028_0}), .out(n6216), .config_in(config_chain[8861:8859]), .config_rst(config_rst)); 
mux6 mux_2954 (.in({n11941_1, n11940_0/**/, n11867_0, n11866_1, n11829_1, n11828_1}), .out(n6217), .config_in(config_chain[8864:8862]), .config_rst(config_rst)); 
mux6 mux_2955 (.in({n13815_0, n13814_0, n13741_0/**/, n13740_1, n13735_0, n13734_1}), .out(n6218), .config_in(config_chain[8867:8865]), .config_rst(config_rst)); 
mux6 mux_2956 (.in({n12181_0, n12180_0/**/, n12173_0, n12172_0, n12091_1, n12090_1}), .out(n6219), .config_in(config_chain[8870:8868]), .config_rst(config_rst)); 
mux6 mux_2957 (.in({n14075_0, n14074_0, n14059_0, n14058_0, n13957_0, n13956_2/**/}), .out(n6220), .config_in(config_chain[8873:8871]), .config_rst(config_rst)); 
mux6 mux_2958 (.in({n11891_0, n11890_0, n11883_1/**/, n11882_1, n11875_0, n11874_1}), .out(n6221), .config_in(config_chain[8876:8874]), .config_rst(config_rst)); 
mux6 mux_2959 (.in({n13773_0, n13772_0, n13765_0, n13764_0, n13757_0, n13756_1}), .out(n6222), .config_in(config_chain[8879:8877]), .config_rst(config_rst)); 
mux6 mux_2960 (.in({n12205_1, n12204_0, n12197_1, n12196_0/**/, n12093_1, n12092_1}), .out(n6223), .config_in(config_chain[8882:8880]), .config_rst(config_rst)); 
mux6 mux_2961 (.in({n14083_0, n14082_0, n14009_0, n14008_1/**/, n13979_0, n13978_1}), .out(n6224), .config_in(config_chain[8885:8883]), .config_rst(config_rst)); 
mux6 mux_2962 (.in({n11913_0, n11912_0, n11905_1, n11904_0, n11899_0, n11898_0}), .out(n6225), .config_in(config_chain[8888:8886]), .config_rst(config_rst)); 
mux6 mux_2963 (.in({n13795_0, n13794_0, n13787_0, n13786_0, n13779_0, n13778_0}), .out(n6226), .config_in(config_chain[8891:8889]), .config_rst(config_rst)); 
mux6 mux_2964 (.in({n12153_0, n12152_0, n12139_0, n12138_1/**/, n12123_1, n12122_1}), .out(n6227), .config_in(config_chain[8894:8892]), .config_rst(config_rst)); 
mux6 mux_2965 (.in({n14031_0, n14030_0, n14023_0, n14022_1/**/, n14017_0, n14016_1}), .out(n6228), .config_in(config_chain[8897:8895]), .config_rst(config_rst)); 
mux6 mux_2966 (.in({n11943_1, n11942_0, n11935_1, n11934_0/**/, n11927_1, n11926_0}), .out(n6229), .config_in(config_chain[8900:8898]), .config_rst(config_rst)); 
mux6 mux_2967 (.in({n13817_0, n13816_0, n13801_0, n13800_0/**/, n13743_0, n13742_1}), .out(n6230), .config_in(config_chain[8903:8901]), .config_rst(config_rst)); 
mux6 mux_2968 (.in({n12199_1, n12198_0, n12191_1, n12190_0, n12183_0, n12182_0}), .out(n6276), .config_in(config_chain[8906:8904]), .config_rst(config_rst)); 
mux6 mux_2969 (.in({n12155_0, n12154_0, n12147_0, n12146_0, n12141_0, n12140_1}), .out(n6279), .config_in(config_chain[8909:8907]), .config_rst(config_rst)); 
mux6 mux_2970 (.in({n12201_1, n12200_0, n12193_1, n12192_0, n12185_0, n12184_0}), .out(n6282), .config_in(config_chain[8912:8910]), .config_rst(config_rst)); 
mux6 mux_2971 (.in({n12157_0, n12156_0, n12149_0, n12148_0, n12143_0, n12142_1}), .out(n6285), .config_in(config_chain[8915:8913]), .config_rst(config_rst)); 
mux6 mux_2972 (.in({n12195_1, n12194_0, n12187_0, n12186_0, n12179_0, n12178_0}), .out(n6288), .config_in(config_chain[8918:8916]), .config_rst(config_rst)); 
mux6 mux_2973 (.in({n12189_1, n12188_0, n12151_0, n12150_0, n12137_0, n12136_1}), .out(n6291), .config_in(config_chain[8921:8919]), .config_rst(config_rst)); 
mux6 mux_2974 (.in({n12197_1, n12196_0, n12181_0, n12180_0, n12093_1, n12092_1}), .out(n6294), .config_in(config_chain[8924:8922]), .config_rst(config_rst)); 
mux6 mux_2975 (.in({n12153_0, n12152_0, n12145_1, n12144_1, n12139_0, n12138_1}), .out(n6297), .config_in(config_chain[8927:8925]), .config_rst(config_rst)); 
mux6 mux_2976 (.in({n9859_0, n9858_0, n9845_0, n9844_0, n9833_0, n9832_0}), .out(n6324), .config_in(config_chain[8930:8928]), .config_rst(config_rst)); 
mux6 mux_2977 (.in({n9875_0, n9874_0, n9807_0, n9806_1, n9799_0, n9798_1}), .out(n6327), .config_in(config_chain[8933:8931]), .config_rst(config_rst)); 
mux6 mux_2978 (.in({n9847_0, n9846_0, n9839_0, n9838_0, n9835_0, n9834_0}), .out(n6330), .config_in(config_chain[8936:8934]), .config_rst(config_rst)); 
mux6 mux_2979 (.in({n9877_0, n9876_0, n9809_0, n9808_1, n9801_0, n9800_1}), .out(n6333), .config_in(config_chain[8939:8937]), .config_rst(config_rst)); 
mux6 mux_2980 (.in({n9849_0, n9848_0, n9841_0, n9840_0, n9837_0, n9836_0}), .out(n6336), .config_in(config_chain[8942:8940]), .config_rst(config_rst)); 
mux6 mux_2981 (.in({n9871_0, n9870_0, n9803_0, n9802_1, n9747_0, n9746_2}), .out(n6339), .config_in(config_chain[8945:8943]), .config_rst(config_rst)); 
mux6 mux_2982 (.in({n9843_0, n9842_0, n9831_0, n9830_0, n9751_0, n9750_2}), .out(n6342), .config_in(config_chain[8948:8946]), .config_rst(config_rst)); 
mux6 mux_2983 (.in({n9873_0, n9872_0, n9805_0, n9804_1, n9755_0, n9754_2}), .out(n6345), .config_in(config_chain[8951:8949]), .config_rst(config_rst)); 
mux6 mux_2984 (.in({n10127_0, n10126_0, n10073_0, n10072_0/**/, n10059_0, n10058_1}), .out(n6373), .config_in(config_chain[8954:8952]), .config_rst(config_rst)); 
mux6 mux_2985 (.in({n14151_1, n14150_0, n14113_0, n14112_0, n14091_0, n14090_0}), .out(n6374), .config_in(config_chain[8957:8955]), .config_rst(config_rst)); 
mux6 mux_2986 (.in({n9859_0, n9858_0, n9853_0, n9852_0, n9845_0, n9844_0}), .out(n6375), .config_in(config_chain[8960:8958]), .config_rst(config_rst)); 
mux6 mux_2987 (.in({n13883_0, n13882_0, n13861_1, n13860_0, n13829_1, n13828_0}), .out(n6376), .config_in(config_chain[8963:8961]), .config_rst(config_rst)); 
mux6 mux_2988 (.in({n10093_0, n10092_0, n10081_0, n10080_0, n10067_0, n10066_1}), .out(n6377), .config_in(config_chain[8966:8964]), .config_rst(config_rst)); 
mux6 mux_2989 (.in({n14155_0, n14154_0, n14123_0, n14122_0, n14093_0, n14092_0}), .out(n6378), .config_in(config_chain[8969:8967]), .config_rst(config_rst)); 
mux6 mux_2990 (.in({n9875_0, n9874_0, n9807_0, n9806_1/**/, n9799_0, n9798_1}), .out(n6379), .config_in(config_chain[8972:8970]), .config_rst(config_rst)); 
mux6 mux_2991 (.in({n13893_1, n13892_0, n13863_0, n13862_0, n13825_0/**/, n13824_0}), .out(n6380), .config_in(config_chain[8975:8973]), .config_rst(config_rst)); 
mux6 mux_2992 (.in({n10113_0, n10112_0, n10109_0, n10108_0, n10101_0, n10100_0}), .out(n6381), .config_in(config_chain[8978:8976]), .config_rst(config_rst)); 
mux6 mux_2993 (.in({n14157_0, n14156_0, n14125_0, n14124_0/**/, n14095_1, n14094_0}), .out(n6382), .config_in(config_chain[8981:8979]), .config_rst(config_rst)); 
mux6 mux_2994 (.in({n9827_0, n9826_0, n9819_0, n9818_0/**/, n9815_0, n9814_1}), .out(n6383), .config_in(config_chain[8984:8982]), .config_rst(config_rst)); 
mux6 mux_2995 (.in({n13895_0, n13894_0, n13857_0, n13856_0, n13827_0, n13826_0}), .out(n6384), .config_in(config_chain[8987:8985]), .config_rst(config_rst)); 
mux6 mux_2996 (.in({n10129_0, n10128_0, n10121_0, n10120_0, n10053_0, n10052_1}), .out(n6385), .config_in(config_chain[8990:8988]), .config_rst(config_rst)); 
mux6 mux_2997 (.in({n14159_1, n14158_0, n14121_0, n14120_0, n14089_0/**/, n14088_0}), .out(n6386), .config_in(config_chain[8993:8991]), .config_rst(config_rst)); 
mux6 mux_2998 (.in({n9861_0, n9860_0, n9847_0, n9846_0, n9835_0, n9834_0}), .out(n6387), .config_in(config_chain[8996:8994]), .config_rst(config_rst)); 
mux6 mux_2999 (.in({n13891_0, n13890_0, n13859_0, n13858_0, n13837_1, n13836_0}), .out(n6388), .config_in(config_chain[8999:8997]), .config_rst(config_rst)); 
mux6 mux_3000 (.in({n10083_0, n10082_0/**/, n10075_0, n10074_0, n10069_0, n10068_1}), .out(n6389), .config_in(config_chain[9002:9000]), .config_rst(config_rst)); 
mux6 mux_3001 (.in({n14153_0, n14152_0, n14131_0, n14130_0, n14101_0, n14100_0}), .out(n6390), .config_in(config_chain[9005:9003]), .config_rst(config_rst)); 
mux6 mux_3002 (.in({n9869_0, n9868_0, n9855_0, n9854_0, n9801_0, n9800_1}), .out(n6391), .config_in(config_chain[9008:9006]), .config_rst(config_rst)); 
mux6 mux_3003 (.in({n13901_1, n13900_0, n13869_1, n13868_0, n13839_0, n13838_0}), .out(n6392), .config_in(config_chain[9011:9009]), .config_rst(config_rst)); 
mux6 mux_3004 (.in({n10103_0, n10102_0, n10095_0, n10094_0, n10091_0, n10090_0/**/}), .out(n6393), .config_in(config_chain[9014:9012]), .config_rst(config_rst)); 
mux6 mux_3005 (.in({n14163_0, n14162_0, n14133_0, n14132_0, n14103_1, n14102_0}), .out(n6394), .config_in(config_chain[9017:9015]), .config_rst(config_rst)); 
mux6 mux_3006 (.in({n9821_0, n9820_0, n9817_0/**/, n9816_1, n9809_0, n9808_1}), .out(n6395), .config_in(config_chain[9020:9018]), .config_rst(config_rst)); 
mux6 mux_3007 (.in({n13903_0/**/, n13902_0, n13865_0, n13864_0, n13833_0, n13832_0}), .out(n6396), .config_in(config_chain[9023:9021]), .config_rst(config_rst)); 
mux6 mux_3008 (.in({n10123_0, n10122_0/**/, n10111_0, n10110_0, n10055_0, n10054_1}), .out(n6397), .config_in(config_chain[9026:9024]), .config_rst(config_rst)); 
mux6 mux_3009 (.in({n14167_1, n14166_0, n14135_1/**/, n14134_0, n14097_0, n14096_0}), .out(n6398), .config_in(config_chain[9029:9027]), .config_rst(config_rst)); 
mux6 mux_3010 (.in({n9849_0, n9848_0, n9841_0, n9840_0, n9837_0, n9836_0}), .out(n6399), .config_in(config_chain[9032:9030]), .config_rst(config_rst)); 
mux6 mux_3011 (.in({n13897_0, n13896_0, n13867_0, n13866_0, n13835_0, n13834_0}), .out(n6400), .config_in(config_chain[9035:9033]), .config_rst(config_rst)); 
mux6 mux_3012 (.in({n10131_0, n10130_0, n10077_0, n10076_0, n10063_0, n10062_1}), .out(n6401), .config_in(config_chain[9038:9036]), .config_rst(config_rst)); 
mux6 mux_3013 (.in({n14161_0, n14160_0, n14129_0, n14128_0, n14107_0, n14106_0}), .out(n6402), .config_in(config_chain[9041:9039]), .config_rst(config_rst)); 
mux6 mux_3014 (.in({n9871_0, n9870_0, n9863_0, n9862_0, n9857_0, n9856_0/**/}), .out(n6403), .config_in(config_chain[9044:9042]), .config_rst(config_rst)); 
mux6 mux_3015 (.in({n13899_0, n13898_0, n13877_1, n13876_0, n13847_0/**/, n13846_0}), .out(n6404), .config_in(config_chain[9047:9045]), .config_rst(config_rst)); 
mux6 mux_3016 (.in({n10097_0, n10096_0, n10085_0/**/, n10084_0, n10011_0, n10010_2}), .out(n6405), .config_in(config_chain[9050:9048]), .config_rst(config_rst)); 
mux6 mux_3017 (.in({n14179_1, n14178_0, n14141_0/**/, n14140_0, n14109_0, n14108_0}), .out(n6406), .config_in(config_chain[9053:9051]), .config_rst(config_rst)); 
mux6 mux_3018 (.in({n9823_0/**/, n9822_0, n9811_0, n9810_1, n9747_0, n9746_2}), .out(n6407), .config_in(config_chain[9056:9054]), .config_rst(config_rst)); 
mux6 mux_3019 (.in({n13905_0, n13904_0, n13879_0, n13878_0, n13841_0, n13840_0/**/}), .out(n6408), .config_in(config_chain[9059:9057]), .config_rst(config_rst)); 
mux6 mux_3020 (.in({n10117_0, n10116_0, n10105_0, n10104_0/**/, n10001_0, n10000_2}), .out(n6409), .config_in(config_chain[9062:9060]), .config_rst(config_rst)); 
mux6 mux_3021 (.in({n14169_0, n14168_0, n14143_1, n14142_0, n14111_1, n14110_0}), .out(n6410), .config_in(config_chain[9065:9063]), .config_rst(config_rst)); 
mux6 mux_3022 (.in({n9843_0, n9842_0, n9831_0, n9830_0, n9749_0, n9748_2}), .out(n6411), .config_in(config_chain[9068:9066]), .config_rst(config_rst)); 
mux6 mux_3023 (.in({n13909_1, n13908_0, n13873_0, n13872_0/**/, n13843_0, n13842_0}), .out(n6412), .config_in(config_chain[9071:9069]), .config_rst(config_rst)); 
mux6 mux_3024 (.in({n10065_0, n10064_1, n10057_0, n10056_1, n10003_0, n10002_2}), .out(n6413), .config_in(config_chain[9074:9072]), .config_rst(config_rst)); 
mux6 mux_3025 (.in({n14171_0, n14170_0, n14137_0/**/, n14136_0, n14115_0, n14114_0}), .out(n6414), .config_in(config_chain[9077:9075]), .config_rst(config_rst)); 
mux6 mux_3026 (.in({n9865_0, n9864_0/**/, n9851_0, n9850_0, n9753_0, n9752_2}), .out(n6415), .config_in(config_chain[9080:9078]), .config_rst(config_rst)); 
mux6 mux_3027 (.in({n13911_1, n13910_0, n13885_1, n13884_0, n13853_1, n13852_0}), .out(n6416), .config_in(config_chain[9083:9081]), .config_rst(config_rst)); 
mux6 mux_3028 (.in({n10087_0, n10086_0, n10079_0, n10078_0, n10005_0, n10004_2}), .out(n6417), .config_in(config_chain[9086:9084]), .config_rst(config_rst)); 
mux6 mux_3029 (.in({n14173_0, n14172_0, n14147_0/**/, n14146_0, n14117_0, n14116_0}), .out(n6418), .config_in(config_chain[9089:9087]), .config_rst(config_rst)); 
mux6 mux_3030 (.in({n9873_0, n9872_0, n9805_0, n9804_1, n9755_0, n9754_2}), .out(n6419), .config_in(config_chain[9092:9090]), .config_rst(config_rst)); 
mux6 mux_3031 (.in({n13913_1, n13912_0, n13887_0, n13886_0, n13855_0, n13854_0}), .out(n6420), .config_in(config_chain[9095:9093]), .config_rst(config_rst)); 
mux6 mux_3032 (.in({n10119_0, n10118_0, n10107_0, n10106_0, n10007_0, n10006_2}), .out(n6421), .config_in(config_chain[9098:9096]), .config_rst(config_rst)); 
mux6 mux_3033 (.in({n14177_1, n14176_0, n14149_0, n14148_0, n14119_1, n14118_0}), .out(n6422), .config_in(config_chain[9101:9099]), .config_rst(config_rst)); 
mux6 mux_3034 (.in({n9833_0, n9832_0/**/, n9825_0, n9824_0, n9757_0, n9756_2}), .out(n6423), .config_in(config_chain[9104:9102]), .config_rst(config_rst)); 
mux6 mux_3035 (.in({n13915_2, n13914_0, n13881_0, n13880_0, n13851_0, n13850_0}), .out(n6424), .config_in(config_chain[9107:9105]), .config_rst(config_rst)); 
mux6 mux_3036 (.in({n10369_0, n10368_0, n10355_0, n10354_0, n10343_0, n10342_0/**/}), .out(n6471), .config_in(config_chain[9110:9108]), .config_rst(config_rst)); 
mux6 mux_3037 (.in({n14181_1, n14180_0, n14149_0, n14148_0, n14119_0, n14118_0}), .out(n6472), .config_in(config_chain[9113:9111]), .config_rst(config_rst)); 
mux6 mux_3038 (.in({n10073_0, n10072_0, n10067_0, n10066_1/**/, n10059_0, n10058_1}), .out(n6473), .config_in(config_chain[9116:9114]), .config_rst(config_rst)); 
mux6 mux_3039 (.in({n13881_0, n13880_0, n13859_0/**/, n13858_0, n13827_0, n13826_0}), .out(n6474), .config_in(config_chain[9119:9117]), .config_rst(config_rst)); 
mux6 mux_3040 (.in({n10377_0, n10376_0, n10363_0, n10362_0, n10309_0, n10308_1}), .out(n6475), .config_in(config_chain[9122:9120]), .config_rst(config_rst)); 
mux6 mux_3041 (.in({n14197_1, n14196_0, n14189_1, n14188_0, n14091_0, n14090_0}), .out(n6476), .config_in(config_chain[9125:9123]), .config_rst(config_rst)); 
mux6 mux_3042 (.in({n10101_0, n10100_0, n10093_0, n10092_0, n10089_0, n10088_0}), .out(n6477), .config_in(config_chain[9128:9126]), .config_rst(config_rst)); 
mux6 mux_3043 (.in({n13917_1, n13916_0, n13891_0, n13890_0, n13861_0, n13860_0}), .out(n6478), .config_in(config_chain[9131:9129]), .config_rst(config_rst)); 
mux6 mux_3044 (.in({n10329_0, n10328_0/**/, n10325_0, n10324_1, n10317_0, n10316_1}), .out(n6479), .config_in(config_chain[9134:9132]), .config_rst(config_rst)); 
mux6 mux_3045 (.in({n14155_0, n14154_0, n14123_0, n14122_0, n14093_0, n14092_0}), .out(n6480), .config_in(config_chain[9137:9135]), .config_rst(config_rst)); 
mux6 mux_3046 (.in({n10121_0, n10120_0, n10113_0, n10112_0, n10109_0, n10108_0}), .out(n6481), .config_in(config_chain[9140:9138]), .config_rst(config_rst)); 
mux6 mux_3047 (.in({n13925_1, n13924_0, n13893_0, n13892_0, n13825_0, n13824_0}), .out(n6482), .config_in(config_chain[9143:9141]), .config_rst(config_rst)); 
mux6 mux_3048 (.in({n10349_0, n10348_0, n10345_0, n10344_0, n10337_0, n10336_0}), .out(n6483), .config_in(config_chain[9146:9144]), .config_rst(config_rst)); 
mux6 mux_3049 (.in({n14157_0, n14156_0, n14127_0, n14126_0, n14095_0/**/, n14094_0}), .out(n6484), .config_in(config_chain[9149:9147]), .config_rst(config_rst)); 
mux6 mux_3050 (.in({n10129_0, n10128_0, n10075_0, n10074_0/**/, n10061_0, n10060_1}), .out(n6485), .config_in(config_chain[9152:9150]), .config_rst(config_rst)); 
mux6 mux_3051 (.in({n13889_0, n13888_0, n13857_0, n13856_0, n13835_0, n13834_0/**/}), .out(n6486), .config_in(config_chain[9155:9153]), .config_rst(config_rst)); 
mux6 mux_3052 (.in({n10379_0, n10378_0, n10371_0, n10370_0/**/, n10365_0, n10364_0}), .out(n6487), .config_in(config_chain[9158:9156]), .config_rst(config_rst)); 
mux6 mux_3053 (.in({n14191_1, n14190_0/**/, n14159_0, n14158_0, n14099_0, n14098_0}), .out(n6488), .config_in(config_chain[9161:9159]), .config_rst(config_rst)); 
mux6 mux_3054 (.in({n10095_0/**/, n10094_0, n10083_0, n10082_0, n10069_0, n10068_1}), .out(n6489), .config_in(config_chain[9164:9162]), .config_rst(config_rst)); 
mux6 mux_3055 (.in({n13899_0, n13898_0, n13867_0, n13866_0, n13837_0, n13836_0}), .out(n6490), .config_in(config_chain[9167:9165]), .config_rst(config_rst)); 
mux6 mux_3056 (.in({n10387_0, n10386_0/**/, n10319_0, n10318_1, n10311_0, n10310_1}), .out(n6491), .config_in(config_chain[9170:9168]), .config_rst(config_rst)); 
mux6 mux_3057 (.in({n14199_1, n14198_0, n14131_0, n14130_0, n14101_0/**/, n14100_0}), .out(n6492), .config_in(config_chain[9173:9171]), .config_rst(config_rst)); 
mux6 mux_3058 (.in({n10115_0, n10114_0/**/, n10111_0, n10110_0, n10103_0, n10102_0}), .out(n6493), .config_in(config_chain[9176:9174]), .config_rst(config_rst)); 
mux6 mux_3059 (.in({n13927_1, n13926_0, n13919_1, n13918_0, n13901_0, n13900_0}), .out(n6494), .config_in(config_chain[9179:9177]), .config_rst(config_rst)); 
mux6 mux_3060 (.in({n10351_0, n10350_0, n10339_0, n10338_0, n10327_0, n10326_1}), .out(n6495), .config_in(config_chain[9182:9180]), .config_rst(config_rst)); 
mux6 mux_3061 (.in({n14165_0, n14164_0, n14133_0, n14132_0, n14103_0, n14102_0}), .out(n6496), .config_in(config_chain[9185:9183]), .config_rst(config_rst)); 
mux6 mux_3062 (.in({n10131_0, n10130_0/**/, n10063_0, n10062_1, n10055_0, n10054_1}), .out(n6497), .config_in(config_chain[9188:9186]), .config_rst(config_rst)); 
mux6 mux_3063 (.in({n13935_1, n13934_0, n13865_0, n13864_0/**/, n13833_0, n13832_0}), .out(n6498), .config_in(config_chain[9191:9189]), .config_rst(config_rst)); 
mux6 mux_3064 (.in({n10373_0, n10372_0, n10359_0, n10358_0, n10347_0/**/, n10346_0}), .out(n6499), .config_in(config_chain[9194:9192]), .config_rst(config_rst)); 
mux6 mux_3065 (.in({n14185_1/**/, n14184_0, n14167_0, n14166_0, n14135_0, n14134_0}), .out(n6500), .config_in(config_chain[9197:9195]), .config_rst(config_rst)); 
mux6 mux_3066 (.in({n10085_0, n10084_0, n10077_0, n10076_0, n10071_0, n10070_1/**/}), .out(n6501), .config_in(config_chain[9200:9198]), .config_rst(config_rst)); 
mux6 mux_3067 (.in({n13897_0, n13896_0/**/, n13875_0, n13874_0, n13845_0, n13844_0}), .out(n6502), .config_in(config_chain[9203:9201]), .config_rst(config_rst)); 
mux6 mux_3068 (.in({n10381_0, n10380_0, n10313_0, n10312_1, n10265_0, n10264_2/**/}), .out(n6503), .config_in(config_chain[9206:9204]), .config_rst(config_rst)); 
mux6 mux_3069 (.in({n14177_1, n14176_0, n14139_0, n14138_0, n14107_0/**/, n14106_0}), .out(n6504), .config_in(config_chain[9209:9207]), .config_rst(config_rst)); 
mux6 mux_3070 (.in({n10117_0, n10116_0, n10105_0, n10104_0, n10011_0, n10010_2}), .out(n6505), .config_in(config_chain[9212:9210]), .config_rst(config_rst)); 
mux6 mux_3071 (.in({n13921_1, n13920_0, n13915_1, n13914_0, n13877_0, n13876_0}), .out(n6506), .config_in(config_chain[9215:9213]), .config_rst(config_rst)); 
mux6 mux_3072 (.in({n10333_0, n10332_0, n10321_0/**/, n10320_1, n10267_0, n10266_2}), .out(n6507), .config_in(config_chain[9218:9216]), .config_rst(config_rst)); 
mux6 mux_3073 (.in({n14179_1, n14178_0, n14141_0, n14140_0, n14109_0/**/, n14108_0}), .out(n6508), .config_in(config_chain[9221:9219]), .config_rst(config_rst)); 
mux6 mux_3074 (.in({n10125_0/**/, n10124_0, n10057_0, n10056_1, n10001_0, n10000_2}), .out(n6509), .config_in(config_chain[9224:9222]), .config_rst(config_rst)); 
mux6 mux_3075 (.in({n13929_1, n13928_0, n13907_0, n13906_0, n13841_0/**/, n13840_0}), .out(n6510), .config_in(config_chain[9227:9225]), .config_rst(config_rst)); 
mux6 mux_3076 (.in({n10389_0, n10388_0, n10361_0, n10360_0, n10353_0/**/, n10352_0}), .out(n6511), .config_in(config_chain[9230:9228]), .config_rst(config_rst)); 
mux6 mux_3077 (.in({n14201_2, n14200_0, n14187_1, n14186_0, n14143_0/**/, n14142_0}), .out(n6512), .config_in(config_chain[9233:9231]), .config_rst(config_rst)); 
mux6 mux_3078 (.in({n10079_0, n10078_0, n10065_0, n10064_1/**/, n10005_0, n10004_2}), .out(n6513), .config_in(config_chain[9236:9234]), .config_rst(config_rst)); 
mux6 mux_3079 (.in({n13909_0, n13908_0, n13883_0, n13882_0, n13851_0/**/, n13850_0}), .out(n6514), .config_in(config_chain[9239:9237]), .config_rst(config_rst)); 
mux6 mux_3080 (.in({n10383_0, n10382_0, n10375_0, n10374_0/**/, n10259_0, n10258_2}), .out(n6515), .config_in(config_chain[9242:9240]), .config_rst(config_rst)); 
mux6 mux_3081 (.in({n14195_1, n14194_0, n14171_0, n14170_0, n14115_0, n14114_0}), .out(n6516), .config_in(config_chain[9245:9243]), .config_rst(config_rst)); 
mux6 mux_3082 (.in({n10099_0, n10098_0, n10087_0, n10086_0/**/, n10007_0, n10006_2}), .out(n6517), .config_in(config_chain[9248:9246]), .config_rst(config_rst)); 
mux6 mux_3083 (.in({n13911_1, n13910_0, n13885_0, n13884_0, n13853_0, n13852_0/**/}), .out(n6518), .config_in(config_chain[9251:9249]), .config_rst(config_rst)); 
mux6 mux_3084 (.in({n10335_0/**/, n10334_0, n10323_0, n10322_1, n10261_0, n10260_2}), .out(n6519), .config_in(config_chain[9254:9252]), .config_rst(config_rst)); 
mux6 mux_3085 (.in({n14175_0, n14174_0, n14147_0, n14146_0, n14117_0/**/, n14116_0}), .out(n6520), .config_in(config_chain[9257:9255]), .config_rst(config_rst)); 
mux6 mux_3086 (.in({n10127_0, n10126_0/**/, n10119_0, n10118_0, n10009_0, n10008_2}), .out(n6521), .config_in(config_chain[9260:9258]), .config_rst(config_rst)); 
mux6 mux_3087 (.in({n13931_1, n13930_0, n13913_1, n13912_0, n13849_0, n13848_0}), .out(n6522), .config_in(config_chain[9263:9261]), .config_rst(config_rst)); 
mux6 mux_3088 (.in({n10643_0/**/, n10642_0, n10587_0, n10586_0, n10573_0, n10572_1}), .out(n6569), .config_in(config_chain[9266:9264]), .config_rst(config_rst)); 
mux6 mux_3089 (.in({n14217_1, n14216_0, n14117_0, n14116_0, n14095_0, n14094_0}), .out(n6570), .config_in(config_chain[9269:9267]), .config_rst(config_rst)); 
mux6 mux_3090 (.in({n10369_0, n10368_0, n10363_0, n10362_0, n10355_0, n10354_0}), .out(n6571), .config_in(config_chain[9272:9270]), .config_rst(config_rst)); 
mux6 mux_3091 (.in({n13945_1, n13944_0, n13937_1, n13936_0, n13931_0, n13930_0}), .out(n6572), .config_in(config_chain[9275:9273]), .config_rst(config_rst)); 
mux6 mux_3092 (.in({n10607_0, n10606_0, n10595_0, n10594_0, n10581_0, n10580_1}), .out(n6573), .config_in(config_chain[9278:9276]), .config_rst(config_rst)); 
mux6 mux_3093 (.in({n14181_0, n14180_0/**/, n14159_0, n14158_0, n14127_0, n14126_0}), .out(n6574), .config_in(config_chain[9281:9279]), .config_rst(config_rst)); 
mux6 mux_3094 (.in({n10385_0, n10384_0, n10317_0, n10316_1, n10309_0, n10308_1}), .out(n6575), .config_in(config_chain[9284:9282]), .config_rst(config_rst)); 
mux6 mux_3095 (.in({n13953_1, n13952_0, n13859_0, n13858_0, n13829_0, n13828_0}), .out(n6576), .config_in(config_chain[9287:9285]), .config_rst(config_rst)); 
mux6 mux_3096 (.in({n10629_0, n10628_0/**/, n10623_0, n10622_0, n10615_0, n10614_0}), .out(n6577), .config_in(config_chain[9290:9288]), .config_rst(config_rst)); 
mux6 mux_3097 (.in({n14203_1, n14202_0, n14197_0, n14196_0, n14189_0, n14188_0}), .out(n6578), .config_in(config_chain[9293:9291]), .config_rst(config_rst)); 
mux6 mux_3098 (.in({n10337_0, n10336_0, n10329_0, n10328_0, n10325_0, n10324_1}), .out(n6579), .config_in(config_chain[9296:9294]), .config_rst(config_rst)); 
mux6 mux_3099 (.in({n13917_0, n13916_0, n13891_0, n13890_0/**/, n13861_0, n13860_0}), .out(n6580), .config_in(config_chain[9299:9297]), .config_rst(config_rst)); 
mux6 mux_3100 (.in({n10645_0/**/, n10644_0, n10637_0, n10636_0, n10567_0, n10566_1}), .out(n6581), .config_in(config_chain[9302:9300]), .config_rst(config_rst)); 
mux6 mux_3101 (.in({n14219_1, n14218_0, n14125_0, n14124_0, n14093_0, n14092_0}), .out(n6582), .config_in(config_chain[9305:9303]), .config_rst(config_rst)); 
mux6 mux_3102 (.in({n10371_0, n10370_0, n10357_0, n10356_0, n10345_0, n10344_0}), .out(n6583), .config_in(config_chain[9308:9306]), .config_rst(config_rst)); 
mux6 mux_3103 (.in({n13939_1, n13938_0, n13933_0, n13932_0, n13925_0/**/, n13924_0}), .out(n6584), .config_in(config_chain[9311:9309]), .config_rst(config_rst)); 
mux6 mux_3104 (.in({n10597_0, n10596_0, n10589_0/**/, n10588_0, n10583_0, n10582_1}), .out(n6585), .config_in(config_chain[9314:9312]), .config_rst(config_rst)); 
mux6 mux_3105 (.in({n14183_0, n14182_0, n14157_0, n14156_0, n14135_0, n14134_0/**/}), .out(n6586), .config_in(config_chain[9317:9315]), .config_rst(config_rst)); 
mux6 mux_3106 (.in({n10379_0, n10378_0/**/, n10365_0, n10364_0, n10311_0, n10310_1}), .out(n6587), .config_in(config_chain[9320:9318]), .config_rst(config_rst)); 
mux6 mux_3107 (.in({n13955_1, n13954_0, n13947_1/**/, n13946_0, n13835_0, n13834_0}), .out(n6588), .config_in(config_chain[9323:9321]), .config_rst(config_rst)); 
mux6 mux_3108 (.in({n10617_0, n10616_0, n10609_0, n10608_0, n10605_0, n10604_0/**/}), .out(n6589), .config_in(config_chain[9326:9324]), .config_rst(config_rst)); 
mux6 mux_3109 (.in({n14205_1, n14204_0, n14191_0, n14190_0/**/, n14167_0, n14166_0}), .out(n6590), .config_in(config_chain[9329:9327]), .config_rst(config_rst)); 
mux6 mux_3110 (.in({n10331_0, n10330_0/**/, n10327_0, n10326_1, n10319_0, n10318_1}), .out(n6591), .config_in(config_chain[9332:9330]), .config_rst(config_rst)); 
mux6 mux_3111 (.in({n13899_0, n13898_0/**/, n13869_0, n13868_0, n13837_0, n13836_0}), .out(n6592), .config_in(config_chain[9335:9333]), .config_rst(config_rst)); 
mux6 mux_3112 (.in({n10639_0, n10638_0, n10625_0, n10624_0, n10569_0/**/, n10568_1}), .out(n6593), .config_in(config_chain[9338:9336]), .config_rst(config_rst)); 
mux6 mux_3113 (.in({n14221_1, n14220_0, n14213_1, n14212_0/**/, n14101_0, n14100_0}), .out(n6594), .config_in(config_chain[9341:9339]), .config_rst(config_rst)); 
mux6 mux_3114 (.in({n10359_0/**/, n10358_0, n10351_0, n10350_0, n10347_0, n10346_0}), .out(n6595), .config_in(config_chain[9344:9342]), .config_rst(config_rst)); 
mux6 mux_3115 (.in({n13927_0, n13926_0, n13919_0, n13918_0, n13901_0, n13900_0}), .out(n6596), .config_in(config_chain[9347:9345]), .config_rst(config_rst)); 
mux6 mux_3116 (.in({n10647_0, n10646_0, n10591_0/**/, n10590_0, n10577_0, n10576_1}), .out(n6597), .config_in(config_chain[9350:9348]), .config_rst(config_rst)); 
mux6 mux_3117 (.in({n14165_0, n14164_0, n14133_0, n14132_0, n14111_0, n14110_0}), .out(n6598), .config_in(config_chain[9353:9351]), .config_rst(config_rst)); 
mux6 mux_3118 (.in({n10381_0, n10380_0, n10373_0, n10372_0/**/, n10367_0, n10366_0}), .out(n6599), .config_in(config_chain[9356:9354]), .config_rst(config_rst)); 
mux6 mux_3119 (.in({n13949_1, n13948_0, n13935_0, n13934_0/**/, n13843_0, n13842_0}), .out(n6600), .config_in(config_chain[9359:9357]), .config_rst(config_rst)); 
mux6 mux_3120 (.in({n10611_0, n10610_0/**/, n10599_0, n10598_0, n10521_0, n10520_2}), .out(n6601), .config_in(config_chain[9362:9360]), .config_rst(config_rst)); 
mux6 mux_3121 (.in({n14193_0, n14192_0, n14185_0, n14184_0, n14175_0, n14174_0/**/}), .out(n6602), .config_in(config_chain[9365:9363]), .config_rst(config_rst)); 
mux6 mux_3122 (.in({n10333_0/**/, n10332_0, n10321_0, n10320_1, n10265_0, n10264_2}), .out(n6603), .config_in(config_chain[9368:9366]), .config_rst(config_rst)); 
mux6 mux_3123 (.in({n13913_1, n13912_0, n13875_0/**/, n13874_0, n13845_0, n13844_0}), .out(n6604), .config_in(config_chain[9371:9369]), .config_rst(config_rst)); 
mux6 mux_3124 (.in({n10633_0, n10632_0, n10619_0/**/, n10618_0, n10523_0, n10522_2}), .out(n6605), .config_in(config_chain[9374:9372]), .config_rst(config_rst)); 
mux6 mux_3125 (.in({n14215_1, n14214_0, n14207_1, n14206_0/**/, n14177_0, n14176_0}), .out(n6606), .config_in(config_chain[9377:9375]), .config_rst(config_rst)); 
mux6 mux_3126 (.in({n10353_0, n10352_0, n10341_0, n10340_0, n10267_0/**/, n10266_2}), .out(n6607), .config_in(config_chain[9380:9378]), .config_rst(config_rst)); 
mux6 mux_3127 (.in({n13957_2, n13956_0, n13921_0, n13920_0, n13877_0, n13876_0}), .out(n6608), .config_in(config_chain[9383:9381]), .config_rst(config_rst)); 
mux6 mux_3128 (.in({n10579_0, n10578_1, n10571_0, n10570_1/**/, n10525_0, n10524_2}), .out(n6609), .config_in(config_chain[9386:9384]), .config_rst(config_rst)); 
mux6 mux_3129 (.in({n14179_1, n14178_0, n14141_0, n14140_0/**/, n14119_0, n14118_0}), .out(n6610), .config_in(config_chain[9389:9387]), .config_rst(config_rst)); 
mux6 mux_3130 (.in({n10375_0, n10374_0, n10361_0, n10360_0/**/, n10259_0, n10258_2}), .out(n6611), .config_in(config_chain[9392:9390]), .config_rst(config_rst)); 
mux6 mux_3131 (.in({n13951_1, n13950_0, n13943_1/**/, n13942_0, n13907_0, n13906_0}), .out(n6612), .config_in(config_chain[9395:9393]), .config_rst(config_rst)); 
mux6 mux_3132 (.in({n10627_0, n10626_0, n10601_0, n10600_0, n10593_0/**/, n10592_0}), .out(n6613), .config_in(config_chain[9398:9396]), .config_rst(config_rst)); 
mux6 mux_3133 (.in({n14201_2, n14200_0, n14187_0/**/, n14186_0, n14151_0, n14150_0}), .out(n6614), .config_in(config_chain[9401:9399]), .config_rst(config_rst)); 
mux6 mux_3134 (.in({n10383_0, n10382_0/**/, n10315_0, n10314_1, n10261_0, n10260_2}), .out(n6615), .config_in(config_chain[9404:9402]), .config_rst(config_rst)); 
mux6 mux_3135 (.in({n13909_0, n13908_0, n13883_0, n13882_0, n13851_0, n13850_0}), .out(n6616), .config_in(config_chain[9407:9405]), .config_rst(config_rst)); 
mux6 mux_3136 (.in({n10649_0, n10648_0, n10635_0, n10634_0, n10621_0, n10620_0/**/}), .out(n6617), .config_in(config_chain[9410:9408]), .config_rst(config_rst)); 
mux6 mux_3137 (.in({n14209_1/**/, n14208_0, n14195_0, n14194_0, n14173_0, n14172_0}), .out(n6618), .config_in(config_chain[9413:9411]), .config_rst(config_rst)); 
mux6 mux_3138 (.in({n10343_0, n10342_0, n10335_0, n10334_0, n10263_0/**/, n10262_2}), .out(n6619), .config_in(config_chain[9416:9414]), .config_rst(config_rst)); 
mux6 mux_3139 (.in({n13923_0, n13922_0, n13911_0, n13910_0, n13885_0, n13884_0}), .out(n6620), .config_in(config_chain[9419:9417]), .config_rst(config_rst)); 
mux6 mux_3140 (.in({n10891_0, n10890_0, n10875_0, n10874_0, n10861_0, n10860_0}), .out(n6667), .config_in(config_chain[9422:9420]), .config_rst(config_rst)); 
mux6 mux_3141 (.in({n14225_1, n14224_0, n14209_0, n14208_0, n14195_0, n14194_0}), .out(n6668), .config_in(config_chain[9425:9423]), .config_rst(config_rst)); 
mux6 mux_3142 (.in({n10587_0, n10586_0, n10581_0, n10580_1, n10573_0, n10572_1}), .out(n6669), .config_in(config_chain[9428:9426]), .config_rst(config_rst)); 
mux6 mux_3143 (.in({n13925_0, n13924_0, n13917_0, n13916_0, n13885_0, n13884_1}), .out(n6670), .config_in(config_chain[9431:9429]), .config_rst(config_rst)); 
mux6 mux_3144 (.in({n10899_0, n10898_0, n10883_0, n10882_0, n10827_0, n10826_1}), .out(n6671), .config_in(config_chain[9434:9432]), .config_rst(config_rst)); 
mux6 mux_3145 (.in({n14241_1, n14240_0, n14233_1, n14232_0, n14095_0, n14094_1}), .out(n6672), .config_in(config_chain[9437:9435]), .config_rst(config_rst)); 
mux6 mux_3146 (.in({n10615_0, n10614_0/**/, n10607_0, n10606_0, n10603_0, n10602_0}), .out(n6673), .config_in(config_chain[9440:9438]), .config_rst(config_rst)); 
mux6 mux_3147 (.in({n13959_1, n13958_0, n13945_0/**/, n13944_0, n13933_0, n13932_0}), .out(n6674), .config_in(config_chain[9443:9441]), .config_rst(config_rst)); 
mux6 mux_3148 (.in({n10847_0, n10846_0, n10843_0, n10842_1, n10835_0, n10834_1}), .out(n6675), .config_in(config_chain[9446:9444]), .config_rst(config_rst)); 
mux6 mux_3149 (.in({n14181_0, n14180_0, n14159_0, n14158_1, n14127_0/**/, n14126_1}), .out(n6676), .config_in(config_chain[9449:9447]), .config_rst(config_rst)); 
mux6 mux_3150 (.in({n10637_0, n10636_0, n10629_0, n10628_0, n10623_0, n10622_0}), .out(n6677), .config_in(config_chain[9452:9450]), .config_rst(config_rst)); 
mux6 mux_3151 (.in({n13967_1, n13966_0, n13953_0, n13952_0, n13829_0, n13828_1/**/}), .out(n6678), .config_in(config_chain[9455:9453]), .config_rst(config_rst)); 
mux6 mux_3152 (.in({n10869_0, n10868_0, n10863_0, n10862_0, n10855_0/**/, n10854_0}), .out(n6679), .config_in(config_chain[9458:9456]), .config_rst(config_rst)); 
mux6 mux_3153 (.in({n14211_0, n14210_0, n14203_0, n14202_0, n14197_0, n14196_0/**/}), .out(n6680), .config_in(config_chain[9461:9459]), .config_rst(config_rst)); 
mux6 mux_3154 (.in({n10645_0, n10644_0, n10589_0, n10588_0, n10575_0, n10574_1/**/}), .out(n6681), .config_in(config_chain[9464:9462]), .config_rst(config_rst)); 
mux6 mux_3155 (.in({n13919_0/**/, n13918_0, n13893_0, n13892_1, n13861_0, n13860_1}), .out(n6682), .config_in(config_chain[9467:9465]), .config_rst(config_rst)); 
mux6 mux_3156 (.in({n10901_0/**/, n10900_0, n10893_0, n10892_0, n10885_0, n10884_0}), .out(n6683), .config_in(config_chain[9470:9468]), .config_rst(config_rst)); 
mux6 mux_3157 (.in({n14235_1/**/, n14234_0, n14219_0, n14218_0, n14103_0, n14102_1}), .out(n6684), .config_in(config_chain[9473:9471]), .config_rst(config_rst)); 
mux6 mux_3158 (.in({n10609_0, n10608_0, n10597_0/**/, n10596_0, n10583_0, n10582_1}), .out(n6685), .config_in(config_chain[9476:9474]), .config_rst(config_rst)); 
mux6 mux_3159 (.in({n13939_0, n13938_0, n13935_0, n13934_0/**/, n13927_0, n13926_0}), .out(n6686), .config_in(config_chain[9479:9477]), .config_rst(config_rst)); 
mux6 mux_3160 (.in({n10909_0, n10908_0, n10837_0, n10836_1, n10829_0, n10828_1}), .out(n6687), .config_in(config_chain[9482:9480]), .config_rst(config_rst)); 
mux6 mux_3161 (.in({n14243_1, n14242_0/**/, n14183_0, n14182_0, n14135_0, n14134_1}), .out(n6688), .config_in(config_chain[9485:9483]), .config_rst(config_rst)); 
mux6 mux_3162 (.in({n10631_0, n10630_0, n10625_0, n10624_0, n10617_0, n10616_0/**/}), .out(n6689), .config_in(config_chain[9488:9486]), .config_rst(config_rst)); 
mux6 mux_3163 (.in({n13969_1/**/, n13968_0, n13961_1, n13960_0, n13955_0, n13954_0}), .out(n6690), .config_in(config_chain[9491:9489]), .config_rst(config_rst)); 
mux6 mux_3164 (.in({n10871_0, n10870_0, n10857_0/**/, n10856_0, n10845_0, n10844_1}), .out(n6691), .config_in(config_chain[9494:9492]), .config_rst(config_rst)); 
mux6 mux_3165 (.in({n14205_0, n14204_0, n14199_0, n14198_0, n14191_0, n14190_0}), .out(n6692), .config_in(config_chain[9497:9495]), .config_rst(config_rst)); 
mux6 mux_3166 (.in({n10647_0, n10646_0/**/, n10577_0, n10576_1, n10569_0, n10568_1}), .out(n6693), .config_in(config_chain[9500:9498]), .config_rst(config_rst)); 
mux6 mux_3167 (.in({n13977_1, n13976_0, n13869_0, n13868_1/**/, n13837_0, n13836_1}), .out(n6694), .config_in(config_chain[9503:9501]), .config_rst(config_rst)); 
mux6 mux_3168 (.in({n10895_0, n10894_0, n10879_0, n10878_0, n10865_0, n10864_0/**/}), .out(n6695), .config_in(config_chain[9506:9504]), .config_rst(config_rst)); 
mux6 mux_3169 (.in({n14229_1, n14228_0, n14221_0, n14220_0/**/, n14213_0, n14212_0}), .out(n6696), .config_in(config_chain[9509:9507]), .config_rst(config_rst)); 
mux6 mux_3170 (.in({n10599_0, n10598_0/**/, n10591_0, n10590_0, n10585_0, n10584_1}), .out(n6697), .config_in(config_chain[9512:9510]), .config_rst(config_rst)); 
mux6 mux_3171 (.in({n13941_0, n13940_0, n13929_0, n13928_0/**/, n13901_0, n13900_1}), .out(n6698), .config_in(config_chain[9515:9513]), .config_rst(config_rst)); 
mux6 mux_3172 (.in({n10911_0, n10910_0, n10903_0, n10902_0, n10831_0, n10830_1/**/}), .out(n6699), .config_in(config_chain[9518:9516]), .config_rst(config_rst)); 
mux6 mux_3173 (.in({n14245_1, n14244_0, n14143_0, n14142_1/**/, n14111_0, n14110_1}), .out(n6700), .config_in(config_chain[9521:9519]), .config_rst(config_rst)); 
mux6 mux_3174 (.in({n10633_0/**/, n10632_0, n10619_0, n10618_0, n10521_0, n10520_2}), .out(n6701), .config_in(config_chain[9524:9522]), .config_rst(config_rst)); 
mux6 mux_3175 (.in({n13963_1, n13962_0, n13949_0, n13948_0, n13911_0, n13910_1}), .out(n6702), .config_in(config_chain[9527:9525]), .config_rst(config_rst)); 
mux6 mux_3176 (.in({n10851_0, n10850_0, n10839_0, n10838_1/**/, n10781_0, n10780_2}), .out(n6703), .config_in(config_chain[9530:9528]), .config_rst(config_rst)); 
mux6 mux_3177 (.in({n14193_0, n14192_0/**/, n14185_0, n14184_0, n14175_0, n14174_1}), .out(n6704), .config_in(config_chain[9533:9531]), .config_rst(config_rst)); 
mux6 mux_3178 (.in({n10641_0, n10640_0, n10571_0/**/, n10570_1, n10523_0, n10522_2}), .out(n6705), .config_in(config_chain[9536:9534]), .config_rst(config_rst)); 
mux6 mux_3179 (.in({n13971_1, n13970_0, n13915_1, n13914_1, n13845_0, n13844_1}), .out(n6706), .config_in(config_chain[9539:9537]), .config_rst(config_rst)); 
mux6 mux_3180 (.in({n10881_0, n10880_0, n10873_0, n10872_0, n10783_0/**/, n10782_2}), .out(n6707), .config_in(config_chain[9542:9540]), .config_rst(config_rst)); 
mux6 mux_3181 (.in({n14231_1, n14230_0/**/, n14215_0, n14214_0, n14177_0, n14176_1}), .out(n6708), .config_in(config_chain[9545:9543]), .config_rst(config_rst)); 
mux6 mux_3182 (.in({n10627_0, n10626_0, n10593_0, n10592_0, n10579_0, n10578_1}), .out(n6709), .config_in(config_chain[9548:9546]), .config_rst(config_rst)); 
mux6 mux_3183 (.in({n13957_1, n13956_0, n13931_0, n13930_0, n13923_0/**/, n13922_0}), .out(n6710), .config_in(config_chain[9551:9549]), .config_rst(config_rst)); 
mux6 mux_3184 (.in({n10905_0, n10904_0/**/, n10897_0, n10896_0, n10785_0, n10784_2}), .out(n6711), .config_in(config_chain[9554:9552]), .config_rst(config_rst)); 
mux6 mux_3185 (.in({n14239_1/**/, n14238_0, n14179_0, n14178_1, n14119_0, n14118_1}), .out(n6712), .config_in(config_chain[9557:9555]), .config_rst(config_rst)); 
mux6 mux_3186 (.in({n10649_0, n10648_0, n10613_0, n10612_0/**/, n10601_0, n10600_0}), .out(n6713), .config_in(config_chain[9560:9558]), .config_rst(config_rst)); 
mux6 mux_3187 (.in({n13979_1, n13978_0, n13951_0/**/, n13950_0, n13943_0, n13942_0}), .out(n6714), .config_in(config_chain[9563:9561]), .config_rst(config_rst)); 
mux6 mux_3188 (.in({n10867_0, n10866_0, n10853_0, n10852_0, n10841_0, n10840_1}), .out(n6715), .config_in(config_chain[9566:9564]), .config_rst(config_rst)); 
mux6 mux_3189 (.in({n14223_1, n14222_0, n14187_0, n14186_0, n14151_0, n14150_1}), .out(n6716), .config_in(config_chain[9569:9567]), .config_rst(config_rst)); 
mux6 mux_3190 (.in({n10643_0, n10642_0/**/, n10635_0, n10634_0, n10519_0, n10518_2}), .out(n6717), .config_in(config_chain[9572:9570]), .config_rst(config_rst)); 
mux6 mux_3191 (.in({n13973_1, n13972_0/**/, n13909_0, n13908_1, n13853_0, n13852_1}), .out(n6718), .config_in(config_chain[9575:9573]), .config_rst(config_rst)); 
mux6 mux_3192 (.in({n11169_0, n11168_0, n11111_0, n11110_0, n11095_0, n11094_1}), .out(n6765), .config_in(config_chain[9578:9576]), .config_rst(config_rst)); 
mux6 mux_3193 (.in({n14261_1, n14260_0, n14203_0, n14202_0, n14187_0, n14186_1}), .out(n6766), .config_in(config_chain[9581:9579]), .config_rst(config_rst)); 
mux6 mux_3194 (.in({n10891_0, n10890_0, n10883_0, n10882_0, n10875_0, n10874_0}), .out(n6767), .config_in(config_chain[9584:9582]), .config_rst(config_rst)); 
mux6 mux_3195 (.in({n13989_1, n13988_0, n13981_1, n13980_0, n13973_0, n13972_0}), .out(n6768), .config_in(config_chain[9587:9585]), .config_rst(config_rst)); 
mux6 mux_3196 (.in({n11133_0, n11132_0, n11119_0, n11118_0, n11103_0, n11102_1}), .out(n6769), .config_in(config_chain[9590:9588]), .config_rst(config_rst)); 
mux6 mux_3197 (.in({n14225_0, n14224_0, n14219_0, n14218_0, n14211_0, n14210_0}), .out(n6770), .config_in(config_chain[9593:9591]), .config_rst(config_rst)); 
mux6 mux_3198 (.in({n10907_0, n10906_0, n10835_0, n10834_1, n10827_0, n10826_1}), .out(n6771), .config_in(config_chain[9596:9594]), .config_rst(config_rst)); 
mux6 mux_3199 (.in({n13997_1, n13996_0, n13937_0, n13936_0, n13925_0, n13924_1}), .out(n6772), .config_in(config_chain[9599:9597]), .config_rst(config_rst)); 
mux6 mux_3200 (.in({n11155_0, n11154_0, n11149_0, n11148_0, n11141_0, n11140_0}), .out(n6773), .config_in(config_chain[9602:9600]), .config_rst(config_rst)); 
mux6 mux_3201 (.in({n14247_1, n14246_0, n14241_0, n14240_0, n14233_0, n14232_0}), .out(n6774), .config_in(config_chain[9605:9603]), .config_rst(config_rst)); 
mux6 mux_3202 (.in({n10855_0, n10854_0, n10847_0, n10846_0, n10843_0, n10842_1}), .out(n6775), .config_in(config_chain[9608:9606]), .config_rst(config_rst)); 
mux6 mux_3203 (.in({n13959_0, n13958_0, n13945_0, n13944_0, n13933_0, n13932_1}), .out(n6776), .config_in(config_chain[9611:9609]), .config_rst(config_rst)); 
mux6 mux_3204 (.in({n11171_0, n11170_0, n11163_0, n11162_0, n11089_0, n11088_1/**/}), .out(n6777), .config_in(config_chain[9614:9612]), .config_rst(config_rst)); 
mux6 mux_3205 (.in({n14263_1/**/, n14262_0, n14189_0, n14188_1, n14181_0, n14180_1}), .out(n6778), .config_in(config_chain[9617:9615]), .config_rst(config_rst)); 
mux6 mux_3206 (.in({n10893_0, n10892_0/**/, n10877_0, n10876_0, n10863_0, n10862_0}), .out(n6779), .config_in(config_chain[9620:9618]), .config_rst(config_rst)); 
mux6 mux_3207 (.in({n13983_1, n13982_0, n13975_0, n13974_0, n13967_0/**/, n13966_0}), .out(n6780), .config_in(config_chain[9623:9621]), .config_rst(config_rst)); 
mux6 mux_3208 (.in({n11121_0, n11120_0, n11113_0, n11112_0, n11105_0, n11104_1/**/}), .out(n6781), .config_in(config_chain[9626:9624]), .config_rst(config_rst)); 
mux6 mux_3209 (.in({n14227_0, n14226_0, n14213_0, n14212_0, n14197_0, n14196_1}), .out(n6782), .config_in(config_chain[9629:9627]), .config_rst(config_rst)); 
mux6 mux_3210 (.in({n10901_0, n10900_0, n10885_0, n10884_0, n10829_0, n10828_1}), .out(n6783), .config_in(config_chain[9632:9630]), .config_rst(config_rst)); 
mux6 mux_3211 (.in({n13999_1, n13998_0, n13991_1, n13990_0, n13919_0, n13918_1}), .out(n6784), .config_in(config_chain[9635:9633]), .config_rst(config_rst)); 
mux6 mux_3212 (.in({n11143_0, n11142_0, n11135_0, n11134_0, n11129_0, n11128_0}), .out(n6785), .config_in(config_chain[9638:9636]), .config_rst(config_rst)); 
mux6 mux_3213 (.in({n14249_1, n14248_0, n14235_0, n14234_0, n14221_0, n14220_0}), .out(n6786), .config_in(config_chain[9641:9639]), .config_rst(config_rst)); 
mux6 mux_3214 (.in({n10849_0, n10848_0, n10845_0, n10844_1/**/, n10837_0, n10836_1}), .out(n6787), .config_in(config_chain[9644:9642]), .config_rst(config_rst)); 
mux6 mux_3215 (.in({n13947_0, n13946_0/**/, n13939_0, n13938_0, n13935_0, n13934_1}), .out(n6788), .config_in(config_chain[9647:9645]), .config_rst(config_rst)); 
mux6 mux_3216 (.in({n11165_0, n11164_0, n11151_0, n11150_0/**/, n11091_0, n11090_1}), .out(n6789), .config_in(config_chain[9650:9648]), .config_rst(config_rst)); 
mux6 mux_3217 (.in({n14265_1, n14264_0, n14257_1/**/, n14256_0, n14183_0, n14182_1}), .out(n6790), .config_in(config_chain[9653:9651]), .config_rst(config_rst)); 
mux6 mux_3218 (.in({n10879_0, n10878_0, n10871_0, n10870_0, n10865_0, n10864_0}), .out(n6791), .config_in(config_chain[9656:9654]), .config_rst(config_rst)); 
mux6 mux_3219 (.in({n13969_0, n13968_0, n13961_0, n13960_0, n13955_0/**/, n13954_0}), .out(n6792), .config_in(config_chain[9659:9657]), .config_rst(config_rst)); 
mux6 mux_3220 (.in({n11173_0/**/, n11172_0, n11115_0, n11114_0, n11099_0, n11098_1}), .out(n6793), .config_in(config_chain[9662:9660]), .config_rst(config_rst)); 
mux6 mux_3221 (.in({n14207_0, n14206_0, n14199_0, n14198_1/**/, n14191_0, n14190_1}), .out(n6794), .config_in(config_chain[9665:9663]), .config_rst(config_rst)); 
mux6 mux_3222 (.in({n10903_0, n10902_0, n10895_0, n10894_0/**/, n10887_0, n10886_0}), .out(n6795), .config_in(config_chain[9668:9666]), .config_rst(config_rst)); 
mux6 mux_3223 (.in({n13993_1, n13992_0, n13977_0, n13976_0, n13921_0, n13920_1/**/}), .out(n6796), .config_in(config_chain[9671:9669]), .config_rst(config_rst)); 
mux6 mux_3224 (.in({n11137_0, n11136_0, n11131_0, n11130_0, n11123_0, n11122_0}), .out(n6797), .config_in(config_chain[9674:9672]), .config_rst(config_rst)); 
mux6 mux_3225 (.in({n14237_0, n14236_0, n14229_0, n14228_0, n14223_1, n14222_0}), .out(n6798), .config_in(config_chain[9677:9675]), .config_rst(config_rst)); 
mux6 mux_3226 (.in({n10911_0, n10910_0, n10851_0, n10850_0, n10839_0, n10838_1/**/}), .out(n6799), .config_in(config_chain[9680:9678]), .config_rst(config_rst)); 
mux6 mux_3227 (.in({n14001_1, n14000_0, n13941_0/**/, n13940_0, n13929_0, n13928_1}), .out(n6800), .config_in(config_chain[9683:9681]), .config_rst(config_rst)); 
mux6 mux_3228 (.in({n11159_0, n11158_0, n11153_0, n11152_0, n11145_0, n11144_0}), .out(n6801), .config_in(config_chain[9686:9684]), .config_rst(config_rst)); 
mux6 mux_3229 (.in({n14259_1, n14258_0, n14251_1, n14250_0, n14245_1, n14244_0}), .out(n6802), .config_in(config_chain[9689:9687]), .config_rst(config_rst)); 
mux6 mux_3230 (.in({n10873_0, n10872_0/**/, n10859_0, n10858_0, n10781_0, n10780_2}), .out(n6803), .config_in(config_chain[9692:9690]), .config_rst(config_rst)); 
mux6 mux_3231 (.in({n13963_0, n13962_0, n13949_0, n13948_0, n13913_0/**/, n13912_1}), .out(n6804), .config_in(config_chain[9695:9693]), .config_rst(config_rst)); 
mux6 mux_3232 (.in({n11175_0, n11174_0, n11101_0, n11100_1, n11093_0, n11092_1/**/}), .out(n6805), .config_in(config_chain[9698:9696]), .config_rst(config_rst)); 
mux6 mux_3233 (.in({n14267_1, n14266_0, n14209_0, n14208_0, n14193_0, n14192_1}), .out(n6806), .config_in(config_chain[9701:9699]), .config_rst(config_rst)); 
mux6 mux_3234 (.in({n10897_0/**/, n10896_0, n10881_0, n10880_0, n10785_0, n10784_2}), .out(n6807), .config_in(config_chain[9704:9702]), .config_rst(config_rst)); 
mux6 mux_3235 (.in({n13995_1, n13994_0, n13987_1, n13986_0, n13915_0, n13914_1}), .out(n6808), .config_in(config_chain[9707:9705]), .config_rst(config_rst)); 
mux6 mux_3236 (.in({n11125_0, n11124_0, n11117_0, n11116_0, n11045_0, n11044_2}), .out(n6809), .config_in(config_chain[9710:9708]), .config_rst(config_rst)); 
mux6 mux_3237 (.in({n14231_0, n14230_0, n14217_0, n14216_0/**/, n14177_0, n14176_1}), .out(n6810), .config_in(config_chain[9713:9711]), .config_rst(config_rst)); 
mux6 mux_3238 (.in({n10905_0, n10904_0, n10867_0, n10866_0, n10833_0/**/, n10832_1}), .out(n6811), .config_in(config_chain[9716:9714]), .config_rst(config_rst)); 
mux6 mux_3239 (.in({n13957_1, n13956_0, n13931_0, n13930_1, n13923_0, n13922_1}), .out(n6812), .config_in(config_chain[9719:9717]), .config_rst(config_rst)); 
mux6 mux_3240 (.in({n11161_0/**/, n11160_0, n11147_0, n11146_0, n11047_0, n11046_2}), .out(n6813), .config_in(config_chain[9722:9720]), .config_rst(config_rst)); 
mux6 mux_3241 (.in({n14253_1, n14252_0, n14239_0, n14238_0, n14201_1, n14200_1}), .out(n6814), .config_in(config_chain[9725:9723]), .config_rst(config_rst)); 
mux6 mux_3242 (.in({n10889_0, n10888_0, n10861_0, n10860_0, n10853_0, n10852_0}), .out(n6815), .config_in(config_chain[9728:9726]), .config_rst(config_rst)); 
mux6 mux_3243 (.in({n13979_1, n13978_0, n13965_0, n13964_0, n13951_0, n13950_0/**/}), .out(n6816), .config_in(config_chain[9731:9729]), .config_rst(config_rst)); 
mux6 mux_3244 (.in({n11421_0, n11420_0, n11405_0, n11404_0, n11391_0, n11390_0}), .out(n6863), .config_in(config_chain[9734:9732]), .config_rst(config_rst)); 
mux6 mux_3245 (.in({n14269_1, n14268_0, n14253_0, n14252_0, n14239_0, n14238_0}), .out(n6864), .config_in(config_chain[9737:9735]), .config_rst(config_rst)); 
mux6 mux_3246 (.in({n11111_0, n11110_0, n11103_0, n11102_1, n11095_0, n11094_1}), .out(n6865), .config_in(config_chain[9740:9738]), .config_rst(config_rst)); 
mux6 mux_3247 (.in({n13967_0, n13966_0, n13959_0, n13958_0, n13951_0/**/, n13950_1}), .out(n6866), .config_in(config_chain[9743:9741]), .config_rst(config_rst)); 
mux6 mux_3248 (.in({n11429_0, n11428_0, n11413_0/**/, n11412_0, n11355_0, n11354_1}), .out(n6867), .config_in(config_chain[9746:9744]), .config_rst(config_rst)); 
mux6 mux_3249 (.in({n14285_1, n14284_0, n14277_1, n14276_0, n14203_0, n14202_1}), .out(n6868), .config_in(config_chain[9749:9747]), .config_rst(config_rst)); 
mux6 mux_3250 (.in({n11141_0, n11140_0, n11133_0, n11132_0, n11127_0, n11126_0}), .out(n6869), .config_in(config_chain[9752:9750]), .config_rst(config_rst)); 
mux6 mux_3251 (.in({n14003_1, n14002_0, n13989_0, n13988_0/**/, n13975_0, n13974_0}), .out(n6870), .config_in(config_chain[9755:9753]), .config_rst(config_rst)); 
mux6 mux_3252 (.in({n11377_0, n11376_0, n11371_0, n11370_1, n11363_0, n11362_1}), .out(n6871), .config_in(config_chain[9758:9756]), .config_rst(config_rst)); 
mux6 mux_3253 (.in({n14225_0, n14224_0, n14219_0, n14218_1, n14211_0, n14210_1}), .out(n6872), .config_in(config_chain[9761:9759]), .config_rst(config_rst)); 
mux6 mux_3254 (.in({n11163_0, n11162_0, n11155_0, n11154_0, n11149_0/**/, n11148_0}), .out(n6873), .config_in(config_chain[9764:9762]), .config_rst(config_rst)); 
mux6 mux_3255 (.in({n14011_1, n14010_0, n13997_0, n13996_0, n13937_0, n13936_1}), .out(n6874), .config_in(config_chain[9767:9765]), .config_rst(config_rst)); 
mux6 mux_3256 (.in({n11399_0, n11398_0, n11393_0, n11392_0, n11385_0/**/, n11384_0}), .out(n6875), .config_in(config_chain[9770:9768]), .config_rst(config_rst)); 
mux6 mux_3257 (.in({n14255_0, n14254_0, n14247_0/**/, n14246_0, n14241_0, n14240_0}), .out(n6876), .config_in(config_chain[9773:9771]), .config_rst(config_rst)); 
mux6 mux_3258 (.in({n11171_0, n11170_0, n11113_0, n11112_0/**/, n11097_0, n11096_1}), .out(n6877), .config_in(config_chain[9776:9774]), .config_rst(config_rst)); 
mux6 mux_3259 (.in({n13961_0/**/, n13960_0, n13953_0, n13952_1, n13945_0, n13944_1}), .out(n6878), .config_in(config_chain[9779:9777]), .config_rst(config_rst)); 
mux6 mux_3260 (.in({n11431_0, n11430_0, n11423_0/**/, n11422_0, n11415_0, n11414_0}), .out(n6879), .config_in(config_chain[9782:9780]), .config_rst(config_rst)); 
mux6 mux_3261 (.in({n14279_1, n14278_0, n14263_0, n14262_0, n14205_0, n14204_1/**/}), .out(n6880), .config_in(config_chain[9785:9783]), .config_rst(config_rst)); 
mux6 mux_3262 (.in({n11135_0, n11134_0, n11121_0, n11120_0/**/, n11105_0, n11104_1}), .out(n6881), .config_in(config_chain[9788:9786]), .config_rst(config_rst)); 
mux6 mux_3263 (.in({n13983_0, n13982_0, n13977_0, n13976_0, n13969_0/**/, n13968_0}), .out(n6882), .config_in(config_chain[9791:9789]), .config_rst(config_rst)); 
mux6 mux_3264 (.in({n11439_0, n11438_0, n11365_0, n11364_1, n11357_0/**/, n11356_1}), .out(n6883), .config_in(config_chain[9794:9792]), .config_rst(config_rst)); 
mux6 mux_3265 (.in({n14287_1/**/, n14286_0, n14227_0, n14226_0, n14213_0, n14212_1}), .out(n6884), .config_in(config_chain[9797:9795]), .config_rst(config_rst)); 
mux6 mux_3266 (.in({n11157_0, n11156_0, n11151_0, n11150_0, n11143_0, n11142_0/**/}), .out(n6885), .config_in(config_chain[9800:9798]), .config_rst(config_rst)); 
mux6 mux_3267 (.in({n14013_1, n14012_0, n14005_1, n14004_0/**/, n13999_0, n13998_0}), .out(n6886), .config_in(config_chain[9803:9801]), .config_rst(config_rst)); 
mux6 mux_3268 (.in({n11401_0, n11400_0/**/, n11387_0, n11386_0, n11373_0, n11372_1}), .out(n6887), .config_in(config_chain[9806:9804]), .config_rst(config_rst)); 
mux6 mux_3269 (.in({n14249_0, n14248_0, n14243_0, n14242_0, n14235_0, n14234_0}), .out(n6888), .config_in(config_chain[9809:9807]), .config_rst(config_rst)); 
mux6 mux_3270 (.in({n11173_0, n11172_0, n11099_0, n11098_1, n11091_0, n11090_1}), .out(n6889), .config_in(config_chain[9812:9810]), .config_rst(config_rst)); 
mux6 mux_3271 (.in({n14021_1, n14020_0, n13947_0, n13946_1, n13939_0, n13938_1}), .out(n6890), .config_in(config_chain[9815:9813]), .config_rst(config_rst)); 
mux6 mux_3272 (.in({n11425_0, n11424_0/**/, n11409_0, n11408_0, n11395_0, n11394_0}), .out(n6891), .config_in(config_chain[9818:9816]), .config_rst(config_rst)); 
mux6 mux_3273 (.in({n14273_1, n14272_0/**/, n14265_0, n14264_0, n14257_0, n14256_0}), .out(n6892), .config_in(config_chain[9821:9819]), .config_rst(config_rst)); 
mux6 mux_3274 (.in({n11123_0, n11122_0, n11115_0, n11114_0, n11107_0, n11106_1/**/}), .out(n6893), .config_in(config_chain[9824:9822]), .config_rst(config_rst)); 
mux6 mux_3275 (.in({n13985_0, n13984_0, n13971_0, n13970_0, n13955_0, n13954_1}), .out(n6894), .config_in(config_chain[9827:9825]), .config_rst(config_rst)); 
mux6 mux_3276 (.in({n11433_0, n11432_0, n11359_0, n11358_1/**/, n11353_0, n11352_1}), .out(n6895), .config_in(config_chain[9830:9828]), .config_rst(config_rst)); 
mux6 mux_3277 (.in({n14215_0/**/, n14214_1, n14207_0, n14206_1, n14201_1, n14200_1}), .out(n6896), .config_in(config_chain[9833:9831]), .config_rst(config_rst)); 
mux6 mux_3278 (.in({n11159_0, n11158_0, n11145_0/**/, n11144_0, n11131_0, n11130_0}), .out(n6897), .config_in(config_chain[9836:9834]), .config_rst(config_rst)); 
mux6 mux_3279 (.in({n14007_1, n14006_0, n13993_0, n13992_0, n13979_1, n13978_0/**/}), .out(n6898), .config_in(config_chain[9839:9837]), .config_rst(config_rst)); 
mux6 mux_3280 (.in({n11381_0, n11380_0, n11375_0, n11374_1, n11367_0, n11366_1/**/}), .out(n6899), .config_in(config_chain[9842:9840]), .config_rst(config_rst)); 
mux6 mux_3281 (.in({n14237_0, n14236_0, n14229_0, n14228_0, n14223_1, n14222_1}), .out(n6900), .config_in(config_chain[9845:9843]), .config_rst(config_rst)); 
mux6 mux_3282 (.in({n11167_0, n11166_0, n11153_0, n11152_0, n11093_0/**/, n11092_1}), .out(n6901), .config_in(config_chain[9848:9846]), .config_rst(config_rst)); 
mux6 mux_3283 (.in({n14023_1, n14022_0, n14015_1, n14014_0, n13941_0, n13940_1}), .out(n6902), .config_in(config_chain[9851:9849]), .config_rst(config_rst)); 
mux6 mux_3284 (.in({n11411_0, n11410_0/**/, n11403_0, n11402_0, n11397_0, n11396_0}), .out(n6903), .config_in(config_chain[9854:9852]), .config_rst(config_rst)); 
mux6 mux_3285 (.in({n14275_1, n14274_0, n14259_0/**/, n14258_0, n14245_1, n14244_0}), .out(n6904), .config_in(config_chain[9857:9855]), .config_rst(config_rst)); 
mux6 mux_3286 (.in({n11117_0, n11116_0/**/, n11101_0, n11100_1, n11045_0, n11044_2}), .out(n6905), .config_in(config_chain[9860:9858]), .config_rst(config_rst)); 
mux6 mux_3287 (.in({n13973_0, n13972_0, n13965_0/**/, n13964_0, n13913_0, n13912_1}), .out(n6906), .config_in(config_chain[9863:9861]), .config_rst(config_rst)); 
mux6 mux_3288 (.in({n11435_0, n11434_0, n11427_0, n11426_0, n11419_0, n11418_0/**/}), .out(n6907), .config_in(config_chain[9866:9864]), .config_rst(config_rst)); 
mux6 mux_3289 (.in({n14283_1, n14282_0, n14267_1, n14266_0, n14209_0, n14208_1}), .out(n6908), .config_in(config_chain[9869:9867]), .config_rst(config_rst)); 
mux6 mux_3290 (.in({n11139_0, n11138_0, n11125_0, n11124_0, n11047_0, n11046_2}), .out(n6909), .config_in(config_chain[9872:9870]), .config_rst(config_rst)); 
mux6 mux_3291 (.in({n13995_0, n13994_0, n13987_0, n13986_0, n13915_0/**/, n13914_1}), .out(n6910), .config_in(config_chain[9875:9873]), .config_rst(config_rst)); 
mux6 mux_3292 (.in({n11441_0, n11440_0, n11383_0, n11382_0, n11369_0, n11368_1/**/}), .out(n6911), .config_in(config_chain[9878:9876]), .config_rst(config_rst)); 
mux6 mux_3293 (.in({n14231_0, n14230_0, n14217_0, n14216_1, n14179_0, n14178_1}), .out(n6912), .config_in(config_chain[9881:9879]), .config_rst(config_rst)); 
mux6 mux_3294 (.in({n11169_0, n11168_0, n11161_0, n11160_0/**/, n11109_0, n11108_1}), .out(n6913), .config_in(config_chain[9884:9882]), .config_rst(config_rst)); 
mux6 mux_3295 (.in({n14017_1, n14016_0, n13957_1, n13956_1, n13943_0, n13942_1/**/}), .out(n6914), .config_in(config_chain[9887:9885]), .config_rst(config_rst)); 
mux6 mux_3296 (.in({n11701_0, n11700_0, n11643_0, n11642_0, n11627_0, n11626_1}), .out(n6961), .config_in(config_chain[9890:9888]), .config_rst(config_rst)); 
mux6 mux_3297 (.in({n14305_0, n14304_0, n14247_0, n14246_0, n14231_0, n14230_1}), .out(n6962), .config_in(config_chain[9893:9891]), .config_rst(config_rst)); 
mux6 mux_3298 (.in({n11421_0, n11420_0, n11413_0, n11412_0, n11405_0, n11404_0}), .out(n6963), .config_in(config_chain[9896:9894]), .config_rst(config_rst)); 
mux6 mux_3299 (.in({n14033_0, n14032_0, n14025_0, n14024_0, n14017_0, n14016_0}), .out(n6964), .config_in(config_chain[9899:9897]), .config_rst(config_rst)); 
mux6 mux_3300 (.in({n11665_0, n11664_0, n11651_0, n11650_0, n11635_0, n11634_1}), .out(n6965), .config_in(config_chain[9902:9900]), .config_rst(config_rst)); 
mux6 mux_3301 (.in({n14269_0, n14268_0, n14263_0, n14262_0/**/, n14255_0, n14254_0}), .out(n6966), .config_in(config_chain[9905:9903]), .config_rst(config_rst)); 
mux6 mux_3302 (.in({n11437_0/**/, n11436_0, n11363_0, n11362_1, n11355_0, n11354_1}), .out(n6967), .config_in(config_chain[9908:9906]), .config_rst(config_rst)); 
mux6 mux_3303 (.in({n14041_0, n14040_0, n13981_0, n13980_0, n13967_0, n13966_1}), .out(n6968), .config_in(config_chain[9911:9909]), .config_rst(config_rst)); 
mux6 mux_3304 (.in({n11687_0, n11686_0, n11681_0, n11680_0, n11673_0, n11672_0}), .out(n6969), .config_in(config_chain[9914:9912]), .config_rst(config_rst)); 
mux6 mux_3305 (.in({n14291_0, n14290_0, n14285_0, n14284_0, n14277_0, n14276_0}), .out(n6970), .config_in(config_chain[9917:9915]), .config_rst(config_rst)); 
mux6 mux_3306 (.in({n11385_0, n11384_0, n11377_0, n11376_0, n11371_0, n11370_1}), .out(n6971), .config_in(config_chain[9920:9918]), .config_rst(config_rst)); 
mux6 mux_3307 (.in({n14003_0, n14002_0, n13989_0, n13988_0, n13975_0, n13974_1}), .out(n6972), .config_in(config_chain[9923:9921]), .config_rst(config_rst)); 
mux6 mux_3308 (.in({n11703_0, n11702_0, n11695_0, n11694_0, n11621_0, n11620_1}), .out(n6973), .config_in(config_chain[9926:9924]), .config_rst(config_rst)); 
mux6 mux_3309 (.in({n14307_0, n14306_0/**/, n14233_0, n14232_1, n14225_0, n14224_1}), .out(n6974), .config_in(config_chain[9929:9927]), .config_rst(config_rst)); 
mux6 mux_3310 (.in({n11423_0, n11422_0/**/, n11407_0, n11406_0, n11393_0, n11392_0}), .out(n6975), .config_in(config_chain[9932:9930]), .config_rst(config_rst)); 
mux6 mux_3311 (.in({n14027_0, n14026_0, n14019_0, n14018_0, n14011_0/**/, n14010_0}), .out(n6976), .config_in(config_chain[9935:9933]), .config_rst(config_rst)); 
mux6 mux_3312 (.in({n11653_0, n11652_0, n11645_0, n11644_0, n11637_0, n11636_1}), .out(n6977), .config_in(config_chain[9938:9936]), .config_rst(config_rst)); 
mux6 mux_3313 (.in({n14271_0, n14270_0/**/, n14257_0, n14256_0, n14241_0, n14240_1}), .out(n6978), .config_in(config_chain[9941:9939]), .config_rst(config_rst)); 
mux6 mux_3314 (.in({n11431_0/**/, n11430_0, n11415_0, n11414_0, n11357_0, n11356_1}), .out(n6979), .config_in(config_chain[9944:9942]), .config_rst(config_rst)); 
mux6 mux_3315 (.in({n14043_0, n14042_0, n14035_0, n14034_0/**/, n13961_0, n13960_1}), .out(n6980), .config_in(config_chain[9947:9945]), .config_rst(config_rst)); 
mux6 mux_3316 (.in({n11675_0, n11674_0, n11667_0, n11666_0, n11661_0, n11660_0}), .out(n6981), .config_in(config_chain[9950:9948]), .config_rst(config_rst)); 
mux6 mux_3317 (.in({n14293_0, n14292_0, n14279_0, n14278_0/**/, n14265_0, n14264_0}), .out(n6982), .config_in(config_chain[9953:9951]), .config_rst(config_rst)); 
mux6 mux_3318 (.in({n11379_0, n11378_0, n11373_0, n11372_1, n11365_0, n11364_1}), .out(n6983), .config_in(config_chain[9956:9954]), .config_rst(config_rst)); 
mux6 mux_3319 (.in({n13991_0, n13990_0, n13983_0/**/, n13982_0, n13977_0, n13976_1}), .out(n6984), .config_in(config_chain[9959:9957]), .config_rst(config_rst)); 
mux6 mux_3320 (.in({n11697_0, n11696_0, n11683_0, n11682_0, n11623_0/**/, n11622_1}), .out(n6985), .config_in(config_chain[9962:9960]), .config_rst(config_rst)); 
mux6 mux_3321 (.in({n14309_0, n14308_0, n14301_0/**/, n14300_0, n14227_0, n14226_1}), .out(n6986), .config_in(config_chain[9965:9963]), .config_rst(config_rst)); 
mux6 mux_3322 (.in({n11409_0, n11408_0, n11401_0, n11400_0, n11395_0, n11394_0}), .out(n6987), .config_in(config_chain[9968:9966]), .config_rst(config_rst)); 
mux6 mux_3323 (.in({n14013_0, n14012_0, n14005_0, n14004_0, n13999_0, n13998_0}), .out(n6988), .config_in(config_chain[9971:9969]), .config_rst(config_rst)); 
mux6 mux_3324 (.in({n11705_0, n11704_0, n11647_0, n11646_0/**/, n11631_0, n11630_1}), .out(n6989), .config_in(config_chain[9974:9972]), .config_rst(config_rst)); 
mux6 mux_3325 (.in({n14251_0/**/, n14250_0, n14243_0, n14242_1, n14235_0, n14234_1}), .out(n6990), .config_in(config_chain[9977:9975]), .config_rst(config_rst)); 
mux6 mux_3326 (.in({n11433_0, n11432_0/**/, n11425_0, n11424_0, n11417_0, n11416_0}), .out(n6991), .config_in(config_chain[9980:9978]), .config_rst(config_rst)); 
mux6 mux_3327 (.in({n14037_0, n14036_0, n14021_0, n14020_0/**/, n13963_0, n13962_1}), .out(n6992), .config_in(config_chain[9983:9981]), .config_rst(config_rst)); 
mux6 mux_3328 (.in({n11707_0, n11706_0, n11669_0, n11668_0/**/, n11655_0, n11654_0}), .out(n6993), .config_in(config_chain[9986:9984]), .config_rst(config_rst)); 
mux6 mux_3329 (.in({n14311_0/**/, n14310_0, n14281_0, n14280_0, n14273_0, n14272_0}), .out(n6994), .config_in(config_chain[9989:9987]), .config_rst(config_rst)); 
mux6 mux_3330 (.in({n11381_0, n11380_0, n11367_0, n11366_1, n11353_0, n11352_1}), .out(n6995), .config_in(config_chain[9992:9990]), .config_rst(config_rst)); 
mux6 mux_3331 (.in({n13985_0, n13984_0, n13971_0, n13970_1, n13957_0, n13956_1}), .out(n6996), .config_in(config_chain[9995:9993]), .config_rst(config_rst)); 
mux6 mux_3332 (.in({n11691_0, n11690_0, n11677_0, n11676_0, n11597_0, n11596_1}), .out(n6997), .config_in(config_chain[9998:9996]), .config_rst(config_rst)); 
mux6 mux_3333 (.in({n14303_0, n14302_0, n14295_0/**/, n14294_0, n14201_0, n14200_1}), .out(n6998), .config_in(config_chain[10001:9999]), .config_rst(config_rst)); 
mux6 mux_3334 (.in({n11403_0, n11402_0, n11389_0, n11388_0, n11375_0, n11374_1}), .out(n6999), .config_in(config_chain[10004:10002]), .config_rst(config_rst)); 
mux6 mux_3335 (.in({n14007_0, n14006_0, n14001_0, n14000_0/**/, n13993_0, n13992_0}), .out(n7000), .config_in(config_chain[10007:10005]), .config_rst(config_rst)); 
mux6 mux_3336 (.in({n11633_0, n11632_1, n11625_0, n11624_1, n11619_0, n11618_1/**/}), .out(n7001), .config_in(config_chain[10010:10008]), .config_rst(config_rst)); 
mux6 mux_3337 (.in({n14253_0/**/, n14252_0, n14237_0, n14236_1, n14223_0, n14222_1}), .out(n7002), .config_in(config_chain[10013:10011]), .config_rst(config_rst)); 
mux6 mux_3338 (.in({n11427_0, n11426_0/**/, n11419_0, n11418_0, n11411_0, n11410_0}), .out(n7003), .config_in(config_chain[10016:10014]), .config_rst(config_rst)); 
mux6 mux_3339 (.in({n14039_0, n14038_0, n14031_0, n14030_0/**/, n14023_0, n14022_0}), .out(n7004), .config_in(config_chain[10019:10017]), .config_rst(config_rst)); 
mux6 mux_3340 (.in({n11657_0/**/, n11656_0, n11649_0, n11648_0, n11641_0, n11640_1}), .out(n7005), .config_in(config_chain[10022:10020]), .config_rst(config_rst)); 
mux6 mux_3341 (.in({n14275_0/**/, n14274_0, n14261_0, n14260_0, n14245_0, n14244_1}), .out(n7006), .config_in(config_chain[10025:10023]), .config_rst(config_rst)); 
mux6 mux_3342 (.in({n11441_0, n11440_0, n11435_0, n11434_0/**/, n11361_0, n11360_1}), .out(n7007), .config_in(config_chain[10028:10026]), .config_rst(config_rst)); 
mux6 mux_3343 (.in({n14045_0, n14044_0/**/, n13973_0, n13972_1, n13965_0, n13964_1}), .out(n7008), .config_in(config_chain[10031:10029]), .config_rst(config_rst)); 
mux6 mux_3344 (.in({n11693_0/**/, n11692_0, n11679_0, n11678_0, n11663_0, n11662_0}), .out(n7009), .config_in(config_chain[10034:10032]), .config_rst(config_rst)); 
mux6 mux_3345 (.in({n14297_0, n14296_0/**/, n14289_0, n14288_0, n14283_0, n14282_0}), .out(n7010), .config_in(config_chain[10037:10035]), .config_rst(config_rst)); 
mux6 mux_3346 (.in({n11391_0, n11390_0, n11383_0, n11382_0/**/, n11311_0, n11310_2}), .out(n7011), .config_in(config_chain[10040:10038]), .config_rst(config_rst)); 
mux6 mux_3347 (.in({n14009_0, n14008_0, n13995_0, n13994_0, n13915_0, n13914_2}), .out(n7012), .config_in(config_chain[10043:10041]), .config_rst(config_rst)); 
mux6 mux_3348 (.in({n11951_0, n11950_0, n11935_0, n11934_0, n11921_0, n11920_0}), .out(n7059), .config_in(config_chain[10046:10044]), .config_rst(config_rst)); 
mux6 mux_3349 (.in({n14313_0, n14312_0, n14297_0, n14296_0, n14283_0, n14282_0}), .out(n7060), .config_in(config_chain[10049:10047]), .config_rst(config_rst)); 
mux6 mux_3350 (.in({n11643_0, n11642_0, n11635_0, n11634_1, n11627_0, n11626_1}), .out(n7061), .config_in(config_chain[10052:10050]), .config_rst(config_rst)); 
mux6 mux_3351 (.in({n14011_0, n14010_0, n14003_0, n14002_0, n13995_0, n13994_1/**/}), .out(n7062), .config_in(config_chain[10055:10053]), .config_rst(config_rst)); 
mux6 mux_3352 (.in({n11959_0, n11958_0, n11943_0, n11942_0, n11885_0, n11884_1}), .out(n7063), .config_in(config_chain[10058:10056]), .config_rst(config_rst)); 
mux6 mux_3353 (.in({n14329_0, n14328_0, n14321_0, n14320_0, n14247_0, n14246_1}), .out(n7064), .config_in(config_chain[10061:10059]), .config_rst(config_rst)); 
mux6 mux_3354 (.in({n11673_0, n11672_0, n11665_0, n11664_0, n11659_0, n11658_0}), .out(n7065), .config_in(config_chain[10064:10062]), .config_rst(config_rst)); 
mux6 mux_3355 (.in({n14047_0/**/, n14046_0, n14033_0, n14032_0, n14019_0, n14018_0}), .out(n7066), .config_in(config_chain[10067:10065]), .config_rst(config_rst)); 
mux6 mux_3356 (.in({n11907_0, n11906_0, n11901_0, n11900_1/**/, n11893_0, n11892_1}), .out(n7067), .config_in(config_chain[10070:10068]), .config_rst(config_rst)); 
mux6 mux_3357 (.in({n14269_0, n14268_0, n14263_0, n14262_1, n14255_0, n14254_1}), .out(n7068), .config_in(config_chain[10073:10071]), .config_rst(config_rst)); 
mux6 mux_3358 (.in({n11695_0, n11694_0, n11687_0, n11686_0, n11681_0, n11680_0}), .out(n7069), .config_in(config_chain[10076:10074]), .config_rst(config_rst)); 
mux6 mux_3359 (.in({n14055_0, n14054_0, n14041_0, n14040_0, n13981_0, n13980_1/**/}), .out(n7070), .config_in(config_chain[10079:10077]), .config_rst(config_rst)); 
mux6 mux_3360 (.in({n11929_0, n11928_0, n11923_0, n11922_0, n11915_0, n11914_0}), .out(n7071), .config_in(config_chain[10082:10080]), .config_rst(config_rst)); 
mux6 mux_3361 (.in({n14299_0/**/, n14298_0, n14291_0, n14290_0, n14285_0, n14284_0}), .out(n7072), .config_in(config_chain[10085:10083]), .config_rst(config_rst)); 
mux6 mux_3362 (.in({n11703_0, n11702_0, n11645_0/**/, n11644_0, n11629_0, n11628_1}), .out(n7073), .config_in(config_chain[10088:10086]), .config_rst(config_rst)); 
mux6 mux_3363 (.in({n14005_0/**/, n14004_0, n13997_0, n13996_1, n13989_0, n13988_1}), .out(n7074), .config_in(config_chain[10091:10089]), .config_rst(config_rst)); 
mux6 mux_3364 (.in({n11961_0, n11960_0/**/, n11953_0, n11952_0, n11945_0, n11944_0}), .out(n7075), .config_in(config_chain[10094:10092]), .config_rst(config_rst)); 
mux6 mux_3365 (.in({n14323_0, n14322_0/**/, n14307_0, n14306_0, n14249_0, n14248_1}), .out(n7076), .config_in(config_chain[10097:10095]), .config_rst(config_rst)); 
mux6 mux_3366 (.in({n11667_0, n11666_0, n11653_0/**/, n11652_0, n11637_0, n11636_1}), .out(n7077), .config_in(config_chain[10100:10098]), .config_rst(config_rst)); 
mux6 mux_3367 (.in({n14027_0, n14026_0, n14021_0, n14020_0, n14013_0, n14012_0}), .out(n7078), .config_in(config_chain[10103:10101]), .config_rst(config_rst)); 
mux6 mux_3368 (.in({n11969_0, n11968_0, n11895_0, n11894_1, n11887_0, n11886_1}), .out(n7079), .config_in(config_chain[10106:10104]), .config_rst(config_rst)); 
mux6 mux_3369 (.in({n14331_0, n14330_0/**/, n14271_0, n14270_0, n14257_0, n14256_1}), .out(n7080), .config_in(config_chain[10109:10107]), .config_rst(config_rst)); 
mux6 mux_3370 (.in({n11689_0, n11688_0/**/, n11683_0, n11682_0, n11675_0, n11674_0}), .out(n7081), .config_in(config_chain[10112:10110]), .config_rst(config_rst)); 
mux6 mux_3371 (.in({n14057_0, n14056_0, n14049_0, n14048_0, n14043_0/**/, n14042_0}), .out(n7082), .config_in(config_chain[10115:10113]), .config_rst(config_rst)); 
mux6 mux_3372 (.in({n11931_0, n11930_0, n11917_0, n11916_0, n11903_0, n11902_1}), .out(n7083), .config_in(config_chain[10118:10116]), .config_rst(config_rst)); 
mux6 mux_3373 (.in({n14293_0, n14292_0, n14287_0, n14286_0, n14279_0/**/, n14278_0}), .out(n7084), .config_in(config_chain[10121:10119]), .config_rst(config_rst)); 
mux6 mux_3374 (.in({n11705_0, n11704_0, n11631_0, n11630_1, n11623_0, n11622_1}), .out(n7085), .config_in(config_chain[10124:10122]), .config_rst(config_rst)); 
mux6 mux_3375 (.in({n14065_0, n14064_0, n13991_0, n13990_1, n13983_0, n13982_1}), .out(n7086), .config_in(config_chain[10127:10125]), .config_rst(config_rst)); 
mux6 mux_3376 (.in({n11955_0, n11954_0, n11939_0, n11938_0, n11925_0/**/, n11924_0}), .out(n7087), .config_in(config_chain[10130:10128]), .config_rst(config_rst)); 
mux6 mux_3377 (.in({n14317_0/**/, n14316_0, n14309_0, n14308_0, n14301_0, n14300_0}), .out(n7088), .config_in(config_chain[10133:10131]), .config_rst(config_rst)); 
mux6 mux_3378 (.in({n11655_0/**/, n11654_0, n11647_0, n11646_0, n11639_0, n11638_1}), .out(n7089), .config_in(config_chain[10136:10134]), .config_rst(config_rst)); 
mux6 mux_3379 (.in({n14029_0, n14028_0, n14015_0, n14014_0/**/, n13999_0, n13998_1}), .out(n7090), .config_in(config_chain[10139:10137]), .config_rst(config_rst)); 
mux6 mux_3380 (.in({n11963_0, n11962_0, n11927_0, n11926_0, n11889_0, n11888_1}), .out(n7091), .config_in(config_chain[10142:10140]), .config_rst(config_rst)); 
mux6 mux_3381 (.in({n14289_0, n14288_0, n14259_0, n14258_1, n14251_0, n14250_1}), .out(n7092), .config_in(config_chain[10145:10143]), .config_rst(config_rst)); 
mux6 mux_3382 (.in({n11707_0, n11706_0/**/, n11691_0, n11690_0, n11677_0, n11676_0}), .out(n7093), .config_in(config_chain[10148:10146]), .config_rst(config_rst)); 
mux6 mux_3383 (.in({n14067_0, n14066_0, n14051_0, n14050_0, n14037_0, n14036_0/**/}), .out(n7094), .config_in(config_chain[10151:10149]), .config_rst(config_rst)); 
mux6 mux_3384 (.in({n11949_0, n11948_0, n11911_0/**/, n11910_0, n11897_0, n11896_1}), .out(n7095), .config_in(config_chain[10154:10152]), .config_rst(config_rst)); 
mux6 mux_3385 (.in({n14311_0, n14310_0, n14281_0, n14280_0, n14273_0, n14272_0}), .out(n7096), .config_in(config_chain[10157:10155]), .config_rst(config_rst)); 
mux6 mux_3386 (.in({n11699_0, n11698_0, n11625_0, n11624_1, n11597_0, n11596_1}), .out(n7097), .config_in(config_chain[10160:10158]), .config_rst(config_rst)); 
mux6 mux_3387 (.in({n14059_0, n14058_0/**/, n13985_0, n13984_1, n13979_0, n13978_1}), .out(n7098), .config_in(config_chain[10163:10161]), .config_rst(config_rst)); 
mux6 mux_3388 (.in({n11941_0, n11940_0, n11933_0, n11932_0, n11829_0, n11828_2}), .out(n7099), .config_in(config_chain[10166:10164]), .config_rst(config_rst)); 
mux6 mux_3389 (.in({n14319_0, n14318_0/**/, n14303_0, n14302_0, n14201_0, n14200_2}), .out(n7100), .config_in(config_chain[10169:10167]), .config_rst(config_rst)); 
mux6 mux_3390 (.in({n11649_0, n11648_0/**/, n11641_0, n11640_1, n11633_0, n11632_1}), .out(n7101), .config_in(config_chain[10172:10170]), .config_rst(config_rst)); 
mux6 mux_3391 (.in({n14017_0, n14016_0, n14009_0, n14008_0/**/, n14001_0, n14000_1}), .out(n7102), .config_in(config_chain[10175:10173]), .config_rst(config_rst)); 
mux6 mux_3392 (.in({n11965_0, n11964_0, n11957_0, n11956_0/**/, n11861_0, n11860_1}), .out(n7103), .config_in(config_chain[10178:10176]), .config_rst(config_rst)); 
mux6 mux_3393 (.in({n14327_0, n14326_0, n14253_0, n14252_1, n14223_0, n14222_1}), .out(n7104), .config_in(config_chain[10181:10179]), .config_rst(config_rst)); 
mux6 mux_3394 (.in({n11671_0, n11670_0, n11663_0, n11662_0, n11657_0, n11656_0/**/}), .out(n7105), .config_in(config_chain[10184:10182]), .config_rst(config_rst)); 
mux6 mux_3395 (.in({n14039_0, n14038_0, n14031_0, n14030_0, n14023_0, n14022_0}), .out(n7106), .config_in(config_chain[10187:10185]), .config_rst(config_rst)); 
mux6 mux_3396 (.in({n11913_0/**/, n11912_0, n11899_0, n11898_1, n11883_0, n11882_1}), .out(n7107), .config_in(config_chain[10190:10188]), .config_rst(config_rst)); 
mux6 mux_3397 (.in({n14275_0, n14274_0, n14267_0, n14266_1, n14261_0/**/, n14260_1}), .out(n7108), .config_in(config_chain[10193:10191]), .config_rst(config_rst)); 
mux6 mux_3398 (.in({n11701_0, n11700_0, n11693_0, n11692_0, n11685_0, n11684_0/**/}), .out(n7109), .config_in(config_chain[10196:10194]), .config_rst(config_rst)); 
mux6 mux_3399 (.in({n14061_0, n14060_0/**/, n14045_0, n14044_0, n13987_0, n13986_1}), .out(n7110), .config_in(config_chain[10199:10197]), .config_rst(config_rst)); 
mux6 mux_3400 (.in({n12225_0, n12224_0, n12169_0, n12168_0, n12153_0, n12152_1}), .out(n7157), .config_in(config_chain[10202:10200]), .config_rst(config_rst)); 
mux6 mux_3401 (.in({n14347_0, n14346_0/**/, n14291_0, n14290_0, n14275_0, n14274_1}), .out(n7158), .config_in(config_chain[10205:10203]), .config_rst(config_rst)); 
mux6 mux_3402 (.in({n11951_0, n11950_0, n11943_0, n11942_0, n11935_0/**/, n11934_0}), .out(n7159), .config_in(config_chain[10208:10206]), .config_rst(config_rst)); 
mux6 mux_3403 (.in({n14077_0, n14076_0, n14069_0, n14068_0, n14061_0, n14060_0}), .out(n7160), .config_in(config_chain[10211:10209]), .config_rst(config_rst)); 
mux6 mux_3404 (.in({n12191_0, n12190_0, n12177_0, n12176_0/**/, n12161_0, n12160_1}), .out(n7161), .config_in(config_chain[10214:10212]), .config_rst(config_rst)); 
mux6 mux_3405 (.in({n14313_0, n14312_0/**/, n14307_0, n14306_0, n14299_0, n14298_0}), .out(n7162), .config_in(config_chain[10217:10215]), .config_rst(config_rst)); 
mux6 mux_3406 (.in({n11967_0, n11966_0, n11893_0, n11892_1, n11885_0, n11884_1}), .out(n7163), .config_in(config_chain[10220:10218]), .config_rst(config_rst)); 
mux6 mux_3407 (.in({n14085_0, n14084_0, n14025_0, n14024_0/**/, n14011_0, n14010_1}), .out(n7164), .config_in(config_chain[10223:10221]), .config_rst(config_rst)); 
mux6 mux_3408 (.in({n12211_0, n12210_0, n12207_0, n12206_0, n12199_0, n12198_0}), .out(n7165), .config_in(config_chain[10226:10224]), .config_rst(config_rst)); 
mux6 mux_3409 (.in({n14333_0, n14332_0, n14329_0, n14328_0, n14321_0, n14320_0}), .out(n7166), .config_in(config_chain[10229:10227]), .config_rst(config_rst)); 
mux6 mux_3410 (.in({n11915_0, n11914_0, n11907_0, n11906_0, n11901_0, n11900_1}), .out(n7167), .config_in(config_chain[10232:10230]), .config_rst(config_rst)); 
mux6 mux_3411 (.in({n14047_0, n14046_0, n14033_0, n14032_0, n14019_0, n14018_1/**/}), .out(n7168), .config_in(config_chain[10235:10233]), .config_rst(config_rst)); 
mux6 mux_3412 (.in({n12227_0, n12226_0, n12219_0, n12218_0, n12147_0, n12146_1}), .out(n7169), .config_in(config_chain[10238:10236]), .config_rst(config_rst)); 
mux6 mux_3413 (.in({n14349_0, n14348_0/**/, n14277_0, n14276_1, n14269_0, n14268_1}), .out(n7170), .config_in(config_chain[10241:10239]), .config_rst(config_rst)); 
mux6 mux_3414 (.in({n11953_0, n11952_0, n11937_0, n11936_0, n11923_0, n11922_0}), .out(n7171), .config_in(config_chain[10244:10242]), .config_rst(config_rst)); 
mux6 mux_3415 (.in({n14071_0, n14070_0, n14063_0/**/, n14062_0, n14055_0, n14054_0}), .out(n7172), .config_in(config_chain[10247:10245]), .config_rst(config_rst)); 
mux6 mux_3416 (.in({n12179_0/**/, n12178_0, n12171_0, n12170_0, n12163_0, n12162_1}), .out(n7173), .config_in(config_chain[10250:10248]), .config_rst(config_rst)); 
mux6 mux_3417 (.in({n14315_0, n14314_0, n14301_0, n14300_0/**/, n14285_0, n14284_1}), .out(n7174), .config_in(config_chain[10253:10251]), .config_rst(config_rst)); 
mux6 mux_3418 (.in({n11961_0, n11960_0, n11945_0, n11944_0, n11887_0, n11886_1}), .out(n7175), .config_in(config_chain[10256:10254]), .config_rst(config_rst)); 
mux6 mux_3419 (.in({n14087_0, n14086_0, n14079_0, n14078_0, n14005_0, n14004_1}), .out(n7176), .config_in(config_chain[10259:10257]), .config_rst(config_rst)); 
mux6 mux_3420 (.in({n12201_0, n12200_0, n12193_0, n12192_0, n12187_0, n12186_0/**/}), .out(n7177), .config_in(config_chain[10262:10260]), .config_rst(config_rst)); 
mux6 mux_3421 (.in({n14335_0, n14334_0, n14323_0, n14322_0, n14309_0, n14308_0}), .out(n7178), .config_in(config_chain[10265:10263]), .config_rst(config_rst)); 
mux6 mux_3422 (.in({n11909_0, n11908_0/**/, n11903_0, n11902_1, n11895_0, n11894_1}), .out(n7179), .config_in(config_chain[10268:10266]), .config_rst(config_rst)); 
mux6 mux_3423 (.in({n14035_0, n14034_0, n14027_0, n14026_0/**/, n14021_0, n14020_1}), .out(n7180), .config_in(config_chain[10271:10269]), .config_rst(config_rst)); 
mux6 mux_3424 (.in({n12221_0, n12220_0, n12209_0, n12208_0, n12149_0, n12148_1}), .out(n7181), .config_in(config_chain[10274:10272]), .config_rst(config_rst)); 
mux6 mux_3425 (.in({n14351_0, n14350_0/**/, n14343_0, n14342_0, n14271_0, n14270_1}), .out(n7182), .config_in(config_chain[10277:10275]), .config_rst(config_rst)); 
mux6 mux_3426 (.in({n11939_0, n11938_0, n11931_0, n11930_0, n11925_0, n11924_0}), .out(n7183), .config_in(config_chain[10280:10278]), .config_rst(config_rst)); 
mux6 mux_3427 (.in({n14057_0, n14056_0, n14049_0/**/, n14048_0, n14043_0, n14042_0}), .out(n7184), .config_in(config_chain[10283:10281]), .config_rst(config_rst)); 
mux6 mux_3428 (.in({n12229_0, n12228_0, n12173_0, n12172_0, n12157_0/**/, n12156_1}), .out(n7185), .config_in(config_chain[10286:10284]), .config_rst(config_rst)); 
mux6 mux_3429 (.in({n14295_0, n14294_0, n14287_0, n14286_1, n14279_0, n14278_1}), .out(n7186), .config_in(config_chain[10289:10287]), .config_rst(config_rst)); 
mux6 mux_3430 (.in({n11963_0, n11962_0/**/, n11955_0, n11954_0, n11947_0, n11946_0}), .out(n7187), .config_in(config_chain[10292:10290]), .config_rst(config_rst)); 
mux6 mux_3431 (.in({n14081_0, n14080_0/**/, n14065_0, n14064_0, n14007_0, n14006_1}), .out(n7188), .config_in(config_chain[10295:10293]), .config_rst(config_rst)); 
mux6 mux_3432 (.in({n12195_0, n12194_0, n12181_0, n12180_0, n12145_0, n12144_1}), .out(n7189), .config_in(config_chain[10298:10296]), .config_rst(config_rst)); 
mux6 mux_3433 (.in({n14325_0, n14324_0, n14317_0, n14316_0, n14267_0, n14266_1/**/}), .out(n7190), .config_in(config_chain[10301:10299]), .config_rst(config_rst)); 
mux6 mux_3434 (.in({n11927_0, n11926_0, n11911_0, n11910_0/**/, n11897_0, n11896_1}), .out(n7191), .config_in(config_chain[10304:10302]), .config_rst(config_rst)); 
mux6 mux_3435 (.in({n14045_0, n14044_0, n14029_0, n14028_0, n14015_0, n14014_1}), .out(n7192), .config_in(config_chain[10307:10305]), .config_rst(config_rst)); 
mux6 mux_3436 (.in({n12215_0, n12214_0, n12203_0, n12202_0, n12167_0, n12166_1}), .out(n7193), .config_in(config_chain[10310:10308]), .config_rst(config_rst)); 
mux6 mux_3437 (.in({n14345_0, n14344_0/**/, n14337_0, n14336_0, n14289_0, n14288_1}), .out(n7194), .config_in(config_chain[10313:10311]), .config_rst(config_rst)); 
mux6 mux_3438 (.in({n11949_0, n11948_0, n11933_0, n11932_0, n11919_0/**/, n11918_0}), .out(n7195), .config_in(config_chain[10316:10314]), .config_rst(config_rst)); 
mux6 mux_3439 (.in({n14051_0, n14050_0, n14037_0, n14036_0/**/, n13957_0, n13956_2}), .out(n7196), .config_in(config_chain[10319:10317]), .config_rst(config_rst)); 
mux6 mux_3440 (.in({n12189_0, n12188_0, n12159_0, n12158_1, n12151_0, n12150_1}), .out(n7197), .config_in(config_chain[10322:10320]), .config_rst(config_rst)); 
mux6 mux_3441 (.in({n14311_0, n14310_0, n14297_0, n14296_0, n14281_0, n14280_1}), .out(n7198), .config_in(config_chain[10325:10323]), .config_rst(config_rst)); 
mux6 mux_3442 (.in({n11957_0, n11956_0, n11941_0, n11940_0, n11861_0, n11860_1/**/}), .out(n7199), .config_in(config_chain[10328:10326]), .config_rst(config_rst)); 
mux6 mux_3443 (.in({n14083_0/**/, n14082_0, n14075_0, n14074_0, n13979_0, n13978_1}), .out(n7200), .config_in(config_chain[10331:10329]), .config_rst(config_rst)); 
mux6 mux_3444 (.in({n12183_0, n12182_0, n12175_0, n12174_0, n12091_0, n12090_2}), .out(n7201), .config_in(config_chain[10334:10332]), .config_rst(config_rst)); 
mux6 mux_3445 (.in({n14319_0, n14318_0, n14305_0, n14304_0, n14201_0, n14200_2}), .out(n7202), .config_in(config_chain[10337:10335]), .config_rst(config_rst)); 
mux6 mux_3446 (.in({n11965_0, n11964_0/**/, n11891_0, n11890_1, n11883_0, n11882_1}), .out(n7203), .config_in(config_chain[10340:10338]), .config_rst(config_rst)); 
mux6 mux_3447 (.in({n14017_0/**/, n14016_1, n14009_0, n14008_1, n14001_0, n14000_1}), .out(n7204), .config_in(config_chain[10343:10341]), .config_rst(config_rst)); 
mux6 mux_3448 (.in({n12217_0, n12216_0/**/, n12205_0, n12204_0, n12093_0, n12092_2}), .out(n7205), .config_in(config_chain[10346:10344]), .config_rst(config_rst)); 
mux6 mux_3449 (.in({n14339_0, n14338_0, n14327_0, n14326_0, n14245_0, n14244_1}), .out(n7206), .config_in(config_chain[10349:10347]), .config_rst(config_rst)); 
mux6 mux_3450 (.in({n11921_0, n11920_0, n11913_0, n11912_0, n11905_0, n11904_1}), .out(n7207), .config_in(config_chain[10352:10350]), .config_rst(config_rst)); 
mux6 mux_3451 (.in({n14053_0, n14052_0, n14039_0, n14038_0, n14023_0, n14022_1}), .out(n7208), .config_in(config_chain[10355:10353]), .config_rst(config_rst)); 
mux6 mux_3452 (.in({n12177_0, n12176_0, n12169_0, n12168_0, n12161_0, n12160_1}), .out(n7254), .config_in(config_chain[10358:10356]), .config_rst(config_rst)); 
mux6 mux_3453 (.in({n12219_0, n12218_0, n12211_0, n12210_0, n12207_0, n12206_0}), .out(n7257), .config_in(config_chain[10361:10359]), .config_rst(config_rst)); 
mux6 mux_3454 (.in({n12179_0, n12178_0, n12171_0, n12170_0, n12163_0, n12162_1/**/}), .out(n7260), .config_in(config_chain[10364:10362]), .config_rst(config_rst)); 
mux6 mux_3455 (.in({n12221_0, n12220_0, n12213_0, n12212_0, n12209_0, n12208_0}), .out(n7263), .config_in(config_chain[10367:10365]), .config_rst(config_rst)); 
mux6 mux_3456 (.in({n12173_0, n12172_0, n12165_0, n12164_1, n12157_0, n12156_1}), .out(n7266), .config_in(config_chain[10370:10368]), .config_rst(config_rst)); 
mux6 mux_3457 (.in({n12215_0, n12214_0, n12203_0, n12202_0, n12167_0, n12166_1}), .out(n7269), .config_in(config_chain[10373:10371]), .config_rst(config_rst)); 
mux6 mux_3458 (.in({n12175_0, n12174_0, n12159_0, n12158_1, n12091_0, n12090_2}), .out(n7272), .config_in(config_chain[10376:10374]), .config_rst(config_rst)); 
mux6 mux_3459 (.in({n12217_0, n12216_0, n12205_0, n12204_0, n12123_0, n12122_1}), .out(n7275), .config_in(config_chain[10379:10377]), .config_rst(config_rst)); 
mux6 mux_3460 (.in({n9893_0, n9892_0, n9839_0, n9838_0, n9825_0, n9824_1}), .out(n7302), .config_in(config_chain[10382:10380]), .config_rst(config_rst)); 
mux6 mux_3461 (.in({n9867_0, n9866_0, n9859_0, n9858_0, n9855_0, n9854_0}), .out(n7305), .config_in(config_chain[10385:10383]), .config_rst(config_rst)); 
mux6 mux_3462 (.in({n9895_0, n9894_0, n9827_0, n9826_1, n9819_0, n9818_1}), .out(n7308), .config_in(config_chain[10388:10386]), .config_rst(config_rst)); 
mux6 mux_3463 (.in({n9869_0, n9868_0, n9861_0, n9860_0, n9857_0, n9856_0}), .out(n7311), .config_in(config_chain[10391:10389]), .config_rst(config_rst)); 
mux6 mux_3464 (.in({n9897_0, n9896_0, n9829_0, n9828_1, n9821_0, n9820_1}), .out(n7314), .config_in(config_chain[10394:10392]), .config_rst(config_rst)); 
mux6 mux_3465 (.in({n9863_0, n9862_0, n9851_0, n9850_0, n9757_0, n9756_2}), .out(n7317), .config_in(config_chain[10397:10395]), .config_rst(config_rst)); 
mux6 mux_3466 (.in({n9891_0, n9890_0, n9823_0, n9822_1, n9749_0, n9748_2}), .out(n7320), .config_in(config_chain[10400:10398]), .config_rst(config_rst)); 
mux6 mux_3467 (.in({n9865_0, n9864_0, n9853_0, n9852_0, n9753_0, n9752_2}), .out(n7323), .config_in(config_chain[10403:10401]), .config_rst(config_rst)); 
mux6 mux_3468 (.in({n10133_0, n10132_0, n10119_0, n10118_0, n10107_0, n10106_0}), .out(n7351), .config_in(config_chain[10406:10404]), .config_rst(config_rst)); 
mux6 mux_3469 (.in({n14413_0, n14412_0, n14383_0, n14382_0, n14353_1, n14352_0}), .out(n7352), .config_in(config_chain[10409:10407]), .config_rst(config_rst)); 
mux6 mux_3470 (.in({n9839_0, n9838_0, n9833_0, n9832_1, n9825_0, n9824_1}), .out(n7353), .config_in(config_chain[10412:10410]), .config_rst(config_rst)); 
mux6 mux_3471 (.in({n14145_0, n14144_0, n14123_0, n14122_0, n14091_0, n14090_0}), .out(n7354), .config_in(config_chain[10415:10413]), .config_rst(config_rst)); 
mux6 mux_3472 (.in({n10141_0, n10140_0, n10127_0, n10126_0, n10073_0, n10072_1}), .out(n7355), .config_in(config_chain[10418:10416]), .config_rst(config_rst)); 
mux6 mux_3473 (.in({n14417_1, n14416_0, n14385_1, n14384_0, n14355_0, n14354_0}), .out(n7356), .config_in(config_chain[10421:10419]), .config_rst(config_rst)); 
mux6 mux_3474 (.in({n9867_0, n9866_0, n9859_0, n9858_0, n9855_0, n9854_0}), .out(n7357), .config_in(config_chain[10424:10422]), .config_rst(config_rst)); 
mux6 mux_3475 (.in({n14155_0, n14154_0, n14125_0, n14124_0, n14095_1, n14094_0}), .out(n7358), .config_in(config_chain[10427:10425]), .config_rst(config_rst)); 
mux6 mux_3476 (.in({n10093_0, n10092_0, n10089_0, n10088_1, n10081_0, n10080_1}), .out(n7359), .config_in(config_chain[10430:10428]), .config_rst(config_rst)); 
mux6 mux_3477 (.in({n14419_0, n14418_0, n14387_0, n14386_0, n14357_0, n14356_0}), .out(n7360), .config_in(config_chain[10433:10431]), .config_rst(config_rst)); 
mux6 mux_3478 (.in({n9887_0, n9886_0, n9879_0, n9878_0, n9875_0, n9874_0}), .out(n7361), .config_in(config_chain[10436:10434]), .config_rst(config_rst)); 
mux6 mux_3479 (.in({n14157_0, n14156_0, n14127_1, n14126_0, n14089_0, n14088_0}), .out(n7362), .config_in(config_chain[10439:10437]), .config_rst(config_rst)); 
mux6 mux_3480 (.in({n10113_0, n10112_0, n10109_0, n10108_0, n10101_0, n10100_0}), .out(n7363), .config_in(config_chain[10442:10440]), .config_rst(config_rst)); 
mux6 mux_3481 (.in({n14421_0, n14420_0, n14391_0, n14390_0, n14359_0, n14358_0}), .out(n7364), .config_in(config_chain[10445:10443]), .config_rst(config_rst)); 
mux6 mux_3482 (.in({n9895_0, n9894_0, n9841_0, n9840_0, n9827_0, n9826_1}), .out(n7365), .config_in(config_chain[10448:10446]), .config_rst(config_rst)); 
mux6 mux_3483 (.in({n14153_0, n14152_0, n14121_0, n14120_0, n14099_0, n14098_0}), .out(n7366), .config_in(config_chain[10451:10449]), .config_rst(config_rst)); 
mux6 mux_3484 (.in({n10143_0, n10142_0, n10135_0, n10134_0, n10129_0, n10128_0}), .out(n7367), .config_in(config_chain[10454:10452]), .config_rst(config_rst)); 
mux6 mux_3485 (.in({n14423_0, n14422_0, n14393_1, n14392_0, n14363_0, n14362_0}), .out(n7368), .config_in(config_chain[10457:10455]), .config_rst(config_rst)); 
mux6 mux_3486 (.in({n9861_0, n9860_0, n9849_0, n9848_0, n9835_0, n9834_1}), .out(n7369), .config_in(config_chain[10460:10458]), .config_rst(config_rst)); 
mux6 mux_3487 (.in({n14163_0, n14162_0, n14131_0, n14130_0, n14101_0, n14100_0}), .out(n7370), .config_in(config_chain[10463:10461]), .config_rst(config_rst)); 
mux6 mux_3488 (.in({n10151_0, n10150_0, n10083_0, n10082_1, n10075_0, n10074_1}), .out(n7371), .config_in(config_chain[10466:10464]), .config_rst(config_rst)); 
mux6 mux_3489 (.in({n14425_1, n14424_0, n14395_0, n14394_0, n14365_0, n14364_0}), .out(n7372), .config_in(config_chain[10469:10467]), .config_rst(config_rst)); 
mux6 mux_3490 (.in({n9881_0, n9880_0, n9877_0, n9876_0, n9869_0, n9868_0}), .out(n7373), .config_in(config_chain[10472:10470]), .config_rst(config_rst)); 
mux6 mux_3491 (.in({n14165_0, n14164_0, n14135_1, n14134_0, n14103_1, n14102_0}), .out(n7374), .config_in(config_chain[10475:10473]), .config_rst(config_rst)); 
mux6 mux_3492 (.in({n10115_0, n10114_0, n10103_0, n10102_0, n10091_0, n10090_1}), .out(n7375), .config_in(config_chain[10478:10476]), .config_rst(config_rst)); 
mux6 mux_3493 (.in({n14429_0, n14428_0, n14397_0, n14396_0, n14367_0, n14366_0}), .out(n7376), .config_in(config_chain[10481:10479]), .config_rst(config_rst)); 
mux6 mux_3494 (.in({n9897_0, n9896_0, n9829_0, n9828_1, n9821_0, n9820_1}), .out(n7377), .config_in(config_chain[10484:10482]), .config_rst(config_rst)); 
mux6 mux_3495 (.in({n14167_1, n14166_0, n14129_0, n14128_0, n14097_0, n14096_0}), .out(n7378), .config_in(config_chain[10487:10485]), .config_rst(config_rst)); 
mux6 mux_3496 (.in({n10137_0, n10136_0, n10123_0, n10122_0, n10111_0, n10110_0}), .out(n7379), .config_in(config_chain[10490:10488]), .config_rst(config_rst)); 
mux6 mux_3497 (.in({n14431_0, n14430_0, n14399_0, n14398_0, n14369_1, n14368_0}), .out(n7380), .config_in(config_chain[10493:10491]), .config_rst(config_rst)); 
mux6 mux_3498 (.in({n9851_0, n9850_0, n9843_0, n9842_0, n9837_0, n9836_1}), .out(n7381), .config_in(config_chain[10496:10494]), .config_rst(config_rst)); 
mux6 mux_3499 (.in({n14161_0, n14160_0, n14139_0, n14138_0, n14109_0, n14108_0}), .out(n7382), .config_in(config_chain[10499:10497]), .config_rst(config_rst)); 
mux6 mux_3500 (.in({n10145_0, n10144_0, n10077_0, n10076_1, n10009_0, n10008_2}), .out(n7383), .config_in(config_chain[10502:10500]), .config_rst(config_rst)); 
mux6 mux_3501 (.in({n14441_1, n14440_0, n14403_0, n14402_0, n14371_0, n14370_0}), .out(n7384), .config_in(config_chain[10505:10503]), .config_rst(config_rst)); 
mux6 mux_3502 (.in({n9883_0, n9882_0, n9871_0, n9870_0, n9757_0, n9756_2}), .out(n7385), .config_in(config_chain[10508:10506]), .config_rst(config_rst)); 
mux6 mux_3503 (.in({n14179_1, n14178_0, n14141_0, n14140_0, n14111_1, n14110_0}), .out(n7386), .config_in(config_chain[10511:10509]), .config_rst(config_rst)); 
mux6 mux_3504 (.in({n10097_0, n10096_0, n10085_0, n10084_1, n10011_0, n10010_2}), .out(n7387), .config_in(config_chain[10514:10512]), .config_rst(config_rst)); 
mux6 mux_3505 (.in({n14443_1, n14442_0, n14405_0, n14404_0, n14373_0, n14372_0}), .out(n7388), .config_in(config_chain[10517:10515]), .config_rst(config_rst)); 
mux6 mux_3506 (.in({n9891_0, n9890_0, n9823_0, n9822_1, n9747_0, n9746_2}), .out(n7389), .config_in(config_chain[10520:10518]), .config_rst(config_rst)); 
mux6 mux_3507 (.in({n14171_0, n14170_0, n14143_1, n14142_0, n14105_0, n14104_0}), .out(n7390), .config_in(config_chain[10523:10521]), .config_rst(config_rst)); 
mux6 mux_3508 (.in({n10153_0, n10152_0, n10125_0, n10124_0, n10117_0, n10116_0}), .out(n7391), .config_in(config_chain[10526:10524]), .config_rst(config_rst)); 
mux6 mux_3509 (.in({n14433_2, n14432_0, n14407_0, n14406_0, n14377_1, n14376_0}), .out(n7392), .config_in(config_chain[10529:10527]), .config_rst(config_rst)); 
mux6 mux_3510 (.in({n9845_0, n9844_0, n9831_0, n9830_1, n9751_0, n9750_2}), .out(n7393), .config_in(config_chain[10532:10530]), .config_rst(config_rst)); 
mux6 mux_3511 (.in({n14173_0, n14172_0, n14147_0, n14146_0, n14115_0, n14114_0}), .out(n7394), .config_in(config_chain[10535:10533]), .config_rst(config_rst)); 
mux6 mux_3512 (.in({n10147_0, n10146_0, n10139_0, n10138_0, n10003_0, n10002_2}), .out(n7395), .config_in(config_chain[10538:10536]), .config_rst(config_rst)); 
mux6 mux_3513 (.in({n14435_0, n14434_0, n14409_1, n14408_0, n14379_0, n14378_0}), .out(n7396), .config_in(config_chain[10541:10539]), .config_rst(config_rst)); 
mux6 mux_3514 (.in({n9865_0, n9864_0, n9853_0, n9852_0, n9753_0, n9752_2}), .out(n7397), .config_in(config_chain[10544:10542]), .config_rst(config_rst)); 
mux6 mux_3515 (.in({n14175_1, n14174_0, n14149_0, n14148_0, n14117_0, n14116_0}), .out(n7398), .config_in(config_chain[10547:10545]), .config_rst(config_rst)); 
mux6 mux_3516 (.in({n10099_0, n10098_0, n10087_0, n10086_1, n10005_0, n10004_2}), .out(n7399), .config_in(config_chain[10550:10548]), .config_rst(config_rst)); 
mux6 mux_3517 (.in({n14439_0, n14438_0, n14411_0, n14410_0, n14381_0, n14380_0}), .out(n7400), .config_in(config_chain[10553:10551]), .config_rst(config_rst)); 
mux6 mux_3518 (.in({n9893_0, n9892_0, n9885_0, n9884_0, n9755_0, n9754_2}), .out(n7401), .config_in(config_chain[10556:10554]), .config_rst(config_rst)); 
mux6 mux_3519 (.in({n14177_1, n14176_0, n14151_1, n14150_0, n14113_0, n14112_0}), .out(n7402), .config_in(config_chain[10559:10557]), .config_rst(config_rst)); 
mux6 mux_3520 (.in({n10405_0, n10404_0, n10349_0, n10348_0, n10335_0, n10334_1}), .out(n7449), .config_in(config_chain[10562:10560]), .config_rst(config_rst)); 
mux6 mux_3521 (.in({n14459_1, n14458_0, n14381_0, n14380_0, n14359_0, n14358_0}), .out(n7450), .config_in(config_chain[10565:10563]), .config_rst(config_rst)); 
mux6 mux_3522 (.in({n10133_0, n10132_0, n10127_0, n10126_0, n10119_0, n10118_0}), .out(n7451), .config_in(config_chain[10568:10566]), .config_rst(config_rst)); 
mux6 mux_3523 (.in({n14189_1, n14188_0, n14181_1, n14180_0, n14151_0, n14150_0}), .out(n7452), .config_in(config_chain[10571:10569]), .config_rst(config_rst)); 
mux6 mux_3524 (.in({n10369_0, n10368_0, n10357_0, n10356_0, n10343_0, n10342_1}), .out(n7453), .config_in(config_chain[10574:10572]), .config_rst(config_rst)); 
mux6 mux_3525 (.in({n14423_0, n14422_0, n14391_0, n14390_0, n14353_0, n14352_0}), .out(n7454), .config_in(config_chain[10577:10575]), .config_rst(config_rst)); 
mux6 mux_3526 (.in({n10149_0, n10148_0, n10081_0, n10080_1, n10073_0, n10072_1/**/}), .out(n7455), .config_in(config_chain[10580:10578]), .config_rst(config_rst)); 
mux6 mux_3527 (.in({n14197_1, n14196_0, n14123_0, n14122_0, n14093_0, n14092_0}), .out(n7456), .config_in(config_chain[10583:10581]), .config_rst(config_rst)); 
mux6 mux_3528 (.in({n10391_0, n10390_0, n10385_0, n10384_0, n10377_0, n10376_0}), .out(n7457), .config_in(config_chain[10586:10584]), .config_rst(config_rst)); 
mux6 mux_3529 (.in({n14445_1, n14444_0, n14417_0, n14416_0, n14385_0, n14384_0}), .out(n7458), .config_in(config_chain[10589:10587]), .config_rst(config_rst)); 
mux6 mux_3530 (.in({n10101_0, n10100_0/**/, n10093_0, n10092_0, n10089_0, n10088_1}), .out(n7459), .config_in(config_chain[10592:10590]), .config_rst(config_rst)); 
mux6 mux_3531 (.in({n14155_0, n14154_0, n14125_0, n14124_0, n14095_0, n14094_0}), .out(n7460), .config_in(config_chain[10595:10593]), .config_rst(config_rst)); 
mux6 mux_3532 (.in({n10407_0, n10406_0, n10399_0, n10398_0, n10329_0/**/, n10328_1}), .out(n7461), .config_in(config_chain[10598:10596]), .config_rst(config_rst)); 
mux6 mux_3533 (.in({n14461_1/**/, n14460_0, n14389_0, n14388_0, n14357_0, n14356_0}), .out(n7462), .config_in(config_chain[10601:10599]), .config_rst(config_rst)); 
mux6 mux_3534 (.in({n10135_0, n10134_0/**/, n10121_0, n10120_0, n10109_0, n10108_0}), .out(n7463), .config_in(config_chain[10604:10602]), .config_rst(config_rst)); 
mux6 mux_3535 (.in({n14183_1, n14182_0, n14159_0, n14158_0/**/, n14127_0, n14126_0}), .out(n7464), .config_in(config_chain[10607:10605]), .config_rst(config_rst)); 
mux6 mux_3536 (.in({n10359_0, n10358_0, n10351_0, n10350_0, n10345_0, n10344_1/**/}), .out(n7465), .config_in(config_chain[10610:10608]), .config_rst(config_rst)); 
mux6 mux_3537 (.in({n14421_0/**/, n14420_0, n14399_0, n14398_0, n14361_0, n14360_0}), .out(n7466), .config_in(config_chain[10613:10611]), .config_rst(config_rst)); 
mux6 mux_3538 (.in({n10143_0, n10142_0, n10129_0, n10128_0, n10075_0/**/, n10074_1}), .out(n7467), .config_in(config_chain[10616:10614]), .config_rst(config_rst)); 
mux6 mux_3539 (.in({n14199_1, n14198_0, n14191_1, n14190_0, n14099_0, n14098_0}), .out(n7468), .config_in(config_chain[10619:10617]), .config_rst(config_rst)); 
mux6 mux_3540 (.in({n10379_0, n10378_0, n10371_0, n10370_0, n10367_0, n10366_0}), .out(n7469), .config_in(config_chain[10622:10620]), .config_rst(config_rst)); 
mux6 mux_3541 (.in({n14447_1/**/, n14446_0, n14431_0, n14430_0, n14393_0, n14392_0}), .out(n7470), .config_in(config_chain[10625:10623]), .config_rst(config_rst)); 
mux6 mux_3542 (.in({n10095_0, n10094_0, n10091_0, n10090_1/**/, n10083_0, n10082_1}), .out(n7471), .config_in(config_chain[10628:10626]), .config_rst(config_rst)); 
mux6 mux_3543 (.in({n14163_0, n14162_0, n14133_0, n14132_0/**/, n14101_0, n14100_0}), .out(n7472), .config_in(config_chain[10631:10629]), .config_rst(config_rst)); 
mux6 mux_3544 (.in({n10401_0, n10400_0, n10387_0, n10386_0, n10331_0, n10330_1}), .out(n7473), .config_in(config_chain[10634:10632]), .config_rst(config_rst)); 
mux6 mux_3545 (.in({n14463_1, n14462_0, n14455_1, n14454_0/**/, n14365_0, n14364_0}), .out(n7474), .config_in(config_chain[10637:10635]), .config_rst(config_rst)); 
mux6 mux_3546 (.in({n10123_0, n10122_0, n10115_0, n10114_0/**/, n10111_0, n10110_0}), .out(n7475), .config_in(config_chain[10640:10638]), .config_rst(config_rst)); 
mux6 mux_3547 (.in({n14165_0, n14164_0, n14135_0, n14134_0, n14103_0, n14102_0/**/}), .out(n7476), .config_in(config_chain[10643:10641]), .config_rst(config_rst)); 
mux6 mux_3548 (.in({n10409_0, n10408_0, n10353_0, n10352_0, n10339_0, n10338_1}), .out(n7477), .config_in(config_chain[10646:10644]), .config_rst(config_rst)); 
mux6 mux_3549 (.in({n14429_0, n14428_0, n14397_0/**/, n14396_0, n14375_0, n14374_0}), .out(n7478), .config_in(config_chain[10649:10647]), .config_rst(config_rst)); 
mux6 mux_3550 (.in({n10145_0, n10144_0/**/, n10137_0, n10136_0, n10131_0, n10130_0}), .out(n7479), .config_in(config_chain[10652:10650]), .config_rst(config_rst)); 
mux6 mux_3551 (.in({n14193_1, n14192_0, n14167_0, n14166_0, n14107_0, n14106_0}), .out(n7480), .config_in(config_chain[10655:10653]), .config_rst(config_rst)); 
mux6 mux_3552 (.in({n10373_0, n10372_0, n10361_0, n10360_0, n10263_0, n10262_2}), .out(n7481), .config_in(config_chain[10658:10656]), .config_rst(config_rst)); 
mux6 mux_3553 (.in({n14439_0, n14438_0, n14401_0, n14400_0/**/, n14369_0, n14368_0}), .out(n7482), .config_in(config_chain[10661:10659]), .config_rst(config_rst)); 
mux6 mux_3554 (.in({n10097_0, n10096_0, n10085_0, n10084_1, n10009_0, n10008_2}), .out(n7483), .config_in(config_chain[10664:10662]), .config_rst(config_rst)); 
mux6 mux_3555 (.in({n14177_1, n14176_0, n14139_0, n14138_0, n14109_0, n14108_0}), .out(n7484), .config_in(config_chain[10667:10665]), .config_rst(config_rst)); 
mux6 mux_3556 (.in({n10395_0, n10394_0, n10381_0, n10380_0, n10265_0, n10264_2}), .out(n7485), .config_in(config_chain[10670:10668]), .config_rst(config_rst)); 
mux6 mux_3557 (.in({n14457_1, n14456_0, n14449_1/**/, n14448_0, n14441_0, n14440_0}), .out(n7486), .config_in(config_chain[10673:10671]), .config_rst(config_rst)); 
mux6 mux_3558 (.in({n10117_0, n10116_0/**/, n10105_0, n10104_0, n10011_0, n10010_2}), .out(n7487), .config_in(config_chain[10676:10674]), .config_rst(config_rst)); 
mux6 mux_3559 (.in({n14201_2, n14200_0, n14141_0, n14140_0, n14111_0, n14110_0}), .out(n7488), .config_in(config_chain[10679:10677]), .config_rst(config_rst)); 
mux6 mux_3560 (.in({n10341_0, n10340_1, n10333_0, n10332_1, n10267_0, n10266_2}), .out(n7489), .config_in(config_chain[10682:10680]), .config_rst(config_rst)); 
mux6 mux_3561 (.in({n14443_1, n14442_0, n14405_0, n14404_0, n14383_0, n14382_0}), .out(n7490), .config_in(config_chain[10685:10683]), .config_rst(config_rst)); 
mux6 mux_3562 (.in({n10139_0, n10138_0, n10125_0, n10124_0, n10003_0, n10002_2}), .out(n7491), .config_in(config_chain[10688:10686]), .config_rst(config_rst)); 
mux6 mux_3563 (.in({n14195_1/**/, n14194_0, n14187_1, n14186_0, n14171_0, n14170_0}), .out(n7492), .config_in(config_chain[10691:10689]), .config_rst(config_rst)); 
mux6 mux_3564 (.in({n10389_0, n10388_0, n10363_0, n10362_0, n10355_0, n10354_0}), .out(n7493), .config_in(config_chain[10694:10692]), .config_rst(config_rst)); 
mux6 mux_3565 (.in({n14433_2, n14432_0, n14415_0/**/, n14414_0, n14377_0, n14376_0}), .out(n7494), .config_in(config_chain[10697:10695]), .config_rst(config_rst)); 
mux6 mux_3566 (.in({n10147_0, n10146_0, n10079_0, n10078_1, n10005_0, n10004_2}), .out(n7495), .config_in(config_chain[10700:10698]), .config_rst(config_rst)); 
mux6 mux_3567 (.in({n14173_0, n14172_0, n14147_0, n14146_0, n14115_0/**/, n14114_0}), .out(n7496), .config_in(config_chain[10703:10701]), .config_rst(config_rst)); 
mux6 mux_3568 (.in({n10411_0, n10410_0, n10397_0, n10396_0, n10383_0, n10382_0}), .out(n7497), .config_in(config_chain[10706:10704]), .config_rst(config_rst)); 
mux6 mux_3569 (.in({n14451_1, n14450_0, n14437_0, n14436_0, n14409_0, n14408_0}), .out(n7498), .config_in(config_chain[10709:10707]), .config_rst(config_rst)); 
mux6 mux_3570 (.in({n10107_0, n10106_0/**/, n10099_0, n10098_0, n10007_0, n10006_2}), .out(n7499), .config_in(config_chain[10712:10710]), .config_rst(config_rst)); 
mux6 mux_3571 (.in({n14175_0, n14174_0, n14149_0/**/, n14148_0, n14119_0, n14118_0}), .out(n7500), .config_in(config_chain[10715:10713]), .config_rst(config_rst)); 
mux6 mux_3572 (.in({n10651_0, n10650_0, n10635_0, n10634_0, n10621_0, n10620_0}), .out(n7547), .config_in(config_chain[10718:10716]), .config_rst(config_rst)); 
mux6 mux_3573 (.in({n14467_1, n14466_0, n14451_0, n14450_0, n14409_0, n14408_0}), .out(n7548), .config_in(config_chain[10721:10719]), .config_rst(config_rst)); 
mux6 mux_3574 (.in({n10349_0, n10348_0, n10343_0, n10342_1, n10335_0, n10334_1}), .out(n7549), .config_in(config_chain[10724:10722]), .config_rst(config_rst)); 
mux6 mux_3575 (.in({n14149_0, n14148_0, n14127_0, n14126_0, n14095_0, n14094_0}), .out(n7550), .config_in(config_chain[10727:10725]), .config_rst(config_rst)); 
mux6 mux_3576 (.in({n10659_0, n10658_0, n10643_0, n10642_0, n10587_0, n10586_1}), .out(n7551), .config_in(config_chain[10730:10728]), .config_rst(config_rst)); 
mux6 mux_3577 (.in({n14483_1, n14482_0, n14475_1, n14474_0, n14359_0, n14358_0}), .out(n7552), .config_in(config_chain[10733:10731]), .config_rst(config_rst)); 
mux6 mux_3578 (.in({n10377_0, n10376_0, n10369_0, n10368_0, n10365_0, n10364_0}), .out(n7553), .config_in(config_chain[10736:10734]), .config_rst(config_rst)); 
mux6 mux_3579 (.in({n14203_1, n14202_0, n14189_0, n14188_0, n14159_0, n14158_0}), .out(n7554), .config_in(config_chain[10739:10737]), .config_rst(config_rst)); 
mux6 mux_3580 (.in({n10607_0, n10606_0/**/, n10603_0, n10602_1, n10595_0, n10594_1}), .out(n7555), .config_in(config_chain[10742:10740]), .config_rst(config_rst)); 
mux6 mux_3581 (.in({n14423_0, n14422_0, n14391_0, n14390_0, n14353_0, n14352_0}), .out(n7556), .config_in(config_chain[10745:10743]), .config_rst(config_rst)); 
mux6 mux_3582 (.in({n10399_0, n10398_0, n10391_0, n10390_0, n10385_0, n10384_0}), .out(n7557), .config_in(config_chain[10748:10746]), .config_rst(config_rst)); 
mux6 mux_3583 (.in({n14211_1, n14210_0, n14197_0, n14196_0, n14093_0, n14092_0}), .out(n7558), .config_in(config_chain[10751:10749]), .config_rst(config_rst)); 
mux6 mux_3584 (.in({n10629_0, n10628_0, n10623_0, n10622_0, n10615_0, n10614_0}), .out(n7559), .config_in(config_chain[10754:10752]), .config_rst(config_rst)); 
mux6 mux_3585 (.in({n14453_0, n14452_0, n14445_0, n14444_0, n14417_0/**/, n14416_0}), .out(n7560), .config_in(config_chain[10757:10755]), .config_rst(config_rst)); 
mux6 mux_3586 (.in({n10407_0, n10406_0/**/, n10351_0, n10350_0, n10337_0, n10336_1}), .out(n7561), .config_in(config_chain[10760:10758]), .config_rst(config_rst)); 
mux6 mux_3587 (.in({n14157_0, n14156_0, n14125_0, n14124_0, n14103_0/**/, n14102_0}), .out(n7562), .config_in(config_chain[10763:10761]), .config_rst(config_rst)); 
mux6 mux_3588 (.in({n10661_0, n10660_0, n10653_0/**/, n10652_0, n10645_0, n10644_0}), .out(n7563), .config_in(config_chain[10766:10764]), .config_rst(config_rst)); 
mux6 mux_3589 (.in({n14477_1, n14476_0, n14461_0/**/, n14460_0, n14367_0, n14366_0}), .out(n7564), .config_in(config_chain[10769:10767]), .config_rst(config_rst)); 
mux6 mux_3590 (.in({n10371_0, n10370_0, n10359_0, n10358_0, n10345_0, n10344_1}), .out(n7565), .config_in(config_chain[10772:10770]), .config_rst(config_rst)); 
mux6 mux_3591 (.in({n14183_0, n14182_0, n14167_0, n14166_0, n14135_0, n14134_0}), .out(n7566), .config_in(config_chain[10775:10773]), .config_rst(config_rst)); 
mux6 mux_3592 (.in({n10669_0, n10668_0, n10597_0, n10596_1, n10589_0, n10588_1}), .out(n7567), .config_in(config_chain[10778:10776]), .config_rst(config_rst)); 
mux6 mux_3593 (.in({n14485_1, n14484_0/**/, n14399_0, n14398_0, n14361_0, n14360_0}), .out(n7568), .config_in(config_chain[10781:10779]), .config_rst(config_rst)); 
mux6 mux_3594 (.in({n10393_0, n10392_0, n10387_0, n10386_0, n10379_0, n10378_0/**/}), .out(n7569), .config_in(config_chain[10784:10782]), .config_rst(config_rst)); 
mux6 mux_3595 (.in({n14213_1, n14212_0, n14205_1/**/, n14204_0, n14199_0, n14198_0}), .out(n7570), .config_in(config_chain[10787:10785]), .config_rst(config_rst)); 
mux6 mux_3596 (.in({n10631_0, n10630_0, n10617_0, n10616_0, n10605_0, n10604_1}), .out(n7571), .config_in(config_chain[10790:10788]), .config_rst(config_rst)); 
mux6 mux_3597 (.in({n14447_0, n14446_0, n14425_0, n14424_0, n14393_0/**/, n14392_0}), .out(n7572), .config_in(config_chain[10793:10791]), .config_rst(config_rst)); 
mux6 mux_3598 (.in({n10409_0, n10408_0/**/, n10339_0, n10338_1, n10331_0, n10330_1}), .out(n7573), .config_in(config_chain[10796:10794]), .config_rst(config_rst)); 
mux6 mux_3599 (.in({n14221_1, n14220_0, n14133_0, n14132_0, n14101_0, n14100_0}), .out(n7574), .config_in(config_chain[10799:10797]), .config_rst(config_rst)); 
mux6 mux_3600 (.in({n10655_0, n10654_0/**/, n10639_0, n10638_0, n10625_0, n10624_0}), .out(n7575), .config_in(config_chain[10802:10800]), .config_rst(config_rst)); 
mux6 mux_3601 (.in({n14471_1, n14470_0, n14463_0, n14462_0/**/, n14455_0, n14454_0}), .out(n7576), .config_in(config_chain[10805:10803]), .config_rst(config_rst)); 
mux6 mux_3602 (.in({n10361_0, n10360_0, n10353_0, n10352_0/**/, n10347_0, n10346_1}), .out(n7577), .config_in(config_chain[10808:10806]), .config_rst(config_rst)); 
mux6 mux_3603 (.in({n14185_0, n14184_0/**/, n14165_0, n14164_0, n14143_0, n14142_0}), .out(n7578), .config_in(config_chain[10811:10809]), .config_rst(config_rst)); 
mux6 mux_3604 (.in({n10671_0, n10670_0, n10663_0/**/, n10662_0, n10591_0, n10590_1}), .out(n7579), .config_in(config_chain[10814:10812]), .config_rst(config_rst)); 
mux6 mux_3605 (.in({n14487_2, n14486_0, n14407_0, n14406_0, n14375_0, n14374_0}), .out(n7580), .config_in(config_chain[10817:10815]), .config_rst(config_rst)); 
mux6 mux_3606 (.in({n10395_0, n10394_0/**/, n10381_0, n10380_0, n10263_0, n10262_2}), .out(n7581), .config_in(config_chain[10820:10818]), .config_rst(config_rst)); 
mux6 mux_3607 (.in({n14207_1/**/, n14206_0, n14193_0, n14192_0, n14175_0, n14174_0}), .out(n7582), .config_in(config_chain[10823:10821]), .config_rst(config_rst)); 
mux6 mux_3608 (.in({n10611_0, n10610_0, n10599_0/**/, n10598_1, n10521_0, n10520_2}), .out(n7583), .config_in(config_chain[10826:10824]), .config_rst(config_rst)); 
mux6 mux_3609 (.in({n14439_0, n14438_0, n14401_0, n14400_0, n14369_0, n14368_0}), .out(n7584), .config_in(config_chain[10829:10827]), .config_rst(config_rst)); 
mux6 mux_3610 (.in({n10403_0, n10402_0, n10333_0, n10332_1, n10265_0, n10264_2}), .out(n7585), .config_in(config_chain[10832:10830]), .config_rst(config_rst)); 
mux6 mux_3611 (.in({n14215_1, n14214_0, n14179_1, n14178_0, n14109_0, n14108_0}), .out(n7586), .config_in(config_chain[10835:10833]), .config_rst(config_rst)); 
mux6 mux_3612 (.in({n10641_0, n10640_0, n10633_0, n10632_0, n10523_0, n10522_2}), .out(n7587), .config_in(config_chain[10838:10836]), .config_rst(config_rst)); 
mux6 mux_3613 (.in({n14473_1, n14472_0, n14457_0, n14456_0, n14441_0/**/, n14440_0}), .out(n7588), .config_in(config_chain[10841:10839]), .config_rst(config_rst)); 
mux6 mux_3614 (.in({n10389_0, n10388_0, n10355_0, n10354_0, n10341_0, n10340_1}), .out(n7589), .config_in(config_chain[10844:10842]), .config_rst(config_rst)); 
mux6 mux_3615 (.in({n14201_2/**/, n14200_0, n14151_0, n14150_0, n14119_0, n14118_0}), .out(n7590), .config_in(config_chain[10847:10845]), .config_rst(config_rst)); 
mux6 mux_3616 (.in({n10665_0, n10664_0, n10657_0, n10656_0, n10525_0, n10524_2}), .out(n7591), .config_in(config_chain[10850:10848]), .config_rst(config_rst)); 
mux6 mux_3617 (.in({n14481_1, n14480_0/**/, n14443_0, n14442_0, n14383_0, n14382_0}), .out(n7592), .config_in(config_chain[10853:10851]), .config_rst(config_rst)); 
mux6 mux_3618 (.in({n10411_0, n10410_0, n10375_0, n10374_0, n10363_0, n10362_0}), .out(n7593), .config_in(config_chain[10856:10854]), .config_rst(config_rst)); 
mux6 mux_3619 (.in({n14223_2, n14222_0, n14195_0, n14194_0, n14187_0, n14186_0/**/}), .out(n7594), .config_in(config_chain[10859:10857]), .config_rst(config_rst)); 
mux6 mux_3620 (.in({n10627_0, n10626_0/**/, n10613_0, n10612_0, n10601_0, n10600_1}), .out(n7595), .config_in(config_chain[10862:10860]), .config_rst(config_rst)); 
mux6 mux_3621 (.in({n14465_2, n14464_0, n14415_0, n14414_0, n14377_0, n14376_0}), .out(n7596), .config_in(config_chain[10865:10863]), .config_rst(config_rst)); 
mux6 mux_3622 (.in({n10405_0, n10404_0, n10397_0, n10396_0, n10261_0, n10260_2}), .out(n7597), .config_in(config_chain[10868:10866]), .config_rst(config_rst)); 
mux6 mux_3623 (.in({n14217_1/**/, n14216_0, n14173_0, n14172_0, n14117_0, n14116_0}), .out(n7598), .config_in(config_chain[10871:10869]), .config_rst(config_rst)); 
mux6 mux_3624 (.in({n10927_0, n10926_0, n10869_0, n10868_0, n10853_0, n10852_1}), .out(n7645), .config_in(config_chain[10874:10872]), .config_rst(config_rst)); 
mux6 mux_3625 (.in({n14503_1, n14502_0, n14445_0, n14444_0/**/, n14377_0, n14376_1}), .out(n7646), .config_in(config_chain[10877:10875]), .config_rst(config_rst)); 
mux6 mux_3626 (.in({n10651_0, n10650_0, n10643_0, n10642_0, n10635_0, n10634_0}), .out(n7647), .config_in(config_chain[10880:10878]), .config_rst(config_rst)); 
mux6 mux_3627 (.in({n14233_1, n14232_0, n14225_1, n14224_0, n14217_0, n14216_0}), .out(n7648), .config_in(config_chain[10883:10881]), .config_rst(config_rst)); 
mux6 mux_3628 (.in({n10891_0, n10890_0, n10877_0, n10876_0, n10861_0, n10860_1}), .out(n7649), .config_in(config_chain[10886:10884]), .config_rst(config_rst)); 
mux6 mux_3629 (.in({n14467_0, n14466_0, n14461_0, n14460_0, n14453_0, n14452_0}), .out(n7650), .config_in(config_chain[10889:10887]), .config_rst(config_rst)); 
mux6 mux_3630 (.in({n10667_0, n10666_0, n10595_0, n10594_1, n10587_0, n10586_1}), .out(n7651), .config_in(config_chain[10892:10890]), .config_rst(config_rst)); 
mux6 mux_3631 (.in({n14241_1, n14240_0, n14181_0, n14180_0, n14127_0/**/, n14126_1}), .out(n7652), .config_in(config_chain[10895:10893]), .config_rst(config_rst)); 
mux6 mux_3632 (.in({n10913_0, n10912_0, n10907_0, n10906_0, n10899_0, n10898_0}), .out(n7653), .config_in(config_chain[10898:10896]), .config_rst(config_rst)); 
mux6 mux_3633 (.in({n14489_1, n14488_0, n14483_0, n14482_0, n14475_0, n14474_0/**/}), .out(n7654), .config_in(config_chain[10901:10899]), .config_rst(config_rst)); 
mux6 mux_3634 (.in({n10615_0, n10614_0, n10607_0, n10606_0, n10603_0, n10602_1}), .out(n7655), .config_in(config_chain[10904:10902]), .config_rst(config_rst)); 
mux6 mux_3635 (.in({n14203_0/**/, n14202_0, n14189_0, n14188_0, n14159_0, n14158_1}), .out(n7656), .config_in(config_chain[10907:10905]), .config_rst(config_rst)); 
mux6 mux_3636 (.in({n10929_0, n10928_0, n10921_0, n10920_0, n10847_0, n10846_1}), .out(n7657), .config_in(config_chain[10910:10908]), .config_rst(config_rst)); 
mux6 mux_3637 (.in({n14505_1, n14504_0, n14385_0, n14384_1/**/, n14353_0, n14352_1}), .out(n7658), .config_in(config_chain[10913:10911]), .config_rst(config_rst)); 
mux6 mux_3638 (.in({n10653_0, n10652_0, n10637_0/**/, n10636_0, n10623_0, n10622_0}), .out(n7659), .config_in(config_chain[10916:10914]), .config_rst(config_rst)); 
mux6 mux_3639 (.in({n14227_1, n14226_0, n14219_0, n14218_0, n14211_0, n14210_0}), .out(n7660), .config_in(config_chain[10919:10917]), .config_rst(config_rst)); 
mux6 mux_3640 (.in({n10879_0, n10878_0/**/, n10871_0, n10870_0, n10863_0, n10862_1}), .out(n7661), .config_in(config_chain[10922:10920]), .config_rst(config_rst)); 
mux6 mux_3641 (.in({n14469_0, n14468_0, n14455_0, n14454_0, n14417_0, n14416_1}), .out(n7662), .config_in(config_chain[10925:10923]), .config_rst(config_rst)); 
mux6 mux_3642 (.in({n10661_0, n10660_0, n10645_0, n10644_0, n10589_0, n10588_1}), .out(n7663), .config_in(config_chain[10928:10926]), .config_rst(config_rst)); 
mux6 mux_3643 (.in({n14243_1, n14242_0, n14235_1, n14234_0/**/, n14103_0, n14102_1}), .out(n7664), .config_in(config_chain[10931:10929]), .config_rst(config_rst)); 
mux6 mux_3644 (.in({n10901_0, n10900_0, n10893_0/**/, n10892_0, n10887_0, n10886_0}), .out(n7665), .config_in(config_chain[10934:10932]), .config_rst(config_rst)); 
mux6 mux_3645 (.in({n14491_1, n14490_0, n14477_0, n14476_0, n14463_0, n14462_0}), .out(n7666), .config_in(config_chain[10937:10935]), .config_rst(config_rst)); 
mux6 mux_3646 (.in({n10609_0, n10608_0, n10605_0, n10604_1, n10597_0, n10596_1}), .out(n7667), .config_in(config_chain[10940:10938]), .config_rst(config_rst)); 
mux6 mux_3647 (.in({n14191_0, n14190_0, n14183_0, n14182_0, n14167_0, n14166_1}), .out(n7668), .config_in(config_chain[10943:10941]), .config_rst(config_rst)); 
mux6 mux_3648 (.in({n10923_0, n10922_0, n10909_0, n10908_0, n10849_0, n10848_1}), .out(n7669), .config_in(config_chain[10946:10944]), .config_rst(config_rst)); 
mux6 mux_3649 (.in({n14507_1, n14506_0, n14499_1, n14498_0, n14361_0/**/, n14360_1}), .out(n7670), .config_in(config_chain[10949:10947]), .config_rst(config_rst)); 
mux6 mux_3650 (.in({n10639_0, n10638_0/**/, n10631_0, n10630_0, n10625_0, n10624_0}), .out(n7671), .config_in(config_chain[10952:10950]), .config_rst(config_rst)); 
mux6 mux_3651 (.in({n14213_0, n14212_0, n14205_0/**/, n14204_0, n14199_0, n14198_0}), .out(n7672), .config_in(config_chain[10955:10953]), .config_rst(config_rst)); 
mux6 mux_3652 (.in({n10931_0, n10930_0/**/, n10873_0, n10872_0, n10857_0, n10856_1}), .out(n7673), .config_in(config_chain[10958:10956]), .config_rst(config_rst)); 
mux6 mux_3653 (.in({n14449_0, n14448_0, n14425_0/**/, n14424_1, n14393_0, n14392_1}), .out(n7674), .config_in(config_chain[10961:10959]), .config_rst(config_rst)); 
mux6 mux_3654 (.in({n10663_0, n10662_0/**/, n10655_0, n10654_0, n10647_0, n10646_0}), .out(n7675), .config_in(config_chain[10964:10962]), .config_rst(config_rst)); 
mux6 mux_3655 (.in({n14237_1, n14236_0, n14221_0, n14220_0, n14111_0, n14110_1}), .out(n7676), .config_in(config_chain[10967:10965]), .config_rst(config_rst)); 
mux6 mux_3656 (.in({n10895_0, n10894_0, n10889_0, n10888_0, n10881_0, n10880_0/**/}), .out(n7677), .config_in(config_chain[10970:10968]), .config_rst(config_rst)); 
mux6 mux_3657 (.in({n14479_0, n14478_0, n14471_0, n14470_0, n14465_1, n14464_0}), .out(n7678), .config_in(config_chain[10973:10971]), .config_rst(config_rst)); 
mux6 mux_3658 (.in({n10671_0, n10670_0, n10611_0, n10610_0, n10599_0, n10598_1}), .out(n7679), .config_in(config_chain[10976:10974]), .config_rst(config_rst)); 
mux6 mux_3659 (.in({n14245_1, n14244_0, n14185_0, n14184_0, n14143_0, n14142_1}), .out(n7680), .config_in(config_chain[10979:10977]), .config_rst(config_rst)); 
mux6 mux_3660 (.in({n10917_0, n10916_0, n10911_0, n10910_0, n10903_0, n10902_0/**/}), .out(n7681), .config_in(config_chain[10982:10980]), .config_rst(config_rst)); 
mux6 mux_3661 (.in({n14501_1, n14500_0, n14493_1/**/, n14492_0, n14487_1, n14486_0}), .out(n7682), .config_in(config_chain[10985:10983]), .config_rst(config_rst)); 
mux6 mux_3662 (.in({n10633_0, n10632_0, n10619_0, n10618_0/**/, n10521_0, n10520_2}), .out(n7683), .config_in(config_chain[10988:10986]), .config_rst(config_rst)); 
mux6 mux_3663 (.in({n14207_0, n14206_0, n14193_0, n14192_0, n14177_0, n14176_1}), .out(n7684), .config_in(config_chain[10991:10989]), .config_rst(config_rst)); 
mux6 mux_3664 (.in({n10933_0, n10932_0, n10859_0, n10858_1, n10851_0, n10850_1}), .out(n7685), .config_in(config_chain[10994:10992]), .config_rst(config_rst)); 
mux6 mux_3665 (.in({n14509_1, n14508_0, n14451_0, n14450_0, n14401_0, n14400_1/**/}), .out(n7686), .config_in(config_chain[10997:10995]), .config_rst(config_rst)); 
mux6 mux_3666 (.in({n10657_0, n10656_0, n10641_0, n10640_0, n10525_0, n10524_2}), .out(n7687), .config_in(config_chain[11000:10998]), .config_rst(config_rst)); 
mux6 mux_3667 (.in({n14239_1/**/, n14238_0, n14231_1, n14230_0, n14179_0, n14178_1}), .out(n7688), .config_in(config_chain[11003:11001]), .config_rst(config_rst)); 
mux6 mux_3668 (.in({n10883_0, n10882_0, n10875_0, n10874_0, n10783_0, n10782_2}), .out(n7689), .config_in(config_chain[11006:11004]), .config_rst(config_rst)); 
mux6 mux_3669 (.in({n14473_0, n14472_0, n14459_0, n14458_0, n14441_0, n14440_1}), .out(n7690), .config_in(config_chain[11009:11007]), .config_rst(config_rst)); 
mux6 mux_3670 (.in({n10665_0, n10664_0, n10627_0, n10626_0, n10593_0/**/, n10592_1}), .out(n7691), .config_in(config_chain[11012:11010]), .config_rst(config_rst)); 
mux6 mux_3671 (.in({n14201_1, n14200_0, n14151_0, n14150_1, n14119_0, n14118_1/**/}), .out(n7692), .config_in(config_chain[11015:11013]), .config_rst(config_rst)); 
mux6 mux_3672 (.in({n10919_0, n10918_0/**/, n10905_0, n10904_0, n10785_0, n10784_2}), .out(n7693), .config_in(config_chain[11018:11016]), .config_rst(config_rst)); 
mux6 mux_3673 (.in({n14495_1, n14494_0, n14481_0, n14480_0/**/, n14433_1, n14432_1}), .out(n7694), .config_in(config_chain[11021:11019]), .config_rst(config_rst)); 
mux6 mux_3674 (.in({n10649_0, n10648_0, n10621_0, n10620_0, n10613_0, n10612_0}), .out(n7695), .config_in(config_chain[11024:11022]), .config_rst(config_rst)); 
mux6 mux_3675 (.in({n14223_1, n14222_0, n14209_0, n14208_0, n14195_0, n14194_0/**/}), .out(n7696), .config_in(config_chain[11027:11025]), .config_rst(config_rst)); 
mux6 mux_3676 (.in({n11177_0, n11176_0, n11161_0, n11160_0, n11147_0, n11146_0}), .out(n7743), .config_in(config_chain[11030:11028]), .config_rst(config_rst)); 
mux6 mux_3677 (.in({n14511_1, n14510_0, n14495_0, n14494_0, n14481_0, n14480_0}), .out(n7744), .config_in(config_chain[11033:11031]), .config_rst(config_rst)); 
mux6 mux_3678 (.in({n10869_0, n10868_0, n10861_0, n10860_1, n10853_0, n10852_1}), .out(n7745), .config_in(config_chain[11036:11034]), .config_rst(config_rst)); 
mux6 mux_3679 (.in({n14211_0, n14210_0/**/, n14203_0, n14202_0, n14195_0, n14194_1}), .out(n7746), .config_in(config_chain[11039:11037]), .config_rst(config_rst)); 
mux6 mux_3680 (.in({n11185_0, n11184_0, n11169_0, n11168_0, n11111_0, n11110_1}), .out(n7747), .config_in(config_chain[11042:11040]), .config_rst(config_rst)); 
mux6 mux_3681 (.in({n14527_1, n14526_0, n14519_1, n14518_0, n14445_0, n14444_1}), .out(n7748), .config_in(config_chain[11045:11043]), .config_rst(config_rst)); 
mux6 mux_3682 (.in({n10899_0, n10898_0, n10891_0, n10890_0, n10885_0, n10884_0}), .out(n7749), .config_in(config_chain[11048:11046]), .config_rst(config_rst)); 
mux6 mux_3683 (.in({n14247_1, n14246_0, n14233_0, n14232_0, n14219_0, n14218_0}), .out(n7750), .config_in(config_chain[11051:11049]), .config_rst(config_rst)); 
mux6 mux_3684 (.in({n11133_0, n11132_0, n11127_0, n11126_1, n11119_0, n11118_1}), .out(n7751), .config_in(config_chain[11054:11052]), .config_rst(config_rst)); 
mux6 mux_3685 (.in({n14467_0, n14466_0, n14461_0, n14460_1, n14453_0, n14452_1}), .out(n7752), .config_in(config_chain[11057:11055]), .config_rst(config_rst)); 
mux6 mux_3686 (.in({n10921_0, n10920_0, n10913_0, n10912_0, n10907_0, n10906_0}), .out(n7753), .config_in(config_chain[11060:11058]), .config_rst(config_rst)); 
mux6 mux_3687 (.in({n14255_1/**/, n14254_0, n14241_0, n14240_0, n14181_0, n14180_1}), .out(n7754), .config_in(config_chain[11063:11061]), .config_rst(config_rst)); 
mux6 mux_3688 (.in({n11155_0, n11154_0, n11149_0, n11148_0, n11141_0, n11140_0}), .out(n7755), .config_in(config_chain[11066:11064]), .config_rst(config_rst)); 
mux6 mux_3689 (.in({n14497_0, n14496_0, n14489_0, n14488_0, n14483_0/**/, n14482_0}), .out(n7756), .config_in(config_chain[11069:11067]), .config_rst(config_rst)); 
mux6 mux_3690 (.in({n10929_0, n10928_0, n10871_0, n10870_0/**/, n10855_0, n10854_1}), .out(n7757), .config_in(config_chain[11072:11070]), .config_rst(config_rst)); 
mux6 mux_3691 (.in({n14205_0, n14204_0, n14197_0/**/, n14196_1, n14189_0, n14188_1}), .out(n7758), .config_in(config_chain[11075:11073]), .config_rst(config_rst)); 
mux6 mux_3692 (.in({n11187_0, n11186_0, n11179_0, n11178_0, n11171_0, n11170_0/**/}), .out(n7759), .config_in(config_chain[11078:11076]), .config_rst(config_rst)); 
mux6 mux_3693 (.in({n14521_1, n14520_0, n14505_0, n14504_0, n14447_0, n14446_1}), .out(n7760), .config_in(config_chain[11081:11079]), .config_rst(config_rst)); 
mux6 mux_3694 (.in({n10893_0/**/, n10892_0, n10879_0, n10878_0, n10863_0, n10862_1}), .out(n7761), .config_in(config_chain[11084:11082]), .config_rst(config_rst)); 
mux6 mux_3695 (.in({n14227_0, n14226_0/**/, n14221_0, n14220_0, n14213_0, n14212_0}), .out(n7762), .config_in(config_chain[11087:11085]), .config_rst(config_rst)); 
mux6 mux_3696 (.in({n11195_0, n11194_0/**/, n11121_0, n11120_1, n11113_0, n11112_1}), .out(n7763), .config_in(config_chain[11090:11088]), .config_rst(config_rst)); 
mux6 mux_3697 (.in({n14529_1, n14528_0/**/, n14469_0, n14468_0, n14455_0, n14454_1}), .out(n7764), .config_in(config_chain[11093:11091]), .config_rst(config_rst)); 
mux6 mux_3698 (.in({n10915_0, n10914_0, n10909_0, n10908_0, n10901_0, n10900_0/**/}), .out(n7765), .config_in(config_chain[11096:11094]), .config_rst(config_rst)); 
mux6 mux_3699 (.in({n14257_1, n14256_0, n14249_1, n14248_0, n14243_0, n14242_0}), .out(n7766), .config_in(config_chain[11099:11097]), .config_rst(config_rst)); 
mux6 mux_3700 (.in({n11157_0, n11156_0, n11143_0, n11142_0, n11129_0, n11128_1}), .out(n7767), .config_in(config_chain[11102:11100]), .config_rst(config_rst)); 
mux6 mux_3701 (.in({n14491_0/**/, n14490_0, n14485_0, n14484_0, n14477_0, n14476_0}), .out(n7768), .config_in(config_chain[11105:11103]), .config_rst(config_rst)); 
mux6 mux_3702 (.in({n10931_0/**/, n10930_0, n10857_0, n10856_1, n10849_0, n10848_1}), .out(n7769), .config_in(config_chain[11108:11106]), .config_rst(config_rst)); 
mux6 mux_3703 (.in({n14265_1, n14264_0, n14191_0, n14190_1, n14183_0, n14182_1}), .out(n7770), .config_in(config_chain[11111:11109]), .config_rst(config_rst)); 
mux6 mux_3704 (.in({n11181_0, n11180_0, n11165_0, n11164_0, n11151_0, n11150_0}), .out(n7771), .config_in(config_chain[11114:11112]), .config_rst(config_rst)); 
mux6 mux_3705 (.in({n14515_1/**/, n14514_0, n14507_0, n14506_0, n14499_0, n14498_0}), .out(n7772), .config_in(config_chain[11117:11115]), .config_rst(config_rst)); 
mux6 mux_3706 (.in({n10881_0, n10880_0/**/, n10873_0, n10872_0, n10865_0, n10864_1}), .out(n7773), .config_in(config_chain[11120:11118]), .config_rst(config_rst)); 
mux6 mux_3707 (.in({n14229_0, n14228_0/**/, n14215_0, n14214_0, n14199_0, n14198_1}), .out(n7774), .config_in(config_chain[11123:11121]), .config_rst(config_rst)); 
mux6 mux_3708 (.in({n11189_0, n11188_0, n11115_0, n11114_1, n11109_0, n11108_1}), .out(n7775), .config_in(config_chain[11126:11124]), .config_rst(config_rst)); 
mux6 mux_3709 (.in({n14457_0, n14456_1, n14449_0/**/, n14448_1, n14433_1, n14432_1}), .out(n7776), .config_in(config_chain[11129:11127]), .config_rst(config_rst)); 
mux6 mux_3710 (.in({n10917_0, n10916_0, n10903_0, n10902_0, n10889_0, n10888_0}), .out(n7777), .config_in(config_chain[11132:11130]), .config_rst(config_rst)); 
mux6 mux_3711 (.in({n14251_1, n14250_0, n14237_0, n14236_0, n14223_1, n14222_0}), .out(n7778), .config_in(config_chain[11135:11133]), .config_rst(config_rst)); 
mux6 mux_3712 (.in({n11137_0/**/, n11136_0, n11131_0, n11130_1, n11123_0, n11122_1}), .out(n7779), .config_in(config_chain[11138:11136]), .config_rst(config_rst)); 
mux6 mux_3713 (.in({n14479_0, n14478_0, n14471_0, n14470_0, n14465_1, n14464_1}), .out(n7780), .config_in(config_chain[11141:11139]), .config_rst(config_rst)); 
mux6 mux_3714 (.in({n10925_0, n10924_0, n10911_0, n10910_0/**/, n10851_0, n10850_1}), .out(n7781), .config_in(config_chain[11144:11142]), .config_rst(config_rst)); 
mux6 mux_3715 (.in({n14267_1, n14266_0, n14259_1, n14258_0, n14185_0, n14184_1}), .out(n7782), .config_in(config_chain[11147:11145]), .config_rst(config_rst)); 
mux6 mux_3716 (.in({n11167_0, n11166_0, n11159_0, n11158_0, n11153_0, n11152_0}), .out(n7783), .config_in(config_chain[11150:11148]), .config_rst(config_rst)); 
mux6 mux_3717 (.in({n14517_1, n14516_0, n14501_0, n14500_0, n14487_1, n14486_0}), .out(n7784), .config_in(config_chain[11153:11151]), .config_rst(config_rst)); 
mux6 mux_3718 (.in({n10875_0, n10874_0, n10859_0/**/, n10858_1, n10783_0, n10782_2}), .out(n7785), .config_in(config_chain[11156:11154]), .config_rst(config_rst)); 
mux6 mux_3719 (.in({n14217_0, n14216_0, n14209_0, n14208_0, n14177_0/**/, n14176_1}), .out(n7786), .config_in(config_chain[11159:11157]), .config_rst(config_rst)); 
mux6 mux_3720 (.in({n11191_0, n11190_0, n11183_0, n11182_0, n11175_0, n11174_0}), .out(n7787), .config_in(config_chain[11162:11160]), .config_rst(config_rst)); 
mux6 mux_3721 (.in({n14525_1, n14524_0/**/, n14509_1, n14508_0, n14451_0, n14450_1}), .out(n7788), .config_in(config_chain[11165:11163]), .config_rst(config_rst)); 
mux6 mux_3722 (.in({n10897_0, n10896_0, n10883_0, n10882_0, n10785_0, n10784_2}), .out(n7789), .config_in(config_chain[11168:11166]), .config_rst(config_rst)); 
mux6 mux_3723 (.in({n14239_0, n14238_0, n14231_0, n14230_0, n14179_0, n14178_1}), .out(n7790), .config_in(config_chain[11171:11169]), .config_rst(config_rst)); 
mux6 mux_3724 (.in({n11197_0, n11196_0, n11139_0, n11138_0/**/, n11125_0, n11124_1}), .out(n7791), .config_in(config_chain[11174:11172]), .config_rst(config_rst)); 
mux6 mux_3725 (.in({n14473_0, n14472_0, n14459_0, n14458_1, n14443_0, n14442_1}), .out(n7792), .config_in(config_chain[11177:11175]), .config_rst(config_rst)); 
mux6 mux_3726 (.in({n10927_0, n10926_0, n10919_0/**/, n10918_0, n10867_0, n10866_1}), .out(n7793), .config_in(config_chain[11180:11178]), .config_rst(config_rst)); 
mux6 mux_3727 (.in({n14261_1, n14260_0, n14201_1, n14200_1/**/, n14187_0, n14186_1}), .out(n7794), .config_in(config_chain[11183:11181]), .config_rst(config_rst)); 
mux6 mux_3728 (.in({n11457_0, n11456_0, n11399_0, n11398_0, n11383_0, n11382_1}), .out(n7841), .config_in(config_chain[11186:11184]), .config_rst(config_rst)); 
mux6 mux_3729 (.in({n14547_1, n14546_0, n14489_0, n14488_0, n14473_0, n14472_1}), .out(n7842), .config_in(config_chain[11189:11187]), .config_rst(config_rst)); 
mux6 mux_3730 (.in({n11177_0, n11176_0, n11169_0, n11168_0, n11161_0, n11160_0/**/}), .out(n7843), .config_in(config_chain[11192:11190]), .config_rst(config_rst)); 
mux6 mux_3731 (.in({n14277_1, n14276_0, n14269_1, n14268_0, n14261_0, n14260_0}), .out(n7844), .config_in(config_chain[11195:11193]), .config_rst(config_rst)); 
mux6 mux_3732 (.in({n11421_0, n11420_0, n11407_0, n11406_0/**/, n11391_0, n11390_1}), .out(n7845), .config_in(config_chain[11198:11196]), .config_rst(config_rst)); 
mux6 mux_3733 (.in({n14511_0, n14510_0, n14505_0, n14504_0, n14497_0, n14496_0}), .out(n7846), .config_in(config_chain[11201:11199]), .config_rst(config_rst)); 
mux6 mux_3734 (.in({n11193_0, n11192_0, n11119_0, n11118_1, n11111_0, n11110_1}), .out(n7847), .config_in(config_chain[11204:11202]), .config_rst(config_rst)); 
mux6 mux_3735 (.in({n14285_1, n14284_0, n14225_0/**/, n14224_0, n14211_0, n14210_1}), .out(n7848), .config_in(config_chain[11207:11205]), .config_rst(config_rst)); 
mux6 mux_3736 (.in({n11443_0, n11442_0, n11437_0, n11436_0, n11429_0, n11428_0}), .out(n7849), .config_in(config_chain[11210:11208]), .config_rst(config_rst)); 
mux6 mux_3737 (.in({n14533_1, n14532_0, n14527_0, n14526_0, n14519_0, n14518_0}), .out(n7850), .config_in(config_chain[11213:11211]), .config_rst(config_rst)); 
mux6 mux_3738 (.in({n11141_0, n11140_0, n11133_0, n11132_0, n11127_0, n11126_1}), .out(n7851), .config_in(config_chain[11216:11214]), .config_rst(config_rst)); 
mux6 mux_3739 (.in({n14247_0, n14246_0, n14233_0, n14232_0, n14219_0, n14218_1}), .out(n7852), .config_in(config_chain[11219:11217]), .config_rst(config_rst)); 
mux6 mux_3740 (.in({n11459_0, n11458_0, n11451_0, n11450_0, n11377_0, n11376_1}), .out(n7853), .config_in(config_chain[11222:11220]), .config_rst(config_rst)); 
mux6 mux_3741 (.in({n14549_1, n14548_0, n14475_0, n14474_1, n14467_0/**/, n14466_1}), .out(n7854), .config_in(config_chain[11225:11223]), .config_rst(config_rst)); 
mux6 mux_3742 (.in({n11179_0, n11178_0/**/, n11163_0, n11162_0, n11149_0, n11148_0}), .out(n7855), .config_in(config_chain[11228:11226]), .config_rst(config_rst)); 
mux6 mux_3743 (.in({n14271_1, n14270_0, n14263_0, n14262_0, n14255_0, n14254_0/**/}), .out(n7856), .config_in(config_chain[11231:11229]), .config_rst(config_rst)); 
mux6 mux_3744 (.in({n11409_0, n11408_0, n11401_0, n11400_0, n11393_0/**/, n11392_1}), .out(n7857), .config_in(config_chain[11234:11232]), .config_rst(config_rst)); 
mux6 mux_3745 (.in({n14513_0, n14512_0/**/, n14499_0, n14498_0, n14483_0, n14482_1}), .out(n7858), .config_in(config_chain[11237:11235]), .config_rst(config_rst)); 
mux6 mux_3746 (.in({n11187_0, n11186_0, n11171_0, n11170_0/**/, n11113_0, n11112_1}), .out(n7859), .config_in(config_chain[11240:11238]), .config_rst(config_rst)); 
mux6 mux_3747 (.in({n14287_1, n14286_0, n14279_1, n14278_0, n14205_0, n14204_1}), .out(n7860), .config_in(config_chain[11243:11241]), .config_rst(config_rst)); 
mux6 mux_3748 (.in({n11431_0, n11430_0, n11423_0, n11422_0, n11417_0, n11416_0}), .out(n7861), .config_in(config_chain[11246:11244]), .config_rst(config_rst)); 
mux6 mux_3749 (.in({n14535_1, n14534_0, n14521_0, n14520_0, n14507_0, n14506_0/**/}), .out(n7862), .config_in(config_chain[11249:11247]), .config_rst(config_rst)); 
mux6 mux_3750 (.in({n11135_0, n11134_0, n11129_0, n11128_1, n11121_0, n11120_1}), .out(n7863), .config_in(config_chain[11252:11250]), .config_rst(config_rst)); 
mux6 mux_3751 (.in({n14235_0, n14234_0, n14227_0/**/, n14226_0, n14221_0, n14220_1}), .out(n7864), .config_in(config_chain[11255:11253]), .config_rst(config_rst)); 
mux6 mux_3752 (.in({n11453_0, n11452_0, n11439_0, n11438_0, n11379_0, n11378_1}), .out(n7865), .config_in(config_chain[11258:11256]), .config_rst(config_rst)); 
mux6 mux_3753 (.in({n14551_1, n14550_0, n14543_1/**/, n14542_0, n14469_0, n14468_1}), .out(n7866), .config_in(config_chain[11261:11259]), .config_rst(config_rst)); 
mux6 mux_3754 (.in({n11165_0, n11164_0/**/, n11157_0, n11156_0, n11151_0, n11150_0}), .out(n7867), .config_in(config_chain[11264:11262]), .config_rst(config_rst)); 
mux6 mux_3755 (.in({n14257_0, n14256_0/**/, n14249_0, n14248_0, n14243_0, n14242_0}), .out(n7868), .config_in(config_chain[11267:11265]), .config_rst(config_rst)); 
mux6 mux_3756 (.in({n11461_0, n11460_0, n11403_0, n11402_0, n11387_0, n11386_1/**/}), .out(n7869), .config_in(config_chain[11270:11268]), .config_rst(config_rst)); 
mux6 mux_3757 (.in({n14493_0, n14492_0, n14485_0, n14484_1/**/, n14477_0, n14476_1}), .out(n7870), .config_in(config_chain[11273:11271]), .config_rst(config_rst)); 
mux6 mux_3758 (.in({n11189_0, n11188_0, n11181_0, n11180_0, n11173_0, n11172_0}), .out(n7871), .config_in(config_chain[11276:11274]), .config_rst(config_rst)); 
mux6 mux_3759 (.in({n14281_1, n14280_0, n14265_0, n14264_0, n14207_0/**/, n14206_1}), .out(n7872), .config_in(config_chain[11279:11277]), .config_rst(config_rst)); 
mux6 mux_3760 (.in({n11463_0, n11462_0, n11425_0, n11424_0, n11411_0, n11410_0}), .out(n7873), .config_in(config_chain[11282:11280]), .config_rst(config_rst)); 
mux6 mux_3761 (.in({n14553_1, n14552_0, n14523_0, n14522_0, n14515_0, n14514_0/**/}), .out(n7874), .config_in(config_chain[11285:11283]), .config_rst(config_rst)); 
mux6 mux_3762 (.in({n11137_0, n11136_0, n11123_0/**/, n11122_1, n11109_0, n11108_1}), .out(n7875), .config_in(config_chain[11288:11286]), .config_rst(config_rst)); 
mux6 mux_3763 (.in({n14229_0, n14228_0, n14215_0, n14214_1, n14201_1, n14200_1}), .out(n7876), .config_in(config_chain[11291:11289]), .config_rst(config_rst)); 
mux6 mux_3764 (.in({n11447_0, n11446_0, n11433_0, n11432_0, n11353_0, n11352_1/**/}), .out(n7877), .config_in(config_chain[11294:11292]), .config_rst(config_rst)); 
mux6 mux_3765 (.in({n14545_1, n14544_0/**/, n14537_1, n14536_0, n14433_1, n14432_1}), .out(n7878), .config_in(config_chain[11297:11295]), .config_rst(config_rst)); 
mux6 mux_3766 (.in({n11159_0, n11158_0, n11145_0, n11144_0, n11131_0, n11130_1}), .out(n7879), .config_in(config_chain[11300:11298]), .config_rst(config_rst)); 
mux6 mux_3767 (.in({n14251_0, n14250_0, n14245_1, n14244_0, n14237_0, n14236_0/**/}), .out(n7880), .config_in(config_chain[11303:11301]), .config_rst(config_rst)); 
mux6 mux_3768 (.in({n11389_0, n11388_1/**/, n11381_0, n11380_1, n11375_0, n11374_1}), .out(n7881), .config_in(config_chain[11306:11304]), .config_rst(config_rst)); 
mux6 mux_3769 (.in({n14495_0, n14494_0, n14479_0, n14478_1/**/, n14465_1, n14464_1}), .out(n7882), .config_in(config_chain[11309:11307]), .config_rst(config_rst)); 
mux6 mux_3770 (.in({n11183_0, n11182_0/**/, n11175_0, n11174_0, n11167_0, n11166_0}), .out(n7883), .config_in(config_chain[11312:11310]), .config_rst(config_rst)); 
mux6 mux_3771 (.in({n14283_1, n14282_0, n14275_1, n14274_0/**/, n14267_1, n14266_0}), .out(n7884), .config_in(config_chain[11315:11313]), .config_rst(config_rst)); 
mux6 mux_3772 (.in({n11413_0, n11412_0, n11405_0, n11404_0, n11397_0, n11396_1}), .out(n7885), .config_in(config_chain[11318:11316]), .config_rst(config_rst)); 
mux6 mux_3773 (.in({n14517_0, n14516_0, n14503_0, n14502_0, n14487_1, n14486_1/**/}), .out(n7886), .config_in(config_chain[11321:11319]), .config_rst(config_rst)); 
mux6 mux_3774 (.in({n11197_0, n11196_0, n11191_0, n11190_0, n11117_0, n11116_1}), .out(n7887), .config_in(config_chain[11324:11322]), .config_rst(config_rst)); 
mux6 mux_3775 (.in({n14289_1, n14288_0, n14217_0, n14216_1, n14209_0/**/, n14208_1}), .out(n7888), .config_in(config_chain[11327:11325]), .config_rst(config_rst)); 
mux6 mux_3776 (.in({n11449_0, n11448_0, n11435_0, n11434_0, n11419_0, n11418_0}), .out(n7889), .config_in(config_chain[11330:11328]), .config_rst(config_rst)); 
mux6 mux_3777 (.in({n14539_1, n14538_0, n14531_1, n14530_0, n14525_0, n14524_0/**/}), .out(n7890), .config_in(config_chain[11333:11331]), .config_rst(config_rst)); 
mux6 mux_3778 (.in({n11147_0, n11146_0, n11139_0, n11138_0, n11047_0, n11046_2}), .out(n7891), .config_in(config_chain[11336:11334]), .config_rst(config_rst)); 
mux6 mux_3779 (.in({n14253_0, n14252_0, n14239_0, n14238_0, n14179_0, n14178_1}), .out(n7892), .config_in(config_chain[11339:11337]), .config_rst(config_rst)); 
mux6 mux_3780 (.in({n11709_0, n11708_0, n11693_0, n11692_0, n11679_0, n11678_0}), .out(n7939), .config_in(config_chain[11342:11340]), .config_rst(config_rst)); 
mux6 mux_3781 (.in({n14555_0, n14554_0, n14539_0, n14538_0, n14525_0, n14524_0}), .out(n7940), .config_in(config_chain[11345:11343]), .config_rst(config_rst)); 
mux6 mux_3782 (.in({n11399_0, n11398_0, n11391_0, n11390_1, n11383_0, n11382_1}), .out(n7941), .config_in(config_chain[11348:11346]), .config_rst(config_rst)); 
mux6 mux_3783 (.in({n14255_0, n14254_0, n14247_0, n14246_0, n14239_0/**/, n14238_1}), .out(n7942), .config_in(config_chain[11351:11349]), .config_rst(config_rst)); 
mux6 mux_3784 (.in({n11717_0, n11716_0, n11701_0, n11700_0, n11643_0, n11642_1/**/}), .out(n7943), .config_in(config_chain[11354:11352]), .config_rst(config_rst)); 
mux6 mux_3785 (.in({n14571_0, n14570_0, n14563_0, n14562_0, n14489_0, n14488_1}), .out(n7944), .config_in(config_chain[11357:11355]), .config_rst(config_rst)); 
mux6 mux_3786 (.in({n11429_0, n11428_0, n11421_0, n11420_0, n11415_0, n11414_0}), .out(n7945), .config_in(config_chain[11360:11358]), .config_rst(config_rst)); 
mux6 mux_3787 (.in({n14291_0, n14290_0, n14277_0, n14276_0, n14263_0, n14262_0}), .out(n7946), .config_in(config_chain[11363:11361]), .config_rst(config_rst)); 
mux6 mux_3788 (.in({n11665_0, n11664_0, n11659_0, n11658_1, n11651_0/**/, n11650_1}), .out(n7947), .config_in(config_chain[11366:11364]), .config_rst(config_rst)); 
mux6 mux_3789 (.in({n14511_0, n14510_0, n14505_0, n14504_1, n14497_0, n14496_1}), .out(n7948), .config_in(config_chain[11369:11367]), .config_rst(config_rst)); 
mux6 mux_3790 (.in({n11451_0, n11450_0, n11443_0, n11442_0, n11437_0, n11436_0}), .out(n7949), .config_in(config_chain[11372:11370]), .config_rst(config_rst)); 
mux6 mux_3791 (.in({n14299_0, n14298_0, n14285_0, n14284_0/**/, n14225_0, n14224_1}), .out(n7950), .config_in(config_chain[11375:11373]), .config_rst(config_rst)); 
mux6 mux_3792 (.in({n11687_0, n11686_0, n11681_0, n11680_0, n11673_0, n11672_0}), .out(n7951), .config_in(config_chain[11378:11376]), .config_rst(config_rst)); 
mux6 mux_3793 (.in({n14541_0, n14540_0/**/, n14533_0, n14532_0, n14527_0, n14526_0}), .out(n7952), .config_in(config_chain[11381:11379]), .config_rst(config_rst)); 
mux6 mux_3794 (.in({n11459_0, n11458_0, n11401_0, n11400_0, n11385_0, n11384_1}), .out(n7953), .config_in(config_chain[11384:11382]), .config_rst(config_rst)); 
mux6 mux_3795 (.in({n14249_0, n14248_0, n14241_0, n14240_1, n14233_0, n14232_1/**/}), .out(n7954), .config_in(config_chain[11387:11385]), .config_rst(config_rst)); 
mux6 mux_3796 (.in({n11719_0, n11718_0, n11711_0, n11710_0, n11703_0/**/, n11702_0}), .out(n7955), .config_in(config_chain[11390:11388]), .config_rst(config_rst)); 
mux6 mux_3797 (.in({n14565_0, n14564_0, n14549_0, n14548_0, n14491_0, n14490_1}), .out(n7956), .config_in(config_chain[11393:11391]), .config_rst(config_rst)); 
mux6 mux_3798 (.in({n11423_0, n11422_0, n11409_0, n11408_0/**/, n11393_0, n11392_1}), .out(n7957), .config_in(config_chain[11396:11394]), .config_rst(config_rst)); 
mux6 mux_3799 (.in({n14271_0, n14270_0, n14265_0/**/, n14264_0, n14257_0, n14256_0}), .out(n7958), .config_in(config_chain[11399:11397]), .config_rst(config_rst)); 
mux6 mux_3800 (.in({n11727_0, n11726_0/**/, n11653_0, n11652_1, n11645_0, n11644_1}), .out(n7959), .config_in(config_chain[11402:11400]), .config_rst(config_rst)); 
mux6 mux_3801 (.in({n14573_0, n14572_0, n14513_0, n14512_0, n14499_0, n14498_1}), .out(n7960), .config_in(config_chain[11405:11403]), .config_rst(config_rst)); 
mux6 mux_3802 (.in({n11445_0, n11444_0, n11439_0, n11438_0, n11431_0, n11430_0/**/}), .out(n7961), .config_in(config_chain[11408:11406]), .config_rst(config_rst)); 
mux6 mux_3803 (.in({n14301_0, n14300_0, n14293_0, n14292_0/**/, n14287_0, n14286_0}), .out(n7962), .config_in(config_chain[11411:11409]), .config_rst(config_rst)); 
mux6 mux_3804 (.in({n11689_0, n11688_0, n11675_0/**/, n11674_0, n11661_0, n11660_1}), .out(n7963), .config_in(config_chain[11414:11412]), .config_rst(config_rst)); 
mux6 mux_3805 (.in({n14535_0, n14534_0, n14529_0/**/, n14528_0, n14521_0, n14520_0}), .out(n7964), .config_in(config_chain[11417:11415]), .config_rst(config_rst)); 
mux6 mux_3806 (.in({n11461_0, n11460_0, n11387_0/**/, n11386_1, n11379_0, n11378_1}), .out(n7965), .config_in(config_chain[11420:11418]), .config_rst(config_rst)); 
mux6 mux_3807 (.in({n14309_0, n14308_0, n14235_0, n14234_1, n14227_0, n14226_1}), .out(n7966), .config_in(config_chain[11423:11421]), .config_rst(config_rst)); 
mux6 mux_3808 (.in({n11713_0, n11712_0, n11697_0, n11696_0/**/, n11683_0, n11682_0}), .out(n7967), .config_in(config_chain[11426:11424]), .config_rst(config_rst)); 
mux6 mux_3809 (.in({n14559_0/**/, n14558_0, n14551_0, n14550_0, n14543_0, n14542_0}), .out(n7968), .config_in(config_chain[11429:11427]), .config_rst(config_rst)); 
mux6 mux_3810 (.in({n11411_0, n11410_0, n11403_0, n11402_0, n11395_0/**/, n11394_1}), .out(n7969), .config_in(config_chain[11432:11430]), .config_rst(config_rst)); 
mux6 mux_3811 (.in({n14273_0, n14272_0, n14259_0, n14258_0, n14243_0, n14242_1}), .out(n7970), .config_in(config_chain[11435:11433]), .config_rst(config_rst)); 
mux6 mux_3812 (.in({n11721_0, n11720_0, n11685_0, n11684_0, n11647_0/**/, n11646_1}), .out(n7971), .config_in(config_chain[11438:11436]), .config_rst(config_rst)); 
mux6 mux_3813 (.in({n14531_0, n14530_0, n14501_0, n14500_1, n14493_0, n14492_1}), .out(n7972), .config_in(config_chain[11441:11439]), .config_rst(config_rst)); 
mux6 mux_3814 (.in({n11463_0, n11462_0, n11447_0, n11446_0, n11433_0, n11432_0/**/}), .out(n7973), .config_in(config_chain[11444:11442]), .config_rst(config_rst)); 
mux6 mux_3815 (.in({n14311_0, n14310_0, n14295_0, n14294_0/**/, n14281_0, n14280_0}), .out(n7974), .config_in(config_chain[11447:11445]), .config_rst(config_rst)); 
mux6 mux_3816 (.in({n11707_0, n11706_0, n11669_0, n11668_0, n11655_0, n11654_1/**/}), .out(n7975), .config_in(config_chain[11450:11448]), .config_rst(config_rst)); 
mux6 mux_3817 (.in({n14553_0, n14552_0, n14523_0, n14522_0/**/, n14515_0, n14514_0}), .out(n7976), .config_in(config_chain[11453:11451]), .config_rst(config_rst)); 
mux6 mux_3818 (.in({n11455_0, n11454_0/**/, n11381_0, n11380_1, n11353_0, n11352_1}), .out(n7977), .config_in(config_chain[11456:11454]), .config_rst(config_rst)); 
mux6 mux_3819 (.in({n14303_0, n14302_0, n14229_0, n14228_1, n14223_0, n14222_1}), .out(n7978), .config_in(config_chain[11459:11457]), .config_rst(config_rst)); 
mux6 mux_3820 (.in({n11699_0, n11698_0, n11691_0, n11690_0, n11597_0, n11596_2}), .out(n7979), .config_in(config_chain[11462:11460]), .config_rst(config_rst)); 
mux6 mux_3821 (.in({n14561_0, n14560_0/**/, n14545_0, n14544_0, n14433_0, n14432_2}), .out(n7980), .config_in(config_chain[11465:11463]), .config_rst(config_rst)); 
mux6 mux_3822 (.in({n11405_0, n11404_0, n11397_0, n11396_1/**/, n11389_0, n11388_1}), .out(n7981), .config_in(config_chain[11468:11466]), .config_rst(config_rst)); 
mux6 mux_3823 (.in({n14261_0, n14260_0, n14253_0, n14252_0/**/, n14245_0, n14244_1}), .out(n7982), .config_in(config_chain[11471:11469]), .config_rst(config_rst)); 
mux6 mux_3824 (.in({n11723_0, n11722_0, n11715_0, n11714_0/**/, n11619_0, n11618_1}), .out(n7983), .config_in(config_chain[11474:11472]), .config_rst(config_rst)); 
mux6 mux_3825 (.in({n14569_0, n14568_0, n14495_0/**/, n14494_1, n14465_0, n14464_1}), .out(n7984), .config_in(config_chain[11477:11475]), .config_rst(config_rst)); 
mux6 mux_3826 (.in({n11427_0, n11426_0, n11419_0, n11418_0, n11413_0/**/, n11412_0}), .out(n7985), .config_in(config_chain[11480:11478]), .config_rst(config_rst)); 
mux6 mux_3827 (.in({n14283_0, n14282_0/**/, n14275_0, n14274_0, n14267_0, n14266_0}), .out(n7986), .config_in(config_chain[11483:11481]), .config_rst(config_rst)); 
mux6 mux_3828 (.in({n11671_0, n11670_0, n11657_0, n11656_1, n11641_0, n11640_1}), .out(n7987), .config_in(config_chain[11486:11484]), .config_rst(config_rst)); 
mux6 mux_3829 (.in({n14517_0/**/, n14516_0, n14509_0, n14508_1, n14503_0, n14502_1}), .out(n7988), .config_in(config_chain[11489:11487]), .config_rst(config_rst)); 
mux6 mux_3830 (.in({n11457_0, n11456_0, n11449_0, n11448_0, n11441_0, n11440_0}), .out(n7989), .config_in(config_chain[11492:11490]), .config_rst(config_rst)); 
mux6 mux_3831 (.in({n14305_0, n14304_0, n14289_0, n14288_0, n14231_0, n14230_1}), .out(n7990), .config_in(config_chain[11495:11493]), .config_rst(config_rst)); 
mux6 mux_3832 (.in({n11985_0, n11984_0, n11929_0, n11928_0/**/, n11913_0, n11912_1}), .out(n8037), .config_in(config_chain[11498:11496]), .config_rst(config_rst)); 
mux6 mux_3833 (.in({n14589_0, n14588_0, n14533_0, n14532_0, n14517_0, n14516_1}), .out(n8038), .config_in(config_chain[11501:11499]), .config_rst(config_rst)); 
mux6 mux_3834 (.in({n11709_0, n11708_0, n11701_0, n11700_0/**/, n11693_0, n11692_0}), .out(n8039), .config_in(config_chain[11504:11502]), .config_rst(config_rst)); 
mux6 mux_3835 (.in({n14321_0, n14320_0, n14313_0, n14312_0, n14305_0, n14304_0}), .out(n8040), .config_in(config_chain[11507:11505]), .config_rst(config_rst)); 
mux6 mux_3836 (.in({n11951_0, n11950_0, n11937_0, n11936_0, n11921_0, n11920_1}), .out(n8041), .config_in(config_chain[11510:11508]), .config_rst(config_rst)); 
mux6 mux_3837 (.in({n14555_0, n14554_0, n14549_0/**/, n14548_0, n14541_0, n14540_0}), .out(n8042), .config_in(config_chain[11513:11511]), .config_rst(config_rst)); 
mux6 mux_3838 (.in({n11725_0, n11724_0, n11651_0, n11650_1, n11643_0, n11642_1}), .out(n8043), .config_in(config_chain[11516:11514]), .config_rst(config_rst)); 
mux6 mux_3839 (.in({n14329_0, n14328_0, n14269_0, n14268_0, n14255_0, n14254_1}), .out(n8044), .config_in(config_chain[11519:11517]), .config_rst(config_rst)); 
mux6 mux_3840 (.in({n11971_0, n11970_0, n11967_0, n11966_0, n11959_0, n11958_0}), .out(n8045), .config_in(config_chain[11522:11520]), .config_rst(config_rst)); 
mux6 mux_3841 (.in({n14575_0, n14574_0, n14571_0, n14570_0, n14563_0, n14562_0}), .out(n8046), .config_in(config_chain[11525:11523]), .config_rst(config_rst)); 
mux6 mux_3842 (.in({n11673_0, n11672_0, n11665_0, n11664_0, n11659_0, n11658_1}), .out(n8047), .config_in(config_chain[11528:11526]), .config_rst(config_rst)); 
mux6 mux_3843 (.in({n14291_0, n14290_0, n14277_0, n14276_0/**/, n14263_0, n14262_1}), .out(n8048), .config_in(config_chain[11531:11529]), .config_rst(config_rst)); 
mux6 mux_3844 (.in({n11987_0, n11986_0, n11979_0, n11978_0, n11907_0, n11906_1}), .out(n8049), .config_in(config_chain[11534:11532]), .config_rst(config_rst)); 
mux6 mux_3845 (.in({n14591_0, n14590_0, n14519_0/**/, n14518_1, n14511_0, n14510_1}), .out(n8050), .config_in(config_chain[11537:11535]), .config_rst(config_rst)); 
mux6 mux_3846 (.in({n11711_0, n11710_0, n11695_0, n11694_0, n11681_0, n11680_0}), .out(n8051), .config_in(config_chain[11540:11538]), .config_rst(config_rst)); 
mux6 mux_3847 (.in({n14315_0, n14314_0, n14307_0, n14306_0, n14299_0, n14298_0}), .out(n8052), .config_in(config_chain[11543:11541]), .config_rst(config_rst)); 
mux6 mux_3848 (.in({n11939_0, n11938_0, n11931_0, n11930_0, n11923_0, n11922_1/**/}), .out(n8053), .config_in(config_chain[11546:11544]), .config_rst(config_rst)); 
mux6 mux_3849 (.in({n14557_0, n14556_0, n14543_0, n14542_0, n14527_0, n14526_1}), .out(n8054), .config_in(config_chain[11549:11547]), .config_rst(config_rst)); 
mux6 mux_3850 (.in({n11719_0/**/, n11718_0, n11703_0, n11702_0, n11645_0, n11644_1}), .out(n8055), .config_in(config_chain[11552:11550]), .config_rst(config_rst)); 
mux6 mux_3851 (.in({n14331_0, n14330_0, n14323_0, n14322_0, n14249_0/**/, n14248_1}), .out(n8056), .config_in(config_chain[11555:11553]), .config_rst(config_rst)); 
mux6 mux_3852 (.in({n11961_0, n11960_0, n11953_0, n11952_0, n11947_0, n11946_0}), .out(n8057), .config_in(config_chain[11558:11556]), .config_rst(config_rst)); 
mux6 mux_3853 (.in({n14577_0, n14576_0/**/, n14565_0, n14564_0, n14551_0, n14550_0}), .out(n8058), .config_in(config_chain[11561:11559]), .config_rst(config_rst)); 
mux6 mux_3854 (.in({n11667_0, n11666_0, n11661_0, n11660_1, n11653_0, n11652_1}), .out(n8059), .config_in(config_chain[11564:11562]), .config_rst(config_rst)); 
mux6 mux_3855 (.in({n14279_0, n14278_0, n14271_0, n14270_0, n14265_0, n14264_1}), .out(n8060), .config_in(config_chain[11567:11565]), .config_rst(config_rst)); 
mux6 mux_3856 (.in({n11981_0, n11980_0, n11969_0, n11968_0, n11909_0/**/, n11908_1}), .out(n8061), .config_in(config_chain[11570:11568]), .config_rst(config_rst)); 
mux6 mux_3857 (.in({n14593_0, n14592_0/**/, n14585_0, n14584_0, n14513_0, n14512_1}), .out(n8062), .config_in(config_chain[11573:11571]), .config_rst(config_rst)); 
mux6 mux_3858 (.in({n11697_0, n11696_0, n11689_0, n11688_0, n11683_0, n11682_0/**/}), .out(n8063), .config_in(config_chain[11576:11574]), .config_rst(config_rst)); 
mux6 mux_3859 (.in({n14301_0, n14300_0, n14293_0, n14292_0, n14287_0, n14286_0/**/}), .out(n8064), .config_in(config_chain[11579:11577]), .config_rst(config_rst)); 
mux6 mux_3860 (.in({n11989_0, n11988_0, n11933_0, n11932_0, n11917_0, n11916_1}), .out(n8065), .config_in(config_chain[11582:11580]), .config_rst(config_rst)); 
mux6 mux_3861 (.in({n14537_0/**/, n14536_0, n14529_0, n14528_1, n14521_0, n14520_1}), .out(n8066), .config_in(config_chain[11585:11583]), .config_rst(config_rst)); 
mux6 mux_3862 (.in({n11721_0, n11720_0, n11713_0, n11712_0/**/, n11705_0, n11704_0}), .out(n8067), .config_in(config_chain[11588:11586]), .config_rst(config_rst)); 
mux6 mux_3863 (.in({n14325_0, n14324_0/**/, n14309_0, n14308_0, n14251_0, n14250_1}), .out(n8068), .config_in(config_chain[11591:11589]), .config_rst(config_rst)); 
mux6 mux_3864 (.in({n11955_0, n11954_0, n11941_0, n11940_0, n11905_0, n11904_1}), .out(n8069), .config_in(config_chain[11594:11592]), .config_rst(config_rst)); 
mux6 mux_3865 (.in({n14567_0, n14566_0, n14559_0, n14558_0, n14509_0, n14508_1}), .out(n8070), .config_in(config_chain[11597:11595]), .config_rst(config_rst)); 
mux6 mux_3866 (.in({n11685_0, n11684_0, n11669_0/**/, n11668_0, n11655_0, n11654_1}), .out(n8071), .config_in(config_chain[11600:11598]), .config_rst(config_rst)); 
mux6 mux_3867 (.in({n14289_0, n14288_0, n14273_0/**/, n14272_0, n14259_0, n14258_1}), .out(n8072), .config_in(config_chain[11603:11601]), .config_rst(config_rst)); 
mux6 mux_3868 (.in({n11975_0, n11974_0, n11963_0, n11962_0, n11927_0, n11926_1}), .out(n8073), .config_in(config_chain[11606:11604]), .config_rst(config_rst)); 
mux6 mux_3869 (.in({n14587_0, n14586_0, n14579_0, n14578_0/**/, n14531_0, n14530_1}), .out(n8074), .config_in(config_chain[11609:11607]), .config_rst(config_rst)); 
mux6 mux_3870 (.in({n11707_0, n11706_0, n11691_0, n11690_0, n11677_0, n11676_0}), .out(n8075), .config_in(config_chain[11612:11610]), .config_rst(config_rst)); 
mux6 mux_3871 (.in({n14295_0, n14294_0, n14281_0, n14280_0/**/, n14201_0, n14200_2}), .out(n8076), .config_in(config_chain[11615:11613]), .config_rst(config_rst)); 
mux6 mux_3872 (.in({n11949_0, n11948_0, n11919_0, n11918_1, n11911_0, n11910_1/**/}), .out(n8077), .config_in(config_chain[11618:11616]), .config_rst(config_rst)); 
mux6 mux_3873 (.in({n14553_0, n14552_0, n14539_0, n14538_0, n14523_0, n14522_1}), .out(n8078), .config_in(config_chain[11621:11619]), .config_rst(config_rst)); 
mux6 mux_3874 (.in({n11715_0, n11714_0, n11699_0, n11698_0, n11619_0, n11618_1}), .out(n8079), .config_in(config_chain[11624:11622]), .config_rst(config_rst)); 
mux6 mux_3875 (.in({n14327_0, n14326_0/**/, n14319_0, n14318_0, n14223_0, n14222_1}), .out(n8080), .config_in(config_chain[11627:11625]), .config_rst(config_rst)); 
mux6 mux_3876 (.in({n11943_0/**/, n11942_0, n11935_0, n11934_0, n11829_0, n11828_2}), .out(n8081), .config_in(config_chain[11630:11628]), .config_rst(config_rst)); 
mux6 mux_3877 (.in({n14561_0, n14560_0, n14547_0, n14546_0, n14433_0, n14432_2}), .out(n8082), .config_in(config_chain[11633:11631]), .config_rst(config_rst)); 
mux6 mux_3878 (.in({n11723_0, n11722_0, n11649_0, n11648_1/**/, n11641_0, n11640_1}), .out(n8083), .config_in(config_chain[11636:11634]), .config_rst(config_rst)); 
mux6 mux_3879 (.in({n14261_0, n14260_1/**/, n14253_0, n14252_1, n14245_0, n14244_1}), .out(n8084), .config_in(config_chain[11639:11637]), .config_rst(config_rst)); 
mux6 mux_3880 (.in({n11977_0, n11976_0/**/, n11965_0, n11964_0, n11861_0, n11860_2}), .out(n8085), .config_in(config_chain[11642:11640]), .config_rst(config_rst)); 
mux6 mux_3881 (.in({n14581_0, n14580_0, n14569_0, n14568_0/**/, n14487_0, n14486_1}), .out(n8086), .config_in(config_chain[11645:11643]), .config_rst(config_rst)); 
mux6 mux_3882 (.in({n11679_0, n11678_0, n11671_0, n11670_0/**/, n11663_0, n11662_1}), .out(n8087), .config_in(config_chain[11648:11646]), .config_rst(config_rst)); 
mux6 mux_3883 (.in({n14297_0, n14296_0, n14283_0, n14282_0/**/, n14267_0, n14266_1}), .out(n8088), .config_in(config_chain[11651:11649]), .config_rst(config_rst)); 
mux6 mux_3884 (.in({n12231_0, n12230_0, n12217_0, n12216_0, n12205_0, n12204_0}), .out(n8135), .config_in(config_chain[11654:11652]), .config_rst(config_rst)); 
mux6 mux_3885 (.in({n14595_0, n14594_0, n14581_0, n14580_0, n14569_0, n14568_0}), .out(n8136), .config_in(config_chain[11657:11655]), .config_rst(config_rst)); 
mux6 mux_3886 (.in({n11929_0, n11928_0, n11921_0, n11920_1, n11913_0, n11912_1}), .out(n8137), .config_in(config_chain[11660:11658]), .config_rst(config_rst)); 
mux6 mux_3887 (.in({n14299_0, n14298_0, n14291_0, n14290_0/**/, n14283_0, n14282_1}), .out(n8138), .config_in(config_chain[11663:11661]), .config_rst(config_rst)); 
mux6 mux_3888 (.in({n12239_0, n12238_0, n12225_0, n12224_0, n12169_0, n12168_1}), .out(n8139), .config_in(config_chain[11666:11664]), .config_rst(config_rst)); 
mux6 mux_3889 (.in({n14611_0, n14610_0, n14603_0, n14602_0, n14533_0, n14532_1}), .out(n8140), .config_in(config_chain[11669:11667]), .config_rst(config_rst)); 
mux6 mux_3890 (.in({n11959_0, n11958_0, n11951_0, n11950_0, n11945_0, n11944_0}), .out(n8141), .config_in(config_chain[11672:11670]), .config_rst(config_rst)); 
mux6 mux_3891 (.in({n14333_0, n14332_0/**/, n14321_0, n14320_0, n14307_0, n14306_0}), .out(n8142), .config_in(config_chain[11675:11673]), .config_rst(config_rst)); 
mux6 mux_3892 (.in({n12191_0, n12190_0, n12185_0, n12184_1, n12177_0, n12176_1}), .out(n8143), .config_in(config_chain[11678:11676]), .config_rst(config_rst)); 
mux6 mux_3893 (.in({n14555_0, n14554_0, n14549_0, n14548_1, n14541_0, n14540_1}), .out(n8144), .config_in(config_chain[11681:11679]), .config_rst(config_rst)); 
mux6 mux_3894 (.in({n11979_0, n11978_0, n11971_0, n11970_0, n11967_0, n11966_0}), .out(n8145), .config_in(config_chain[11684:11682]), .config_rst(config_rst)); 
mux6 mux_3895 (.in({n14341_0, n14340_0, n14329_0, n14328_0, n14269_0, n14268_1}), .out(n8146), .config_in(config_chain[11687:11685]), .config_rst(config_rst)); 
mux6 mux_3896 (.in({n12211_0, n12210_0, n12207_0, n12206_0, n12199_0, n12198_0}), .out(n8147), .config_in(config_chain[11690:11688]), .config_rst(config_rst)); 
mux6 mux_3897 (.in({n14583_0, n14582_0, n14575_0, n14574_0, n14571_0, n14570_0}), .out(n8148), .config_in(config_chain[11693:11691]), .config_rst(config_rst)); 
mux6 mux_3898 (.in({n11987_0, n11986_0/**/, n11931_0, n11930_0, n11915_0, n11914_1}), .out(n8149), .config_in(config_chain[11696:11694]), .config_rst(config_rst)); 
mux6 mux_3899 (.in({n14293_0, n14292_0, n14285_0, n14284_1, n14277_0, n14276_1/**/}), .out(n8150), .config_in(config_chain[11699:11697]), .config_rst(config_rst)); 
mux6 mux_3900 (.in({n12241_0, n12240_0, n12233_0, n12232_0, n12227_0, n12226_0}), .out(n8151), .config_in(config_chain[11702:11700]), .config_rst(config_rst)); 
mux6 mux_3901 (.in({n14605_0, n14604_0/**/, n14591_0, n14590_0, n14535_0, n14534_1}), .out(n8152), .config_in(config_chain[11705:11703]), .config_rst(config_rst)); 
mux6 mux_3902 (.in({n11953_0, n11952_0/**/, n11939_0, n11938_0, n11923_0, n11922_1}), .out(n8153), .config_in(config_chain[11708:11706]), .config_rst(config_rst)); 
mux6 mux_3903 (.in({n14315_0, n14314_0, n14309_0, n14308_0, n14301_0, n14300_0}), .out(n8154), .config_in(config_chain[11711:11709]), .config_rst(config_rst)); 
mux6 mux_3904 (.in({n12249_0, n12248_0, n12179_0, n12178_1/**/, n12171_0, n12170_1}), .out(n8155), .config_in(config_chain[11714:11712]), .config_rst(config_rst)); 
mux6 mux_3905 (.in({n14613_0, n14612_0, n14557_0, n14556_0, n14543_0, n14542_1}), .out(n8156), .config_in(config_chain[11717:11715]), .config_rst(config_rst)); 
mux6 mux_3906 (.in({n11973_0, n11972_0, n11969_0, n11968_0/**/, n11961_0, n11960_0}), .out(n8157), .config_in(config_chain[11720:11718]), .config_rst(config_rst)); 
mux6 mux_3907 (.in({n14343_0, n14342_0, n14335_0, n14334_0/**/, n14331_0, n14330_0}), .out(n8158), .config_in(config_chain[11723:11721]), .config_rst(config_rst)); 
mux6 mux_3908 (.in({n12213_0, n12212_0, n12201_0, n12200_0, n12187_0, n12186_1}), .out(n8159), .config_in(config_chain[11726:11724]), .config_rst(config_rst)); 
mux6 mux_3909 (.in({n14577_0, n14576_0, n14573_0, n14572_0, n14565_0, n14564_0}), .out(n8160), .config_in(config_chain[11729:11727]), .config_rst(config_rst)); 
mux6 mux_3910 (.in({n11989_0, n11988_0, n11917_0, n11916_1, n11909_0, n11908_1}), .out(n8161), .config_in(config_chain[11732:11730]), .config_rst(config_rst)); 
mux6 mux_3911 (.in({n14351_0, n14350_0, n14279_0, n14278_1, n14271_0, n14270_1}), .out(n8162), .config_in(config_chain[11735:11733]), .config_rst(config_rst)); 
mux6 mux_3912 (.in({n12235_0, n12234_0, n12221_0, n12220_0, n12209_0, n12208_0}), .out(n8163), .config_in(config_chain[11738:11736]), .config_rst(config_rst)); 
mux6 mux_3913 (.in({n14599_0, n14598_0, n14593_0, n14592_0, n14585_0, n14584_0}), .out(n8164), .config_in(config_chain[11741:11739]), .config_rst(config_rst)); 
mux6 mux_3914 (.in({n11941_0, n11940_0, n11933_0, n11932_0, n11925_0, n11924_1/**/}), .out(n8165), .config_in(config_chain[11744:11742]), .config_rst(config_rst)); 
mux6 mux_3915 (.in({n14317_0, n14316_0, n14303_0, n14302_0, n14287_0, n14286_1}), .out(n8166), .config_in(config_chain[11747:11745]), .config_rst(config_rst)); 
mux6 mux_3916 (.in({n12243_0, n12242_0, n12173_0, n12172_1, n12123_0, n12122_2}), .out(n8167), .config_in(config_chain[11750:11748]), .config_rst(config_rst)); 
mux6 mux_3917 (.in({n14545_0, n14544_1, n14537_0, n14536_1, n14487_0, n14486_2}), .out(n8168), .config_in(config_chain[11753:11751]), .config_rst(config_rst)); 
mux6 mux_3918 (.in({n11975_0, n11974_0, n11963_0, n11962_0, n11905_0, n11904_1}), .out(n8169), .config_in(config_chain[11756:11754]), .config_rst(config_rst)); 
mux6 mux_3919 (.in({n14337_0, n14336_0/**/, n14325_0, n14324_0, n14267_0, n14266_1}), .out(n8170), .config_in(config_chain[11759:11757]), .config_rst(config_rst)); 
mux6 mux_3920 (.in({n12195_0, n12194_0, n12181_0, n12180_1, n12145_0, n12144_1}), .out(n8171), .config_in(config_chain[11762:11760]), .config_rst(config_rst)); 
mux6 mux_3921 (.in({n14567_0, n14566_0, n14559_0, n14558_0/**/, n14509_0, n14508_1}), .out(n8172), .config_in(config_chain[11765:11763]), .config_rst(config_rst)); 
mux6 mux_3922 (.in({n11983_0, n11982_0, n11927_0, n11926_1, n11911_0, n11910_1/**/}), .out(n8173), .config_in(config_chain[11768:11766]), .config_rst(config_rst)); 
mux6 mux_3923 (.in({n14345_0, n14344_0/**/, n14311_0, n14310_0, n14273_0, n14272_1}), .out(n8174), .config_in(config_chain[11771:11769]), .config_rst(config_rst)); 
mux6 mux_3924 (.in({n12223_0, n12222_0, n12215_0, n12214_0/**/, n12167_0, n12166_1}), .out(n8175), .config_in(config_chain[11774:11772]), .config_rst(config_rst)); 
mux6 mux_3925 (.in({n14601_0, n14600_0/**/, n14587_0, n14586_0, n14531_0, n14530_1}), .out(n8176), .config_in(config_chain[11777:11775]), .config_rst(config_rst)); 
mux6 mux_3926 (.in({n11935_0, n11934_0, n11919_0, n11918_1/**/, n11829_0, n11828_2}), .out(n8177), .config_in(config_chain[11780:11778]), .config_rst(config_rst)); 
mux6 mux_3927 (.in({n14305_0, n14304_0, n14297_0, n14296_0, n14201_0, n14200_2}), .out(n8178), .config_in(config_chain[11783:11781]), .config_rst(config_rst)); 
mux6 mux_3928 (.in({n12245_0, n12244_0, n12237_0, n12236_0, n12189_0, n12188_1}), .out(n8179), .config_in(config_chain[11786:11784]), .config_rst(config_rst)); 
mux6 mux_3929 (.in({n14609_0, n14608_0, n14553_0, n14552_1, n14539_0, n14538_1/**/}), .out(n8180), .config_in(config_chain[11789:11787]), .config_rst(config_rst)); 
mux6 mux_3930 (.in({n11957_0, n11956_0, n11943_0, n11942_0, n11861_0, n11860_2}), .out(n8181), .config_in(config_chain[11792:11790]), .config_rst(config_rst)); 
mux6 mux_3931 (.in({n14327_0, n14326_0, n14319_0, n14318_0, n14223_0, n14222_2}), .out(n8182), .config_in(config_chain[11795:11793]), .config_rst(config_rst)); 
mux6 mux_3932 (.in({n12197_0, n12196_0, n12183_0, n12182_1, n12091_0, n12090_2}), .out(n8183), .config_in(config_chain[11798:11796]), .config_rst(config_rst)); 
mux6 mux_3933 (.in({n14561_0, n14560_0, n14547_0, n14546_1, n14465_0, n14464_2}), .out(n8184), .config_in(config_chain[11801:11799]), .config_rst(config_rst)); 
mux6 mux_3934 (.in({n11985_0, n11984_0, n11977_0, n11976_0, n11883_0, n11882_1}), .out(n8185), .config_in(config_chain[11804:11802]), .config_rst(config_rst)); 
mux6 mux_3935 (.in({n14347_0, n14346_0, n14275_0, n14274_1, n14245_0, n14244_1}), .out(n8186), .config_in(config_chain[11807:11805]), .config_rst(config_rst)); 
mux6 mux_3936 (.in({n12239_0, n12238_0, n12231_0, n12230_0, n12225_0, n12224_0}), .out(n8232), .config_in(config_chain[11810:11808]), .config_rst(config_rst)); 
mux6 mux_3937 (.in({n12199_0, n12198_0, n12191_0, n12190_0, n12185_0, n12184_1}), .out(n8235), .config_in(config_chain[11813:11811]), .config_rst(config_rst)); 
mux6 mux_3938 (.in({n12241_0, n12240_0, n12233_0, n12232_0, n12227_0, n12226_0}), .out(n8238), .config_in(config_chain[11816:11814]), .config_rst(config_rst)); 
mux6 mux_3939 (.in({n12201_0, n12200_0, n12193_0, n12192_0, n12187_0, n12186_1}), .out(n8241), .config_in(config_chain[11819:11817]), .config_rst(config_rst)); 
mux6 mux_3940 (.in({n12235_0, n12234_0, n12229_0, n12228_0, n12221_0, n12220_0}), .out(n8244), .config_in(config_chain[11822:11820]), .config_rst(config_rst)); 
mux6 mux_3941 (.in({n12195_0, n12194_0, n12181_0, n12180_1, n12145_0, n12144_1}), .out(n8247), .config_in(config_chain[11825:11823]), .config_rst(config_rst)); 
mux6 mux_3942 (.in({n12237_0, n12236_0, n12223_0, n12222_0, n12189_0, n12188_1}), .out(n8250), .config_in(config_chain[11828:11826]), .config_rst(config_rst)); 
mux6 mux_3943 (.in({n12197_0, n12196_0, n12183_0, n12182_1, n12093_0, n12092_2}), .out(n8253), .config_in(config_chain[11831:11829]), .config_rst(config_rst)); 
mux6 mux_3944 (.in({n9899_0, n9898_0, n9885_0, n9884_0, n9873_0, n9872_0}), .out(n8280), .config_in(config_chain[11834:11832]), .config_rst(config_rst)); 
mux6 mux_3945 (.in({n9915_0, n9914_0, n9847_0, n9846_1, n9839_0, n9838_1}), .out(n8283), .config_in(config_chain[11837:11835]), .config_rst(config_rst)); 
mux6 mux_3946 (.in({n9887_0, n9886_0, n9879_0, n9878_0, n9875_0, n9874_0}), .out(n8286), .config_in(config_chain[11840:11838]), .config_rst(config_rst)); 
mux6 mux_3947 (.in({n9917_0, n9916_0, n9849_0, n9848_1, n9841_0, n9840_1}), .out(n8289), .config_in(config_chain[11843:11841]), .config_rst(config_rst)); 
mux6 mux_3948 (.in({n9889_0, n9888_0, n9881_0, n9880_0, n9877_0, n9876_0}), .out(n8292), .config_in(config_chain[11846:11844]), .config_rst(config_rst)); 
mux6 mux_3949 (.in({n9911_0, n9910_0, n9843_0, n9842_1, n9755_0, n9754_2}), .out(n8295), .config_in(config_chain[11849:11847]), .config_rst(config_rst)); 
mux6 mux_3950 (.in({n9919_0, n9918_0, n9883_0, n9882_0, n9871_0, n9870_0}), .out(n8298), .config_in(config_chain[11852:11850]), .config_rst(config_rst)); 
mux6 mux_3951 (.in({n9913_0, n9912_0, n9845_0, n9844_1, n9751_0, n9750_2}), .out(n8301), .config_in(config_chain[11855:11853]), .config_rst(config_rst)); 
mux6 mux_3952 (.in({n10169_0, n10168_0, n10113_0, n10112_0, n10099_0, n10098_1}), .out(n8329), .config_in(config_chain[11858:11856]), .config_rst(config_rst)); 
mux6 mux_3953 (.in({n14673_1, n14672_0, n14643_0, n14642_0, n14621_0, n14620_0}), .out(n8330), .config_in(config_chain[11861:11859]), .config_rst(config_rst)); 
mux6 mux_3954 (.in({n9899_0, n9898_0, n9893_0, n9892_0, n9885_0, n9884_0}), .out(n8331), .config_in(config_chain[11864:11862]), .config_rst(config_rst)); 
mux6 mux_3955 (.in({n14415_0, n14414_0, n14385_1, n14384_0, n14353_1, n14352_0}), .out(n8332), .config_in(config_chain[11867:11865]), .config_rst(config_rst)); 
mux6 mux_3956 (.in({n10133_0, n10132_0, n10121_0, n10120_0, n10107_0, n10106_1}), .out(n8333), .config_in(config_chain[11870:11868]), .config_rst(config_rst)); 
mux6 mux_3957 (.in({n14685_0, n14684_0, n14653_0, n14652_0, n14615_0, n14614_0}), .out(n8334), .config_in(config_chain[11873:11871]), .config_rst(config_rst)); 
mux6 mux_3958 (.in({n9915_0, n9914_0, n9847_0, n9846_1, n9839_0, n9838_1}), .out(n8335), .config_in(config_chain[11876:11874]), .config_rst(config_rst)); 
mux6 mux_3959 (.in({n14417_1, n14416_0, n14387_0, n14386_0, n14357_0, n14356_0}), .out(n8336), .config_in(config_chain[11879:11877]), .config_rst(config_rst)); 
mux6 mux_3960 (.in({n10155_0, n10154_0, n10149_0, n10148_0, n10141_0, n10140_0}), .out(n8337), .config_in(config_chain[11882:11880]), .config_rst(config_rst)); 
mux6 mux_3961 (.in({n14679_0, n14678_0, n14647_0, n14646_0, n14617_1, n14616_0}), .out(n8338), .config_in(config_chain[11885:11883]), .config_rst(config_rst)); 
mux6 mux_3962 (.in({n9867_0, n9866_0, n9859_0, n9858_0, n9855_0, n9854_1}), .out(n8339), .config_in(config_chain[11888:11886]), .config_rst(config_rst)); 
mux6 mux_3963 (.in({n14419_0, n14418_0, n14389_0, n14388_0, n14359_0, n14358_0}), .out(n8340), .config_in(config_chain[11891:11889]), .config_rst(config_rst)); 
mux6 mux_3964 (.in({n10171_0, n10170_0, n10163_0, n10162_0, n10093_0, n10092_1}), .out(n8341), .config_in(config_chain[11894:11892]), .config_rst(config_rst)); 
mux6 mux_3965 (.in({n14681_1, n14680_0, n14651_0, n14650_0, n14619_0, n14618_0}), .out(n8342), .config_in(config_chain[11897:11895]), .config_rst(config_rst)); 
mux6 mux_3966 (.in({n9901_0, n9900_0, n9887_0, n9886_0, n9875_0, n9874_0}), .out(n8343), .config_in(config_chain[11900:11898]), .config_rst(config_rst)); 
mux6 mux_3967 (.in({n14423_0, n14422_0, n14391_0, n14390_0, n14361_1, n14360_0}), .out(n8344), .config_in(config_chain[11903:11901]), .config_rst(config_rst)); 
mux6 mux_3968 (.in({n10123_0, n10122_0, n10115_0, n10114_0, n10109_0, n10108_1}), .out(n8345), .config_in(config_chain[11906:11904]), .config_rst(config_rst)); 
mux6 mux_3969 (.in({n14683_0, n14682_0, n14661_0, n14660_0, n14623_0, n14622_0}), .out(n8346), .config_in(config_chain[11909:11907]), .config_rst(config_rst)); 
mux6 mux_3970 (.in({n9909_0, n9908_0, n9895_0, n9894_0, n9841_0, n9840_1}), .out(n8347), .config_in(config_chain[11912:11910]), .config_rst(config_rst)); 
mux6 mux_3971 (.in({n14425_1, n14424_0, n14393_1, n14392_0, n14363_0, n14362_0}), .out(n8348), .config_in(config_chain[11915:11913]), .config_rst(config_rst)); 
mux6 mux_3972 (.in({n10143_0, n10142_0, n10135_0, n10134_0, n10131_0, n10130_0}), .out(n8349), .config_in(config_chain[11918:11916]), .config_rst(config_rst)); 
mux6 mux_3973 (.in({n14693_0, n14692_0, n14655_0, n14654_0, n14625_1, n14624_0}), .out(n8350), .config_in(config_chain[11921:11919]), .config_rst(config_rst)); 
mux6 mux_3974 (.in({n9861_0, n9860_0, n9857_0, n9856_1, n9849_0, n9848_1}), .out(n8351), .config_in(config_chain[11924:11922]), .config_rst(config_rst)); 
mux6 mux_3975 (.in({n14427_0, n14426_0, n14397_0, n14396_0, n14365_0, n14364_0}), .out(n8352), .config_in(config_chain[11927:11925]), .config_rst(config_rst)); 
mux6 mux_3976 (.in({n10165_0, n10164_0, n10151_0, n10150_0, n10095_0, n10094_1}), .out(n8353), .config_in(config_chain[11930:11928]), .config_rst(config_rst)); 
mux6 mux_3977 (.in({n14689_1, n14688_0, n14657_1, n14656_0, n14627_0, n14626_0}), .out(n8354), .config_in(config_chain[11933:11931]), .config_rst(config_rst)); 
mux6 mux_3978 (.in({n9889_0, n9888_0, n9881_0, n9880_0, n9877_0, n9876_0}), .out(n8355), .config_in(config_chain[11936:11934]), .config_rst(config_rst)); 
mux6 mux_3979 (.in({n14429_0, n14428_0, n14399_0, n14398_0, n14367_0, n14366_0}), .out(n8356), .config_in(config_chain[11939:11937]), .config_rst(config_rst)); 
mux6 mux_3980 (.in({n10173_0, n10172_0, n10117_0, n10116_0, n10103_0, n10102_1}), .out(n8357), .config_in(config_chain[11942:11940]), .config_rst(config_rst)); 
mux6 mux_3981 (.in({n14691_0, n14690_0, n14659_0, n14658_0, n14637_0, n14636_0}), .out(n8358), .config_in(config_chain[11945:11943]), .config_rst(config_rst)); 
mux6 mux_3982 (.in({n9911_0, n9910_0, n9903_0, n9902_0, n9897_0, n9896_0}), .out(n8359), .config_in(config_chain[11948:11946]), .config_rst(config_rst)); 
mux6 mux_3983 (.in({n14431_0, n14430_0, n14401_1, n14400_0, n14371_0, n14370_0}), .out(n8360), .config_in(config_chain[11951:11949]), .config_rst(config_rst)); 
mux6 mux_3984 (.in({n10137_0, n10136_0, n10125_0, n10124_0, n10007_0, n10006_2}), .out(n8361), .config_in(config_chain[11954:11952]), .config_rst(config_rst)); 
mux6 mux_3985 (.in({n14701_0, n14700_0, n14663_0, n14662_0, n14631_0, n14630_0}), .out(n8362), .config_in(config_chain[11957:11955]), .config_rst(config_rst)); 
mux6 mux_3986 (.in({n9863_0, n9862_0, n9851_0, n9850_1, n9755_0, n9754_2}), .out(n8363), .config_in(config_chain[11960:11958]), .config_rst(config_rst)); 
mux6 mux_3987 (.in({n14441_1, n14440_0, n14403_0, n14402_0, n14373_0, n14372_0}), .out(n8364), .config_in(config_chain[11963:11961]), .config_rst(config_rst)); 
mux6 mux_3988 (.in({n10159_0, n10158_0, n10145_0, n10144_0, n10009_0, n10008_2}), .out(n8365), .config_in(config_chain[11966:11964]), .config_rst(config_rst)); 
mux6 mux_3989 (.in({n14703_0, n14702_0, n14665_1, n14664_0, n14633_1, n14632_0}), .out(n8366), .config_in(config_chain[11969:11967]), .config_rst(config_rst)); 
mux6 mux_3990 (.in({n9883_0, n9882_0, n9871_0, n9870_0, n9757_0, n9756_2}), .out(n8367), .config_in(config_chain[11972:11970]), .config_rst(config_rst)); 
mux6 mux_3991 (.in({n14433_2, n14432_0, n14405_0, n14404_0, n14375_0, n14374_0}), .out(n8368), .config_in(config_chain[11975:11973]), .config_rst(config_rst)); 
mux6 mux_3992 (.in({n10105_0, n10104_1, n10097_0, n10096_1, n10011_0, n10010_2}), .out(n8369), .config_in(config_chain[11978:11976]), .config_rst(config_rst)); 
mux6 mux_3993 (.in({n14705_1, n14704_0, n14667_0, n14666_0, n14645_0, n14644_0}), .out(n8370), .config_in(config_chain[11981:11979]), .config_rst(config_rst)); 
mux6 mux_3994 (.in({n9905_0, n9904_0, n9891_0, n9890_0, n9749_0, n9748_2}), .out(n8371), .config_in(config_chain[11984:11982]), .config_rst(config_rst)); 
mux6 mux_3995 (.in({n14435_0, n14434_0, n14409_1, n14408_0, n14377_1, n14376_0}), .out(n8372), .config_in(config_chain[11987:11985]), .config_rst(config_rst)); 
mux6 mux_3996 (.in({n10153_0, n10152_0, n10127_0, n10126_0, n10119_0, n10118_0}), .out(n8373), .config_in(config_chain[11990:11988]), .config_rst(config_rst)); 
mux6 mux_3997 (.in({n14695_2, n14694_0, n14677_0, n14676_0, n14639_0, n14638_0}), .out(n8374), .config_in(config_chain[11993:11991]), .config_rst(config_rst)); 
mux6 mux_3998 (.in({n9913_0, n9912_0, n9845_0, n9844_1, n9751_0, n9750_2}), .out(n8375), .config_in(config_chain[11996:11994]), .config_rst(config_rst)); 
mux6 mux_3999 (.in({n14437_0, n14436_0, n14411_0, n14410_0, n14379_0, n14378_0}), .out(n8376), .config_in(config_chain[11999:11997]), .config_rst(config_rst)); 
mux6 mux_4000 (.in({n10175_0, n10174_0, n10161_0, n10160_0, n10147_0, n10146_0}), .out(n8377), .config_in(config_chain[12002:12000]), .config_rst(config_rst)); 
mux6 mux_4001 (.in({n14699_0, n14698_0, n14671_0, n14670_0, n14641_1, n14640_0}), .out(n8378), .config_in(config_chain[12005:12003]), .config_rst(config_rst)); 
mux6 mux_4002 (.in({n9873_0, n9872_0, n9865_0, n9864_0, n9753_0, n9752_2}), .out(n8379), .config_in(config_chain[12008:12006]), .config_rst(config_rst)); 
mux6 mux_4003 (.in({n14439_0, n14438_0, n14413_0, n14412_0, n14383_0, n14382_0}), .out(n8380), .config_in(config_chain[12011:12009]), .config_rst(config_rst)); 
mux6 mux_4004 (.in({n10413_0, n10412_0, n10397_0, n10396_0, n10383_0, n10382_0}), .out(n8427), .config_in(config_chain[12014:12012]), .config_rst(config_rst)); 
mux6 mux_4005 (.in({n14707_1, n14706_0, n14671_0, n14670_0, n14641_0, n14640_0}), .out(n8428), .config_in(config_chain[12017:12015]), .config_rst(config_rst)); 
mux6 mux_4006 (.in({n10113_0, n10112_0, n10107_0, n10106_1, n10099_0, n10098_1}), .out(n8429), .config_in(config_chain[12020:12018]), .config_rst(config_rst)); 
mux6 mux_4007 (.in({n14413_0, n14412_0, n14391_0, n14390_0, n14359_0, n14358_0}), .out(n8430), .config_in(config_chain[12023:12021]), .config_rst(config_rst)); 
mux6 mux_4008 (.in({n10421_0, n10420_0, n10405_0, n10404_0, n10349_0, n10348_1}), .out(n8431), .config_in(config_chain[12026:12024]), .config_rst(config_rst)); 
mux6 mux_4009 (.in({n14723_1, n14722_0, n14715_1, n14714_0, n14621_0, n14620_0}), .out(n8432), .config_in(config_chain[12029:12027]), .config_rst(config_rst)); 
mux6 mux_4010 (.in({n10141_0, n10140_0, n10133_0, n10132_0, n10129_0, n10128_0}), .out(n8433), .config_in(config_chain[12032:12030]), .config_rst(config_rst)); 
mux6 mux_4011 (.in({n14445_1, n14444_0, n14423_0, n14422_0, n14385_0, n14384_0}), .out(n8434), .config_in(config_chain[12035:12033]), .config_rst(config_rst)); 
mux6 mux_4012 (.in({n10369_0, n10368_0, n10365_0, n10364_1, n10357_0, n10356_1}), .out(n8435), .config_in(config_chain[12038:12036]), .config_rst(config_rst)); 
mux6 mux_4013 (.in({n14685_0, n14684_0, n14653_0, n14652_0, n14615_0, n14614_0}), .out(n8436), .config_in(config_chain[12041:12039]), .config_rst(config_rst)); 
mux6 mux_4014 (.in({n10163_0, n10162_0, n10155_0, n10154_0, n10149_0, n10148_0}), .out(n8437), .config_in(config_chain[12044:12042]), .config_rst(config_rst)); 
mux6 mux_4015 (.in({n14453_1, n14452_0, n14417_0, n14416_0, n14357_0, n14356_0}), .out(n8438), .config_in(config_chain[12047:12045]), .config_rst(config_rst)); 
mux6 mux_4016 (.in({n10391_0, n10390_0, n10385_0, n10384_0, n10377_0, n10376_0}), .out(n8439), .config_in(config_chain[12050:12048]), .config_rst(config_rst)); 
mux6 mux_4017 (.in({n14679_0, n14678_0, n14649_0, n14648_0, n14617_0, n14616_0}), .out(n8440), .config_in(config_chain[12053:12051]), .config_rst(config_rst)); 
mux6 mux_4018 (.in({n10171_0, n10170_0, n10115_0, n10114_0, n10101_0, n10100_1}), .out(n8441), .config_in(config_chain[12056:12054]), .config_rst(config_rst)); 
mux6 mux_4019 (.in({n14421_0, n14420_0, n14389_0, n14388_0, n14367_0, n14366_0}), .out(n8442), .config_in(config_chain[12059:12057]), .config_rst(config_rst)); 
mux6 mux_4020 (.in({n10423_0, n10422_0, n10415_0, n10414_0, n10407_0, n10406_0}), .out(n8443), .config_in(config_chain[12062:12060]), .config_rst(config_rst)); 
mux6 mux_4021 (.in({n14717_1, n14716_0, n14681_0, n14680_0, n14629_0, n14628_0}), .out(n8444), .config_in(config_chain[12065:12063]), .config_rst(config_rst)); 
mux6 mux_4022 (.in({n10135_0, n10134_0, n10123_0, n10122_0, n10109_0, n10108_1}), .out(n8445), .config_in(config_chain[12068:12066]), .config_rst(config_rst)); 
mux6 mux_4023 (.in({n14431_0, n14430_0, n14399_0, n14398_0, n14361_0, n14360_0}), .out(n8446), .config_in(config_chain[12071:12069]), .config_rst(config_rst)); 
mux6 mux_4024 (.in({n10431_0, n10430_0, n10359_0, n10358_1, n10351_0, n10350_1}), .out(n8447), .config_in(config_chain[12074:12072]), .config_rst(config_rst)); 
mux6 mux_4025 (.in({n14725_1, n14724_0, n14661_0, n14660_0, n14623_0, n14622_0}), .out(n8448), .config_in(config_chain[12077:12075]), .config_rst(config_rst)); 
mux6 mux_4026 (.in({n10157_0, n10156_0, n10151_0, n10150_0, n10143_0, n10142_0}), .out(n8449), .config_in(config_chain[12080:12078]), .config_rst(config_rst)); 
mux6 mux_4027 (.in({n14455_1, n14454_0, n14447_1, n14446_0, n14425_0, n14424_0}), .out(n8450), .config_in(config_chain[12083:12081]), .config_rst(config_rst)); 
mux6 mux_4028 (.in({n10393_0, n10392_0, n10379_0, n10378_0, n10367_0, n10366_1}), .out(n8451), .config_in(config_chain[12086:12084]), .config_rst(config_rst)); 
mux6 mux_4029 (.in({n14687_0, n14686_0, n14655_0, n14654_0, n14625_0, n14624_0}), .out(n8452), .config_in(config_chain[12089:12087]), .config_rst(config_rst)); 
mux6 mux_4030 (.in({n10173_0, n10172_0, n10103_0, n10102_1, n10095_0, n10094_1}), .out(n8453), .config_in(config_chain[12092:12090]), .config_rst(config_rst)); 
mux6 mux_4031 (.in({n14463_1, n14462_0, n14397_0, n14396_0, n14365_0, n14364_0}), .out(n8454), .config_in(config_chain[12095:12093]), .config_rst(config_rst)); 
mux6 mux_4032 (.in({n10417_0, n10416_0, n10401_0, n10400_0, n10387_0, n10386_0}), .out(n8455), .config_in(config_chain[12098:12096]), .config_rst(config_rst)); 
mux6 mux_4033 (.in({n14711_1, n14710_0, n14689_0, n14688_0, n14657_0, n14656_0}), .out(n8456), .config_in(config_chain[12101:12099]), .config_rst(config_rst)); 
mux6 mux_4034 (.in({n10125_0, n10124_0, n10117_0, n10116_0, n10111_0, n10110_1}), .out(n8457), .config_in(config_chain[12104:12102]), .config_rst(config_rst)); 
mux6 mux_4035 (.in({n14429_0, n14428_0, n14407_0, n14406_0, n14369_0, n14368_0}), .out(n8458), .config_in(config_chain[12107:12105]), .config_rst(config_rst)); 
mux6 mux_4036 (.in({n10433_0, n10432_0, n10425_0, n10424_0, n10353_0, n10352_1}), .out(n8459), .config_in(config_chain[12110:12108]), .config_rst(config_rst)); 
mux6 mux_4037 (.in({n14727_2, n14726_0, n14669_0, n14668_0, n14637_0, n14636_0}), .out(n8460), .config_in(config_chain[12113:12111]), .config_rst(config_rst)); 
mux6 mux_4038 (.in({n10159_0, n10158_0, n10145_0, n10144_0, n10007_0, n10006_2}), .out(n8461), .config_in(config_chain[12116:12114]), .config_rst(config_rst)); 
mux6 mux_4039 (.in({n14449_1, n14448_0, n14439_0, n14438_0, n14401_0, n14400_0}), .out(n8462), .config_in(config_chain[12119:12117]), .config_rst(config_rst)); 
mux6 mux_4040 (.in({n10373_0, n10372_0, n10361_0, n10360_1, n10263_0, n10262_2}), .out(n8463), .config_in(config_chain[12122:12120]), .config_rst(config_rst)); 
mux6 mux_4041 (.in({n14701_0, n14700_0, n14663_0, n14662_0, n14631_0, n14630_0}), .out(n8464), .config_in(config_chain[12125:12123]), .config_rst(config_rst)); 
mux6 mux_4042 (.in({n10167_0, n10166_0, n10097_0, n10096_1, n10009_0, n10008_2}), .out(n8465), .config_in(config_chain[12128:12126]), .config_rst(config_rst)); 
mux6 mux_4043 (.in({n14457_1, n14456_0, n14443_1, n14442_0, n14373_0, n14372_0}), .out(n8466), .config_in(config_chain[12131:12129]), .config_rst(config_rst)); 
mux6 mux_4044 (.in({n10403_0, n10402_0, n10395_0, n10394_0, n10265_0, n10264_2}), .out(n8467), .config_in(config_chain[12134:12132]), .config_rst(config_rst)); 
mux6 mux_4045 (.in({n14713_1, n14712_0, n14703_0, n14702_0, n14665_0, n14664_0}), .out(n8468), .config_in(config_chain[12137:12135]), .config_rst(config_rst)); 
mux6 mux_4046 (.in({n10153_0, n10152_0, n10119_0, n10118_0, n10105_0, n10104_1}), .out(n8469), .config_in(config_chain[12140:12138]), .config_rst(config_rst)); 
mux6 mux_4047 (.in({n14433_2, n14432_0, n14415_0, n14414_0, n14383_0, n14382_0}), .out(n8470), .config_in(config_chain[12143:12141]), .config_rst(config_rst)); 
mux6 mux_4048 (.in({n10427_0, n10426_0, n10419_0, n10418_0, n10267_0, n10266_2}), .out(n8471), .config_in(config_chain[12146:12144]), .config_rst(config_rst)); 
mux6 mux_4049 (.in({n14721_1, n14720_0, n14705_0, n14704_0, n14645_0, n14644_0}), .out(n8472), .config_in(config_chain[12149:12147]), .config_rst(config_rst)); 
mux6 mux_4050 (.in({n10175_0, n10174_0, n10139_0, n10138_0, n10127_0, n10126_0}), .out(n8473), .config_in(config_chain[12152:12150]), .config_rst(config_rst)); 
mux6 mux_4051 (.in({n14465_2, n14464_0, n14409_0, n14408_0, n14377_0, n14376_0}), .out(n8474), .config_in(config_chain[12155:12153]), .config_rst(config_rst)); 
mux6 mux_4052 (.in({n10389_0, n10388_0, n10375_0, n10374_0, n10363_0, n10362_1}), .out(n8475), .config_in(config_chain[12158:12156]), .config_rst(config_rst)); 
mux6 mux_4053 (.in({n14697_2, n14696_0, n14677_0, n14676_0, n14639_0, n14638_0}), .out(n8476), .config_in(config_chain[12161:12159]), .config_rst(config_rst)); 
mux6 mux_4054 (.in({n10169_0, n10168_0, n10161_0, n10160_0, n10005_0, n10004_2}), .out(n8477), .config_in(config_chain[12164:12162]), .config_rst(config_rst)); 
mux6 mux_4055 (.in({n14459_1, n14458_0, n14437_0, n14436_0, n14381_0, n14380_0}), .out(n8478), .config_in(config_chain[12167:12165]), .config_rst(config_rst)); 
mux6 mux_4056 (.in({n10687_0, n10686_0, n10629_0, n10628_0, n10613_0, n10612_1}), .out(n8525), .config_in(config_chain[12170:12168]), .config_rst(config_rst)); 
mux6 mux_4057 (.in({n14743_1, n14742_0, n14639_0, n14638_0, n14617_0, n14616_0}), .out(n8526), .config_in(config_chain[12173:12171]), .config_rst(config_rst)); 
mux6 mux_4058 (.in({n10413_0, n10412_0, n10405_0, n10404_0/**/, n10397_0, n10396_0}), .out(n8527), .config_in(config_chain[12176:12174]), .config_rst(config_rst)); 
mux6 mux_4059 (.in({n14475_1, n14474_0, n14467_1, n14466_0, n14459_0, n14458_0}), .out(n8528), .config_in(config_chain[12179:12177]), .config_rst(config_rst)); 
mux6 mux_4060 (.in({n10651_0, n10650_0, n10637_0, n10636_0, n10621_0, n10620_1}), .out(n8529), .config_in(config_chain[12182:12180]), .config_rst(config_rst)); 
mux6 mux_4061 (.in({n14707_0, n14706_0, n14681_0, n14680_0, n14649_0, n14648_0}), .out(n8530), .config_in(config_chain[12185:12183]), .config_rst(config_rst)); 
mux6 mux_4062 (.in({n10429_0, n10428_0, n10357_0, n10356_1, n10349_0, n10348_1}), .out(n8531), .config_in(config_chain[12188:12186]), .config_rst(config_rst)); 
mux6 mux_4063 (.in({n14483_1, n14482_0, n14391_0, n14390_0, n14353_0, n14352_0}), .out(n8532), .config_in(config_chain[12191:12189]), .config_rst(config_rst)); 
mux6 mux_4064 (.in({n10673_0, n10672_0, n10667_0, n10666_0, n10659_0, n10658_0/**/}), .out(n8533), .config_in(config_chain[12194:12192]), .config_rst(config_rst)); 
mux6 mux_4065 (.in({n14729_1, n14728_0, n14723_0, n14722_0, n14715_0, n14714_0}), .out(n8534), .config_in(config_chain[12197:12195]), .config_rst(config_rst)); 
mux6 mux_4066 (.in({n10377_0, n10376_0, n10369_0, n10368_0, n10365_0, n10364_1}), .out(n8535), .config_in(config_chain[12200:12198]), .config_rst(config_rst)); 
mux6 mux_4067 (.in({n14445_0, n14444_0, n14423_0, n14422_0, n14385_0, n14384_0}), .out(n8536), .config_in(config_chain[12203:12201]), .config_rst(config_rst)); 
mux6 mux_4068 (.in({n10689_0, n10688_0, n10681_0, n10680_0, n10607_0, n10606_1}), .out(n8537), .config_in(config_chain[12206:12204]), .config_rst(config_rst)); 
mux6 mux_4069 (.in({n14745_1, n14744_0, n14647_0/**/, n14646_0, n14615_0, n14614_0}), .out(n8538), .config_in(config_chain[12209:12207]), .config_rst(config_rst)); 
mux6 mux_4070 (.in({n10415_0, n10414_0/**/, n10399_0, n10398_0, n10385_0, n10384_0}), .out(n8539), .config_in(config_chain[12212:12210]), .config_rst(config_rst)); 
mux6 mux_4071 (.in({n14469_1, n14468_0, n14461_0, n14460_0, n14453_0, n14452_0}), .out(n8540), .config_in(config_chain[12215:12213]), .config_rst(config_rst)); 
mux6 mux_4072 (.in({n10639_0, n10638_0, n10631_0, n10630_0, n10623_0, n10622_1/**/}), .out(n8541), .config_in(config_chain[12218:12216]), .config_rst(config_rst)); 
mux6 mux_4073 (.in({n14709_0/**/, n14708_0, n14679_0, n14678_0, n14657_0, n14656_0}), .out(n8542), .config_in(config_chain[12221:12219]), .config_rst(config_rst)); 
mux6 mux_4074 (.in({n10423_0, n10422_0, n10407_0, n10406_0, n10351_0, n10350_1}), .out(n8543), .config_in(config_chain[12224:12222]), .config_rst(config_rst)); 
mux6 mux_4075 (.in({n14485_1, n14484_0, n14477_1, n14476_0, n14367_0, n14366_0/**/}), .out(n8544), .config_in(config_chain[12227:12225]), .config_rst(config_rst)); 
mux6 mux_4076 (.in({n10661_0, n10660_0, n10653_0, n10652_0/**/, n10647_0, n10646_0}), .out(n8545), .config_in(config_chain[12230:12228]), .config_rst(config_rst)); 
mux6 mux_4077 (.in({n14731_1, n14730_0, n14717_0, n14716_0, n14689_0, n14688_0}), .out(n8546), .config_in(config_chain[12233:12231]), .config_rst(config_rst)); 
mux6 mux_4078 (.in({n10371_0, n10370_0, n10367_0, n10366_1, n10359_0, n10358_1/**/}), .out(n8547), .config_in(config_chain[12236:12234]), .config_rst(config_rst)); 
mux6 mux_4079 (.in({n14431_0, n14430_0, n14393_0, n14392_0, n14361_0, n14360_0}), .out(n8548), .config_in(config_chain[12239:12237]), .config_rst(config_rst)); 
mux6 mux_4080 (.in({n10683_0, n10682_0/**/, n10669_0, n10668_0, n10609_0, n10608_1}), .out(n8549), .config_in(config_chain[12242:12240]), .config_rst(config_rst)); 
mux6 mux_4081 (.in({n14747_1, n14746_0, n14739_1, n14738_0, n14623_0, n14622_0}), .out(n8550), .config_in(config_chain[12245:12243]), .config_rst(config_rst)); 
mux6 mux_4082 (.in({n10401_0/**/, n10400_0, n10393_0, n10392_0, n10387_0, n10386_0}), .out(n8551), .config_in(config_chain[12248:12246]), .config_rst(config_rst)); 
mux6 mux_4083 (.in({n14455_0/**/, n14454_0, n14447_0, n14446_0, n14425_0, n14424_0}), .out(n8552), .config_in(config_chain[12251:12249]), .config_rst(config_rst)); 
mux6 mux_4084 (.in({n10691_0, n10690_0, n10633_0, n10632_0/**/, n10617_0, n10616_1}), .out(n8553), .config_in(config_chain[12254:12252]), .config_rst(config_rst)); 
mux6 mux_4085 (.in({n14687_0, n14686_0, n14655_0, n14654_0, n14633_0, n14632_0}), .out(n8554), .config_in(config_chain[12257:12255]), .config_rst(config_rst)); 
mux6 mux_4086 (.in({n10425_0, n10424_0/**/, n10417_0, n10416_0, n10409_0, n10408_0}), .out(n8555), .config_in(config_chain[12260:12258]), .config_rst(config_rst)); 
mux6 mux_4087 (.in({n14479_1/**/, n14478_0, n14463_0, n14462_0, n14375_0, n14374_0}), .out(n8556), .config_in(config_chain[12263:12261]), .config_rst(config_rst)); 
mux6 mux_4088 (.in({n10655_0, n10654_0, n10649_0, n10648_0, n10641_0, n10640_0}), .out(n8557), .config_in(config_chain[12266:12264]), .config_rst(config_rst)); 
mux6 mux_4089 (.in({n14719_0/**/, n14718_0, n14711_0, n14710_0, n14697_2, n14696_0}), .out(n8558), .config_in(config_chain[12269:12267]), .config_rst(config_rst)); 
mux6 mux_4090 (.in({n10433_0, n10432_0/**/, n10373_0, n10372_0, n10361_0, n10360_1}), .out(n8559), .config_in(config_chain[12272:12270]), .config_rst(config_rst)); 
mux6 mux_4091 (.in({n14487_2, n14486_0, n14407_0/**/, n14406_0, n14369_0, n14368_0}), .out(n8560), .config_in(config_chain[12275:12273]), .config_rst(config_rst)); 
mux6 mux_4092 (.in({n10677_0, n10676_0, n10671_0, n10670_0, n10663_0, n10662_0}), .out(n8561), .config_in(config_chain[12278:12276]), .config_rst(config_rst)); 
mux6 mux_4093 (.in({n14741_1, n14740_0, n14733_1/**/, n14732_0, n14727_2, n14726_0}), .out(n8562), .config_in(config_chain[12281:12279]), .config_rst(config_rst)); 
mux6 mux_4094 (.in({n10395_0, n10394_0, n10381_0, n10380_0/**/, n10263_0, n10262_2}), .out(n8563), .config_in(config_chain[12284:12282]), .config_rst(config_rst)); 
mux6 mux_4095 (.in({n14449_0, n14448_0, n14441_0, n14440_0, n14401_0, n14400_0/**/}), .out(n8564), .config_in(config_chain[12287:12285]), .config_rst(config_rst)); 
mux6 mux_4096 (.in({n10693_0/**/, n10692_0, n10619_0, n10618_1, n10611_0, n10610_1}), .out(n8565), .config_in(config_chain[12290:12288]), .config_rst(config_rst)); 
mux6 mux_4097 (.in({n14749_2, n14748_0, n14663_0/**/, n14662_0, n14641_0, n14640_0}), .out(n8566), .config_in(config_chain[12293:12291]), .config_rst(config_rst)); 
mux6 mux_4098 (.in({n10419_0, n10418_0/**/, n10403_0, n10402_0, n10267_0, n10266_2}), .out(n8567), .config_in(config_chain[12296:12294]), .config_rst(config_rst)); 
mux6 mux_4099 (.in({n14481_1, n14480_0, n14473_1/**/, n14472_0, n14443_0, n14442_0}), .out(n8568), .config_in(config_chain[12299:12297]), .config_rst(config_rst)); 
mux6 mux_4100 (.in({n10643_0, n10642_0, n10635_0, n10634_0, n10523_0, n10522_2}), .out(n8569), .config_in(config_chain[12302:12300]), .config_rst(config_rst)); 
mux6 mux_4101 (.in({n14713_0, n14712_0/**/, n14703_0, n14702_0, n14673_0, n14672_0}), .out(n8570), .config_in(config_chain[12305:12303]), .config_rst(config_rst)); 
mux6 mux_4102 (.in({n10427_0, n10426_0, n10389_0, n10388_0, n10355_0, n10354_1}), .out(n8571), .config_in(config_chain[12308:12306]), .config_rst(config_rst)); 
mux6 mux_4103 (.in({n14433_2, n14432_0, n14415_0, n14414_0, n14383_0/**/, n14382_0}), .out(n8572), .config_in(config_chain[12311:12309]), .config_rst(config_rst)); 
mux6 mux_4104 (.in({n10679_0, n10678_0, n10665_0, n10664_0, n10525_0, n10524_2}), .out(n8573), .config_in(config_chain[12314:12312]), .config_rst(config_rst)); 
mux6 mux_4105 (.in({n14735_1, n14734_0, n14721_0, n14720_0, n14695_2, n14694_0}), .out(n8574), .config_in(config_chain[12317:12315]), .config_rst(config_rst)); 
mux6 mux_4106 (.in({n10411_0, n10410_0, n10383_0, n10382_0, n10375_0, n10374_0}), .out(n8575), .config_in(config_chain[12320:12318]), .config_rst(config_rst)); 
mux6 mux_4107 (.in({n14465_2, n14464_0, n14451_0, n14450_0, n14409_0, n14408_0/**/}), .out(n8576), .config_in(config_chain[12323:12321]), .config_rst(config_rst)); 
mux6 mux_4108 (.in({n10935_0, n10934_0, n10919_0, n10918_0, n10905_0, n10904_0}), .out(n8623), .config_in(config_chain[12326:12324]), .config_rst(config_rst)); 
mux6 mux_4109 (.in({n14751_1, n14750_0, n14735_0, n14734_0, n14721_0, n14720_0}), .out(n8624), .config_in(config_chain[12329:12327]), .config_rst(config_rst)); 
mux6 mux_4110 (.in({n10629_0, n10628_0, n10621_0, n10620_1, n10613_0, n10612_1}), .out(n8625), .config_in(config_chain[12332:12330]), .config_rst(config_rst)); 
mux6 mux_4111 (.in({n14453_0, n14452_0, n14445_0, n14444_0, n14409_0, n14408_1}), .out(n8626), .config_in(config_chain[12335:12333]), .config_rst(config_rst)); 
mux6 mux_4112 (.in({n10943_0, n10942_0/**/, n10927_0, n10926_0, n10869_0, n10868_1}), .out(n8627), .config_in(config_chain[12338:12336]), .config_rst(config_rst)); 
mux6 mux_4113 (.in({n14767_1, n14766_0, n14759_1, n14758_0, n14617_0, n14616_1}), .out(n8628), .config_in(config_chain[12341:12339]), .config_rst(config_rst)); 
mux6 mux_4114 (.in({n10659_0, n10658_0, n10651_0, n10650_0, n10645_0, n10644_0}), .out(n8629), .config_in(config_chain[12344:12342]), .config_rst(config_rst)); 
mux6 mux_4115 (.in({n14489_1, n14488_0, n14475_0, n14474_0, n14461_0/**/, n14460_0}), .out(n8630), .config_in(config_chain[12347:12345]), .config_rst(config_rst)); 
mux6 mux_4116 (.in({n10891_0, n10890_0, n10885_0, n10884_1, n10877_0, n10876_1/**/}), .out(n8631), .config_in(config_chain[12350:12348]), .config_rst(config_rst)); 
mux6 mux_4117 (.in({n14707_0, n14706_0, n14681_0, n14680_1, n14649_0, n14648_1}), .out(n8632), .config_in(config_chain[12353:12351]), .config_rst(config_rst)); 
mux6 mux_4118 (.in({n10681_0, n10680_0, n10673_0, n10672_0, n10667_0, n10666_0}), .out(n8633), .config_in(config_chain[12356:12354]), .config_rst(config_rst)); 
mux6 mux_4119 (.in({n14497_1, n14496_0, n14483_0, n14482_0, n14353_0, n14352_1}), .out(n8634), .config_in(config_chain[12359:12357]), .config_rst(config_rst)); 
mux6 mux_4120 (.in({n10913_0, n10912_0, n10907_0, n10906_0, n10899_0, n10898_0/**/}), .out(n8635), .config_in(config_chain[12362:12360]), .config_rst(config_rst)); 
mux6 mux_4121 (.in({n14737_0/**/, n14736_0, n14729_0, n14728_0, n14723_0, n14722_0}), .out(n8636), .config_in(config_chain[12365:12363]), .config_rst(config_rst)); 
mux6 mux_4122 (.in({n10689_0, n10688_0, n10631_0, n10630_0, n10615_0, n10614_1}), .out(n8637), .config_in(config_chain[12368:12366]), .config_rst(config_rst)); 
mux6 mux_4123 (.in({n14447_0, n14446_0, n14417_0, n14416_1, n14385_0, n14384_1}), .out(n8638), .config_in(config_chain[12371:12369]), .config_rst(config_rst)); 
mux6 mux_4124 (.in({n10945_0, n10944_0, n10937_0, n10936_0/**/, n10929_0, n10928_0}), .out(n8639), .config_in(config_chain[12374:12372]), .config_rst(config_rst)); 
mux6 mux_4125 (.in({n14761_1, n14760_0, n14745_0/**/, n14744_0, n14625_0, n14624_1}), .out(n8640), .config_in(config_chain[12377:12375]), .config_rst(config_rst)); 
mux6 mux_4126 (.in({n10653_0, n10652_0, n10639_0, n10638_0, n10623_0, n10622_1}), .out(n8641), .config_in(config_chain[12380:12378]), .config_rst(config_rst)); 
mux6 mux_4127 (.in({n14469_0, n14468_0, n14463_0, n14462_0, n14455_0, n14454_0}), .out(n8642), .config_in(config_chain[12383:12381]), .config_rst(config_rst)); 
mux6 mux_4128 (.in({n10953_0, n10952_0, n10879_0, n10878_1, n10871_0, n10870_1/**/}), .out(n8643), .config_in(config_chain[12386:12384]), .config_rst(config_rst)); 
mux6 mux_4129 (.in({n14769_1, n14768_0, n14709_0, n14708_0/**/, n14657_0, n14656_1}), .out(n8644), .config_in(config_chain[12389:12387]), .config_rst(config_rst)); 
mux6 mux_4130 (.in({n10675_0, n10674_0, n10669_0, n10668_0, n10661_0, n10660_0}), .out(n8645), .config_in(config_chain[12392:12390]), .config_rst(config_rst)); 
mux6 mux_4131 (.in({n14499_1, n14498_0, n14491_1, n14490_0, n14485_0/**/, n14484_0}), .out(n8646), .config_in(config_chain[12395:12393]), .config_rst(config_rst)); 
mux6 mux_4132 (.in({n10915_0, n10914_0, n10901_0, n10900_0, n10887_0, n10886_1}), .out(n8647), .config_in(config_chain[12398:12396]), .config_rst(config_rst)); 
mux6 mux_4133 (.in({n14731_0, n14730_0/**/, n14725_0, n14724_0, n14717_0, n14716_0}), .out(n8648), .config_in(config_chain[12401:12399]), .config_rst(config_rst)); 
mux6 mux_4134 (.in({n10691_0, n10690_0/**/, n10617_0, n10616_1, n10609_0, n10608_1}), .out(n8649), .config_in(config_chain[12404:12402]), .config_rst(config_rst)); 
mux6 mux_4135 (.in({n14507_1, n14506_0, n14393_0, n14392_1, n14361_0, n14360_1/**/}), .out(n8650), .config_in(config_chain[12407:12405]), .config_rst(config_rst)); 
mux6 mux_4136 (.in({n10939_0, n10938_0/**/, n10923_0, n10922_0, n10909_0, n10908_0}), .out(n8651), .config_in(config_chain[12410:12408]), .config_rst(config_rst)); 
mux6 mux_4137 (.in({n14755_1, n14754_0, n14747_0, n14746_0, n14739_0, n14738_0/**/}), .out(n8652), .config_in(config_chain[12413:12411]), .config_rst(config_rst)); 
mux6 mux_4138 (.in({n10641_0, n10640_0/**/, n10633_0, n10632_0, n10625_0, n10624_1}), .out(n8653), .config_in(config_chain[12416:12414]), .config_rst(config_rst)); 
mux6 mux_4139 (.in({n14471_0, n14470_0, n14457_0, n14456_0, n14425_0, n14424_1}), .out(n8654), .config_in(config_chain[12419:12417]), .config_rst(config_rst)); 
mux6 mux_4140 (.in({n10947_0/**/, n10946_0, n10873_0, n10872_1, n10867_0, n10866_1}), .out(n8655), .config_in(config_chain[12422:12420]), .config_rst(config_rst)); 
mux6 mux_4141 (.in({n14695_1, n14694_1, n14665_0, n14664_1, n14633_0, n14632_1}), .out(n8656), .config_in(config_chain[12425:12423]), .config_rst(config_rst)); 
mux6 mux_4142 (.in({n10677_0, n10676_0/**/, n10663_0, n10662_0, n10649_0, n10648_0}), .out(n8657), .config_in(config_chain[12428:12426]), .config_rst(config_rst)); 
mux6 mux_4143 (.in({n14493_1, n14492_0, n14479_0, n14478_0, n14465_1, n14464_0}), .out(n8658), .config_in(config_chain[12431:12429]), .config_rst(config_rst)); 
mux6 mux_4144 (.in({n10895_0, n10894_0, n10889_0, n10888_1, n10881_0, n10880_1}), .out(n8659), .config_in(config_chain[12434:12432]), .config_rst(config_rst)); 
mux6 mux_4145 (.in({n14719_0, n14718_0, n14711_0, n14710_0, n14697_1, n14696_1}), .out(n8660), .config_in(config_chain[12437:12435]), .config_rst(config_rst)); 
mux6 mux_4146 (.in({n10685_0/**/, n10684_0, n10671_0, n10670_0, n10611_0, n10610_1}), .out(n8661), .config_in(config_chain[12440:12438]), .config_rst(config_rst)); 
mux6 mux_4147 (.in({n14509_1/**/, n14508_0, n14501_1, n14500_0, n14369_0, n14368_1}), .out(n8662), .config_in(config_chain[12443:12441]), .config_rst(config_rst)); 
mux6 mux_4148 (.in({n10925_0, n10924_0/**/, n10917_0, n10916_0, n10911_0, n10910_0}), .out(n8663), .config_in(config_chain[12446:12444]), .config_rst(config_rst)); 
mux6 mux_4149 (.in({n14757_1, n14756_0, n14741_0, n14740_0, n14727_1, n14726_0}), .out(n8664), .config_in(config_chain[12449:12447]), .config_rst(config_rst)); 
mux6 mux_4150 (.in({n10635_0, n10634_0/**/, n10619_0, n10618_1, n10523_0, n10522_2}), .out(n8665), .config_in(config_chain[12452:12450]), .config_rst(config_rst)); 
mux6 mux_4151 (.in({n14459_0, n14458_0, n14451_0, n14450_0/**/, n14441_0, n14440_1}), .out(n8666), .config_in(config_chain[12455:12453]), .config_rst(config_rst)); 
mux6 mux_4152 (.in({n10949_0, n10948_0, n10941_0, n10940_0/**/, n10933_0, n10932_0}), .out(n8667), .config_in(config_chain[12458:12456]), .config_rst(config_rst)); 
mux6 mux_4153 (.in({n14765_1, n14764_0, n14749_1, n14748_0, n14641_0/**/, n14640_1}), .out(n8668), .config_in(config_chain[12461:12459]), .config_rst(config_rst)); 
mux6 mux_4154 (.in({n10657_0, n10656_0, n10643_0, n10642_0, n10525_0, n10524_2}), .out(n8669), .config_in(config_chain[12464:12462]), .config_rst(config_rst)); 
mux6 mux_4155 (.in({n14481_0, n14480_0, n14473_0, n14472_0, n14443_0, n14442_1}), .out(n8670), .config_in(config_chain[12467:12465]), .config_rst(config_rst)); 
mux6 mux_4156 (.in({n10955_0, n10954_0, n10897_0, n10896_0, n10883_0, n10882_1/**/}), .out(n8671), .config_in(config_chain[12470:12468]), .config_rst(config_rst)); 
mux6 mux_4157 (.in({n14713_0/**/, n14712_0, n14705_0, n14704_1, n14673_0, n14672_1}), .out(n8672), .config_in(config_chain[12473:12471]), .config_rst(config_rst)); 
mux6 mux_4158 (.in({n10687_0, n10686_0, n10679_0, n10678_0, n10627_0, n10626_1}), .out(n8673), .config_in(config_chain[12476:12474]), .config_rst(config_rst)); 
mux6 mux_4159 (.in({n14503_1, n14502_0, n14433_1, n14432_1, n14377_0, n14376_1}), .out(n8674), .config_in(config_chain[12479:12477]), .config_rst(config_rst)); 
mux6 mux_4160 (.in({n11213_0, n11212_0, n11155_0, n11154_0, n11139_0, n11138_1}), .out(n8721), .config_in(config_chain[12482:12480]), .config_rst(config_rst)); 
mux6 mux_4161 (.in({n14787_1, n14786_0/**/, n14729_0, n14728_0, n14713_0, n14712_1}), .out(n8722), .config_in(config_chain[12485:12483]), .config_rst(config_rst)); 
mux6 mux_4162 (.in({n10935_0, n10934_0, n10927_0, n10926_0, n10919_0, n10918_0}), .out(n8723), .config_in(config_chain[12488:12486]), .config_rst(config_rst)); 
mux6 mux_4163 (.in({n14519_1, n14518_0, n14511_1, n14510_0, n14503_0, n14502_0}), .out(n8724), .config_in(config_chain[12491:12489]), .config_rst(config_rst)); 
mux6 mux_4164 (.in({n11177_0, n11176_0, n11163_0, n11162_0, n11147_0, n11146_1}), .out(n8725), .config_in(config_chain[12494:12492]), .config_rst(config_rst)); 
mux6 mux_4165 (.in({n14751_0, n14750_0, n14745_0, n14744_0, n14737_0, n14736_0}), .out(n8726), .config_in(config_chain[12497:12495]), .config_rst(config_rst)); 
mux6 mux_4166 (.in({n10951_0, n10950_0, n10877_0, n10876_1, n10869_0, n10868_1}), .out(n8727), .config_in(config_chain[12500:12498]), .config_rst(config_rst)); 
mux6 mux_4167 (.in({n14527_1, n14526_0/**/, n14467_0, n14466_0, n14453_0, n14452_1}), .out(n8728), .config_in(config_chain[12503:12501]), .config_rst(config_rst)); 
mux6 mux_4168 (.in({n11199_0, n11198_0, n11193_0, n11192_0, n11185_0, n11184_0}), .out(n8729), .config_in(config_chain[12506:12504]), .config_rst(config_rst)); 
mux6 mux_4169 (.in({n14773_1, n14772_0, n14767_0, n14766_0/**/, n14759_0, n14758_0}), .out(n8730), .config_in(config_chain[12509:12507]), .config_rst(config_rst)); 
mux6 mux_4170 (.in({n10899_0, n10898_0, n10891_0, n10890_0, n10885_0, n10884_1}), .out(n8731), .config_in(config_chain[12512:12510]), .config_rst(config_rst)); 
mux6 mux_4171 (.in({n14489_0, n14488_0, n14475_0, n14474_0, n14461_0, n14460_1}), .out(n8732), .config_in(config_chain[12515:12513]), .config_rst(config_rst)); 
mux6 mux_4172 (.in({n11215_0, n11214_0, n11207_0, n11206_0/**/, n11133_0, n11132_1}), .out(n8733), .config_in(config_chain[12518:12516]), .config_rst(config_rst)); 
mux6 mux_4173 (.in({n14789_1, n14788_0, n14715_0, n14714_1/**/, n14707_0, n14706_1}), .out(n8734), .config_in(config_chain[12521:12519]), .config_rst(config_rst)); 
mux6 mux_4174 (.in({n10937_0, n10936_0, n10921_0, n10920_0, n10907_0, n10906_0/**/}), .out(n8735), .config_in(config_chain[12524:12522]), .config_rst(config_rst)); 
mux6 mux_4175 (.in({n14513_1, n14512_0, n14505_0, n14504_0/**/, n14497_0, n14496_0}), .out(n8736), .config_in(config_chain[12527:12525]), .config_rst(config_rst)); 
mux6 mux_4176 (.in({n11165_0, n11164_0, n11157_0, n11156_0/**/, n11149_0, n11148_1}), .out(n8737), .config_in(config_chain[12530:12528]), .config_rst(config_rst)); 
mux6 mux_4177 (.in({n14753_0, n14752_0, n14739_0, n14738_0, n14723_0, n14722_1}), .out(n8738), .config_in(config_chain[12533:12531]), .config_rst(config_rst)); 
mux6 mux_4178 (.in({n10945_0, n10944_0/**/, n10929_0, n10928_0, n10871_0, n10870_1}), .out(n8739), .config_in(config_chain[12536:12534]), .config_rst(config_rst)); 
mux6 mux_4179 (.in({n14529_1, n14528_0, n14521_1, n14520_0, n14447_0, n14446_1}), .out(n8740), .config_in(config_chain[12539:12537]), .config_rst(config_rst)); 
mux6 mux_4180 (.in({n11187_0, n11186_0/**/, n11179_0, n11178_0, n11173_0, n11172_0}), .out(n8741), .config_in(config_chain[12542:12540]), .config_rst(config_rst)); 
mux6 mux_4181 (.in({n14775_1, n14774_0, n14761_0/**/, n14760_0, n14747_0, n14746_0}), .out(n8742), .config_in(config_chain[12545:12543]), .config_rst(config_rst)); 
mux6 mux_4182 (.in({n10893_0, n10892_0/**/, n10887_0, n10886_1, n10879_0, n10878_1}), .out(n8743), .config_in(config_chain[12548:12546]), .config_rst(config_rst)); 
mux6 mux_4183 (.in({n14477_0, n14476_0, n14469_0, n14468_0, n14463_0/**/, n14462_1}), .out(n8744), .config_in(config_chain[12551:12549]), .config_rst(config_rst)); 
mux6 mux_4184 (.in({n11209_0, n11208_0, n11195_0/**/, n11194_0, n11135_0, n11134_1}), .out(n8745), .config_in(config_chain[12554:12552]), .config_rst(config_rst)); 
mux6 mux_4185 (.in({n14791_1, n14790_0, n14783_1/**/, n14782_0, n14709_0, n14708_1}), .out(n8746), .config_in(config_chain[12557:12555]), .config_rst(config_rst)); 
mux6 mux_4186 (.in({n10923_0, n10922_0/**/, n10915_0, n10914_0, n10909_0, n10908_0}), .out(n8747), .config_in(config_chain[12560:12558]), .config_rst(config_rst)); 
mux6 mux_4187 (.in({n14499_0, n14498_0, n14491_0, n14490_0, n14485_0, n14484_0}), .out(n8748), .config_in(config_chain[12563:12561]), .config_rst(config_rst)); 
mux6 mux_4188 (.in({n11217_0, n11216_0/**/, n11159_0, n11158_0, n11143_0, n11142_1}), .out(n8749), .config_in(config_chain[12566:12564]), .config_rst(config_rst)); 
mux6 mux_4189 (.in({n14733_0, n14732_0, n14725_0, n14724_1, n14717_0, n14716_1/**/}), .out(n8750), .config_in(config_chain[12569:12567]), .config_rst(config_rst)); 
mux6 mux_4190 (.in({n10947_0, n10946_0/**/, n10939_0, n10938_0, n10931_0, n10930_0}), .out(n8751), .config_in(config_chain[12572:12570]), .config_rst(config_rst)); 
mux6 mux_4191 (.in({n14523_1, n14522_0, n14507_0, n14506_0, n14449_0/**/, n14448_1}), .out(n8752), .config_in(config_chain[12575:12573]), .config_rst(config_rst)); 
mux6 mux_4192 (.in({n11219_0, n11218_0, n11181_0, n11180_0, n11167_0/**/, n11166_0}), .out(n8753), .config_in(config_chain[12578:12576]), .config_rst(config_rst)); 
mux6 mux_4193 (.in({n14793_1, n14792_0, n14763_0, n14762_0, n14755_0, n14754_0}), .out(n8754), .config_in(config_chain[12581:12579]), .config_rst(config_rst)); 
mux6 mux_4194 (.in({n10895_0, n10894_0, n10881_0, n10880_1, n10867_0, n10866_1/**/}), .out(n8755), .config_in(config_chain[12584:12582]), .config_rst(config_rst)); 
mux6 mux_4195 (.in({n14471_0, n14470_0, n14457_0/**/, n14456_1, n14433_1, n14432_1}), .out(n8756), .config_in(config_chain[12587:12585]), .config_rst(config_rst)); 
mux6 mux_4196 (.in({n11203_0, n11202_0, n11189_0, n11188_0/**/, n11109_0, n11108_1}), .out(n8757), .config_in(config_chain[12590:12588]), .config_rst(config_rst)); 
mux6 mux_4197 (.in({n14785_1, n14784_0, n14777_1, n14776_0/**/, n14695_1, n14694_1}), .out(n8758), .config_in(config_chain[12593:12591]), .config_rst(config_rst)); 
mux6 mux_4198 (.in({n10917_0, n10916_0, n10903_0, n10902_0/**/, n10889_0, n10888_1}), .out(n8759), .config_in(config_chain[12596:12594]), .config_rst(config_rst)); 
mux6 mux_4199 (.in({n14493_0, n14492_0/**/, n14487_1, n14486_0, n14479_0, n14478_0}), .out(n8760), .config_in(config_chain[12599:12597]), .config_rst(config_rst)); 
mux6 mux_4200 (.in({n11145_0, n11144_1/**/, n11137_0, n11136_1, n11131_0, n11130_1}), .out(n8761), .config_in(config_chain[12602:12600]), .config_rst(config_rst)); 
mux6 mux_4201 (.in({n14735_0, n14734_0, n14719_0, n14718_1, n14697_1, n14696_1}), .out(n8762), .config_in(config_chain[12605:12603]), .config_rst(config_rst)); 
mux6 mux_4202 (.in({n10941_0, n10940_0, n10933_0, n10932_0, n10925_0/**/, n10924_0}), .out(n8763), .config_in(config_chain[12608:12606]), .config_rst(config_rst)); 
mux6 mux_4203 (.in({n14525_1/**/, n14524_0, n14517_1, n14516_0, n14509_1, n14508_0}), .out(n8764), .config_in(config_chain[12611:12609]), .config_rst(config_rst)); 
mux6 mux_4204 (.in({n11169_0, n11168_0, n11161_0, n11160_0, n11153_0, n11152_1/**/}), .out(n8765), .config_in(config_chain[12614:12612]), .config_rst(config_rst)); 
mux6 mux_4205 (.in({n14757_0, n14756_0, n14743_0/**/, n14742_0, n14727_1, n14726_1}), .out(n8766), .config_in(config_chain[12617:12615]), .config_rst(config_rst)); 
mux6 mux_4206 (.in({n10955_0, n10954_0, n10949_0, n10948_0, n10875_0, n10874_1}), .out(n8767), .config_in(config_chain[12620:12618]), .config_rst(config_rst)); 
mux6 mux_4207 (.in({n14531_1, n14530_0, n14459_0, n14458_1/**/, n14451_0, n14450_1}), .out(n8768), .config_in(config_chain[12623:12621]), .config_rst(config_rst)); 
mux6 mux_4208 (.in({n11205_0, n11204_0/**/, n11191_0, n11190_0, n11175_0, n11174_0}), .out(n8769), .config_in(config_chain[12626:12624]), .config_rst(config_rst)); 
mux6 mux_4209 (.in({n14779_1, n14778_0, n14771_1, n14770_0, n14765_0, n14764_0}), .out(n8770), .config_in(config_chain[12629:12627]), .config_rst(config_rst)); 
mux6 mux_4210 (.in({n10905_0, n10904_0, n10897_0, n10896_0, n10785_0, n10784_2}), .out(n8771), .config_in(config_chain[12632:12630]), .config_rst(config_rst)); 
mux6 mux_4211 (.in({n14495_0, n14494_0, n14481_0, n14480_0, n14443_0, n14442_1}), .out(n8772), .config_in(config_chain[12635:12633]), .config_rst(config_rst)); 
mux6 mux_4212 (.in({n11465_0, n11464_0/**/, n11449_0, n11448_0, n11435_0, n11434_0}), .out(n8819), .config_in(config_chain[12638:12636]), .config_rst(config_rst)); 
mux6 mux_4213 (.in({n14795_1, n14794_0, n14779_0, n14778_0, n14765_0, n14764_0}), .out(n8820), .config_in(config_chain[12641:12639]), .config_rst(config_rst)); 
mux6 mux_4214 (.in({n11155_0, n11154_0, n11147_0, n11146_1, n11139_0, n11138_1}), .out(n8821), .config_in(config_chain[12644:12642]), .config_rst(config_rst)); 
mux6 mux_4215 (.in({n14497_0, n14496_0, n14489_0, n14488_0, n14481_0, n14480_1}), .out(n8822), .config_in(config_chain[12647:12645]), .config_rst(config_rst)); 
mux6 mux_4216 (.in({n11473_0, n11472_0, n11457_0, n11456_0, n11399_0, n11398_1}), .out(n8823), .config_in(config_chain[12650:12648]), .config_rst(config_rst)); 
mux6 mux_4217 (.in({n14811_1, n14810_0, n14803_1, n14802_0, n14729_0, n14728_1}), .out(n8824), .config_in(config_chain[12653:12651]), .config_rst(config_rst)); 
mux6 mux_4218 (.in({n11185_0, n11184_0, n11177_0, n11176_0, n11171_0, n11170_0}), .out(n8825), .config_in(config_chain[12656:12654]), .config_rst(config_rst)); 
mux6 mux_4219 (.in({n14533_1, n14532_0, n14519_0, n14518_0, n14505_0, n14504_0}), .out(n8826), .config_in(config_chain[12659:12657]), .config_rst(config_rst)); 
mux6 mux_4220 (.in({n11421_0, n11420_0, n11415_0, n11414_1, n11407_0, n11406_1}), .out(n8827), .config_in(config_chain[12662:12660]), .config_rst(config_rst)); 
mux6 mux_4221 (.in({n14751_0, n14750_0, n14745_0, n14744_1, n14737_0, n14736_1}), .out(n8828), .config_in(config_chain[12665:12663]), .config_rst(config_rst)); 
mux6 mux_4222 (.in({n11207_0, n11206_0, n11199_0, n11198_0, n11193_0, n11192_0}), .out(n8829), .config_in(config_chain[12668:12666]), .config_rst(config_rst)); 
mux6 mux_4223 (.in({n14541_1/**/, n14540_0, n14527_0, n14526_0, n14467_0, n14466_1}), .out(n8830), .config_in(config_chain[12671:12669]), .config_rst(config_rst)); 
mux6 mux_4224 (.in({n11443_0, n11442_0, n11437_0, n11436_0, n11429_0, n11428_0}), .out(n8831), .config_in(config_chain[12674:12672]), .config_rst(config_rst)); 
mux6 mux_4225 (.in({n14781_0, n14780_0, n14773_0, n14772_0, n14767_0, n14766_0}), .out(n8832), .config_in(config_chain[12677:12675]), .config_rst(config_rst)); 
mux6 mux_4226 (.in({n11215_0, n11214_0, n11157_0, n11156_0, n11141_0, n11140_1/**/}), .out(n8833), .config_in(config_chain[12680:12678]), .config_rst(config_rst)); 
mux6 mux_4227 (.in({n14491_0, n14490_0, n14483_0/**/, n14482_1, n14475_0, n14474_1}), .out(n8834), .config_in(config_chain[12683:12681]), .config_rst(config_rst)); 
mux6 mux_4228 (.in({n11475_0/**/, n11474_0, n11467_0, n11466_0, n11459_0, n11458_0}), .out(n8835), .config_in(config_chain[12686:12684]), .config_rst(config_rst)); 
mux6 mux_4229 (.in({n14805_1, n14804_0, n14789_0/**/, n14788_0, n14731_0, n14730_1}), .out(n8836), .config_in(config_chain[12689:12687]), .config_rst(config_rst)); 
mux6 mux_4230 (.in({n11179_0, n11178_0, n11165_0, n11164_0, n11149_0, n11148_1}), .out(n8837), .config_in(config_chain[12692:12690]), .config_rst(config_rst)); 
mux6 mux_4231 (.in({n14513_0, n14512_0, n14507_0/**/, n14506_0, n14499_0, n14498_0}), .out(n8838), .config_in(config_chain[12695:12693]), .config_rst(config_rst)); 
mux6 mux_4232 (.in({n11483_0, n11482_0, n11409_0, n11408_1/**/, n11401_0, n11400_1}), .out(n8839), .config_in(config_chain[12698:12696]), .config_rst(config_rst)); 
mux6 mux_4233 (.in({n14813_1/**/, n14812_0, n14753_0, n14752_0, n14739_0, n14738_1}), .out(n8840), .config_in(config_chain[12701:12699]), .config_rst(config_rst)); 
mux6 mux_4234 (.in({n11201_0, n11200_0, n11195_0, n11194_0, n11187_0, n11186_0}), .out(n8841), .config_in(config_chain[12704:12702]), .config_rst(config_rst)); 
mux6 mux_4235 (.in({n14543_1, n14542_0, n14535_1, n14534_0, n14529_0, n14528_0}), .out(n8842), .config_in(config_chain[12707:12705]), .config_rst(config_rst)); 
mux6 mux_4236 (.in({n11445_0, n11444_0, n11431_0, n11430_0, n11417_0, n11416_1}), .out(n8843), .config_in(config_chain[12710:12708]), .config_rst(config_rst)); 
mux6 mux_4237 (.in({n14775_0, n14774_0, n14769_0, n14768_0, n14761_0/**/, n14760_0}), .out(n8844), .config_in(config_chain[12713:12711]), .config_rst(config_rst)); 
mux6 mux_4238 (.in({n11217_0, n11216_0, n11143_0, n11142_1, n11135_0, n11134_1}), .out(n8845), .config_in(config_chain[12716:12714]), .config_rst(config_rst)); 
mux6 mux_4239 (.in({n14551_1/**/, n14550_0, n14477_0, n14476_1, n14469_0, n14468_1}), .out(n8846), .config_in(config_chain[12719:12717]), .config_rst(config_rst)); 
mux6 mux_4240 (.in({n11469_0, n11468_0, n11453_0, n11452_0, n11439_0, n11438_0}), .out(n8847), .config_in(config_chain[12722:12720]), .config_rst(config_rst)); 
mux6 mux_4241 (.in({n14799_1, n14798_0, n14791_0, n14790_0, n14783_0, n14782_0/**/}), .out(n8848), .config_in(config_chain[12725:12723]), .config_rst(config_rst)); 
mux6 mux_4242 (.in({n11167_0, n11166_0, n11159_0, n11158_0, n11151_0/**/, n11150_1}), .out(n8849), .config_in(config_chain[12728:12726]), .config_rst(config_rst)); 
mux6 mux_4243 (.in({n14515_0, n14514_0, n14501_0, n14500_0, n14485_0, n14484_1}), .out(n8850), .config_in(config_chain[12731:12729]), .config_rst(config_rst)); 
mux6 mux_4244 (.in({n11477_0, n11476_0, n11441_0, n11440_0/**/, n11403_0, n11402_1}), .out(n8851), .config_in(config_chain[12734:12732]), .config_rst(config_rst)); 
mux6 mux_4245 (.in({n14771_1, n14770_0, n14741_0, n14740_1, n14733_0/**/, n14732_1}), .out(n8852), .config_in(config_chain[12737:12735]), .config_rst(config_rst)); 
mux6 mux_4246 (.in({n11219_0, n11218_0, n11203_0, n11202_0/**/, n11189_0, n11188_0}), .out(n8853), .config_in(config_chain[12740:12738]), .config_rst(config_rst)); 
mux6 mux_4247 (.in({n14553_1, n14552_0/**/, n14537_1, n14536_0, n14523_0, n14522_0}), .out(n8854), .config_in(config_chain[12743:12741]), .config_rst(config_rst)); 
mux6 mux_4248 (.in({n11463_0, n11462_0, n11425_0, n11424_0, n11411_0, n11410_1}), .out(n8855), .config_in(config_chain[12746:12744]), .config_rst(config_rst)); 
mux6 mux_4249 (.in({n14793_1, n14792_0, n14763_0/**/, n14762_0, n14755_0, n14754_0}), .out(n8856), .config_in(config_chain[12749:12747]), .config_rst(config_rst)); 
mux6 mux_4250 (.in({n11211_0, n11210_0/**/, n11137_0, n11136_1, n11109_0, n11108_1}), .out(n8857), .config_in(config_chain[12752:12750]), .config_rst(config_rst)); 
mux6 mux_4251 (.in({n14545_1/**/, n14544_0, n14471_0, n14470_1, n14465_1, n14464_1}), .out(n8858), .config_in(config_chain[12755:12753]), .config_rst(config_rst)); 
mux6 mux_4252 (.in({n11455_0, n11454_0, n11447_0, n11446_0, n11353_0, n11352_2}), .out(n8859), .config_in(config_chain[12758:12756]), .config_rst(config_rst)); 
mux6 mux_4253 (.in({n14801_1, n14800_0, n14785_0/**/, n14784_0, n14695_1, n14694_1}), .out(n8860), .config_in(config_chain[12761:12759]), .config_rst(config_rst)); 
mux6 mux_4254 (.in({n11161_0, n11160_0, n11153_0, n11152_1/**/, n11145_0, n11144_1}), .out(n8861), .config_in(config_chain[12764:12762]), .config_rst(config_rst)); 
mux6 mux_4255 (.in({n14503_0, n14502_0, n14495_0, n14494_0, n14487_1, n14486_1}), .out(n8862), .config_in(config_chain[12767:12765]), .config_rst(config_rst)); 
mux6 mux_4256 (.in({n11479_0, n11478_0, n11471_0, n11470_0, n11375_0, n11374_1}), .out(n8863), .config_in(config_chain[12770:12768]), .config_rst(config_rst)); 
mux6 mux_4257 (.in({n14809_1, n14808_0/**/, n14735_0, n14734_1, n14697_1, n14696_1}), .out(n8864), .config_in(config_chain[12773:12771]), .config_rst(config_rst)); 
mux6 mux_4258 (.in({n11183_0, n11182_0, n11175_0, n11174_0, n11169_0, n11168_0}), .out(n8865), .config_in(config_chain[12776:12774]), .config_rst(config_rst)); 
mux6 mux_4259 (.in({n14525_0, n14524_0/**/, n14517_0, n14516_0, n14509_1, n14508_0}), .out(n8866), .config_in(config_chain[12779:12777]), .config_rst(config_rst)); 
mux6 mux_4260 (.in({n11427_0, n11426_0, n11413_0, n11412_1, n11397_0, n11396_1}), .out(n8867), .config_in(config_chain[12782:12780]), .config_rst(config_rst)); 
mux6 mux_4261 (.in({n14757_0, n14756_0/**/, n14749_1, n14748_1, n14743_0, n14742_1}), .out(n8868), .config_in(config_chain[12785:12783]), .config_rst(config_rst)); 
mux6 mux_4262 (.in({n11213_0, n11212_0, n11205_0, n11204_0, n11197_0, n11196_0}), .out(n8869), .config_in(config_chain[12788:12786]), .config_rst(config_rst)); 
mux6 mux_4263 (.in({n14547_1, n14546_0, n14531_1, n14530_0, n14473_0, n14472_1}), .out(n8870), .config_in(config_chain[12791:12789]), .config_rst(config_rst)); 
mux6 mux_4264 (.in({n11743_0, n11742_0, n11687_0, n11686_0, n11671_0, n11670_1}), .out(n8917), .config_in(config_chain[12794:12792]), .config_rst(config_rst)); 
mux6 mux_4265 (.in({n14829_0, n14828_0, n14773_0, n14772_0, n14757_0, n14756_1}), .out(n8918), .config_in(config_chain[12797:12795]), .config_rst(config_rst)); 
mux6 mux_4266 (.in({n11465_0, n11464_0, n11457_0, n11456_0, n11449_0, n11448_0}), .out(n8919), .config_in(config_chain[12800:12798]), .config_rst(config_rst)); 
mux6 mux_4267 (.in({n14563_0, n14562_0, n14555_0, n14554_0, n14547_0, n14546_0}), .out(n8920), .config_in(config_chain[12803:12801]), .config_rst(config_rst)); 
mux6 mux_4268 (.in({n11709_0, n11708_0, n11695_0, n11694_0, n11679_0, n11678_1}), .out(n8921), .config_in(config_chain[12806:12804]), .config_rst(config_rst)); 
mux6 mux_4269 (.in({n14795_0, n14794_0, n14789_0, n14788_0/**/, n14781_0, n14780_0}), .out(n8922), .config_in(config_chain[12809:12807]), .config_rst(config_rst)); 
mux6 mux_4270 (.in({n11481_0, n11480_0/**/, n11407_0, n11406_1, n11399_0, n11398_1}), .out(n8923), .config_in(config_chain[12812:12810]), .config_rst(config_rst)); 
mux6 mux_4271 (.in({n14571_0, n14570_0, n14511_0, n14510_0, n14497_0, n14496_1}), .out(n8924), .config_in(config_chain[12815:12813]), .config_rst(config_rst)); 
mux6 mux_4272 (.in({n11729_0, n11728_0, n11725_0, n11724_0/**/, n11717_0, n11716_0}), .out(n8925), .config_in(config_chain[12818:12816]), .config_rst(config_rst)); 
mux6 mux_4273 (.in({n14815_0, n14814_0, n14811_0, n14810_0/**/, n14803_0, n14802_0}), .out(n8926), .config_in(config_chain[12821:12819]), .config_rst(config_rst)); 
mux6 mux_4274 (.in({n11429_0, n11428_0, n11421_0, n11420_0, n11415_0, n11414_1}), .out(n8927), .config_in(config_chain[12824:12822]), .config_rst(config_rst)); 
mux6 mux_4275 (.in({n14533_0, n14532_0, n14519_0, n14518_0, n14505_0, n14504_1}), .out(n8928), .config_in(config_chain[12827:12825]), .config_rst(config_rst)); 
mux6 mux_4276 (.in({n11745_0, n11744_0, n11737_0, n11736_0, n11665_0, n11664_1}), .out(n8929), .config_in(config_chain[12830:12828]), .config_rst(config_rst)); 
mux6 mux_4277 (.in({n14831_0, n14830_0, n14759_0, n14758_1, n14751_0, n14750_1/**/}), .out(n8930), .config_in(config_chain[12833:12831]), .config_rst(config_rst)); 
mux6 mux_4278 (.in({n11467_0, n11466_0, n11451_0, n11450_0, n11437_0, n11436_0/**/}), .out(n8931), .config_in(config_chain[12836:12834]), .config_rst(config_rst)); 
mux6 mux_4279 (.in({n14557_0, n14556_0, n14549_0, n14548_0, n14541_0, n14540_0}), .out(n8932), .config_in(config_chain[12839:12837]), .config_rst(config_rst)); 
mux6 mux_4280 (.in({n11697_0, n11696_0, n11689_0, n11688_0, n11681_0, n11680_1}), .out(n8933), .config_in(config_chain[12842:12840]), .config_rst(config_rst)); 
mux6 mux_4281 (.in({n14797_0, n14796_0, n14783_0, n14782_0, n14767_0, n14766_1}), .out(n8934), .config_in(config_chain[12845:12843]), .config_rst(config_rst)); 
mux6 mux_4282 (.in({n11475_0, n11474_0, n11459_0, n11458_0, n11401_0, n11400_1}), .out(n8935), .config_in(config_chain[12848:12846]), .config_rst(config_rst)); 
mux6 mux_4283 (.in({n14573_0/**/, n14572_0, n14565_0, n14564_0, n14491_0, n14490_1}), .out(n8936), .config_in(config_chain[12851:12849]), .config_rst(config_rst)); 
mux6 mux_4284 (.in({n11719_0, n11718_0, n11711_0, n11710_0, n11705_0, n11704_0}), .out(n8937), .config_in(config_chain[12854:12852]), .config_rst(config_rst)); 
mux6 mux_4285 (.in({n14817_0, n14816_0, n14805_0, n14804_0/**/, n14791_0, n14790_0}), .out(n8938), .config_in(config_chain[12857:12855]), .config_rst(config_rst)); 
mux6 mux_4286 (.in({n11423_0, n11422_0, n11417_0, n11416_1, n11409_0, n11408_1}), .out(n8939), .config_in(config_chain[12860:12858]), .config_rst(config_rst)); 
mux6 mux_4287 (.in({n14521_0/**/, n14520_0, n14513_0, n14512_0, n14507_0, n14506_1}), .out(n8940), .config_in(config_chain[12863:12861]), .config_rst(config_rst)); 
mux6 mux_4288 (.in({n11739_0, n11738_0/**/, n11727_0, n11726_0, n11667_0, n11666_1}), .out(n8941), .config_in(config_chain[12866:12864]), .config_rst(config_rst)); 
mux6 mux_4289 (.in({n14833_0, n14832_0, n14825_0, n14824_0, n14753_0, n14752_1}), .out(n8942), .config_in(config_chain[12869:12867]), .config_rst(config_rst)); 
mux6 mux_4290 (.in({n11453_0, n11452_0, n11445_0, n11444_0, n11439_0, n11438_0/**/}), .out(n8943), .config_in(config_chain[12872:12870]), .config_rst(config_rst)); 
mux6 mux_4291 (.in({n14543_0/**/, n14542_0, n14535_0, n14534_0, n14529_0, n14528_0}), .out(n8944), .config_in(config_chain[12875:12873]), .config_rst(config_rst)); 
mux6 mux_4292 (.in({n11747_0, n11746_0, n11691_0, n11690_0, n11675_0, n11674_1}), .out(n8945), .config_in(config_chain[12878:12876]), .config_rst(config_rst)); 
mux6 mux_4293 (.in({n14777_0, n14776_0, n14769_0, n14768_1, n14761_0, n14760_1}), .out(n8946), .config_in(config_chain[12881:12879]), .config_rst(config_rst)); 
mux6 mux_4294 (.in({n11477_0, n11476_0/**/, n11469_0, n11468_0, n11461_0, n11460_0}), .out(n8947), .config_in(config_chain[12884:12882]), .config_rst(config_rst)); 
mux6 mux_4295 (.in({n14567_0, n14566_0, n14551_0, n14550_0, n14493_0, n14492_1}), .out(n8948), .config_in(config_chain[12887:12885]), .config_rst(config_rst)); 
mux6 mux_4296 (.in({n11713_0, n11712_0, n11699_0, n11698_0, n11663_0, n11662_1}), .out(n8949), .config_in(config_chain[12890:12888]), .config_rst(config_rst)); 
mux6 mux_4297 (.in({n14807_0, n14806_0, n14799_0, n14798_0, n14749_0, n14748_1}), .out(n8950), .config_in(config_chain[12893:12891]), .config_rst(config_rst)); 
mux6 mux_4298 (.in({n11441_0, n11440_0/**/, n11425_0, n11424_0, n11411_0, n11410_1}), .out(n8951), .config_in(config_chain[12896:12894]), .config_rst(config_rst)); 
mux6 mux_4299 (.in({n14531_0, n14530_0/**/, n14515_0, n14514_0, n14501_0, n14500_1}), .out(n8952), .config_in(config_chain[12899:12897]), .config_rst(config_rst)); 
mux6 mux_4300 (.in({n11733_0, n11732_0/**/, n11721_0, n11720_0, n11685_0, n11684_1}), .out(n8953), .config_in(config_chain[12902:12900]), .config_rst(config_rst)); 
mux6 mux_4301 (.in({n14827_0, n14826_0/**/, n14819_0, n14818_0, n14771_0, n14770_1}), .out(n8954), .config_in(config_chain[12905:12903]), .config_rst(config_rst)); 
mux6 mux_4302 (.in({n11463_0/**/, n11462_0, n11447_0, n11446_0, n11433_0, n11432_0}), .out(n8955), .config_in(config_chain[12908:12906]), .config_rst(config_rst)); 
mux6 mux_4303 (.in({n14537_0, n14536_0, n14523_0, n14522_0, n14433_0, n14432_2}), .out(n8956), .config_in(config_chain[12911:12909]), .config_rst(config_rst)); 
mux6 mux_4304 (.in({n11707_0, n11706_0, n11677_0, n11676_1/**/, n11669_0, n11668_1}), .out(n8957), .config_in(config_chain[12914:12912]), .config_rst(config_rst)); 
mux6 mux_4305 (.in({n14793_0, n14792_0, n14779_0, n14778_0, n14763_0, n14762_1}), .out(n8958), .config_in(config_chain[12917:12915]), .config_rst(config_rst)); 
mux6 mux_4306 (.in({n11471_0, n11470_0/**/, n11455_0, n11454_0, n11375_0, n11374_1}), .out(n8959), .config_in(config_chain[12920:12918]), .config_rst(config_rst)); 
mux6 mux_4307 (.in({n14569_0, n14568_0, n14561_0, n14560_0, n14465_0, n14464_1}), .out(n8960), .config_in(config_chain[12923:12921]), .config_rst(config_rst)); 
mux6 mux_4308 (.in({n11701_0, n11700_0, n11693_0, n11692_0, n11597_0, n11596_2}), .out(n8961), .config_in(config_chain[12926:12924]), .config_rst(config_rst)); 
mux6 mux_4309 (.in({n14801_0, n14800_0, n14787_0, n14786_0, n14695_0, n14694_2}), .out(n8962), .config_in(config_chain[12929:12927]), .config_rst(config_rst)); 
mux6 mux_4310 (.in({n11479_0, n11478_0, n11405_0, n11404_1/**/, n11397_0, n11396_1}), .out(n8963), .config_in(config_chain[12932:12930]), .config_rst(config_rst)); 
mux6 mux_4311 (.in({n14503_0/**/, n14502_1, n14495_0, n14494_1, n14487_0, n14486_1}), .out(n8964), .config_in(config_chain[12935:12933]), .config_rst(config_rst)); 
mux6 mux_4312 (.in({n11735_0, n11734_0, n11723_0, n11722_0, n11619_0, n11618_2}), .out(n8965), .config_in(config_chain[12938:12936]), .config_rst(config_rst)); 
mux6 mux_4313 (.in({n14821_0, n14820_0, n14809_0, n14808_0, n14727_0, n14726_1}), .out(n8966), .config_in(config_chain[12941:12939]), .config_rst(config_rst)); 
mux6 mux_4314 (.in({n11435_0, n11434_0, n11427_0, n11426_0, n11419_0, n11418_1/**/}), .out(n8967), .config_in(config_chain[12944:12942]), .config_rst(config_rst)); 
mux6 mux_4315 (.in({n14539_0, n14538_0, n14525_0, n14524_0/**/, n14509_0, n14508_1}), .out(n8968), .config_in(config_chain[12947:12945]), .config_rst(config_rst)); 
mux6 mux_4316 (.in({n11991_0, n11990_0, n11977_0, n11976_0, n11965_0, n11964_0}), .out(n9015), .config_in(config_chain[12950:12948]), .config_rst(config_rst)); 
mux6 mux_4317 (.in({n14835_0, n14834_0/**/, n14821_0, n14820_0, n14809_0, n14808_0}), .out(n9016), .config_in(config_chain[12953:12951]), .config_rst(config_rst)); 
mux6 mux_4318 (.in({n11687_0, n11686_0, n11679_0, n11678_1, n11671_0, n11670_1}), .out(n9017), .config_in(config_chain[12956:12954]), .config_rst(config_rst)); 
mux6 mux_4319 (.in({n14541_0, n14540_0, n14533_0, n14532_0, n14525_0, n14524_1}), .out(n9018), .config_in(config_chain[12959:12957]), .config_rst(config_rst)); 
mux6 mux_4320 (.in({n11999_0, n11998_0, n11985_0, n11984_0, n11929_0, n11928_1}), .out(n9019), .config_in(config_chain[12962:12960]), .config_rst(config_rst)); 
mux6 mux_4321 (.in({n14851_0, n14850_0, n14843_0, n14842_0, n14773_0, n14772_1}), .out(n9020), .config_in(config_chain[12965:12963]), .config_rst(config_rst)); 
mux6 mux_4322 (.in({n11717_0, n11716_0, n11709_0, n11708_0, n11703_0, n11702_0}), .out(n9021), .config_in(config_chain[12968:12966]), .config_rst(config_rst)); 
mux6 mux_4323 (.in({n14575_0, n14574_0, n14563_0, n14562_0, n14549_0, n14548_0}), .out(n9022), .config_in(config_chain[12971:12969]), .config_rst(config_rst)); 
mux6 mux_4324 (.in({n11951_0, n11950_0, n11945_0, n11944_1, n11937_0, n11936_1}), .out(n9023), .config_in(config_chain[12974:12972]), .config_rst(config_rst)); 
mux6 mux_4325 (.in({n14795_0, n14794_0/**/, n14789_0, n14788_1, n14781_0, n14780_1}), .out(n9024), .config_in(config_chain[12977:12975]), .config_rst(config_rst)); 
mux6 mux_4326 (.in({n11737_0, n11736_0, n11729_0, n11728_0, n11725_0, n11724_0}), .out(n9025), .config_in(config_chain[12980:12978]), .config_rst(config_rst)); 
mux6 mux_4327 (.in({n14583_0, n14582_0, n14571_0, n14570_0, n14511_0, n14510_1}), .out(n9026), .config_in(config_chain[12983:12981]), .config_rst(config_rst)); 
mux6 mux_4328 (.in({n11971_0, n11970_0, n11967_0, n11966_0, n11959_0, n11958_0}), .out(n9027), .config_in(config_chain[12986:12984]), .config_rst(config_rst)); 
mux6 mux_4329 (.in({n14823_0, n14822_0, n14815_0, n14814_0, n14811_0, n14810_0}), .out(n9028), .config_in(config_chain[12989:12987]), .config_rst(config_rst)); 
mux6 mux_4330 (.in({n11745_0, n11744_0/**/, n11689_0, n11688_0, n11673_0, n11672_1}), .out(n9029), .config_in(config_chain[12992:12990]), .config_rst(config_rst)); 
mux6 mux_4331 (.in({n14535_0, n14534_0, n14527_0/**/, n14526_1, n14519_0, n14518_1}), .out(n9030), .config_in(config_chain[12995:12993]), .config_rst(config_rst)); 
mux6 mux_4332 (.in({n12001_0, n12000_0, n11993_0, n11992_0/**/, n11987_0, n11986_0}), .out(n9031), .config_in(config_chain[12998:12996]), .config_rst(config_rst)); 
mux6 mux_4333 (.in({n14845_0, n14844_0, n14831_0, n14830_0, n14775_0, n14774_1}), .out(n9032), .config_in(config_chain[13001:12999]), .config_rst(config_rst)); 
mux6 mux_4334 (.in({n11711_0, n11710_0, n11697_0, n11696_0, n11681_0, n11680_1}), .out(n9033), .config_in(config_chain[13004:13002]), .config_rst(config_rst)); 
mux6 mux_4335 (.in({n14557_0, n14556_0, n14551_0, n14550_0, n14543_0, n14542_0/**/}), .out(n9034), .config_in(config_chain[13007:13005]), .config_rst(config_rst)); 
mux6 mux_4336 (.in({n12009_0, n12008_0, n11939_0, n11938_1, n11931_0, n11930_1}), .out(n9035), .config_in(config_chain[13010:13008]), .config_rst(config_rst)); 
mux6 mux_4337 (.in({n14853_0, n14852_0, n14797_0, n14796_0, n14783_0, n14782_1}), .out(n9036), .config_in(config_chain[13013:13011]), .config_rst(config_rst)); 
mux6 mux_4338 (.in({n11731_0, n11730_0/**/, n11727_0, n11726_0, n11719_0, n11718_0}), .out(n9037), .config_in(config_chain[13016:13014]), .config_rst(config_rst)); 
mux6 mux_4339 (.in({n14585_0, n14584_0, n14577_0, n14576_0, n14573_0, n14572_0}), .out(n9038), .config_in(config_chain[13019:13017]), .config_rst(config_rst)); 
mux6 mux_4340 (.in({n11973_0, n11972_0, n11961_0, n11960_0, n11947_0, n11946_1}), .out(n9039), .config_in(config_chain[13022:13020]), .config_rst(config_rst)); 
mux6 mux_4341 (.in({n14817_0, n14816_0, n14813_0, n14812_0, n14805_0, n14804_0}), .out(n9040), .config_in(config_chain[13025:13023]), .config_rst(config_rst)); 
mux6 mux_4342 (.in({n11747_0, n11746_0/**/, n11675_0, n11674_1, n11667_0, n11666_1}), .out(n9041), .config_in(config_chain[13028:13026]), .config_rst(config_rst)); 
mux6 mux_4343 (.in({n14593_0, n14592_0, n14521_0, n14520_1, n14513_0, n14512_1}), .out(n9042), .config_in(config_chain[13031:13029]), .config_rst(config_rst)); 
mux6 mux_4344 (.in({n11995_0, n11994_0/**/, n11981_0, n11980_0, n11969_0, n11968_0}), .out(n9043), .config_in(config_chain[13034:13032]), .config_rst(config_rst)); 
mux6 mux_4345 (.in({n14839_0, n14838_0, n14833_0, n14832_0, n14825_0, n14824_0}), .out(n9044), .config_in(config_chain[13037:13035]), .config_rst(config_rst)); 
mux6 mux_4346 (.in({n11699_0, n11698_0, n11691_0, n11690_0, n11683_0, n11682_1}), .out(n9045), .config_in(config_chain[13040:13038]), .config_rst(config_rst)); 
mux6 mux_4347 (.in({n14559_0, n14558_0, n14545_0, n14544_0, n14529_0/**/, n14528_1}), .out(n9046), .config_in(config_chain[13043:13041]), .config_rst(config_rst)); 
mux6 mux_4348 (.in({n12003_0, n12002_0, n11933_0, n11932_1, n11883_0, n11882_2/**/}), .out(n9047), .config_in(config_chain[13046:13044]), .config_rst(config_rst)); 
mux6 mux_4349 (.in({n14785_0, n14784_1/**/, n14777_0, n14776_1, n14727_0, n14726_2}), .out(n9048), .config_in(config_chain[13049:13047]), .config_rst(config_rst)); 
mux6 mux_4350 (.in({n11733_0, n11732_0, n11721_0, n11720_0, n11663_0, n11662_1}), .out(n9049), .config_in(config_chain[13052:13050]), .config_rst(config_rst)); 
mux6 mux_4351 (.in({n14579_0, n14578_0, n14567_0, n14566_0, n14509_0, n14508_1}), .out(n9050), .config_in(config_chain[13055:13053]), .config_rst(config_rst)); 
mux6 mux_4352 (.in({n11955_0/**/, n11954_0, n11941_0, n11940_1, n11905_0, n11904_1}), .out(n9051), .config_in(config_chain[13058:13056]), .config_rst(config_rst)); 
mux6 mux_4353 (.in({n14807_0/**/, n14806_0, n14799_0, n14798_0, n14749_0, n14748_1}), .out(n9052), .config_in(config_chain[13061:13059]), .config_rst(config_rst)); 
mux6 mux_4354 (.in({n11741_0, n11740_0/**/, n11685_0, n11684_1, n11669_0, n11668_1}), .out(n9053), .config_in(config_chain[13064:13062]), .config_rst(config_rst)); 
mux6 mux_4355 (.in({n14587_0, n14586_0, n14553_0, n14552_0, n14515_0, n14514_1}), .out(n9054), .config_in(config_chain[13067:13065]), .config_rst(config_rst)); 
mux6 mux_4356 (.in({n11983_0, n11982_0/**/, n11975_0, n11974_0, n11927_0, n11926_1}), .out(n9055), .config_in(config_chain[13070:13068]), .config_rst(config_rst)); 
mux6 mux_4357 (.in({n14841_0, n14840_0, n14827_0, n14826_0, n14771_0, n14770_1}), .out(n9056), .config_in(config_chain[13073:13071]), .config_rst(config_rst)); 
mux6 mux_4358 (.in({n11693_0, n11692_0, n11677_0, n11676_1, n11597_0, n11596_2}), .out(n9057), .config_in(config_chain[13076:13074]), .config_rst(config_rst)); 
mux6 mux_4359 (.in({n14547_0, n14546_0, n14539_0, n14538_0, n14433_0, n14432_2/**/}), .out(n9058), .config_in(config_chain[13079:13077]), .config_rst(config_rst)); 
mux6 mux_4360 (.in({n12005_0, n12004_0, n11997_0, n11996_0/**/, n11949_0, n11948_1}), .out(n9059), .config_in(config_chain[13082:13080]), .config_rst(config_rst)); 
mux6 mux_4361 (.in({n14849_0, n14848_0, n14793_0, n14792_1, n14779_0/**/, n14778_1}), .out(n9060), .config_in(config_chain[13085:13083]), .config_rst(config_rst)); 
mux6 mux_4362 (.in({n11715_0, n11714_0, n11701_0, n11700_0/**/, n11619_0, n11618_2}), .out(n9061), .config_in(config_chain[13088:13086]), .config_rst(config_rst)); 
mux6 mux_4363 (.in({n14569_0, n14568_0, n14561_0, n14560_0, n14465_0, n14464_2}), .out(n9062), .config_in(config_chain[13091:13089]), .config_rst(config_rst)); 
mux6 mux_4364 (.in({n11957_0, n11956_0, n11943_0, n11942_1, n11829_0, n11828_2}), .out(n9063), .config_in(config_chain[13094:13092]), .config_rst(config_rst)); 
mux6 mux_4365 (.in({n14801_0, n14800_0, n14787_0, n14786_1/**/, n14697_0, n14696_2}), .out(n9064), .config_in(config_chain[13097:13095]), .config_rst(config_rst)); 
mux6 mux_4366 (.in({n11743_0, n11742_0, n11735_0, n11734_0/**/, n11641_0, n11640_1}), .out(n9065), .config_in(config_chain[13100:13098]), .config_rst(config_rst)); 
mux6 mux_4367 (.in({n14589_0, n14588_0, n14517_0, n14516_1, n14487_0, n14486_1}), .out(n9066), .config_in(config_chain[13103:13101]), .config_rst(config_rst)); 
mux6 mux_4368 (.in({n12265_0, n12264_0, n12211_0, n12210_0, n12197_0, n12196_1}), .out(n9113), .config_in(config_chain[13106:13104]), .config_rst(config_rst)); 
mux6 mux_4369 (.in({n14869_0, n14868_0, n14815_0, n14814_0, n14801_0, n14800_1}), .out(n9114), .config_in(config_chain[13109:13107]), .config_rst(config_rst)); 
mux6 mux_4370 (.in({n11991_0, n11990_0, n11985_0, n11984_0, n11977_0, n11976_0}), .out(n9115), .config_in(config_chain[13112:13110]), .config_rst(config_rst)); 
mux6 mux_4371 (.in({n14603_0, n14602_0, n14595_0, n14594_0, n14589_0, n14588_0}), .out(n9116), .config_in(config_chain[13115:13113]), .config_rst(config_rst)); 
mux6 mux_4372 (.in({n12231_0, n12230_0, n12219_0, n12218_0, n12205_0, n12204_1}), .out(n9117), .config_in(config_chain[13118:13116]), .config_rst(config_rst)); 
mux6 mux_4373 (.in({n14835_0, n14834_0, n14831_0, n14830_0, n14823_0, n14822_0}), .out(n9118), .config_in(config_chain[13121:13119]), .config_rst(config_rst)); 
mux6 mux_4374 (.in({n12007_0, n12006_0, n11937_0, n11936_1, n11929_0, n11928_1}), .out(n9119), .config_in(config_chain[13124:13122]), .config_rst(config_rst)); 
mux6 mux_4375 (.in({n14611_0, n14610_0, n14555_0, n14554_0, n14541_0, n14540_1}), .out(n9120), .config_in(config_chain[13127:13125]), .config_rst(config_rst)); 
mux6 mux_4376 (.in({n12251_0, n12250_0, n12247_0, n12246_0, n12239_0, n12238_0}), .out(n9121), .config_in(config_chain[13130:13128]), .config_rst(config_rst)); 
mux6 mux_4377 (.in({n14855_0, n14854_0, n14851_0, n14850_0, n14843_0, n14842_0}), .out(n9122), .config_in(config_chain[13133:13131]), .config_rst(config_rst)); 
mux6 mux_4378 (.in({n11959_0, n11958_0, n11951_0, n11950_0, n11945_0, n11944_1}), .out(n9123), .config_in(config_chain[13136:13134]), .config_rst(config_rst)); 
mux6 mux_4379 (.in({n14575_0, n14574_0, n14563_0, n14562_0, n14549_0, n14548_1}), .out(n9124), .config_in(config_chain[13139:13137]), .config_rst(config_rst)); 
mux6 mux_4380 (.in({n12267_0, n12266_0, n12259_0, n12258_0, n12191_0, n12190_1}), .out(n9125), .config_in(config_chain[13142:13140]), .config_rst(config_rst)); 
mux6 mux_4381 (.in({n14871_0, n14870_0, n14803_0, n14802_1, n14795_0, n14794_1}), .out(n9126), .config_in(config_chain[13145:13143]), .config_rst(config_rst)); 
mux6 mux_4382 (.in({n11993_0, n11992_0, n11979_0, n11978_0, n11967_0, n11966_0}), .out(n9127), .config_in(config_chain[13148:13146]), .config_rst(config_rst)); 
mux6 mux_4383 (.in({n14597_0, n14596_0, n14591_0, n14590_0, n14583_0, n14582_0}), .out(n9128), .config_in(config_chain[13151:13149]), .config_rst(config_rst)); 
mux6 mux_4384 (.in({n12221_0, n12220_0, n12213_0, n12212_0, n12207_0, n12206_1}), .out(n9129), .config_in(config_chain[13154:13152]), .config_rst(config_rst)); 
mux6 mux_4385 (.in({n14837_0, n14836_0, n14825_0, n14824_0, n14811_0, n14810_1}), .out(n9130), .config_in(config_chain[13157:13155]), .config_rst(config_rst)); 
mux6 mux_4386 (.in({n12001_0, n12000_0, n11987_0, n11986_0, n11931_0, n11930_1}), .out(n9131), .config_in(config_chain[13160:13158]), .config_rst(config_rst)); 
mux6 mux_4387 (.in({n14613_0, n14612_0, n14605_0, n14604_0, n14535_0, n14534_1}), .out(n9132), .config_in(config_chain[13163:13161]), .config_rst(config_rst)); 
mux6 mux_4388 (.in({n12241_0, n12240_0, n12233_0, n12232_0, n12229_0, n12228_0}), .out(n9133), .config_in(config_chain[13166:13164]), .config_rst(config_rst)); 
mux6 mux_4389 (.in({n14857_0, n14856_0, n14845_0, n14844_0, n14833_0, n14832_0}), .out(n9134), .config_in(config_chain[13169:13167]), .config_rst(config_rst)); 
mux6 mux_4390 (.in({n11953_0, n11952_0, n11947_0, n11946_1, n11939_0, n11938_1}), .out(n9135), .config_in(config_chain[13172:13170]), .config_rst(config_rst)); 
mux6 mux_4391 (.in({n14565_0, n14564_0, n14557_0, n14556_0, n14551_0, n14550_1}), .out(n9136), .config_in(config_chain[13175:13173]), .config_rst(config_rst)); 
mux6 mux_4392 (.in({n12261_0, n12260_0, n12249_0, n12248_0, n12193_0, n12192_1}), .out(n9137), .config_in(config_chain[13178:13176]), .config_rst(config_rst)); 
mux6 mux_4393 (.in({n14873_0, n14872_0, n14865_0, n14864_0, n14797_0, n14796_1}), .out(n9138), .config_in(config_chain[13181:13179]), .config_rst(config_rst)); 
mux6 mux_4394 (.in({n11981_0, n11980_0, n11973_0, n11972_0, n11969_0, n11968_0}), .out(n9139), .config_in(config_chain[13184:13182]), .config_rst(config_rst)); 
mux6 mux_4395 (.in({n14585_0, n14584_0, n14577_0, n14576_0, n14573_0, n14572_0}), .out(n9140), .config_in(config_chain[13187:13185]), .config_rst(config_rst)); 
mux6 mux_4396 (.in({n12269_0, n12268_0, n12215_0, n12214_0, n12201_0, n12200_1}), .out(n9141), .config_in(config_chain[13190:13188]), .config_rst(config_rst)); 
mux6 mux_4397 (.in({n14819_0, n14818_0, n14813_0, n14812_1, n14805_0, n14804_1}), .out(n9142), .config_in(config_chain[13193:13191]), .config_rst(config_rst)); 
mux6 mux_4398 (.in({n12003_0, n12002_0, n11995_0, n11994_0, n11989_0, n11988_0}), .out(n9143), .config_in(config_chain[13196:13194]), .config_rst(config_rst)); 
mux6 mux_4399 (.in({n14607_0, n14606_0, n14593_0, n14592_0, n14537_0, n14536_1}), .out(n9144), .config_in(config_chain[13199:13197]), .config_rst(config_rst)); 
mux6 mux_4400 (.in({n12235_0, n12234_0, n12223_0, n12222_0, n12093_0, n12092_2}), .out(n9145), .config_in(config_chain[13202:13200]), .config_rst(config_rst)); 
mux6 mux_4401 (.in({n14847_0, n14846_0, n14839_0, n14838_0, n14697_0, n14696_2}), .out(n9146), .config_in(config_chain[13205:13203]), .config_rst(config_rst)); 
mux6 mux_4402 (.in({n11955_0, n11954_0, n11941_0, n11940_1, n11883_0, n11882_2}), .out(n9147), .config_in(config_chain[13208:13206]), .config_rst(config_rst)); 
mux6 mux_4403 (.in({n14559_0, n14558_0, n14545_0, n14544_1, n14487_0, n14486_2}), .out(n9148), .config_in(config_chain[13211:13209]), .config_rst(config_rst)); 
mux6 mux_4404 (.in({n12255_0, n12254_0, n12243_0, n12242_0, n12123_0, n12122_2}), .out(n9149), .config_in(config_chain[13214:13212]), .config_rst(config_rst)); 
mux6 mux_4405 (.in({n14867_0, n14866_0, n14859_0, n14858_0, n14727_0, n14726_2}), .out(n9150), .config_in(config_chain[13217:13215]), .config_rst(config_rst)); 
mux6 mux_4406 (.in({n11975_0, n11974_0, n11963_0, n11962_0, n11905_0, n11904_1}), .out(n9151), .config_in(config_chain[13220:13218]), .config_rst(config_rst)); 
mux6 mux_4407 (.in({n14579_0, n14578_0, n14567_0, n14566_0, n14531_0, n14530_1}), .out(n9152), .config_in(config_chain[13223:13221]), .config_rst(config_rst)); 
mux6 mux_4408 (.in({n12203_0, n12202_1, n12195_0, n12194_1, n12145_0, n12144_2}), .out(n9153), .config_in(config_chain[13226:13224]), .config_rst(config_rst)); 
mux6 mux_4409 (.in({n14821_0, n14820_0, n14807_0, n14806_1, n14749_0, n14748_2}), .out(n9154), .config_in(config_chain[13229:13227]), .config_rst(config_rst)); 
mux6 mux_4410 (.in({n11997_0, n11996_0, n11983_0, n11982_0, n11949_0, n11948_1}), .out(n9155), .config_in(config_chain[13232:13230]), .config_rst(config_rst)); 
mux6 mux_4411 (.in({n14609_0, n14608_0, n14601_0, n14600_0, n14553_0, n14552_1}), .out(n9156), .config_in(config_chain[13235:13233]), .config_rst(config_rst)); 
mux6 mux_4412 (.in({n12225_0, n12224_0, n12217_0, n12216_0, n12167_0, n12166_1}), .out(n9157), .config_in(config_chain[13238:13236]), .config_rst(config_rst)); 
mux6 mux_4413 (.in({n14841_0, n14840_0, n14829_0, n14828_0, n14771_0, n14770_1}), .out(n9158), .config_in(config_chain[13241:13239]), .config_rst(config_rst)); 
mux6 mux_4414 (.in({n12005_0, n12004_0, n11935_0, n11934_1, n11829_0, n11828_2}), .out(n9159), .config_in(config_chain[13244:13242]), .config_rst(config_rst)); 
mux6 mux_4415 (.in({n14547_0, n14546_1, n14539_0, n14538_1, n14433_0, n14432_2}), .out(n9160), .config_in(config_chain[13247:13245]), .config_rst(config_rst)); 
mux6 mux_4416 (.in({n12257_0, n12256_0, n12245_0, n12244_0, n12189_0, n12188_1}), .out(n9161), .config_in(config_chain[13250:13248]), .config_rst(config_rst)); 
mux6 mux_4417 (.in({n14861_0, n14860_0, n14849_0, n14848_0, n14695_0, n14694_2}), .out(n9162), .config_in(config_chain[13253:13251]), .config_rst(config_rst)); 
mux6 mux_4418 (.in({n11965_0, n11964_0, n11957_0, n11956_0, n11861_0, n11860_2}), .out(n9163), .config_in(config_chain[13256:13254]), .config_rst(config_rst)); 
mux6 mux_4419 (.in({n14581_0, n14580_0, n14569_0, n14568_0, n14465_0, n14464_2}), .out(n9164), .config_in(config_chain[13259:13257]), .config_rst(config_rst)); 
mux6 mux_4420 (.in({n12219_0, n12218_0, n12211_0, n12210_0, n12205_0, n12204_1}), .out(n9210), .config_in(config_chain[13262:13260]), .config_rst(config_rst)); 
mux6 mux_4421 (.in({n12259_0, n12258_0, n12251_0, n12250_0, n12247_0, n12246_0}), .out(n9213), .config_in(config_chain[13265:13263]), .config_rst(config_rst)); 
mux6 mux_4422 (.in({n12221_0, n12220_0, n12213_0, n12212_0, n12207_0, n12206_1}), .out(n9216), .config_in(config_chain[13268:13266]), .config_rst(config_rst)); 
mux6 mux_4423 (.in({n12261_0, n12260_0, n12253_0, n12252_0, n12249_0, n12248_0}), .out(n9219), .config_in(config_chain[13271:13269]), .config_rst(config_rst)); 
mux6 mux_4424 (.in({n12215_0, n12214_0, n12209_0, n12208_1, n12201_0, n12200_1}), .out(n9222), .config_in(config_chain[13274:13272]), .config_rst(config_rst)); 
mux6 mux_4425 (.in({n12255_0, n12254_0, n12243_0, n12242_0, n12123_0, n12122_2}), .out(n9225), .config_in(config_chain[13277:13275]), .config_rst(config_rst)); 
mux6 mux_4426 (.in({n12217_0, n12216_0, n12203_0, n12202_1, n12167_0, n12166_1}), .out(n9228), .config_in(config_chain[13280:13278]), .config_rst(config_rst)); 
mux6 mux_4427 (.in({n12257_0, n12256_0, n12245_0, n12244_0, n12091_0, n12090_2}), .out(n9231), .config_in(config_chain[13283:13281]), .config_rst(config_rst)); 
mux6 mux_4428 (.in({n14685_0, n14684_0, n14653_0, n14652_0, n14615_0, n14614_0}), .out(n9258), .config_in(config_chain[13286:13284]), .config_rst(config_rst)); 
mux6 mux_4429 (.in({n14681_1, n14680_0, n14649_1, n14648_0, n14619_0, n14618_0}), .out(n9261), .config_in(config_chain[13289:13287]), .config_rst(config_rst)); 
mux6 mux_4430 (.in({n14683_0, n14682_0, n14661_0, n14660_0, n14623_0, n14622_0}), .out(n9264), .config_in(config_chain[13292:13290]), .config_rst(config_rst)); 
mux6 mux_4431 (.in({n14687_0, n14686_0, n14657_1, n14656_0, n14627_0, n14626_0}), .out(n9267), .config_in(config_chain[13295:13293]), .config_rst(config_rst)); 
mux6 mux_4432 (.in({n14691_0, n14690_0, n14669_0, n14668_0, n14631_0, n14630_0}), .out(n9270), .config_in(config_chain[13298:13296]), .config_rst(config_rst)); 
mux6 mux_4433 (.in({n14703_0, n14702_0, n14665_1, n14664_0, n14635_0, n14634_0}), .out(n9273), .config_in(config_chain[13301:13299]), .config_rst(config_rst)); 
mux6 mux_4434 (.in({n14695_2, n14694_0, n14677_0, n14676_0, n14645_0, n14644_0}), .out(n9276), .config_in(config_chain[13304:13302]), .config_rst(config_rst)); 
mux6 mux_4435 (.in({n14699_0, n14698_0, n14673_1, n14672_0, n14641_1, n14640_0}), .out(n9279), .config_in(config_chain[13307:13305]), .config_rst(config_rst)); 
mux6 mux_4436 (.in({n14723_1, n14722_0, n14715_1, n14714_0, n14621_0, n14620_0}), .out(n9306), .config_in(config_chain[13310:13308]), .config_rst(config_rst)); 
mux6 mux_4437 (.in({n14679_0, n14678_0, n14647_0, n14646_0, n14617_0, n14616_0}), .out(n9309), .config_in(config_chain[13313:13311]), .config_rst(config_rst)); 
mux6 mux_4438 (.in({n14717_1, n14716_0, n14681_0, n14680_0, n14629_0, n14628_0}), .out(n9312), .config_in(config_chain[13316:13314]), .config_rst(config_rst)); 
mux6 mux_4439 (.in({n14693_0, n14692_0, n14655_0, n14654_0, n14625_0, n14624_0}), .out(n9315), .config_in(config_chain[13319:13317]), .config_rst(config_rst)); 
mux6 mux_4440 (.in({n14719_1, n14718_0, n14689_0, n14688_0, n14637_0, n14636_0}), .out(n9318), .config_in(config_chain[13322:13320]), .config_rst(config_rst)); 
mux6 mux_4441 (.in({n14701_0, n14700_0, n14663_0, n14662_0, n14633_0, n14632_0}), .out(n9321), .config_in(config_chain[13325:13323]), .config_rst(config_rst)); 
mux6 mux_4442 (.in({n14721_1, n14720_0, n14713_1, n14712_0, n14705_0, n14704_0}), .out(n9324), .config_in(config_chain[13328:13326]), .config_rst(config_rst)); 
mux6 mux_4443 (.in({n14697_2, n14696_0, n14671_0, n14670_0, n14639_0, n14638_0}), .out(n9327), .config_in(config_chain[13331:13329]), .config_rst(config_rst)); 
mux6 mux_4444 (.in({n14707_0, n14706_0, n14681_0, n14680_0, n14649_0, n14648_0}), .out(n9354), .config_in(config_chain[13334:13332]), .config_rst(config_rst)); 
mux6 mux_4445 (.in({n14745_1, n14744_0, n14737_1, n14736_0, n14615_0, n14614_0}), .out(n9357), .config_in(config_chain[13337:13335]), .config_rst(config_rst)); 
mux6 mux_4446 (.in({n14709_0, n14708_0, n14679_0, n14678_0, n14657_0, n14656_0}), .out(n9360), .config_in(config_chain[13340:13338]), .config_rst(config_rst)); 
mux6 mux_4447 (.in({n14739_1, n14738_0, n14725_0, n14724_0, n14623_0, n14622_0}), .out(n9363), .config_in(config_chain[13343:13341]), .config_rst(config_rst)); 
mux6 mux_4448 (.in({n14711_0, n14710_0, n14687_0, n14686_0, n14665_0, n14664_0}), .out(n9366), .config_in(config_chain[13346:13344]), .config_rst(config_rst)); 
mux6 mux_4449 (.in({n14741_1, n14740_0, n14727_2, n14726_0, n14631_0, n14630_0/**/}), .out(n9369), .config_in(config_chain[13349:13347]), .config_rst(config_rst)); 
mux6 mux_4450 (.in({n14703_0, n14702_0, n14673_0, n14672_0/**/, n14641_0, n14640_0}), .out(n9372), .config_in(config_chain[13352:13350]), .config_rst(config_rst)); 
mux6 mux_4451 (.in({n14743_1, n14742_0, n14735_1, n14734_0, n14695_2, n14694_0}), .out(n9375), .config_in(config_chain[13355:13353]), .config_rst(config_rst)); 
mux6 mux_4452 (.in({n14767_1, n14766_0, n14759_1, n14758_0, n14617_0, n14616_1}), .out(n9402), .config_in(config_chain[13358:13356]), .config_rst(config_rst)); 
mux6 mux_4453 (.in({n14729_0, n14728_0, n14723_0, n14722_0, n14715_0, n14714_0}), .out(n9405), .config_in(config_chain[13361:13359]), .config_rst(config_rst)); 
mux6 mux_4454 (.in({n14761_1, n14760_0, n14745_0, n14744_0, n14625_0, n14624_1}), .out(n9408), .config_in(config_chain[13364:13362]), .config_rst(config_rst)); 
mux6 mux_4455 (.in({n14731_0, n14730_0, n14717_0, n14716_0, n14689_0, n14688_1}), .out(n9411), .config_in(config_chain[13367:13365]), .config_rst(config_rst)); 
mux6 mux_4456 (.in({n14763_1, n14762_0, n14747_0, n14746_0, n14633_0, n14632_1}), .out(n9414), .config_in(config_chain[13370:13368]), .config_rst(config_rst)); 
mux6 mux_4457 (.in({n14733_0, n14732_0, n14719_0, n14718_0, n14697_1, n14696_1}), .out(n9417), .config_in(config_chain[13373:13371]), .config_rst(config_rst)); 
mux6 mux_4458 (.in({n14765_1, n14764_0, n14757_1, n14756_0, n14749_1, n14748_0}), .out(n9420), .config_in(config_chain[13376:13374]), .config_rst(config_rst)); 
mux6 mux_4459 (.in({n14721_0, n14720_0, n14713_0, n14712_0, n14705_0, n14704_1}), .out(n9423), .config_in(config_chain[13379:13377]), .config_rst(config_rst)); 
mux6 mux_4460 (.in({n14751_0, n14750_0, n14745_0, n14744_0, n14737_0, n14736_0}), .out(n9450), .config_in(config_chain[13382:13380]), .config_rst(config_rst)); 
mux6 mux_4461 (.in({n14789_1, n14788_0, n14781_1, n14780_0, n14707_0, n14706_1}), .out(n9453), .config_in(config_chain[13385:13383]), .config_rst(config_rst)); 
mux6 mux_4462 (.in({n14753_0, n14752_0, n14739_0, n14738_0, n14723_0, n14722_1}), .out(n9456), .config_in(config_chain[13388:13386]), .config_rst(config_rst)); 
mux6 mux_4463 (.in({n14783_1, n14782_0, n14769_0, n14768_0, n14709_0, n14708_1}), .out(n9459), .config_in(config_chain[13391:13389]), .config_rst(config_rst)); 
mux6 mux_4464 (.in({n14755_0, n14754_0, n14741_0, n14740_0, n14725_0, n14724_1}), .out(n9462), .config_in(config_chain[13394:13392]), .config_rst(config_rst)); 
mux6 mux_4465 (.in({n14785_1, n14784_0, n14711_0, n14710_1, n14695_1, n14694_1}), .out(n9465), .config_in(config_chain[13397:13395]), .config_rst(config_rst)); 
mux6 mux_4466 (.in({n14743_0, n14742_0, n14735_0, n14734_0, n14727_1, n14726_1}), .out(n9468), .config_in(config_chain[13400:13398]), .config_rst(config_rst)); 
mux6 mux_4467 (.in({n14787_1, n14786_0, n14779_1, n14778_0, n14771_1, n14770_0}), .out(n9471), .config_in(config_chain[13403:13401]), .config_rst(config_rst)); 
mux6 mux_4468 (.in({n14811_1, n14810_0, n14803_1, n14802_0, n14729_0/**/, n14728_1}), .out(n9498), .config_in(config_chain[13406:13404]), .config_rst(config_rst)); 
mux6 mux_4469 (.in({n14773_0, n14772_0, n14767_0, n14766_0, n14759_0, n14758_0}), .out(n9501), .config_in(config_chain[13409:13407]), .config_rst(config_rst)); 
mux6 mux_4470 (.in({n14805_1, n14804_0, n14789_0, n14788_0, n14731_0, n14730_1}), .out(n9504), .config_in(config_chain[13412:13410]), .config_rst(config_rst)); 
mux6 mux_4471 (.in({n14775_0, n14774_0, n14761_0, n14760_0, n14747_0, n14746_1}), .out(n9507), .config_in(config_chain[13415:13413]), .config_rst(config_rst)); 
mux6 mux_4472 (.in({n14807_1, n14806_0, n14791_0, n14790_0, n14733_0, n14732_1}), .out(n9510), .config_in(config_chain[13418:13416]), .config_rst(config_rst)); 
mux6 mux_4473 (.in({n14793_1, n14792_0, n14777_0, n14776_0, n14763_0, n14762_0}), .out(n9513), .config_in(config_chain[13421:13419]), .config_rst(config_rst)); 
mux6 mux_4474 (.in({n14809_1, n14808_0, n14801_1, n14800_0, n14697_1, n14696_1}), .out(n9516), .config_in(config_chain[13424:13422]), .config_rst(config_rst)); 
mux6 mux_4475 (.in({n14765_0, n14764_0, n14757_0, n14756_0, n14749_1, n14748_1}), .out(n9519), .config_in(config_chain[13427:13425]), .config_rst(config_rst)); 
mux6 mux_4476 (.in({n14795_0, n14794_0, n14789_0, n14788_0, n14781_0, n14780_0}), .out(n9546), .config_in(config_chain[13430:13428]), .config_rst(config_rst)); 
mux6 mux_4477 (.in({n14831_0, n14830_0, n14823_0, n14822_0, n14751_0, n14750_1}), .out(n9549), .config_in(config_chain[13433:13431]), .config_rst(config_rst)); 
mux6 mux_4478 (.in({n14797_0, n14796_0, n14783_0, n14782_0, n14767_0, n14766_1}), .out(n9552), .config_in(config_chain[13436:13434]), .config_rst(config_rst)); 
mux6 mux_4479 (.in({n14825_0, n14824_0, n14813_0, n14812_0, n14753_0, n14752_1}), .out(n9555), .config_in(config_chain[13439:13437]), .config_rst(config_rst)); 
mux6 mux_4480 (.in({n14799_0, n14798_0, n14785_0, n14784_0, n14769_0, n14768_1}), .out(n9558), .config_in(config_chain[13442:13440]), .config_rst(config_rst)); 
mux6 mux_4481 (.in({n14827_0, n14826_0, n14771_0, n14770_1, n14755_0, n14754_1}), .out(n9561), .config_in(config_chain[13445:13443]), .config_rst(config_rst)); 
mux6 mux_4482 (.in({n14787_0, n14786_0, n14779_0, n14778_0, n14695_0, n14694_2}), .out(n9564), .config_in(config_chain[13448:13446]), .config_rst(config_rst)); 
mux6 mux_4483 (.in({n14829_0, n14828_0, n14821_0, n14820_0, n14727_0, n14726_1}), .out(n9567), .config_in(config_chain[13451:13449]), .config_rst(config_rst)); 
mux6 mux_4484 (.in({n14851_0, n14850_0, n14843_0, n14842_0, n14773_0, n14772_1}), .out(n9594), .config_in(config_chain[13454:13452]), .config_rst(config_rst)); 
mux6 mux_4485 (.in({n14815_0, n14814_0, n14811_0, n14810_0, n14803_0, n14802_0}), .out(n9597), .config_in(config_chain[13457:13455]), .config_rst(config_rst)); 
mux6 mux_4486 (.in({n14845_0, n14844_0, n14831_0, n14830_0, n14775_0, n14774_1}), .out(n9600), .config_in(config_chain[13460:13458]), .config_rst(config_rst)); 
mux6 mux_4487 (.in({n14817_0, n14816_0, n14805_0, n14804_0, n14791_0, n14790_1}), .out(n9603), .config_in(config_chain[13463:13461]), .config_rst(config_rst)); 
mux6 mux_4488 (.in({n14847_0, n14846_0, n14833_0, n14832_0, n14777_0/**/, n14776_1}), .out(n9606), .config_in(config_chain[13466:13464]), .config_rst(config_rst)); 
mux6 mux_4489 (.in({n14819_0, n14818_0, n14807_0, n14806_0/**/, n14749_0, n14748_1}), .out(n9609), .config_in(config_chain[13469:13467]), .config_rst(config_rst)); 
mux6 mux_4490 (.in({n14849_0, n14848_0, n14841_0, n14840_0, n14793_0, n14792_1}), .out(n9612), .config_in(config_chain[13472:13470]), .config_rst(config_rst)); 
mux6 mux_4491 (.in({n14809_0, n14808_0, n14801_0, n14800_0, n14697_0, n14696_2}), .out(n9615), .config_in(config_chain[13475:13473]), .config_rst(config_rst)); 
mux6 mux_4492 (.in({n14835_0, n14834_0, n14831_0, n14830_0, n14823_0, n14822_0}), .out(n9642), .config_in(config_chain[13478:13476]), .config_rst(config_rst)); 
mux6 mux_4493 (.in({n14871_0, n14870_0, n14863_0, n14862_0, n14795_0, n14794_1}), .out(n9645), .config_in(config_chain[13481:13479]), .config_rst(config_rst)); 
mux6 mux_4494 (.in({n14837_0, n14836_0, n14825_0, n14824_0, n14811_0, n14810_1}), .out(n9648), .config_in(config_chain[13484:13482]), .config_rst(config_rst)); 
mux6 mux_4495 (.in({n14865_0, n14864_0, n14853_0, n14852_0, n14797_0, n14796_1}), .out(n9651), .config_in(config_chain[13487:13485]), .config_rst(config_rst)); 
mux6 mux_4496 (.in({n14839_0, n14838_0, n14827_0, n14826_0, n14813_0, n14812_1}), .out(n9654), .config_in(config_chain[13490:13488]), .config_rst(config_rst)); 
mux6 mux_4497 (.in({n14867_0, n14866_0, n14799_0, n14798_1, n14727_0, n14726_2}), .out(n9657), .config_in(config_chain[13493:13491]), .config_rst(config_rst)); 
mux6 mux_4498 (.in({n14829_0, n14828_0, n14821_0, n14820_0, n14771_0, n14770_1}), .out(n9660), .config_in(config_chain[13496:13494]), .config_rst(config_rst)); 
mux6 mux_4499 (.in({n14869_0, n14868_0, n14861_0, n14860_0, n14695_0, n14694_2}), .out(n9663), .config_in(config_chain[13499:13497]), .config_rst(config_rst)); 
mux3 mux_4500 (.in({n12361_2, n563, n457}), .out(n9666), .config_in(config_chain[13501:13500]), .config_rst(config_rst)); 
buffer_wire buffer_9666 (.in(n9666), .out(n9666_0));
mux13 mux_4501 (.in({n13379_1, n13359_0/**/, n13339_1, n13319_0, n13299_1, n9819_1, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9667), .config_in(config_chain[13507:13502]), .config_rst(config_rst)); 
buffer_wire buffer_9667 (.in(n9667), .out(n9667_0));
mux3 mux_4502 (.in({n12271_1, n563, n457}), .out(n9668), .config_in(config_chain[13509:13508]), .config_rst(config_rst)); 
buffer_wire buffer_9668 (.in(n9668), .out(n9668_0));
mux13 mux_4503 (.in({n12605_2, n12585_0, n12565_0, n12545_0, n12525_0, n9759_1, n575, n567, n559, n475, n469, n463, n457}), .out(n9669), .config_in(config_chain[13515:13510]), .config_rst(config_rst)); 
buffer_wire buffer_9669 (.in(n9669), .out(n9669_0));
mux3 mux_4504 (.in({n12273_0, n563, n457}), .out(n9670), .config_in(config_chain[13517:13516]), .config_rst(config_rst)); 
buffer_wire buffer_9670 (.in(n9670), .out(n9670_0));
mux13 mux_4505 (.in({n12861_1, n12841_1, n12821_0/**/, n12801_1, n12781_0, n9779_1, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9671), .config_in(config_chain[13523:13518]), .config_rst(config_rst)); 
buffer_wire buffer_9671 (.in(n9671), .out(n9671_0));
mux3 mux_4506 (.in({n12275_0, n563, n457}), .out(n9672), .config_in(config_chain[13525:13524]), .config_rst(config_rst)); 
buffer_wire buffer_9672 (.in(n9672), .out(n9672_0));
mux13 mux_4507 (.in({n13119_1, n13099_0, n13079_0, n13059_0, n13039_0/**/, n9799_1, n2531, n2523, n2515, n2431, n2425, n2419, n2413}), .out(n9673), .config_in(config_chain[13531:13526]), .config_rst(config_rst)); 
buffer_wire buffer_9673 (.in(n9673), .out(n9673_0));
mux3 mux_4508 (.in({n12277_0/**/, n567, n457}), .out(n9674), .config_in(config_chain[13533:13532]), .config_rst(config_rst)); 
buffer_wire buffer_9674 (.in(n9674), .out(n9674_0));
mux13 mux_4509 (.in({n13381_1, n13361_0, n13341_0/**/, n13321_0, n13301_0, n9821_1, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9675), .config_in(config_chain[13539:13534]), .config_rst(config_rst)); 
buffer_wire buffer_9675 (.in(n9675), .out(n9675_0));
mux3 mux_4510 (.in({n12279_1, n567, n460}), .out(n9676), .config_in(config_chain[13541:13540]), .config_rst(config_rst)); 
buffer_wire buffer_9676 (.in(n9676), .out(n9676_0));
mux13 mux_4511 (.in({n12607_2, n12587_0, n12567_1, n12547_0, n12527_1, n9761_1, n575, n567, n559, n475, n469, n463, n457}), .out(n9677), .config_in(config_chain[13547:13542]), .config_rst(config_rst)); 
buffer_wire buffer_9677 (.in(n9677), .out(n9677_0));
mux3 mux_4512 (.in({n12281_0/**/, n567, n460}), .out(n9678), .config_in(config_chain[13549:13548]), .config_rst(config_rst)); 
buffer_wire buffer_9678 (.in(n9678), .out(n9678_0));
mux13 mux_4513 (.in({n12863_2, n12843_0, n12823_0, n12803_0, n12783_0, n9781_1, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9679), .config_in(config_chain[13555:13550]), .config_rst(config_rst)); 
buffer_wire buffer_9679 (.in(n9679), .out(n9679_0));
mux3 mux_4514 (.in({n12283_0, n567, n460}), .out(n9680), .config_in(config_chain[13557:13556]), .config_rst(config_rst)); 
buffer_wire buffer_9680 (.in(n9680), .out(n9680_0));
mux13 mux_4515 (.in({n13121_1, n13101_1, n13081_0, n13061_1, n13041_0, n9801_1, n2531, n2523, n2515/**/, n2431, n2425, n2419, n2413}), .out(n9681), .config_in(config_chain[13563:13558]), .config_rst(config_rst)); 
buffer_wire buffer_9681 (.in(n9681), .out(n9681_0));
mux3 mux_4516 (.in({n12285_0/**/, n567, n460}), .out(n9682), .config_in(config_chain[13565:13564]), .config_rst(config_rst)); 
buffer_wire buffer_9682 (.in(n9682), .out(n9682_0));
mux13 mux_4517 (.in({n13383_1, n13363_1, n13343_0, n13323_1, n13303_0/**/, n9823_1, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9683), .config_in(config_chain[13571:13566]), .config_rst(config_rst)); 
buffer_wire buffer_9683 (.in(n9683), .out(n9683_0));
mux3 mux_4518 (.in({n12287_1/**/, n571, n460}), .out(n9684), .config_in(config_chain[13573:13572]), .config_rst(config_rst)); 
buffer_wire buffer_9684 (.in(n9684), .out(n9684_0));
mux13 mux_4519 (.in({n12609_2, n12589_0, n12569_0/**/, n12549_0, n12529_0, n9763_1, n575, n567, n559, n475, n469, n463, n457}), .out(n9685), .config_in(config_chain[13579:13574]), .config_rst(config_rst)); 
buffer_wire buffer_9685 (.in(n9685), .out(n9685_0));
mux3 mux_4520 (.in({n12289_0/**/, n571, n463}), .out(n9686), .config_in(config_chain[13581:13580]), .config_rst(config_rst)); 
buffer_wire buffer_9686 (.in(n9686), .out(n9686_0));
mux13 mux_4521 (.in({n12865_2, n12845_0, n12825_1, n12805_0, n12785_1, n9783_1, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9687), .config_in(config_chain[13587:13582]), .config_rst(config_rst)); 
buffer_wire buffer_9687 (.in(n9687), .out(n9687_0));
mux3 mux_4522 (.in({n12291_0, n571, n463}), .out(n9688), .config_in(config_chain[13589:13588]), .config_rst(config_rst)); 
buffer_wire buffer_9688 (.in(n9688), .out(n9688_0));
mux13 mux_4523 (.in({n13123_2, n13103_0, n13083_0, n13063_0, n13043_0, n9803_1, n2531, n2523, n2515/**/, n2431, n2425, n2419, n2413}), .out(n9689), .config_in(config_chain[13595:13590]), .config_rst(config_rst)); 
buffer_wire buffer_9689 (.in(n9689), .out(n9689_0));
mux3 mux_4524 (.in({n12293_0, n571, n463}), .out(n9690), .config_in(config_chain[13597:13596]), .config_rst(config_rst)); 
buffer_wire buffer_9690 (.in(n9690), .out(n9690_0));
mux13 mux_4525 (.in({n13385_2, n13365_0, n13345_0, n13325_0, n13305_0, n9825_1, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9691), .config_in(config_chain[13603:13598]), .config_rst(config_rst)); 
buffer_wire buffer_9691 (.in(n9691), .out(n9691_0));
mux3 mux_4526 (.in({n12295_1, n571, n463}), .out(n9692), .config_in(config_chain[13605:13604]), .config_rst(config_rst)); 
buffer_wire buffer_9692 (.in(n9692), .out(n9692_0));
mux13 mux_4527 (.in({n12611_2, n12591_1, n12571_0, n12551_1, n12531_0, n9765_1, n575, n567, n559, n475, n469, n463, n457}), .out(n9693), .config_in(config_chain[13611:13606]), .config_rst(config_rst)); 
buffer_wire buffer_9693 (.in(n9693), .out(n9693_0));
mux3 mux_4528 (.in({n12297_0/**/, n575, n463}), .out(n9694), .config_in(config_chain[13613:13612]), .config_rst(config_rst)); 
buffer_wire buffer_9694 (.in(n9694), .out(n9694_0));
mux13 mux_4529 (.in({n12867_2, n12847_0, n12827_0, n12807_0, n12787_0, n9785_1, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9695), .config_in(config_chain[13619:13614]), .config_rst(config_rst)); 
buffer_wire buffer_9695 (.in(n9695), .out(n9695_0));
mux3 mux_4530 (.in({n12299_0, n575, n466}), .out(n9696), .config_in(config_chain[13621:13620]), .config_rst(config_rst)); 
buffer_wire buffer_9696 (.in(n9696), .out(n9696_0));
mux13 mux_4531 (.in({n13125_2, n13105_0, n13085_1/**/, n13065_0, n13045_1, n9805_1, n2531, n2523, n2515, n2431, n2425, n2419, n2413}), .out(n9697), .config_in(config_chain[13627:13622]), .config_rst(config_rst)); 
buffer_wire buffer_9697 (.in(n9697), .out(n9697_0));
mux3 mux_4532 (.in({n12301_0, n575, n466}), .out(n9698), .config_in(config_chain[13629:13628]), .config_rst(config_rst)); 
buffer_wire buffer_9698 (.in(n9698), .out(n9698_0));
mux13 mux_4533 (.in({n13387_2, n13367_0, n13347_1, n13327_0, n13307_1, n9827_1, n3509, n3501, n3493/**/, n3409, n3403, n3397, n3391}), .out(n9699), .config_in(config_chain[13635:13630]), .config_rst(config_rst)); 
buffer_wire buffer_9699 (.in(n9699), .out(n9699_0));
mux3 mux_4534 (.in({n12303_1, n575, n466}), .out(n9700), .config_in(config_chain[13637:13636]), .config_rst(config_rst)); 
buffer_wire buffer_9700 (.in(n9700), .out(n9700_0));
mux13 mux_4535 (.in({n12613_2, n12593_0, n12573_0, n12553_0/**/, n12533_0, n9767_1, n575, n567, n559, n475, n469, n463, n457}), .out(n9701), .config_in(config_chain[13643:13638]), .config_rst(config_rst)); 
buffer_wire buffer_9701 (.in(n9701), .out(n9701_0));
mux3 mux_4536 (.in({n12305_0, n575, n466}), .out(n9702), .config_in(config_chain[13645:13644]), .config_rst(config_rst)); 
buffer_wire buffer_9702 (.in(n9702), .out(n9702_0));
mux13 mux_4537 (.in({n12869_2, n12849_1, n12829_0, n12809_1, n12789_0, n9787_1, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9703), .config_in(config_chain[13651:13646]), .config_rst(config_rst)); 
buffer_wire buffer_9703 (.in(n9703), .out(n9703_0));
mux2 mux_4538 (.in({n12307_0, n466}), .out(n9704), .config_in(config_chain[13652:13652]), .config_rst(config_rst)); 
buffer_wire buffer_9704 (.in(n9704), .out(n9704_0));
mux13 mux_4539 (.in({n13127_2, n13107_0, n13087_0, n13067_0, n13047_0, n9807_1, n2531, n2523, n2515/**/, n2431, n2425, n2419, n2413}), .out(n9705), .config_in(config_chain[13658:13653]), .config_rst(config_rst)); 
buffer_wire buffer_9705 (.in(n9705), .out(n9705_0));
mux2 mux_4540 (.in({n12309_0/**/, n469}), .out(n9706), .config_in(config_chain[13659:13659]), .config_rst(config_rst)); 
buffer_wire buffer_9706 (.in(n9706), .out(n9706_0));
mux12 mux_4541 (.in({n13389_2, n13369_0, n13349_0/**/, n13329_0, n13309_0, n9829_1, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9707), .config_in(config_chain[13665:13660]), .config_rst(config_rst)); 
buffer_wire buffer_9707 (.in(n9707), .out(n9707_0));
mux2 mux_4542 (.in({n12311_1, n469}), .out(n9708), .config_in(config_chain[13666:13666]), .config_rst(config_rst)); 
buffer_wire buffer_9708 (.in(n9708), .out(n9708_0));
mux12 mux_4543 (.in({n12615_2, n12595_0/**/, n12575_1, n12555_0, n12535_1, n9769_1, n571, n563, n478, n472, n466, n460}), .out(n9709), .config_in(config_chain[13672:13667]), .config_rst(config_rst)); 
buffer_wire buffer_9709 (.in(n9709), .out(n9709_0));
mux2 mux_4544 (.in({n12313_0/**/, n469}), .out(n9710), .config_in(config_chain[13673:13673]), .config_rst(config_rst)); 
buffer_wire buffer_9710 (.in(n9710), .out(n9710_0));
mux12 mux_4545 (.in({n12871_2, n12851_0, n12831_0, n12811_0, n12791_0, n9789_1, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9711), .config_in(config_chain[13679:13674]), .config_rst(config_rst)); 
buffer_wire buffer_9711 (.in(n9711), .out(n9711_0));
mux2 mux_4546 (.in({n12315_0, n469}), .out(n9712), .config_in(config_chain[13680:13680]), .config_rst(config_rst)); 
buffer_wire buffer_9712 (.in(n9712), .out(n9712_0));
mux12 mux_4547 (.in({n13129_2, n13109_1, n13089_0, n13069_1, n13049_0, n9809_1, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9713), .config_in(config_chain[13686:13681]), .config_rst(config_rst)); 
buffer_wire buffer_9713 (.in(n9713), .out(n9713_0));
mux2 mux_4548 (.in({n12317_0, n469}), .out(n9714), .config_in(config_chain[13687:13687]), .config_rst(config_rst)); 
buffer_wire buffer_9714 (.in(n9714), .out(n9714_0));
mux11 mux_4549 (.in({n13371_1, n13351_0, n13331_1, n13311_0, n9831_1, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9715), .config_in(config_chain[13693:13688]), .config_rst(config_rst)); 
buffer_wire buffer_9715 (.in(n9715), .out(n9715_0));
mux2 mux_4550 (.in({n12319_1, n472}), .out(n9716), .config_in(config_chain[13694:13694]), .config_rst(config_rst)); 
buffer_wire buffer_9716 (.in(n9716), .out(n9716_0));
mux11 mux_4551 (.in({n12597_0, n12577_0, n12557_0, n12537_0/**/, n9771_1, n571, n563, n478, n472, n466, n460}), .out(n9717), .config_in(config_chain[13700:13695]), .config_rst(config_rst)); 
buffer_wire buffer_9717 (.in(n9717), .out(n9717_0));
mux2 mux_4552 (.in({n12321_0/**/, n472}), .out(n9718), .config_in(config_chain[13701:13701]), .config_rst(config_rst)); 
buffer_wire buffer_9718 (.in(n9718), .out(n9718_0));
mux11 mux_4553 (.in({n12853_0, n12833_1, n12813_0, n12793_1, n9791_1, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9719), .config_in(config_chain[13707:13702]), .config_rst(config_rst)); 
buffer_wire buffer_9719 (.in(n9719), .out(n9719_0));
mux2 mux_4554 (.in({n12323_0/**/, n472}), .out(n9720), .config_in(config_chain[13708:13708]), .config_rst(config_rst)); 
buffer_wire buffer_9720 (.in(n9720), .out(n9720_0));
mux11 mux_4555 (.in({n13111_0, n13091_0, n13071_0, n13051_0/**/, n9811_1, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9721), .config_in(config_chain[13714:13709]), .config_rst(config_rst)); 
buffer_wire buffer_9721 (.in(n9721), .out(n9721_0));
mux2 mux_4556 (.in({n12325_0/**/, n472}), .out(n9722), .config_in(config_chain[13715:13715]), .config_rst(config_rst)); 
buffer_wire buffer_9722 (.in(n9722), .out(n9722_0));
mux11 mux_4557 (.in({n13373_0/**/, n13353_0, n13333_0, n13313_0, n9833_1, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9723), .config_in(config_chain[13721:13716]), .config_rst(config_rst)); 
buffer_wire buffer_9723 (.in(n9723), .out(n9723_0));
mux2 mux_4558 (.in({n12327_1, n472}), .out(n9724), .config_in(config_chain[13722:13722]), .config_rst(config_rst)); 
buffer_wire buffer_9724 (.in(n9724), .out(n9724_0));
mux11 mux_4559 (.in({n12599_1, n12579_0, n12559_1, n12539_0, n9773_1, n571, n563, n478, n472, n466, n460}), .out(n9725), .config_in(config_chain[13728:13723]), .config_rst(config_rst)); 
buffer_wire buffer_9725 (.in(n9725), .out(n9725_0));
mux2 mux_4560 (.in({n12329_0/**/, n475}), .out(n9726), .config_in(config_chain[13729:13729]), .config_rst(config_rst)); 
buffer_wire buffer_9726 (.in(n9726), .out(n9726_0));
mux11 mux_4561 (.in({n12855_0, n12835_0, n12815_0, n12795_0, n9793_1, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9727), .config_in(config_chain[13735:13730]), .config_rst(config_rst)); 
buffer_wire buffer_9727 (.in(n9727), .out(n9727_0));
mux2 mux_4562 (.in({n12331_0, n475}), .out(n9728), .config_in(config_chain[13736:13736]), .config_rst(config_rst)); 
buffer_wire buffer_9728 (.in(n9728), .out(n9728_0));
mux11 mux_4563 (.in({n13113_0, n13093_1, n13073_0, n13053_1, n9813_1, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9729), .config_in(config_chain[13742:13737]), .config_rst(config_rst)); 
buffer_wire buffer_9729 (.in(n9729), .out(n9729_0));
mux2 mux_4564 (.in({n12333_0, n475}), .out(n9730), .config_in(config_chain[13743:13743]), .config_rst(config_rst)); 
buffer_wire buffer_9730 (.in(n9730), .out(n9730_0));
mux11 mux_4565 (.in({n13375_0, n13355_1, n13335_0, n13315_1, n9835_1, n3505, n3497/**/, n3412, n3406, n3400, n3394}), .out(n9731), .config_in(config_chain[13749:13744]), .config_rst(config_rst)); 
buffer_wire buffer_9731 (.in(n9731), .out(n9731_0));
mux2 mux_4566 (.in({n12335_1/**/, n475}), .out(n9732), .config_in(config_chain[13750:13750]), .config_rst(config_rst)); 
buffer_wire buffer_9732 (.in(n9732), .out(n9732_0));
mux11 mux_4567 (.in({n12601_0, n12581_0, n12561_0/**/, n12541_0, n9775_1, n571, n563, n478, n472, n466, n460}), .out(n9733), .config_in(config_chain[13756:13751]), .config_rst(config_rst)); 
buffer_wire buffer_9733 (.in(n9733), .out(n9733_0));
mux2 mux_4568 (.in({n12337_0, n475}), .out(n9734), .config_in(config_chain[13757:13757]), .config_rst(config_rst)); 
buffer_wire buffer_9734 (.in(n9734), .out(n9734_0));
mux11 mux_4569 (.in({n12857_1, n12837_0, n12817_1, n12797_0, n9795_1, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9735), .config_in(config_chain[13763:13758]), .config_rst(config_rst)); 
buffer_wire buffer_9735 (.in(n9735), .out(n9735_0));
mux2 mux_4570 (.in({n12339_0, n478}), .out(n9736), .config_in(config_chain[13764:13764]), .config_rst(config_rst)); 
buffer_wire buffer_9736 (.in(n9736), .out(n9736_0));
mux11 mux_4571 (.in({n13115_0, n13095_0, n13075_0, n13055_0, n9815_1, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9737), .config_in(config_chain[13770:13765]), .config_rst(config_rst)); 
buffer_wire buffer_9737 (.in(n9737), .out(n9737_0));
mux2 mux_4572 (.in({n12341_0/**/, n478}), .out(n9738), .config_in(config_chain[13771:13771]), .config_rst(config_rst)); 
buffer_wire buffer_9738 (.in(n9738), .out(n9738_0));
mux11 mux_4573 (.in({n13377_0, n13357_0, n13337_0, n13317_0, n9837_1, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9739), .config_in(config_chain[13777:13772]), .config_rst(config_rst)); 
buffer_wire buffer_9739 (.in(n9739), .out(n9739_0));
mux2 mux_4574 (.in({n12343_1/**/, n478}), .out(n9740), .config_in(config_chain[13778:13778]), .config_rst(config_rst)); 
buffer_wire buffer_9740 (.in(n9740), .out(n9740_0));
mux11 mux_4575 (.in({n12603_0, n12583_1, n12563_0, n12543_1, n9777_1, n571, n563, n478, n472, n466, n460}), .out(n9741), .config_in(config_chain[13784:13779]), .config_rst(config_rst)); 
buffer_wire buffer_9741 (.in(n9741), .out(n9741_0));
mux2 mux_4576 (.in({n12345_0/**/, n478}), .out(n9742), .config_in(config_chain[13785:13785]), .config_rst(config_rst)); 
buffer_wire buffer_9742 (.in(n9742), .out(n9742_0));
mux11 mux_4577 (.in({n12859_0, n12839_0, n12819_0, n12799_0, n9797_1, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9743), .config_in(config_chain[13791:13786]), .config_rst(config_rst)); 
buffer_wire buffer_9743 (.in(n9743), .out(n9743_0));
mux2 mux_4578 (.in({n12347_0, n478}), .out(n9744), .config_in(config_chain[13792:13792]), .config_rst(config_rst)); 
buffer_wire buffer_9744 (.in(n9744), .out(n9744_0));
mux11 mux_4579 (.in({n13117_1, n13097_0, n13077_1, n13057_0, n9817_1, n2527, n2519/**/, n2434, n2428, n2422, n2416}), .out(n9745), .config_in(config_chain[13798:13793]), .config_rst(config_rst)); 
buffer_wire buffer_9745 (.in(n9745), .out(n9745_0));
mux2 mux_4580 (.in({n12349_0/**/, n559}), .out(n9746), .config_in(config_chain[13799:13799]), .config_rst(config_rst)); 
buffer_wire buffer_9746 (.in(n9746), .out(n9746_0));
mux10 mux_4581 (.in({n14439_0, n14417_1, n14395_0, n14373_0, n9919_0, n7413, n7405, n7321, n7315, n7309}), .out(n9747), .config_in(config_chain[13805:13800]), .config_rst(config_rst)); 
buffer_wire buffer_9747 (.in(n9747), .out(n9747_0));
mux2 mux_4582 (.in({n12351_2, n559}), .out(n9748), .config_in(config_chain[13806:13806]), .config_rst(config_rst)); 
buffer_wire buffer_9748 (.in(n9748), .out(n9748_0));
mux2 mux_4583 (.in({n14625_1, n8383}), .out(n9749), .config_in(config_chain[13807:13807]), .config_rst(config_rst)); 
buffer_wire buffer_9749 (.in(n9749), .out(n9749_0));
mux2 mux_4584 (.in({n12353_2, n559}), .out(n9750), .config_in(config_chain[13808:13808]), .config_rst(config_rst)); 
buffer_wire buffer_9750 (.in(n9750), .out(n9750_0));
mux2 mux_4585 (.in({n14623_0, n8383}), .out(n9751), .config_in(config_chain[13809:13809]), .config_rst(config_rst)); 
buffer_wire buffer_9751 (.in(n9751), .out(n9751_0));
mux2 mux_4586 (.in({n12355_2, n559}), .out(n9752), .config_in(config_chain[13810:13810]), .config_rst(config_rst)); 
buffer_wire buffer_9752 (.in(n9752), .out(n9752_0));
mux2 mux_4587 (.in({n14621_0/**/, n8383}), .out(n9753), .config_in(config_chain[13811:13811]), .config_rst(config_rst)); 
buffer_wire buffer_9753 (.in(n9753), .out(n9753_0));
mux2 mux_4588 (.in({n12357_2, n559}), .out(n9754), .config_in(config_chain[13812:13812]), .config_rst(config_rst)); 
buffer_wire buffer_9754 (.in(n9754), .out(n9754_0));
mux2 mux_4589 (.in({n14619_0/**/, n8383}), .out(n9755), .config_in(config_chain[13813:13813]), .config_rst(config_rst)); 
buffer_wire buffer_9755 (.in(n9755), .out(n9755_0));
mux2 mux_4590 (.in({n12359_2, n563}), .out(n9756), .config_in(config_chain[13814:13814]), .config_rst(config_rst)); 
buffer_wire buffer_9756 (.in(n9756), .out(n9756_0));
mux2 mux_4591 (.in({n14617_1, n8387}), .out(n9757), .config_in(config_chain[13815:13815]), .config_rst(config_rst)); 
buffer_wire buffer_9757 (.in(n9757), .out(n9757_0));
mux13 mux_4592 (.in({n12605_2, n12585_0, n12565_0, n12545_0/**/, n12525_0, n9668_0, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9758), .config_in(config_chain[13821:13816]), .config_rst(config_rst)); 
buffer_wire buffer_9758 (.in(n9758), .out(n9758_0));
mux13 mux_4593 (.in({n13641_0, n13621_0, n13601_0, n13581_0, n13561_0, n9839_1, n4487, n4479, n4471, n4387, n4381/**/, n4375, n4369}), .out(n9759), .config_in(config_chain[13827:13822]), .config_rst(config_rst)); 
buffer_wire buffer_9759 (.in(n9759), .out(n9759_0));
mux13 mux_4594 (.in({n12607_2, n12587_0, n12567_1, n12547_0, n12527_1, n9676_0, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9760), .config_in(config_chain[13833:13828]), .config_rst(config_rst)); 
buffer_wire buffer_9760 (.in(n9760), .out(n9760_0));
mux13 mux_4595 (.in({n13643_1, n13623_0, n13603_1, n13583_0, n13563_1, n9841_1, n4487, n4479/**/, n4471, n4387, n4381, n4375, n4369}), .out(n9761), .config_in(config_chain[13839:13834]), .config_rst(config_rst)); 
buffer_wire buffer_9761 (.in(n9761), .out(n9761_0));
mux13 mux_4596 (.in({n12609_2, n12589_0, n12569_0, n12549_0, n12529_0, n9684_0/**/, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9762), .config_in(config_chain[13845:13840]), .config_rst(config_rst)); 
buffer_wire buffer_9762 (.in(n9762), .out(n9762_0));
mux13 mux_4597 (.in({n13645_1, n13625_0, n13605_0, n13585_0, n13565_0, n9843_1, n4487, n4479, n4471, n4387, n4381/**/, n4375, n4369}), .out(n9763), .config_in(config_chain[13851:13846]), .config_rst(config_rst)); 
buffer_wire buffer_9763 (.in(n9763), .out(n9763_0));
mux13 mux_4598 (.in({n12611_2, n12591_1, n12571_0, n12551_1, n12531_0, n9692_0, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9764), .config_in(config_chain[13857:13852]), .config_rst(config_rst)); 
buffer_wire buffer_9764 (.in(n9764), .out(n9764_0));
mux13 mux_4599 (.in({n13647_1, n13627_1, n13607_0, n13587_1, n13567_0, n9845_1, n4487, n4479, n4471, n4387, n4381/**/, n4375, n4369}), .out(n9765), .config_in(config_chain[13863:13858]), .config_rst(config_rst)); 
buffer_wire buffer_9765 (.in(n9765), .out(n9765_0));
mux13 mux_4600 (.in({n12613_2, n12593_0, n12573_0/**/, n12553_0, n12533_0, n9700_0, n1553, n1545, n1537, n1453, n1447, n1441, n1435}), .out(n9766), .config_in(config_chain[13869:13864]), .config_rst(config_rst)); 
buffer_wire buffer_9766 (.in(n9766), .out(n9766_0));
mux13 mux_4601 (.in({n13649_2, n13629_0, n13609_0, n13589_0, n13569_0, n9847_1, n4487, n4479, n4471, n4387, n4381, n4375, n4369/**/}), .out(n9767), .config_in(config_chain[13875:13870]), .config_rst(config_rst)); 
buffer_wire buffer_9767 (.in(n9767), .out(n9767_0));
mux12 mux_4602 (.in({n12615_2, n12595_0, n12575_1, n12555_0, n12535_1, n9708_0, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9768), .config_in(config_chain[13881:13876]), .config_rst(config_rst)); 
buffer_wire buffer_9768 (.in(n9768), .out(n9768_0));
mux12 mux_4603 (.in({n13651_2, n13631_0, n13611_1, n13591_0, n13571_1, n9849_1, n4483, n4475, n4390/**/, n4384, n4378, n4372}), .out(n9769), .config_in(config_chain[13887:13882]), .config_rst(config_rst)); 
buffer_wire buffer_9769 (.in(n9769), .out(n9769_0));
mux11 mux_4604 (.in({n12597_0, n12577_0/**/, n12557_0, n12537_0, n9716_0, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9770), .config_in(config_chain[13893:13888]), .config_rst(config_rst)); 
buffer_wire buffer_9770 (.in(n9770), .out(n9770_0));
mux11 mux_4605 (.in({n13633_0, n13613_0, n13593_0, n13573_0, n9851_1, n4483, n4475, n4390/**/, n4384, n4378, n4372}), .out(n9771), .config_in(config_chain[13899:13894]), .config_rst(config_rst)); 
buffer_wire buffer_9771 (.in(n9771), .out(n9771_0));
mux11 mux_4606 (.in({n12599_1, n12579_0, n12559_1/**/, n12539_0, n9724_0, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9772), .config_in(config_chain[13905:13900]), .config_rst(config_rst)); 
buffer_wire buffer_9772 (.in(n9772), .out(n9772_0));
mux11 mux_4607 (.in({n13635_1, n13615_0, n13595_1, n13575_0, n9853_1, n4483, n4475, n4390/**/, n4384, n4378, n4372}), .out(n9773), .config_in(config_chain[13911:13906]), .config_rst(config_rst)); 
buffer_wire buffer_9773 (.in(n9773), .out(n9773_0));
mux11 mux_4608 (.in({n12601_0, n12581_0, n12561_0, n12541_0, n9732_0/**/, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9774), .config_in(config_chain[13917:13912]), .config_rst(config_rst)); 
buffer_wire buffer_9774 (.in(n9774), .out(n9774_0));
mux11 mux_4609 (.in({n13637_0, n13617_0, n13597_0, n13577_0, n9855_1, n4483, n4475, n4390, n4384, n4378/**/, n4372}), .out(n9775), .config_in(config_chain[13923:13918]), .config_rst(config_rst)); 
buffer_wire buffer_9775 (.in(n9775), .out(n9775_0));
mux11 mux_4610 (.in({n12603_0, n12583_1, n12563_0, n12543_1, n9740_0/**/, n1549, n1541, n1456, n1450, n1444, n1438}), .out(n9776), .config_in(config_chain[13929:13924]), .config_rst(config_rst)); 
buffer_wire buffer_9776 (.in(n9776), .out(n9776_0));
mux11 mux_4611 (.in({n13639_0, n13619_1, n13599_0, n13579_1, n9857_1, n4483, n4475, n4390, n4384, n4378, n4372/**/}), .out(n9777), .config_in(config_chain[13935:13930]), .config_rst(config_rst)); 
buffer_wire buffer_9777 (.in(n9777), .out(n9777_0));
mux13 mux_4612 (.in({n12861_1, n12841_1, n12821_0, n12801_1/**/, n12781_0, n9670_0, n2531, n2523, n2515, n2431, n2425, n2419, n2413}), .out(n9778), .config_in(config_chain[13941:13936]), .config_rst(config_rst)); 
buffer_wire buffer_9778 (.in(n9778), .out(n9778_0));
mux13 mux_4613 (.in({n13905_0, n13885_1, n13865_0, n13845_1, n13825_0, n9859_0, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9779), .config_in(config_chain[13947:13942]), .config_rst(config_rst)); 
buffer_wire buffer_9779 (.in(n9779), .out(n9779_0));
mux13 mux_4614 (.in({n12863_2, n12843_0, n12823_0, n12803_0/**/, n12783_0, n9678_0, n2531, n2523, n2515, n2431, n2425, n2419, n2413}), .out(n9780), .config_in(config_chain[13953:13948]), .config_rst(config_rst)); 
buffer_wire buffer_9780 (.in(n9780), .out(n9780_0));
mux13 mux_4615 (.in({n13907_0, n13887_0, n13867_0, n13847_0, n13827_0, n9861_0, n5465, n5457, n5449/**/, n5365, n5359, n5353, n5347}), .out(n9781), .config_in(config_chain[13959:13954]), .config_rst(config_rst)); 
buffer_wire buffer_9781 (.in(n9781), .out(n9781_0));
mux13 mux_4616 (.in({n12865_2, n12845_0, n12825_1, n12805_0, n12785_1, n9686_0, n2531, n2523, n2515/**/, n2431, n2425, n2419, n2413}), .out(n9782), .config_in(config_chain[13965:13960]), .config_rst(config_rst)); 
buffer_wire buffer_9782 (.in(n9782), .out(n9782_0));
mux13 mux_4617 (.in({n13909_1, n13889_0, n13869_1, n13849_0, n13829_1, n9863_0, n5465, n5457, n5449/**/, n5365, n5359, n5353, n5347}), .out(n9783), .config_in(config_chain[13971:13966]), .config_rst(config_rst)); 
buffer_wire buffer_9783 (.in(n9783), .out(n9783_0));
mux13 mux_4618 (.in({n12867_2, n12847_0, n12827_0/**/, n12807_0, n12787_0, n9694_0, n2531, n2523, n2515, n2431, n2425, n2419, n2413}), .out(n9784), .config_in(config_chain[13977:13972]), .config_rst(config_rst)); 
buffer_wire buffer_9784 (.in(n9784), .out(n9784_0));
mux13 mux_4619 (.in({n13911_1, n13891_0, n13871_0, n13851_0, n13831_0/**/, n9865_0, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9785), .config_in(config_chain[13983:13978]), .config_rst(config_rst)); 
buffer_wire buffer_9785 (.in(n9785), .out(n9785_0));
mux13 mux_4620 (.in({n12869_2, n12849_1, n12829_0, n12809_1, n12789_0, n9702_0, n2531, n2523, n2515/**/, n2431, n2425, n2419, n2413}), .out(n9786), .config_in(config_chain[13989:13984]), .config_rst(config_rst)); 
buffer_wire buffer_9786 (.in(n9786), .out(n9786_0));
mux13 mux_4621 (.in({n13913_1, n13893_1, n13873_0/**/, n13853_1, n13833_0, n9867_0, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9787), .config_in(config_chain[13995:13990]), .config_rst(config_rst)); 
buffer_wire buffer_9787 (.in(n9787), .out(n9787_0));
mux12 mux_4622 (.in({n12871_2, n12851_0, n12831_0, n12811_0, n12791_0, n9710_0/**/, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9788), .config_in(config_chain[14001:13996]), .config_rst(config_rst)); 
buffer_wire buffer_9788 (.in(n9788), .out(n9788_0));
mux12 mux_4623 (.in({n13915_2, n13895_0/**/, n13875_0, n13855_0, n13835_0, n9869_0, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9789), .config_in(config_chain[14007:14002]), .config_rst(config_rst)); 
buffer_wire buffer_9789 (.in(n9789), .out(n9789_0));
mux11 mux_4624 (.in({n12853_0, n12833_1, n12813_0, n12793_1/**/, n9718_0, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9790), .config_in(config_chain[14013:14008]), .config_rst(config_rst)); 
buffer_wire buffer_9790 (.in(n9790), .out(n9790_0));
mux11 mux_4625 (.in({n13897_0, n13877_1, n13857_0, n13837_1, n9871_0, n5461, n5453/**/, n5368, n5362, n5356, n5350}), .out(n9791), .config_in(config_chain[14019:14014]), .config_rst(config_rst)); 
buffer_wire buffer_9791 (.in(n9791), .out(n9791_0));
mux11 mux_4626 (.in({n12855_0, n12835_0, n12815_0, n12795_0, n9726_0/**/, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9792), .config_in(config_chain[14025:14020]), .config_rst(config_rst)); 
buffer_wire buffer_9792 (.in(n9792), .out(n9792_0));
mux11 mux_4627 (.in({n13899_0, n13879_0, n13859_0, n13839_0, n9873_0, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9793), .config_in(config_chain[14031:14026]), .config_rst(config_rst)); 
buffer_wire buffer_9793 (.in(n9793), .out(n9793_0));
mux11 mux_4628 (.in({n12857_1, n12837_0, n12817_1/**/, n12797_0, n9734_0, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9794), .config_in(config_chain[14037:14032]), .config_rst(config_rst)); 
buffer_wire buffer_9794 (.in(n9794), .out(n9794_0));
mux11 mux_4629 (.in({n13901_1, n13881_0, n13861_1, n13841_0, n9875_0, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9795), .config_in(config_chain[14043:14038]), .config_rst(config_rst)); 
buffer_wire buffer_9795 (.in(n9795), .out(n9795_0));
mux11 mux_4630 (.in({n12859_0, n12839_0, n12819_0/**/, n12799_0, n9742_0, n2527, n2519, n2434, n2428, n2422, n2416}), .out(n9796), .config_in(config_chain[14049:14044]), .config_rst(config_rst)); 
buffer_wire buffer_9796 (.in(n9796), .out(n9796_0));
mux11 mux_4631 (.in({n13903_0, n13883_0/**/, n13863_0, n13843_0, n9877_0, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9797), .config_in(config_chain[14055:14050]), .config_rst(config_rst)); 
buffer_wire buffer_9797 (.in(n9797), .out(n9797_0));
mux13 mux_4632 (.in({n13119_1, n13099_0, n13079_0, n13059_0, n13039_0, n9672_0, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9798), .config_in(config_chain[14061:14056]), .config_rst(config_rst)); 
buffer_wire buffer_9798 (.in(n9798), .out(n9798_0));
mux13 mux_4633 (.in({n14169_0/**/, n14149_0, n14129_0, n14109_0, n14089_0, n9879_0, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9799), .config_in(config_chain[14067:14062]), .config_rst(config_rst)); 
buffer_wire buffer_9799 (.in(n9799), .out(n9799_0));
mux13 mux_4634 (.in({n13121_1, n13101_1/**/, n13081_0, n13061_1, n13041_0, n9680_0, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9800), .config_in(config_chain[14073:14068]), .config_rst(config_rst)); 
buffer_wire buffer_9800 (.in(n9800), .out(n9800_0));
mux13 mux_4635 (.in({n14171_0, n14151_1/**/, n14131_0, n14111_1, n14091_0, n9881_0, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9801), .config_in(config_chain[14079:14074]), .config_rst(config_rst)); 
buffer_wire buffer_9801 (.in(n9801), .out(n9801_0));
mux13 mux_4636 (.in({n13123_2, n13103_0, n13083_0, n13063_0/**/, n13043_0, n9688_0, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9802), .config_in(config_chain[14085:14080]), .config_rst(config_rst)); 
buffer_wire buffer_9802 (.in(n9802), .out(n9802_0));
mux13 mux_4637 (.in({n14173_0, n14153_0, n14133_0, n14113_0/**/, n14093_0, n9883_0, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9803), .config_in(config_chain[14091:14086]), .config_rst(config_rst)); 
buffer_wire buffer_9803 (.in(n9803), .out(n9803_0));
mux13 mux_4638 (.in({n13125_2, n13105_0, n13085_1, n13065_0, n13045_1/**/, n9696_0, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9804), .config_in(config_chain[14097:14092]), .config_rst(config_rst)); 
buffer_wire buffer_9804 (.in(n9804), .out(n9804_0));
mux13 mux_4639 (.in({n14175_1, n14155_0, n14135_1, n14115_0, n14095_1, n9885_0, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9805), .config_in(config_chain[14103:14098]), .config_rst(config_rst)); 
buffer_wire buffer_9805 (.in(n9805), .out(n9805_0));
mux13 mux_4640 (.in({n13127_2, n13107_0, n13087_0, n13067_0, n13047_0/**/, n9704_0, n3509, n3501, n3493, n3409, n3403, n3397, n3391}), .out(n9806), .config_in(config_chain[14109:14104]), .config_rst(config_rst)); 
buffer_wire buffer_9806 (.in(n9806), .out(n9806_0));
mux13 mux_4641 (.in({n14177_1, n14157_0, n14137_0, n14117_0, n14097_0, n9887_0, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9807), .config_in(config_chain[14115:14110]), .config_rst(config_rst)); 
buffer_wire buffer_9807 (.in(n9807), .out(n9807_0));
mux12 mux_4642 (.in({n13129_2, n13109_1, n13089_0/**/, n13069_1, n13049_0, n9712_0, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9808), .config_in(config_chain[14121:14116]), .config_rst(config_rst)); 
buffer_wire buffer_9808 (.in(n9808), .out(n9808_0));
mux12 mux_4643 (.in({n14179_1, n14159_1, n14139_0, n14119_1, n14099_0, n9889_0/**/, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9809), .config_in(config_chain[14127:14122]), .config_rst(config_rst)); 
buffer_wire buffer_9809 (.in(n9809), .out(n9809_0));
mux11 mux_4644 (.in({n13111_0, n13091_0/**/, n13071_0, n13051_0, n9720_0, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9810), .config_in(config_chain[14133:14128]), .config_rst(config_rst)); 
buffer_wire buffer_9810 (.in(n9810), .out(n9810_0));
mux11 mux_4645 (.in({n14161_0/**/, n14141_0, n14121_0, n14101_0, n9891_0, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9811), .config_in(config_chain[14139:14134]), .config_rst(config_rst)); 
buffer_wire buffer_9811 (.in(n9811), .out(n9811_0));
mux11 mux_4646 (.in({n13113_0/**/, n13093_1, n13073_0, n13053_1, n9728_0, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9812), .config_in(config_chain[14145:14140]), .config_rst(config_rst)); 
buffer_wire buffer_9812 (.in(n9812), .out(n9812_0));
mux11 mux_4647 (.in({n14163_0, n14143_1, n14123_0/**/, n14103_1, n9893_0, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9813), .config_in(config_chain[14151:14146]), .config_rst(config_rst)); 
buffer_wire buffer_9813 (.in(n9813), .out(n9813_0));
mux11 mux_4648 (.in({n13115_0, n13095_0/**/, n13075_0, n13055_0, n9736_0, n3505, n3497, n3412, n3406, n3400, n3394}), .out(n9814), .config_in(config_chain[14157:14152]), .config_rst(config_rst)); 
buffer_wire buffer_9814 (.in(n9814), .out(n9814_0));
mux11 mux_4649 (.in({n14165_0, n14145_0, n14125_0, n14105_0, n9895_0, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9815), .config_in(config_chain[14163:14158]), .config_rst(config_rst)); 
buffer_wire buffer_9815 (.in(n9815), .out(n9815_0));
mux11 mux_4650 (.in({n13117_1, n13097_0, n13077_1, n13057_0, n9744_0, n3505, n3497/**/, n3412, n3406, n3400, n3394}), .out(n9816), .config_in(config_chain[14169:14164]), .config_rst(config_rst)); 
buffer_wire buffer_9816 (.in(n9816), .out(n9816_0));
mux11 mux_4651 (.in({n14167_1, n14147_0, n14127_1/**/, n14107_0, n9897_0, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9817), .config_in(config_chain[14175:14170]), .config_rst(config_rst)); 
buffer_wire buffer_9817 (.in(n9817), .out(n9817_0));
mux13 mux_4652 (.in({n13379_1, n13359_0, n13339_1, n13319_0/**/, n13299_1, n9666_1, n4487, n4479, n4471, n4387, n4381, n4375, n4369}), .out(n9818), .config_in(config_chain[14181:14176]), .config_rst(config_rst)); 
buffer_wire buffer_9818 (.in(n9818), .out(n9818_0));
mux12 mux_4653 (.in({n14441_1, n14419_0, n14397_0, n14375_0/**/, n14353_1, n9899_0, n7417, n7405, n7321, n7315, n7309, n7303}), .out(n9819), .config_in(config_chain[14187:14182]), .config_rst(config_rst)); 
buffer_wire buffer_9819 (.in(n9819), .out(n9819_0));
mux13 mux_4654 (.in({n13381_1, n13361_0, n13341_0, n13321_0, n13301_0, n9674_1, n4487, n4479, n4471, n4387, n4381/**/, n4375, n4369}), .out(n9820), .config_in(config_chain[14193:14188]), .config_rst(config_rst)); 
buffer_wire buffer_9820 (.in(n9820), .out(n9820_0));
mux12 mux_4655 (.in({n14443_1, n14421_0, n14399_0, n14377_1, n14355_0, n9901_0/**/, n7417, n7409, n7321, n7315, n7309, n7303}), .out(n9821), .config_in(config_chain[14199:14194]), .config_rst(config_rst)); 
buffer_wire buffer_9821 (.in(n9821), .out(n9821_0));
mux13 mux_4656 (.in({n13383_1, n13363_1/**/, n13343_0, n13323_1, n13303_0, n9682_1, n4487, n4479, n4471, n4387, n4381, n4375, n4369}), .out(n9822), .config_in(config_chain[14205:14200]), .config_rst(config_rst)); 
buffer_wire buffer_9822 (.in(n9822), .out(n9822_0));
mux11 mux_4657 (.in({n14423_0, n14401_1, n14379_0/**/, n14357_0, n9903_0, n7417, n7409, n7324, n7315, n7309, n7303}), .out(n9823), .config_in(config_chain[14211:14206]), .config_rst(config_rst)); 
buffer_wire buffer_9823 (.in(n9823), .out(n9823_0));
mux13 mux_4658 (.in({n13385_2, n13365_0, n13345_0, n13325_0, n13305_0, n9690_1, n4487, n4479, n4471, n4387, n4381, n4375, n4369/**/}), .out(n9824), .config_in(config_chain[14217:14212]), .config_rst(config_rst)); 
buffer_wire buffer_9824 (.in(n9824), .out(n9824_0));
mux11 mux_4659 (.in({n14425_1, n14403_0, n14381_0/**/, n14359_0, n9905_0, n7417, n7409, n7324, n7318, n7309, n7303}), .out(n9825), .config_in(config_chain[14223:14218]), .config_rst(config_rst)); 
buffer_wire buffer_9825 (.in(n9825), .out(n9825_0));
mux13 mux_4660 (.in({n13387_2, n13367_0, n13347_1, n13327_0, n13307_1, n9698_1, n4487, n4479, n4471, n4387, n4381/**/, n4375, n4369}), .out(n9826), .config_in(config_chain[14229:14224]), .config_rst(config_rst)); 
buffer_wire buffer_9826 (.in(n9826), .out(n9826_0));
mux11 mux_4661 (.in({n14427_0, n14405_0, n14383_0, n14361_1, n9907_0, n7417, n7409, n7324, n7318, n7312, n7303}), .out(n9827), .config_in(config_chain[14235:14230]), .config_rst(config_rst)); 
buffer_wire buffer_9827 (.in(n9827), .out(n9827_0));
mux12 mux_4662 (.in({n13389_2, n13369_0, n13349_0, n13329_0, n13309_0, n9706_1, n4483, n4475, n4390, n4384, n4378/**/, n4372}), .out(n9828), .config_in(config_chain[14241:14236]), .config_rst(config_rst)); 
buffer_wire buffer_9828 (.in(n9828), .out(n9828_0));
mux11 mux_4663 (.in({n14429_0/**/, n14407_0, n14385_1, n14363_0, n9909_0, n7421, n7409, n7324, n7318, n7312, n7306}), .out(n9829), .config_in(config_chain[14247:14242]), .config_rst(config_rst)); 
buffer_wire buffer_9829 (.in(n9829), .out(n9829_0));
mux11 mux_4664 (.in({n13371_1, n13351_0, n13331_1, n13311_0, n9714_1, n4483, n4475, n4390, n4384, n4378, n4372/**/}), .out(n9830), .config_in(config_chain[14253:14248]), .config_rst(config_rst)); 
buffer_wire buffer_9830 (.in(n9830), .out(n9830_0));
mux11 mux_4665 (.in({n14431_0, n14409_1, n14387_0, n14365_0/**/, n9911_0, n7421, n7413, n7324, n7318, n7312, n7306}), .out(n9831), .config_in(config_chain[14259:14254]), .config_rst(config_rst)); 
buffer_wire buffer_9831 (.in(n9831), .out(n9831_0));
mux11 mux_4666 (.in({n13373_0, n13353_0, n13333_0, n13313_0, n9722_1, n4483, n4475, n4390/**/, n4384, n4378, n4372}), .out(n9832), .config_in(config_chain[14265:14260]), .config_rst(config_rst)); 
buffer_wire buffer_9832 (.in(n9832), .out(n9832_0));
mux11 mux_4667 (.in({n14433_2, n14411_0, n14389_0, n14367_0, n9913_0, n7421, n7413, n7405, n7318, n7312, n7306}), .out(n9833), .config_in(config_chain[14271:14266]), .config_rst(config_rst)); 
buffer_wire buffer_9833 (.in(n9833), .out(n9833_0));
mux11 mux_4668 (.in({n13375_0, n13355_1, n13335_0, n13315_1, n9730_1, n4483, n4475/**/, n4390, n4384, n4378, n4372}), .out(n9834), .config_in(config_chain[14277:14272]), .config_rst(config_rst)); 
buffer_wire buffer_9834 (.in(n9834), .out(n9834_0));
mux11 mux_4669 (.in({n14435_0, n14413_0, n14391_0, n14369_1, n9915_0, n7421, n7413, n7405, n7321, n7312, n7306}), .out(n9835), .config_in(config_chain[14283:14278]), .config_rst(config_rst)); 
buffer_wire buffer_9835 (.in(n9835), .out(n9835_0));
mux11 mux_4670 (.in({n13377_0, n13357_0, n13337_0, n13317_0, n9738_1, n4483, n4475, n4390, n4384, n4378, n4372/**/}), .out(n9836), .config_in(config_chain[14289:14284]), .config_rst(config_rst)); 
buffer_wire buffer_9836 (.in(n9836), .out(n9836_0));
mux11 mux_4671 (.in({n14437_0, n14415_0, n14393_1, n14371_0, n9917_0, n7421, n7413, n7405, n7321, n7315, n7306}), .out(n9837), .config_in(config_chain[14295:14290]), .config_rst(config_rst)); 
buffer_wire buffer_9837 (.in(n9837), .out(n9837_0));
mux13 mux_4672 (.in({n13641_0, n13621_0/**/, n13601_0, n13581_0, n13561_0, n9758_1, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9838), .config_in(config_chain[14301:14296]), .config_rst(config_rst)); 
buffer_wire buffer_9838 (.in(n9838), .out(n9838_0));
mux3 mux_4673 (.in({n14705_1, n8387, n8281}), .out(n9839), .config_in(config_chain[14303:14302]), .config_rst(config_rst)); 
buffer_wire buffer_9839 (.in(n9839), .out(n9839_0));
mux13 mux_4674 (.in({n13643_1, n13623_0, n13603_1, n13583_0, n13563_1, n9760_1, n5465, n5457, n5449/**/, n5365, n5359, n5353, n5347}), .out(n9840), .config_in(config_chain[14309:14304]), .config_rst(config_rst)); 
buffer_wire buffer_9840 (.in(n9840), .out(n9840_0));
mux3 mux_4675 (.in({n14697_2, n8391, n8284}), .out(n9841), .config_in(config_chain[14311:14310]), .config_rst(config_rst)); 
buffer_wire buffer_9841 (.in(n9841), .out(n9841_0));
mux13 mux_4676 (.in({n13645_1, n13625_0, n13605_0, n13585_0, n13565_0/**/, n9762_1, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9842), .config_in(config_chain[14317:14312]), .config_rst(config_rst)); 
buffer_wire buffer_9842 (.in(n9842), .out(n9842_0));
mux3 mux_4677 (.in({n14689_1, n8395, n8284}), .out(n9843), .config_in(config_chain[14319:14318]), .config_rst(config_rst)); 
buffer_wire buffer_9843 (.in(n9843), .out(n9843_0));
mux13 mux_4678 (.in({n13647_1, n13627_1, n13607_0, n13587_1, n13567_0, n9764_1, n5465, n5457, n5449/**/, n5365, n5359, n5353, n5347}), .out(n9844), .config_in(config_chain[14325:14320]), .config_rst(config_rst)); 
buffer_wire buffer_9844 (.in(n9844), .out(n9844_0));
mux3 mux_4679 (.in({n14681_1, n8395, n8287}), .out(n9845), .config_in(config_chain[14327:14326]), .config_rst(config_rst)); 
buffer_wire buffer_9845 (.in(n9845), .out(n9845_0));
mux13 mux_4680 (.in({n13649_2, n13629_0, n13609_0, n13589_0, n13569_0, n9766_1/**/, n5465, n5457, n5449, n5365, n5359, n5353, n5347}), .out(n9846), .config_in(config_chain[14333:14328]), .config_rst(config_rst)); 
buffer_wire buffer_9846 (.in(n9846), .out(n9846_0));
mux3 mux_4681 (.in({n14673_1, n8399, n8290}), .out(n9847), .config_in(config_chain[14335:14334]), .config_rst(config_rst)); 
buffer_wire buffer_9847 (.in(n9847), .out(n9847_0));
mux12 mux_4682 (.in({n13651_2, n13631_0, n13611_1, n13591_0, n13571_1, n9768_1, n5461, n5453/**/, n5368, n5362, n5356, n5350}), .out(n9848), .config_in(config_chain[14341:14336]), .config_rst(config_rst)); 
buffer_wire buffer_9848 (.in(n9848), .out(n9848_0));
mux2 mux_4683 (.in({n14665_1, n8293}), .out(n9849), .config_in(config_chain[14342:14342]), .config_rst(config_rst)); 
buffer_wire buffer_9849 (.in(n9849), .out(n9849_0));
mux11 mux_4684 (.in({n13633_0, n13613_0, n13593_0, n13573_0/**/, n9770_1, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9850), .config_in(config_chain[14348:14343]), .config_rst(config_rst)); 
buffer_wire buffer_9850 (.in(n9850), .out(n9850_0));
mux2 mux_4685 (.in({n14657_1, n8296}), .out(n9851), .config_in(config_chain[14349:14349]), .config_rst(config_rst)); 
buffer_wire buffer_9851 (.in(n9851), .out(n9851_0));
mux11 mux_4686 (.in({n13635_1, n13615_0, n13595_1, n13575_0, n9772_1/**/, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9852), .config_in(config_chain[14355:14350]), .config_rst(config_rst)); 
buffer_wire buffer_9852 (.in(n9852), .out(n9852_0));
mux2 mux_4687 (.in({n14649_1/**/, n8296}), .out(n9853), .config_in(config_chain[14356:14356]), .config_rst(config_rst)); 
buffer_wire buffer_9853 (.in(n9853), .out(n9853_0));
mux11 mux_4688 (.in({n13637_0/**/, n13617_0, n13597_0, n13577_0, n9774_1, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9854), .config_in(config_chain[14362:14357]), .config_rst(config_rst)); 
buffer_wire buffer_9854 (.in(n9854), .out(n9854_0));
mux2 mux_4689 (.in({n14641_1, n8299}), .out(n9855), .config_in(config_chain[14363:14363]), .config_rst(config_rst)); 
buffer_wire buffer_9855 (.in(n9855), .out(n9855_0));
mux11 mux_4690 (.in({n13639_0, n13619_1, n13599_0, n13579_1, n9776_1/**/, n5461, n5453, n5368, n5362, n5356, n5350}), .out(n9856), .config_in(config_chain[14369:14364]), .config_rst(config_rst)); 
buffer_wire buffer_9856 (.in(n9856), .out(n9856_0));
mux2 mux_4691 (.in({n14633_1, n8302}), .out(n9857), .config_in(config_chain[14370:14370]), .config_rst(config_rst)); 
buffer_wire buffer_9857 (.in(n9857), .out(n9857_0));
mux13 mux_4692 (.in({n13905_0, n13885_1, n13865_0/**/, n13845_1, n13825_0, n9778_1, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9858), .config_in(config_chain[14376:14371]), .config_rst(config_rst)); 
buffer_wire buffer_9858 (.in(n9858), .out(n9858_0));
mux3 mux_4693 (.in({n14703_0, n8387, n8281}), .out(n9859), .config_in(config_chain[14378:14377]), .config_rst(config_rst)); 
buffer_wire buffer_9859 (.in(n9859), .out(n9859_0));
mux13 mux_4694 (.in({n13907_0, n13887_0, n13867_0, n13847_0, n13827_0, n9780_1/**/, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9860), .config_in(config_chain[14384:14379]), .config_rst(config_rst)); 
buffer_wire buffer_9860 (.in(n9860), .out(n9860_0));
mux3 mux_4695 (.in({n14695_2, n8391, n8284}), .out(n9861), .config_in(config_chain[14386:14385]), .config_rst(config_rst)); 
buffer_wire buffer_9861 (.in(n9861), .out(n9861_0));
mux13 mux_4696 (.in({n13909_1, n13889_0/**/, n13869_1, n13849_0, n13829_1, n9782_1, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9862), .config_in(config_chain[14392:14387]), .config_rst(config_rst)); 
buffer_wire buffer_9862 (.in(n9862), .out(n9862_0));
mux3 mux_4697 (.in({n14687_0, n8395, n8287}), .out(n9863), .config_in(config_chain[14394:14393]), .config_rst(config_rst)); 
buffer_wire buffer_9863 (.in(n9863), .out(n9863_0));
mux13 mux_4698 (.in({n13911_1, n13891_0, n13871_0/**/, n13851_0, n13831_0, n9784_1, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9864), .config_in(config_chain[14400:14395]), .config_rst(config_rst)); 
buffer_wire buffer_9864 (.in(n9864), .out(n9864_0));
mux3 mux_4699 (.in({n14679_0/**/, n8399, n8287}), .out(n9865), .config_in(config_chain[14402:14401]), .config_rst(config_rst)); 
buffer_wire buffer_9865 (.in(n9865), .out(n9865_0));
mux13 mux_4700 (.in({n13913_1/**/, n13893_1, n13873_0, n13853_1, n13833_0, n9786_1, n6443, n6435, n6427, n6343, n6337, n6331, n6325}), .out(n9866), .config_in(config_chain[14408:14403]), .config_rst(config_rst)); 
buffer_wire buffer_9866 (.in(n9866), .out(n9866_0));
mux3 mux_4701 (.in({n14671_0, n8399, n8290}), .out(n9867), .config_in(config_chain[14410:14409]), .config_rst(config_rst)); 
buffer_wire buffer_9867 (.in(n9867), .out(n9867_0));
mux12 mux_4702 (.in({n13915_2, n13895_0, n13875_0, n13855_0/**/, n13835_0, n9788_1, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9868), .config_in(config_chain[14416:14411]), .config_rst(config_rst)); 
buffer_wire buffer_9868 (.in(n9868), .out(n9868_0));
mux2 mux_4703 (.in({n14663_0, n8293}), .out(n9869), .config_in(config_chain[14417:14417]), .config_rst(config_rst)); 
buffer_wire buffer_9869 (.in(n9869), .out(n9869_0));
mux11 mux_4704 (.in({n13897_0, n13877_1, n13857_0/**/, n13837_1, n9790_1, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9870), .config_in(config_chain[14423:14418]), .config_rst(config_rst)); 
buffer_wire buffer_9870 (.in(n9870), .out(n9870_0));
mux2 mux_4705 (.in({n14655_0, n8296}), .out(n9871), .config_in(config_chain[14424:14424]), .config_rst(config_rst)); 
buffer_wire buffer_9871 (.in(n9871), .out(n9871_0));
mux11 mux_4706 (.in({n13899_0, n13879_0, n13859_0, n13839_0, n9792_1, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9872), .config_in(config_chain[14430:14425]), .config_rst(config_rst)); 
buffer_wire buffer_9872 (.in(n9872), .out(n9872_0));
mux2 mux_4707 (.in({n14647_0, n8299}), .out(n9873), .config_in(config_chain[14431:14431]), .config_rst(config_rst)); 
buffer_wire buffer_9873 (.in(n9873), .out(n9873_0));
mux11 mux_4708 (.in({n13901_1, n13881_0/**/, n13861_1, n13841_0, n9794_1, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9874), .config_in(config_chain[14437:14432]), .config_rst(config_rst)); 
buffer_wire buffer_9874 (.in(n9874), .out(n9874_0));
mux2 mux_4709 (.in({n14639_0, n8299}), .out(n9875), .config_in(config_chain[14438:14438]), .config_rst(config_rst)); 
buffer_wire buffer_9875 (.in(n9875), .out(n9875_0));
mux11 mux_4710 (.in({n13903_0, n13883_0, n13863_0, n13843_0/**/, n9796_1, n6439, n6431, n6346, n6340, n6334, n6328}), .out(n9876), .config_in(config_chain[14444:14439]), .config_rst(config_rst)); 
buffer_wire buffer_9876 (.in(n9876), .out(n9876_0));
mux2 mux_4711 (.in({n14631_0, n8302}), .out(n9877), .config_in(config_chain[14445:14445]), .config_rst(config_rst)); 
buffer_wire buffer_9877 (.in(n9877), .out(n9877_0));
mux13 mux_4712 (.in({n14169_0, n14149_0, n14129_0/**/, n14109_0, n14089_0, n9798_1, n7421, n7413, n7405, n7321, n7315, n7309, n7303}), .out(n9878), .config_in(config_chain[14451:14446]), .config_rst(config_rst)); 
buffer_wire buffer_9878 (.in(n9878), .out(n9878_0));
mux3 mux_4713 (.in({n14701_0, n8387, n8281}), .out(n9879), .config_in(config_chain[14453:14452]), .config_rst(config_rst)); 
buffer_wire buffer_9879 (.in(n9879), .out(n9879_0));
mux13 mux_4714 (.in({n14171_0, n14151_1, n14131_0/**/, n14111_1, n14091_0, n9800_1, n7421, n7413, n7405, n7321, n7315, n7309, n7303}), .out(n9880), .config_in(config_chain[14459:14454]), .config_rst(config_rst)); 
buffer_wire buffer_9880 (.in(n9880), .out(n9880_0));
mux3 mux_4715 (.in({n14693_0, n8391, n8284}), .out(n9881), .config_in(config_chain[14461:14460]), .config_rst(config_rst)); 
buffer_wire buffer_9881 (.in(n9881), .out(n9881_0));
mux13 mux_4716 (.in({n14173_0/**/, n14153_0, n14133_0, n14113_0, n14093_0, n9802_1, n7421, n7413, n7405, n7321, n7315, n7309, n7303}), .out(n9882), .config_in(config_chain[14467:14462]), .config_rst(config_rst)); 
buffer_wire buffer_9882 (.in(n9882), .out(n9882_0));
mux3 mux_4717 (.in({n14685_0, n8395, n8287}), .out(n9883), .config_in(config_chain[14469:14468]), .config_rst(config_rst)); 
buffer_wire buffer_9883 (.in(n9883), .out(n9883_0));
mux13 mux_4718 (.in({n14175_1, n14155_0, n14135_1, n14115_0/**/, n14095_1, n9804_1, n7421, n7413, n7405, n7321, n7315, n7309, n7303}), .out(n9884), .config_in(config_chain[14475:14470]), .config_rst(config_rst)); 
buffer_wire buffer_9884 (.in(n9884), .out(n9884_0));
mux3 mux_4719 (.in({n14677_0, n8399, n8290}), .out(n9885), .config_in(config_chain[14477:14476]), .config_rst(config_rst)); 
buffer_wire buffer_9885 (.in(n9885), .out(n9885_0));
mux13 mux_4720 (.in({n14177_1, n14157_0, n14137_0, n14117_0, n14097_0/**/, n9806_1, n7421, n7413, n7405, n7321, n7315, n7309, n7303}), .out(n9886), .config_in(config_chain[14483:14478]), .config_rst(config_rst)); 
buffer_wire buffer_9886 (.in(n9886), .out(n9886_0));
mux2 mux_4721 (.in({n14669_0, n8290}), .out(n9887), .config_in(config_chain[14484:14484]), .config_rst(config_rst)); 
buffer_wire buffer_9887 (.in(n9887), .out(n9887_0));
mux12 mux_4722 (.in({n14179_1, n14159_1, n14139_0, n14119_1/**/, n14099_0, n9808_1, n7417, n7409, n7324, n7318, n7312, n7306}), .out(n9888), .config_in(config_chain[14490:14485]), .config_rst(config_rst)); 
buffer_wire buffer_9888 (.in(n9888), .out(n9888_0));
mux2 mux_4723 (.in({n14661_0/**/, n8293}), .out(n9889), .config_in(config_chain[14491:14491]), .config_rst(config_rst)); 
buffer_wire buffer_9889 (.in(n9889), .out(n9889_0));
mux11 mux_4724 (.in({n14161_0, n14141_0, n14121_0, n14101_0, n9810_1, n7417, n7409, n7324, n7318, n7312, n7306}), .out(n9890), .config_in(config_chain[14497:14492]), .config_rst(config_rst)); 
buffer_wire buffer_9890 (.in(n9890), .out(n9890_0));
mux2 mux_4725 (.in({n14653_0, n8296}), .out(n9891), .config_in(config_chain[14498:14498]), .config_rst(config_rst)); 
buffer_wire buffer_9891 (.in(n9891), .out(n9891_0));
mux11 mux_4726 (.in({n14163_0, n14143_1, n14123_0, n14103_1, n9812_1/**/, n7417, n7409, n7324, n7318, n7312, n7306}), .out(n9892), .config_in(config_chain[14504:14499]), .config_rst(config_rst)); 
buffer_wire buffer_9892 (.in(n9892), .out(n9892_0));
mux2 mux_4727 (.in({n14645_0/**/, n8299}), .out(n9893), .config_in(config_chain[14505:14505]), .config_rst(config_rst)); 
buffer_wire buffer_9893 (.in(n9893), .out(n9893_0));
mux11 mux_4728 (.in({n14165_0, n14145_0, n14125_0, n14105_0/**/, n9814_1, n7417, n7409, n7324, n7318, n7312, n7306}), .out(n9894), .config_in(config_chain[14511:14506]), .config_rst(config_rst)); 
buffer_wire buffer_9894 (.in(n9894), .out(n9894_0));
mux2 mux_4729 (.in({n14637_0, n8302}), .out(n9895), .config_in(config_chain[14512:14512]), .config_rst(config_rst)); 
buffer_wire buffer_9895 (.in(n9895), .out(n9895_0));
mux11 mux_4730 (.in({n14167_1, n14147_0, n14127_1, n14107_0, n9816_1/**/, n7417, n7409, n7324, n7318, n7312, n7306}), .out(n9896), .config_in(config_chain[14518:14513]), .config_rst(config_rst)); 
buffer_wire buffer_9896 (.in(n9896), .out(n9896_0));
mux2 mux_4731 (.in({n14629_0/**/, n8302}), .out(n9897), .config_in(config_chain[14519:14519]), .config_rst(config_rst)); 
buffer_wire buffer_9897 (.in(n9897), .out(n9897_0));
mux12 mux_4732 (.in({n14441_1, n14419_0/**/, n14397_0, n14375_0, n14353_1, n9818_1, n8395, n8383, n8299, n8293, n8287, n8281}), .out(n9898), .config_in(config_chain[14525:14520]), .config_rst(config_rst)); 
buffer_wire buffer_9898 (.in(n9898), .out(n9898_0));
mux3 mux_4733 (.in({n14615_0, n8387, n8281}), .out(n9899), .config_in(config_chain[14527:14526]), .config_rst(config_rst)); 
buffer_wire buffer_9899 (.in(n9899), .out(n9899_0));
mux12 mux_4734 (.in({n14443_1, n14421_0, n14399_0, n14377_1, n14355_0, n9820_1, n8395, n8387, n8299, n8293, n8287, n8281}), .out(n9900), .config_in(config_chain[14533:14528]), .config_rst(config_rst)); 
buffer_wire buffer_9900 (.in(n9900), .out(n9900_0));
mux3 mux_4735 (.in({n14699_0/**/, n8391, n8281}), .out(n9901), .config_in(config_chain[14535:14534]), .config_rst(config_rst)); 
buffer_wire buffer_9901 (.in(n9901), .out(n9901_0));
mux11 mux_4736 (.in({n14423_0, n14401_1, n14379_0, n14357_0, n9822_1, n8395, n8387, n8302, n8293, n8287, n8281}), .out(n9902), .config_in(config_chain[14541:14536]), .config_rst(config_rst)); 
buffer_wire buffer_9902 (.in(n9902), .out(n9902_0));
mux3 mux_4737 (.in({n14691_0, n8391, n8284}), .out(n9903), .config_in(config_chain[14543:14542]), .config_rst(config_rst)); 
buffer_wire buffer_9903 (.in(n9903), .out(n9903_0));
mux11 mux_4738 (.in({n14425_1, n14403_0, n14381_0, n14359_0, n9824_1/**/, n8395, n8387, n8302, n8296, n8287, n8281}), .out(n9904), .config_in(config_chain[14549:14544]), .config_rst(config_rst)); 
buffer_wire buffer_9904 (.in(n9904), .out(n9904_0));
mux3 mux_4739 (.in({n14683_0, n8395, n8287}), .out(n9905), .config_in(config_chain[14551:14550]), .config_rst(config_rst)); 
buffer_wire buffer_9905 (.in(n9905), .out(n9905_0));
mux11 mux_4740 (.in({n14427_0, n14405_0, n14383_0, n14361_1, n9826_1, n8395, n8387, n8302, n8296, n8290, n8281}), .out(n9906), .config_in(config_chain[14557:14552]), .config_rst(config_rst)); 
buffer_wire buffer_9906 (.in(n9906), .out(n9906_0));
mux3 mux_4741 (.in({n14675_0, n8399, n8290}), .out(n9907), .config_in(config_chain[14559:14558]), .config_rst(config_rst)); 
buffer_wire buffer_9907 (.in(n9907), .out(n9907_0));
mux11 mux_4742 (.in({n14429_0, n14407_0, n14385_1, n14363_0, n9828_1/**/, n8399, n8387, n8302, n8296, n8290, n8284}), .out(n9908), .config_in(config_chain[14565:14560]), .config_rst(config_rst)); 
buffer_wire buffer_9908 (.in(n9908), .out(n9908_0));
mux2 mux_4743 (.in({n14667_0, n8293}), .out(n9909), .config_in(config_chain[14566:14566]), .config_rst(config_rst)); 
buffer_wire buffer_9909 (.in(n9909), .out(n9909_0));
mux11 mux_4744 (.in({n14431_0, n14409_1, n14387_0, n14365_0, n9830_1/**/, n8399, n8391, n8302, n8296, n8290, n8284}), .out(n9910), .config_in(config_chain[14572:14567]), .config_rst(config_rst)); 
buffer_wire buffer_9910 (.in(n9910), .out(n9910_0));
mux2 mux_4745 (.in({n14659_0, n8293}), .out(n9911), .config_in(config_chain[14573:14573]), .config_rst(config_rst)); 
buffer_wire buffer_9911 (.in(n9911), .out(n9911_0));
mux11 mux_4746 (.in({n14433_2, n14411_0, n14389_0, n14367_0, n9832_1/**/, n8399, n8391, n8383, n8296, n8290, n8284}), .out(n9912), .config_in(config_chain[14579:14574]), .config_rst(config_rst)); 
buffer_wire buffer_9912 (.in(n9912), .out(n9912_0));
mux2 mux_4747 (.in({n14651_0, n8296}), .out(n9913), .config_in(config_chain[14580:14580]), .config_rst(config_rst)); 
buffer_wire buffer_9913 (.in(n9913), .out(n9913_0));
mux11 mux_4748 (.in({n14435_0, n14413_0/**/, n14391_0, n14369_1, n9834_1, n8399, n8391, n8383, n8299, n8290, n8284}), .out(n9914), .config_in(config_chain[14586:14581]), .config_rst(config_rst)); 
buffer_wire buffer_9914 (.in(n9914), .out(n9914_0));
mux2 mux_4749 (.in({n14643_0, n8299}), .out(n9915), .config_in(config_chain[14587:14587]), .config_rst(config_rst)); 
buffer_wire buffer_9915 (.in(n9915), .out(n9915_0));
mux11 mux_4750 (.in({n14437_0, n14415_0, n14393_1, n14371_0, n9836_1, n8399, n8391, n8383, n8299, n8293, n8284}), .out(n9916), .config_in(config_chain[14593:14588]), .config_rst(config_rst)); 
buffer_wire buffer_9916 (.in(n9916), .out(n9916_0));
mux2 mux_4751 (.in({n14635_0, n8302}), .out(n9917), .config_in(config_chain[14594:14594]), .config_rst(config_rst)); 
buffer_wire buffer_9917 (.in(n9917), .out(n9917_0));
mux10 mux_4752 (.in({n14439_0, n14417_1, n14395_0, n14373_0, n9746_2, n8391, n8383, n8299, n8293, n8287}), .out(n9918), .config_in(config_chain[14600:14595]), .config_rst(config_rst)); 
buffer_wire buffer_9918 (.in(n9918), .out(n9918_0));
mux2 mux_4753 (.in({n14627_0/**/, n8383}), .out(n9919), .config_in(config_chain[14601:14601]), .config_rst(config_rst)); 
buffer_wire buffer_9919 (.in(n9919), .out(n9919_0));
mux4 mux_4754 (.in({n12271_0, n12270_0, n673, n557}), .out(n9920), .config_in(config_chain[14603:14602]), .config_rst(config_rst)); 
buffer_wire buffer_9920 (.in(n9920), .out(n9920_0));
mux16 mux_4755 (.in({n13131_1, n13126_0, n13119_1, n13110_0, n13104_0/**/, n13093_0, n13076_0, n13067_0, n13050_0, n13041_0, n10053_1, n2625, n2617, n2529, n2521, n2513}), .out(n9921), .config_in(config_chain[14609:14604]), .config_rst(config_rst)); 
buffer_wire buffer_9921 (.in(n9921), .out(n9921_0));
mux4 mux_4756 (.in({n12363_1, n12272_0/**/, n673, n557}), .out(n9922), .config_in(config_chain[14611:14610]), .config_rst(config_rst)); 
buffer_wire buffer_9922 (.in(n9922), .out(n9922_0));
mux16 mux_4757 (.in({n13391_1, n13386_0, n13379_0, n13372_0, n13362_0, n13353_0, n13336_0, n13327_0/**/, n13310_0, n13299_0, n10073_1, n3603, n3595, n3507, n3499, n3491}), .out(n9923), .config_in(config_chain[14617:14612]), .config_rst(config_rst)); 
buffer_wire buffer_9923 (.in(n9923), .out(n9923_0));
mux4 mux_4758 (.in({n12275_0, n12274_0, n673, n557}), .out(n9924), .config_in(config_chain[14619:14618]), .config_rst(config_rst)); 
buffer_wire buffer_9924 (.in(n9924), .out(n9924_0));
mux16 mux_4759 (.in({n12617_1, n12612_0, n12605_1, n12600_0, n12588_0, n12579_0, n12562_0, n12551_0, n12534_0, n12525_0, n10013_1, n669, n661, n573, n565, n557}), .out(n9925), .config_in(config_chain[14625:14620]), .config_rst(config_rst)); 
buffer_wire buffer_9925 (.in(n9925), .out(n9925_0));
mux4 mux_4760 (.in({n12277_0, n12276_0, n673, n557}), .out(n9926), .config_in(config_chain[14627:14626]), .config_rst(config_rst)); 
buffer_wire buffer_9926 (.in(n9926), .out(n9926_0));
mux16 mux_4761 (.in({n12873_1, n12868_0, n12861_1, n12858_0, n12844_0, n12833_0, n12816_0, n12807_0, n12790_0, n12781_0, n10033_1, n1647, n1639, n1551, n1543, n1535}), .out(n9927), .config_in(config_chain[14633:14628]), .config_rst(config_rst)); 
buffer_wire buffer_9927 (.in(n9927), .out(n9927_0));
mux3 mux_4762 (.in({n12279_0, n12278_0, n557}), .out(n9928), .config_in(config_chain[14635:14634]), .config_rst(config_rst)); 
buffer_wire buffer_9928 (.in(n9928), .out(n9928_0));
mux16 mux_4763 (.in({n13149_1, n13128_0, n13121_1, n13106_0, n13097_0, n13080_0, n13069_0, n13052_0/**/, n13043_0, n13038_0, n10055_1, n2625, n2617, n2529, n2521, n2513}), .out(n9929), .config_in(config_chain[14641:14636]), .config_rst(config_rst)); 
buffer_wire buffer_9929 (.in(n9929), .out(n9929_0));
mux3 mux_4764 (.in({n12365_1/**/, n12280_0, n561}), .out(n9930), .config_in(config_chain[14643:14642]), .config_rst(config_rst)); 
buffer_wire buffer_9930 (.in(n9930), .out(n9930_0));
mux16 mux_4765 (.in({n13409_1, n13388_0, n13381_1, n13366_0, n13355_0, n13338_0, n13329_0, n13312_0, n13303_0/**/, n13300_0, n10075_1, n3603, n3595, n3507, n3499, n3491}), .out(n9931), .config_in(config_chain[14649:14644]), .config_rst(config_rst)); 
buffer_wire buffer_9931 (.in(n9931), .out(n9931_0));
mux3 mux_4766 (.in({n12283_0, n12282_0, n561}), .out(n9932), .config_in(config_chain[14651:14650]), .config_rst(config_rst)); 
buffer_wire buffer_9932 (.in(n9932), .out(n9932_0));
mux16 mux_4767 (.in({n12635_1, n12614_0, n12607_2, n12590_0/**/, n12581_0, n12564_0, n12555_0, n12538_0, n12528_0, n12527_0, n10015_1, n669, n661, n573, n565, n557}), .out(n9933), .config_in(config_chain[14657:14652]), .config_rst(config_rst)); 
buffer_wire buffer_9933 (.in(n9933), .out(n9933_0));
mux3 mux_4768 (.in({n12285_0, n12284_0, n561}), .out(n9934), .config_in(config_chain[14659:14658]), .config_rst(config_rst)); 
buffer_wire buffer_9934 (.in(n9934), .out(n9934_0));
mux16 mux_4769 (.in({n12891_1, n12870_0, n12863_1, n12846_0, n12837_0/**/, n12820_0, n12809_0, n12792_0, n12786_0, n12783_0, n10035_1, n1647, n1639, n1551, n1543, n1535}), .out(n9935), .config_in(config_chain[14665:14660]), .config_rst(config_rst)); 
buffer_wire buffer_9935 (.in(n9935), .out(n9935_0));
mux3 mux_4770 (.in({n12287_0, n12286_0, n561}), .out(n9936), .config_in(config_chain[14667:14666]), .config_rst(config_rst)); 
buffer_wire buffer_9936 (.in(n9936), .out(n9936_0));
mux15 mux_4771 (.in({n13147_1, n13123_1, n13108_0, n13099_0, n13082_0, n13073_0, n13056_0, n13046_0, n13045_0, n10057_1, n2625, n2617, n2529, n2521, n2513}), .out(n9937), .config_in(config_chain[14673:14668]), .config_rst(config_rst)); 
buffer_wire buffer_9937 (.in(n9937), .out(n9937_0));
mux3 mux_4772 (.in({n12367_1/**/, n12288_0, n561}), .out(n9938), .config_in(config_chain[14675:14674]), .config_rst(config_rst)); 
buffer_wire buffer_9938 (.in(n9938), .out(n9938_0));
mux15 mux_4773 (.in({n13407_1, n13383_1, n13368_0, n13359_0, n13342_0, n13331_0, n13314_0, n13308_0, n13305_0, n10077_1, n3603, n3595, n3507, n3499, n3491}), .out(n9939), .config_in(config_chain[14681:14676]), .config_rst(config_rst)); 
buffer_wire buffer_9939 (.in(n9939), .out(n9939_0));
mux3 mux_4774 (.in({n12291_0, n12290_0, n565}), .out(n9940), .config_in(config_chain[14683:14682]), .config_rst(config_rst)); 
buffer_wire buffer_9940 (.in(n9940), .out(n9940_0));
mux15 mux_4775 (.in({n12633_1, n12609_2, n12594_0, n12583_0, n12566_0, n12557_0, n12540_0, n12536_0, n12531_0, n10017_1, n669, n661, n573, n565, n557}), .out(n9941), .config_in(config_chain[14689:14684]), .config_rst(config_rst)); 
buffer_wire buffer_9941 (.in(n9941), .out(n9941_0));
mux3 mux_4776 (.in({n12293_0, n12292_0, n565}), .out(n9942), .config_in(config_chain[14691:14690]), .config_rst(config_rst)); 
buffer_wire buffer_9942 (.in(n9942), .out(n9942_0));
mux15 mux_4777 (.in({n12889_1, n12865_2, n12848_0, n12839_0, n12822_0, n12813_0, n12796_0, n12794_0, n12785_0, n10037_1, n1647, n1639, n1551, n1543, n1535}), .out(n9943), .config_in(config_chain[14697:14692]), .config_rst(config_rst)); 
buffer_wire buffer_9943 (.in(n9943), .out(n9943_0));
mux3 mux_4778 (.in({n12295_0, n12294_0, n565}), .out(n9944), .config_in(config_chain[14699:14698]), .config_rst(config_rst)); 
buffer_wire buffer_9944 (.in(n9944), .out(n9944_0));
mux15 mux_4779 (.in({n13145_1, n13125_2, n13112_0/**/, n13101_0, n13084_0, n13075_0, n13058_0, n13054_0, n13049_0, n10059_1, n2625, n2617, n2529, n2521, n2513}), .out(n9945), .config_in(config_chain[14705:14700]), .config_rst(config_rst)); 
buffer_wire buffer_9945 (.in(n9945), .out(n9945_0));
mux3 mux_4780 (.in({n12369_1/**/, n12296_0, n565}), .out(n9946), .config_in(config_chain[14707:14706]), .config_rst(config_rst)); 
buffer_wire buffer_9946 (.in(n9946), .out(n9946_0));
mux15 mux_4781 (.in({n13405_1, n13385_1, n13370_0, n13361_0, n13344_0, n13335_0, n13318_0, n13316_0, n13307_0, n10079_1, n3603, n3595, n3507, n3499/**/, n3491}), .out(n9947), .config_in(config_chain[14713:14708]), .config_rst(config_rst)); 
buffer_wire buffer_9947 (.in(n9947), .out(n9947_0));
mux3 mux_4782 (.in({n12299_0, n12298_0/**/, n565}), .out(n9948), .config_in(config_chain[14715:14714]), .config_rst(config_rst)); 
buffer_wire buffer_9948 (.in(n9948), .out(n9948_0));
mux15 mux_4783 (.in({n12631_1, n12611_2, n12596_0, n12587_0, n12570_0, n12559_0, n12544_0, n12542_0, n12533_0, n10019_1, n669, n661, n573, n565, n557}), .out(n9949), .config_in(config_chain[14721:14716]), .config_rst(config_rst)); 
buffer_wire buffer_9949 (.in(n9949), .out(n9949_0));
mux3 mux_4784 (.in({n12301_0, n12300_0, n569}), .out(n9950), .config_in(config_chain[14723:14722]), .config_rst(config_rst)); 
buffer_wire buffer_9950 (.in(n9950), .out(n9950_0));
mux15 mux_4785 (.in({n12887_1, n12867_2, n12852_0, n12841_0, n12824_0, n12815_0, n12802_0, n12798_0, n12789_0, n10039_1, n1647, n1639, n1551, n1543, n1535}), .out(n9951), .config_in(config_chain[14729:14724]), .config_rst(config_rst)); 
buffer_wire buffer_9951 (.in(n9951), .out(n9951_0));
mux3 mux_4786 (.in({n12303_0, n12302_0, n569}), .out(n9952), .config_in(config_chain[14731:14730]), .config_rst(config_rst)); 
buffer_wire buffer_9952 (.in(n9952), .out(n9952_0));
mux15 mux_4787 (.in({n13143_1, n13127_2, n13114_0, n13105_0/**/, n13088_0, n13077_0, n13062_0, n13060_0, n13051_0, n10061_1, n2625, n2617, n2529, n2521, n2513}), .out(n9953), .config_in(config_chain[14737:14732]), .config_rst(config_rst)); 
buffer_wire buffer_9953 (.in(n9953), .out(n9953_0));
mux3 mux_4788 (.in({n12371_1/**/, n12304_0, n569}), .out(n9954), .config_in(config_chain[14739:14738]), .config_rst(config_rst)); 
buffer_wire buffer_9954 (.in(n9954), .out(n9954_0));
mux15 mux_4789 (.in({n13403_1, n13387_2, n13374_0, n13363_0, n13346_0, n13337_0, n13324_0, n13320_0, n13311_0, n10081_1, n3603, n3595, n3507, n3499, n3491}), .out(n9955), .config_in(config_chain[14745:14740]), .config_rst(config_rst)); 
buffer_wire buffer_9955 (.in(n9955), .out(n9955_0));
mux3 mux_4790 (.in({n12307_0, n12306_0, n569}), .out(n9956), .config_in(config_chain[14747:14746]), .config_rst(config_rst)); 
buffer_wire buffer_9956 (.in(n9956), .out(n9956_0));
mux15 mux_4791 (.in({n12629_1, n12613_2, n12598_0, n12589_0/**/, n12572_0, n12563_0, n12552_0, n12546_0, n12535_0, n10021_1, n669, n661, n573, n565, n557}), .out(n9957), .config_in(config_chain[14753:14748]), .config_rst(config_rst)); 
buffer_wire buffer_9957 (.in(n9957), .out(n9957_0));
mux3 mux_4792 (.in({n12309_0, n12308_0, n569}), .out(n9958), .config_in(config_chain[14755:14754]), .config_rst(config_rst)); 
buffer_wire buffer_9958 (.in(n9958), .out(n9958_0));
mux15 mux_4793 (.in({n12885_1, n12869_2, n12854_0, n12845_0/**/, n12828_0, n12817_0, n12810_0, n12800_0, n12791_0, n10041_1, n1647, n1639, n1551, n1543, n1535}), .out(n9959), .config_in(config_chain[14761:14756]), .config_rst(config_rst)); 
buffer_wire buffer_9959 (.in(n9959), .out(n9959_0));
mux3 mux_4794 (.in({n12311_0, n12310_0, n573}), .out(n9960), .config_in(config_chain[14763:14762]), .config_rst(config_rst)); 
buffer_wire buffer_9960 (.in(n9960), .out(n9960_0));
mux15 mux_4795 (.in({n13141_1, n13129_2, n13116_0, n13107_0, n13090_0, n13081_0, n13070_0, n13064_0, n13053_0, n10063_1, n2629, n2621, n2613, n2525, n2517}), .out(n9961), .config_in(config_chain[14769:14764]), .config_rst(config_rst)); 
buffer_wire buffer_9961 (.in(n9961), .out(n9961_0));
mux3 mux_4796 (.in({n12373_1, n12312_0, n573}), .out(n9962), .config_in(config_chain[14771:14770]), .config_rst(config_rst)); 
buffer_wire buffer_9962 (.in(n9962), .out(n9962_0));
mux15 mux_4797 (.in({n13401_1, n13389_2, n13376_0, n13367_0, n13350_0, n13339_0, n13332_0/**/, n13322_0, n13313_0, n10083_1, n3607, n3599, n3591, n3503, n3495}), .out(n9963), .config_in(config_chain[14777:14772]), .config_rst(config_rst)); 
buffer_wire buffer_9963 (.in(n9963), .out(n9963_0));
mux3 mux_4798 (.in({n12315_0, n12314_0, n573}), .out(n9964), .config_in(config_chain[14779:14778]), .config_rst(config_rst)); 
buffer_wire buffer_9964 (.in(n9964), .out(n9964_0));
mux15 mux_4799 (.in({n12627_1, n12615_2, n12602_0, n12591_0, n12574_0, n12565_0, n12560_0, n12548_0, n12539_0, n10023_1, n673, n665, n657, n569, n561}), .out(n9965), .config_in(config_chain[14785:14780]), .config_rst(config_rst)); 
buffer_wire buffer_9965 (.in(n9965), .out(n9965_0));
mux3 mux_4800 (.in({n12317_0, n12316_0, n573}), .out(n9966), .config_in(config_chain[14787:14786]), .config_rst(config_rst)); 
buffer_wire buffer_9966 (.in(n9966), .out(n9966_0));
mux15 mux_4801 (.in({n12883_1, n12871_2, n12856_0, n12847_0, n12830_0, n12821_0, n12818_0, n12804_0, n12793_0, n10043_1, n1651, n1643, n1635, n1547, n1539}), .out(n9967), .config_in(config_chain[14793:14788]), .config_rst(config_rst)); 
buffer_wire buffer_9967 (.in(n9967), .out(n9967_0));
mux3 mux_4802 (.in({n12319_0/**/, n12318_0, n573}), .out(n9968), .config_in(config_chain[14795:14794]), .config_rst(config_rst)); 
buffer_wire buffer_9968 (.in(n9968), .out(n9968_0));
mux15 mux_4803 (.in({n13139_1, n13118_0, n13109_0, n13092_0, n13083_0, n13078_0, n13066_0, n13057_0, n13040_0, n10065_1, n2629, n2621, n2613, n2525, n2517/**/}), .out(n9969), .config_in(config_chain[14801:14796]), .config_rst(config_rst)); 
buffer_wire buffer_9969 (.in(n9969), .out(n9969_0));
mux3 mux_4804 (.in({n12375_1/**/, n12320_0, n657}), .out(n9970), .config_in(config_chain[14803:14802]), .config_rst(config_rst)); 
buffer_wire buffer_9970 (.in(n9970), .out(n9970_0));
mux15 mux_4805 (.in({n13399_1, n13378_0, n13369_0, n13352_0, n13343_0, n13340_0, n13326_0, n13315_0/**/, n13298_0, n10085_1, n3607, n3599, n3591, n3503, n3495}), .out(n9971), .config_in(config_chain[14809:14804]), .config_rst(config_rst)); 
buffer_wire buffer_9971 (.in(n9971), .out(n9971_0));
mux3 mux_4806 (.in({n12323_0, n12322_0, n657}), .out(n9972), .config_in(config_chain[14811:14810]), .config_rst(config_rst)); 
buffer_wire buffer_9972 (.in(n9972), .out(n9972_0));
mux15 mux_4807 (.in({n12625_1, n12604_0, n12595_0, n12578_0, n12568_0, n12567_0, n12550_0, n12541_0, n12524_0, n10025_1, n673, n665, n657, n569, n561}), .out(n9973), .config_in(config_chain[14817:14812]), .config_rst(config_rst)); 
buffer_wire buffer_9973 (.in(n9973), .out(n9973_0));
mux3 mux_4808 (.in({n12325_0, n12324_0, n657}), .out(n9974), .config_in(config_chain[14819:14818]), .config_rst(config_rst)); 
buffer_wire buffer_9974 (.in(n9974), .out(n9974_0));
mux15 mux_4809 (.in({n12881_1, n12860_0, n12849_0, n12832_0, n12826_0, n12823_0, n12806_0, n12797_0/**/, n12780_0, n10045_1, n1651, n1643, n1635, n1547, n1539}), .out(n9975), .config_in(config_chain[14825:14820]), .config_rst(config_rst)); 
buffer_wire buffer_9975 (.in(n9975), .out(n9975_0));
mux3 mux_4810 (.in({n12327_0/**/, n12326_0, n657}), .out(n9976), .config_in(config_chain[14827:14826]), .config_rst(config_rst)); 
buffer_wire buffer_9976 (.in(n9976), .out(n9976_0));
mux15 mux_4811 (.in({n13137_1, n13120_0, n13113_0, n13096_0, n13086_0, n13085_0, n13068_0, n13059_0, n13042_0, n10067_1, n2629, n2621, n2613, n2525, n2517/**/}), .out(n9977), .config_in(config_chain[14833:14828]), .config_rst(config_rst)); 
buffer_wire buffer_9977 (.in(n9977), .out(n9977_0));
mux3 mux_4812 (.in({n12377_1/**/, n12328_0, n657}), .out(n9978), .config_in(config_chain[14835:14834]), .config_rst(config_rst)); 
buffer_wire buffer_9978 (.in(n9978), .out(n9978_0));
mux15 mux_4813 (.in({n13397_1, n13380_0, n13371_0, n13354_0, n13348_0, n13345_0, n13328_0, n13319_0, n13302_0, n10087_1, n3607, n3599, n3591, n3503, n3495}), .out(n9979), .config_in(config_chain[14841:14836]), .config_rst(config_rst)); 
buffer_wire buffer_9979 (.in(n9979), .out(n9979_0));
mux3 mux_4814 (.in({n12331_0, n12330_0, n661}), .out(n9980), .config_in(config_chain[14843:14842]), .config_rst(config_rst)); 
buffer_wire buffer_9980 (.in(n9980), .out(n9980_0));
mux15 mux_4815 (.in({n12623_1, n12606_0, n12597_0, n12580_0, n12576_0, n12571_0, n12554_0, n12543_0, n12526_0, n10027_1, n673, n665, n657, n569, n561}), .out(n9981), .config_in(config_chain[14849:14844]), .config_rst(config_rst)); 
buffer_wire buffer_9981 (.in(n9981), .out(n9981_0));
mux3 mux_4816 (.in({n12333_0, n12332_0, n661}), .out(n9982), .config_in(config_chain[14851:14850]), .config_rst(config_rst)); 
buffer_wire buffer_9982 (.in(n9982), .out(n9982_0));
mux15 mux_4817 (.in({n12879_1, n12862_0, n12853_0, n12836_0, n12834_0, n12825_0, n12808_0, n12799_0, n12782_0, n10047_1, n1651, n1643, n1635, n1547, n1539}), .out(n9983), .config_in(config_chain[14857:14852]), .config_rst(config_rst)); 
buffer_wire buffer_9983 (.in(n9983), .out(n9983_0));
mux3 mux_4818 (.in({n12335_0/**/, n12334_0, n661}), .out(n9984), .config_in(config_chain[14859:14858]), .config_rst(config_rst)); 
buffer_wire buffer_9984 (.in(n9984), .out(n9984_0));
mux15 mux_4819 (.in({n13135_1, n13122_0, n13115_0, n13098_0, n13094_0, n13089_0, n13072_0, n13061_0, n13044_0, n10069_1, n2629, n2621, n2613, n2525, n2517/**/}), .out(n9985), .config_in(config_chain[14865:14860]), .config_rst(config_rst)); 
buffer_wire buffer_9985 (.in(n9985), .out(n9985_0));
mux3 mux_4820 (.in({n12379_1/**/, n12336_0, n661}), .out(n9986), .config_in(config_chain[14867:14866]), .config_rst(config_rst)); 
buffer_wire buffer_9986 (.in(n9986), .out(n9986_0));
mux15 mux_4821 (.in({n13395_1, n13382_0, n13375_0, n13358_0, n13356_0, n13347_0, n13330_0, n13321_0, n13304_0, n10089_1, n3607, n3599/**/, n3591, n3503, n3495}), .out(n9987), .config_in(config_chain[14873:14868]), .config_rst(config_rst)); 
buffer_wire buffer_9987 (.in(n9987), .out(n9987_0));
mux3 mux_4822 (.in({n12339_0, n12338_0, n661}), .out(n9988), .config_in(config_chain[14875:14874]), .config_rst(config_rst)); 
buffer_wire buffer_9988 (.in(n9988), .out(n9988_0));
mux15 mux_4823 (.in({n12621_1, n12608_0, n12599_0, n12584_0, n12582_0, n12573_0, n12556_0, n12547_0, n12530_0, n10029_1, n673, n665, n657, n569, n561}), .out(n9989), .config_in(config_chain[14881:14876]), .config_rst(config_rst)); 
buffer_wire buffer_9989 (.in(n9989), .out(n9989_0));
mux3 mux_4824 (.in({n12341_0, n12340_0, n665}), .out(n9990), .config_in(config_chain[14883:14882]), .config_rst(config_rst)); 
buffer_wire buffer_9990 (.in(n9990), .out(n9990_0));
mux15 mux_4825 (.in({n12877_1, n12864_0, n12855_0, n12842_0, n12838_0, n12829_0, n12812_0, n12801_0, n12784_0, n10049_1, n1651, n1643, n1635, n1547, n1539}), .out(n9991), .config_in(config_chain[14889:14884]), .config_rst(config_rst)); 
buffer_wire buffer_9991 (.in(n9991), .out(n9991_0));
mux3 mux_4826 (.in({n12343_0/**/, n12342_0, n665}), .out(n9992), .config_in(config_chain[14891:14890]), .config_rst(config_rst)); 
buffer_wire buffer_9992 (.in(n9992), .out(n9992_0));
mux15 mux_4827 (.in({n13133_1, n13124_0, n13117_0, n13102_0, n13100_0, n13091_0, n13074_0, n13065_0, n13048_0, n10071_1, n2629, n2621/**/, n2613, n2525, n2517}), .out(n9993), .config_in(config_chain[14897:14892]), .config_rst(config_rst)); 
buffer_wire buffer_9993 (.in(n9993), .out(n9993_0));
mux3 mux_4828 (.in({n12381_1/**/, n12344_0, n665}), .out(n9994), .config_in(config_chain[14899:14898]), .config_rst(config_rst)); 
buffer_wire buffer_9994 (.in(n9994), .out(n9994_0));
mux15 mux_4829 (.in({n13393_1, n13384_0, n13377_0, n13364_0, n13360_0, n13351_0, n13334_0, n13323_0, n13306_0, n10091_1, n3607, n3599, n3591, n3503, n3495}), .out(n9995), .config_in(config_chain[14905:14900]), .config_rst(config_rst)); 
buffer_wire buffer_9995 (.in(n9995), .out(n9995_0));
mux3 mux_4830 (.in({n12347_0, n12346_0, n665}), .out(n9996), .config_in(config_chain[14907:14906]), .config_rst(config_rst)); 
buffer_wire buffer_9996 (.in(n9996), .out(n9996_0));
mux15 mux_4831 (.in({n12619_1, n12610_0, n12603_0, n12592_0, n12586_0, n12575_0, n12558_0, n12549_0, n12532_0, n10031_1, n673, n665, n657, n569, n561}), .out(n9997), .config_in(config_chain[14913:14908]), .config_rst(config_rst)); 
buffer_wire buffer_9997 (.in(n9997), .out(n9997_0));
mux3 mux_4832 (.in({n12349_0, n12348_0, n665}), .out(n9998), .config_in(config_chain[14915:14914]), .config_rst(config_rst)); 
buffer_wire buffer_9998 (.in(n9998), .out(n9998_0));
mux15 mux_4833 (.in({n12875_1, n12866_0, n12857_0, n12850_0, n12840_0, n12831_0, n12814_0/**/, n12805_0, n12788_0, n10051_1, n1651, n1643, n1635, n1547, n1539}), .out(n9999), .config_in(config_chain[14921:14916]), .config_rst(config_rst)); 
buffer_wire buffer_9999 (.in(n9999), .out(n9999_0));
mux3 mux_4834 (.in({n12351_2, n12350_0, n669}), .out(n10000), .config_in(config_chain[14923:14922]), .config_rst(config_rst)); 
buffer_wire buffer_10000 (.in(n10000), .out(n10000_0));
mux13 mux_4835 (.in({n14183_1, n14175_0/**/, n14170_0, n14160_0, n14147_0, n14140_0, n14117_0, n14110_0, n10153_0, n6537, n6529, n6441, n6433}), .out(n10001), .config_in(config_chain[14929:14924]), .config_rst(config_rst)); 
buffer_wire buffer_10001 (.in(n10001), .out(n10001_0));
mux3 mux_4836 (.in({n12353_2, n12352_0, n669}), .out(n10002), .config_in(config_chain[14931:14930]), .config_rst(config_rst)); 
buffer_wire buffer_10002 (.in(n10002), .out(n10002_0));
mux13 mux_4837 (.in({n14447_1, n14439_0, n14432_0, n14426_0, n14409_0, n14404_0, n14381_0, n14374_0/**/, n10175_0, n7515, n7507, n7419, n7411}), .out(n10003), .config_in(config_chain[14937:14932]), .config_rst(config_rst)); 
buffer_wire buffer_10003 (.in(n10003), .out(n10003_0));
mux3 mux_4838 (.in({n12355_2, n12354_0, n669}), .out(n10004), .config_in(config_chain[14939:14938]), .config_rst(config_rst)); 
buffer_wire buffer_10004 (.in(n10004), .out(n10004_0));
mux3 mux_4839 (.in({n14727_2, n14698_0, n8493}), .out(n10005), .config_in(config_chain[14941:14940]), .config_rst(config_rst)); 
buffer_wire buffer_10005 (.in(n10005), .out(n10005_0));
mux3 mux_4840 (.in({n12357_2, n12356_0, n669}), .out(n10006), .config_in(config_chain[14943:14942]), .config_rst(config_rst)); 
buffer_wire buffer_10006 (.in(n10006), .out(n10006_0));
mux3 mux_4841 (.in({n14701_0, n14700_0, n8493}), .out(n10007), .config_in(config_chain[14945:14944]), .config_rst(config_rst)); 
buffer_wire buffer_10007 (.in(n10007), .out(n10007_0));
mux3 mux_4842 (.in({n12359_2, n12358_0, n669}), .out(n10008), .config_in(config_chain[14947:14946]), .config_rst(config_rst)); 
buffer_wire buffer_10008 (.in(n10008), .out(n10008_0));
mux3 mux_4843 (.in({n14703_0, n14702_0, n8493}), .out(n10009), .config_in(config_chain[14949:14948]), .config_rst(config_rst)); 
buffer_wire buffer_10009 (.in(n10009), .out(n10009_0));
mux3 mux_4844 (.in({n12361_2, n12360_0, n673}), .out(n10010), .config_in(config_chain[14951:14950]), .config_rst(config_rst)); 
buffer_wire buffer_10010 (.in(n10010), .out(n10010_0));
mux3 mux_4845 (.in({n14705_0, n14704_0, n8497}), .out(n10011), .config_in(config_chain[14953:14952]), .config_rst(config_rst)); 
buffer_wire buffer_10011 (.in(n10011), .out(n10011_0));
mux16 mux_4846 (.in({n12635_1, n12613_2, n12604_0, n12592_0, n12589_0, n12578_0, n12563_0, n12550_0, n12535_0, n12524_0, n9924_0, n1647, n1639, n1551, n1543, n1535}), .out(n10012), .config_in(config_chain[14959:14954]), .config_rst(config_rst)); 
buffer_wire buffer_10012 (.in(n10012), .out(n10012_0));
mux16 mux_4847 (.in({n13653_1, n13648_0, n13641_0, n13636_0, n13624_0, n13615_0, n13598_0, n13587_0, n13570_0, n13561_0, n10093_1/**/, n4581, n4573, n4485, n4477, n4469}), .out(n10013), .config_in(config_chain[14965:14960]), .config_rst(config_rst)); 
buffer_wire buffer_10013 (.in(n10013), .out(n10013_0));
mux16 mux_4848 (.in({n12617_1, n12615_2, n12606_0, n12591_0, n12584_0, n12580_0, n12565_0, n12554_0, n12539_0, n12526_0, n9932_0, n1647, n1639, n1551, n1543, n1535}), .out(n10014), .config_in(config_chain[14971:14966]), .config_rst(config_rst)); 
buffer_wire buffer_10014 (.in(n10014), .out(n10014_0));
mux16 mux_4849 (.in({n13671_1, n13650_0, n13643_0, n13626_0, n13617_0, n13600_0, n13591_0, n13574_0, n13564_0, n13563_0, n10095_1/**/, n4581, n4573, n4485, n4477, n4469}), .out(n10015), .config_in(config_chain[14977:14972]), .config_rst(config_rst)); 
buffer_wire buffer_10015 (.in(n10015), .out(n10015_0));
mux15 mux_4850 (.in({n12619_1, n12608_0, n12595_0, n12582_0, n12576_0, n12567_0, n12556_0/**/, n12541_0, n12530_0, n9940_0, n1647, n1639, n1551, n1543, n1535}), .out(n10016), .config_in(config_chain[14983:14978]), .config_rst(config_rst)); 
buffer_wire buffer_10016 (.in(n10016), .out(n10016_0));
mux15 mux_4851 (.in({n13669_1, n13645_1, n13630_0, n13619_0, n13602_0, n13593_0, n13576_0, n13572_0, n13567_0, n10097_1/**/, n4581, n4573, n4485, n4477, n4469}), .out(n10017), .config_in(config_chain[14989:14984]), .config_rst(config_rst)); 
buffer_wire buffer_10017 (.in(n10017), .out(n10017_0));
mux15 mux_4852 (.in({n12621_1, n12610_0, n12597_0, n12586_0, n12571_0/**/, n12568_0, n12558_0, n12543_0, n12532_0, n9948_0, n1647, n1639, n1551, n1543, n1535}), .out(n10018), .config_in(config_chain[14995:14990]), .config_rst(config_rst)); 
buffer_wire buffer_10018 (.in(n10018), .out(n10018_0));
mux15 mux_4853 (.in({n13667_1, n13647_1, n13632_0, n13623_0, n13606_0, n13595_0, n13580_0, n13578_0, n13569_0, n10099_1, n4581/**/, n4573, n4485, n4477, n4469}), .out(n10019), .config_in(config_chain[15001:14996]), .config_rst(config_rst)); 
buffer_wire buffer_10019 (.in(n10019), .out(n10019_0));
mux15 mux_4854 (.in({n12623_1, n12612_0, n12599_0, n12588_0, n12573_0, n12562_0, n12560_0, n12547_0, n12534_0, n9956_0, n1647, n1639, n1551, n1543, n1535}), .out(n10020), .config_in(config_chain[15007:15002]), .config_rst(config_rst)); 
buffer_wire buffer_10020 (.in(n10020), .out(n10020_0));
mux15 mux_4855 (.in({n13665_1, n13649_1, n13634_0, n13625_0, n13608_0, n13599_0, n13588_0, n13582_0, n13571_0, n10101_1/**/, n4581, n4573, n4485, n4477, n4469}), .out(n10021), .config_in(config_chain[15013:15008]), .config_rst(config_rst)); 
buffer_wire buffer_10021 (.in(n10021), .out(n10021_0));
mux15 mux_4856 (.in({n12625_1, n12614_0, n12603_0, n12590_0, n12575_0, n12564_0, n12552_0/**/, n12549_0, n12538_0, n9964_0, n1651, n1643, n1635, n1547, n1539}), .out(n10022), .config_in(config_chain[15019:15014]), .config_rst(config_rst)); 
buffer_wire buffer_10022 (.in(n10022), .out(n10022_0));
mux15 mux_4857 (.in({n13663_1, n13651_2, n13638_0/**/, n13627_0, n13610_0, n13601_0, n13596_0, n13584_0, n13575_0, n10103_1, n4585, n4577, n4569, n4481, n4473}), .out(n10023), .config_in(config_chain[15025:15020]), .config_rst(config_rst)); 
buffer_wire buffer_10023 (.in(n10023), .out(n10023_0));
mux15 mux_4858 (.in({n12627_1, n12605_1, n12594_0, n12579_0, n12566_0/**/, n12551_0, n12544_0, n12540_0, n12525_0, n9972_0, n1651, n1643, n1635, n1547, n1539}), .out(n10024), .config_in(config_chain[15031:15026]), .config_rst(config_rst)); 
buffer_wire buffer_10024 (.in(n10024), .out(n10024_0));
mux15 mux_4859 (.in({n13661_1/**/, n13640_0, n13631_0, n13614_0, n13604_0, n13603_0, n13586_0, n13577_0, n13560_0, n10105_1, n4585, n4577, n4569, n4481, n4473}), .out(n10025), .config_in(config_chain[15037:15032]), .config_rst(config_rst)); 
buffer_wire buffer_10025 (.in(n10025), .out(n10025_0));
mux15 mux_4860 (.in({n12629_1, n12607_2, n12596_0, n12581_0, n12570_0, n12555_0, n12542_0, n12536_0/**/, n12527_0, n9980_0, n1651, n1643, n1635, n1547, n1539}), .out(n10026), .config_in(config_chain[15043:15038]), .config_rst(config_rst)); 
buffer_wire buffer_10026 (.in(n10026), .out(n10026_0));
mux15 mux_4861 (.in({n13659_1, n13642_0, n13633_0/**/, n13616_0, n13612_0, n13607_0, n13590_0, n13579_0, n13562_0, n10107_1, n4585, n4577, n4569, n4481, n4473}), .out(n10027), .config_in(config_chain[15049:15044]), .config_rst(config_rst)); 
buffer_wire buffer_10027 (.in(n10027), .out(n10027_0));
mux15 mux_4862 (.in({n12631_1, n12609_2, n12598_0, n12583_0/**/, n12572_0, n12557_0, n12546_0, n12531_0, n12528_0, n9988_0, n1651, n1643, n1635, n1547, n1539}), .out(n10028), .config_in(config_chain[15055:15050]), .config_rst(config_rst)); 
buffer_wire buffer_10028 (.in(n10028), .out(n10028_0));
mux15 mux_4863 (.in({n13657_1, n13644_0, n13635_0, n13620_0, n13618_0, n13609_0, n13592_0, n13583_0, n13566_0, n10109_1, n4585, n4577/**/, n4569, n4481, n4473}), .out(n10029), .config_in(config_chain[15061:15056]), .config_rst(config_rst)); 
buffer_wire buffer_10029 (.in(n10029), .out(n10029_0));
mux15 mux_4864 (.in({n12633_1/**/, n12611_2, n12602_0, n12600_0, n12587_0, n12574_0, n12559_0, n12548_0, n12533_0, n9996_0, n1651, n1643, n1635, n1547, n1539}), .out(n10030), .config_in(config_chain[15067:15062]), .config_rst(config_rst)); 
buffer_wire buffer_10030 (.in(n10030), .out(n10030_0));
mux15 mux_4865 (.in({n13655_1, n13646_0, n13639_0, n13628_0, n13622_0, n13611_0, n13594_0, n13585_0, n13568_0/**/, n10111_1, n4585, n4577, n4569, n4481, n4473}), .out(n10031), .config_in(config_chain[15073:15068]), .config_rst(config_rst)); 
buffer_wire buffer_10031 (.in(n10031), .out(n10031_0));
mux16 mux_4866 (.in({n12891_1, n12869_2, n12860_0, n12850_0, n12845_0, n12832_0, n12817_0, n12806_0, n12791_0, n12780_0, n9926_0, n2625/**/, n2617, n2529, n2521, n2513}), .out(n10032), .config_in(config_chain[15079:15074]), .config_rst(config_rst)); 
buffer_wire buffer_10032 (.in(n10032), .out(n10032_0));
mux16 mux_4867 (.in({n13917_1, n13912_0, n13905_0, n13902_0, n13888_0, n13877_0, n13860_0, n13851_0, n13834_0, n13825_0, n10113_0, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10033), .config_in(config_chain[15085:15080]), .config_rst(config_rst)); 
buffer_wire buffer_10033 (.in(n10033), .out(n10033_0));
mux16 mux_4868 (.in({n12873_1/**/, n12871_2, n12862_0, n12847_0, n12842_0, n12836_0, n12821_0, n12808_0, n12793_0, n12782_0, n9934_0, n2625, n2617, n2529, n2521, n2513}), .out(n10034), .config_in(config_chain[15091:15086]), .config_rst(config_rst)); 
buffer_wire buffer_10034 (.in(n10034), .out(n10034_0));
mux16 mux_4869 (.in({n13935_1, n13914_0, n13907_0, n13890_0, n13881_0, n13864_0, n13853_0, n13836_0, n13830_0, n13827_0, n10115_0, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10035), .config_in(config_chain[15097:15092]), .config_rst(config_rst)); 
buffer_wire buffer_10035 (.in(n10035), .out(n10035_0));
mux15 mux_4870 (.in({n12875_1, n12864_0, n12849_0/**/, n12838_0, n12834_0, n12823_0, n12812_0, n12797_0, n12784_0, n9942_0, n2625, n2617, n2529, n2521, n2513}), .out(n10036), .config_in(config_chain[15103:15098]), .config_rst(config_rst)); 
buffer_wire buffer_10036 (.in(n10036), .out(n10036_0));
mux15 mux_4871 (.in({n13933_1, n13909_0, n13892_0, n13883_0, n13866_0, n13857_0, n13840_0, n13838_0, n13829_0, n10117_0, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10037), .config_in(config_chain[15109:15104]), .config_rst(config_rst)); 
buffer_wire buffer_10037 (.in(n10037), .out(n10037_0));
mux15 mux_4872 (.in({n12877_1, n12866_0, n12853_0/**/, n12840_0, n12826_0, n12825_0, n12814_0, n12799_0, n12788_0, n9950_0, n2625, n2617, n2529, n2521, n2513}), .out(n10038), .config_in(config_chain[15115:15110]), .config_rst(config_rst)); 
buffer_wire buffer_10038 (.in(n10038), .out(n10038_0));
mux15 mux_4873 (.in({n13931_1, n13911_1, n13896_0, n13885_0, n13868_0, n13859_0, n13846_0, n13842_0, n13833_0, n10119_0, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10039), .config_in(config_chain[15121:15116]), .config_rst(config_rst)); 
buffer_wire buffer_10039 (.in(n10039), .out(n10039_0));
mux15 mux_4874 (.in({n12879_1, n12868_0, n12855_0, n12844_0, n12829_0, n12818_0, n12816_0, n12801_0, n12790_0/**/, n9958_0, n2625, n2617, n2529, n2521, n2513}), .out(n10040), .config_in(config_chain[15127:15122]), .config_rst(config_rst)); 
buffer_wire buffer_10040 (.in(n10040), .out(n10040_0));
mux15 mux_4875 (.in({n13929_1, n13913_1, n13898_0, n13889_0, n13872_0/**/, n13861_0, n13854_0, n13844_0, n13835_0, n10121_0, n5559, n5551, n5463, n5455, n5447}), .out(n10041), .config_in(config_chain[15133:15128]), .config_rst(config_rst)); 
buffer_wire buffer_10041 (.in(n10041), .out(n10041_0));
mux15 mux_4876 (.in({n12881_1, n12870_0, n12857_0, n12846_0, n12831_0, n12820_0, n12810_0, n12805_0, n12792_0, n9966_0, n2629, n2621, n2613, n2525, n2517}), .out(n10042), .config_in(config_chain[15139:15134]), .config_rst(config_rst)); 
buffer_wire buffer_10042 (.in(n10042), .out(n10042_0));
mux15 mux_4877 (.in({n13927_1, n13915_1, n13900_0, n13891_0, n13874_0, n13865_0, n13862_0, n13848_0/**/, n13837_0, n10123_0, n5563, n5555, n5547, n5459, n5451}), .out(n10043), .config_in(config_chain[15145:15140]), .config_rst(config_rst)); 
buffer_wire buffer_10043 (.in(n10043), .out(n10043_0));
mux15 mux_4878 (.in({n12883_1, n12861_1, n12848_0, n12833_0, n12822_0, n12807_0, n12802_0, n12796_0, n12781_0/**/, n9974_0, n2629, n2621, n2613, n2525, n2517}), .out(n10044), .config_in(config_chain[15151:15146]), .config_rst(config_rst)); 
buffer_wire buffer_10044 (.in(n10044), .out(n10044_0));
mux15 mux_4879 (.in({n13925_1, n13904_0, n13893_0, n13876_0, n13870_0, n13867_0/**/, n13850_0, n13841_0, n13824_0, n10125_0, n5563, n5555, n5547, n5459, n5451}), .out(n10045), .config_in(config_chain[15157:15152]), .config_rst(config_rst)); 
buffer_wire buffer_10045 (.in(n10045), .out(n10045_0));
mux15 mux_4880 (.in({n12885_1, n12863_1, n12852_0, n12837_0, n12824_0, n12809_0, n12798_0, n12794_0, n12783_0/**/, n9982_0, n2629, n2621, n2613, n2525, n2517}), .out(n10046), .config_in(config_chain[15163:15158]), .config_rst(config_rst)); 
buffer_wire buffer_10046 (.in(n10046), .out(n10046_0));
mux15 mux_4881 (.in({n13923_1, n13906_0, n13897_0/**/, n13880_0, n13878_0, n13869_0, n13852_0, n13843_0, n13826_0, n10127_0, n5563, n5555, n5547, n5459, n5451}), .out(n10047), .config_in(config_chain[15169:15164]), .config_rst(config_rst)); 
buffer_wire buffer_10047 (.in(n10047), .out(n10047_0));
mux15 mux_4882 (.in({n12887_1, n12865_2, n12854_0, n12839_0, n12828_0, n12813_0, n12800_0, n12786_0/**/, n12785_0, n9990_0, n2629, n2621, n2613, n2525, n2517}), .out(n10048), .config_in(config_chain[15175:15170]), .config_rst(config_rst)); 
buffer_wire buffer_10048 (.in(n10048), .out(n10048_0));
mux15 mux_4883 (.in({n13921_1, n13908_0, n13899_0, n13886_0, n13882_0, n13873_0, n13856_0, n13845_0, n13828_0, n10129_0, n5563, n5555, n5547, n5459, n5451}), .out(n10049), .config_in(config_chain[15181:15176]), .config_rst(config_rst)); 
buffer_wire buffer_10049 (.in(n10049), .out(n10049_0));
mux15 mux_4884 (.in({n12889_1, n12867_2, n12858_0, n12856_0, n12841_0, n12830_0, n12815_0, n12804_0, n12789_0, n9998_0, n2629, n2621, n2613/**/, n2525, n2517}), .out(n10050), .config_in(config_chain[15187:15182]), .config_rst(config_rst)); 
buffer_wire buffer_10050 (.in(n10050), .out(n10050_0));
mux15 mux_4885 (.in({n13919_1, n13910_0, n13901_0, n13894_0, n13884_0, n13875_0, n13858_0, n13849_0/**/, n13832_0, n10131_0, n5563, n5555, n5547, n5459, n5451}), .out(n10051), .config_in(config_chain[15193:15188]), .config_rst(config_rst)); 
buffer_wire buffer_10051 (.in(n10051), .out(n10051_0));
mux16 mux_4886 (.in({n13149_1, n13127_2, n13118_0, n13105_0, n13102_0, n13092_0, n13077_0, n13066_0, n13051_0, n13040_0, n9920_0, n3603, n3595, n3507, n3499/**/, n3491}), .out(n10052), .config_in(config_chain[15199:15194]), .config_rst(config_rst)); 
buffer_wire buffer_10052 (.in(n10052), .out(n10052_0));
mux15 mux_4887 (.in({n14181_1, n14177_1, n14172_0, n14168_0, n14149_0, n14142_0, n14119_0, n14114_0, n14091_0, n10133_0, n6537/**/, n6529, n6441, n6433, n6425}), .out(n10053), .config_in(config_chain[15205:15200]), .config_rst(config_rst)); 
buffer_wire buffer_10053 (.in(n10053), .out(n10053_0));
mux16 mux_4888 (.in({n13131_1, n13129_2, n13120_0, n13107_0, n13096_0, n13094_0, n13081_0/**/, n13068_0, n13053_0, n13042_0, n9928_0, n3603, n3595, n3507, n3499, n3491}), .out(n10054), .config_in(config_chain[15211:15206]), .config_rst(config_rst)); 
buffer_wire buffer_10054 (.in(n10054), .out(n10054_0));
mux15 mux_4889 (.in({n14201_2, n14179_1, n14174_0, n14151_0, n14146_0, n14123_0, n14116_0, n14093_0, n14088_0, n10135_0, n6541, n6529, n6441, n6433, n6425/**/}), .out(n10055), .config_in(config_chain[15217:15212]), .config_rst(config_rst)); 
buffer_wire buffer_10055 (.in(n10055), .out(n10055_0));
mux15 mux_4890 (.in({n13133_1, n13122_0, n13109_0, n13098_0/**/, n13086_0, n13083_0, n13072_0, n13057_0, n13044_0, n9936_0, n3603, n3595, n3507, n3499, n3491}), .out(n10056), .config_in(config_chain[15223:15218]), .config_rst(config_rst)); 
buffer_wire buffer_10056 (.in(n10056), .out(n10056_0));
mux15 mux_4891 (.in({n14199_1, n14176_0, n14155_0, n14148_0, n14125_0, n14118_0, n14096_0/**/, n14095_0, n14090_0, n10137_0, n6541, n6533, n6441, n6433, n6425}), .out(n10057), .config_in(config_chain[15229:15224]), .config_rst(config_rst)); 
buffer_wire buffer_10057 (.in(n10057), .out(n10057_0));
mux15 mux_4892 (.in({n13135_1, n13124_0, n13113_0, n13100_0, n13085_0, n13078_0, n13074_0, n13059_0/**/, n13048_0, n9944_0, n3603, n3595, n3507, n3499, n3491}), .out(n10058), .config_in(config_chain[15235:15230]), .config_rst(config_rst)); 
buffer_wire buffer_10058 (.in(n10058), .out(n10058_0));
mux15 mux_4893 (.in({n14197_1, n14178_0, n14157_0, n14150_0, n14127_0, n14122_0, n14104_0, n14099_0, n14092_0, n10139_0, n6541, n6533, n6525, n6433, n6425/**/}), .out(n10059), .config_in(config_chain[15241:15236]), .config_rst(config_rst)); 
buffer_wire buffer_10059 (.in(n10059), .out(n10059_0));
mux15 mux_4894 (.in({n13137_1, n13126_0, n13115_0, n13104_0/**/, n13089_0, n13076_0, n13070_0, n13061_0, n13050_0, n9952_0, n3603, n3595, n3507, n3499, n3491}), .out(n10060), .config_in(config_chain[15247:15242]), .config_rst(config_rst)); 
buffer_wire buffer_10060 (.in(n10060), .out(n10060_0));
mux14 mux_4895 (.in({n14195_1, n14159_0, n14154_0, n14131_0, n14124_0, n14112_0/**/, n14101_0, n14094_0, n10141_0, n6541, n6533, n6525, n6437, n6425}), .out(n10061), .config_in(config_chain[15253:15248]), .config_rst(config_rst)); 
buffer_wire buffer_10061 (.in(n10061), .out(n10061_0));
mux15 mux_4896 (.in({n13139_1, n13128_0, n13117_0, n13106_0, n13091_0, n13080_0, n13065_0, n13062_0, n13052_0, n9960_0, n3607, n3599/**/, n3591, n3503, n3495}), .out(n10062), .config_in(config_chain[15259:15254]), .config_rst(config_rst)); 
buffer_wire buffer_10062 (.in(n10062), .out(n10062_0));
mux14 mux_4897 (.in({n14193_1, n14163_0, n14156_0, n14133_0, n14126_0, n14120_0, n14103_0, n14098_0, n10143_0, n6541, n6533, n6525, n6437, n6429/**/}), .out(n10063), .config_in(config_chain[15265:15260]), .config_rst(config_rst)); 
buffer_wire buffer_10063 (.in(n10063), .out(n10063_0));
mux15 mux_4898 (.in({n13141_1, n13119_1, n13108_0, n13093_0, n13082_0, n13067_0, n13056_0, n13054_0, n13041_0, n9968_0/**/, n3607, n3599, n3591, n3503, n3495}), .out(n10064), .config_in(config_chain[15271:15266]), .config_rst(config_rst)); 
buffer_wire buffer_10064 (.in(n10064), .out(n10064_0));
mux13 mux_4899 (.in({n14191_1, n14165_0, n14158_0, n14135_0, n14130_0, n14128_0, n14107_0, n14100_0, n10145_0, n6533, n6525, n6437, n6429}), .out(n10065), .config_in(config_chain[15277:15272]), .config_rst(config_rst)); 
buffer_wire buffer_10065 (.in(n10065), .out(n10065_0));
mux15 mux_4900 (.in({n13143_1, n13121_1, n13112_0, n13097_0, n13084_0, n13069_0, n13058_0, n13046_0, n13043_0/**/, n9976_0, n3607, n3599, n3591, n3503, n3495}), .out(n10066), .config_in(config_chain[15283:15278]), .config_rst(config_rst)); 
buffer_wire buffer_10066 (.in(n10066), .out(n10066_0));
mux13 mux_4901 (.in({n14189_1, n14167_0, n14162_0, n14139_0, n14136_0, n14132_0, n14109_0, n14102_0, n10147_0, n6537, n6525, n6437, n6429}), .out(n10067), .config_in(config_chain[15289:15284]), .config_rst(config_rst)); 
buffer_wire buffer_10067 (.in(n10067), .out(n10067_0));
mux15 mux_4902 (.in({n13145_1, n13123_1, n13114_0, n13099_0, n13088_0, n13073_0, n13060_0, n13045_0, n13038_0, n9984_0, n3607, n3599/**/, n3591, n3503, n3495}), .out(n10068), .config_in(config_chain[15295:15290]), .config_rst(config_rst)); 
buffer_wire buffer_10068 (.in(n10068), .out(n10068_0));
mux13 mux_4903 (.in({n14187_1, n14171_0, n14164_0, n14144_0, n14141_0, n14134_0, n14111_0, n14106_0, n10149_0, n6537, n6529, n6437, n6429/**/}), .out(n10069), .config_in(config_chain[15301:15296]), .config_rst(config_rst)); 
buffer_wire buffer_10069 (.in(n10069), .out(n10069_0));
mux15 mux_4904 (.in({n13147_1, n13125_2, n13116_0, n13110_0, n13101_0, n13090_0, n13075_0, n13064_0, n13049_0, n9992_0/**/, n3607, n3599, n3591, n3503, n3495}), .out(n10070), .config_in(config_chain[15307:15302]), .config_rst(config_rst)); 
buffer_wire buffer_10070 (.in(n10070), .out(n10070_0));
mux13 mux_4905 (.in({n14185_1, n14173_0, n14166_0, n14152_0, n14143_0, n14138_0, n14115_0, n14108_0, n10151_0, n6537/**/, n6529, n6441, n6429}), .out(n10071), .config_in(config_chain[15313:15308]), .config_rst(config_rst)); 
buffer_wire buffer_10071 (.in(n10071), .out(n10071_0));
mux16 mux_4906 (.in({n13409_1, n13387_2, n13378_0, n13364_0/**/, n13363_0, n13352_0, n13337_0, n13326_0, n13311_0, n13298_0, n9922_1, n4581, n4573, n4485, n4477, n4469}), .out(n10072), .config_in(config_chain[15319:15314]), .config_rst(config_rst)); 
buffer_wire buffer_10072 (.in(n10072), .out(n10072_0));
mux15 mux_4907 (.in({n14445_1, n14441_0, n14436_0, n14434_0, n14413_0, n14406_0, n14383_0, n14376_0, n14353_0, n10155_0, n7515, n7507, n7419, n7411, n7403}), .out(n10073), .config_in(config_chain[15325:15320]), .config_rst(config_rst)); 
buffer_wire buffer_10073 (.in(n10073), .out(n10073_0));
mux16 mux_4908 (.in({n13391_1, n13389_2, n13380_0, n13367_0, n13356_0, n13354_0, n13339_0, n13328_0, n13313_0, n13302_0, n9930_1, n4581, n4573, n4485, n4477, n4469/**/}), .out(n10074), .config_in(config_chain[15331:15326]), .config_rst(config_rst)); 
buffer_wire buffer_10074 (.in(n10074), .out(n10074_0));
mux15 mux_4909 (.in({n14465_2, n14443_1, n14438_0, n14415_0, n14408_0/**/, n14385_0, n14380_0, n14357_0, n14354_0, n10157_0, n7519, n7507, n7419, n7411, n7403}), .out(n10075), .config_in(config_chain[15337:15332]), .config_rst(config_rst)); 
buffer_wire buffer_10075 (.in(n10075), .out(n10075_0));
mux15 mux_4910 (.in({n13393_1, n13382_0, n13369_0, n13358_0, n13348_0, n13343_0, n13330_0, n13315_0, n13304_0, n9938_1, n4581, n4573, n4485, n4477, n4469/**/}), .out(n10076), .config_in(config_chain[15343:15338]), .config_rst(config_rst)); 
buffer_wire buffer_10076 (.in(n10076), .out(n10076_0));
mux15 mux_4911 (.in({n14463_1, n14440_0, n14417_0, n14412_0, n14389_0, n14382_0, n14362_0, n14359_0, n14352_0, n10159_0, n7519, n7511, n7419, n7411, n7403}), .out(n10077), .config_in(config_chain[15349:15344]), .config_rst(config_rst)); 
buffer_wire buffer_10077 (.in(n10077), .out(n10077_0));
mux15 mux_4912 (.in({n13395_1, n13384_0, n13371_0, n13360_0, n13345_0, n13340_0, n13334_0, n13319_0, n13306_0, n9946_1, n4581, n4573, n4485, n4477, n4469/**/}), .out(n10078), .config_in(config_chain[15355:15350]), .config_rst(config_rst)); 
buffer_wire buffer_10078 (.in(n10078), .out(n10078_0));
mux15 mux_4913 (.in({n14461_1/**/, n14442_0, n14421_0, n14414_0, n14391_0, n14384_0, n14370_0, n14361_0, n14356_0, n10161_0, n7519, n7511, n7503, n7411, n7403}), .out(n10079), .config_in(config_chain[15361:15356]), .config_rst(config_rst)); 
buffer_wire buffer_10079 (.in(n10079), .out(n10079_0));
mux15 mux_4914 (.in({n13397_1, n13386_0, n13375_0, n13362_0, n13347_0, n13336_0, n13332_0, n13321_0, n13310_0, n9954_1/**/, n4581, n4573, n4485, n4477, n4469}), .out(n10080), .config_in(config_chain[15367:15362]), .config_rst(config_rst)); 
buffer_wire buffer_10080 (.in(n10080), .out(n10080_0));
mux14 mux_4915 (.in({n14459_1, n14423_0, n14416_0, n14393_0, n14388_0, n14378_0, n14365_0, n14358_0/**/, n10163_0, n7519, n7511, n7503, n7415, n7403}), .out(n10081), .config_in(config_chain[15373:15368]), .config_rst(config_rst)); 
buffer_wire buffer_10081 (.in(n10081), .out(n10081_0));
mux15 mux_4916 (.in({n13399_1, n13388_0, n13377_0, n13366_0, n13351_0, n13338_0, n13324_0, n13323_0, n13312_0/**/, n9962_1, n4585, n4577, n4569, n4481, n4473}), .out(n10082), .config_in(config_chain[15379:15374]), .config_rst(config_rst)); 
buffer_wire buffer_10082 (.in(n10082), .out(n10082_0));
mux14 mux_4917 (.in({n14457_1, n14425_0, n14420_0, n14397_0, n14390_0, n14386_0, n14367_0, n14360_0, n10165_0, n7519, n7511, n7503, n7415, n7407}), .out(n10083), .config_in(config_chain[15385:15380]), .config_rst(config_rst)); 
buffer_wire buffer_10083 (.in(n10083), .out(n10083_0));
mux15 mux_4918 (.in({n13401_1, n13379_0, n13368_0, n13353_0, n13342_0, n13327_0, n13316_0, n13314_0, n13299_0, n9970_1, n4585, n4577, n4569, n4481/**/, n4473}), .out(n10084), .config_in(config_chain[15391:15386]), .config_rst(config_rst)); 
buffer_wire buffer_10084 (.in(n10084), .out(n10084_0));
mux13 mux_4919 (.in({n14455_1, n14429_0/**/, n14422_0, n14399_0, n14394_0, n14392_0, n14369_0, n14364_0, n10167_0, n7511, n7503, n7415, n7407}), .out(n10085), .config_in(config_chain[15397:15392]), .config_rst(config_rst)); 
buffer_wire buffer_10085 (.in(n10085), .out(n10085_0));
mux15 mux_4920 (.in({n13403_1, n13381_1, n13370_0/**/, n13355_0, n13344_0, n13329_0, n13318_0, n13308_0, n13303_0, n9978_1, n4585, n4577, n4569, n4481, n4473}), .out(n10086), .config_in(config_chain[15403:15398]), .config_rst(config_rst)); 
buffer_wire buffer_10086 (.in(n10086), .out(n10086_0));
mux13 mux_4921 (.in({n14453_1/**/, n14431_0, n14424_0, n14402_0, n14401_0, n14396_0, n14373_0, n14366_0, n10169_0, n7515, n7503, n7415, n7407}), .out(n10087), .config_in(config_chain[15409:15404]), .config_rst(config_rst)); 
buffer_wire buffer_10087 (.in(n10087), .out(n10087_0));
mux15 mux_4922 (.in({n13405_1, n13383_1, n13374_0, n13359_0, n13346_0, n13331_0, n13320_0, n13305_0, n13300_0, n9986_1/**/, n4585, n4577, n4569, n4481, n4473}), .out(n10088), .config_in(config_chain[15415:15410]), .config_rst(config_rst)); 
buffer_wire buffer_10088 (.in(n10088), .out(n10088_0));
mux13 mux_4923 (.in({n14451_1, n14433_2, n14428_0, n14410_0, n14405_0, n14398_0, n14375_0, n14368_0, n10171_0, n7515, n7507, n7415, n7407}), .out(n10089), .config_in(config_chain[15421:15416]), .config_rst(config_rst)); 
buffer_wire buffer_10089 (.in(n10089), .out(n10089_0));
mux15 mux_4924 (.in({n13407_1, n13385_1, n13376_0, n13372_0, n13361_0, n13350_0, n13335_0, n13322_0, n13307_0, n9994_1/**/, n4585, n4577, n4569, n4481, n4473}), .out(n10090), .config_in(config_chain[15427:15422]), .config_rst(config_rst)); 
buffer_wire buffer_10090 (.in(n10090), .out(n10090_0));
mux13 mux_4925 (.in({n14449_1, n14437_0, n14430_0, n14418_0, n14407_0, n14400_0, n14377_0, n14372_0, n10173_0, n7515, n7507, n7419, n7407}), .out(n10091), .config_in(config_chain[15433:15428]), .config_rst(config_rst)); 
buffer_wire buffer_10091 (.in(n10091), .out(n10091_0));
mux16 mux_4926 (.in({n13671_1, n13649_1, n13640_0, n13628_0, n13625_0, n13614_0, n13599_0/**/, n13586_0, n13571_0, n13560_0, n10012_1, n5559, n5551, n5463, n5455, n5447}), .out(n10092), .config_in(config_chain[15439:15434]), .config_rst(config_rst)); 
buffer_wire buffer_10092 (.in(n10092), .out(n10092_0));
mux4 mux_4927 (.in({n14707_1/**/, n14618_0, n8497, n8381}), .out(n10093), .config_in(config_chain[15441:15440]), .config_rst(config_rst)); 
buffer_wire buffer_10093 (.in(n10093), .out(n10093_0));
mux16 mux_4928 (.in({n13653_1, n13651_2, n13642_0, n13627_0, n13620_0, n13616_0, n13601_0, n13590_0, n13575_0, n13562_0, n10014_1, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10094), .config_in(config_chain[15447:15442]), .config_rst(config_rst)); 
buffer_wire buffer_10094 (.in(n10094), .out(n10094_0));
mux3 mux_4929 (.in({n14709_1/**/, n14626_0, n8385}), .out(n10095), .config_in(config_chain[15449:15448]), .config_rst(config_rst)); 
buffer_wire buffer_10095 (.in(n10095), .out(n10095_0));
mux15 mux_4930 (.in({n13655_1, n13644_0, n13631_0, n13618_0, n13612_0, n13603_0, n13592_0, n13577_0, n13566_0, n10016_1, n5559, n5551, n5463/**/, n5455, n5447}), .out(n10096), .config_in(config_chain[15455:15450]), .config_rst(config_rst)); 
buffer_wire buffer_10096 (.in(n10096), .out(n10096_0));
mux3 mux_4931 (.in({n14711_1/**/, n14634_0, n8389}), .out(n10097), .config_in(config_chain[15457:15456]), .config_rst(config_rst)); 
buffer_wire buffer_10097 (.in(n10097), .out(n10097_0));
mux15 mux_4932 (.in({n13657_1, n13646_0, n13633_0, n13622_0, n13607_0, n13604_0, n13594_0, n13579_0, n13568_0, n10018_1, n5559, n5551, n5463, n5455/**/, n5447}), .out(n10098), .config_in(config_chain[15463:15458]), .config_rst(config_rst)); 
buffer_wire buffer_10098 (.in(n10098), .out(n10098_0));
mux3 mux_4933 (.in({n14713_1, n14642_0/**/, n8389}), .out(n10099), .config_in(config_chain[15465:15464]), .config_rst(config_rst)); 
buffer_wire buffer_10099 (.in(n10099), .out(n10099_0));
mux15 mux_4934 (.in({n13659_1, n13648_0, n13635_0, n13624_0, n13609_0, n13598_0, n13596_0/**/, n13583_0, n13570_0, n10020_1, n5559, n5551, n5463, n5455, n5447}), .out(n10100), .config_in(config_chain[15471:15466]), .config_rst(config_rst)); 
buffer_wire buffer_10100 (.in(n10100), .out(n10100_0));
mux3 mux_4935 (.in({n14715_1/**/, n14650_0, n8393}), .out(n10101), .config_in(config_chain[15473:15472]), .config_rst(config_rst)); 
buffer_wire buffer_10101 (.in(n10101), .out(n10101_0));
mux15 mux_4936 (.in({n13661_1, n13650_0, n13639_0, n13626_0, n13611_0, n13600_0, n13588_0, n13585_0, n13574_0/**/, n10022_1, n5563, n5555, n5547, n5459, n5451}), .out(n10102), .config_in(config_chain[15479:15474]), .config_rst(config_rst)); 
buffer_wire buffer_10102 (.in(n10102), .out(n10102_0));
mux3 mux_4937 (.in({n14717_1, n14658_0/**/, n8397}), .out(n10103), .config_in(config_chain[15481:15480]), .config_rst(config_rst)); 
buffer_wire buffer_10103 (.in(n10103), .out(n10103_0));
mux15 mux_4938 (.in({n13663_1, n13641_0/**/, n13630_0, n13615_0, n13602_0, n13587_0, n13580_0, n13576_0, n13561_0, n10024_1, n5563, n5555, n5547, n5459, n5451}), .out(n10104), .config_in(config_chain[15487:15482]), .config_rst(config_rst)); 
buffer_wire buffer_10104 (.in(n10104), .out(n10104_0));
mux3 mux_4939 (.in({n14719_1, n14666_0/**/, n8481}), .out(n10105), .config_in(config_chain[15489:15488]), .config_rst(config_rst)); 
buffer_wire buffer_10105 (.in(n10105), .out(n10105_0));
mux15 mux_4940 (.in({n13665_1, n13643_0, n13632_0, n13617_0, n13606_0, n13591_0, n13578_0, n13572_0, n13563_0, n10026_1/**/, n5563, n5555, n5547, n5459, n5451}), .out(n10106), .config_in(config_chain[15495:15490]), .config_rst(config_rst)); 
buffer_wire buffer_10106 (.in(n10106), .out(n10106_0));
mux3 mux_4941 (.in({n14721_1/**/, n14674_0, n8485}), .out(n10107), .config_in(config_chain[15497:15496]), .config_rst(config_rst)); 
buffer_wire buffer_10107 (.in(n10107), .out(n10107_0));
mux15 mux_4942 (.in({n13667_1, n13645_1, n13634_0, n13619_0, n13608_0, n13593_0, n13582_0, n13567_0, n13564_0/**/, n10028_1, n5563, n5555, n5547, n5459, n5451}), .out(n10108), .config_in(config_chain[15503:15498]), .config_rst(config_rst)); 
buffer_wire buffer_10108 (.in(n10108), .out(n10108_0));
mux3 mux_4943 (.in({n14723_1, n14682_0, n8485}), .out(n10109), .config_in(config_chain[15505:15504]), .config_rst(config_rst)); 
buffer_wire buffer_10109 (.in(n10109), .out(n10109_0));
mux15 mux_4944 (.in({n13669_1, n13647_1, n13638_0, n13636_0, n13623_0, n13610_0, n13595_0, n13584_0/**/, n13569_0, n10030_1, n5563, n5555, n5547, n5459, n5451}), .out(n10110), .config_in(config_chain[15511:15506]), .config_rst(config_rst)); 
buffer_wire buffer_10110 (.in(n10110), .out(n10110_0));
mux3 mux_4945 (.in({n14725_1, n14690_0, n8489}), .out(n10111), .config_in(config_chain[15513:15512]), .config_rst(config_rst)); 
buffer_wire buffer_10111 (.in(n10111), .out(n10111_0));
mux16 mux_4946 (.in({n13935_1, n13913_1, n13904_0, n13894_0, n13889_0, n13876_0, n13861_0, n13850_0, n13835_0, n13824_0, n10032_1/**/, n6537, n6529, n6441, n6433, n6425}), .out(n10112), .config_in(config_chain[15519:15514]), .config_rst(config_rst)); 
buffer_wire buffer_10112 (.in(n10112), .out(n10112_0));
mux4 mux_4947 (.in({n14621_0, n14620_0, n8497, n8381}), .out(n10113), .config_in(config_chain[15521:15520]), .config_rst(config_rst)); 
buffer_wire buffer_10113 (.in(n10113), .out(n10113_0));
mux16 mux_4948 (.in({n13917_1, n13915_1, n13906_0, n13891_0, n13886_0, n13880_0/**/, n13865_0, n13852_0, n13837_0, n13826_0, n10034_1, n6537, n6529, n6441, n6433, n6425}), .out(n10114), .config_in(config_chain[15527:15522]), .config_rst(config_rst)); 
buffer_wire buffer_10114 (.in(n10114), .out(n10114_0));
mux3 mux_4949 (.in({n14629_0, n14628_0, n8385}), .out(n10115), .config_in(config_chain[15529:15528]), .config_rst(config_rst)); 
buffer_wire buffer_10115 (.in(n10115), .out(n10115_0));
mux15 mux_4950 (.in({n13919_1, n13908_0, n13893_0, n13882_0, n13878_0, n13867_0, n13856_0/**/, n13841_0, n13828_0, n10036_1, n6537, n6529, n6441, n6433, n6425}), .out(n10116), .config_in(config_chain[15535:15530]), .config_rst(config_rst)); 
buffer_wire buffer_10116 (.in(n10116), .out(n10116_0));
mux3 mux_4951 (.in({n14637_0, n14636_0, n8389}), .out(n10117), .config_in(config_chain[15537:15536]), .config_rst(config_rst)); 
buffer_wire buffer_10117 (.in(n10117), .out(n10117_0));
mux15 mux_4952 (.in({n13921_1, n13910_0, n13897_0, n13884_0, n13870_0, n13869_0, n13858_0, n13843_0, n13832_0, n10038_1, n6537, n6529, n6441/**/, n6433, n6425}), .out(n10118), .config_in(config_chain[15543:15538]), .config_rst(config_rst)); 
buffer_wire buffer_10118 (.in(n10118), .out(n10118_0));
mux3 mux_4953 (.in({n14645_0, n14644_0, n8393}), .out(n10119), .config_in(config_chain[15545:15544]), .config_rst(config_rst)); 
buffer_wire buffer_10119 (.in(n10119), .out(n10119_0));
mux15 mux_4954 (.in({n13923_1, n13912_0, n13899_0, n13888_0, n13873_0, n13862_0, n13860_0, n13845_0, n13834_0, n10040_1, n6537, n6529, n6441, n6433, n6425/**/}), .out(n10120), .config_in(config_chain[15551:15546]), .config_rst(config_rst)); 
buffer_wire buffer_10120 (.in(n10120), .out(n10120_0));
mux3 mux_4955 (.in({n14653_0, n14652_0, n8393}), .out(n10121), .config_in(config_chain[15553:15552]), .config_rst(config_rst)); 
buffer_wire buffer_10121 (.in(n10121), .out(n10121_0));
mux15 mux_4956 (.in({n13925_1/**/, n13914_0, n13901_0, n13890_0, n13875_0, n13864_0, n13854_0, n13849_0, n13836_0, n10042_1, n6541, n6533, n6525, n6437, n6429}), .out(n10122), .config_in(config_chain[15559:15554]), .config_rst(config_rst)); 
buffer_wire buffer_10122 (.in(n10122), .out(n10122_0));
mux3 mux_4957 (.in({n14661_0, n14660_0, n8397}), .out(n10123), .config_in(config_chain[15561:15560]), .config_rst(config_rst)); 
buffer_wire buffer_10123 (.in(n10123), .out(n10123_0));
mux15 mux_4958 (.in({n13927_1, n13905_0, n13892_0, n13877_0, n13866_0, n13851_0, n13846_0, n13840_0, n13825_0, n10044_1, n6541, n6533/**/, n6525, n6437, n6429}), .out(n10124), .config_in(config_chain[15567:15562]), .config_rst(config_rst)); 
buffer_wire buffer_10124 (.in(n10124), .out(n10124_0));
mux3 mux_4959 (.in({n14669_0, n14668_0/**/, n8481}), .out(n10125), .config_in(config_chain[15569:15568]), .config_rst(config_rst)); 
buffer_wire buffer_10125 (.in(n10125), .out(n10125_0));
mux15 mux_4960 (.in({n13929_1, n13907_0, n13896_0, n13881_0, n13868_0, n13853_0, n13842_0/**/, n13838_0, n13827_0, n10046_1, n6541, n6533, n6525, n6437, n6429}), .out(n10126), .config_in(config_chain[15575:15570]), .config_rst(config_rst)); 
buffer_wire buffer_10126 (.in(n10126), .out(n10126_0));
mux3 mux_4961 (.in({n14677_0/**/, n14676_0, n8485}), .out(n10127), .config_in(config_chain[15577:15576]), .config_rst(config_rst)); 
buffer_wire buffer_10127 (.in(n10127), .out(n10127_0));
mux15 mux_4962 (.in({n13931_1, n13909_0, n13898_0, n13883_0, n13872_0, n13857_0, n13844_0, n13830_0, n13829_0, n10048_1, n6541, n6533, n6525, n6437, n6429/**/}), .out(n10128), .config_in(config_chain[15583:15578]), .config_rst(config_rst)); 
buffer_wire buffer_10128 (.in(n10128), .out(n10128_0));
mux3 mux_4963 (.in({n14685_0, n14684_0, n8489}), .out(n10129), .config_in(config_chain[15585:15584]), .config_rst(config_rst)); 
buffer_wire buffer_10129 (.in(n10129), .out(n10129_0));
mux15 mux_4964 (.in({n13933_1, n13911_1, n13902_0, n13900_0, n13885_0, n13874_0, n13859_0, n13848_0/**/, n13833_0, n10050_1, n6541, n6533, n6525, n6437, n6429}), .out(n10130), .config_in(config_chain[15591:15586]), .config_rst(config_rst)); 
buffer_wire buffer_10130 (.in(n10130), .out(n10130_0));
mux3 mux_4965 (.in({n14693_0, n14692_0, n8489}), .out(n10131), .config_in(config_chain[15593:15592]), .config_rst(config_rst)); 
buffer_wire buffer_10131 (.in(n10131), .out(n10131_0));
mux15 mux_4966 (.in({n14201_2, n14176_0, n14173_0, n14160_0, n14148_0, n14143_0, n14118_0, n14115_0, n14090_0, n10052_1/**/, n7515, n7507, n7419, n7411, n7403}), .out(n10132), .config_in(config_chain[15599:15594]), .config_rst(config_rst)); 
buffer_wire buffer_10132 (.in(n10132), .out(n10132_0));
mux4 mux_4967 (.in({n14615_0, n14614_0, n8497, n8381}), .out(n10133), .config_in(config_chain[15601:15600]), .config_rst(config_rst)); 
buffer_wire buffer_10133 (.in(n10133), .out(n10133_0));
mux15 mux_4968 (.in({n14181_1, n14178_0, n14175_0, n14152_0, n14150_0, n14147_0/**/, n14122_0, n14117_0, n14092_0, n10054_1, n7519, n7507, n7419, n7411, n7403}), .out(n10134), .config_in(config_chain[15607:15602]), .config_rst(config_rst)); 
buffer_wire buffer_10134 (.in(n10134), .out(n10134_0));
mux3 mux_4969 (.in({n14623_0, n14622_0, n8381}), .out(n10135), .config_in(config_chain[15609:15608]), .config_rst(config_rst)); 
buffer_wire buffer_10135 (.in(n10135), .out(n10135_0));
mux15 mux_4970 (.in({n14183_1, n14177_1, n14154_0, n14149_0, n14144_0/**/, n14124_0, n14119_0, n14094_0, n14091_0, n10056_1, n7519, n7511, n7419, n7411, n7403}), .out(n10136), .config_in(config_chain[15615:15610]), .config_rst(config_rst)); 
buffer_wire buffer_10136 (.in(n10136), .out(n10136_0));
mux3 mux_4971 (.in({n14631_0, n14630_0, n8385}), .out(n10137), .config_in(config_chain[15617:15616]), .config_rst(config_rst)); 
buffer_wire buffer_10137 (.in(n10137), .out(n10137_0));
mux15 mux_4972 (.in({n14185_1, n14179_1, n14156_0, n14151_0, n14136_0/**/, n14126_0, n14123_0, n14098_0, n14093_0, n10058_1, n7519, n7511, n7503, n7411, n7403}), .out(n10138), .config_in(config_chain[15623:15618]), .config_rst(config_rst)); 
buffer_wire buffer_10138 (.in(n10138), .out(n10138_0));
mux3 mux_4973 (.in({n14639_0/**/, n14638_0, n8389}), .out(n10139), .config_in(config_chain[15625:15624]), .config_rst(config_rst)); 
buffer_wire buffer_10139 (.in(n10139), .out(n10139_0));
mux14 mux_4974 (.in({n14187_1, n14158_0, n14155_0, n14130_0, n14128_0/**/, n14125_0, n14100_0, n14095_0, n10060_1, n7519, n7511, n7503, n7415, n7403}), .out(n10140), .config_in(config_chain[15631:15626]), .config_rst(config_rst)); 
buffer_wire buffer_10140 (.in(n10140), .out(n10140_0));
mux3 mux_4975 (.in({n14647_0, n14646_0, n8393}), .out(n10141), .config_in(config_chain[15633:15632]), .config_rst(config_rst)); 
buffer_wire buffer_10141 (.in(n10141), .out(n10141_0));
mux14 mux_4976 (.in({n14189_1, n14162_0, n14157_0, n14132_0, n14127_0, n14120_0, n14102_0, n14099_0/**/, n10062_1, n7519, n7511, n7503, n7415, n7407}), .out(n10142), .config_in(config_chain[15639:15634]), .config_rst(config_rst)); 
buffer_wire buffer_10142 (.in(n10142), .out(n10142_0));
mux3 mux_4977 (.in({n14655_0, n14654_0, n8397}), .out(n10143), .config_in(config_chain[15641:15640]), .config_rst(config_rst)); 
buffer_wire buffer_10143 (.in(n10143), .out(n10143_0));
mux13 mux_4978 (.in({n14191_1, n14164_0, n14159_0, n14134_0, n14131_0, n14112_0/**/, n14106_0, n14101_0, n10064_1, n7511, n7503, n7415, n7407}), .out(n10144), .config_in(config_chain[15647:15642]), .config_rst(config_rst)); 
buffer_wire buffer_10144 (.in(n10144), .out(n10144_0));
mux3 mux_4979 (.in({n14663_0, n14662_0, n8397}), .out(n10145), .config_in(config_chain[15649:15648]), .config_rst(config_rst)); 
buffer_wire buffer_10145 (.in(n10145), .out(n10145_0));
mux13 mux_4980 (.in({n14193_1, n14166_0, n14163_0, n14138_0, n14133_0, n14108_0, n14104_0, n14103_0, n10066_1, n7515, n7503, n7415, n7407}), .out(n10146), .config_in(config_chain[15655:15650]), .config_rst(config_rst)); 
buffer_wire buffer_10146 (.in(n10146), .out(n10146_0));
mux3 mux_4981 (.in({n14671_0/**/, n14670_0, n8481}), .out(n10147), .config_in(config_chain[15657:15656]), .config_rst(config_rst)); 
buffer_wire buffer_10147 (.in(n10147), .out(n10147_0));
mux13 mux_4982 (.in({n14195_1, n14170_0, n14165_0, n14140_0, n14135_0, n14110_0, n14107_0, n14096_0, n10068_1, n7515/**/, n7507, n7415, n7407}), .out(n10148), .config_in(config_chain[15663:15658]), .config_rst(config_rst)); 
buffer_wire buffer_10148 (.in(n10148), .out(n10148_0));
mux3 mux_4983 (.in({n14679_0, n14678_0, n8485}), .out(n10149), .config_in(config_chain[15665:15664]), .config_rst(config_rst)); 
buffer_wire buffer_10149 (.in(n10149), .out(n10149_0));
mux13 mux_4984 (.in({n14197_1, n14172_0, n14167_0, n14142_0, n14139_0, n14114_0, n14109_0, n14088_0, n10070_1, n7515, n7507/**/, n7419, n7407}), .out(n10150), .config_in(config_chain[15671:15666]), .config_rst(config_rst)); 
buffer_wire buffer_10150 (.in(n10150), .out(n10150_0));
mux3 mux_4985 (.in({n14687_0, n14686_0, n8489}), .out(n10151), .config_in(config_chain[15673:15672]), .config_rst(config_rst)); 
buffer_wire buffer_10151 (.in(n10151), .out(n10151_0));
mux13 mux_4986 (.in({n14199_1, n14174_0, n14171_0, n14168_0, n14146_0, n14141_0, n14116_0, n14111_0, n10000_2, n7515, n7507, n7419, n7411}), .out(n10152), .config_in(config_chain[15679:15674]), .config_rst(config_rst)); 
buffer_wire buffer_10152 (.in(n10152), .out(n10152_0));
mux3 mux_4987 (.in({n14695_2, n14694_0, n8493}), .out(n10153), .config_in(config_chain[15681:15680]), .config_rst(config_rst)); 
buffer_wire buffer_10153 (.in(n10153), .out(n10153_0));
mux15 mux_4988 (.in({n14465_2, n14440_0, n14437_0, n14426_0, n14412_0, n14407_0, n14382_0, n14377_0, n14352_0, n10072_1, n8493, n8485, n8397, n8389, n8381}), .out(n10154), .config_in(config_chain[15687:15682]), .config_rst(config_rst)); 
buffer_wire buffer_10154 (.in(n10154), .out(n10154_0));
mux4 mux_4989 (.in({n14617_0, n14616_0, n8497, n8381}), .out(n10155), .config_in(config_chain[15689:15688]), .config_rst(config_rst)); 
buffer_wire buffer_10155 (.in(n10155), .out(n10155_0));
mux15 mux_4990 (.in({n14445_1, n14442_0, n14439_0, n14418_0, n14414_0, n14409_0, n14384_0, n14381_0, n14356_0, n10074_1, n8497, n8485, n8397, n8389, n8381}), .out(n10156), .config_in(config_chain[15695:15690]), .config_rst(config_rst)); 
buffer_wire buffer_10156 (.in(n10156), .out(n10156_0));
mux3 mux_4991 (.in({n14625_0, n14624_0, n8385}), .out(n10157), .config_in(config_chain[15697:15696]), .config_rst(config_rst)); 
buffer_wire buffer_10157 (.in(n10157), .out(n10157_0));
mux15 mux_4992 (.in({n14447_1, n14441_0, n14416_0, n14413_0, n14410_0, n14388_0, n14383_0, n14358_0, n14353_0, n10076_1, n8497, n8489, n8397, n8389, n8381}), .out(n10158), .config_in(config_chain[15703:15698]), .config_rst(config_rst)); 
buffer_wire buffer_10158 (.in(n10158), .out(n10158_0));
mux3 mux_4993 (.in({n14633_0, n14632_0, n8385}), .out(n10159), .config_in(config_chain[15705:15704]), .config_rst(config_rst)); 
buffer_wire buffer_10159 (.in(n10159), .out(n10159_0));
mux15 mux_4994 (.in({n14449_1, n14443_1, n14420_0, n14415_0, n14402_0, n14390_0, n14385_0, n14360_0, n14357_0, n10078_1, n8497, n8489, n8481, n8389, n8381}), .out(n10160), .config_in(config_chain[15711:15706]), .config_rst(config_rst)); 
buffer_wire buffer_10160 (.in(n10160), .out(n10160_0));
mux3 mux_4995 (.in({n14641_0, n14640_0, n8389}), .out(n10161), .config_in(config_chain[15713:15712]), .config_rst(config_rst)); 
buffer_wire buffer_10161 (.in(n10161), .out(n10161_0));
mux14 mux_4996 (.in({n14451_1, n14422_0, n14417_0, n14394_0, n14392_0, n14389_0, n14364_0, n14359_0, n10080_1, n8497, n8489, n8481, n8393, n8381}), .out(n10162), .config_in(config_chain[15719:15714]), .config_rst(config_rst)); 
buffer_wire buffer_10162 (.in(n10162), .out(n10162_0));
mux3 mux_4997 (.in({n14649_0, n14648_0, n8393}), .out(n10163), .config_in(config_chain[15721:15720]), .config_rst(config_rst)); 
buffer_wire buffer_10163 (.in(n10163), .out(n10163_0));
mux14 mux_4998 (.in({n14453_1, n14424_0/**/, n14421_0, n14396_0, n14391_0, n14386_0, n14366_0, n14361_0, n10082_1, n8497, n8489, n8481, n8393, n8385}), .out(n10164), .config_in(config_chain[15727:15722]), .config_rst(config_rst)); 
buffer_wire buffer_10164 (.in(n10164), .out(n10164_0));
mux3 mux_4999 (.in({n14657_0, n14656_0, n8397}), .out(n10165), .config_in(config_chain[15729:15728]), .config_rst(config_rst)); 
buffer_wire buffer_10165 (.in(n10165), .out(n10165_0));
mux13 mux_5000 (.in({n14455_1, n14428_0, n14423_0, n14398_0, n14393_0, n14378_0, n14368_0, n14365_0, n10084_1, n8489, n8481, n8393, n8385}), .out(n10166), .config_in(config_chain[15735:15730]), .config_rst(config_rst)); 
buffer_wire buffer_10166 (.in(n10166), .out(n10166_0));
mux3 mux_5001 (.in({n14665_0, n14664_0, n8481}), .out(n10167), .config_in(config_chain[15737:15736]), .config_rst(config_rst)); 
buffer_wire buffer_10167 (.in(n10167), .out(n10167_0));
mux13 mux_5002 (.in({n14457_1, n14430_0, n14425_0, n14400_0/**/, n14397_0, n14372_0, n14370_0, n14367_0, n10086_1, n8493, n8481, n8393, n8385}), .out(n10168), .config_in(config_chain[15743:15738]), .config_rst(config_rst)); 
buffer_wire buffer_10168 (.in(n10168), .out(n10168_0));
mux3 mux_5003 (.in({n14673_0, n14672_0, n8481}), .out(n10169), .config_in(config_chain[15745:15744]), .config_rst(config_rst)); 
buffer_wire buffer_10169 (.in(n10169), .out(n10169_0));
mux13 mux_5004 (.in({n14459_1, n14432_0, n14429_0, n14404_0, n14399_0, n14374_0, n14369_0, n14362_0, n10088_1, n8493, n8485, n8393, n8385}), .out(n10170), .config_in(config_chain[15751:15746]), .config_rst(config_rst)); 
buffer_wire buffer_10170 (.in(n10170), .out(n10170_0));
mux3 mux_5005 (.in({n14681_0, n14680_0, n8485}), .out(n10171), .config_in(config_chain[15753:15752]), .config_rst(config_rst)); 
buffer_wire buffer_10171 (.in(n10171), .out(n10171_0));
mux13 mux_5006 (.in({n14461_1, n14436_0, n14431_0, n14406_0, n14401_0, n14376_0, n14373_0, n14354_0, n10090_1, n8493, n8485, n8397, n8385}), .out(n10172), .config_in(config_chain[15759:15754]), .config_rst(config_rst)); 
buffer_wire buffer_10172 (.in(n10172), .out(n10172_0));
mux3 mux_5007 (.in({n14689_0, n14688_0, n8489}), .out(n10173), .config_in(config_chain[15761:15760]), .config_rst(config_rst)); 
buffer_wire buffer_10173 (.in(n10173), .out(n10173_0));
mux13 mux_5008 (.in({n14463_1, n14438_0, n14434_0, n14433_2, n14408_0, n14405_0, n14380_0, n14375_0, n10002_2, n8493, n8485, n8397, n8389}), .out(n10174), .config_in(config_chain[15767:15762]), .config_rst(config_rst)); 
buffer_wire buffer_10174 (.in(n10174), .out(n10174_0));
mux3 mux_5009 (.in({n14697_2, n14696_0, n8493}), .out(n10175), .config_in(config_chain[15769:15768]), .config_rst(config_rst)); 
buffer_wire buffer_10175 (.in(n10175), .out(n10175_0));
mux4 mux_5010 (.in({n12271_0, n12270_0, n771, n655}), .out(n10176), .config_in(config_chain[15771:15770]), .config_rst(config_rst)); 
buffer_wire buffer_10176 (.in(n10176), .out(n10176_0));
mux16 mux_5011 (.in({n12893_1, n12885_0, n12880_0, n12868_0, n12861_1, n12852_0, n12846_0, n12809_0, n12792_0, n12783_0/**/, n10289_1, n1745, n1737, n1649, n1641, n1633}), .out(n10177), .config_in(config_chain[15777:15772]), .config_rst(config_rst)); 
buffer_wire buffer_10177 (.in(n10177), .out(n10177_0));
mux4 mux_5012 (.in({n12363_0, n12362_0, n771, n655}), .out(n10178), .config_in(config_chain[15779:15778]), .config_rst(config_rst)); 
buffer_wire buffer_10178 (.in(n10178), .out(n10178_0));
mux16 mux_5013 (.in({n13151_1, n13146_0, n13131_0, n13126_0, n13119_0, n13112_0/**/, n13093_0, n13076_0, n13067_0, n13050_0, n10309_1, n2723, n2715, n2627, n2619, n2611}), .out(n10179), .config_in(config_chain[15785:15780]), .config_rst(config_rst)); 
buffer_wire buffer_10179 (.in(n10179), .out(n10179_0));
mux4 mux_5014 (.in({n12383_1, n12274_0, n771, n655}), .out(n10180), .config_in(config_chain[15787:15786]), .config_rst(config_rst)); 
buffer_wire buffer_10180 (.in(n10180), .out(n10180_0));
mux16 mux_5015 (.in({n13411_1, n13397_0, n13392_0, n13386_0, n13379_0, n13374_0, n13362_0, n13353_0, n13336_0, n13299_0, n10329_1, n3701, n3693, n3605, n3597, n3589}), .out(n10181), .config_in(config_chain[15793:15788]), .config_rst(config_rst)); 
buffer_wire buffer_10181 (.in(n10181), .out(n10181_0));
mux4 mux_5016 (.in({n12277_0, n12276_0, n771, n655}), .out(n10182), .config_in(config_chain[15795:15794]), .config_rst(config_rst)); 
buffer_wire buffer_10182 (.in(n10182), .out(n10182_0));
mux16 mux_5017 (.in({n12637_1, n12629_0, n12624_0, n12612_0, n12605_1, n12602_0, n12588_0, n12551_0, n12534_0, n12525_0, n10269_1/**/, n767, n759, n671, n663, n655}), .out(n10183), .config_in(config_chain[15801:15796]), .config_rst(config_rst)); 
buffer_wire buffer_10183 (.in(n10183), .out(n10183_0));
mux3 mux_5018 (.in({n12279_0, n12278_0, n655}), .out(n10184), .config_in(config_chain[15803:15802]), .config_rst(config_rst)); 
buffer_wire buffer_10184 (.in(n10184), .out(n10184_0));
mux16 mux_5019 (.in({n12911_1, n12879_0, n12874_0, n12870_0, n12863_1, n12848_0, n12839_0, n12822_0, n12785_0, n12780_0/**/, n10291_1, n1745, n1737, n1649, n1641, n1633}), .out(n10185), .config_in(config_chain[15809:15804]), .config_rst(config_rst)); 
buffer_wire buffer_10185 (.in(n10185), .out(n10185_0));
mux3 mux_5020 (.in({n12365_0, n12364_0, n659}), .out(n10186), .config_in(config_chain[15811:15810]), .config_rst(config_rst)); 
buffer_wire buffer_10186 (.in(n10186), .out(n10186_0));
mux16 mux_5021 (.in({n13169_1, n13145_0, n13140_0, n13128_0, n13121_1, n13106_0, n13069_0, n13052_0, n13043_0, n13040_0, n10311_1, n2723, n2715, n2627, n2619/**/, n2611}), .out(n10187), .config_in(config_chain[15817:15812]), .config_rst(config_rst)); 
buffer_wire buffer_10187 (.in(n10187), .out(n10187_0));
mux3 mux_5022 (.in({n12385_1, n12282_0/**/, n659}), .out(n10188), .config_in(config_chain[15819:15818]), .config_rst(config_rst)); 
buffer_wire buffer_10188 (.in(n10188), .out(n10188_0));
mux16 mux_5023 (.in({n13429_1, n13406_0, n13391_0/**/, n13388_0, n13381_0, n13355_0, n13338_0, n13329_0, n13312_0, n13302_0, n10331_1, n3701, n3693, n3605, n3597, n3589}), .out(n10189), .config_in(config_chain[15825:15820]), .config_rst(config_rst)); 
buffer_wire buffer_10189 (.in(n10189), .out(n10189_0));
mux3 mux_5024 (.in({n12285_0, n12284_0, n659}), .out(n10190), .config_in(config_chain[15827:15826]), .config_rst(config_rst)); 
buffer_wire buffer_10190 (.in(n10190), .out(n10190_0));
mux16 mux_5025 (.in({n12655_1, n12623_0, n12618_0, n12614_0, n12607_1, n12590_0/**/, n12581_0, n12564_0, n12530_0, n12527_0, n10271_1, n767, n759, n671, n663, n655}), .out(n10191), .config_in(config_chain[15833:15828]), .config_rst(config_rst)); 
buffer_wire buffer_10191 (.in(n10191), .out(n10191_0));
mux3 mux_5026 (.in({n12287_0, n12286_0, n659}), .out(n10192), .config_in(config_chain[15835:15834]), .config_rst(config_rst)); 
buffer_wire buffer_10192 (.in(n10192), .out(n10192_0));
mux15 mux_5027 (.in({n12909_1, n12888_0, n12873_0, n12865_1, n12841_0, n12824_0, n12815_0, n12798_0, n12788_0, n10293_1, n1745, n1737, n1649, n1641, n1633}), .out(n10193), .config_in(config_chain[15841:15836]), .config_rst(config_rst)); 
buffer_wire buffer_10193 (.in(n10193), .out(n10193_0));
mux3 mux_5028 (.in({n12367_0, n12366_0, n659}), .out(n10194), .config_in(config_chain[15843:15842]), .config_rst(config_rst)); 
buffer_wire buffer_10194 (.in(n10194), .out(n10194_0));
mux15 mux_5029 (.in({n13167_1/**/, n13139_0, n13134_0, n13123_1, n13108_0, n13099_0, n13082_0, n13048_0, n13045_0, n10313_1, n2723, n2715, n2627, n2619, n2611}), .out(n10195), .config_in(config_chain[15849:15844]), .config_rst(config_rst)); 
buffer_wire buffer_10195 (.in(n10195), .out(n10195_0));
mux3 mux_5030 (.in({n12387_1, n12290_0, n663}), .out(n10196), .config_in(config_chain[15851:15850]), .config_rst(config_rst)); 
buffer_wire buffer_10196 (.in(n10196), .out(n10196_0));
mux15 mux_5031 (.in({n13427_1, n13405_0, n13400_0, n13383_1, n13368_0, n13331_0, n13314_0, n13310_0, n13305_0, n10333_1/**/, n3701, n3693, n3605, n3597, n3589}), .out(n10197), .config_in(config_chain[15857:15852]), .config_rst(config_rst)); 
buffer_wire buffer_10197 (.in(n10197), .out(n10197_0));
mux3 mux_5032 (.in({n12293_0/**/, n12292_0, n663}), .out(n10198), .config_in(config_chain[15859:15858]), .config_rst(config_rst)); 
buffer_wire buffer_10198 (.in(n10198), .out(n10198_0));
mux15 mux_5033 (.in({n12653_1, n12632_0, n12617_0, n12609_2, n12583_0, n12566_0, n12557_0, n12540_0, n12538_0, n10273_1, n767, n759, n671, n663, n655}), .out(n10199), .config_in(config_chain[15865:15860]), .config_rst(config_rst)); 
buffer_wire buffer_10199 (.in(n10199), .out(n10199_0));
mux3 mux_5034 (.in({n12295_0, n12294_0, n663}), .out(n10200), .config_in(config_chain[15867:15866]), .config_rst(config_rst)); 
buffer_wire buffer_10200 (.in(n10200), .out(n10200_0));
mux15 mux_5035 (.in({n12907_1, n12887_0, n12882_0, n12867_2, n12854_0, n12817_0/**/, n12800_0, n12796_0, n12791_0, n10295_1, n1745, n1737, n1649, n1641, n1633}), .out(n10201), .config_in(config_chain[15873:15868]), .config_rst(config_rst)); 
buffer_wire buffer_10201 (.in(n10201), .out(n10201_0));
mux3 mux_5036 (.in({n12369_0/**/, n12368_0, n663}), .out(n10202), .config_in(config_chain[15875:15874]), .config_rst(config_rst)); 
buffer_wire buffer_10202 (.in(n10202), .out(n10202_0));
mux15 mux_5037 (.in({n13165_1, n13148_0, n13133_0, n13125_1, n13101_0, n13084_0, n13075_0/**/, n13058_0, n13056_0, n10315_1, n2723, n2715, n2627, n2619, n2611}), .out(n10203), .config_in(config_chain[15881:15876]), .config_rst(config_rst)); 
buffer_wire buffer_10203 (.in(n10203), .out(n10203_0));
mux3 mux_5038 (.in({n12389_1, n12298_0, n663}), .out(n10204), .config_in(config_chain[15883:15882]), .config_rst(config_rst)); 
buffer_wire buffer_10204 (.in(n10204), .out(n10204_0));
mux15 mux_5039 (.in({n13425_1/**/, n13399_0, n13394_0, n13385_1, n13370_0, n13361_0, n13344_0, n13318_0, n13307_0, n10335_1, n3701, n3693, n3605, n3597, n3589}), .out(n10205), .config_in(config_chain[15889:15884]), .config_rst(config_rst)); 
buffer_wire buffer_10205 (.in(n10205), .out(n10205_0));
mux3 mux_5040 (.in({n12301_0, n12300_0, n667}), .out(n10206), .config_in(config_chain[15891:15890]), .config_rst(config_rst)); 
buffer_wire buffer_10206 (.in(n10206), .out(n10206_0));
mux15 mux_5041 (.in({n12651_1, n12631_0, n12626_0, n12611_2, n12596_0, n12559_0, n12546_0, n12542_0/**/, n12533_0, n10275_1, n767, n759, n671, n663, n655}), .out(n10207), .config_in(config_chain[15897:15892]), .config_rst(config_rst)); 
buffer_wire buffer_10207 (.in(n10207), .out(n10207_0));
mux3 mux_5042 (.in({n12303_0, n12302_0, n667}), .out(n10208), .config_in(config_chain[15899:15898]), .config_rst(config_rst)); 
buffer_wire buffer_10208 (.in(n10208), .out(n10208_0));
mux15 mux_5043 (.in({n12905_1, n12881_0, n12876_0, n12869_2, n12856_0, n12847_0, n12830_0, n12804_0, n12793_0, n10297_1, n1745, n1737, n1649, n1641, n1633}), .out(n10209), .config_in(config_chain[15905:15900]), .config_rst(config_rst)); 
buffer_wire buffer_10209 (.in(n10209), .out(n10209_0));
mux3 mux_5044 (.in({n12371_0/**/, n12370_0, n667}), .out(n10210), .config_in(config_chain[15907:15906]), .config_rst(config_rst)); 
buffer_wire buffer_10210 (.in(n10210), .out(n10210_0));
mux15 mux_5045 (.in({n13163_1/**/, n13147_0, n13142_0, n13127_2, n13114_0, n13077_0, n13064_0, n13060_0, n13051_0, n10317_1, n2723, n2715, n2627, n2619, n2611}), .out(n10211), .config_in(config_chain[15913:15908]), .config_rst(config_rst)); 
buffer_wire buffer_10211 (.in(n10211), .out(n10211_0));
mux3 mux_5046 (.in({n12391_1, n12306_0, n667}), .out(n10212), .config_in(config_chain[15915:15914]), .config_rst(config_rst)); 
buffer_wire buffer_10212 (.in(n10212), .out(n10212_0));
mux15 mux_5047 (.in({n13423_1, n13408_0, n13393_0, n13387_1, n13363_0, n13346_0, n13337_0, n13326_0, n13320_0, n10337_1/**/, n3701, n3693, n3605, n3597, n3589}), .out(n10213), .config_in(config_chain[15921:15916]), .config_rst(config_rst)); 
buffer_wire buffer_10213 (.in(n10213), .out(n10213_0));
mux3 mux_5048 (.in({n12309_0, n12308_0, n667}), .out(n10214), .config_in(config_chain[15923:15922]), .config_rst(config_rst)); 
buffer_wire buffer_10214 (.in(n10214), .out(n10214_0));
mux15 mux_5049 (.in({n12649_1, n12625_0, n12620_0, n12613_2, n12598_0, n12589_0, n12572_0, n12554_0, n12535_0, n10277_1, n767, n759, n671, n663, n655}), .out(n10215), .config_in(config_chain[15929:15924]), .config_rst(config_rst)); 
buffer_wire buffer_10215 (.in(n10215), .out(n10215_0));
mux3 mux_5050 (.in({n12311_0/**/, n12310_0, n671}), .out(n10216), .config_in(config_chain[15931:15930]), .config_rst(config_rst)); 
buffer_wire buffer_10216 (.in(n10216), .out(n10216_0));
mux15 mux_5051 (.in({n12903_1, n12890_0, n12875_0, n12871_2, n12849_0, n12832_0, n12823_0, n12812_0, n12806_0, n10299_1, n1749, n1741, n1733, n1645, n1637/**/}), .out(n10217), .config_in(config_chain[15937:15932]), .config_rst(config_rst)); 
buffer_wire buffer_10217 (.in(n10217), .out(n10217_0));
mux3 mux_5052 (.in({n12373_0, n12372_0, n671}), .out(n10218), .config_in(config_chain[15939:15938]), .config_rst(config_rst)); 
buffer_wire buffer_10218 (.in(n10218), .out(n10218_0));
mux15 mux_5053 (.in({n13161_1, n13141_0, n13136_0, n13129_2, n13116_0, n13107_0/**/, n13090_0, n13072_0, n13053_0, n10319_1, n2727, n2719, n2711, n2623, n2615}), .out(n10219), .config_in(config_chain[15945:15940]), .config_rst(config_rst)); 
buffer_wire buffer_10219 (.in(n10219), .out(n10219_0));
mux3 mux_5054 (.in({n12393_1, n12314_0, n671}), .out(n10220), .config_in(config_chain[15947:15946]), .config_rst(config_rst)); 
buffer_wire buffer_10220 (.in(n10220), .out(n10220_0));
mux15 mux_5055 (.in({n13421_1, n13407_0, n13402_0, n13389_2, n13376_0, n13339_0, n13334_0, n13322_0, n13313_0, n10339_1, n3705, n3697/**/, n3689, n3601, n3593}), .out(n10221), .config_in(config_chain[15953:15948]), .config_rst(config_rst)); 
buffer_wire buffer_10221 (.in(n10221), .out(n10221_0));
mux3 mux_5056 (.in({n12317_0, n12316_0, n671}), .out(n10222), .config_in(config_chain[15955:15954]), .config_rst(config_rst)); 
buffer_wire buffer_10222 (.in(n10222), .out(n10222_0));
mux15 mux_5057 (.in({n12647_1, n12634_0/**/, n12619_0, n12615_2, n12591_0, n12574_0, n12565_0, n12562_0, n12548_0, n10279_1, n771, n763, n755, n667, n659}), .out(n10223), .config_in(config_chain[15961:15956]), .config_rst(config_rst)); 
buffer_wire buffer_10223 (.in(n10223), .out(n10223_0));
mux3 mux_5058 (.in({n12319_0/**/, n12318_0, n671}), .out(n10224), .config_in(config_chain[15963:15962]), .config_rst(config_rst)); 
buffer_wire buffer_10224 (.in(n10224), .out(n10224_0));
mux15 mux_5059 (.in({n12901_1, n12889_0, n12884_0, n12860_0, n12825_0/**/, n12820_0, n12808_0, n12799_0, n12782_0, n10301_1, n1749, n1741, n1733, n1645, n1637}), .out(n10225), .config_in(config_chain[15969:15964]), .config_rst(config_rst)); 
buffer_wire buffer_10225 (.in(n10225), .out(n10225_0));
mux3 mux_5060 (.in({n12375_0/**/, n12374_0, n755}), .out(n10226), .config_in(config_chain[15971:15970]), .config_rst(config_rst)); 
buffer_wire buffer_10226 (.in(n10226), .out(n10226_0));
mux15 mux_5061 (.in({n13159_1, n13135_0, n13130_0, n13118_0, n13109_0, n13092_0, n13083_0, n13080_0, n13066_0, n10321_1, n2727, n2719, n2711, n2623, n2615}), .out(n10227), .config_in(config_chain[15977:15972]), .config_rst(config_rst)); 
buffer_wire buffer_10227 (.in(n10227), .out(n10227_0));
mux3 mux_5062 (.in({n12395_1, n12322_0/**/, n755}), .out(n10228), .config_in(config_chain[15979:15978]), .config_rst(config_rst)); 
buffer_wire buffer_10228 (.in(n10228), .out(n10228_0));
mux15 mux_5063 (.in({n13419_1, n13401_0, n13396_0, n13378_0, n13369_0, n13352_0, n13342_0, n13315_0, n13298_0, n10341_1, n3705, n3697/**/, n3689, n3601, n3593}), .out(n10229), .config_in(config_chain[15985:15980]), .config_rst(config_rst)); 
buffer_wire buffer_10229 (.in(n10229), .out(n10229_0));
mux3 mux_5064 (.in({n12325_0, n12324_0, n755}), .out(n10230), .config_in(config_chain[15987:15986]), .config_rst(config_rst)); 
buffer_wire buffer_10230 (.in(n10230), .out(n10230_0));
mux15 mux_5065 (.in({n12645_1, n12633_0, n12628_0, n12604_0, n12570_0, n12567_0, n12550_0, n12541_0, n12524_0, n10281_1, n771, n763/**/, n755, n667, n659}), .out(n10231), .config_in(config_chain[15993:15988]), .config_rst(config_rst)); 
buffer_wire buffer_10231 (.in(n10231), .out(n10231_0));
mux3 mux_5066 (.in({n12327_0/**/, n12326_0, n755}), .out(n10232), .config_in(config_chain[15995:15994]), .config_rst(config_rst)); 
buffer_wire buffer_10232 (.in(n10232), .out(n10232_0));
mux15 mux_5067 (.in({n12899_1, n12883_0, n12878_0, n12862_0, n12855_0/**/, n12838_0, n12828_0, n12801_0, n12784_0, n10303_1, n1749, n1741, n1733, n1645, n1637}), .out(n10233), .config_in(config_chain[16001:15996]), .config_rst(config_rst)); 
buffer_wire buffer_10233 (.in(n10233), .out(n10233_0));
mux3 mux_5068 (.in({n12377_0, n12376_0, n755}), .out(n10234), .config_in(config_chain[16003:16002]), .config_rst(config_rst)); 
buffer_wire buffer_10234 (.in(n10234), .out(n10234_0));
mux15 mux_5069 (.in({n13157_1/**/, n13149_0, n13144_0, n13120_0, n13088_0, n13085_0, n13068_0, n13059_0, n13042_0, n10323_1, n2727, n2719, n2711, n2623, n2615}), .out(n10235), .config_in(config_chain[16009:16004]), .config_rst(config_rst)); 
buffer_wire buffer_10235 (.in(n10235), .out(n10235_0));
mux3 mux_5070 (.in({n12397_1, n12330_0, n759/**/}), .out(n10236), .config_in(config_chain[16011:16010]), .config_rst(config_rst)); 
buffer_wire buffer_10236 (.in(n10236), .out(n10236_0));
mux15 mux_5071 (.in({n13417_1, n13395_0, n13390_0, n13380_0, n13371_0, n13354_0, n13350_0, n13345_0, n13328_0, n10343_1, n3705, n3697, n3689, n3601/**/, n3593}), .out(n10237), .config_in(config_chain[16017:16012]), .config_rst(config_rst)); 
buffer_wire buffer_10237 (.in(n10237), .out(n10237_0));
mux3 mux_5072 (.in({n12333_0, n12332_0, n759}), .out(n10238), .config_in(config_chain[16019:16018]), .config_rst(config_rst)); 
buffer_wire buffer_10238 (.in(n10238), .out(n10238_0));
mux15 mux_5073 (.in({n12643_1, n12627_0, n12622_0, n12606_0, n12597_0, n12580_0/**/, n12578_0, n12543_0, n12526_0, n10283_1, n771, n763, n755, n667, n659}), .out(n10239), .config_in(config_chain[16025:16020]), .config_rst(config_rst)); 
buffer_wire buffer_10239 (.in(n10239), .out(n10239_0));
mux3 mux_5074 (.in({n12335_0/**/, n12334_0, n759}), .out(n10240), .config_in(config_chain[16027:16026]), .config_rst(config_rst)); 
buffer_wire buffer_10240 (.in(n10240), .out(n10240_0));
mux15 mux_5075 (.in({n12897_1, n12877_0, n12872_0, n12864_0, n12857_0, n12840_0, n12836_0, n12831_0, n12814_0/**/, n10305_1, n1749, n1741, n1733, n1645, n1637}), .out(n10241), .config_in(config_chain[16033:16028]), .config_rst(config_rst)); 
buffer_wire buffer_10241 (.in(n10241), .out(n10241_0));
mux3 mux_5076 (.in({n12379_0/**/, n12378_0, n759}), .out(n10242), .config_in(config_chain[16035:16034]), .config_rst(config_rst)); 
buffer_wire buffer_10242 (.in(n10242), .out(n10242_0));
mux15 mux_5077 (.in({n13155_1, n13143_0, n13138_0, n13122_0, n13115_0, n13098_0, n13096_0, n13061_0, n13044_0, n10325_1, n2727, n2719, n2711, n2623, n2615}), .out(n10243), .config_in(config_chain[16041:16036]), .config_rst(config_rst)); 
buffer_wire buffer_10243 (.in(n10243), .out(n10243_0));
mux3 mux_5078 (.in({n12399_1, n12338_0, n759}), .out(n10244), .config_in(config_chain[16043:16042]), .config_rst(config_rst)); 
buffer_wire buffer_10244 (.in(n10244), .out(n10244_0));
mux15 mux_5079 (.in({n13415_1, n13409_0, n13404_0, n13382_0, n13358_0, n13347_0, n13330_0, n13321_0, n13304_0, n10345_1/**/, n3705, n3697, n3689, n3601, n3593}), .out(n10245), .config_in(config_chain[16049:16044]), .config_rst(config_rst)); 
buffer_wire buffer_10245 (.in(n10245), .out(n10245_0));
mux3 mux_5080 (.in({n12341_0, n12340_0, n763}), .out(n10246), .config_in(config_chain[16051:16050]), .config_rst(config_rst)); 
buffer_wire buffer_10246 (.in(n10246), .out(n10246_0));
mux15 mux_5081 (.in({n12641_1, n12621_0, n12616_0, n12608_0, n12599_0/**/, n12586_0, n12582_0, n12573_0, n12556_0, n10285_1, n771, n763, n755, n667, n659}), .out(n10247), .config_in(config_chain[16057:16052]), .config_rst(config_rst)); 
buffer_wire buffer_10247 (.in(n10247), .out(n10247_0));
mux3 mux_5082 (.in({n12343_0, n12342_0, n763}), .out(n10248), .config_in(config_chain[16059:16058]), .config_rst(config_rst)); 
buffer_wire buffer_10248 (.in(n10248), .out(n10248_0));
mux15 mux_5083 (.in({n12895_1, n12891_0, n12886_0, n12866_0, n12844_0, n12833_0, n12816_0, n12807_0, n12790_0, n10307_1, n1749, n1741, n1733/**/, n1645, n1637}), .out(n10249), .config_in(config_chain[16065:16060]), .config_rst(config_rst)); 
buffer_wire buffer_10249 (.in(n10249), .out(n10249_0));
mux3 mux_5084 (.in({n12381_0/**/, n12380_0, n763}), .out(n10250), .config_in(config_chain[16067:16066]), .config_rst(config_rst)); 
buffer_wire buffer_10250 (.in(n10250), .out(n10250_0));
mux15 mux_5085 (.in({n13153_1, n13137_0, n13132_0, n13124_0, n13117_0, n13104_0, n13100_0, n13091_0, n13074_0, n10327_1, n2727/**/, n2719, n2711, n2623, n2615}), .out(n10251), .config_in(config_chain[16073:16068]), .config_rst(config_rst)); 
buffer_wire buffer_10251 (.in(n10251), .out(n10251_0));
mux3 mux_5086 (.in({n12401_1/**/, n12346_0, n763}), .out(n10252), .config_in(config_chain[16075:16074]), .config_rst(config_rst)); 
buffer_wire buffer_10252 (.in(n10252), .out(n10252_0));
mux15 mux_5087 (.in({n13413_1, n13403_0, n13398_0, n13384_0, n13377_0, n13366_0, n13360_0, n13323_0, n13306_0, n10347_1, n3705, n3697, n3689/**/, n3601, n3593}), .out(n10253), .config_in(config_chain[16081:16076]), .config_rst(config_rst)); 
buffer_wire buffer_10253 (.in(n10253), .out(n10253_0));
mux3 mux_5088 (.in({n12349_0, n12348_0, n763/**/}), .out(n10254), .config_in(config_chain[16083:16082]), .config_rst(config_rst)); 
buffer_wire buffer_10254 (.in(n10254), .out(n10254_0));
mux15 mux_5089 (.in({n12639_1, n12635_0, n12630_0, n12610_0, n12594_0, n12575_0, n12558_0, n12549_0, n12532_0, n10287_1, n771, n763/**/, n755, n667, n659}), .out(n10255), .config_in(config_chain[16089:16084]), .config_rst(config_rst)); 
buffer_wire buffer_10255 (.in(n10255), .out(n10255_0));
mux3 mux_5090 (.in({n12351_1, n12350_0, n767}), .out(n10256), .config_in(config_chain[16091:16090]), .config_rst(config_rst)); 
buffer_wire buffer_10256 (.in(n10256), .out(n10256_0));
mux13 mux_5091 (.in({n13939_1, n13920_0, n13911_0, n13906_0, n13896_0, n13883_0, n13876_0, n13853_0, n10389_0, n5657, n5649, n5561, n5553}), .out(n10257), .config_in(config_chain[16097:16092]), .config_rst(config_rst)); 
buffer_wire buffer_10257 (.in(n10257), .out(n10257_0));
mux3 mux_5092 (.in({n12353_2, n12352_0, n767}), .out(n10258), .config_in(config_chain[16099:16098]), .config_rst(config_rst)); 
buffer_wire buffer_10258 (.in(n10258), .out(n10258_0));
mux13 mux_5093 (.in({n14205_1, n14200_0, n14195_0, n14175_0, n14162_0, n14140_0, n14117_0, n14110_0, n10411_0, n6635, n6627, n6539, n6531}), .out(n10259), .config_in(config_chain[16105:16100]), .config_rst(config_rst)); 
buffer_wire buffer_10259 (.in(n10259), .out(n10259_0));
mux3 mux_5094 (.in({n12355_2, n12354_0, n767}), .out(n10260), .config_in(config_chain[16107:16106]), .config_rst(config_rst)); 
buffer_wire buffer_10260 (.in(n10260), .out(n10260_0));
mux13 mux_5095 (.in({n14469_1/**/, n14456_0, n14451_0, n14439_0, n14432_0, n14428_0, n14409_0, n14374_0, n10433_0, n7613, n7605, n7517, n7509}), .out(n10261), .config_in(config_chain[16113:16108]), .config_rst(config_rst)); 
buffer_wire buffer_10261 (.in(n10261), .out(n10261_0));
mux3 mux_5096 (.in({n12357_2, n12356_0, n767}), .out(n10262), .config_in(config_chain[16115:16114]), .config_rst(config_rst)); 
buffer_wire buffer_10262 (.in(n10262), .out(n10262_0));
mux3 mux_5097 (.in({n14749_2/**/, n14700_0, n8591}), .out(n10263), .config_in(config_chain[16117:16116]), .config_rst(config_rst)); 
buffer_wire buffer_10263 (.in(n10263), .out(n10263_0));
mux3 mux_5098 (.in({n12359_2/**/, n12358_0, n767}), .out(n10264), .config_in(config_chain[16119:16118]), .config_rst(config_rst)); 
buffer_wire buffer_10264 (.in(n10264), .out(n10264_0));
mux3 mux_5099 (.in({n14703_0, n14702_0, n8591}), .out(n10265), .config_in(config_chain[16121:16120]), .config_rst(config_rst)); 
buffer_wire buffer_10265 (.in(n10265), .out(n10265_0));
mux3 mux_5100 (.in({n12361_2, n12360_0, n771}), .out(n10266), .config_in(config_chain[16123:16122]), .config_rst(config_rst)); 
buffer_wire buffer_10266 (.in(n10266), .out(n10266_0));
mux3 mux_5101 (.in({n14705_0, n14704_0/**/, n8595}), .out(n10267), .config_in(config_chain[16125:16124]), .config_rst(config_rst)); 
buffer_wire buffer_10267 (.in(n10267), .out(n10267_0));
mux16 mux_5102 (.in({n12655_1/**/, n12628_0, n12625_0, n12613_2, n12604_0, n12594_0, n12589_0, n12550_0, n12535_0, n12524_0, n10182_0, n1745, n1737, n1649, n1641, n1633}), .out(n10268), .config_in(config_chain[16131:16126]), .config_rst(config_rst)); 
buffer_wire buffer_10268 (.in(n10268), .out(n10268_0));
mux16 mux_5103 (.in({n13673_1, n13665_0, n13660_0, n13648_0, n13641_0, n13638_0, n13624_0, n13587_0, n13570_0/**/, n13561_0, n10349_1, n4679, n4671, n4583, n4575, n4567}), .out(n10269), .config_in(config_chain[16137:16132]), .config_rst(config_rst)); 
buffer_wire buffer_10269 (.in(n10269), .out(n10269_0));
mux16 mux_5104 (.in({n12637_1, n12622_0, n12619_0, n12615_2, n12606_0, n12591_0/**/, n12586_0, n12580_0, n12565_0, n12526_0, n10190_0, n1745, n1737, n1649, n1641, n1633}), .out(n10270), .config_in(config_chain[16143:16138]), .config_rst(config_rst)); 
buffer_wire buffer_10270 (.in(n10270), .out(n10270_0));
mux16 mux_5105 (.in({n13691_1, n13659_0, n13654_0, n13650_0, n13643_0, n13626_0, n13617_0, n13600_0, n13566_0, n13563_0, n10351_1, n4679, n4671, n4583, n4575/**/, n4567}), .out(n10271), .config_in(config_chain[16149:16144]), .config_rst(config_rst)); 
buffer_wire buffer_10271 (.in(n10271), .out(n10271_0));
mux15 mux_5106 (.in({n12639_1, n12633_0, n12616_0, n12608_0, n12582_0, n12578_0, n12567_0/**/, n12556_0, n12541_0, n10198_0, n1745, n1737, n1649, n1641, n1633}), .out(n10272), .config_in(config_chain[16155:16150]), .config_rst(config_rst)); 
buffer_wire buffer_10272 (.in(n10272), .out(n10272_0));
mux15 mux_5107 (.in({n13689_1, n13668_0, n13653_0, n13645_0, n13619_0, n13602_0, n13593_0, n13576_0, n13574_0, n10353_1, n4679, n4671, n4583/**/, n4575, n4567}), .out(n10273), .config_in(config_chain[16161:16156]), .config_rst(config_rst)); 
buffer_wire buffer_10273 (.in(n10273), .out(n10273_0));
mux15 mux_5108 (.in({n12641_1, n12630_0, n12627_0, n12610_0, n12597_0, n12570_0, n12558_0/**/, n12543_0, n12532_0, n10206_0, n1745, n1737, n1649, n1641, n1633}), .out(n10274), .config_in(config_chain[16167:16162]), .config_rst(config_rst)); 
buffer_wire buffer_10274 (.in(n10274), .out(n10274_0));
mux15 mux_5109 (.in({n13687_1, n13667_0, n13662_0, n13647_1, n13632_0, n13595_0, n13582_0, n13578_0, n13569_0, n10355_1, n4679, n4671, n4583, n4575, n4567}), .out(n10275), .config_in(config_chain[16173:16168]), .config_rst(config_rst)); 
buffer_wire buffer_10275 (.in(n10275), .out(n10275_0));
mux15 mux_5110 (.in({n12643_1, n12624_0, n12621_0, n12612_0, n12599_0, n12588_0, n12573_0, n12562_0, n12534_0, n10214_0, n1745, n1737, n1649, n1641, n1633}), .out(n10276), .config_in(config_chain[16179:16174]), .config_rst(config_rst)); 
buffer_wire buffer_10276 (.in(n10276), .out(n10276_0));
mux15 mux_5111 (.in({n13685_1, n13661_0, n13656_0, n13649_1, n13634_0, n13625_0, n13608_0, n13590_0, n13571_0, n10357_1, n4679, n4671, n4583, n4575, n4567}), .out(n10277), .config_in(config_chain[16185:16180]), .config_rst(config_rst)); 
buffer_wire buffer_10277 (.in(n10277), .out(n10277_0));
mux15 mux_5112 (.in({n12645_1, n12635_0, n12618_0, n12614_0, n12590_0, n12575_0, n12564_0, n12554_0, n12549_0/**/, n10222_0, n1749, n1741, n1733, n1645, n1637}), .out(n10278), .config_in(config_chain[16191:16186]), .config_rst(config_rst)); 
buffer_wire buffer_10278 (.in(n10278), .out(n10278_0));
mux15 mux_5113 (.in({n13683_1, n13670_0, n13655_0, n13651_1, n13627_0, n13610_0, n13601_0, n13598_0, n13584_0/**/, n10359_1, n4683, n4675, n4667, n4579, n4571}), .out(n10279), .config_in(config_chain[16197:16192]), .config_rst(config_rst)); 
buffer_wire buffer_10279 (.in(n10279), .out(n10279_0));
mux15 mux_5114 (.in({n12647_1, n12632_0, n12629_0, n12605_1, n12566_0, n12551_0, n12546_0, n12540_0, n12525_0, n10230_0, n1749, n1741, n1733, n1645, n1637/**/}), .out(n10280), .config_in(config_chain[16203:16198]), .config_rst(config_rst)); 
buffer_wire buffer_10280 (.in(n10280), .out(n10280_0));
mux15 mux_5115 (.in({n13681_1, n13669_0, n13664_0, n13640_0, n13606_0, n13603_0, n13586_0, n13577_0, n13560_0, n10361_1, n4683, n4675/**/, n4667, n4579, n4571}), .out(n10281), .config_in(config_chain[16209:16204]), .config_rst(config_rst)); 
buffer_wire buffer_10281 (.in(n10281), .out(n10281_0));
mux15 mux_5116 (.in({n12649_1, n12626_0, n12623_0, n12607_1, n12596_0, n12581_0, n12542_0, n12538_0, n12527_0/**/, n10238_0, n1749, n1741, n1733, n1645, n1637}), .out(n10282), .config_in(config_chain[16215:16210]), .config_rst(config_rst)); 
buffer_wire buffer_10282 (.in(n10282), .out(n10282_0));
mux15 mux_5117 (.in({n13679_1, n13663_0, n13658_0, n13642_0, n13633_0, n13616_0, n13614_0, n13579_0, n13562_0, n10363_1, n4683, n4675, n4667/**/, n4579, n4571}), .out(n10283), .config_in(config_chain[16221:16216]), .config_rst(config_rst)); 
buffer_wire buffer_10283 (.in(n10283), .out(n10283_0));
mux15 mux_5118 (.in({n12651_1, n12620_0, n12617_0, n12609_2, n12598_0, n12583_0, n12572_0, n12557_0, n12530_0, n10246_0, n1749, n1741, n1733/**/, n1645, n1637}), .out(n10284), .config_in(config_chain[16227:16222]), .config_rst(config_rst)); 
buffer_wire buffer_10284 (.in(n10284), .out(n10284_0));
mux15 mux_5119 (.in({n13677_1, n13657_0, n13652_0, n13644_0, n13635_0, n13622_0, n13618_0, n13609_0, n13592_0, n10365_1, n4683, n4675, n4667, n4579, n4571}), .out(n10285), .config_in(config_chain[16233:16228]), .config_rst(config_rst)); 
buffer_wire buffer_10285 (.in(n10285), .out(n10285_0));
mux15 mux_5120 (.in({n12653_1, n12634_0, n12631_0, n12611_2, n12602_0, n12574_0, n12559_0, n12548_0, n12533_0/**/, n10254_0, n1749, n1741, n1733, n1645, n1637}), .out(n10286), .config_in(config_chain[16239:16234]), .config_rst(config_rst)); 
buffer_wire buffer_10286 (.in(n10286), .out(n10286_0));
mux15 mux_5121 (.in({n13675_1, n13671_0, n13666_0, n13646_0, n13630_0, n13611_0, n13594_0, n13585_0, n13568_0, n10367_1, n4683, n4675, n4667, n4579, n4571}), .out(n10287), .config_in(config_chain[16245:16240]), .config_rst(config_rst)); 
buffer_wire buffer_10287 (.in(n10287), .out(n10287_0));
mux16 mux_5122 (.in({n12911_1, n12884_0, n12881_0, n12869_2, n12860_0, n12847_0, n12844_0, n12808_0, n12793_0, n12782_0, n10176_0, n2723, n2715, n2627, n2619/**/, n2611}), .out(n10288), .config_in(config_chain[16251:16246]), .config_rst(config_rst)); 
buffer_wire buffer_10288 (.in(n10288), .out(n10288_0));
mux15 mux_5123 (.in({n13937_1, n13928_0, n13923_0, n13913_1/**/, n13908_0, n13904_0, n13885_0, n13850_0, n13827_0, n10369_0, n5657, n5649, n5561, n5553, n5545}), .out(n10289), .config_in(config_chain[16257:16252]), .config_rst(config_rst)); 
buffer_wire buffer_10289 (.in(n10289), .out(n10289_0));
mux16 mux_5124 (.in({n12893_1, n12878_0, n12875_0, n12871_2, n12862_0, n12849_0, n12838_0, n12836_0, n12823_0, n12784_0, n10184_0, n2723, n2715, n2627, n2619/**/, n2611}), .out(n10290), .config_in(config_chain[16263:16258]), .config_rst(config_rst)); 
buffer_wire buffer_10290 (.in(n10290), .out(n10290_0));
mux15 mux_5125 (.in({n13957_2, n13931_0, n13915_1, n13910_0, n13882_0, n13859_0, n13852_0, n13829_0, n13824_0, n10371_0, n5661, n5649, n5561, n5553, n5545/**/}), .out(n10291), .config_in(config_chain[16269:16264]), .config_rst(config_rst)); 
buffer_wire buffer_10291 (.in(n10291), .out(n10291_0));
mux15 mux_5126 (.in({n12895_1, n12889_0/**/, n12872_0, n12864_0, n12840_0, n12828_0, n12825_0, n12814_0, n12799_0, n10192_0, n2723, n2715, n2627, n2619, n2611}), .out(n10292), .config_in(config_chain[16275:16270]), .config_rst(config_rst)); 
buffer_wire buffer_10292 (.in(n10292), .out(n10292_0));
mux15 mux_5127 (.in({n13955_1, n13922_0, n13917_0, n13912_0, n13891_0, n13884_0, n13861_0, n13832_0, n13826_0, n10373_0, n5661, n5653, n5561, n5553, n5545/**/}), .out(n10293), .config_in(config_chain[16281:16276]), .config_rst(config_rst)); 
buffer_wire buffer_10293 (.in(n10293), .out(n10293_0));
mux15 mux_5128 (.in({n12897_1, n12886_0, n12883_0, n12866_0, n12855_0, n12820_0, n12816_0, n12801_0, n12790_0, n10200_0, n2723, n2715/**/, n2627, n2619, n2611}), .out(n10294), .config_in(config_chain[16287:16282]), .config_rst(config_rst)); 
buffer_wire buffer_10294 (.in(n10294), .out(n10294_0));
mux15 mux_5129 (.in({n13953_1, n13930_0, n13925_0/**/, n13914_0, n13893_0, n13858_0, n13840_0, n13835_0, n13828_0, n10375_0, n5661, n5653, n5645, n5553, n5545}), .out(n10295), .config_in(config_chain[16293:16288]), .config_rst(config_rst)); 
buffer_wire buffer_10295 (.in(n10295), .out(n10295_0));
mux15 mux_5130 (.in({n12899_1, n12880_0, n12877_0, n12868_0, n12857_0, n12846_0, n12831_0, n12812_0, n12792_0, n10208_0, n2723, n2715/**/, n2627, n2619, n2611}), .out(n10296), .config_in(config_chain[16299:16294]), .config_rst(config_rst)); 
buffer_wire buffer_10296 (.in(n10296), .out(n10296_0));
mux14 mux_5131 (.in({n13951_1, n13933_0, n13916_0, n13890_0, n13867_0, n13860_0, n13848_0/**/, n13837_0, n10377_0, n5661, n5653, n5645, n5557, n5545}), .out(n10297), .config_in(config_chain[16305:16300]), .config_rst(config_rst)); 
buffer_wire buffer_10297 (.in(n10297), .out(n10297_0));
mux15 mux_5132 (.in({n12901_1, n12891_0, n12874_0, n12870_0, n12848_0, n12833_0, n12822_0, n12807_0, n12804_0, n10216_0/**/, n2727, n2719, n2711, n2623, n2615}), .out(n10298), .config_in(config_chain[16311:16306]), .config_rst(config_rst)); 
buffer_wire buffer_10298 (.in(n10298), .out(n10298_0));
mux14 mux_5133 (.in({n13949_1, n13924_0, n13919_0, n13899_0/**/, n13892_0, n13869_0, n13856_0, n13834_0, n10379_0, n5661, n5653, n5645, n5557, n5549}), .out(n10299), .config_in(config_chain[16317:16312]), .config_rst(config_rst)); 
buffer_wire buffer_10299 (.in(n10299), .out(n10299_0));
mux15 mux_5134 (.in({n12903_1, n12888_0, n12885_0, n12861_1, n12824_0, n12809_0, n12798_0, n12796_0, n12783_0/**/, n10224_0, n2727, n2719, n2711, n2623, n2615}), .out(n10300), .config_in(config_chain[16323:16318]), .config_rst(config_rst)); 
buffer_wire buffer_10300 (.in(n10300), .out(n10300_0));
mux13 mux_5135 (.in({n13947_1, n13932_0, n13927_0, n13901_0, n13866_0, n13864_0/**/, n13843_0, n13836_0, n10381_0, n5653, n5645, n5557, n5549}), .out(n10301), .config_in(config_chain[16329:16324]), .config_rst(config_rst)); 
buffer_wire buffer_10301 (.in(n10301), .out(n10301_0));
mux15 mux_5136 (.in({n12905_1, n12882_0, n12879_0, n12863_1, n12854_0/**/, n12839_0, n12800_0, n12788_0, n12785_0, n10232_0, n2727, n2719, n2711, n2623, n2615}), .out(n10302), .config_in(config_chain[16335:16330]), .config_rst(config_rst)); 
buffer_wire buffer_10302 (.in(n10302), .out(n10302_0));
mux13 mux_5137 (.in({n13945_1, n13935_0/**/, n13918_0, n13898_0, n13875_0, n13872_0, n13868_0, n13845_0, n10383_0, n5657, n5645, n5557, n5549}), .out(n10303), .config_in(config_chain[16341:16336]), .config_rst(config_rst)); 
buffer_wire buffer_10303 (.in(n10303), .out(n10303_0));
mux15 mux_5138 (.in({n12907_1, n12876_0, n12873_0, n12865_1, n12856_0, n12841_0, n12830_0, n12815_0, n12780_0, n10240_0/**/, n2727, n2719, n2711, n2623, n2615}), .out(n10304), .config_in(config_chain[16347:16342]), .config_rst(config_rst)); 
buffer_wire buffer_10304 (.in(n10304), .out(n10304_0));
mux13 mux_5139 (.in({n13943_1, n13926_0, n13921_0, n13907_0, n13900_0, n13880_0, n13877_0, n13842_0, n10385_0, n5657, n5649/**/, n5557, n5549}), .out(n10305), .config_in(config_chain[16353:16348]), .config_rst(config_rst)); 
buffer_wire buffer_10305 (.in(n10305), .out(n10305_0));
mux15 mux_5140 (.in({n12909_1, n12890_0, n12887_0, n12867_2, n12852_0, n12832_0, n12817_0, n12806_0/**/, n12791_0, n10248_0, n2727, n2719, n2711, n2623, n2615}), .out(n10306), .config_in(config_chain[16359:16354]), .config_rst(config_rst)); 
buffer_wire buffer_10306 (.in(n10306), .out(n10306_0));
mux13 mux_5141 (.in({n13941_1, n13934_0, n13929_0, n13909_0, n13888_0, n13874_0, n13851_0, n13844_0, n10387_0, n5657, n5649, n5561, n5549}), .out(n10307), .config_in(config_chain[16365:16360]), .config_rst(config_rst)); 
buffer_wire buffer_10307 (.in(n10307), .out(n10307_0));
mux16 mux_5142 (.in({n13169_1, n13147_0/**/, n13130_0, n13127_2, n13118_0, n13104_0, n13092_0, n13077_0, n13066_0, n13051_0, n10178_0, n3701, n3693, n3605, n3597, n3589}), .out(n10308), .config_in(config_chain[16371:16366]), .config_rst(config_rst)); 
buffer_wire buffer_10308 (.in(n10308), .out(n10308_0));
mux15 mux_5143 (.in({n14203_1, n14186_0, n14181_0/**/, n14177_0, n14172_0, n14170_0, n14149_0, n14142_0, n14119_0, n10391_0, n6635, n6627, n6539, n6531, n6523}), .out(n10309), .config_in(config_chain[16377:16372]), .config_rst(config_rst)); 
buffer_wire buffer_10309 (.in(n10309), .out(n10309_0));
mux16 mux_5144 (.in({n13151_1, n13144_0, n13141_0, n13129_2, n13120_0, n13107_0, n13096_0, n13068_0, n13053_0, n13042_0, n10186_0, n3701, n3693, n3605, n3597, n3589/**/}), .out(n10310), .config_in(config_chain[16383:16378]), .config_rst(config_rst)); 
buffer_wire buffer_10310 (.in(n10310), .out(n10310_0));
mux15 mux_5145 (.in({n14223_2, n14194_0, n14189_0, n14179_1, n14174_0, n14151_0/**/, n14116_0, n14093_0, n14090_0, n10393_0, n6639, n6627, n6539, n6531, n6523}), .out(n10311), .config_in(config_chain[16389:16384]), .config_rst(config_rst)); 
buffer_wire buffer_10311 (.in(n10311), .out(n10311_0));
mux15 mux_5146 (.in({n13153_1, n13138_0, n13135_0, n13122_0, n13109_0, n13098_0/**/, n13088_0, n13083_0, n13044_0, n10194_0, n3701, n3693, n3605, n3597, n3589}), .out(n10312), .config_in(config_chain[16395:16390]), .config_rst(config_rst)); 
buffer_wire buffer_10312 (.in(n10312), .out(n10312_0));
mux15 mux_5147 (.in({n14221_1/**/, n14197_0, n14180_0, n14176_0, n14148_0, n14125_0, n14118_0, n14098_0, n14095_0, n10395_0, n6639, n6631, n6539, n6531, n6523}), .out(n10313), .config_in(config_chain[16401:16396]), .config_rst(config_rst)); 
buffer_wire buffer_10313 (.in(n10313), .out(n10313_0));
mux15 mux_5148 (.in({n13155_1, n13149_0, n13132_0, n13124_0, n13100_0, n13085_0, n13080_0, n13074_0, n13059_0, n10202_0, n3701, n3693/**/, n3605, n3597, n3589}), .out(n10314), .config_in(config_chain[16407:16402]), .config_rst(config_rst)); 
buffer_wire buffer_10314 (.in(n10314), .out(n10314_0));
mux15 mux_5149 (.in({n14219_1, n14188_0/**/, n14183_0, n14178_0, n14157_0, n14150_0, n14127_0, n14106_0, n14092_0, n10397_0, n6639, n6631, n6623, n6531, n6523}), .out(n10315), .config_in(config_chain[16413:16408]), .config_rst(config_rst)); 
buffer_wire buffer_10315 (.in(n10315), .out(n10315_0));
mux15 mux_5150 (.in({n13157_1, n13146_0, n13143_0, n13126_0, n13115_0, n13076_0, n13072_0, n13061_0, n13050_0, n10210_0, n3701, n3693, n3605, n3597, n3589/**/}), .out(n10316), .config_in(config_chain[16419:16414]), .config_rst(config_rst)); 
buffer_wire buffer_10316 (.in(n10316), .out(n10316_0));
mux14 mux_5151 (.in({n14217_1, n14196_0, n14191_0, n14159_0, n14124_0, n14114_0, n14101_0, n14094_0, n10399_0, n6639, n6631, n6623, n6535, n6523}), .out(n10317), .config_in(config_chain[16425:16420]), .config_rst(config_rst)); 
buffer_wire buffer_10317 (.in(n10317), .out(n10317_0));
mux15 mux_5152 (.in({n13159_1, n13140_0, n13137_0/**/, n13128_0, n13117_0, n13106_0, n13091_0, n13064_0, n13052_0, n10218_0, n3705, n3697, n3689, n3601, n3593}), .out(n10318), .config_in(config_chain[16431:16426]), .config_rst(config_rst)); 
buffer_wire buffer_10318 (.in(n10318), .out(n10318_0));
mux14 mux_5153 (.in({n14215_1, n14199_0, n14182_0/**/, n14156_0, n14133_0, n14126_0, n14122_0, n14103_0, n10401_0, n6639, n6631, n6623, n6535, n6527}), .out(n10319), .config_in(config_chain[16437:16432]), .config_rst(config_rst)); 
buffer_wire buffer_10319 (.in(n10319), .out(n10319_0));
mux15 mux_5154 (.in({n13161_1, n13134_0, n13131_0, n13119_0, n13108_0, n13093_0, n13082_0, n13067_0, n13056_0, n10226_0/**/, n3705, n3697, n3689, n3601, n3593}), .out(n10320), .config_in(config_chain[16443:16438]), .config_rst(config_rst)); 
buffer_wire buffer_10320 (.in(n10320), .out(n10320_0));
mux13 mux_5155 (.in({n14213_1, n14190_0, n14185_0, n14165_0, n14158_0, n14135_0, n14130_0/**/, n14100_0, n10403_0, n6631, n6623, n6535, n6527}), .out(n10321), .config_in(config_chain[16449:16444]), .config_rst(config_rst)); 
buffer_wire buffer_10321 (.in(n10321), .out(n10321_0));
mux15 mux_5156 (.in({n13163_1/**/, n13148_0, n13145_0, n13121_1, n13084_0, n13069_0, n13058_0, n13048_0, n13043_0, n10234_0, n3705, n3697, n3689, n3601, n3593}), .out(n10322), .config_in(config_chain[16455:16450]), .config_rst(config_rst)); 
buffer_wire buffer_10322 (.in(n10322), .out(n10322_0));
mux13 mux_5157 (.in({n14211_1, n14198_0, n14193_0, n14167_0, n14138_0, n14132_0, n14109_0, n14102_0, n10405_0, n6635, n6623, n6535/**/, n6527}), .out(n10323), .config_in(config_chain[16461:16456]), .config_rst(config_rst)); 
buffer_wire buffer_10323 (.in(n10323), .out(n10323_0));
mux15 mux_5158 (.in({n13165_1, n13142_0, n13139_0, n13123_1, n13114_0, n13099_0, n13060_0, n13045_0, n13040_0, n10242_0/**/, n3705, n3697, n3689, n3601, n3593}), .out(n10324), .config_in(config_chain[16467:16462]), .config_rst(config_rst)); 
buffer_wire buffer_10324 (.in(n10324), .out(n10324_0));
mux13 mux_5159 (.in({n14209_1, n14201_2, n14184_0, n14164_0, n14146_0, n14141_0, n14134_0, n14111_0, n10407_0, n6635, n6627, n6535, n6527/**/}), .out(n10325), .config_in(config_chain[16473:16468]), .config_rst(config_rst)); 
buffer_wire buffer_10325 (.in(n10325), .out(n10325_0));
mux15 mux_5160 (.in({n13167_1, n13136_0, n13133_0, n13125_1, n13116_0, n13112_0, n13101_0, n13090_0/**/, n13075_0, n10250_0, n3705, n3697, n3689, n3601, n3593}), .out(n10326), .config_in(config_chain[16479:16474]), .config_rst(config_rst)); 
buffer_wire buffer_10326 (.in(n10326), .out(n10326_0));
mux13 mux_5161 (.in({n14207_1/**/, n14192_0, n14187_0, n14173_0, n14166_0, n14154_0, n14143_0, n14108_0, n10409_0, n6635, n6627, n6539, n6527}), .out(n10327), .config_in(config_chain[16485:16480]), .config_rst(config_rst)); 
buffer_wire buffer_10327 (.in(n10327), .out(n10327_0));
mux16 mux_5162 (.in({n13429_1, n13396_0/**/, n13393_0, n13387_1, n13378_0, n13366_0, n13363_0, n13352_0, n13337_0, n13298_0, n10180_1, n4679, n4671, n4583, n4575, n4567}), .out(n10328), .config_in(config_chain[16491:16486]), .config_rst(config_rst)); 
buffer_wire buffer_10328 (.in(n10328), .out(n10328_0));
mux15 mux_5163 (.in({n14467_1, n14464_0, n14459_0, n14441_0, n14436_0, n14406_0, n14383_0, n14376_0/**/, n14353_0, n10413_0, n7613, n7605, n7517, n7509, n7501}), .out(n10329), .config_in(config_chain[16497:16492]), .config_rst(config_rst)); 
buffer_wire buffer_10329 (.in(n10329), .out(n10329_0));
mux16 mux_5164 (.in({n13411_1, n13407_0/**/, n13390_0, n13389_2, n13380_0, n13358_0, n13354_0, n13339_0, n13328_0, n13313_0, n10188_1, n4679, n4671, n4583, n4575, n4567}), .out(n10330), .config_in(config_chain[16503:16498]), .config_rst(config_rst)); 
buffer_wire buffer_10330 (.in(n10330), .out(n10330_0));
mux15 mux_5165 (.in({n14487_2, n14450_0, n14445_0, n14443_0, n14438_0, n14415_0, n14408_0/**/, n14385_0, n14356_0, n10415_0, n7617, n7605, n7517, n7509, n7501}), .out(n10331), .config_in(config_chain[16509:16504]), .config_rst(config_rst)); 
buffer_wire buffer_10331 (.in(n10331), .out(n10331_0));
mux15 mux_5166 (.in({n13413_1, n13404_0, n13401_0, n13382_0, n13369_0, n13350_0, n13330_0, n13315_0, n13304_0/**/, n10196_1, n4679, n4671, n4583, n4575, n4567}), .out(n10332), .config_in(config_chain[16515:16510]), .config_rst(config_rst)); 
buffer_wire buffer_10332 (.in(n10332), .out(n10332_0));
mux15 mux_5167 (.in({n14485_1, n14458_0, n14453_0, n14440_0, n14417_0, n14382_0, n14364_0, n14359_0, n14352_0, n10417_0/**/, n7617, n7609, n7517, n7509, n7501}), .out(n10333), .config_in(config_chain[16521:16516]), .config_rst(config_rst)); 
buffer_wire buffer_10333 (.in(n10333), .out(n10333_0));
mux15 mux_5168 (.in({n13415_1, n13398_0, n13395_0, n13384_0, n13371_0, n13360_0, n13345_0, n13342_0, n13306_0, n10204_1, n4679, n4671/**/, n4583, n4575, n4567}), .out(n10334), .config_in(config_chain[16527:16522]), .config_rst(config_rst)); 
buffer_wire buffer_10334 (.in(n10334), .out(n10334_0));
mux15 mux_5169 (.in({n14483_1, n14461_0, n14444_0, n14442_0, n14414_0, n14391_0, n14384_0, n14372_0, n14361_0, n10419_0/**/, n7617, n7609, n7601, n7509, n7501}), .out(n10335), .config_in(config_chain[16533:16528]), .config_rst(config_rst)); 
buffer_wire buffer_10335 (.in(n10335), .out(n10335_0));
mux15 mux_5170 (.in({n13417_1, n13409_0, n13392_0, n13386_0, n13362_0, n13347_0, n13336_0, n13334_0, n13321_0/**/, n10212_1, n4679, n4671, n4583, n4575, n4567}), .out(n10336), .config_in(config_chain[16539:16534]), .config_rst(config_rst)); 
buffer_wire buffer_10336 (.in(n10336), .out(n10336_0));
mux14 mux_5171 (.in({n14481_1, n14452_0, n14447_0, n14423_0, n14416_0, n14393_0, n14380_0, n14358_0, n10421_0, n7617, n7609/**/, n7601, n7513, n7501}), .out(n10337), .config_in(config_chain[16545:16540]), .config_rst(config_rst)); 
buffer_wire buffer_10337 (.in(n10337), .out(n10337_0));
mux15 mux_5172 (.in({n13419_1, n13406_0, n13403_0, n13388_0, n13377_0, n13338_0, n13326_0, n13323_0, n13312_0, n10220_1, n4683, n4675, n4667/**/, n4579, n4571}), .out(n10338), .config_in(config_chain[16551:16546]), .config_rst(config_rst)); 
buffer_wire buffer_10338 (.in(n10338), .out(n10338_0));
mux14 mux_5173 (.in({n14479_1, n14460_0, n14455_0, n14425_0, n14390_0, n14388_0, n14367_0, n14360_0, n10423_0, n7617, n7609, n7601/**/, n7513, n7505}), .out(n10339), .config_in(config_chain[16557:16552]), .config_rst(config_rst)); 
buffer_wire buffer_10339 (.in(n10339), .out(n10339_0));
mux15 mux_5174 (.in({n13421_1, n13400_0, n13397_0, n13379_0, n13368_0, n13353_0, n13318_0, n13314_0, n13299_0, n10228_1, n4683, n4675, n4667, n4579/**/, n4571}), .out(n10340), .config_in(config_chain[16563:16558]), .config_rst(config_rst)); 
buffer_wire buffer_10340 (.in(n10340), .out(n10340_0));
mux13 mux_5175 (.in({n14477_1, n14463_0, n14446_0, n14422_0, n14399_0, n14396_0, n14392_0, n14369_0, n10425_0, n7609, n7601/**/, n7513, n7505}), .out(n10341), .config_in(config_chain[16569:16564]), .config_rst(config_rst)); 
buffer_wire buffer_10341 (.in(n10341), .out(n10341_0));
mux15 mux_5176 (.in({n13423_1, n13394_0, n13391_0, n13381_0, n13370_0, n13355_0, n13344_0, n13329_0, n13310_0, n10236_1, n4683, n4675, n4667/**/, n4579, n4571}), .out(n10342), .config_in(config_chain[16575:16570]), .config_rst(config_rst)); 
buffer_wire buffer_10342 (.in(n10342), .out(n10342_0));
mux13 mux_5177 (.in({n14475_1, n14454_0, n14449_0, n14431_0, n14424_0, n14404_0, n14401_0, n14366_0, n10427_0, n7613, n7601, n7513/**/, n7505}), .out(n10343), .config_in(config_chain[16581:16576]), .config_rst(config_rst)); 
buffer_wire buffer_10343 (.in(n10343), .out(n10343_0));
mux15 mux_5178 (.in({n13425_1, n13408_0/**/, n13405_0, n13383_1, n13346_0, n13331_0, n13320_0, n13305_0, n13302_0, n10244_1, n4683, n4675, n4667, n4579, n4571}), .out(n10344), .config_in(config_chain[16587:16582]), .config_rst(config_rst)); 
buffer_wire buffer_10344 (.in(n10344), .out(n10344_0));
mux13 mux_5179 (.in({n14473_1, n14462_0, n14457_0, n14433_2, n14412_0, n14398_0, n14375_0, n14368_0, n10429_0/**/, n7613, n7605, n7513, n7505}), .out(n10345), .config_in(config_chain[16593:16588]), .config_rst(config_rst)); 
buffer_wire buffer_10345 (.in(n10345), .out(n10345_0));
mux15 mux_5180 (.in({n13427_1, n13402_0, n13399_0, n13385_1, n13376_0, n13374_0/**/, n13361_0, n13322_0, n13307_0, n10252_1, n4683, n4675, n4667, n4579, n4571}), .out(n10346), .config_in(config_chain[16599:16594]), .config_rst(config_rst)); 
buffer_wire buffer_10346 (.in(n10346), .out(n10346_0));
mux13 mux_5181 (.in({n14471_1, n14465_2, n14448_0, n14430_0, n14420_0, n14407_0, n14400_0, n14377_0, n10431_0/**/, n7613, n7605, n7517, n7505}), .out(n10347), .config_in(config_chain[16605:16600]), .config_rst(config_rst)); 
buffer_wire buffer_10347 (.in(n10347), .out(n10347_0));
mux16 mux_5182 (.in({n13691_1, n13664_0, n13661_0, n13649_1, n13640_0, n13630_0, n13625_0/**/, n13586_0, n13571_0, n13560_0, n10268_1, n5657, n5649, n5561, n5553, n5545}), .out(n10348), .config_in(config_chain[16611:16606]), .config_rst(config_rst)); 
buffer_wire buffer_10348 (.in(n10348), .out(n10348_0));
mux4 mux_5183 (.in({n14729_1, n14620_0, n8595, n8479}), .out(n10349), .config_in(config_chain[16613:16612]), .config_rst(config_rst)); 
buffer_wire buffer_10349 (.in(n10349), .out(n10349_0));
mux16 mux_5184 (.in({n13673_1, n13658_0, n13655_0, n13651_1, n13642_0, n13627_0, n13622_0, n13616_0, n13601_0, n13562_0, n10270_1, n5657, n5649, n5561, n5553, n5545/**/}), .out(n10350), .config_in(config_chain[16619:16614]), .config_rst(config_rst)); 
buffer_wire buffer_10350 (.in(n10350), .out(n10350_0));
mux3 mux_5185 (.in({n14731_1, n14628_0, n8483}), .out(n10351), .config_in(config_chain[16621:16620]), .config_rst(config_rst)); 
buffer_wire buffer_10351 (.in(n10351), .out(n10351_0));
mux15 mux_5186 (.in({n13675_1, n13669_0, n13652_0, n13644_0, n13618_0, n13614_0, n13603_0, n13592_0/**/, n13577_0, n10272_1, n5657, n5649, n5561, n5553, n5545}), .out(n10352), .config_in(config_chain[16627:16622]), .config_rst(config_rst)); 
buffer_wire buffer_10352 (.in(n10352), .out(n10352_0));
mux3 mux_5187 (.in({n14733_1, n14636_0/**/, n8487}), .out(n10353), .config_in(config_chain[16629:16628]), .config_rst(config_rst)); 
buffer_wire buffer_10353 (.in(n10353), .out(n10353_0));
mux15 mux_5188 (.in({n13677_1, n13666_0, n13663_0, n13646_0, n13633_0, n13606_0, n13594_0, n13579_0, n13568_0, n10274_1, n5657, n5649/**/, n5561, n5553, n5545}), .out(n10354), .config_in(config_chain[16635:16630]), .config_rst(config_rst)); 
buffer_wire buffer_10354 (.in(n10354), .out(n10354_0));
mux3 mux_5189 (.in({n14735_1, n14644_0/**/, n8491}), .out(n10355), .config_in(config_chain[16637:16636]), .config_rst(config_rst)); 
buffer_wire buffer_10355 (.in(n10355), .out(n10355_0));
mux15 mux_5190 (.in({n13679_1, n13660_0, n13657_0, n13648_0, n13635_0, n13624_0, n13609_0, n13598_0, n13570_0/**/, n10276_1, n5657, n5649, n5561, n5553, n5545}), .out(n10356), .config_in(config_chain[16643:16638]), .config_rst(config_rst)); 
buffer_wire buffer_10356 (.in(n10356), .out(n10356_0));
mux3 mux_5191 (.in({n14737_1, n14652_0, n8491}), .out(n10357), .config_in(config_chain[16645:16644]), .config_rst(config_rst)); 
buffer_wire buffer_10357 (.in(n10357), .out(n10357_0));
mux15 mux_5192 (.in({n13681_1, n13671_0, n13654_0, n13650_0, n13626_0, n13611_0, n13600_0, n13590_0, n13585_0/**/, n10278_1, n5661, n5653, n5645, n5557, n5549}), .out(n10358), .config_in(config_chain[16651:16646]), .config_rst(config_rst)); 
buffer_wire buffer_10358 (.in(n10358), .out(n10358_0));
mux3 mux_5193 (.in({n14739_1, n14660_0/**/, n8495}), .out(n10359), .config_in(config_chain[16653:16652]), .config_rst(config_rst)); 
buffer_wire buffer_10359 (.in(n10359), .out(n10359_0));
mux15 mux_5194 (.in({n13683_1, n13668_0/**/, n13665_0, n13641_0, n13602_0, n13587_0, n13582_0, n13576_0, n13561_0, n10280_1, n5661, n5653, n5645, n5557, n5549}), .out(n10360), .config_in(config_chain[16659:16654]), .config_rst(config_rst)); 
buffer_wire buffer_10360 (.in(n10360), .out(n10360_0));
mux3 mux_5195 (.in({n14741_1, n14668_0, n8579/**/}), .out(n10361), .config_in(config_chain[16661:16660]), .config_rst(config_rst)); 
buffer_wire buffer_10361 (.in(n10361), .out(n10361_0));
mux15 mux_5196 (.in({n13685_1, n13662_0, n13659_0, n13643_0, n13632_0/**/, n13617_0, n13578_0, n13574_0, n13563_0, n10282_1, n5661, n5653, n5645, n5557, n5549}), .out(n10362), .config_in(config_chain[16667:16662]), .config_rst(config_rst)); 
buffer_wire buffer_10362 (.in(n10362), .out(n10362_0));
mux3 mux_5197 (.in({n14743_1, n14676_0/**/, n8583}), .out(n10363), .config_in(config_chain[16669:16668]), .config_rst(config_rst)); 
buffer_wire buffer_10363 (.in(n10363), .out(n10363_0));
mux15 mux_5198 (.in({n13687_1, n13656_0, n13653_0, n13645_0, n13634_0, n13619_0, n13608_0, n13593_0, n13566_0/**/, n10284_1, n5661, n5653, n5645, n5557, n5549}), .out(n10364), .config_in(config_chain[16675:16670]), .config_rst(config_rst)); 
buffer_wire buffer_10364 (.in(n10364), .out(n10364_0));
mux3 mux_5199 (.in({n14745_1, n14684_0, n8587}), .out(n10365), .config_in(config_chain[16677:16676]), .config_rst(config_rst)); 
buffer_wire buffer_10365 (.in(n10365), .out(n10365_0));
mux15 mux_5200 (.in({n13689_1, n13670_0, n13667_0, n13647_1, n13638_0, n13610_0, n13595_0, n13584_0, n13569_0, n10286_1/**/, n5661, n5653, n5645, n5557, n5549}), .out(n10366), .config_in(config_chain[16683:16678]), .config_rst(config_rst)); 
buffer_wire buffer_10366 (.in(n10366), .out(n10366_0));
mux3 mux_5201 (.in({n14747_1, n14692_0, n8587}), .out(n10367), .config_in(config_chain[16685:16684]), .config_rst(config_rst)); 
buffer_wire buffer_10367 (.in(n10367), .out(n10367_0));
mux15 mux_5202 (.in({n13957_2, n13929_0, n13922_0, n13912_0, n13909_0, n13896_0, n13884_0, n13851_0, n13826_0, n10288_1/**/, n6635, n6627, n6539, n6531, n6523}), .out(n10368), .config_in(config_chain[16691:16686]), .config_rst(config_rst)); 
buffer_wire buffer_10368 (.in(n10368), .out(n10368_0));
mux4 mux_5203 (.in({n14615_0, n14614_0, n8595, n8479}), .out(n10369), .config_in(config_chain[16693:16692]), .config_rst(config_rst)); 
buffer_wire buffer_10369 (.in(n10369), .out(n10369_0));
mux15 mux_5204 (.in({n13937_1, n13930_0, n13914_0, n13911_0, n13888_0, n13883_0/**/, n13858_0, n13853_0, n13828_0, n10290_1, n6639, n6627, n6539, n6531, n6523}), .out(n10370), .config_in(config_chain[16699:16694]), .config_rst(config_rst)); 
buffer_wire buffer_10370 (.in(n10370), .out(n10370_0));
mux3 mux_5205 (.in({n14623_0/**/, n14622_0, n8479}), .out(n10371), .config_in(config_chain[16701:16700]), .config_rst(config_rst)); 
buffer_wire buffer_10371 (.in(n10371), .out(n10371_0));
mux15 mux_5206 (.in({n13939_1/**/, n13923_0, n13916_0, n13913_1, n13890_0, n13885_0, n13880_0, n13860_0, n13827_0, n10292_1, n6639, n6631, n6539, n6531, n6523}), .out(n10372), .config_in(config_chain[16707:16702]), .config_rst(config_rst)); 
buffer_wire buffer_10372 (.in(n10372), .out(n10372_0));
mux3 mux_5207 (.in({n14631_0, n14630_0, n8483}), .out(n10373), .config_in(config_chain[16709:16708]), .config_rst(config_rst)); 
buffer_wire buffer_10373 (.in(n10373), .out(n10373_0));
mux15 mux_5208 (.in({n13941_1, n13931_0, n13924_0, n13915_1, n13892_0, n13872_0, n13859_0, n13834_0, n13829_0/**/, n10294_1, n6639, n6631, n6623, n6531, n6523}), .out(n10374), .config_in(config_chain[16715:16710]), .config_rst(config_rst)); 
buffer_wire buffer_10374 (.in(n10374), .out(n10374_0));
mux3 mux_5209 (.in({n14639_0, n14638_0/**/, n8487}), .out(n10375), .config_in(config_chain[16717:16716]), .config_rst(config_rst)); 
buffer_wire buffer_10375 (.in(n10375), .out(n10375_0));
mux14 mux_5210 (.in({n13943_1, n13932_0, n13917_0, n13891_0, n13866_0, n13864_0, n13861_0, n13836_0, n10296_1/**/, n6639, n6631, n6623, n6535, n6523}), .out(n10376), .config_in(config_chain[16723:16718]), .config_rst(config_rst)); 
buffer_wire buffer_10376 (.in(n10376), .out(n10376_0));
mux3 mux_5211 (.in({n14647_0, n14646_0, n8491}), .out(n10377), .config_in(config_chain[16725:16724]), .config_rst(config_rst)); 
buffer_wire buffer_10377 (.in(n10377), .out(n10377_0));
mux14 mux_5212 (.in({n13945_1, n13925_0, n13918_0, n13898_0, n13893_0, n13868_0, n13856_0, n13835_0, n10298_1/**/, n6639, n6631, n6623, n6535, n6527}), .out(n10378), .config_in(config_chain[16731:16726]), .config_rst(config_rst)); 
buffer_wire buffer_10378 (.in(n10378), .out(n10378_0));
mux3 mux_5213 (.in({n14655_0, n14654_0, n8495}), .out(n10379), .config_in(config_chain[16733:16732]), .config_rst(config_rst)); 
buffer_wire buffer_10379 (.in(n10379), .out(n10379_0));
mux13 mux_5214 (.in({n13947_1, n13933_0, n13926_0, n13900_0, n13867_0, n13848_0/**/, n13842_0, n13837_0, n10300_1, n6631, n6623, n6535, n6527}), .out(n10380), .config_in(config_chain[16739:16734]), .config_rst(config_rst)); 
buffer_wire buffer_10380 (.in(n10380), .out(n10380_0));
mux3 mux_5215 (.in({n14663_0, n14662_0, n8495}), .out(n10381), .config_in(config_chain[16741:16740]), .config_rst(config_rst)); 
buffer_wire buffer_10381 (.in(n10381), .out(n10381_0));
mux13 mux_5216 (.in({n13949_1, n13934_0, n13919_0, n13899_0, n13874_0, n13869_0/**/, n13844_0, n13840_0, n10302_1, n6635, n6623, n6535, n6527}), .out(n10382), .config_in(config_chain[16747:16742]), .config_rst(config_rst)); 
buffer_wire buffer_10382 (.in(n10382), .out(n10382_0));
mux3 mux_5217 (.in({n14671_0, n14670_0, n8579}), .out(n10383), .config_in(config_chain[16749:16748]), .config_rst(config_rst)); 
buffer_wire buffer_10383 (.in(n10383), .out(n10383_0));
mux13 mux_5218 (.in({n13951_1, n13927_0, n13920_0, n13906_0, n13901_0, n13876_0, n13843_0, n13832_0, n10304_1, n6635, n6627, n6535, n6527}), .out(n10384), .config_in(config_chain[16755:16750]), .config_rst(config_rst)); 
buffer_wire buffer_10384 (.in(n10384), .out(n10384_0));
mux3 mux_5219 (.in({n14679_0, n14678_0, n8583}), .out(n10385), .config_in(config_chain[16757:16756]), .config_rst(config_rst)); 
buffer_wire buffer_10385 (.in(n10385), .out(n10385_0));
mux13 mux_5220 (.in({n13953_1, n13935_0, n13928_0, n13908_0, n13875_0, n13850_0, n13845_0, n13824_0, n10306_1/**/, n6635, n6627, n6539, n6527}), .out(n10386), .config_in(config_chain[16763:16758]), .config_rst(config_rst)); 
buffer_wire buffer_10386 (.in(n10386), .out(n10386_0));
mux3 mux_5221 (.in({n14687_0, n14686_0, n8587}), .out(n10387), .config_in(config_chain[16765:16764]), .config_rst(config_rst)); 
buffer_wire buffer_10387 (.in(n10387), .out(n10387_0));
mux13 mux_5222 (.in({n13955_1, n13921_0, n13910_0, n13907_0/**/, n13904_0, n13882_0, n13877_0, n13852_0, n10256_1, n6635, n6627, n6539, n6531}), .out(n10388), .config_in(config_chain[16771:16766]), .config_rst(config_rst)); 
buffer_wire buffer_10388 (.in(n10388), .out(n10388_0));
mux3 mux_5223 (.in({n14695_2, n14694_0, n8591}), .out(n10389), .config_in(config_chain[16773:16772]), .config_rst(config_rst)); 
buffer_wire buffer_10389 (.in(n10389), .out(n10389_0));
mux15 mux_5224 (.in({n14223_2, n14187_0, n14180_0, n14176_0, n14173_0, n14162_0, n14148_0, n14143_0, n14118_0, n10308_1, n7613, n7605, n7517, n7509, n7501/**/}), .out(n10390), .config_in(config_chain[16779:16774]), .config_rst(config_rst)); 
buffer_wire buffer_10390 (.in(n10390), .out(n10390_0));
mux4 mux_5225 (.in({n14617_0/**/, n14616_0, n8595, n8479}), .out(n10391), .config_in(config_chain[16781:16780]), .config_rst(config_rst)); 
buffer_wire buffer_10391 (.in(n10391), .out(n10391_0));
mux15 mux_5226 (.in({n14203_1, n14195_0, n14188_0/**/, n14178_0, n14175_0, n14154_0, n14150_0, n14117_0, n14092_0, n10310_1, n7617, n7605, n7517, n7509, n7501}), .out(n10392), .config_in(config_chain[16787:16782]), .config_rst(config_rst)); 
buffer_wire buffer_10392 (.in(n10392), .out(n10392_0));
mux3 mux_5227 (.in({n14625_0, n14624_0, n8483}), .out(n10393), .config_in(config_chain[16789:16788]), .config_rst(config_rst)); 
buffer_wire buffer_10393 (.in(n10393), .out(n10393_0));
mux15 mux_5228 (.in({n14205_1, n14196_0, n14181_0, n14177_0, n14149_0, n14146_0, n14124_0, n14119_0, n14094_0, n10312_1, n7617, n7609, n7517, n7509, n7501/**/}), .out(n10394), .config_in(config_chain[16795:16790]), .config_rst(config_rst)); 
buffer_wire buffer_10394 (.in(n10394), .out(n10394_0));
mux3 mux_5229 (.in({n14633_0, n14632_0, n8483}), .out(n10395), .config_in(config_chain[16797:16796]), .config_rst(config_rst)); 
buffer_wire buffer_10395 (.in(n10395), .out(n10395_0));
mux15 mux_5230 (.in({n14207_1, n14189_0, n14182_0, n14179_1, n14156_0, n14151_0, n14138_0, n14126_0, n14093_0, n10314_1, n7617, n7609, n7601, n7509, n7501}), .out(n10396), .config_in(config_chain[16803:16798]), .config_rst(config_rst)); 
buffer_wire buffer_10396 (.in(n10396), .out(n10396_0));
mux3 mux_5231 (.in({n14641_0, n14640_0, n8487}), .out(n10397), .config_in(config_chain[16805:16804]), .config_rst(config_rst)); 
buffer_wire buffer_10397 (.in(n10397), .out(n10397_0));
mux14 mux_5232 (.in({n14209_1, n14197_0, n14190_0, n14158_0, n14130_0, n14125_0, n14100_0, n14095_0, n10316_1, n7617, n7609/**/, n7601, n7513, n7501}), .out(n10398), .config_in(config_chain[16811:16806]), .config_rst(config_rst)); 
buffer_wire buffer_10398 (.in(n10398), .out(n10398_0));
mux3 mux_5233 (.in({n14649_0, n14648_0, n8491}), .out(n10399), .config_in(config_chain[16813:16812]), .config_rst(config_rst)); 
buffer_wire buffer_10399 (.in(n10399), .out(n10399_0));
mux14 mux_5234 (.in({n14211_1, n14198_0, n14183_0, n14157_0, n14132_0, n14127_0, n14122_0, n14102_0, n10318_1, n7617, n7609/**/, n7601, n7513, n7505}), .out(n10400), .config_in(config_chain[16819:16814]), .config_rst(config_rst)); 
buffer_wire buffer_10400 (.in(n10400), .out(n10400_0));
mux3 mux_5235 (.in({n14657_0/**/, n14656_0, n8495}), .out(n10401), .config_in(config_chain[16821:16820]), .config_rst(config_rst)); 
buffer_wire buffer_10401 (.in(n10401), .out(n10401_0));
mux13 mux_5236 (.in({n14213_1, n14191_0, n14184_0, n14164_0, n14159_0, n14134_0, n14114_0, n14101_0, n10320_1, n7609, n7601/**/, n7513, n7505}), .out(n10402), .config_in(config_chain[16827:16822]), .config_rst(config_rst)); 
buffer_wire buffer_10402 (.in(n10402), .out(n10402_0));
mux3 mux_5237 (.in({n14665_0, n14664_0, n8579}), .out(n10403), .config_in(config_chain[16829:16828]), .config_rst(config_rst)); 
buffer_wire buffer_10403 (.in(n10403), .out(n10403_0));
mux13 mux_5238 (.in({n14215_1, n14199_0, n14192_0, n14166_0, n14133_0/**/, n14108_0, n14106_0, n14103_0, n10322_1, n7613, n7601, n7513, n7505}), .out(n10404), .config_in(config_chain[16835:16830]), .config_rst(config_rst)); 
buffer_wire buffer_10404 (.in(n10404), .out(n10404_0));
mux3 mux_5239 (.in({n14673_0, n14672_0, n8579}), .out(n10405), .config_in(config_chain[16837:16836]), .config_rst(config_rst)); 
buffer_wire buffer_10405 (.in(n10405), .out(n10405_0));
mux13 mux_5240 (.in({n14217_1, n14200_0, n14185_0, n14165_0, n14140_0, n14135_0, n14110_0, n14098_0, n10324_1/**/, n7613, n7605, n7513, n7505}), .out(n10406), .config_in(config_chain[16843:16838]), .config_rst(config_rst)); 
buffer_wire buffer_10406 (.in(n10406), .out(n10406_0));
mux3 mux_5241 (.in({n14681_0, n14680_0, n8583}), .out(n10407), .config_in(config_chain[16845:16844]), .config_rst(config_rst)); 
buffer_wire buffer_10407 (.in(n10407), .out(n10407_0));
mux13 mux_5242 (.in({n14219_1, n14193_0, n14186_0, n14172_0, n14167_0, n14142_0, n14109_0, n14090_0, n10326_1/**/, n7613, n7605, n7517, n7505}), .out(n10408), .config_in(config_chain[16851:16846]), .config_rst(config_rst)); 
buffer_wire buffer_10408 (.in(n10408), .out(n10408_0));
mux3 mux_5243 (.in({n14689_0, n14688_0, n8587}), .out(n10409), .config_in(config_chain[16853:16852]), .config_rst(config_rst)); 
buffer_wire buffer_10409 (.in(n10409), .out(n10409_0));
mux13 mux_5244 (.in({n14221_1, n14201_2, n14194_0, n14174_0, n14170_0, n14141_0, n14116_0, n14111_0, n10258_2, n7613, n7605, n7517, n7509}), .out(n10410), .config_in(config_chain[16859:16854]), .config_rst(config_rst)); 
buffer_wire buffer_10410 (.in(n10410), .out(n10410_0));
mux3 mux_5245 (.in({n14697_2, n14696_0, n8591}), .out(n10411), .config_in(config_chain[16861:16860]), .config_rst(config_rst)); 
buffer_wire buffer_10411 (.in(n10411), .out(n10411_0));
mux15 mux_5246 (.in({n14487_2, n14465_2, n14458_0, n14440_0, n14428_0, n14407_0, n14382_0, n14377_0, n14352_0, n10328_1, n8591, n8583/**/, n8495, n8487, n8479}), .out(n10412), .config_in(config_chain[16867:16862]), .config_rst(config_rst)); 
buffer_wire buffer_10412 (.in(n10412), .out(n10412_0));
mux4 mux_5247 (.in({n14707_0/**/, n14706_0, n8595, n8479}), .out(n10413), .config_in(config_chain[16869:16868]), .config_rst(config_rst)); 
buffer_wire buffer_10413 (.in(n10413), .out(n10413_0));
mux15 mux_5248 (.in({n14467_1, n14451_0, n14444_0, n14442_0, n14439_0, n14420_0, n14414_0, n14409_0, n14384_0/**/, n10330_1, n8595, n8583, n8495, n8487, n8479}), .out(n10414), .config_in(config_chain[16875:16870]), .config_rst(config_rst)); 
buffer_wire buffer_10414 (.in(n10414), .out(n10414_0));
mux3 mux_5249 (.in({n14709_0/**/, n14708_0, n8483}), .out(n10415), .config_in(config_chain[16877:16876]), .config_rst(config_rst)); 
buffer_wire buffer_10415 (.in(n10415), .out(n10415_0));
mux15 mux_5250 (.in({n14469_1, n14459_0, n14452_0, n14441_0, n14416_0, n14412_0, n14383_0, n14358_0, n14353_0, n10332_1, n8595, n8587, n8495, n8487, n8479}), .out(n10416), .config_in(config_chain[16883:16878]), .config_rst(config_rst)); 
buffer_wire buffer_10416 (.in(n10416), .out(n10416_0));
mux3 mux_5251 (.in({n14711_0/**/, n14710_0, n8487}), .out(n10417), .config_in(config_chain[16885:16884]), .config_rst(config_rst)); 
buffer_wire buffer_10417 (.in(n10417), .out(n10417_0));
mux15 mux_5252 (.in({n14471_1, n14460_0, n14445_0/**/, n14443_0, n14415_0, n14404_0, n14390_0, n14385_0, n14360_0, n10334_1, n8595, n8587, n8579, n8487, n8479}), .out(n10418), .config_in(config_chain[16891:16886]), .config_rst(config_rst)); 
buffer_wire buffer_10418 (.in(n10418), .out(n10418_0));
mux3 mux_5253 (.in({n14713_0/**/, n14712_0, n8487}), .out(n10419), .config_in(config_chain[16893:16892]), .config_rst(config_rst)); 
buffer_wire buffer_10419 (.in(n10419), .out(n10419_0));
mux14 mux_5254 (.in({n14473_1, n14453_0, n14446_0, n14422_0, n14417_0, n14396_0, n14392_0/**/, n14359_0, n10336_1, n8595, n8587, n8579, n8491, n8479}), .out(n10420), .config_in(config_chain[16899:16894]), .config_rst(config_rst)); 
buffer_wire buffer_10420 (.in(n10420), .out(n10420_0));
mux3 mux_5255 (.in({n14715_0, n14714_0, n8491}), .out(n10421), .config_in(config_chain[16901:16900]), .config_rst(config_rst)); 
buffer_wire buffer_10421 (.in(n10421), .out(n10421_0));
mux14 mux_5256 (.in({n14475_1, n14461_0, n14454_0, n14424_0/**/, n14391_0, n14388_0, n14366_0, n14361_0, n10338_1, n8595, n8587, n8579, n8491, n8483}), .out(n10422), .config_in(config_chain[16907:16902]), .config_rst(config_rst)); 
buffer_wire buffer_10422 (.in(n10422), .out(n10422_0));
mux3 mux_5257 (.in({n14717_0, n14716_0, n8495}), .out(n10423), .config_in(config_chain[16909:16908]), .config_rst(config_rst)); 
buffer_wire buffer_10423 (.in(n10423), .out(n10423_0));
mux13 mux_5258 (.in({n14477_1, n14462_0, n14447_0, n14423_0, n14398_0, n14393_0, n14380_0, n14368_0, n10340_1, n8587/**/, n8579, n8491, n8483}), .out(n10424), .config_in(config_chain[16915:16910]), .config_rst(config_rst)); 
buffer_wire buffer_10424 (.in(n10424), .out(n10424_0));
mux3 mux_5259 (.in({n14719_0, n14718_0, n8579/**/}), .out(n10425), .config_in(config_chain[16917:16916]), .config_rst(config_rst)); 
buffer_wire buffer_10425 (.in(n10425), .out(n10425_0));
mux13 mux_5260 (.in({n14479_1, n14455_0, n14448_0, n14430_0, n14425_0, n14400_0, n14372_0, n14367_0, n10342_1/**/, n8591, n8579, n8491, n8483}), .out(n10426), .config_in(config_chain[16923:16918]), .config_rst(config_rst)); 
buffer_wire buffer_10426 (.in(n10426), .out(n10426_0));
mux3 mux_5261 (.in({n14721_0, n14720_0, n8583}), .out(n10427), .config_in(config_chain[16925:16924]), .config_rst(config_rst)); 
buffer_wire buffer_10427 (.in(n10427), .out(n10427_0));
mux13 mux_5262 (.in({n14481_1, n14463_0, n14456_0, n14432_0, n14399_0/**/, n14374_0, n14369_0, n14364_0, n10344_1, n8591, n8583, n8491, n8483}), .out(n10428), .config_in(config_chain[16931:16926]), .config_rst(config_rst)); 
buffer_wire buffer_10428 (.in(n10428), .out(n10428_0));
mux3 mux_5263 (.in({n14723_0/**/, n14722_0, n8583}), .out(n10429), .config_in(config_chain[16933:16932]), .config_rst(config_rst)); 
buffer_wire buffer_10429 (.in(n10429), .out(n10429_0));
mux13 mux_5264 (.in({n14483_1, n14464_0, n14449_0, n14431_0, n14406_0, n14401_0, n14376_0, n14356_0, n10346_1, n8591, n8583, n8495, n8483}), .out(n10430), .config_in(config_chain[16939:16934]), .config_rst(config_rst)); 
buffer_wire buffer_10430 (.in(n10430), .out(n10430_0));
mux3 mux_5265 (.in({n14725_0/**/, n14724_0, n8587}), .out(n10431), .config_in(config_chain[16941:16940]), .config_rst(config_rst)); 
buffer_wire buffer_10431 (.in(n10431), .out(n10431_0));
mux13 mux_5266 (.in({n14485_1, n14457_0, n14450_0/**/, n14438_0, n14436_0, n14433_2, n14408_0, n14375_0, n10260_2, n8591, n8583, n8495, n8487}), .out(n10432), .config_in(config_chain[16947:16942]), .config_rst(config_rst)); 
buffer_wire buffer_10432 (.in(n10432), .out(n10432_0));
mux3 mux_5267 (.in({n14727_2, n14726_0, n8591}), .out(n10433), .config_in(config_chain[16949:16948]), .config_rst(config_rst)); 
buffer_wire buffer_10433 (.in(n10433), .out(n10433_0));
mux4 mux_5268 (.in({n12271_0, n12270_0, n869, n753/**/}), .out(n10434), .config_in(config_chain[16951:16950]), .config_rst(config_rst)); 
buffer_wire buffer_10434 (.in(n10434), .out(n10434_0));
mux16 mux_5269 (.in({n12657_1, n12649_0, n12644_0, n12623_0, n12618_0, n12612_0, n12605_1, n12596_0, n12590_0, n12527_0, n10527_1, n865/**/, n857, n769, n761, n753}), .out(n10435), .config_in(config_chain[16957:16952]), .config_rst(config_rst)); 
buffer_wire buffer_10435 (.in(n10435), .out(n10435_0));
mux4 mux_5270 (.in({n12363_0/**/, n12362_0, n869, n753}), .out(n10436), .config_in(config_chain[16959:16958]), .config_rst(config_rst)); 
buffer_wire buffer_10436 (.in(n10436), .out(n10436_0));
mux16 mux_5271 (.in({n12913_1, n12908_0, n12893_0, n12885_0, n12880_0, n12868_0, n12861_0, n12854_0, n12809_0, n12792_0, n10547_1, n1843, n1835, n1747, n1739/**/, n1731}), .out(n10437), .config_in(config_chain[16965:16960]), .config_rst(config_rst)); 
buffer_wire buffer_10437 (.in(n10437), .out(n10437_0));
mux4 mux_5272 (.in({n12383_0/**/, n12382_0, n869, n753}), .out(n10438), .config_in(config_chain[16967:16966]), .config_rst(config_rst)); 
buffer_wire buffer_10438 (.in(n10438), .out(n10438_0));
mux16 mux_5273 (.in({n13171_1, n13157_0, n13152_0, n13146_0, n13131_0, n13126_0, n13119_0, n13114_0, n13093_0, n13076_0, n10567_1, n2821, n2813, n2725, n2717, n2709}), .out(n10439), .config_in(config_chain[16973:16968]), .config_rst(config_rst)); 
buffer_wire buffer_10439 (.in(n10439), .out(n10439_0));
mux4 mux_5274 (.in({n12403_1, n12276_0, n869, n753}), .out(n10440), .config_in(config_chain[16975:16974]), .config_rst(config_rst)); 
buffer_wire buffer_10440 (.in(n10440), .out(n10440_0));
mux16 mux_5275 (.in({n13431_1, n13423_0, n13418_0, n13397_0, n13392_0, n13386_0, n13379_0, n13376_0, n13362_0, n13299_0, n10587_1, n3799, n3791/**/, n3703, n3695, n3687}), .out(n10441), .config_in(config_chain[16981:16976]), .config_rst(config_rst)); 
buffer_wire buffer_10441 (.in(n10441), .out(n10441_0));
mux3 mux_5276 (.in({n12279_0, n12278_0, n753}), .out(n10442), .config_in(config_chain[16983:16982]), .config_rst(config_rst)); 
buffer_wire buffer_10442 (.in(n10442), .out(n10442_0));
mux16 mux_5277 (.in({n12675_1, n12643_0, n12638_0, n12632_0, n12617_0, n12614_0, n12607_1, n12583_0, n12566_0, n12524_0, n10529_1, n865, n857/**/, n769, n761, n753}), .out(n10443), .config_in(config_chain[16989:16984]), .config_rst(config_rst)); 
buffer_wire buffer_10443 (.in(n10443), .out(n10443_0));
mux3 mux_5278 (.in({n12365_0/**/, n12364_0, n757}), .out(n10444), .config_in(config_chain[16991:16990]), .config_rst(config_rst)); 
buffer_wire buffer_10444 (.in(n10444), .out(n10444_0));
mux16 mux_5279 (.in({n12931_1, n12907_0, n12902_0, n12879_0, n12874_0, n12870_0, n12863_1, n12848_0, n12785_0, n12782_0/**/, n10549_1, n1843, n1835, n1747, n1739, n1731}), .out(n10445), .config_in(config_chain[16997:16992]), .config_rst(config_rst)); 
buffer_wire buffer_10445 (.in(n10445), .out(n10445_0));
mux3 mux_5280 (.in({n12385_0, n12384_0, n757/**/}), .out(n10446), .config_in(config_chain[16999:16998]), .config_rst(config_rst)); 
buffer_wire buffer_10446 (.in(n10446), .out(n10446_0));
mux16 mux_5281 (.in({n13189_1, n13166_0, n13151_0, n13145_0, n13140_0, n13128_0, n13121_0, n13069_0, n13052_0, n13042_0, n10569_1, n2821/**/, n2813, n2725, n2717, n2709}), .out(n10447), .config_in(config_chain[17005:17000]), .config_rst(config_rst)); 
buffer_wire buffer_10447 (.in(n10447), .out(n10447_0));
mux3 mux_5282 (.in({n12405_1, n12284_0, n757}), .out(n10448), .config_in(config_chain[17007:17006]), .config_rst(config_rst)); 
buffer_wire buffer_10448 (.in(n10448), .out(n10448_0));
mux16 mux_5283 (.in({n13449_1, n13417_0, n13412_0, n13406_0, n13391_0, n13388_0, n13381_0, n13355_0, n13338_0, n13304_0, n10589_1, n3799, n3791, n3703, n3695, n3687/**/}), .out(n10449), .config_in(config_chain[17013:17008]), .config_rst(config_rst)); 
buffer_wire buffer_10449 (.in(n10449), .out(n10449_0));
mux3 mux_5284 (.in({n12287_0, n12286_0, n757/**/}), .out(n10450), .config_in(config_chain[17015:17014]), .config_rst(config_rst)); 
buffer_wire buffer_10450 (.in(n10450), .out(n10450_0));
mux15 mux_5285 (.in({n12673_1/**/, n12652_0, n12637_0, n12631_0, n12626_0, n12609_1, n12559_0, n12542_0, n12532_0, n10531_1, n865, n857, n769, n761, n753}), .out(n10451), .config_in(config_chain[17021:17016]), .config_rst(config_rst)); 
buffer_wire buffer_10451 (.in(n10451), .out(n10451_0));
mux3 mux_5286 (.in({n12367_0/**/, n12366_0, n757}), .out(n10452), .config_in(config_chain[17023:17022]), .config_rst(config_rst)); 
buffer_wire buffer_10452 (.in(n10452), .out(n10452_0));
mux15 mux_5287 (.in({n12929_1, n12901_0, n12896_0, n12888_0, n12873_0, n12865_1, n12841_0, n12824_0, n12790_0, n10551_1/**/, n1843, n1835, n1747, n1739, n1731}), .out(n10453), .config_in(config_chain[17029:17024]), .config_rst(config_rst)); 
buffer_wire buffer_10453 (.in(n10453), .out(n10453_0));
mux3 mux_5288 (.in({n12387_0/**/, n12386_0, n761}), .out(n10454), .config_in(config_chain[17031:17030]), .config_rst(config_rst)); 
buffer_wire buffer_10454 (.in(n10454), .out(n10454_0));
mux15 mux_5289 (.in({n13187_1, n13165_0, n13160_0, n13139_0, n13134_0, n13123_1, n13108_0, n13050_0, n13045_0, n10571_1, n2821, n2813, n2725, n2717, n2709}), .out(n10455), .config_in(config_chain[17037:17032]), .config_rst(config_rst)); 
buffer_wire buffer_10455 (.in(n10455), .out(n10455_0));
mux3 mux_5290 (.in({n12407_1, n12292_0, n761/**/}), .out(n10456), .config_in(config_chain[17039:17038]), .config_rst(config_rst)); 
buffer_wire buffer_10456 (.in(n10456), .out(n10456_0));
mux15 mux_5291 (.in({n13447_1, n13426_0, n13411_0, n13405_0/**/, n13400_0, n13383_0, n13331_0, n13314_0, n13312_0, n10591_1, n3799, n3791, n3703, n3695, n3687}), .out(n10457), .config_in(config_chain[17045:17040]), .config_rst(config_rst)); 
buffer_wire buffer_10457 (.in(n10457), .out(n10457_0));
mux3 mux_5292 (.in({n12295_0/**/, n12294_0, n761}), .out(n10458), .config_in(config_chain[17047:17046]), .config_rst(config_rst)); 
buffer_wire buffer_10458 (.in(n10458), .out(n10458_0));
mux15 mux_5293 (.in({n12671_1, n12651_0, n12646_0, n12625_0, n12620_0, n12611_1, n12598_0, n12540_0, n12535_0, n10533_1, n865/**/, n857, n769, n761, n753}), .out(n10459), .config_in(config_chain[17053:17048]), .config_rst(config_rst)); 
buffer_wire buffer_10459 (.in(n10459), .out(n10459_0));
mux3 mux_5294 (.in({n12369_0/**/, n12368_0, n761}), .out(n10460), .config_in(config_chain[17055:17054]), .config_rst(config_rst)); 
buffer_wire buffer_10460 (.in(n10460), .out(n10460_0));
mux15 mux_5295 (.in({n12927_1, n12910_0, n12895_0, n12887_0, n12882_0, n12867_1, n12817_0, n12800_0, n12798_0, n10553_1, n1843, n1835, n1747, n1739, n1731}), .out(n10461), .config_in(config_chain[17061:17056]), .config_rst(config_rst)); 
buffer_wire buffer_10461 (.in(n10461), .out(n10461_0));
mux3 mux_5296 (.in({n12389_0, n12388_0, n761/**/}), .out(n10462), .config_in(config_chain[17063:17062]), .config_rst(config_rst)); 
buffer_wire buffer_10462 (.in(n10462), .out(n10462_0));
mux15 mux_5297 (.in({n13185_1, n13159_0, n13154_0, n13148_0/**/, n13133_0, n13125_1, n13101_0, n13084_0, n13058_0, n10573_1, n2821, n2813, n2725, n2717, n2709}), .out(n10463), .config_in(config_chain[17069:17064]), .config_rst(config_rst)); 
buffer_wire buffer_10463 (.in(n10463), .out(n10463_0));
mux3 mux_5298 (.in({n12409_1, n12300_0, n765}), .out(n10464), .config_in(config_chain[17071:17070]), .config_rst(config_rst)); 
buffer_wire buffer_10464 (.in(n10464), .out(n10464_0));
mux15 mux_5299 (.in({n13445_1, n13425_0, n13420_0, n13399_0, n13394_0, n13385_1, n13370_0, n13320_0, n13307_0, n10593_1, n3799, n3791/**/, n3703, n3695, n3687}), .out(n10465), .config_in(config_chain[17077:17072]), .config_rst(config_rst)); 
buffer_wire buffer_10465 (.in(n10465), .out(n10465_0));
mux3 mux_5300 (.in({n12303_0/**/, n12302_0, n765}), .out(n10466), .config_in(config_chain[17079:17078]), .config_rst(config_rst)); 
buffer_wire buffer_10466 (.in(n10466), .out(n10466_0));
mux15 mux_5301 (.in({n12669_1, n12645_0, n12640_0, n12634_0, n12619_0, n12613_1, n12591_0, n12574_0, n12548_0, n10535_1, n865, n857, n769, n761/**/, n753}), .out(n10467), .config_in(config_chain[17085:17080]), .config_rst(config_rst)); 
buffer_wire buffer_10467 (.in(n10467), .out(n10467_0));
mux3 mux_5302 (.in({n12371_0, n12370_0, n765}), .out(n10468), .config_in(config_chain[17087:17086]), .config_rst(config_rst)); 
buffer_wire buffer_10468 (.in(n10468), .out(n10468_0));
mux15 mux_5303 (.in({n12925_1, n12909_0, n12904_0, n12881_0, n12876_0, n12869_1, n12856_0, n12806_0, n12793_0, n10555_1, n1843, n1835, n1747, n1739, n1731}), .out(n10469), .config_in(config_chain[17093:17088]), .config_rst(config_rst)); 
buffer_wire buffer_10469 (.in(n10469), .out(n10469_0));
mux3 mux_5304 (.in({n12391_0, n12390_0, n765}), .out(n10470), .config_in(config_chain[17095:17094]), .config_rst(config_rst)); 
buffer_wire buffer_10470 (.in(n10470), .out(n10470_0));
mux15 mux_5305 (.in({n13183_1, n13168_0, n13153_0, n13147_0, n13142_0, n13127_1, n13077_0, n13066_0, n13060_0, n10575_1/**/, n2821, n2813, n2725, n2717, n2709}), .out(n10471), .config_in(config_chain[17101:17096]), .config_rst(config_rst)); 
buffer_wire buffer_10471 (.in(n10471), .out(n10471_0));
mux3 mux_5306 (.in({n12411_1, n12308_0, n765}), .out(n10472), .config_in(config_chain[17103:17102]), .config_rst(config_rst)); 
buffer_wire buffer_10472 (.in(n10472), .out(n10472_0));
mux15 mux_5307 (.in({n13443_1, n13419_0, n13414_0, n13408_0, n13393_0, n13387_1, n13363_0, n13346_0, n13328_0, n10595_1, n3799, n3791, n3703, n3695, n3687/**/}), .out(n10473), .config_in(config_chain[17109:17104]), .config_rst(config_rst)); 
buffer_wire buffer_10473 (.in(n10473), .out(n10473_0));
mux3 mux_5308 (.in({n12311_0, n12310_0, n769}), .out(n10474), .config_in(config_chain[17111:17110]), .config_rst(config_rst)); 
buffer_wire buffer_10474 (.in(n10474), .out(n10474_0));
mux15 mux_5309 (.in({n12667_1, n12654_0, n12639_0, n12633_0, n12628_0, n12615_1, n12567_0, n12556_0, n12550_0, n10537_1, n869, n861, n853, n765, n757}), .out(n10475), .config_in(config_chain[17117:17112]), .config_rst(config_rst)); 
buffer_wire buffer_10475 (.in(n10475), .out(n10475_0));
mux3 mux_5310 (.in({n12373_0, n12372_0, n769}), .out(n10476), .config_in(config_chain[17119:17118]), .config_rst(config_rst)); 
buffer_wire buffer_10476 (.in(n10476), .out(n10476_0));
mux15 mux_5311 (.in({n12923_1, n12903_0, n12898_0, n12890_0, n12875_0/**/, n12871_1, n12849_0, n12832_0, n12814_0, n10557_1, n1847, n1839, n1831, n1743, n1735}), .out(n10477), .config_in(config_chain[17125:17120]), .config_rst(config_rst)); 
buffer_wire buffer_10477 (.in(n10477), .out(n10477_0));
mux3 mux_5312 (.in({n12393_0, n12392_0, n769}), .out(n10478), .config_in(config_chain[17127:17126]), .config_rst(config_rst)); 
buffer_wire buffer_10478 (.in(n10478), .out(n10478_0));
mux15 mux_5313 (.in({n13181_1, n13167_0, n13162_0, n13141_0, n13136_0, n13129_1, n13116_0, n13074_0, n13053_0, n10577_1, n2825, n2817, n2809, n2721, n2713}), .out(n10479), .config_in(config_chain[17133:17128]), .config_rst(config_rst)); 
buffer_wire buffer_10479 (.in(n10479), .out(n10479_0));
mux3 mux_5314 (.in({n12413_1, n12316_0, n769}), .out(n10480), .config_in(config_chain[17135:17134]), .config_rst(config_rst)); 
buffer_wire buffer_10480 (.in(n10480), .out(n10480_0));
mux15 mux_5315 (.in({n13441_1, n13428_0, n13413_0, n13407_0, n13402_0, n13389_1, n13339_0, n13336_0, n13322_0, n10597_1, n3803, n3795, n3787/**/, n3699, n3691}), .out(n10481), .config_in(config_chain[17141:17136]), .config_rst(config_rst)); 
buffer_wire buffer_10481 (.in(n10481), .out(n10481_0));
mux3 mux_5316 (.in({n12319_0, n12318_0, n769}), .out(n10482), .config_in(config_chain[17143:17142]), .config_rst(config_rst)); 
buffer_wire buffer_10482 (.in(n10482), .out(n10482_0));
mux15 mux_5317 (.in({n12665_1, n12653_0/**/, n12648_0, n12627_0, n12622_0, n12604_0, n12564_0, n12543_0, n12526_0, n10539_1, n869, n861, n853, n765, n757}), .out(n10483), .config_in(config_chain[17149:17144]), .config_rst(config_rst)); 
buffer_wire buffer_10483 (.in(n10483), .out(n10483_0));
mux3 mux_5318 (.in({n12375_0/**/, n12374_0, n853}), .out(n10484), .config_in(config_chain[17151:17150]), .config_rst(config_rst)); 
buffer_wire buffer_10484 (.in(n10484), .out(n10484_0));
mux15 mux_5319 (.in({n12921_1, n12897_0, n12892_0, n12889_0, n12884_0, n12860_0, n12825_0, n12822_0, n12808_0, n10559_1, n1847, n1839, n1831, n1743, n1735}), .out(n10485), .config_in(config_chain[17157:17152]), .config_rst(config_rst)); 
buffer_wire buffer_10485 (.in(n10485), .out(n10485_0));
mux3 mux_5320 (.in({n12395_0, n12394_0, n853}), .out(n10486), .config_in(config_chain[17159:17158]), .config_rst(config_rst)); 
buffer_wire buffer_10486 (.in(n10486), .out(n10486_0));
mux15 mux_5321 (.in({n13179_1, n13161_0, n13156_0, n13135_0, n13130_0/**/, n13118_0, n13109_0, n13092_0, n13082_0, n10579_1, n2825, n2817, n2809, n2721, n2713}), .out(n10487), .config_in(config_chain[17165:17160]), .config_rst(config_rst)); 
buffer_wire buffer_10487 (.in(n10487), .out(n10487_0));
mux3 mux_5322 (.in({n12415_1, n12324_0/**/, n853}), .out(n10488), .config_in(config_chain[17167:17166]), .config_rst(config_rst)); 
buffer_wire buffer_10488 (.in(n10488), .out(n10488_0));
mux15 mux_5323 (.in({n13439_1, n13427_0, n13422_0, n13401_0, n13396_0/**/, n13378_0, n13344_0, n13315_0, n13298_0, n10599_1, n3803, n3795, n3787, n3699, n3691}), .out(n10489), .config_in(config_chain[17173:17168]), .config_rst(config_rst)); 
buffer_wire buffer_10489 (.in(n10489), .out(n10489_0));
mux3 mux_5324 (.in({n12327_0/**/, n12326_0, n853}), .out(n10490), .config_in(config_chain[17175:17174]), .config_rst(config_rst)); 
buffer_wire buffer_10490 (.in(n10490), .out(n10490_0));
mux15 mux_5325 (.in({n12663_1, n12647_0, n12642_0, n12621_0, n12616_0, n12606_0, n12599_0, n12582_0, n12572_0, n10541_1, n869, n861, n853, n765, n757}), .out(n10491), .config_in(config_chain[17181:17176]), .config_rst(config_rst)); 
buffer_wire buffer_10491 (.in(n10491), .out(n10491_0));
mux3 mux_5326 (.in({n12377_0, n12376_0, n853}), .out(n10492), .config_in(config_chain[17183:17182]), .config_rst(config_rst)); 
buffer_wire buffer_10492 (.in(n10492), .out(n10492_0));
mux15 mux_5327 (.in({n12919_1, n12911_0, n12906_0, n12883_0, n12878_0/**/, n12862_0, n12830_0, n12801_0, n12784_0, n10561_1, n1847, n1839, n1831, n1743, n1735}), .out(n10493), .config_in(config_chain[17189:17184]), .config_rst(config_rst)); 
buffer_wire buffer_10493 (.in(n10493), .out(n10493_0));
mux3 mux_5328 (.in({n12397_0, n12396_0, n857}), .out(n10494), .config_in(config_chain[17191:17190]), .config_rst(config_rst)); 
buffer_wire buffer_10494 (.in(n10494), .out(n10494_0));
mux15 mux_5329 (.in({n13177_1, n13155_0, n13150_0, n13149_0, n13144_0/**/, n13120_0, n13090_0, n13085_0, n13068_0, n10581_1, n2825, n2817, n2809, n2721, n2713}), .out(n10495), .config_in(config_chain[17197:17192]), .config_rst(config_rst)); 
buffer_wire buffer_10495 (.in(n10495), .out(n10495_0));
mux3 mux_5330 (.in({n12417_1, n12332_0, n857}), .out(n10496), .config_in(config_chain[17199:17198]), .config_rst(config_rst)); 
buffer_wire buffer_10496 (.in(n10496), .out(n10496_0));
mux15 mux_5331 (.in({n13437_1, n13421_0, n13416_0, n13395_0, n13390_0, n13380_0, n13371_0, n13354_0, n13352_0, n10601_1, n3803, n3795, n3787/**/, n3699, n3691}), .out(n10497), .config_in(config_chain[17205:17200]), .config_rst(config_rst)); 
buffer_wire buffer_10497 (.in(n10497), .out(n10497_0));
mux3 mux_5332 (.in({n12335_0, n12334_0, n857}), .out(n10498), .config_in(config_chain[17207:17206]), .config_rst(config_rst)); 
buffer_wire buffer_10498 (.in(n10498), .out(n10498_0));
mux15 mux_5333 (.in({n12661_1, n12641_0, n12636_0, n12635_0, n12630_0, n12608_0, n12580_0, n12575_0, n12558_0, n10543_1, n869, n861, n853, n765, n757/**/}), .out(n10499), .config_in(config_chain[17213:17208]), .config_rst(config_rst)); 
buffer_wire buffer_10499 (.in(n10499), .out(n10499_0));
mux3 mux_5334 (.in({n12379_0/**/, n12378_0, n857}), .out(n10500), .config_in(config_chain[17215:17214]), .config_rst(config_rst)); 
buffer_wire buffer_10500 (.in(n10500), .out(n10500_0));
mux15 mux_5335 (.in({n12917_1, n12905_0, n12900_0, n12877_0, n12872_0/**/, n12864_0, n12857_0, n12840_0, n12838_0, n10563_1, n1847, n1839, n1831, n1743, n1735}), .out(n10501), .config_in(config_chain[17221:17216]), .config_rst(config_rst)); 
buffer_wire buffer_10501 (.in(n10501), .out(n10501_0));
mux3 mux_5336 (.in({n12399_0/**/, n12398_0, n857}), .out(n10502), .config_in(config_chain[17223:17222]), .config_rst(config_rst)); 
buffer_wire buffer_10502 (.in(n10502), .out(n10502_0));
mux15 mux_5337 (.in({n13175_1, n13169_0, n13164_0, n13143_0, n13138_0, n13122_0, n13098_0, n13061_0, n13044_0, n10583_1, n2825/**/, n2817, n2809, n2721, n2713}), .out(n10503), .config_in(config_chain[17229:17224]), .config_rst(config_rst)); 
buffer_wire buffer_10503 (.in(n10503), .out(n10503_0));
mux3 mux_5338 (.in({n12419_1/**/, n12340_0, n861}), .out(n10504), .config_in(config_chain[17231:17230]), .config_rst(config_rst)); 
buffer_wire buffer_10504 (.in(n10504), .out(n10504_0));
mux15 mux_5339 (.in({n13435_1, n13415_0, n13410_0, n13409_0, n13404_0, n13382_0, n13360_0, n13347_0, n13330_0, n10603_1, n3803, n3795, n3787, n3699, n3691}), .out(n10505), .config_in(config_chain[17237:17232]), .config_rst(config_rst)); 
buffer_wire buffer_10505 (.in(n10505), .out(n10505_0));
mux3 mux_5340 (.in({n12343_0, n12342_0, n861}), .out(n10506), .config_in(config_chain[17239:17238]), .config_rst(config_rst)); 
buffer_wire buffer_10506 (.in(n10506), .out(n10506_0));
mux15 mux_5341 (.in({n12659_1, n12655_0, n12650_0, n12629_0, n12624_0, n12610_0, n12588_0, n12551_0, n12534_0, n10545_1, n869, n861, n853, n765, n757}), .out(n10507), .config_in(config_chain[17245:17240]), .config_rst(config_rst)); 
buffer_wire buffer_10507 (.in(n10507), .out(n10507_0));
mux3 mux_5342 (.in({n12381_0/**/, n12380_0, n861}), .out(n10508), .config_in(config_chain[17247:17246]), .config_rst(config_rst)); 
buffer_wire buffer_10508 (.in(n10508), .out(n10508_0));
mux15 mux_5343 (.in({n12915_1, n12899_0/**/, n12894_0, n12891_0, n12886_0, n12866_0, n12846_0, n12833_0, n12816_0, n10565_1, n1847, n1839, n1831, n1743, n1735}), .out(n10509), .config_in(config_chain[17253:17248]), .config_rst(config_rst)); 
buffer_wire buffer_10509 (.in(n10509), .out(n10509_0));
mux3 mux_5344 (.in({n12401_0, n12400_0, n861}), .out(n10510), .config_in(config_chain[17255:17254]), .config_rst(config_rst)); 
buffer_wire buffer_10510 (.in(n10510), .out(n10510_0));
mux15 mux_5345 (.in({n13173_1, n13163_0, n13158_0, n13137_0, n13132_0, n13124_0, n13117_0/**/, n13106_0, n13100_0, n10585_1, n2825, n2817, n2809, n2721, n2713}), .out(n10511), .config_in(config_chain[17261:17256]), .config_rst(config_rst)); 
buffer_wire buffer_10511 (.in(n10511), .out(n10511_0));
mux3 mux_5346 (.in({n12421_1, n12348_0, n861}), .out(n10512), .config_in(config_chain[17263:17262]), .config_rst(config_rst)); 
buffer_wire buffer_10512 (.in(n10512), .out(n10512_0));
mux15 mux_5347 (.in({n13433_1, n13429_0, n13424_0, n13403_0, n13398_0, n13384_0, n13368_0, n13323_0, n13306_0, n10605_1, n3803/**/, n3795, n3787, n3699, n3691}), .out(n10513), .config_in(config_chain[17269:17264]), .config_rst(config_rst)); 
buffer_wire buffer_10513 (.in(n10513), .out(n10513_0));
mux3 mux_5348 (.in({n12351_1, n12350_0, n865}), .out(n10514), .config_in(config_chain[17271:17270]), .config_rst(config_rst)); 
buffer_wire buffer_10514 (.in(n10514), .out(n10514_0));
mux13 mux_5349 (.in({n13695_1, n13676_0, n13664_0, n13659_0, n13647_0, n13642_0, n13632_0/**/, n13619_0, n10627_1, n4777, n4769, n4681, n4673}), .out(n10515), .config_in(config_chain[17277:17272]), .config_rst(config_rst)); 
buffer_wire buffer_10515 (.in(n10515), .out(n10515_0));
mux3 mux_5350 (.in({n12353_1, n12352_0, n865}), .out(n10516), .config_in(config_chain[17279:17278]), .config_rst(config_rst)); 
buffer_wire buffer_10516 (.in(n10516), .out(n10516_0));
mux13 mux_5351 (.in({n13961_1, n13956_0, n13951_0, n13920_0, n13911_0/**/, n13898_0, n13876_0, n13853_0, n10649_0, n5755, n5747, n5659, n5651}), .out(n10517), .config_in(config_chain[17285:17280]), .config_rst(config_rst)); 
buffer_wire buffer_10517 (.in(n10517), .out(n10517_0));
mux3 mux_5352 (.in({n12355_1, n12354_0, n865}), .out(n10518), .config_in(config_chain[17287:17286]), .config_rst(config_rst)); 
buffer_wire buffer_10518 (.in(n10518), .out(n10518_0));
mux13 mux_5353 (.in({n14227_1, n14214_0, n14209_0, n14200_0/**/, n14195_0, n14175_0, n14164_0, n14110_0, n10671_0, n6733, n6725, n6637, n6629}), .out(n10519), .config_in(config_chain[17293:17288]), .config_rst(config_rst)); 
buffer_wire buffer_10519 (.in(n10519), .out(n10519_0));
mux3 mux_5354 (.in({n12357_1, n12356_0, n865}), .out(n10520), .config_in(config_chain[17295:17294]), .config_rst(config_rst)); 
buffer_wire buffer_10520 (.in(n10520), .out(n10520_0));
mux13 mux_5355 (.in({n14491_1, n14487_1, n14470_0, n14456_0/**/, n14451_0, n14432_0, n14430_0, n14409_0, n10693_0, n7711, n7703, n7615, n7607}), .out(n10521), .config_in(config_chain[17301:17296]), .config_rst(config_rst)); 
buffer_wire buffer_10521 (.in(n10521), .out(n10521_0));
mux3 mux_5356 (.in({n12359_1, n12358_0, n865}), .out(n10522), .config_in(config_chain[17303:17302]), .config_rst(config_rst)); 
buffer_wire buffer_10522 (.in(n10522), .out(n10522_0));
mux3 mux_5357 (.in({n14771_1, n14702_0, n8689}), .out(n10523), .config_in(config_chain[17305:17304]), .config_rst(config_rst)); 
buffer_wire buffer_10523 (.in(n10523), .out(n10523_0));
mux3 mux_5358 (.in({n12361_1, n12360_0, n869}), .out(n10524), .config_in(config_chain[17307:17306]), .config_rst(config_rst)); 
buffer_wire buffer_10524 (.in(n10524), .out(n10524_0));
mux3 mux_5359 (.in({n14705_0/**/, n14704_0, n8693}), .out(n10525), .config_in(config_chain[17309:17308]), .config_rst(config_rst)); 
buffer_wire buffer_10525 (.in(n10525), .out(n10525_0));
mux16 mux_5360 (.in({n12675_1, n12648_0, n12645_0/**/, n12622_0, n12619_0, n12613_1, n12604_0, n12591_0, n12588_0, n12526_0, n10434_0, n1843, n1835, n1747, n1739, n1731}), .out(n10526), .config_in(config_chain[17315:17310]), .config_rst(config_rst)); 
buffer_wire buffer_10526 (.in(n10526), .out(n10526_0));
mux15 mux_5361 (.in({n13693_1, n13684_0, n13679_0, n13667_0, n13649_1, n13644_0, n13640_0, n13586_0, n13563_0, n10607_1, n4777, n4769, n4681, n4673, n4665}), .out(n10527), .config_in(config_chain[17321:17316]), .config_rst(config_rst)); 
buffer_wire buffer_10527 (.in(n10527), .out(n10527_0));
mux16 mux_5362 (.in({n12657_1, n12642_0/**/, n12639_0, n12633_0, n12616_0, n12615_1, n12606_0, n12582_0, n12580_0, n12567_0, n10442_0, n1843, n1835, n1747, n1739, n1731}), .out(n10528), .config_in(config_chain[17327:17322]), .config_rst(config_rst)); 
buffer_wire buffer_10528 (.in(n10528), .out(n10528_0));
mux15 mux_5363 (.in({n13713_1, n13687_0, n13658_0, n13653_0, n13651_1, n13646_0, n13618_0, n13595_0, n13560_0, n10609_1, n4781, n4769, n4681, n4673/**/, n4665}), .out(n10529), .config_in(config_chain[17333:17328]), .config_rst(config_rst)); 
buffer_wire buffer_10529 (.in(n10529), .out(n10529_0));
mux15 mux_5364 (.in({n12659_1, n12653_0, n12636_0, n12630_0, n12627_0, n12608_0, n12572_0, n12558_0/**/, n12543_0, n10450_0, n1843, n1835, n1747, n1739, n1731}), .out(n10530), .config_in(config_chain[17339:17334]), .config_rst(config_rst)); 
buffer_wire buffer_10530 (.in(n10530), .out(n10530_0));
mux15 mux_5365 (.in({n13711_1, n13678_0, n13673_0, n13666_0, n13661_0, n13648_0, n13627_0, n13568_0, n13562_0, n10611_1, n4781, n4773, n4681, n4673/**/, n4665}), .out(n10531), .config_in(config_chain[17345:17340]), .config_rst(config_rst)); 
buffer_wire buffer_10531 (.in(n10531), .out(n10531_0));
mux15 mux_5366 (.in({n12661_1, n12650_0, n12647_0, n12624_0, n12621_0, n12610_0, n12599_0, n12564_0, n12534_0, n10458_0, n1843, n1835, n1747, n1739, n1731}), .out(n10532), .config_in(config_chain[17351:17346]), .config_rst(config_rst)); 
buffer_wire buffer_10532 (.in(n10532), .out(n10532_0));
mux15 mux_5367 (.in({n13709_1, n13686_0, n13681_0, n13669_0/**/, n13652_0, n13650_0, n13594_0, n13576_0, n13571_0, n10613_1, n4781, n4773, n4765, n4673, n4665}), .out(n10533), .config_in(config_chain[17357:17352]), .config_rst(config_rst)); 
buffer_wire buffer_10533 (.in(n10533), .out(n10533_0));
mux15 mux_5368 (.in({n12663_1, n12644_0, n12641_0, n12635_0/**/, n12618_0, n12612_0, n12590_0, n12575_0, n12556_0, n10466_0, n1843, n1835, n1747, n1739, n1731}), .out(n10534), .config_in(config_chain[17363:17358]), .config_rst(config_rst)); 
buffer_wire buffer_10534 (.in(n10534), .out(n10534_0));
mux14 mux_5369 (.in({n13707_1, n13689_0, n13672_0, n13660_0, n13655_0, n13626_0, n13603_0, n13584_0, n10615_1, n4781, n4773/**/, n4765, n4677, n4665}), .out(n10535), .config_in(config_chain[17369:17364]), .config_rst(config_rst)); 
buffer_wire buffer_10535 (.in(n10535), .out(n10535_0));
mux15 mux_5370 (.in({n12665_1, n12655_0, n12638_0, n12632_0/**/, n12629_0, n12614_0, n12566_0, n12551_0, n12548_0, n10474_0, n1847, n1839, n1831, n1743, n1735}), .out(n10536), .config_in(config_chain[17375:17370]), .config_rst(config_rst)); 
buffer_wire buffer_10536 (.in(n10536), .out(n10536_0));
mux14 mux_5371 (.in({n13705_1, n13680_0/**/, n13675_0, n13668_0, n13663_0, n13635_0, n13592_0, n13570_0, n10617_1, n4781, n4773, n4765, n4677, n4669}), .out(n10537), .config_in(config_chain[17381:17376]), .config_rst(config_rst)); 
buffer_wire buffer_10537 (.in(n10537), .out(n10537_0));
mux15 mux_5372 (.in({n12667_1/**/, n12652_0, n12649_0, n12626_0, n12623_0, n12605_1, n12542_0, n12540_0, n12527_0, n10482_0, n1847, n1839, n1831, n1743, n1735}), .out(n10538), .config_in(config_chain[17387:17382]), .config_rst(config_rst)); 
buffer_wire buffer_10538 (.in(n10538), .out(n10538_0));
mux13 mux_5373 (.in({n13703_1, n13688_0, n13683_0, n13671_0, n13654_0, n13602_0, n13600_0/**/, n13579_0, n10619_1, n4773, n4765, n4677, n4669}), .out(n10539), .config_in(config_chain[17393:17388]), .config_rst(config_rst)); 
buffer_wire buffer_10539 (.in(n10539), .out(n10539_0));
mux15 mux_5374 (.in({n12669_1/**/, n12646_0, n12643_0, n12620_0, n12617_0, n12607_1, n12598_0, n12583_0, n12532_0, n10490_0, n1847, n1839, n1831, n1743, n1735}), .out(n10540), .config_in(config_chain[17399:17394]), .config_rst(config_rst)); 
buffer_wire buffer_10540 (.in(n10540), .out(n10540_0));
mux13 mux_5375 (.in({n13701_1, n13691_0, n13674_0, n13662_0, n13657_0, n13634_0, n13611_0, n13608_0/**/, n10621_1, n4777, n4765, n4677, n4669}), .out(n10541), .config_in(config_chain[17405:17400]), .config_rst(config_rst)); 
buffer_wire buffer_10541 (.in(n10541), .out(n10541_0));
mux15 mux_5376 (.in({n12671_1, n12640_0, n12637_0, n12634_0, n12631_0/**/, n12609_1, n12574_0, n12559_0, n12524_0, n10498_0, n1847, n1839, n1831, n1743, n1735}), .out(n10542), .config_in(config_chain[17411:17406]), .config_rst(config_rst)); 
buffer_wire buffer_10542 (.in(n10542), .out(n10542_0));
mux13 mux_5377 (.in({n13699_1, n13682_0, n13677_0, n13670_0, n13665_0, n13643_0, n13616_0/**/, n13578_0, n10623_1, n4777, n4769, n4677, n4669}), .out(n10543), .config_in(config_chain[17417:17412]), .config_rst(config_rst)); 
buffer_wire buffer_10543 (.in(n10543), .out(n10543_0));
mux15 mux_5378 (.in({n12673_1, n12654_0, n12651_0, n12628_0, n12625_0, n12611_1, n12596_0, n12550_0, n12535_0, n10506_0, n1847, n1839/**/, n1831, n1743, n1735}), .out(n10544), .config_in(config_chain[17423:17418]), .config_rst(config_rst)); 
buffer_wire buffer_10544 (.in(n10544), .out(n10544_0));
mux13 mux_5379 (.in({n13697_1, n13690_0/**/, n13685_0, n13656_0, n13645_0, n13624_0, n13610_0, n13587_0, n10625_1, n4777, n4769, n4681, n4669}), .out(n10545), .config_in(config_chain[17429:17424]), .config_rst(config_rst)); 
buffer_wire buffer_10545 (.in(n10545), .out(n10545_0));
mux16 mux_5380 (.in({n12931_1, n12909_0, n12892_0, n12884_0, n12881_0, n12869_1, n12860_0, n12846_0, n12808_0, n12793_0, n10436_0/**/, n2821, n2813, n2725, n2717, n2709}), .out(n10546), .config_in(config_chain[17435:17430]), .config_rst(config_rst)); 
buffer_wire buffer_10546 (.in(n10546), .out(n10546_0));
mux15 mux_5381 (.in({n13959_1, n13942_0, n13937_0, n13928_0, n13923_0, n13913_0, n13908_0, n13906_0, n13885_0, n10629_0, n5755, n5747, n5659, n5651, n5643}), .out(n10547), .config_in(config_chain[17441:17436]), .config_rst(config_rst)); 
buffer_wire buffer_10547 (.in(n10547), .out(n10547_0));
mux16 mux_5382 (.in({n12913_1, n12906_0/**/, n12903_0, n12878_0, n12875_0, n12871_1, n12862_0, n12849_0, n12838_0, n12784_0, n10444_0, n2821, n2813, n2725, n2717, n2709}), .out(n10548), .config_in(config_chain[17447:17442]), .config_rst(config_rst)); 
buffer_wire buffer_10548 (.in(n10548), .out(n10548_0));
mux15 mux_5383 (.in({n13979_1, n13950_0, n13945_0, n13931_0, n13915_1, n13910_0, n13852_0, n13829_0, n13826_0, n10631_0/**/, n5759, n5747, n5659, n5651, n5643}), .out(n10549), .config_in(config_chain[17453:17448]), .config_rst(config_rst)); 
buffer_wire buffer_10549 (.in(n10549), .out(n10549_0));
mux15 mux_5384 (.in({n12915_1, n12900_0, n12897_0, n12889_0, n12872_0, n12864_0, n12840_0, n12830_0, n12825_0/**/, n10452_0, n2821, n2813, n2725, n2717, n2709}), .out(n10550), .config_in(config_chain[17459:17454]), .config_rst(config_rst)); 
buffer_wire buffer_10550 (.in(n10550), .out(n10550_0));
mux15 mux_5385 (.in({n13977_1, n13953_0/**/, n13936_0, n13922_0, n13917_0, n13912_0, n13884_0, n13861_0, n13834_0, n10633_0, n5759, n5751, n5659, n5651, n5643}), .out(n10551), .config_in(config_chain[17465:17460]), .config_rst(config_rst)); 
buffer_wire buffer_10551 (.in(n10551), .out(n10551_0));
mux15 mux_5386 (.in({n12917_1, n12911_0, n12894_0, n12886_0, n12883_0, n12866_0, n12822_0, n12816_0, n12801_0, n10460_0/**/, n2821, n2813, n2725, n2717, n2709}), .out(n10552), .config_in(config_chain[17471:17466]), .config_rst(config_rst)); 
buffer_wire buffer_10552 (.in(n10552), .out(n10552_0));
mux15 mux_5387 (.in({n13975_1, n13944_0, n13939_0, n13930_0, n13925_0, n13914_0, n13893_0, n13842_0, n13828_0, n10635_0, n5759, n5751, n5743, n5651, n5643}), .out(n10553), .config_in(config_chain[17477:17472]), .config_rst(config_rst)); 
buffer_wire buffer_10553 (.in(n10553), .out(n10553_0));
mux15 mux_5388 (.in({n12919_1, n12908_0, n12905_0, n12880_0, n12877_0, n12868_0, n12857_0, n12814_0/**/, n12792_0, n10468_0, n2821, n2813, n2725, n2717, n2709}), .out(n10554), .config_in(config_chain[17483:17478]), .config_rst(config_rst)); 
buffer_wire buffer_10554 (.in(n10554), .out(n10554_0));
mux14 mux_5389 (.in({n13973_1, n13952_0, n13947_0, n13933_0, n13916_0/**/, n13860_0, n13850_0, n13837_0, n10637_0, n5759, n5751, n5743, n5655, n5643}), .out(n10555), .config_in(config_chain[17489:17484]), .config_rst(config_rst)); 
buffer_wire buffer_10555 (.in(n10555), .out(n10555_0));
mux15 mux_5390 (.in({n12921_1, n12902_0, n12899_0, n12891_0, n12874_0, n12870_0, n12848_0, n12833_0, n12806_0/**/, n10476_0, n2825, n2817, n2809, n2721, n2713}), .out(n10556), .config_in(config_chain[17495:17490]), .config_rst(config_rst)); 
buffer_wire buffer_10556 (.in(n10556), .out(n10556_0));
mux14 mux_5391 (.in({n13971_1, n13955_0, n13938_0, n13924_0, n13919_0/**/, n13892_0, n13869_0, n13858_0, n10639_0, n5759, n5751, n5743, n5655, n5647}), .out(n10557), .config_in(config_chain[17501:17496]), .config_rst(config_rst)); 
buffer_wire buffer_10557 (.in(n10557), .out(n10557_0));
mux15 mux_5392 (.in({n12923_1, n12896_0, n12893_0, n12888_0, n12885_0, n12861_0, n12824_0, n12809_0/**/, n12798_0, n10484_0, n2825, n2817, n2809, n2721, n2713}), .out(n10558), .config_in(config_chain[17507:17502]), .config_rst(config_rst)); 
buffer_wire buffer_10558 (.in(n10558), .out(n10558_0));
mux13 mux_5393 (.in({n13969_1/**/, n13946_0, n13941_0, n13932_0, n13927_0, n13901_0, n13866_0, n13836_0, n10641_0, n5751, n5743, n5655, n5647}), .out(n10559), .config_in(config_chain[17513:17508]), .config_rst(config_rst)); 
buffer_wire buffer_10559 (.in(n10559), .out(n10559_0));
mux15 mux_5394 (.in({n12925_1, n12910_0, n12907_0, n12882_0, n12879_0, n12863_1, n12800_0, n12790_0/**/, n12785_0, n10492_0, n2825, n2817, n2809, n2721, n2713}), .out(n10560), .config_in(config_chain[17519:17514]), .config_rst(config_rst)); 
buffer_wire buffer_10560 (.in(n10560), .out(n10560_0));
mux13 mux_5395 (.in({n13967_1/**/, n13954_0, n13949_0, n13935_0, n13918_0, n13874_0, n13868_0, n13845_0, n10643_0, n5755, n5743, n5655, n5647}), .out(n10561), .config_in(config_chain[17525:17520]), .config_rst(config_rst)); 
buffer_wire buffer_10561 (.in(n10561), .out(n10561_0));
mux15 mux_5396 (.in({n12927_1, n12904_0, n12901_0, n12876_0, n12873_0, n12865_1, n12856_0, n12841_0/**/, n12782_0, n10500_0, n2825, n2817, n2809, n2721, n2713}), .out(n10562), .config_in(config_chain[17531:17526]), .config_rst(config_rst)); 
buffer_wire buffer_10562 (.in(n10562), .out(n10562_0));
mux13 mux_5397 (.in({n13965_1, n13957_1, n13940_0, n13926_0, n13921_0, n13900_0, n13882_0, n13877_0, n10645_0, n5755, n5747, n5655, n5647}), .out(n10563), .config_in(config_chain[17537:17532]), .config_rst(config_rst)); 
buffer_wire buffer_10563 (.in(n10563), .out(n10563_0));
mux15 mux_5398 (.in({n12929_1, n12898_0, n12895_0, n12890_0, n12887_0, n12867_1, n12854_0, n12832_0, n12817_0, n10508_0/**/, n2825, n2817, n2809, n2721, n2713}), .out(n10564), .config_in(config_chain[17543:17538]), .config_rst(config_rst)); 
buffer_wire buffer_10564 (.in(n10564), .out(n10564_0));
mux13 mux_5399 (.in({n13963_1, n13948_0, n13943_0, n13934_0, n13929_0, n13909_0, n13890_0, n13844_0/**/, n10647_0, n5755, n5747, n5659, n5647}), .out(n10565), .config_in(config_chain[17549:17544]), .config_rst(config_rst)); 
buffer_wire buffer_10565 (.in(n10565), .out(n10565_0));
mux16 mux_5400 (.in({n13189_1, n13156_0, n13153_0, n13147_0, n13130_0, n13127_1, n13118_0, n13106_0, n13092_0, n13077_0, n10438_0, n3799, n3791/**/, n3703, n3695, n3687}), .out(n10566), .config_in(config_chain[17555:17550]), .config_rst(config_rst)); 
buffer_wire buffer_10566 (.in(n10566), .out(n10566_0));
mux15 mux_5401 (.in({n14225_1, n14222_0, n14217_0, n14186_0, n14181_0, n14177_0, n14172_0, n14142_0, n14119_0, n10651_0, n6733, n6725, n6637, n6629/**/, n6621}), .out(n10567), .config_in(config_chain[17561:17556]), .config_rst(config_rst)); 
buffer_wire buffer_10567 (.in(n10567), .out(n10567_0));
mux16 mux_5402 (.in({n13171_1, n13167_0, n13150_0, n13144_0, n13141_0, n13129_1, n13120_0, n13098_0, n13068_0, n13053_0, n10446_0, n3799, n3791, n3703/**/, n3695, n3687}), .out(n10568), .config_in(config_chain[17567:17562]), .config_rst(config_rst)); 
buffer_wire buffer_10568 (.in(n10568), .out(n10568_0));
mux15 mux_5403 (.in({n14245_1, n14208_0, n14203_0, n14194_0, n14189_0, n14179_0, n14174_0, n14151_0, n14092_0, n10653_0, n6737, n6725, n6637/**/, n6629, n6621}), .out(n10569), .config_in(config_chain[17573:17568]), .config_rst(config_rst)); 
buffer_wire buffer_10569 (.in(n10569), .out(n10569_0));
mux15 mux_5404 (.in({n13173_1, n13164_0, n13161_0, n13138_0, n13135_0, n13122_0, n13109_0, n13090_0, n13044_0/**/, n10454_0, n3799, n3791, n3703, n3695, n3687}), .out(n10570), .config_in(config_chain[17579:17574]), .config_rst(config_rst)); 
buffer_wire buffer_10570 (.in(n10570), .out(n10570_0));
mux15 mux_5405 (.in({n14243_1, n14216_0, n14211_0, n14197_0, n14180_0, n14176_0, n14118_0, n14100_0, n14095_0, n10655_0, n6737, n6729, n6637, n6629/**/, n6621}), .out(n10571), .config_in(config_chain[17585:17580]), .config_rst(config_rst)); 
buffer_wire buffer_10571 (.in(n10571), .out(n10571_0));
mux15 mux_5406 (.in({n13175_1, n13158_0, n13155_0, n13149_0, n13132_0, n13124_0, n13100_0, n13085_0, n13082_0, n10462_0, n3799, n3791, n3703, n3695, n3687/**/}), .out(n10572), .config_in(config_chain[17591:17586]), .config_rst(config_rst)); 
buffer_wire buffer_10572 (.in(n10572), .out(n10572_0));
mux15 mux_5407 (.in({n14241_1, n14219_0, n14202_0, n14188_0, n14183_0, n14178_0, n14150_0, n14127_0, n14108_0, n10657_0/**/, n6737, n6729, n6721, n6629, n6621}), .out(n10573), .config_in(config_chain[17597:17592]), .config_rst(config_rst)); 
buffer_wire buffer_10573 (.in(n10573), .out(n10573_0));
mux15 mux_5408 (.in({n13177_1, n13169_0, n13152_0, n13146_0, n13143_0, n13126_0, n13076_0, n13074_0, n13061_0, n10470_0, n3799/**/, n3791, n3703, n3695, n3687}), .out(n10574), .config_in(config_chain[17603:17598]), .config_rst(config_rst)); 
buffer_wire buffer_10574 (.in(n10574), .out(n10574_0));
mux14 mux_5409 (.in({n14239_1, n14210_0, n14205_0, n14196_0, n14191_0, n14159_0/**/, n14116_0, n14094_0, n10659_0, n6737, n6729, n6721, n6633, n6621}), .out(n10575), .config_in(config_chain[17609:17604]), .config_rst(config_rst)); 
buffer_wire buffer_10575 (.in(n10575), .out(n10575_0));
mux15 mux_5410 (.in({n13179_1, n13166_0/**/, n13163_0, n13140_0, n13137_0, n13128_0, n13117_0, n13066_0, n13052_0, n10478_0, n3803, n3795, n3787, n3699, n3691}), .out(n10576), .config_in(config_chain[17615:17610]), .config_rst(config_rst)); 
buffer_wire buffer_10576 (.in(n10576), .out(n10576_0));
mux14 mux_5411 (.in({n14237_1, n14218_0, n14213_0, n14199_0, n14182_0, n14126_0, n14124_0, n14103_0, n10661_0, n6737, n6729, n6721, n6633, n6625/**/}), .out(n10577), .config_in(config_chain[17621:17616]), .config_rst(config_rst)); 
buffer_wire buffer_10577 (.in(n10577), .out(n10577_0));
mux15 mux_5412 (.in({n13181_1, n13160_0, n13157_0, n13134_0, n13131_0, n13119_0, n13108_0, n13093_0/**/, n13058_0, n10486_0, n3803, n3795, n3787, n3699, n3691}), .out(n10578), .config_in(config_chain[17627:17622]), .config_rst(config_rst)); 
buffer_wire buffer_10578 (.in(n10578), .out(n10578_0));
mux13 mux_5413 (.in({n14235_1, n14221_0, n14204_0, n14190_0, n14185_0, n14158_0, n14135_0, n14132_0, n10663_0, n6729, n6721/**/, n6633, n6625}), .out(n10579), .config_in(config_chain[17633:17628]), .config_rst(config_rst)); 
buffer_wire buffer_10579 (.in(n10579), .out(n10579_0));
mux15 mux_5414 (.in({n13183_1, n13154_0, n13151_0, n13148_0, n13145_0/**/, n13121_0, n13084_0, n13069_0, n13050_0, n10494_0, n3803, n3795, n3787, n3699, n3691}), .out(n10580), .config_in(config_chain[17639:17634]), .config_rst(config_rst)); 
buffer_wire buffer_10580 (.in(n10580), .out(n10580_0));
mux13 mux_5415 (.in({n14233_1, n14212_0/**/, n14207_0, n14198_0, n14193_0, n14167_0, n14140_0, n14102_0, n10665_0, n6733, n6721, n6633, n6625}), .out(n10581), .config_in(config_chain[17645:17640]), .config_rst(config_rst)); 
buffer_wire buffer_10581 (.in(n10581), .out(n10581_0));
mux15 mux_5416 (.in({n13185_1, n13168_0, n13165_0, n13142_0, n13139_0, n13123_1, n13060_0, n13045_0, n13042_0, n10502_0, n3803, n3795/**/, n3787, n3699, n3691}), .out(n10582), .config_in(config_chain[17651:17646]), .config_rst(config_rst)); 
buffer_wire buffer_10582 (.in(n10582), .out(n10582_0));
mux13 mux_5417 (.in({n14231_1, n14220_0, n14215_0, n14201_1, n14184_0, n14148_0, n14134_0, n14111_0, n10667_0/**/, n6733, n6725, n6633, n6625}), .out(n10583), .config_in(config_chain[17657:17652]), .config_rst(config_rst)); 
buffer_wire buffer_10583 (.in(n10583), .out(n10583_0));
mux15 mux_5418 (.in({n13187_1, n13162_0, n13159_0, n13136_0, n13133_0/**/, n13125_1, n13116_0, n13114_0, n13101_0, n10510_0, n3803, n3795, n3787, n3699, n3691}), .out(n10584), .config_in(config_chain[17663:17658]), .config_rst(config_rst)); 
buffer_wire buffer_10584 (.in(n10584), .out(n10584_0));
mux13 mux_5419 (.in({n14229_1, n14223_1, n14206_0, n14192_0, n14187_0, n14166_0/**/, n14156_0, n14143_0, n10669_0, n6733, n6725, n6637, n6625}), .out(n10585), .config_in(config_chain[17669:17664]), .config_rst(config_rst)); 
buffer_wire buffer_10585 (.in(n10585), .out(n10585_0));
mux16 mux_5420 (.in({n13449_1, n13422_0, n13419_0, n13396_0, n13393_0, n13387_1, n13378_0, n13368_0, n13363_0, n13298_0, n10440_1, n4777, n4769, n4681, n4673, n4665}), .out(n10586), .config_in(config_chain[17675:17670]), .config_rst(config_rst)); 
buffer_wire buffer_10586 (.in(n10586), .out(n10586_0));
mux15 mux_5421 (.in({n14489_1, n14478_0, n14473_0, n14464_0, n14459_0, n14441_0, n14438_0, n14376_0, n14353_0, n10673_0, n7711/**/, n7703, n7615, n7607, n7599}), .out(n10587), .config_in(config_chain[17681:17676]), .config_rst(config_rst)); 
buffer_wire buffer_10587 (.in(n10587), .out(n10587_0));
mux16 mux_5422 (.in({n13431_1, n13416_0, n13413_0, n13407_0, n13390_0, n13389_1, n13380_0, n13360_0, n13354_0, n13339_0, n10448_1, n4777, n4769, n4681/**/, n4673, n4665}), .out(n10588), .config_in(config_chain[17687:17682]), .config_rst(config_rst)); 
buffer_wire buffer_10588 (.in(n10588), .out(n10588_0));
mux15 mux_5423 (.in({n14509_1, n14486_0, n14481_0, n14450_0, n14445_0, n14443_0, n14408_0, n14385_0, n14358_0, n10675_0, n7715, n7703, n7615, n7607, n7599/**/}), .out(n10589), .config_in(config_chain[17693:17688]), .config_rst(config_rst)); 
buffer_wire buffer_10589 (.in(n10589), .out(n10589_0));
mux15 mux_5424 (.in({n13433_1, n13427_0, n13410_0, n13404_0, n13401_0, n13382_0, n13352_0, n13330_0, n13315_0, n10456_1/**/, n4777, n4769, n4681, n4673, n4665}), .out(n10590), .config_in(config_chain[17699:17694]), .config_rst(config_rst)); 
buffer_wire buffer_10590 (.in(n10590), .out(n10590_0));
mux15 mux_5425 (.in({n14507_1, n14472_0/**/, n14467_0, n14458_0, n14453_0, n14440_0, n14417_0, n14366_0, n14352_0, n10677_0, n7715, n7707, n7615, n7607, n7599}), .out(n10591), .config_in(config_chain[17705:17700]), .config_rst(config_rst)); 
buffer_wire buffer_10591 (.in(n10591), .out(n10591_0));
mux15 mux_5426 (.in({n13435_1, n13424_0, n13421_0, n13398_0, n13395_0, n13384_0, n13371_0, n13344_0, n13306_0, n10464_1, n4777, n4769/**/, n4681, n4673, n4665}), .out(n10592), .config_in(config_chain[17711:17706]), .config_rst(config_rst)); 
buffer_wire buffer_10592 (.in(n10592), .out(n10592_0));
mux15 mux_5427 (.in({n14505_1, n14480_0, n14475_0, n14461_0, n14444_0, n14442_0, n14384_0/**/, n14374_0, n14361_0, n10679_0, n7715, n7707, n7699, n7607, n7599}), .out(n10593), .config_in(config_chain[17717:17712]), .config_rst(config_rst)); 
buffer_wire buffer_10593 (.in(n10593), .out(n10593_0));
mux15 mux_5428 (.in({n13437_1, n13418_0, n13415_0, n13409_0, n13392_0, n13386_0, n13362_0/**/, n13347_0, n13336_0, n10472_1, n4777, n4769, n4681, n4673, n4665}), .out(n10594), .config_in(config_chain[17723:17718]), .config_rst(config_rst)); 
buffer_wire buffer_10594 (.in(n10594), .out(n10594_0));
mux14 mux_5429 (.in({n14503_1, n14483_0, n14466_0, n14452_0, n14447_0, n14416_0, n14393_0, n14382_0, n10681_0, n7715, n7707, n7699/**/, n7611, n7599}), .out(n10595), .config_in(config_chain[17729:17724]), .config_rst(config_rst)); 
buffer_wire buffer_10595 (.in(n10595), .out(n10595_0));
mux15 mux_5430 (.in({n13439_1, n13429_0, n13412_0, n13406_0, n13403_0, n13388_0, n13338_0, n13328_0, n13323_0, n10480_1, n4781, n4773, n4765, n4677/**/, n4669}), .out(n10596), .config_in(config_chain[17735:17730]), .config_rst(config_rst)); 
buffer_wire buffer_10596 (.in(n10596), .out(n10596_0));
mux14 mux_5431 (.in({n14501_1, n14474_0, n14469_0, n14460_0, n14455_0, n14425_0, n14390_0, n14360_0, n10683_0, n7715, n7707, n7699, n7611/**/, n7603}), .out(n10597), .config_in(config_chain[17741:17736]), .config_rst(config_rst)); 
buffer_wire buffer_10597 (.in(n10597), .out(n10597_0));
mux15 mux_5432 (.in({n13441_1/**/, n13426_0, n13423_0, n13400_0, n13397_0, n13379_0, n13320_0, n13314_0, n13299_0, n10488_1, n4781, n4773, n4765, n4677, n4669}), .out(n10598), .config_in(config_chain[17747:17742]), .config_rst(config_rst)); 
buffer_wire buffer_10598 (.in(n10598), .out(n10598_0));
mux13 mux_5433 (.in({n14499_1, n14482_0, n14477_0, n14463_0, n14446_0, n14398_0, n14392_0/**/, n14369_0, n10685_0, n7707, n7699, n7611, n7603}), .out(n10599), .config_in(config_chain[17753:17748]), .config_rst(config_rst)); 
buffer_wire buffer_10599 (.in(n10599), .out(n10599_0));
mux15 mux_5434 (.in({n13443_1, n13420_0, n13417_0, n13394_0, n13391_0, n13381_0, n13370_0, n13355_0, n13312_0/**/, n10496_1, n4781, n4773, n4765, n4677, n4669}), .out(n10600), .config_in(config_chain[17759:17754]), .config_rst(config_rst)); 
buffer_wire buffer_10600 (.in(n10600), .out(n10600_0));
mux13 mux_5435 (.in({n14497_1, n14485_0, n14468_0, n14454_0, n14449_0, n14424_0, n14406_0, n14401_0, n10687_0, n7711, n7699, n7611, n7603}), .out(n10601), .config_in(config_chain[17765:17760]), .config_rst(config_rst)); 
buffer_wire buffer_10601 (.in(n10601), .out(n10601_0));
mux15 mux_5436 (.in({n13445_1, n13414_0, n13411_0, n13408_0, n13405_0/**/, n13383_0, n13346_0, n13331_0, n13304_0, n10504_1, n4781, n4773, n4765, n4677, n4669}), .out(n10602), .config_in(config_chain[17771:17766]), .config_rst(config_rst)); 
buffer_wire buffer_10602 (.in(n10602), .out(n10602_0));
mux13 mux_5437 (.in({n14495_1, n14476_0/**/, n14471_0, n14462_0, n14457_0, n14433_1, n14414_0, n14368_0, n10689_0, n7711, n7703, n7611, n7603}), .out(n10603), .config_in(config_chain[17777:17772]), .config_rst(config_rst)); 
buffer_wire buffer_10603 (.in(n10603), .out(n10603_0));
mux15 mux_5438 (.in({n13447_1, n13428_0/**/, n13425_0, n13402_0, n13399_0, n13385_1, n13376_0, n13322_0, n13307_0, n10512_1, n4781, n4773, n4765, n4677, n4669}), .out(n10604), .config_in(config_chain[17783:17778]), .config_rst(config_rst)); 
buffer_wire buffer_10604 (.in(n10604), .out(n10604_0));
mux13 mux_5439 (.in({n14493_1, n14484_0, n14479_0, n14465_1, n14448_0, n14422_0, n14400_0, n14377_0/**/, n10691_0, n7711, n7703, n7615, n7603}), .out(n10605), .config_in(config_chain[17789:17784]), .config_rst(config_rst)); 
buffer_wire buffer_10605 (.in(n10605), .out(n10605_0));
mux15 mux_5440 (.in({n13713_1, n13685_0, n13678_0, n13666_0, n13648_0, n13645_0, n13632_0/**/, n13587_0, n13562_0, n10526_1, n5755, n5747, n5659, n5651, n5643}), .out(n10606), .config_in(config_chain[17795:17790]), .config_rst(config_rst)); 
buffer_wire buffer_10606 (.in(n10606), .out(n10606_0));
mux4 mux_5441 (.in({n14751_1/**/, n14614_0, n8693, n8577}), .out(n10607), .config_in(config_chain[17797:17796]), .config_rst(config_rst)); 
buffer_wire buffer_10607 (.in(n10607), .out(n10607_0));
mux15 mux_5442 (.in({n13693_1, n13686_0, n13659_0, n13652_0, n13650_0, n13647_0, n13624_0, n13619_0, n13594_0, n10528_1, n5759, n5747, n5659, n5651, n5643/**/}), .out(n10608), .config_in(config_chain[17803:17798]), .config_rst(config_rst)); 
buffer_wire buffer_10608 (.in(n10608), .out(n10608_0));
mux3 mux_5443 (.in({n14753_1/**/, n14622_0, n8577}), .out(n10609), .config_in(config_chain[17805:17804]), .config_rst(config_rst)); 
buffer_wire buffer_10609 (.in(n10609), .out(n10609_0));
mux15 mux_5444 (.in({n13695_1/**/, n13679_0, n13672_0, n13667_0, n13660_0, n13649_1, n13626_0, n13616_0, n13563_0, n10530_1, n5759, n5751, n5659, n5651, n5643}), .out(n10610), .config_in(config_chain[17811:17806]), .config_rst(config_rst)); 
buffer_wire buffer_10610 (.in(n10610), .out(n10610_0));
mux3 mux_5445 (.in({n14755_1/**/, n14630_0, n8581}), .out(n10611), .config_in(config_chain[17813:17812]), .config_rst(config_rst)); 
buffer_wire buffer_10611 (.in(n10611), .out(n10611_0));
mux15 mux_5446 (.in({n13697_1, n13687_0, n13680_0, n13668_0, n13653_0, n13651_1, n13608_0, n13595_0/**/, n13570_0, n10532_1, n5759, n5751, n5743, n5651, n5643}), .out(n10612), .config_in(config_chain[17819:17814]), .config_rst(config_rst)); 
buffer_wire buffer_10612 (.in(n10612), .out(n10612_0));
mux3 mux_5447 (.in({n14757_1/**/, n14638_0, n8585}), .out(n10613), .config_in(config_chain[17821:17820]), .config_rst(config_rst)); 
buffer_wire buffer_10613 (.in(n10613), .out(n10613_0));
mux14 mux_5448 (.in({n13699_1/**/, n13688_0, n13673_0, n13661_0, n13654_0, n13627_0, n13602_0, n13600_0, n10534_1, n5759, n5751, n5743, n5655, n5643}), .out(n10614), .config_in(config_chain[17827:17822]), .config_rst(config_rst)); 
buffer_wire buffer_10614 (.in(n10614), .out(n10614_0));
mux3 mux_5449 (.in({n14759_1, n14646_0, n8589/**/}), .out(n10615), .config_in(config_chain[17829:17828]), .config_rst(config_rst)); 
buffer_wire buffer_10615 (.in(n10615), .out(n10615_0));
mux14 mux_5450 (.in({n13701_1, n13681_0, n13674_0, n13669_0, n13662_0, n13634_0, n13592_0, n13571_0, n10536_1, n5759, n5751/**/, n5743, n5655, n5647}), .out(n10616), .config_in(config_chain[17835:17830]), .config_rst(config_rst)); 
buffer_wire buffer_10616 (.in(n10616), .out(n10616_0));
mux3 mux_5451 (.in({n14761_1, n14654_0, n8593}), .out(n10617), .config_in(config_chain[17837:17836]), .config_rst(config_rst)); 
buffer_wire buffer_10617 (.in(n10617), .out(n10617_0));
mux13 mux_5452 (.in({n13703_1, n13689_0, n13682_0, n13670_0, n13655_0/**/, n13603_0, n13584_0, n13578_0, n10538_1, n5751, n5743, n5655, n5647}), .out(n10618), .config_in(config_chain[17843:17838]), .config_rst(config_rst)); 
buffer_wire buffer_10618 (.in(n10618), .out(n10618_0));
mux3 mux_5453 (.in({n14763_1/**/, n14662_0, n8593}), .out(n10619), .config_in(config_chain[17845:17844]), .config_rst(config_rst)); 
buffer_wire buffer_10619 (.in(n10619), .out(n10619_0));
mux13 mux_5454 (.in({n13705_1, n13690_0/**/, n13675_0, n13663_0, n13656_0, n13635_0, n13610_0, n13576_0, n10540_1, n5755, n5743, n5655, n5647}), .out(n10620), .config_in(config_chain[17851:17846]), .config_rst(config_rst)); 
buffer_wire buffer_10620 (.in(n10620), .out(n10620_0));
mux3 mux_5455 (.in({n14765_1, n14670_0, n8677}), .out(n10621), .config_in(config_chain[17853:17852]), .config_rst(config_rst)); 
buffer_wire buffer_10621 (.in(n10621), .out(n10621_0));
mux13 mux_5456 (.in({n13707_1, n13683_0, n13676_0, n13671_0, n13664_0, n13642_0, n13579_0, n13568_0, n10542_1/**/, n5755, n5747, n5655, n5647}), .out(n10622), .config_in(config_chain[17859:17854]), .config_rst(config_rst)); 
buffer_wire buffer_10622 (.in(n10622), .out(n10622_0));
mux3 mux_5457 (.in({n14767_1, n14678_0, n8681/**/}), .out(n10623), .config_in(config_chain[17861:17860]), .config_rst(config_rst)); 
buffer_wire buffer_10623 (.in(n10623), .out(n10623_0));
mux13 mux_5458 (.in({n13709_1, n13691_0, n13684_0, n13657_0, n13644_0, n13611_0, n13586_0, n13560_0, n10544_1, n5755, n5747, n5659, n5647}), .out(n10624), .config_in(config_chain[17867:17862]), .config_rst(config_rst)); 
buffer_wire buffer_10624 (.in(n10624), .out(n10624_0));
mux3 mux_5459 (.in({n14769_1, n14686_0/**/, n8685}), .out(n10625), .config_in(config_chain[17869:17868]), .config_rst(config_rst)); 
buffer_wire buffer_10625 (.in(n10625), .out(n10625_0));
mux13 mux_5460 (.in({n13711_1/**/, n13677_0, n13665_0, n13658_0, n13646_0, n13643_0, n13640_0, n13618_0, n10514_1, n5755, n5747, n5659, n5651}), .out(n10626), .config_in(config_chain[17875:17870]), .config_rst(config_rst)); 
buffer_wire buffer_10626 (.in(n10626), .out(n10626_0));
mux3 mux_5461 (.in({n14695_1, n14694_0, n8689}), .out(n10627), .config_in(config_chain[17877:17876]), .config_rst(config_rst)); 
buffer_wire buffer_10627 (.in(n10627), .out(n10627_0));
mux15 mux_5462 (.in({n13979_1, n13943_0, n13936_0, n13929_0, n13922_0, n13912_0, n13909_0/**/, n13898_0, n13884_0, n10546_1, n6733, n6725, n6637, n6629, n6621}), .out(n10628), .config_in(config_chain[17883:17878]), .config_rst(config_rst)); 
buffer_wire buffer_10628 (.in(n10628), .out(n10628_0));
mux4 mux_5463 (.in({n14617_0, n14616_0, n8693, n8577}), .out(n10629), .config_in(config_chain[17885:17884]), .config_rst(config_rst)); 
buffer_wire buffer_10629 (.in(n10629), .out(n10629_0));
mux15 mux_5464 (.in({n13959_1, n13951_0, n13944_0, n13930_0, n13914_0, n13911_0, n13890_0, n13853_0, n13828_0, n10548_1/**/, n6737, n6725, n6637, n6629, n6621}), .out(n10630), .config_in(config_chain[17891:17886]), .config_rst(config_rst)); 
buffer_wire buffer_10630 (.in(n10630), .out(n10630_0));
mux3 mux_5465 (.in({n14625_0/**/, n14624_0, n8581}), .out(n10631), .config_in(config_chain[17893:17892]), .config_rst(config_rst)); 
buffer_wire buffer_10631 (.in(n10631), .out(n10631_0));
mux15 mux_5466 (.in({n13961_1, n13952_0, n13937_0/**/, n13923_0, n13916_0, n13913_0, n13885_0, n13882_0, n13860_0, n10550_1, n6737, n6729, n6637, n6629, n6621}), .out(n10632), .config_in(config_chain[17899:17894]), .config_rst(config_rst)); 
buffer_wire buffer_10632 (.in(n10632), .out(n10632_0));
mux3 mux_5467 (.in({n14633_0/**/, n14632_0, n8581}), .out(n10633), .config_in(config_chain[17901:17900]), .config_rst(config_rst)); 
buffer_wire buffer_10633 (.in(n10633), .out(n10633_0));
mux15 mux_5468 (.in({n13963_1, n13945_0, n13938_0, n13931_0/**/, n13924_0, n13915_1, n13892_0, n13874_0, n13829_0, n10552_1, n6737, n6729, n6721, n6629, n6621}), .out(n10634), .config_in(config_chain[17907:17902]), .config_rst(config_rst)); 
buffer_wire buffer_10634 (.in(n10634), .out(n10634_0));
mux3 mux_5469 (.in({n14641_0/**/, n14640_0, n8585}), .out(n10635), .config_in(config_chain[17909:17908]), .config_rst(config_rst)); 
buffer_wire buffer_10635 (.in(n10635), .out(n10635_0));
mux14 mux_5470 (.in({n13965_1, n13953_0, n13946_0, n13932_0, n13917_0, n13866_0, n13861_0, n13836_0, n10554_1/**/, n6737, n6729, n6721, n6633, n6621}), .out(n10636), .config_in(config_chain[17915:17910]), .config_rst(config_rst)); 
buffer_wire buffer_10636 (.in(n10636), .out(n10636_0));
mux3 mux_5471 (.in({n14649_0, n14648_0/**/, n8589}), .out(n10637), .config_in(config_chain[17917:17916]), .config_rst(config_rst)); 
buffer_wire buffer_10637 (.in(n10637), .out(n10637_0));
mux14 mux_5472 (.in({n13967_1/**/, n13954_0, n13939_0, n13925_0, n13918_0, n13893_0, n13868_0, n13858_0, n10556_1, n6737, n6729, n6721, n6633, n6625}), .out(n10638), .config_in(config_chain[17923:17918]), .config_rst(config_rst)); 
buffer_wire buffer_10638 (.in(n10638), .out(n10638_0));
mux3 mux_5473 (.in({n14657_0/**/, n14656_0, n8593}), .out(n10639), .config_in(config_chain[17925:17924]), .config_rst(config_rst)); 
buffer_wire buffer_10639 (.in(n10639), .out(n10639_0));
mux13 mux_5474 (.in({n13969_1, n13947_0, n13940_0, n13933_0, n13926_0, n13900_0, n13850_0, n13837_0, n10558_1/**/, n6729, n6721, n6633, n6625}), .out(n10640), .config_in(config_chain[17931:17926]), .config_rst(config_rst)); 
buffer_wire buffer_10640 (.in(n10640), .out(n10640_0));
mux3 mux_5475 (.in({n14665_0/**/, n14664_0, n8677}), .out(n10641), .config_in(config_chain[17933:17932]), .config_rst(config_rst)); 
buffer_wire buffer_10641 (.in(n10641), .out(n10641_0));
mux13 mux_5476 (.in({n13971_1, n13955_0, n13948_0/**/, n13934_0, n13919_0, n13869_0, n13844_0, n13842_0, n10560_1, n6733, n6721, n6633, n6625}), .out(n10642), .config_in(config_chain[17939:17934]), .config_rst(config_rst)); 
buffer_wire buffer_10642 (.in(n10642), .out(n10642_0));
mux3 mux_5477 (.in({n14673_0/**/, n14672_0, n8677}), .out(n10643), .config_in(config_chain[17941:17940]), .config_rst(config_rst)); 
buffer_wire buffer_10643 (.in(n10643), .out(n10643_0));
mux13 mux_5478 (.in({n13973_1, n13956_0, n13941_0, n13927_0, n13920_0, n13901_0, n13876_0, n13834_0, n10562_1/**/, n6733, n6725, n6633, n6625}), .out(n10644), .config_in(config_chain[17947:17942]), .config_rst(config_rst)); 
buffer_wire buffer_10644 (.in(n10644), .out(n10644_0));
mux3 mux_5479 (.in({n14681_0/**/, n14680_0, n8681}), .out(n10645), .config_in(config_chain[17949:17948]), .config_rst(config_rst)); 
buffer_wire buffer_10645 (.in(n10645), .out(n10645_0));
mux13 mux_5480 (.in({n13975_1, n13949_0, n13942_0, n13935_0, n13928_0, n13908_0, n13845_0, n13826_0/**/, n10564_1, n6733, n6725, n6637, n6625}), .out(n10646), .config_in(config_chain[17955:17950]), .config_rst(config_rst)); 
buffer_wire buffer_10646 (.in(n10646), .out(n10646_0));
mux3 mux_5481 (.in({n14689_0, n14688_0, n8685}), .out(n10647), .config_in(config_chain[17957:17956]), .config_rst(config_rst)); 
buffer_wire buffer_10647 (.in(n10647), .out(n10647_0));
mux13 mux_5482 (.in({n13977_1, n13957_1, n13950_0, n13921_0, n13910_0, n13906_0, n13877_0, n13852_0, n10516_1, n6733, n6725, n6637, n6629/**/}), .out(n10648), .config_in(config_chain[17963:17958]), .config_rst(config_rst)); 
buffer_wire buffer_10648 (.in(n10648), .out(n10648_0));
mux3 mux_5483 (.in({n14697_1, n14696_0, n8689}), .out(n10649), .config_in(config_chain[17965:17964]), .config_rst(config_rst)); 
buffer_wire buffer_10649 (.in(n10649), .out(n10649_0));
mux15 mux_5484 (.in({n14245_1, n14223_1, n14216_0, n14187_0, n14180_0, n14176_0, n14164_0, n14143_0, n14118_0, n10566_1, n7711, n7703, n7615, n7607, n7599/**/}), .out(n10650), .config_in(config_chain[17971:17966]), .config_rst(config_rst)); 
buffer_wire buffer_10650 (.in(n10650), .out(n10650_0));
mux4 mux_5485 (.in({n14707_0, n14706_0, n8693, n8577}), .out(n10651), .config_in(config_chain[17973:17972]), .config_rst(config_rst)); 
buffer_wire buffer_10651 (.in(n10651), .out(n10651_0));
mux15 mux_5486 (.in({n14225_1, n14209_0, n14202_0, n14195_0, n14188_0, n14178_0, n14175_0, n14156_0, n14150_0, n10568_1, n7715, n7703, n7615, n7607, n7599/**/}), .out(n10652), .config_in(config_chain[17979:17974]), .config_rst(config_rst)); 
buffer_wire buffer_10652 (.in(n10652), .out(n10652_0));
mux3 mux_5487 (.in({n14709_0/**/, n14708_0, n8581}), .out(n10653), .config_in(config_chain[17981:17980]), .config_rst(config_rst)); 
buffer_wire buffer_10653 (.in(n10653), .out(n10653_0));
mux15 mux_5488 (.in({n14227_1, n14217_0, n14210_0, n14196_0, n14181_0, n14177_0/**/, n14148_0, n14119_0, n14094_0, n10570_1, n7715, n7707, n7615, n7607, n7599}), .out(n10654), .config_in(config_chain[17987:17982]), .config_rst(config_rst)); 
buffer_wire buffer_10654 (.in(n10654), .out(n10654_0));
mux3 mux_5489 (.in({n14711_0, n14710_0, n8585}), .out(n10655), .config_in(config_chain[17989:17988]), .config_rst(config_rst)); 
buffer_wire buffer_10655 (.in(n10655), .out(n10655_0));
mux15 mux_5490 (.in({n14229_1, n14218_0, n14203_0, n14189_0, n14182_0, n14179_0, n14151_0, n14140_0, n14126_0, n10572_1, n7715, n7707, n7699, n7607, n7599/**/}), .out(n10656), .config_in(config_chain[17995:17990]), .config_rst(config_rst)); 
buffer_wire buffer_10656 (.in(n10656), .out(n10656_0));
mux3 mux_5491 (.in({n14713_0/**/, n14712_0, n8585}), .out(n10657), .config_in(config_chain[17997:17996]), .config_rst(config_rst)); 
buffer_wire buffer_10657 (.in(n10657), .out(n10657_0));
mux14 mux_5492 (.in({n14231_1, n14211_0, n14204_0, n14197_0, n14190_0, n14158_0/**/, n14132_0, n14095_0, n10574_1, n7715, n7707, n7699, n7611, n7599}), .out(n10658), .config_in(config_chain[18003:17998]), .config_rst(config_rst)); 
buffer_wire buffer_10658 (.in(n10658), .out(n10658_0));
mux3 mux_5493 (.in({n14715_0, n14714_0/**/, n8589}), .out(n10659), .config_in(config_chain[18005:18004]), .config_rst(config_rst)); 
buffer_wire buffer_10659 (.in(n10659), .out(n10659_0));
mux14 mux_5494 (.in({n14233_1, n14219_0, n14212_0, n14198_0, n14183_0, n14127_0, n14124_0, n14102_0, n10576_1, n7715, n7707, n7699, n7611, n7603/**/}), .out(n10660), .config_in(config_chain[18011:18006]), .config_rst(config_rst)); 
buffer_wire buffer_10660 (.in(n10660), .out(n10660_0));
mux3 mux_5495 (.in({n14717_0, n14716_0, n8593}), .out(n10661), .config_in(config_chain[18013:18012]), .config_rst(config_rst)); 
buffer_wire buffer_10661 (.in(n10661), .out(n10661_0));
mux13 mux_5496 (.in({n14235_1, n14220_0, n14205_0, n14191_0/**/, n14184_0, n14159_0, n14134_0, n14116_0, n10578_1, n7707, n7699, n7611, n7603}), .out(n10662), .config_in(config_chain[18019:18014]), .config_rst(config_rst)); 
buffer_wire buffer_10662 (.in(n10662), .out(n10662_0));
mux3 mux_5497 (.in({n14719_0/**/, n14718_0, n8677}), .out(n10663), .config_in(config_chain[18021:18020]), .config_rst(config_rst)); 
buffer_wire buffer_10663 (.in(n10663), .out(n10663_0));
mux13 mux_5498 (.in({n14237_1/**/, n14213_0, n14206_0, n14199_0, n14192_0, n14166_0, n14108_0, n14103_0, n10580_1, n7711, n7699, n7611, n7603}), .out(n10664), .config_in(config_chain[18027:18022]), .config_rst(config_rst)); 
buffer_wire buffer_10664 (.in(n10664), .out(n10664_0));
mux3 mux_5499 (.in({n14721_0, n14720_0, n8681}), .out(n10665), .config_in(config_chain[18029:18028]), .config_rst(config_rst)); 
buffer_wire buffer_10665 (.in(n10665), .out(n10665_0));
mux13 mux_5500 (.in({n14239_1, n14221_0, n14214_0, n14200_0, n14185_0, n14135_0, n14110_0, n14100_0, n10582_1, n7711, n7703, n7611/**/, n7603}), .out(n10666), .config_in(config_chain[18035:18030]), .config_rst(config_rst)); 
buffer_wire buffer_10666 (.in(n10666), .out(n10666_0));
mux3 mux_5501 (.in({n14723_0, n14722_0, n8681/**/}), .out(n10667), .config_in(config_chain[18037:18036]), .config_rst(config_rst)); 
buffer_wire buffer_10667 (.in(n10667), .out(n10667_0));
mux13 mux_5502 (.in({n14241_1, n14222_0, n14207_0, n14193_0, n14186_0, n14167_0, n14142_0, n14092_0/**/, n10584_1, n7711, n7703, n7615, n7603}), .out(n10668), .config_in(config_chain[18043:18038]), .config_rst(config_rst)); 
buffer_wire buffer_10668 (.in(n10668), .out(n10668_0));
mux3 mux_5503 (.in({n14725_0, n14724_0, n8685}), .out(n10669), .config_in(config_chain[18045:18044]), .config_rst(config_rst)); 
buffer_wire buffer_10669 (.in(n10669), .out(n10669_0));
mux13 mux_5504 (.in({n14243_1, n14215_0, n14208_0, n14201_1, n14194_0, n14174_0, n14172_0, n14111_0, n10518_2, n7711/**/, n7703, n7615, n7607}), .out(n10670), .config_in(config_chain[18051:18046]), .config_rst(config_rst)); 
buffer_wire buffer_10670 (.in(n10670), .out(n10670_0));
mux3 mux_5505 (.in({n14727_1, n14726_0, n8689}), .out(n10671), .config_in(config_chain[18053:18052]), .config_rst(config_rst)); 
buffer_wire buffer_10671 (.in(n10671), .out(n10671_0));
mux15 mux_5506 (.in({n14509_1, n14479_0, n14472_0, n14465_1, n14458_0, n14440_0, n14430_0, n14377_0, n14352_0, n10586_1, n8689, n8681, n8593, n8585, n8577}), .out(n10672), .config_in(config_chain[18059:18054]), .config_rst(config_rst)); 
buffer_wire buffer_10672 (.in(n10672), .out(n10672_0));
mux4 mux_5507 (.in({n14729_0, n14728_0, n8693, n8577}), .out(n10673), .config_in(config_chain[18061:18060]), .config_rst(config_rst)); 
buffer_wire buffer_10673 (.in(n10673), .out(n10673_0));
mux15 mux_5508 (.in({n14489_1, n14487_1, n14480_0, n14451_0, n14444_0, n14442_0, n14422_0, n14409_0/**/, n14384_0, n10588_1, n8693, n8681, n8593, n8585, n8577}), .out(n10674), .config_in(config_chain[18067:18062]), .config_rst(config_rst)); 
buffer_wire buffer_10674 (.in(n10674), .out(n10674_0));
mux3 mux_5509 (.in({n14731_0, n14730_0, n8581}), .out(n10675), .config_in(config_chain[18069:18068]), .config_rst(config_rst)); 
buffer_wire buffer_10675 (.in(n10675), .out(n10675_0));
mux15 mux_5510 (.in({n14491_1, n14473_0, n14466_0, n14459_0/**/, n14452_0, n14441_0, n14416_0, n14414_0, n14353_0, n10590_1, n8693, n8685, n8593, n8585, n8577}), .out(n10676), .config_in(config_chain[18075:18070]), .config_rst(config_rst)); 
buffer_wire buffer_10676 (.in(n10676), .out(n10676_0));
mux3 mux_5511 (.in({n14733_0, n14732_0, n8585}), .out(n10677), .config_in(config_chain[18077:18076]), .config_rst(config_rst)); 
buffer_wire buffer_10677 (.in(n10677), .out(n10677_0));
mux15 mux_5512 (.in({n14493_1, n14481_0, n14474_0, n14460_0, n14445_0, n14443_0, n14406_0, n14385_0/**/, n14360_0, n10592_1, n8693, n8685, n8677, n8585, n8577}), .out(n10678), .config_in(config_chain[18083:18078]), .config_rst(config_rst)); 
buffer_wire buffer_10678 (.in(n10678), .out(n10678_0));
mux3 mux_5513 (.in({n14735_0, n14734_0, n8589}), .out(n10679), .config_in(config_chain[18085:18084]), .config_rst(config_rst)); 
buffer_wire buffer_10679 (.in(n10679), .out(n10679_0));
mux14 mux_5514 (.in({n14495_1, n14482_0, n14467_0, n14453_0, n14446_0/**/, n14417_0, n14398_0, n14392_0, n10594_1, n8693, n8685, n8677, n8589, n8577}), .out(n10680), .config_in(config_chain[18091:18086]), .config_rst(config_rst)); 
buffer_wire buffer_10680 (.in(n10680), .out(n10680_0));
mux3 mux_5515 (.in({n14737_0, n14736_0, n8589}), .out(n10681), .config_in(config_chain[18093:18092]), .config_rst(config_rst)); 
buffer_wire buffer_10681 (.in(n10681), .out(n10681_0));
mux14 mux_5516 (.in({n14497_1, n14475_0/**/, n14468_0, n14461_0, n14454_0, n14424_0, n14390_0, n14361_0, n10596_1, n8693, n8685, n8677, n8589, n8581}), .out(n10682), .config_in(config_chain[18099:18094]), .config_rst(config_rst)); 
buffer_wire buffer_10682 (.in(n10682), .out(n10682_0));
mux3 mux_5517 (.in({n14739_0, n14738_0, n8593}), .out(n10683), .config_in(config_chain[18101:18100]), .config_rst(config_rst)); 
buffer_wire buffer_10683 (.in(n10683), .out(n10683_0));
mux13 mux_5518 (.in({n14499_1/**/, n14483_0, n14476_0, n14462_0, n14447_0, n14393_0, n14382_0, n14368_0, n10598_1, n8685, n8677, n8589, n8581}), .out(n10684), .config_in(config_chain[18107:18102]), .config_rst(config_rst)); 
buffer_wire buffer_10684 (.in(n10684), .out(n10684_0));
mux3 mux_5519 (.in({n14741_0/**/, n14740_0, n8677}), .out(n10685), .config_in(config_chain[18109:18108]), .config_rst(config_rst)); 
buffer_wire buffer_10685 (.in(n10685), .out(n10685_0));
mux13 mux_5520 (.in({n14501_1, n14484_0, n14469_0, n14455_0, n14448_0, n14425_0, n14400_0, n14374_0, n10600_1, n8689, n8677, n8589, n8581}), .out(n10686), .config_in(config_chain[18115:18110]), .config_rst(config_rst)); 
buffer_wire buffer_10686 (.in(n10686), .out(n10686_0));
mux3 mux_5521 (.in({n14743_0, n14742_0, n8681}), .out(n10687), .config_in(config_chain[18117:18116]), .config_rst(config_rst)); 
buffer_wire buffer_10687 (.in(n10687), .out(n10687_0));
mux13 mux_5522 (.in({n14503_1, n14477_0, n14470_0, n14463_0, n14456_0, n14432_0, n14369_0, n14366_0, n10602_1, n8689, n8681/**/, n8589, n8581}), .out(n10688), .config_in(config_chain[18123:18118]), .config_rst(config_rst)); 
buffer_wire buffer_10688 (.in(n10688), .out(n10688_0));
mux3 mux_5523 (.in({n14745_0, n14744_0, n8685}), .out(n10689), .config_in(config_chain[18125:18124]), .config_rst(config_rst)); 
buffer_wire buffer_10689 (.in(n10689), .out(n10689_0));
mux13 mux_5524 (.in({n14505_1, n14485_0, n14478_0, n14464_0, n14449_0, n14401_0, n14376_0/**/, n14358_0, n10604_1, n8689, n8681, n8593, n8581}), .out(n10690), .config_in(config_chain[18131:18126]), .config_rst(config_rst)); 
buffer_wire buffer_10690 (.in(n10690), .out(n10690_0));
mux3 mux_5525 (.in({n14747_0, n14746_0, n8685/**/}), .out(n10691), .config_in(config_chain[18133:18132]), .config_rst(config_rst)); 
buffer_wire buffer_10691 (.in(n10691), .out(n10691_0));
mux13 mux_5526 (.in({n14507_1, n14486_0, n14471_0, n14457_0, n14450_0, n14438_0, n14433_1, n14408_0/**/, n10520_2, n8689, n8681, n8593, n8585}), .out(n10692), .config_in(config_chain[18139:18134]), .config_rst(config_rst)); 
buffer_wire buffer_10692 (.in(n10692), .out(n10692_0));
mux3 mux_5527 (.in({n14749_1/**/, n14748_0, n8689}), .out(n10693), .config_in(config_chain[18141:18140]), .config_rst(config_rst)); 
buffer_wire buffer_10693 (.in(n10693), .out(n10693_0));
mux4 mux_5528 (.in({n12423_1, n12270_1, n967, n851}), .out(n10694), .config_in(config_chain[18143:18142]), .config_rst(config_rst)); 
buffer_wire buffer_10694 (.in(n10694), .out(n10694_0));
mux15 mux_5529 (.in({n13451_1, n13442_0, n13437_0, n13425_0, n13396_0/**/, n13391_0, n13387_1, n13382_1, n13378_1, n10847_1, n3897, n3889, n3801, n3793, n3785}), .out(n10695), .config_in(config_chain[18149:18144]), .config_rst(config_rst)); 
buffer_wire buffer_10695 (.in(n10695), .out(n10695_0));
mux4 mux_5530 (.in({n12363_0, n12362_0, n967, n851}), .out(n10696), .config_in(config_chain[18151:18150]), .config_rst(config_rst)); 
buffer_wire buffer_10696 (.in(n10696), .out(n10696_0));
mux16 mux_5531 (.in({n12677_1, n12672_0, n12657_0, n12649_0, n12644_0, n12623_0, n12618_0, n12612_1, n12605_0, n12598_1/**/, n10787_1, n963, n955, n867, n859, n851}), .out(n10697), .config_in(config_chain[18157:18152]), .config_rst(config_rst)); 
buffer_wire buffer_10697 (.in(n10697), .out(n10697_0));
mux4 mux_5532 (.in({n12383_0, n12382_0, n967, n851}), .out(n10698), .config_in(config_chain[18159:18158]), .config_rst(config_rst)); 
buffer_wire buffer_10698 (.in(n10698), .out(n10698_0));
mux16 mux_5533 (.in({n12933_1, n12919_0, n12914_0, n12908_0, n12893_0, n12885_0, n12880_0, n12868_1, n12861_0, n12856_1, n10807_1, n1941, n1933, n1845, n1837, n1829}), .out(n10699), .config_in(config_chain[18165:18160]), .config_rst(config_rst)); 
buffer_wire buffer_10699 (.in(n10699), .out(n10699_0));
mux4 mux_5534 (.in({n12403_0, n12402_0, n967, n851}), .out(n10700), .config_in(config_chain[18167:18166]), .config_rst(config_rst)); 
buffer_wire buffer_10700 (.in(n10700), .out(n10700_0));
mux16 mux_5535 (.in({n13191_1, n13183_0, n13178_0, n13157_0, n13152_0, n13146_0/**/, n13131_0, n13126_1, n13119_0, n13116_1, n10827_1, n2919, n2911, n2823, n2815, n2807}), .out(n10701), .config_in(config_chain[18173:18168]), .config_rst(config_rst)); 
buffer_wire buffer_10701 (.in(n10701), .out(n10701_0));
mux3 mux_5536 (.in({n12425_1/**/, n12278_1, n851}), .out(n10702), .config_in(config_chain[18175:18174]), .config_rst(config_rst)); 
buffer_wire buffer_10702 (.in(n10702), .out(n10702_0));
mux15 mux_5537 (.in({n13471_1, n13445_0, n13416_0, n13411_0, n13404_0, n13399_0, n13389_1, n13384_1, n13298_1, n10849_1, n3901, n3889, n3801, n3793, n3785}), .out(n10703), .config_in(config_chain[18181:18176]), .config_rst(config_rst)); 
buffer_wire buffer_10703 (.in(n10703), .out(n10703_0));
mux3 mux_5538 (.in({n12365_0/**/, n12364_0, n855}), .out(n10704), .config_in(config_chain[18183:18182]), .config_rst(config_rst)); 
buffer_wire buffer_10704 (.in(n10704), .out(n10704_0));
mux16 mux_5539 (.in({n12695_1, n12671_0, n12666_0, n12643_0, n12638_0, n12632_0, n12617_0/**/, n12614_1, n12607_1, n12526_1, n10789_1, n963, n955, n867, n859, n851}), .out(n10705), .config_in(config_chain[18189:18184]), .config_rst(config_rst)); 
buffer_wire buffer_10705 (.in(n10705), .out(n10705_0));
mux3 mux_5540 (.in({n12385_0, n12384_0, n855}), .out(n10706), .config_in(config_chain[18191:18190]), .config_rst(config_rst)); 
buffer_wire buffer_10706 (.in(n10706), .out(n10706_0));
mux16 mux_5541 (.in({n12951_1, n12928_0, n12913_0, n12907_0, n12902_0, n12879_0, n12874_0, n12870_1, n12863_0, n12784_1, n10809_1, n1941, n1933, n1845/**/, n1837, n1829}), .out(n10707), .config_in(config_chain[18197:18192]), .config_rst(config_rst)); 
buffer_wire buffer_10707 (.in(n10707), .out(n10707_0));
mux3 mux_5542 (.in({n12405_0, n12404_0, n855/**/}), .out(n10708), .config_in(config_chain[18199:18198]), .config_rst(config_rst)); 
buffer_wire buffer_10708 (.in(n10708), .out(n10708_0));
mux16 mux_5543 (.in({n13209_1, n13177_0, n13172_0, n13166_0, n13151_0, n13145_0, n13140_0, n13128_1, n13121_0, n13044_1, n10829_1, n2919/**/, n2911, n2823, n2815, n2807}), .out(n10709), .config_in(config_chain[18205:18200]), .config_rst(config_rst)); 
buffer_wire buffer_10709 (.in(n10709), .out(n10709_0));
mux3 mux_5544 (.in({n12427_1, n12286_1/**/, n855}), .out(n10710), .config_in(config_chain[18207:18206]), .config_rst(config_rst)); 
buffer_wire buffer_10710 (.in(n10710), .out(n10710_0));
mux15 mux_5545 (.in({n13469_1, n13436_0, n13431_0, n13424_0, n13419_0, n13407_0, n13390_0, n13386_1, n13306_1, n10851_1/**/, n3901, n3893, n3801, n3793, n3785}), .out(n10711), .config_in(config_chain[18213:18208]), .config_rst(config_rst)); 
buffer_wire buffer_10711 (.in(n10711), .out(n10711_0));
mux3 mux_5546 (.in({n12367_0, n12366_0, n855}), .out(n10712), .config_in(config_chain[18215:18214]), .config_rst(config_rst)); 
buffer_wire buffer_10712 (.in(n10712), .out(n10712_0));
mux15 mux_5547 (.in({n12693_1, n12665_0, n12660_0, n12652_0, n12637_0, n12631_0, n12626_0, n12609_1, n12534_1, n10791_1, n963, n955, n867, n859, n851}), .out(n10713), .config_in(config_chain[18221:18216]), .config_rst(config_rst)); 
buffer_wire buffer_10713 (.in(n10713), .out(n10713_0));
mux3 mux_5548 (.in({n12387_0, n12386_0/**/, n859}), .out(n10714), .config_in(config_chain[18223:18222]), .config_rst(config_rst)); 
buffer_wire buffer_10714 (.in(n10714), .out(n10714_0));
mux15 mux_5549 (.in({n12949_1, n12927_0, n12922_0, n12901_0, n12896_0, n12888_0, n12873_0, n12865_1, n12792_1, n10811_1, n1941, n1933, n1845, n1837, n1829}), .out(n10715), .config_in(config_chain[18229:18224]), .config_rst(config_rst)); 
buffer_wire buffer_10715 (.in(n10715), .out(n10715_0));
mux3 mux_5550 (.in({n12407_0, n12406_0, n859}), .out(n10716), .config_in(config_chain[18231:18230]), .config_rst(config_rst)); 
buffer_wire buffer_10716 (.in(n10716), .out(n10716_0));
mux15 mux_5551 (.in({n13207_1, n13186_0, n13171_0, n13165_0, n13160_0, n13139_0/**/, n13134_0, n13123_0, n13052_1, n10831_1, n2919, n2911, n2823, n2815, n2807}), .out(n10717), .config_in(config_chain[18237:18232]), .config_rst(config_rst)); 
buffer_wire buffer_10717 (.in(n10717), .out(n10717_0));
mux3 mux_5552 (.in({n12429_1/**/, n12294_1, n859}), .out(n10718), .config_in(config_chain[18239:18238]), .config_rst(config_rst)); 
buffer_wire buffer_10718 (.in(n10718), .out(n10718_0));
mux15 mux_5553 (.in({n13467_1, n13444_0, n13439_0, n13427_0, n13410_0, n13398_0, n13393_0, n13388_1, n13314_1, n10853_1/**/, n3901, n3893, n3885, n3793, n3785}), .out(n10719), .config_in(config_chain[18245:18240]), .config_rst(config_rst)); 
buffer_wire buffer_10719 (.in(n10719), .out(n10719_0));
mux3 mux_5554 (.in({n12369_0, n12368_0, n859}), .out(n10720), .config_in(config_chain[18247:18246]), .config_rst(config_rst)); 
buffer_wire buffer_10720 (.in(n10720), .out(n10720_0));
mux15 mux_5555 (.in({n12691_1, n12674_0, n12659_0, n12651_0, n12646_0, n12625_0, n12620_0, n12611_1, n12542_1/**/, n10793_1, n963, n955, n867, n859, n851}), .out(n10721), .config_in(config_chain[18253:18248]), .config_rst(config_rst)); 
buffer_wire buffer_10721 (.in(n10721), .out(n10721_0));
mux3 mux_5556 (.in({n12389_0, n12388_0/**/, n859}), .out(n10722), .config_in(config_chain[18255:18254]), .config_rst(config_rst)); 
buffer_wire buffer_10722 (.in(n10722), .out(n10722_0));
mux15 mux_5557 (.in({n12947_1/**/, n12921_0, n12916_0, n12910_0, n12895_0, n12887_0, n12882_0, n12867_1, n12800_1, n10813_1, n1941, n1933, n1845, n1837, n1829}), .out(n10723), .config_in(config_chain[18261:18256]), .config_rst(config_rst)); 
buffer_wire buffer_10723 (.in(n10723), .out(n10723_0));
mux3 mux_5558 (.in({n12409_0, n12408_0, n863}), .out(n10724), .config_in(config_chain[18263:18262]), .config_rst(config_rst)); 
buffer_wire buffer_10724 (.in(n10724), .out(n10724_0));
mux15 mux_5559 (.in({n13205_1, n13185_0/**/, n13180_0, n13159_0, n13154_0, n13148_0, n13133_0, n13125_1, n13060_1, n10833_1, n2919, n2911, n2823, n2815, n2807}), .out(n10725), .config_in(config_chain[18269:18264]), .config_rst(config_rst)); 
buffer_wire buffer_10725 (.in(n10725), .out(n10725_0));
mux3 mux_5560 (.in({n12431_1, n12302_1/**/, n863}), .out(n10726), .config_in(config_chain[18271:18270]), .config_rst(config_rst)); 
buffer_wire buffer_10726 (.in(n10726), .out(n10726_0));
mux14 mux_5561 (.in({n13465_1, n13447_0, n13430_0, n13418_0, n13413_0, n13406_0, n13401_0, n13322_1, n10855_1, n3901, n3893, n3885, n3797, n3785}), .out(n10727), .config_in(config_chain[18277:18272]), .config_rst(config_rst)); 
buffer_wire buffer_10727 (.in(n10727), .out(n10727_0));
mux3 mux_5562 (.in({n12371_0/**/, n12370_0, n863}), .out(n10728), .config_in(config_chain[18279:18278]), .config_rst(config_rst)); 
buffer_wire buffer_10728 (.in(n10728), .out(n10728_0));
mux15 mux_5563 (.in({n12689_1, n12673_0, n12668_0, n12645_0, n12640_0, n12634_0, n12619_0, n12613_1, n12550_1, n10795_1, n963, n955, n867, n859, n851}), .out(n10729), .config_in(config_chain[18285:18280]), .config_rst(config_rst)); 
buffer_wire buffer_10729 (.in(n10729), .out(n10729_0));
mux3 mux_5564 (.in({n12391_0, n12390_0, n863}), .out(n10730), .config_in(config_chain[18287:18286]), .config_rst(config_rst)); 
buffer_wire buffer_10730 (.in(n10730), .out(n10730_0));
mux15 mux_5565 (.in({n12945_1, n12930_0, n12915_0, n12909_0, n12904_0, n12881_0, n12876_0/**/, n12869_1, n12808_1, n10815_1, n1941, n1933, n1845, n1837, n1829}), .out(n10731), .config_in(config_chain[18293:18288]), .config_rst(config_rst)); 
buffer_wire buffer_10731 (.in(n10731), .out(n10731_0));
mux3 mux_5566 (.in({n12411_0, n12410_0, n863}), .out(n10732), .config_in(config_chain[18295:18294]), .config_rst(config_rst)); 
buffer_wire buffer_10732 (.in(n10732), .out(n10732_0));
mux15 mux_5567 (.in({n13203_1, n13179_0, n13174_0, n13168_0, n13153_0, n13147_0, n13142_0, n13127_1, n13068_1, n10835_1, n2919, n2911, n2823, n2815, n2807}), .out(n10733), .config_in(config_chain[18301:18296]), .config_rst(config_rst)); 
buffer_wire buffer_10733 (.in(n10733), .out(n10733_0));
mux3 mux_5568 (.in({n12433_1, n12310_1/**/, n867}), .out(n10734), .config_in(config_chain[18303:18302]), .config_rst(config_rst)); 
buffer_wire buffer_10734 (.in(n10734), .out(n10734_0));
mux14 mux_5569 (.in({n13463_1, n13438_0, n13433_0, n13426_0, n13421_0, n13409_0, n13392_0, n13330_1, n10857_1, n3901, n3893, n3885, n3797/**/, n3789}), .out(n10735), .config_in(config_chain[18309:18304]), .config_rst(config_rst)); 
buffer_wire buffer_10735 (.in(n10735), .out(n10735_0));
mux3 mux_5570 (.in({n12373_0, n12372_0, n867}), .out(n10736), .config_in(config_chain[18311:18310]), .config_rst(config_rst)); 
buffer_wire buffer_10736 (.in(n10736), .out(n10736_0));
mux15 mux_5571 (.in({n12687_1, n12667_0, n12662_0, n12654_0, n12639_0, n12633_0, n12628_0, n12615_1, n12558_1, n10797_1, n967, n959, n951, n863, n855}), .out(n10737), .config_in(config_chain[18317:18312]), .config_rst(config_rst)); 
buffer_wire buffer_10737 (.in(n10737), .out(n10737_0));
mux3 mux_5572 (.in({n12393_0/**/, n12392_0, n867}), .out(n10738), .config_in(config_chain[18319:18318]), .config_rst(config_rst)); 
buffer_wire buffer_10738 (.in(n10738), .out(n10738_0));
mux15 mux_5573 (.in({n12943_1/**/, n12929_0, n12924_0, n12903_0, n12898_0, n12890_0, n12875_0, n12871_1, n12816_1, n10817_1, n1945, n1937, n1929, n1841, n1833}), .out(n10739), .config_in(config_chain[18325:18320]), .config_rst(config_rst)); 
buffer_wire buffer_10739 (.in(n10739), .out(n10739_0));
mux3 mux_5574 (.in({n12413_0, n12412_0/**/, n867}), .out(n10740), .config_in(config_chain[18327:18326]), .config_rst(config_rst)); 
buffer_wire buffer_10740 (.in(n10740), .out(n10740_0));
mux15 mux_5575 (.in({n13201_1, n13188_0/**/, n13173_0, n13167_0, n13162_0, n13141_0, n13136_0, n13129_1, n13076_1, n10837_1, n2923, n2915, n2907, n2819, n2811}), .out(n10741), .config_in(config_chain[18333:18328]), .config_rst(config_rst)); 
buffer_wire buffer_10741 (.in(n10741), .out(n10741_0));
mux3 mux_5576 (.in({n12435_1, n12318_1/**/, n867}), .out(n10742), .config_in(config_chain[18335:18334]), .config_rst(config_rst)); 
buffer_wire buffer_10742 (.in(n10742), .out(n10742_0));
mux13 mux_5577 (.in({n13461_1, n13446_0, n13441_0, n13429_0, n13412_0, n13400_0, n13395_0, n13338_1, n10859_1/**/, n3893, n3885, n3797, n3789}), .out(n10743), .config_in(config_chain[18341:18336]), .config_rst(config_rst)); 
buffer_wire buffer_10743 (.in(n10743), .out(n10743_0));
mux3 mux_5578 (.in({n12375_0/**/, n12374_0, n951}), .out(n10744), .config_in(config_chain[18343:18342]), .config_rst(config_rst)); 
buffer_wire buffer_10744 (.in(n10744), .out(n10744_0));
mux15 mux_5579 (.in({n12685_1, n12661_0, n12656_0, n12653_0, n12648_0, n12627_0, n12622_0, n12604_1, n12566_1/**/, n10799_1, n967, n959, n951, n863, n855}), .out(n10745), .config_in(config_chain[18349:18344]), .config_rst(config_rst)); 
buffer_wire buffer_10745 (.in(n10745), .out(n10745_0));
mux3 mux_5580 (.in({n12395_0, n12394_0/**/, n951}), .out(n10746), .config_in(config_chain[18351:18350]), .config_rst(config_rst)); 
buffer_wire buffer_10746 (.in(n10746), .out(n10746_0));
mux15 mux_5581 (.in({n12941_1, n12923_0, n12918_0, n12897_0, n12892_0, n12889_0, n12884_0/**/, n12860_1, n12824_1, n10819_1, n1945, n1937, n1929, n1841, n1833}), .out(n10747), .config_in(config_chain[18357:18352]), .config_rst(config_rst)); 
buffer_wire buffer_10747 (.in(n10747), .out(n10747_0));
mux3 mux_5582 (.in({n12415_0, n12414_0/**/, n951}), .out(n10748), .config_in(config_chain[18359:18358]), .config_rst(config_rst)); 
buffer_wire buffer_10748 (.in(n10748), .out(n10748_0));
mux15 mux_5583 (.in({n13199_1, n13187_0, n13182_0, n13161_0, n13156_0, n13135_0/**/, n13130_0, n13118_1, n13084_1, n10839_1, n2923, n2915, n2907, n2819, n2811}), .out(n10749), .config_in(config_chain[18365:18360]), .config_rst(config_rst)); 
buffer_wire buffer_10749 (.in(n10749), .out(n10749_0));
mux3 mux_5584 (.in({n12437_1, n12326_1, n951/**/}), .out(n10750), .config_in(config_chain[18367:18366]), .config_rst(config_rst)); 
buffer_wire buffer_10750 (.in(n10750), .out(n10750_0));
mux13 mux_5585 (.in({n13459_1, n13449_0, n13432_0, n13420_0/**/, n13415_0, n13408_0, n13403_0, n13346_1, n10861_1, n3897, n3885, n3797, n3789}), .out(n10751), .config_in(config_chain[18373:18368]), .config_rst(config_rst)); 
buffer_wire buffer_10751 (.in(n10751), .out(n10751_0));
mux3 mux_5586 (.in({n12377_0, n12376_0, n951}), .out(n10752), .config_in(config_chain[18375:18374]), .config_rst(config_rst)); 
buffer_wire buffer_10752 (.in(n10752), .out(n10752_0));
mux15 mux_5587 (.in({n12683_1, n12675_0, n12670_0, n12647_0, n12642_0, n12621_0, n12616_0, n12606_1, n12574_1, n10801_1, n967, n959, n951, n863, n855}), .out(n10753), .config_in(config_chain[18381:18376]), .config_rst(config_rst)); 
buffer_wire buffer_10753 (.in(n10753), .out(n10753_0));
mux3 mux_5588 (.in({n12397_0, n12396_0, n955}), .out(n10754), .config_in(config_chain[18383:18382]), .config_rst(config_rst)); 
buffer_wire buffer_10754 (.in(n10754), .out(n10754_0));
mux15 mux_5589 (.in({n12939_1, n12917_0, n12912_0, n12911_0, n12906_0, n12883_0, n12878_0, n12862_1, n12832_1, n10821_1, n1945, n1937, n1929, n1841/**/, n1833}), .out(n10755), .config_in(config_chain[18389:18384]), .config_rst(config_rst)); 
buffer_wire buffer_10755 (.in(n10755), .out(n10755_0));
mux3 mux_5590 (.in({n12417_0, n12416_0, n955}), .out(n10756), .config_in(config_chain[18391:18390]), .config_rst(config_rst)); 
buffer_wire buffer_10756 (.in(n10756), .out(n10756_0));
mux15 mux_5591 (.in({n13197_1, n13181_0, n13176_0/**/, n13155_0, n13150_0, n13149_0, n13144_0, n13120_1, n13092_1, n10841_1, n2923, n2915, n2907, n2819, n2811}), .out(n10757), .config_in(config_chain[18397:18392]), .config_rst(config_rst)); 
buffer_wire buffer_10757 (.in(n10757), .out(n10757_0));
mux3 mux_5592 (.in({n12439_1, n12334_1/**/, n955}), .out(n10758), .config_in(config_chain[18399:18398]), .config_rst(config_rst)); 
buffer_wire buffer_10758 (.in(n10758), .out(n10758_0));
mux13 mux_5593 (.in({n13457_1, n13440_0, n13435_0, n13428_0, n13423_0, n13394_0, n13381_0, n13354_1, n10863_1, n3897, n3889, n3797, n3789}), .out(n10759), .config_in(config_chain[18405:18400]), .config_rst(config_rst)); 
buffer_wire buffer_10759 (.in(n10759), .out(n10759_0));
mux3 mux_5594 (.in({n12379_0/**/, n12378_0, n955}), .out(n10760), .config_in(config_chain[18407:18406]), .config_rst(config_rst)); 
buffer_wire buffer_10760 (.in(n10760), .out(n10760_0));
mux15 mux_5595 (.in({n12681_1, n12669_0, n12664_0, n12641_0, n12636_0, n12635_0, n12630_0, n12608_1, n12582_1, n10803_1, n967, n959, n951, n863, n855}), .out(n10761), .config_in(config_chain[18413:18408]), .config_rst(config_rst)); 
buffer_wire buffer_10761 (.in(n10761), .out(n10761_0));
mux3 mux_5596 (.in({n12399_0, n12398_0, n955}), .out(n10762), .config_in(config_chain[18415:18414]), .config_rst(config_rst)); 
buffer_wire buffer_10762 (.in(n10762), .out(n10762_0));
mux15 mux_5597 (.in({n12937_1, n12931_0, n12926_0, n12905_0, n12900_0, n12877_0, n12872_0, n12864_1, n12840_1, n10823_1/**/, n1945, n1937, n1929, n1841, n1833}), .out(n10763), .config_in(config_chain[18421:18416]), .config_rst(config_rst)); 
buffer_wire buffer_10763 (.in(n10763), .out(n10763_0));
mux3 mux_5598 (.in({n12419_0, n12418_0/**/, n959}), .out(n10764), .config_in(config_chain[18423:18422]), .config_rst(config_rst)); 
buffer_wire buffer_10764 (.in(n10764), .out(n10764_0));
mux15 mux_5599 (.in({n13195_1, n13175_0, n13170_0, n13169_0, n13164_0, n13143_0, n13138_0, n13122_1, n13100_1, n10843_1, n2923, n2915, n2907, n2819, n2811}), .out(n10765), .config_in(config_chain[18429:18424]), .config_rst(config_rst)); 
buffer_wire buffer_10765 (.in(n10765), .out(n10765_0));
mux3 mux_5600 (.in({n12441_1, n12342_1, n959/**/}), .out(n10766), .config_in(config_chain[18431:18430]), .config_rst(config_rst)); 
buffer_wire buffer_10766 (.in(n10766), .out(n10766_0));
mux13 mux_5601 (.in({n13455_1, n13448_0, n13443_0, n13414_0, n13402_0, n13397_0, n13383_0, n13362_1, n10865_1/**/, n3897, n3889, n3801, n3789}), .out(n10767), .config_in(config_chain[18437:18432]), .config_rst(config_rst)); 
buffer_wire buffer_10767 (.in(n10767), .out(n10767_0));
mux3 mux_5602 (.in({n12381_0, n12380_0, n959/**/}), .out(n10768), .config_in(config_chain[18439:18438]), .config_rst(config_rst)); 
buffer_wire buffer_10768 (.in(n10768), .out(n10768_0));
mux15 mux_5603 (.in({n12679_1, n12663_0, n12658_0, n12655_0, n12650_0, n12629_0, n12624_0, n12610_1, n12590_1, n10805_1, n967, n959, n951, n863, n855}), .out(n10769), .config_in(config_chain[18445:18440]), .config_rst(config_rst)); 
buffer_wire buffer_10769 (.in(n10769), .out(n10769_0));
mux3 mux_5604 (.in({n12401_0, n12400_0, n959}), .out(n10770), .config_in(config_chain[18447:18446]), .config_rst(config_rst)); 
buffer_wire buffer_10770 (.in(n10770), .out(n10770_0));
mux15 mux_5605 (.in({n12935_1, n12925_0, n12920_0, n12899_0, n12894_0, n12891_0, n12886_0, n12866_1, n12848_1, n10825_1, n1945, n1937/**/, n1929, n1841, n1833}), .out(n10771), .config_in(config_chain[18453:18448]), .config_rst(config_rst)); 
buffer_wire buffer_10771 (.in(n10771), .out(n10771_0));
mux3 mux_5606 (.in({n12421_0, n12420_0, n959}), .out(n10772), .config_in(config_chain[18455:18454]), .config_rst(config_rst)); 
buffer_wire buffer_10772 (.in(n10772), .out(n10772_0));
mux15 mux_5607 (.in({n13193_1, n13189_0, n13184_0, n13163_0, n13158_0, n13137_0, n13132_0, n13124_1, n13108_1, n10845_1, n2923, n2915, n2907, n2819/**/, n2811}), .out(n10773), .config_in(config_chain[18461:18456]), .config_rst(config_rst)); 
buffer_wire buffer_10773 (.in(n10773), .out(n10773_0));
mux3 mux_5608 (.in({n12351_1, n12350_1, n963}), .out(n10774), .config_in(config_chain[18463:18462]), .config_rst(config_rst)); 
buffer_wire buffer_10774 (.in(n10774), .out(n10774_0));
mux13 mux_5609 (.in({n13453_1, n13434_0, n13422_0, n13417_0, n13405_0, n13385_0, n13380_1, n13370_1, n10867_1, n3897, n3889, n3801, n3793}), .out(n10775), .config_in(config_chain[18469:18464]), .config_rst(config_rst)); 
buffer_wire buffer_10775 (.in(n10775), .out(n10775_0));
mux3 mux_5610 (.in({n12353_1, n12352_1, n963}), .out(n10776), .config_in(config_chain[18471:18470]), .config_rst(config_rst)); 
buffer_wire buffer_10776 (.in(n10776), .out(n10776_0));
mux13 mux_5611 (.in({n13717_1/**/, n13712_0, n13707_0, n13676_0, n13664_0, n13659_0, n13647_0, n13634_1, n10889_1, n4875, n4867, n4779, n4771}), .out(n10777), .config_in(config_chain[18477:18472]), .config_rst(config_rst)); 
buffer_wire buffer_10777 (.in(n10777), .out(n10777_0));
mux3 mux_5612 (.in({n12355_1, n12354_1, n963}), .out(n10778), .config_in(config_chain[18479:18478]), .config_rst(config_rst)); 
buffer_wire buffer_10778 (.in(n10778), .out(n10778_0));
mux13 mux_5613 (.in({n13983_1, n13970_0/**/, n13965_0, n13956_0, n13951_0, n13920_0, n13911_0, n13900_1, n10911_0, n5853, n5845, n5757, n5749}), .out(n10779), .config_in(config_chain[18485:18480]), .config_rst(config_rst)); 
buffer_wire buffer_10779 (.in(n10779), .out(n10779_0));
mux3 mux_5614 (.in({n12357_1, n12356_1, n963}), .out(n10780), .config_in(config_chain[18487:18486]), .config_rst(config_rst)); 
buffer_wire buffer_10780 (.in(n10780), .out(n10780_0));
mux13 mux_5615 (.in({n14249_1, n14245_1, n14228_0, n14214_0, n14209_0, n14200_0, n14195_0/**/, n14166_1, n10933_0, n6831, n6823, n6735, n6727}), .out(n10781), .config_in(config_chain[18493:18488]), .config_rst(config_rst)); 
buffer_wire buffer_10781 (.in(n10781), .out(n10781_0));
mux3 mux_5616 (.in({n12359_1/**/, n12358_1, n963}), .out(n10782), .config_in(config_chain[18495:18494]), .config_rst(config_rst)); 
buffer_wire buffer_10782 (.in(n10782), .out(n10782_0));
mux13 mux_5617 (.in({n14513_1/**/, n14492_0, n14487_1, n14478_0, n14473_0, n14459_0, n14432_1, n14424_1, n10955_0, n7809, n7801, n7713, n7705}), .out(n10783), .config_in(config_chain[18501:18496]), .config_rst(config_rst)); 
buffer_wire buffer_10783 (.in(n10783), .out(n10783_0));
mux3 mux_5618 (.in({n12361_1, n12360_1, n967}), .out(n10784), .config_in(config_chain[18503:18502]), .config_rst(config_rst)); 
buffer_wire buffer_10784 (.in(n10784), .out(n10784_0));
mux3 mux_5619 (.in({n14793_1/**/, n14704_1, n8791}), .out(n10785), .config_in(config_chain[18505:18504]), .config_rst(config_rst)); 
buffer_wire buffer_10785 (.in(n10785), .out(n10785_0));
mux16 mux_5620 (.in({n12695_1, n12673_0, n12656_0, n12648_0, n12645_0, n12622_0, n12619_0, n12613_1, n12604_1, n12590_1, n10696_0, n1941, n1933/**/, n1845, n1837, n1829}), .out(n10786), .config_in(config_chain[18511:18506]), .config_rst(config_rst)); 
buffer_wire buffer_10786 (.in(n10786), .out(n10786_0));
mux15 mux_5621 (.in({n13715_1, n13698_0, n13693_0, n13684_0, n13679_0, n13667_0, n13649_0, n13644_1, n13642_1, n10869_1, n4875, n4867, n4779, n4771, n4763}), .out(n10787), .config_in(config_chain[18517:18512]), .config_rst(config_rst)); 
buffer_wire buffer_10787 (.in(n10787), .out(n10787_0));
mux16 mux_5622 (.in({n12677_1, n12670_0, n12667_0, n12642_0, n12639_0, n12633_0, n12616_0, n12615_1, n12606_1, n12582_1, n10704_0/**/, n1941, n1933, n1845, n1837, n1829}), .out(n10788), .config_in(config_chain[18523:18518]), .config_rst(config_rst)); 
buffer_wire buffer_10788 (.in(n10788), .out(n10788_0));
mux15 mux_5623 (.in({n13735_1, n13706_0, n13701_0, n13687_0, n13658_0, n13653_0, n13651_1, n13646_1, n13562_1, n10871_1, n4879, n4867, n4779, n4771, n4763}), .out(n10789), .config_in(config_chain[18529:18524]), .config_rst(config_rst)); 
buffer_wire buffer_10789 (.in(n10789), .out(n10789_0));
mux15 mux_5624 (.in({n12679_1, n12664_0, n12661_0, n12653_0, n12636_0, n12630_0, n12627_0, n12608_1, n12574_1/**/, n10712_0, n1941, n1933, n1845, n1837, n1829}), .out(n10790), .config_in(config_chain[18535:18530]), .config_rst(config_rst)); 
buffer_wire buffer_10790 (.in(n10790), .out(n10790_0));
mux15 mux_5625 (.in({n13733_1, n13709_0, n13692_0, n13678_0, n13673_0, n13666_0, n13661_0, n13648_1, n13570_1, n10873_1, n4879, n4871, n4779/**/, n4771, n4763}), .out(n10791), .config_in(config_chain[18541:18536]), .config_rst(config_rst)); 
buffer_wire buffer_10791 (.in(n10791), .out(n10791_0));
mux15 mux_5626 (.in({n12681_1, n12675_0, n12658_0, n12650_0, n12647_0, n12624_0, n12621_0, n12610_1, n12566_1/**/, n10720_0, n1941, n1933, n1845, n1837, n1829}), .out(n10792), .config_in(config_chain[18547:18542]), .config_rst(config_rst)); 
buffer_wire buffer_10792 (.in(n10792), .out(n10792_0));
mux15 mux_5627 (.in({n13731_1, n13700_0, n13695_0, n13686_0, n13681_0/**/, n13669_0, n13652_0, n13650_1, n13578_1, n10875_1, n4879, n4871, n4863, n4771, n4763}), .out(n10793), .config_in(config_chain[18553:18548]), .config_rst(config_rst)); 
buffer_wire buffer_10793 (.in(n10793), .out(n10793_0));
mux15 mux_5628 (.in({n12683_1, n12672_0, n12669_0, n12644_0, n12641_0, n12635_0, n12618_0, n12612_1, n12558_1, n10728_0/**/, n1941, n1933, n1845, n1837, n1829}), .out(n10794), .config_in(config_chain[18559:18554]), .config_rst(config_rst)); 
buffer_wire buffer_10794 (.in(n10794), .out(n10794_0));
mux14 mux_5629 (.in({n13729_1, n13708_0, n13703_0, n13689_0, n13672_0, n13660_0, n13655_0, n13586_1, n10877_1, n4879, n4871/**/, n4863, n4775, n4763}), .out(n10795), .config_in(config_chain[18565:18560]), .config_rst(config_rst)); 
buffer_wire buffer_10795 (.in(n10795), .out(n10795_0));
mux15 mux_5630 (.in({n12685_1, n12666_0, n12663_0, n12655_0, n12638_0, n12632_0, n12629_0, n12614_1, n12550_1, n10736_0, n1945, n1937/**/, n1929, n1841, n1833}), .out(n10796), .config_in(config_chain[18571:18566]), .config_rst(config_rst)); 
buffer_wire buffer_10796 (.in(n10796), .out(n10796_0));
mux14 mux_5631 (.in({n13727_1, n13711_0, n13694_0, n13680_0, n13675_0, n13668_0, n13663_0/**/, n13594_1, n10879_1, n4879, n4871, n4863, n4775, n4767}), .out(n10797), .config_in(config_chain[18577:18572]), .config_rst(config_rst)); 
buffer_wire buffer_10797 (.in(n10797), .out(n10797_0));
mux15 mux_5632 (.in({n12687_1, n12660_0, n12657_0, n12652_0, n12649_0, n12626_0, n12623_0, n12605_0, n12542_1, n10744_0/**/, n1945, n1937, n1929, n1841, n1833}), .out(n10798), .config_in(config_chain[18583:18578]), .config_rst(config_rst)); 
buffer_wire buffer_10798 (.in(n10798), .out(n10798_0));
mux13 mux_5633 (.in({n13725_1, n13702_0, n13697_0/**/, n13688_0, n13683_0, n13671_0, n13654_0, n13602_1, n10881_1, n4871, n4863, n4775, n4767}), .out(n10799), .config_in(config_chain[18589:18584]), .config_rst(config_rst)); 
buffer_wire buffer_10799 (.in(n10799), .out(n10799_0));
mux15 mux_5634 (.in({n12689_1, n12674_0/**/, n12671_0, n12646_0, n12643_0, n12620_0, n12617_0, n12607_1, n12534_1, n10752_0, n1945, n1937, n1929, n1841, n1833}), .out(n10800), .config_in(config_chain[18595:18590]), .config_rst(config_rst)); 
buffer_wire buffer_10800 (.in(n10800), .out(n10800_0));
mux13 mux_5635 (.in({n13723_1, n13710_0, n13705_0, n13691_0, n13674_0, n13662_0, n13657_0/**/, n13610_1, n10883_1, n4875, n4863, n4775, n4767}), .out(n10801), .config_in(config_chain[18601:18596]), .config_rst(config_rst)); 
buffer_wire buffer_10801 (.in(n10801), .out(n10801_0));
mux15 mux_5636 (.in({n12691_1, n12668_0, n12665_0, n12640_0, n12637_0, n12634_0, n12631_0, n12609_1, n12526_1, n10760_0/**/, n1945, n1937, n1929, n1841, n1833}), .out(n10802), .config_in(config_chain[18607:18602]), .config_rst(config_rst)); 
buffer_wire buffer_10802 (.in(n10802), .out(n10802_0));
mux13 mux_5637 (.in({n13721_1, n13713_1, n13696_0, n13682_0, n13677_0, n13670_0/**/, n13665_0, n13618_1, n10885_1, n4875, n4867, n4775, n4767}), .out(n10803), .config_in(config_chain[18613:18608]), .config_rst(config_rst)); 
buffer_wire buffer_10803 (.in(n10803), .out(n10803_0));
mux15 mux_5638 (.in({n12693_1, n12662_0, n12659_0, n12654_0, n12651_0, n12628_0, n12625_0/**/, n12611_1, n12598_1, n10768_0, n1945, n1937, n1929, n1841, n1833}), .out(n10804), .config_in(config_chain[18619:18614]), .config_rst(config_rst)); 
buffer_wire buffer_10804 (.in(n10804), .out(n10804_0));
mux13 mux_5639 (.in({n13719_1/**/, n13704_0, n13699_0, n13690_0, n13685_0, n13656_0, n13645_0, n13626_1, n10887_1, n4875, n4867, n4779, n4767}), .out(n10805), .config_in(config_chain[18625:18620]), .config_rst(config_rst)); 
buffer_wire buffer_10805 (.in(n10805), .out(n10805_0));
mux16 mux_5640 (.in({n12951_1, n12918_0/**/, n12915_0, n12909_0, n12892_0, n12884_0, n12881_0, n12869_1, n12860_1, n12848_1, n10698_0, n2919, n2911, n2823, n2815, n2807}), .out(n10806), .config_in(config_chain[18631:18626]), .config_rst(config_rst)); 
buffer_wire buffer_10806 (.in(n10806), .out(n10806_0));
mux15 mux_5641 (.in({n13981_1, n13978_0, n13973_0, n13942_0, n13937_0, n13928_0, n13923_0, n13913_0, n13908_1, n10891_0, n5853, n5845, n5757, n5749, n5741}), .out(n10807), .config_in(config_chain[18637:18632]), .config_rst(config_rst)); 
buffer_wire buffer_10807 (.in(n10807), .out(n10807_0));
mux16 mux_5642 (.in({n12933_1, n12929_0, n12912_0, n12906_0, n12903_0/**/, n12878_0, n12875_0, n12871_1, n12862_1, n12840_1, n10706_0, n2919, n2911, n2823, n2815, n2807}), .out(n10808), .config_in(config_chain[18643:18638]), .config_rst(config_rst)); 
buffer_wire buffer_10808 (.in(n10808), .out(n10808_0));
mux15 mux_5643 (.in({n14001_1, n13964_0, n13959_0, n13950_0, n13945_0, n13931_0, n13915_0, n13910_1, n13828_1, n10893_0/**/, n5857, n5845, n5757, n5749, n5741}), .out(n10809), .config_in(config_chain[18649:18644]), .config_rst(config_rst)); 
buffer_wire buffer_10809 (.in(n10809), .out(n10809_0));
mux15 mux_5644 (.in({n12935_1, n12926_0, n12923_0, n12900_0, n12897_0, n12889_0, n12872_0/**/, n12864_1, n12832_1, n10714_0, n2919, n2911, n2823, n2815, n2807}), .out(n10810), .config_in(config_chain[18655:18650]), .config_rst(config_rst)); 
buffer_wire buffer_10810 (.in(n10810), .out(n10810_0));
mux15 mux_5645 (.in({n13999_1, n13972_0, n13967_0, n13953_0, n13936_0, n13922_0, n13917_0, n13912_1, n13836_1, n10895_0/**/, n5857, n5849, n5757, n5749, n5741}), .out(n10811), .config_in(config_chain[18661:18656]), .config_rst(config_rst)); 
buffer_wire buffer_10811 (.in(n10811), .out(n10811_0));
mux15 mux_5646 (.in({n12937_1, n12920_0, n12917_0, n12911_0, n12894_0, n12886_0/**/, n12883_0, n12866_1, n12824_1, n10722_0, n2919, n2911, n2823, n2815, n2807}), .out(n10812), .config_in(config_chain[18667:18662]), .config_rst(config_rst)); 
buffer_wire buffer_10812 (.in(n10812), .out(n10812_0));
mux15 mux_5647 (.in({n13997_1, n13975_0, n13958_0, n13944_0, n13939_0, n13930_0/**/, n13925_0, n13914_1, n13844_1, n10897_0, n5857, n5849, n5841, n5749, n5741}), .out(n10813), .config_in(config_chain[18673:18668]), .config_rst(config_rst)); 
buffer_wire buffer_10813 (.in(n10813), .out(n10813_0));
mux15 mux_5648 (.in({n12939_1/**/, n12931_0, n12914_0, n12908_0, n12905_0, n12880_0, n12877_0, n12868_1, n12816_1, n10730_0, n2919, n2911, n2823, n2815, n2807}), .out(n10814), .config_in(config_chain[18679:18674]), .config_rst(config_rst)); 
buffer_wire buffer_10814 (.in(n10814), .out(n10814_0));
mux14 mux_5649 (.in({n13995_1, n13966_0/**/, n13961_0, n13952_0, n13947_0, n13933_0, n13916_0, n13852_1, n10899_0, n5857, n5849, n5841, n5753, n5741}), .out(n10815), .config_in(config_chain[18685:18680]), .config_rst(config_rst)); 
buffer_wire buffer_10815 (.in(n10815), .out(n10815_0));
mux15 mux_5650 (.in({n12941_1, n12928_0, n12925_0, n12902_0/**/, n12899_0, n12891_0, n12874_0, n12870_1, n12808_1, n10738_0, n2923, n2915, n2907, n2819, n2811}), .out(n10816), .config_in(config_chain[18691:18686]), .config_rst(config_rst)); 
buffer_wire buffer_10816 (.in(n10816), .out(n10816_0));
mux14 mux_5651 (.in({n13993_1, n13974_0, n13969_0, n13955_0, n13938_0, n13924_0/**/, n13919_0, n13860_1, n10901_0, n5857, n5849, n5841, n5753, n5745}), .out(n10817), .config_in(config_chain[18697:18692]), .config_rst(config_rst)); 
buffer_wire buffer_10817 (.in(n10817), .out(n10817_0));
mux15 mux_5652 (.in({n12943_1, n12922_0, n12919_0, n12896_0, n12893_0, n12888_0, n12885_0, n12861_0, n12800_1, n10746_0, n2923, n2915/**/, n2907, n2819, n2811}), .out(n10818), .config_in(config_chain[18703:18698]), .config_rst(config_rst)); 
buffer_wire buffer_10818 (.in(n10818), .out(n10818_0));
mux13 mux_5653 (.in({n13991_1, n13977_0, n13960_0, n13946_0, n13941_0, n13932_0/**/, n13927_0, n13868_1, n10903_0, n5849, n5841, n5753, n5745}), .out(n10819), .config_in(config_chain[18709:18704]), .config_rst(config_rst)); 
buffer_wire buffer_10819 (.in(n10819), .out(n10819_0));
mux15 mux_5654 (.in({n12945_1, n12916_0, n12913_0, n12910_0, n12907_0, n12882_0, n12879_0, n12863_0, n12792_1, n10754_0, n2923/**/, n2915, n2907, n2819, n2811}), .out(n10820), .config_in(config_chain[18715:18710]), .config_rst(config_rst)); 
buffer_wire buffer_10820 (.in(n10820), .out(n10820_0));
mux13 mux_5655 (.in({n13989_1, n13968_0, n13963_0, n13954_0, n13949_0, n13935_0, n13918_0, n13876_1, n10905_0, n5853, n5841, n5753/**/, n5745}), .out(n10821), .config_in(config_chain[18721:18716]), .config_rst(config_rst)); 
buffer_wire buffer_10821 (.in(n10821), .out(n10821_0));
mux15 mux_5656 (.in({n12947_1, n12930_0, n12927_0, n12904_0, n12901_0, n12876_0, n12873_0/**/, n12865_1, n12784_1, n10762_0, n2923, n2915, n2907, n2819, n2811}), .out(n10822), .config_in(config_chain[18727:18722]), .config_rst(config_rst)); 
buffer_wire buffer_10822 (.in(n10822), .out(n10822_0));
mux13 mux_5657 (.in({n13987_1, n13976_0, n13971_0, n13957_1, n13940_0, n13926_0, n13921_0/**/, n13884_1, n10907_0, n5853, n5845, n5753, n5745}), .out(n10823), .config_in(config_chain[18733:18728]), .config_rst(config_rst)); 
buffer_wire buffer_10823 (.in(n10823), .out(n10823_0));
mux15 mux_5658 (.in({n12949_1, n12924_0, n12921_0, n12898_0, n12895_0, n12890_0/**/, n12887_0, n12867_1, n12856_1, n10770_0, n2923, n2915, n2907, n2819, n2811}), .out(n10824), .config_in(config_chain[18739:18734]), .config_rst(config_rst)); 
buffer_wire buffer_10824 (.in(n10824), .out(n10824_0));
mux13 mux_5659 (.in({n13985_1, n13979_1, n13962_0, n13948_0/**/, n13943_0, n13934_0, n13929_0, n13892_1, n10909_0, n5853, n5845, n5757, n5745}), .out(n10825), .config_in(config_chain[18745:18740]), .config_rst(config_rst)); 
buffer_wire buffer_10825 (.in(n10825), .out(n10825_0));
mux16 mux_5660 (.in({n13209_1, n13182_0/**/, n13179_0, n13156_0, n13153_0, n13147_0, n13130_0, n13127_1, n13118_1, n13108_1, n10700_0, n3897, n3889, n3801, n3793, n3785}), .out(n10826), .config_in(config_chain[18751:18746]), .config_rst(config_rst)); 
buffer_wire buffer_10826 (.in(n10826), .out(n10826_0));
mux15 mux_5661 (.in({n14247_1, n14236_0, n14231_0, n14222_0, n14217_0, n14186_0, n14181_0, n14177_0, n14174_1, n10913_0, n6831/**/, n6823, n6735, n6727, n6719}), .out(n10827), .config_in(config_chain[18757:18752]), .config_rst(config_rst)); 
buffer_wire buffer_10827 (.in(n10827), .out(n10827_0));
mux16 mux_5662 (.in({n13191_1, n13176_0, n13173_0, n13167_0, n13150_0, n13144_0, n13141_0, n13129_1, n13120_1, n13100_1, n10708_0/**/, n3897, n3889, n3801, n3793, n3785}), .out(n10828), .config_in(config_chain[18763:18758]), .config_rst(config_rst)); 
buffer_wire buffer_10828 (.in(n10828), .out(n10828_0));
mux15 mux_5663 (.in({n14267_1, n14244_0, n14239_0/**/, n14208_0, n14203_0, n14194_0, n14189_0, n14179_0, n14094_1, n10915_0, n6835, n6823, n6735, n6727, n6719}), .out(n10829), .config_in(config_chain[18769:18764]), .config_rst(config_rst)); 
buffer_wire buffer_10829 (.in(n10829), .out(n10829_0));
mux15 mux_5664 (.in({n13193_1, n13187_0, n13170_0, n13164_0/**/, n13161_0, n13138_0, n13135_0, n13122_1, n13092_1, n10716_0, n3897, n3889, n3801, n3793, n3785}), .out(n10830), .config_in(config_chain[18775:18770]), .config_rst(config_rst)); 
buffer_wire buffer_10830 (.in(n10830), .out(n10830_0));
mux15 mux_5665 (.in({n14265_1, n14230_0, n14225_0, n14216_0, n14211_0, n14197_0, n14180_0, n14176_1, n14102_1, n10917_0, n6835/**/, n6827, n6735, n6727, n6719}), .out(n10831), .config_in(config_chain[18781:18776]), .config_rst(config_rst)); 
buffer_wire buffer_10831 (.in(n10831), .out(n10831_0));
mux15 mux_5666 (.in({n13195_1, n13184_0, n13181_0, n13158_0, n13155_0, n13149_0/**/, n13132_0, n13124_1, n13084_1, n10724_0, n3897, n3889, n3801, n3793, n3785}), .out(n10832), .config_in(config_chain[18787:18782]), .config_rst(config_rst)); 
buffer_wire buffer_10832 (.in(n10832), .out(n10832_0));
mux15 mux_5667 (.in({n14263_1, n14238_0, n14233_0, n14219_0, n14202_0, n14188_0/**/, n14183_0, n14178_1, n14110_1, n10919_0, n6835, n6827, n6819, n6727, n6719}), .out(n10833), .config_in(config_chain[18793:18788]), .config_rst(config_rst)); 
buffer_wire buffer_10833 (.in(n10833), .out(n10833_0));
mux15 mux_5668 (.in({n13197_1, n13178_0, n13175_0, n13169_0/**/, n13152_0, n13146_0, n13143_0, n13126_1, n13076_1, n10732_0, n3897, n3889, n3801, n3793, n3785}), .out(n10834), .config_in(config_chain[18799:18794]), .config_rst(config_rst)); 
buffer_wire buffer_10834 (.in(n10834), .out(n10834_0));
mux14 mux_5669 (.in({n14261_1, n14241_0, n14224_0, n14210_0, n14205_0, n14196_0, n14191_0, n14118_1, n10921_0, n6835, n6827, n6819, n6731/**/, n6719}), .out(n10835), .config_in(config_chain[18805:18800]), .config_rst(config_rst)); 
buffer_wire buffer_10835 (.in(n10835), .out(n10835_0));
mux15 mux_5670 (.in({n13199_1, n13189_0, n13172_0/**/, n13166_0, n13163_0, n13140_0, n13137_0, n13128_1, n13068_1, n10740_0, n3901, n3893, n3885, n3797, n3789}), .out(n10836), .config_in(config_chain[18811:18806]), .config_rst(config_rst)); 
buffer_wire buffer_10836 (.in(n10836), .out(n10836_0));
mux14 mux_5671 (.in({n14259_1, n14232_0, n14227_0, n14218_0, n14213_0, n14199_0, n14182_0, n14126_1, n10923_0, n6835, n6827/**/, n6819, n6731, n6723}), .out(n10837), .config_in(config_chain[18817:18812]), .config_rst(config_rst)); 
buffer_wire buffer_10837 (.in(n10837), .out(n10837_0));
mux15 mux_5672 (.in({n13201_1, n13186_0, n13183_0, n13160_0, n13157_0, n13134_0, n13131_0, n13119_0, n13060_1, n10748_0/**/, n3901, n3893, n3885, n3797, n3789}), .out(n10838), .config_in(config_chain[18823:18818]), .config_rst(config_rst)); 
buffer_wire buffer_10838 (.in(n10838), .out(n10838_0));
mux13 mux_5673 (.in({n14257_1, n14240_0/**/, n14235_0, n14221_0, n14204_0, n14190_0, n14185_0, n14134_1, n10925_0, n6827, n6819, n6731, n6723}), .out(n10839), .config_in(config_chain[18829:18824]), .config_rst(config_rst)); 
buffer_wire buffer_10839 (.in(n10839), .out(n10839_0));
mux15 mux_5674 (.in({n13203_1, n13180_0, n13177_0, n13154_0, n13151_0, n13148_0, n13145_0, n13121_0, n13052_1, n10756_0, n3901, n3893, n3885, n3797, n3789/**/}), .out(n10840), .config_in(config_chain[18835:18830]), .config_rst(config_rst)); 
buffer_wire buffer_10840 (.in(n10840), .out(n10840_0));
mux13 mux_5675 (.in({n14255_1, n14243_0, n14226_0, n14212_0, n14207_0, n14198_0, n14193_0/**/, n14142_1, n10927_0, n6831, n6819, n6731, n6723}), .out(n10841), .config_in(config_chain[18841:18836]), .config_rst(config_rst)); 
buffer_wire buffer_10841 (.in(n10841), .out(n10841_0));
mux15 mux_5676 (.in({n13205_1, n13174_0, n13171_0, n13168_0, n13165_0, n13142_0, n13139_0, n13123_0, n13044_1, n10764_0/**/, n3901, n3893, n3885, n3797, n3789}), .out(n10842), .config_in(config_chain[18847:18842]), .config_rst(config_rst)); 
buffer_wire buffer_10842 (.in(n10842), .out(n10842_0));
mux13 mux_5677 (.in({n14253_1, n14234_0, n14229_0, n14220_0, n14215_0, n14201_1, n14184_0, n14150_1/**/, n10929_0, n6831, n6823, n6731, n6723}), .out(n10843), .config_in(config_chain[18853:18848]), .config_rst(config_rst)); 
buffer_wire buffer_10843 (.in(n10843), .out(n10843_0));
mux15 mux_5678 (.in({n13207_1, n13188_0, n13185_0, n13162_0, n13159_0, n13136_0/**/, n13133_0, n13125_1, n13116_1, n10772_0, n3901, n3893, n3885, n3797, n3789}), .out(n10844), .config_in(config_chain[18859:18854]), .config_rst(config_rst)); 
buffer_wire buffer_10844 (.in(n10844), .out(n10844_0));
mux13 mux_5679 (.in({n14251_1, n14242_0, n14237_0, n14223_1, n14206_0, n14192_0, n14187_0, n14158_1, n10931_0, n6831/**/, n6823, n6735, n6723}), .out(n10845), .config_in(config_chain[18865:18860]), .config_rst(config_rst)); 
buffer_wire buffer_10845 (.in(n10845), .out(n10845_0));
mux15 mux_5680 (.in({n13471_1, n13443_0, n13436_0, n13424_0, n13397_0/**/, n13390_0, n13386_1, n13383_0, n13370_1, n10694_1, n4875, n4867, n4779, n4771, n4763}), .out(n10846), .config_in(config_chain[18871:18866]), .config_rst(config_rst)); 
buffer_wire buffer_10846 (.in(n10846), .out(n10846_0));
mux15 mux_5681 (.in({n14511_1, n14509_1, n14500_0/**/, n14495_0, n14481_0, n14464_0, n14450_0, n14445_0, n14440_1, n10935_0, n7809, n7801, n7713, n7705, n7697}), .out(n10847), .config_in(config_chain[18877:18872]), .config_rst(config_rst)); 
buffer_wire buffer_10847 (.in(n10847), .out(n10847_0));
mux15 mux_5682 (.in({n13451_1, n13444_0, n13417_0, n13410_0, n13405_0, n13398_0, n13388_1, n13385_0, n13362_1, n10702_1, n4879, n4867, n4779, n4771, n4763/**/}), .out(n10848), .config_in(config_chain[18883:18878]), .config_rst(config_rst)); 
buffer_wire buffer_10848 (.in(n10848), .out(n10848_0));
mux15 mux_5683 (.in({n14531_1, n14503_0, n14486_0, n14472_0, n14467_0, n14458_0, n14453_0, n14443_0/**/, n14352_1, n10937_0, n7813, n7801, n7713, n7705, n7697}), .out(n10849), .config_in(config_chain[18889:18884]), .config_rst(config_rst)); 
buffer_wire buffer_10849 (.in(n10849), .out(n10849_0));
mux15 mux_5684 (.in({n13453_1, n13437_0, n13430_0, n13425_0, n13418_0, n13406_0, n13391_0/**/, n13387_1, n13354_1, n10710_1, n4879, n4871, n4779, n4771, n4763}), .out(n10850), .config_in(config_chain[18895:18890]), .config_rst(config_rst)); 
buffer_wire buffer_10850 (.in(n10850), .out(n10850_0));
mux15 mux_5685 (.in({n14529_1, n14508_0, n14494_0/**/, n14489_0, n14480_0, n14475_0, n14461_0, n14444_0, n14360_1, n10939_0, n7813, n7805, n7713, n7705, n7697}), .out(n10851), .config_in(config_chain[18901:18896]), .config_rst(config_rst)); 
buffer_wire buffer_10851 (.in(n10851), .out(n10851_0));
mux15 mux_5686 (.in({n13455_1, n13445_0, n13438_0, n13426_0, n13411_0, n13399_0, n13392_0, n13389_1, n13346_1, n10718_1/**/, n4879, n4871, n4863, n4771, n4763}), .out(n10852), .config_in(config_chain[18907:18902]), .config_rst(config_rst)); 
buffer_wire buffer_10852 (.in(n10852), .out(n10852_0));
mux15 mux_5687 (.in({n14527_1, n14502_0, n14497_0, n14483_0, n14466_0, n14452_0, n14447_0, n14442_1, n14368_1, n10941_0, n7813, n7805/**/, n7797, n7705, n7697}), .out(n10853), .config_in(config_chain[18913:18908]), .config_rst(config_rst)); 
buffer_wire buffer_10853 (.in(n10853), .out(n10853_0));
mux14 mux_5688 (.in({n13457_1, n13446_0, n13431_0/**/, n13419_0, n13412_0, n13407_0, n13400_0, n13338_1, n10726_1, n4879, n4871, n4863, n4775, n4763}), .out(n10854), .config_in(config_chain[18919:18914]), .config_rst(config_rst)); 
buffer_wire buffer_10854 (.in(n10854), .out(n10854_0));
mux14 mux_5689 (.in({n14525_1, n14505_0, n14488_0, n14474_0, n14469_0, n14460_0, n14455_0, n14376_1/**/, n10943_0, n7813, n7805, n7797, n7709, n7697}), .out(n10855), .config_in(config_chain[18925:18920]), .config_rst(config_rst)); 
buffer_wire buffer_10855 (.in(n10855), .out(n10855_0));
mux14 mux_5690 (.in({n13459_1, n13439_0, n13432_0, n13427_0, n13420_0, n13408_0, n13393_0, n13330_1, n10734_1, n4879/**/, n4871, n4863, n4775, n4767}), .out(n10856), .config_in(config_chain[18931:18926]), .config_rst(config_rst)); 
buffer_wire buffer_10856 (.in(n10856), .out(n10856_0));
mux14 mux_5691 (.in({n14523_1, n14496_0, n14491_0, n14482_0/**/, n14477_0, n14463_0, n14446_0, n14384_1, n10945_0, n7813, n7805, n7797, n7709, n7701}), .out(n10857), .config_in(config_chain[18937:18932]), .config_rst(config_rst)); 
buffer_wire buffer_10857 (.in(n10857), .out(n10857_0));
mux13 mux_5692 (.in({n13461_1, n13447_0, n13440_0/**/, n13428_0, n13413_0, n13401_0, n13394_0, n13322_1, n10742_1, n4871, n4863, n4775, n4767}), .out(n10858), .config_in(config_chain[18943:18938]), .config_rst(config_rst)); 
buffer_wire buffer_10858 (.in(n10858), .out(n10858_0));
mux13 mux_5693 (.in({n14521_1, n14504_0, n14499_0, n14485_0, n14468_0, n14454_0, n14449_0, n14392_1/**/, n10947_0, n7805, n7797, n7709, n7701}), .out(n10859), .config_in(config_chain[18949:18944]), .config_rst(config_rst)); 
buffer_wire buffer_10859 (.in(n10859), .out(n10859_0));
mux13 mux_5694 (.in({n13463_1, n13448_0, n13433_0, n13421_0, n13414_0, n13409_0, n13402_0, n13314_1, n10750_1/**/, n4875, n4863, n4775, n4767}), .out(n10860), .config_in(config_chain[18955:18950]), .config_rst(config_rst)); 
buffer_wire buffer_10860 (.in(n10860), .out(n10860_0));
mux13 mux_5695 (.in({n14519_1, n14507_0, n14490_0, n14476_0, n14471_0, n14462_0, n14457_0, n14400_1/**/, n10949_0, n7809, n7797, n7709, n7701}), .out(n10861), .config_in(config_chain[18961:18956]), .config_rst(config_rst)); 
buffer_wire buffer_10861 (.in(n10861), .out(n10861_0));
mux13 mux_5696 (.in({n13465_1, n13441_0, n13434_0, n13429_0, n13422_0, n13395_0, n13380_1, n13306_1, n10758_1, n4875, n4867, n4775, n4767/**/}), .out(n10862), .config_in(config_chain[18967:18962]), .config_rst(config_rst)); 
buffer_wire buffer_10862 (.in(n10862), .out(n10862_0));
mux13 mux_5697 (.in({n14517_1, n14498_0, n14493_0, n14484_0, n14479_0, n14448_0/**/, n14433_1, n14408_1, n10951_0, n7809, n7801, n7709, n7701}), .out(n10863), .config_in(config_chain[18973:18968]), .config_rst(config_rst)); 
buffer_wire buffer_10863 (.in(n10863), .out(n10863_0));
mux13 mux_5698 (.in({n13467_1, n13449_0, n13442_0, n13415_0, n13403_0, n13396_0/**/, n13382_1, n13298_1, n10766_1, n4875, n4867, n4779, n4767}), .out(n10864), .config_in(config_chain[18979:18974]), .config_rst(config_rst)); 
buffer_wire buffer_10864 (.in(n10864), .out(n10864_0));
mux13 mux_5699 (.in({n14515_1, n14506_0, n14501_0, n14470_0, n14465_1, n14456_0, n14451_0/**/, n14416_1, n10953_0, n7809, n7801, n7713, n7701}), .out(n10865), .config_in(config_chain[18985:18980]), .config_rst(config_rst)); 
buffer_wire buffer_10865 (.in(n10865), .out(n10865_0));
mux13 mux_5700 (.in({n13469_1, n13435_0, n13423_0, n13416_0, n13404_0, n13384_1, n13381_0/**/, n13378_1, n10774_1, n4875, n4867, n4779, n4771}), .out(n10866), .config_in(config_chain[18991:18986]), .config_rst(config_rst)); 
buffer_wire buffer_10866 (.in(n10866), .out(n10866_0));
mux3 mux_5701 (.in({n14695_1, n14694_1, n8787}), .out(n10867), .config_in(config_chain[18993:18992]), .config_rst(config_rst)); 
buffer_wire buffer_10867 (.in(n10867), .out(n10867_0));
mux15 mux_5702 (.in({n13735_1, n13699_0, n13692_0, n13685_0, n13678_0, n13666_0, n13648_1, n13645_0, n13634_1, n10786_1/**/, n5853, n5845, n5757, n5749, n5741}), .out(n10868), .config_in(config_chain[18999:18994]), .config_rst(config_rst)); 
buffer_wire buffer_10868 (.in(n10868), .out(n10868_0));
mux4 mux_5703 (.in({n14773_1, n14616_1, n8791, n8675}), .out(n10869), .config_in(config_chain[19001:19000]), .config_rst(config_rst)); 
buffer_wire buffer_10869 (.in(n10869), .out(n10869_0));
mux15 mux_5704 (.in({n13715_1, n13707_0, n13700_0, n13686_0, n13659_0, n13652_0, n13650_1, n13647_0, n13626_1, n10788_1/**/, n5857, n5845, n5757, n5749, n5741}), .out(n10870), .config_in(config_chain[19007:19002]), .config_rst(config_rst)); 
buffer_wire buffer_10870 (.in(n10870), .out(n10870_0));
mux3 mux_5705 (.in({n14775_1/**/, n14624_1, n8679}), .out(n10871), .config_in(config_chain[19009:19008]), .config_rst(config_rst)); 
buffer_wire buffer_10871 (.in(n10871), .out(n10871_0));
mux15 mux_5706 (.in({n13717_1, n13708_0, n13693_0/**/, n13679_0, n13672_0, n13667_0, n13660_0, n13649_0, n13618_1, n10790_1, n5857, n5849, n5757, n5749, n5741}), .out(n10872), .config_in(config_chain[19015:19010]), .config_rst(config_rst)); 
buffer_wire buffer_10872 (.in(n10872), .out(n10872_0));
mux3 mux_5707 (.in({n14777_1, n14632_1, n8679}), .out(n10873), .config_in(config_chain[19017:19016]), .config_rst(config_rst)); 
buffer_wire buffer_10873 (.in(n10873), .out(n10873_0));
mux15 mux_5708 (.in({n13719_1, n13701_0, n13694_0, n13687_0, n13680_0, n13668_0, n13653_0, n13651_1, n13610_1, n10792_1/**/, n5857, n5849, n5841, n5749, n5741}), .out(n10874), .config_in(config_chain[19023:19018]), .config_rst(config_rst)); 
buffer_wire buffer_10874 (.in(n10874), .out(n10874_0));
mux3 mux_5709 (.in({n14779_1, n14640_1, n8683}), .out(n10875), .config_in(config_chain[19025:19024]), .config_rst(config_rst)); 
buffer_wire buffer_10875 (.in(n10875), .out(n10875_0));
mux14 mux_5710 (.in({n13721_1, n13709_0/**/, n13702_0, n13688_0, n13673_0, n13661_0, n13654_0, n13602_1, n10794_1, n5857, n5849, n5841, n5753, n5741}), .out(n10876), .config_in(config_chain[19031:19026]), .config_rst(config_rst)); 
buffer_wire buffer_10876 (.in(n10876), .out(n10876_0));
mux3 mux_5711 (.in({n14781_1, n14648_1, n8687}), .out(n10877), .config_in(config_chain[19033:19032]), .config_rst(config_rst)); 
buffer_wire buffer_10877 (.in(n10877), .out(n10877_0));
mux14 mux_5712 (.in({n13723_1, n13710_0, n13695_0, n13681_0, n13674_0, n13669_0, n13662_0, n13594_1, n10796_1, n5857, n5849, n5841, n5753/**/, n5745}), .out(n10878), .config_in(config_chain[19039:19034]), .config_rst(config_rst)); 
buffer_wire buffer_10878 (.in(n10878), .out(n10878_0));
mux3 mux_5713 (.in({n14783_1, n14656_1/**/, n8691}), .out(n10879), .config_in(config_chain[19041:19040]), .config_rst(config_rst)); 
buffer_wire buffer_10879 (.in(n10879), .out(n10879_0));
mux13 mux_5714 (.in({n13725_1, n13703_0, n13696_0, n13689_0, n13682_0, n13670_0, n13655_0, n13586_1, n10798_1/**/, n5849, n5841, n5753, n5745}), .out(n10880), .config_in(config_chain[19047:19042]), .config_rst(config_rst)); 
buffer_wire buffer_10880 (.in(n10880), .out(n10880_0));
mux3 mux_5715 (.in({n14785_1, n14664_1, n8775}), .out(n10881), .config_in(config_chain[19049:19048]), .config_rst(config_rst)); 
buffer_wire buffer_10881 (.in(n10881), .out(n10881_0));
mux13 mux_5716 (.in({n13727_1, n13711_0, n13704_0, n13690_0, n13675_0, n13663_0, n13656_0, n13578_1, n10800_1/**/, n5853, n5841, n5753, n5745}), .out(n10882), .config_in(config_chain[19055:19050]), .config_rst(config_rst)); 
buffer_wire buffer_10882 (.in(n10882), .out(n10882_0));
mux3 mux_5717 (.in({n14787_1, n14672_1, n8775}), .out(n10883), .config_in(config_chain[19057:19056]), .config_rst(config_rst)); 
buffer_wire buffer_10883 (.in(n10883), .out(n10883_0));
mux13 mux_5718 (.in({n13729_1, n13712_0, n13697_0/**/, n13683_0, n13676_0, n13671_0, n13664_0, n13570_1, n10802_1, n5853, n5845, n5753, n5745}), .out(n10884), .config_in(config_chain[19063:19058]), .config_rst(config_rst)); 
buffer_wire buffer_10884 (.in(n10884), .out(n10884_0));
mux3 mux_5719 (.in({n14789_1, n14680_1, n8779}), .out(n10885), .config_in(config_chain[19065:19064]), .config_rst(config_rst)); 
buffer_wire buffer_10885 (.in(n10885), .out(n10885_0));
mux13 mux_5720 (.in({n13731_1, n13705_0, n13698_0, n13691_0, n13684_0, n13657_0, n13644_1, n13562_1, n10804_1, n5853, n5845, n5757, n5745/**/}), .out(n10886), .config_in(config_chain[19071:19066]), .config_rst(config_rst)); 
buffer_wire buffer_10886 (.in(n10886), .out(n10886_0));
mux3 mux_5721 (.in({n14791_1, n14688_1, n8783}), .out(n10887), .config_in(config_chain[19073:19072]), .config_rst(config_rst)); 
buffer_wire buffer_10887 (.in(n10887), .out(n10887_0));
mux13 mux_5722 (.in({n13733_1/**/, n13713_1, n13706_0, n13677_0, n13665_0, n13658_0, n13646_1, n13642_1, n10776_1, n5853, n5845, n5757, n5749}), .out(n10888), .config_in(config_chain[19079:19074]), .config_rst(config_rst)); 
buffer_wire buffer_10888 (.in(n10888), .out(n10888_0));
mux3 mux_5723 (.in({n14697_1, n14696_1, n8787}), .out(n10889), .config_in(config_chain[19081:19080]), .config_rst(config_rst)); 
buffer_wire buffer_10889 (.in(n10889), .out(n10889_0));
mux15 mux_5724 (.in({n14001_1, n13979_1, n13972_0, n13943_0, n13936_0, n13929_0, n13922_0, n13912_1, n13900_1, n10806_1, n6831, n6823, n6735, n6727, n6719}), .out(n10890), .config_in(config_chain[19087:19082]), .config_rst(config_rst)); 
buffer_wire buffer_10890 (.in(n10890), .out(n10890_0));
mux4 mux_5725 (.in({n14707_0/**/, n14706_0, n8791, n8675}), .out(n10891), .config_in(config_chain[19089:19088]), .config_rst(config_rst)); 
buffer_wire buffer_10891 (.in(n10891), .out(n10891_0));
mux15 mux_5726 (.in({n13981_1/**/, n13965_0, n13958_0, n13951_0, n13944_0, n13930_0, n13914_1, n13911_0, n13892_1, n10808_1, n6835, n6823, n6735, n6727, n6719}), .out(n10892), .config_in(config_chain[19095:19090]), .config_rst(config_rst)); 
buffer_wire buffer_10892 (.in(n10892), .out(n10892_0));
mux3 mux_5727 (.in({n14709_0/**/, n14708_0, n8679}), .out(n10893), .config_in(config_chain[19097:19096]), .config_rst(config_rst)); 
buffer_wire buffer_10893 (.in(n10893), .out(n10893_0));
mux15 mux_5728 (.in({n13983_1, n13973_0/**/, n13966_0, n13952_0, n13937_0, n13923_0, n13916_0, n13913_0, n13884_1, n10810_1, n6835, n6827, n6735, n6727, n6719}), .out(n10894), .config_in(config_chain[19103:19098]), .config_rst(config_rst)); 
buffer_wire buffer_10894 (.in(n10894), .out(n10894_0));
mux3 mux_5729 (.in({n14711_0/**/, n14710_0, n8683}), .out(n10895), .config_in(config_chain[19105:19104]), .config_rst(config_rst)); 
buffer_wire buffer_10895 (.in(n10895), .out(n10895_0));
mux15 mux_5730 (.in({n13985_1, n13974_0, n13959_0, n13945_0, n13938_0, n13931_0, n13924_0, n13915_0, n13876_1, n10812_1, n6835, n6827, n6819/**/, n6727, n6719}), .out(n10896), .config_in(config_chain[19111:19106]), .config_rst(config_rst)); 
buffer_wire buffer_10896 (.in(n10896), .out(n10896_0));
mux3 mux_5731 (.in({n14713_0/**/, n14712_0, n8683}), .out(n10897), .config_in(config_chain[19113:19112]), .config_rst(config_rst)); 
buffer_wire buffer_10897 (.in(n10897), .out(n10897_0));
mux14 mux_5732 (.in({n13987_1, n13967_0, n13960_0, n13953_0, n13946_0, n13932_0, n13917_0, n13868_1, n10814_1/**/, n6835, n6827, n6819, n6731, n6719}), .out(n10898), .config_in(config_chain[19119:19114]), .config_rst(config_rst)); 
buffer_wire buffer_10898 (.in(n10898), .out(n10898_0));
mux3 mux_5733 (.in({n14715_0, n14714_0, n8687}), .out(n10899), .config_in(config_chain[19121:19120]), .config_rst(config_rst)); 
buffer_wire buffer_10899 (.in(n10899), .out(n10899_0));
mux14 mux_5734 (.in({n13989_1, n13975_0, n13968_0/**/, n13954_0, n13939_0, n13925_0, n13918_0, n13860_1, n10816_1, n6835, n6827, n6819, n6731, n6723}), .out(n10900), .config_in(config_chain[19127:19122]), .config_rst(config_rst)); 
buffer_wire buffer_10900 (.in(n10900), .out(n10900_0));
mux3 mux_5735 (.in({n14717_0/**/, n14716_0, n8691}), .out(n10901), .config_in(config_chain[19129:19128]), .config_rst(config_rst)); 
buffer_wire buffer_10901 (.in(n10901), .out(n10901_0));
mux13 mux_5736 (.in({n13991_1, n13976_0, n13961_0, n13947_0/**/, n13940_0, n13933_0, n13926_0, n13852_1, n10818_1, n6827, n6819, n6731, n6723}), .out(n10902), .config_in(config_chain[19135:19130]), .config_rst(config_rst)); 
buffer_wire buffer_10902 (.in(n10902), .out(n10902_0));
mux3 mux_5737 (.in({n14719_0, n14718_0, n8775}), .out(n10903), .config_in(config_chain[19137:19136]), .config_rst(config_rst)); 
buffer_wire buffer_10903 (.in(n10903), .out(n10903_0));
mux13 mux_5738 (.in({n13993_1, n13969_0/**/, n13962_0, n13955_0, n13948_0, n13934_0, n13919_0, n13844_1, n10820_1, n6831, n6819, n6731, n6723}), .out(n10904), .config_in(config_chain[19143:19138]), .config_rst(config_rst)); 
buffer_wire buffer_10904 (.in(n10904), .out(n10904_0));
mux3 mux_5739 (.in({n14721_0, n14720_0, n8779/**/}), .out(n10905), .config_in(config_chain[19145:19144]), .config_rst(config_rst)); 
buffer_wire buffer_10905 (.in(n10905), .out(n10905_0));
mux13 mux_5740 (.in({n13995_1, n13977_0, n13970_0, n13956_0, n13941_0, n13927_0, n13920_0, n13836_1, n10822_1, n6831, n6823, n6731/**/, n6723}), .out(n10906), .config_in(config_chain[19151:19146]), .config_rst(config_rst)); 
buffer_wire buffer_10906 (.in(n10906), .out(n10906_0));
mux3 mux_5741 (.in({n14723_0, n14722_0, n8779/**/}), .out(n10907), .config_in(config_chain[19153:19152]), .config_rst(config_rst)); 
buffer_wire buffer_10907 (.in(n10907), .out(n10907_0));
mux13 mux_5742 (.in({n13997_1, n13978_0, n13963_0, n13949_0, n13942_0, n13935_0, n13928_0, n13828_1, n10824_1, n6831, n6823, n6735, n6723}), .out(n10908), .config_in(config_chain[19159:19154]), .config_rst(config_rst)); 
buffer_wire buffer_10908 (.in(n10908), .out(n10908_0));
mux3 mux_5743 (.in({n14725_0, n14724_0, n8783}), .out(n10909), .config_in(config_chain[19161:19160]), .config_rst(config_rst)); 
buffer_wire buffer_10909 (.in(n10909), .out(n10909_0));
mux13 mux_5744 (.in({n13999_1, n13971_0, n13964_0, n13957_1, n13950_0, n13921_0/**/, n13910_1, n13908_1, n10778_1, n6831, n6823, n6735, n6727}), .out(n10910), .config_in(config_chain[19167:19162]), .config_rst(config_rst)); 
buffer_wire buffer_10910 (.in(n10910), .out(n10910_0));
mux3 mux_5745 (.in({n14727_1, n14726_0, n8787}), .out(n10911), .config_in(config_chain[19169:19168]), .config_rst(config_rst)); 
buffer_wire buffer_10911 (.in(n10911), .out(n10911_0));
mux15 mux_5746 (.in({n14267_1, n14237_0, n14230_0, n14223_1, n14216_0, n14187_0, n14180_0, n14176_1, n14166_1, n10826_1, n7809/**/, n7801, n7713, n7705, n7697}), .out(n10912), .config_in(config_chain[19175:19170]), .config_rst(config_rst)); 
buffer_wire buffer_10912 (.in(n10912), .out(n10912_0));
mux4 mux_5747 (.in({n14729_0, n14728_0, n8791, n8675}), .out(n10913), .config_in(config_chain[19177:19176]), .config_rst(config_rst)); 
buffer_wire buffer_10913 (.in(n10913), .out(n10913_0));
mux15 mux_5748 (.in({n14247_1, n14245_1, n14238_0, n14209_0, n14202_0, n14195_0/**/, n14188_0, n14178_1, n14158_1, n10828_1, n7813, n7801, n7713, n7705, n7697}), .out(n10914), .config_in(config_chain[19183:19178]), .config_rst(config_rst)); 
buffer_wire buffer_10914 (.in(n10914), .out(n10914_0));
mux3 mux_5749 (.in({n14731_0, n14730_0, n8679}), .out(n10915), .config_in(config_chain[19185:19184]), .config_rst(config_rst)); 
buffer_wire buffer_10915 (.in(n10915), .out(n10915_0));
mux15 mux_5750 (.in({n14249_1, n14231_0, n14224_0, n14217_0, n14210_0, n14196_0, n14181_0, n14177_0, n14150_1, n10830_1, n7813, n7805, n7713, n7705, n7697}), .out(n10916), .config_in(config_chain[19191:19186]), .config_rst(config_rst)); 
buffer_wire buffer_10916 (.in(n10916), .out(n10916_0));
mux3 mux_5751 (.in({n14733_0, n14732_0, n8683}), .out(n10917), .config_in(config_chain[19193:19192]), .config_rst(config_rst)); 
buffer_wire buffer_10917 (.in(n10917), .out(n10917_0));
mux15 mux_5752 (.in({n14251_1, n14239_0, n14232_0/**/, n14218_0, n14203_0, n14189_0, n14182_0, n14179_0, n14142_1, n10832_1, n7813, n7805, n7797, n7705, n7697}), .out(n10918), .config_in(config_chain[19199:19194]), .config_rst(config_rst)); 
buffer_wire buffer_10918 (.in(n10918), .out(n10918_0));
mux3 mux_5753 (.in({n14735_0/**/, n14734_0, n8687}), .out(n10919), .config_in(config_chain[19201:19200]), .config_rst(config_rst)); 
buffer_wire buffer_10919 (.in(n10919), .out(n10919_0));
mux14 mux_5754 (.in({n14253_1, n14240_0, n14225_0, n14211_0, n14204_0, n14197_0, n14190_0, n14134_1, n10834_1, n7813, n7805, n7797, n7709, n7697}), .out(n10920), .config_in(config_chain[19207:19202]), .config_rst(config_rst)); 
buffer_wire buffer_10920 (.in(n10920), .out(n10920_0));
mux3 mux_5755 (.in({n14737_0, n14736_0, n8687}), .out(n10921), .config_in(config_chain[19209:19208]), .config_rst(config_rst)); 
buffer_wire buffer_10921 (.in(n10921), .out(n10921_0));
mux14 mux_5756 (.in({n14255_1, n14233_0, n14226_0, n14219_0, n14212_0, n14198_0, n14183_0/**/, n14126_1, n10836_1, n7813, n7805, n7797, n7709, n7701}), .out(n10922), .config_in(config_chain[19215:19210]), .config_rst(config_rst)); 
buffer_wire buffer_10922 (.in(n10922), .out(n10922_0));
mux3 mux_5757 (.in({n14739_0, n14738_0, n8691}), .out(n10923), .config_in(config_chain[19217:19216]), .config_rst(config_rst)); 
buffer_wire buffer_10923 (.in(n10923), .out(n10923_0));
mux13 mux_5758 (.in({n14257_1, n14241_0, n14234_0, n14220_0, n14205_0, n14191_0, n14184_0, n14118_1, n10838_1/**/, n7805, n7797, n7709, n7701}), .out(n10924), .config_in(config_chain[19223:19218]), .config_rst(config_rst)); 
buffer_wire buffer_10924 (.in(n10924), .out(n10924_0));
mux3 mux_5759 (.in({n14741_0/**/, n14740_0, n8775}), .out(n10925), .config_in(config_chain[19225:19224]), .config_rst(config_rst)); 
buffer_wire buffer_10925 (.in(n10925), .out(n10925_0));
mux13 mux_5760 (.in({n14259_1, n14242_0, n14227_0, n14213_0, n14206_0, n14199_0, n14192_0, n14110_1, n10840_1/**/, n7809, n7797, n7709, n7701}), .out(n10926), .config_in(config_chain[19231:19226]), .config_rst(config_rst)); 
buffer_wire buffer_10926 (.in(n10926), .out(n10926_0));
mux3 mux_5761 (.in({n14743_0, n14742_0, n8779}), .out(n10927), .config_in(config_chain[19233:19232]), .config_rst(config_rst)); 
buffer_wire buffer_10927 (.in(n10927), .out(n10927_0));
mux13 mux_5762 (.in({n14261_1, n14235_0, n14228_0, n14221_0, n14214_0/**/, n14200_0, n14185_0, n14102_1, n10842_1, n7809, n7801, n7709, n7701}), .out(n10928), .config_in(config_chain[19239:19234]), .config_rst(config_rst)); 
buffer_wire buffer_10928 (.in(n10928), .out(n10928_0));
mux3 mux_5763 (.in({n14745_0, n14744_0/**/, n8783}), .out(n10929), .config_in(config_chain[19241:19240]), .config_rst(config_rst)); 
buffer_wire buffer_10929 (.in(n10929), .out(n10929_0));
mux13 mux_5764 (.in({n14263_1, n14243_0, n14236_0, n14222_0, n14207_0, n14193_0, n14186_0, n14094_1, n10844_1, n7809, n7801, n7713/**/, n7701}), .out(n10930), .config_in(config_chain[19247:19242]), .config_rst(config_rst)); 
buffer_wire buffer_10930 (.in(n10930), .out(n10930_0));
mux3 mux_5765 (.in({n14747_0, n14746_0/**/, n8783}), .out(n10931), .config_in(config_chain[19249:19248]), .config_rst(config_rst)); 
buffer_wire buffer_10931 (.in(n10931), .out(n10931_0));
mux13 mux_5766 (.in({n14265_1, n14244_0, n14229_0, n14215_0, n14208_0, n14201_1, n14194_0, n14174_1, n10780_2, n7809, n7801, n7713, n7705}), .out(n10932), .config_in(config_chain[19255:19250]), .config_rst(config_rst)); 
buffer_wire buffer_10932 (.in(n10932), .out(n10932_0));
mux3 mux_5767 (.in({n14749_1, n14748_0, n8787}), .out(n10933), .config_in(config_chain[19257:19256]), .config_rst(config_rst)); 
buffer_wire buffer_10933 (.in(n10933), .out(n10933_0));
mux15 mux_5768 (.in({n14531_1, n14508_0, n14501_0/**/, n14494_0, n14480_0, n14465_1, n14451_0, n14444_0, n14424_1, n10846_1, n8787, n8779, n8691, n8683, n8675}), .out(n10934), .config_in(config_chain[19263:19258]), .config_rst(config_rst)); 
buffer_wire buffer_10934 (.in(n10934), .out(n10934_0));
mux4 mux_5769 (.in({n14751_0, n14750_0/**/, n8791, n8675}), .out(n10935), .config_in(config_chain[19265:19264]), .config_rst(config_rst)); 
buffer_wire buffer_10935 (.in(n10935), .out(n10935_0));
mux15 mux_5770 (.in({n14511_1, n14502_0, n14487_1, n14473_0, n14466_0, n14459_0, n14452_0, n14442_1, n14416_1, n10848_1, n8791, n8779, n8691/**/, n8683, n8675}), .out(n10936), .config_in(config_chain[19271:19266]), .config_rst(config_rst)); 
buffer_wire buffer_10936 (.in(n10936), .out(n10936_0));
mux3 mux_5771 (.in({n14753_0, n14752_0, n8675}), .out(n10937), .config_in(config_chain[19273:19272]), .config_rst(config_rst)); 
buffer_wire buffer_10937 (.in(n10937), .out(n10937_0));
mux15 mux_5772 (.in({n14513_1, n14509_1, n14495_0, n14488_0, n14481_0, n14474_0, n14460_0, n14445_0, n14408_1/**/, n10850_1, n8791, n8783, n8691, n8683, n8675}), .out(n10938), .config_in(config_chain[19279:19274]), .config_rst(config_rst)); 
buffer_wire buffer_10938 (.in(n10938), .out(n10938_0));
mux3 mux_5773 (.in({n14755_0, n14754_0, n8679}), .out(n10939), .config_in(config_chain[19281:19280]), .config_rst(config_rst)); 
buffer_wire buffer_10939 (.in(n10939), .out(n10939_0));
mux15 mux_5774 (.in({n14515_1, n14503_0, n14496_0, n14482_0, n14467_0, n14453_0, n14446_0, n14443_0, n14400_1/**/, n10852_1, n8791, n8783, n8775, n8683, n8675}), .out(n10940), .config_in(config_chain[19287:19282]), .config_rst(config_rst)); 
buffer_wire buffer_10940 (.in(n10940), .out(n10940_0));
mux3 mux_5775 (.in({n14757_0, n14756_0, n8683}), .out(n10941), .config_in(config_chain[19289:19288]), .config_rst(config_rst)); 
buffer_wire buffer_10941 (.in(n10941), .out(n10941_0));
mux14 mux_5776 (.in({n14517_1, n14504_0, n14489_0, n14475_0/**/, n14468_0, n14461_0, n14454_0, n14392_1, n10854_1, n8791, n8783, n8775, n8687, n8675}), .out(n10942), .config_in(config_chain[19295:19290]), .config_rst(config_rst)); 
buffer_wire buffer_10942 (.in(n10942), .out(n10942_0));
mux3 mux_5777 (.in({n14759_0, n14758_0, n8687}), .out(n10943), .config_in(config_chain[19297:19296]), .config_rst(config_rst)); 
buffer_wire buffer_10943 (.in(n10943), .out(n10943_0));
mux14 mux_5778 (.in({n14519_1, n14497_0, n14490_0, n14483_0, n14476_0, n14462_0, n14447_0, n14384_1, n10856_1, n8791/**/, n8783, n8775, n8687, n8679}), .out(n10944), .config_in(config_chain[19303:19298]), .config_rst(config_rst)); 
buffer_wire buffer_10944 (.in(n10944), .out(n10944_0));
mux3 mux_5779 (.in({n14761_0, n14760_0, n8691}), .out(n10945), .config_in(config_chain[19305:19304]), .config_rst(config_rst)); 
buffer_wire buffer_10945 (.in(n10945), .out(n10945_0));
mux13 mux_5780 (.in({n14521_1, n14505_0, n14498_0, n14484_0, n14469_0, n14455_0, n14448_0, n14376_1/**/, n10858_1, n8783, n8775, n8687, n8679}), .out(n10946), .config_in(config_chain[19311:19306]), .config_rst(config_rst)); 
buffer_wire buffer_10946 (.in(n10946), .out(n10946_0));
mux3 mux_5781 (.in({n14763_0/**/, n14762_0, n8691}), .out(n10947), .config_in(config_chain[19313:19312]), .config_rst(config_rst)); 
buffer_wire buffer_10947 (.in(n10947), .out(n10947_0));
mux13 mux_5782 (.in({n14523_1, n14506_0, n14491_0, n14477_0, n14470_0, n14463_0, n14456_0, n14368_1, n10860_1/**/, n8787, n8775, n8687, n8679}), .out(n10948), .config_in(config_chain[19319:19314]), .config_rst(config_rst)); 
buffer_wire buffer_10948 (.in(n10948), .out(n10948_0));
mux3 mux_5783 (.in({n14765_0, n14764_0, n8775}), .out(n10949), .config_in(config_chain[19321:19320]), .config_rst(config_rst)); 
buffer_wire buffer_10949 (.in(n10949), .out(n10949_0));
mux13 mux_5784 (.in({n14525_1, n14499_0, n14492_0, n14485_0, n14478_0, n14449_0, n14432_1, n14360_1/**/, n10862_1, n8787, n8779, n8687, n8679}), .out(n10950), .config_in(config_chain[19327:19322]), .config_rst(config_rst)); 
buffer_wire buffer_10950 (.in(n10950), .out(n10950_0));
mux3 mux_5785 (.in({n14767_0, n14766_0, n8779}), .out(n10951), .config_in(config_chain[19329:19328]), .config_rst(config_rst)); 
buffer_wire buffer_10951 (.in(n10951), .out(n10951_0));
mux13 mux_5786 (.in({n14527_1, n14507_0, n14500_0, n14471_0, n14464_0, n14457_0, n14450_0, n14352_1, n10864_1, n8787, n8779, n8691, n8679}), .out(n10952), .config_in(config_chain[19335:19330]), .config_rst(config_rst)); 
buffer_wire buffer_10952 (.in(n10952), .out(n10952_0));
mux3 mux_5787 (.in({n14769_0, n14768_0, n8783}), .out(n10953), .config_in(config_chain[19337:19336]), .config_rst(config_rst)); 
buffer_wire buffer_10953 (.in(n10953), .out(n10953_0));
mux13 mux_5788 (.in({n14529_1, n14493_0, n14486_0, n14479_0, n14472_0, n14458_0, n14440_1, n14433_1, n10782_2, n8787, n8779, n8691, n8683}), .out(n10954), .config_in(config_chain[19343:19338]), .config_rst(config_rst)); 
buffer_wire buffer_10954 (.in(n10954), .out(n10954_0));
mux3 mux_5789 (.in({n14771_1, n14770_0, n8787}), .out(n10955), .config_in(config_chain[19345:19344]), .config_rst(config_rst)); 
buffer_wire buffer_10955 (.in(n10955), .out(n10955_0));
mux4 mux_5790 (.in({n12423_0, n12422_0/**/, n1065, n949}), .out(n10956), .config_in(config_chain[19347:19346]), .config_rst(config_rst)); 
buffer_wire buffer_10956 (.in(n10956), .out(n10956_0));
mux15 mux_5791 (.in({n13211_1, n13202_0, n13197_0, n13185_0, n13156_0, n13151_0, n13127_1, n13122_1, n13118_1, n11089_1/**/, n3017, n3009, n2921, n2913, n2905}), .out(n10957), .config_in(config_chain[19353:19348]), .config_rst(config_rst)); 
buffer_wire buffer_10957 (.in(n10957), .out(n10957_0));
mux4 mux_5792 (.in({n12443_1, n12362_1, n1065, n949/**/}), .out(n10958), .config_in(config_chain[19355:19354]), .config_rst(config_rst)); 
buffer_wire buffer_10958 (.in(n10958), .out(n10958_0));
mux15 mux_5793 (.in({n13473_1, n13456_0, n13451_0, n13442_0, n13437_0, n13425_0, n13387_0, n13382_1, n13380_1, n11111_1, n3995, n3987, n3899, n3891, n3883}), .out(n10959), .config_in(config_chain[19361:19356]), .config_rst(config_rst)); 
buffer_wire buffer_10959 (.in(n10959), .out(n10959_0));
mux4 mux_5794 (.in({n12383_0, n12382_0, n1065, n949/**/}), .out(n10960), .config_in(config_chain[19363:19362]), .config_rst(config_rst)); 
buffer_wire buffer_10960 (.in(n10960), .out(n10960_0));
mux16 mux_5795 (.in({n12697_1, n12683_0, n12678_0, n12672_0, n12657_0, n12649_0, n12644_0, n12634_1, n12612_1, n12605_0, n11049_1, n1061, n1053, n965, n957, n949}), .out(n10961), .config_in(config_chain[19369:19364]), .config_rst(config_rst)); 
buffer_wire buffer_10961 (.in(n10961), .out(n10961_0));
mux4 mux_5796 (.in({n12403_0, n12402_0, n1065, n949}), .out(n10962), .config_in(config_chain[19371:19370]), .config_rst(config_rst)); 
buffer_wire buffer_10962 (.in(n10962), .out(n10962_0));
mux16 mux_5797 (.in({n12953_1, n12945_0, n12940_0, n12919_0, n12914_0, n12908_0, n12893_0, n12890_1, n12868_1, n12861_0, n11069_1, n2039, n2031, n1943, n1935, n1927}), .out(n10963), .config_in(config_chain[19377:19372]), .config_rst(config_rst)); 
buffer_wire buffer_10963 (.in(n10963), .out(n10963_0));
mux3 mux_5798 (.in({n12425_0, n12424_0, n949/**/}), .out(n10964), .config_in(config_chain[19379:19378]), .config_rst(config_rst)); 
buffer_wire buffer_10964 (.in(n10964), .out(n10964_0));
mux15 mux_5799 (.in({n13231_1, n13205_0, n13176_0, n13171_0, n13164_0/**/, n13159_0, n13130_1, n13129_1, n13124_1, n11091_1, n3021, n3009, n2921, n2913, n2905}), .out(n10965), .config_in(config_chain[19385:19380]), .config_rst(config_rst)); 
buffer_wire buffer_10965 (.in(n10965), .out(n10965_0));
mux3 mux_5800 (.in({n12445_1, n12364_1/**/, n953}), .out(n10966), .config_in(config_chain[19387:19386]), .config_rst(config_rst)); 
buffer_wire buffer_10966 (.in(n10966), .out(n10966_0));
mux15 mux_5801 (.in({n13493_1, n13464_0, n13459_0, n13445_0, n13416_0, n13411_0, n13390_1, n13389_1, n13384_1, n11113_1, n3999, n3987, n3899, n3891, n3883}), .out(n10967), .config_in(config_chain[19393:19388]), .config_rst(config_rst)); 
buffer_wire buffer_10967 (.in(n10967), .out(n10967_0));
mux3 mux_5802 (.in({n12385_0, n12384_0, n953}), .out(n10968), .config_in(config_chain[19395:19394]), .config_rst(config_rst)); 
buffer_wire buffer_10968 (.in(n10968), .out(n10968_0));
mux16 mux_5803 (.in({n12715_1, n12692_0, n12677_0, n12671_0, n12666_0, n12643_0, n12638_0, n12616_1, n12614_1, n12607_0, n11051_1, n1061, n1053, n965, n957, n949/**/}), .out(n10969), .config_in(config_chain[19401:19396]), .config_rst(config_rst)); 
buffer_wire buffer_10969 (.in(n10969), .out(n10969_0));
mux3 mux_5804 (.in({n12405_0/**/, n12404_0, n953}), .out(n10970), .config_in(config_chain[19403:19402]), .config_rst(config_rst)); 
buffer_wire buffer_10970 (.in(n10970), .out(n10970_0));
mux16 mux_5805 (.in({n12971_1, n12939_0, n12934_0, n12928_0, n12913_0, n12907_0, n12902_0, n12872_1, n12870_1, n12863_0, n11071_1, n2039, n2031, n1943/**/, n1935, n1927}), .out(n10971), .config_in(config_chain[19409:19404]), .config_rst(config_rst)); 
buffer_wire buffer_10971 (.in(n10971), .out(n10971_0));
mux3 mux_5806 (.in({n12427_0, n12426_0/**/, n953}), .out(n10972), .config_in(config_chain[19411:19410]), .config_rst(config_rst)); 
buffer_wire buffer_10972 (.in(n10972), .out(n10972_0));
mux15 mux_5807 (.in({n13229_1, n13196_0, n13191_0, n13184_0, n13179_0, n13167_0, n13150_0, n13132_1, n13126_1, n11093_1, n3021, n3013, n2921, n2913, n2905}), .out(n10973), .config_in(config_chain[19417:19412]), .config_rst(config_rst)); 
buffer_wire buffer_10973 (.in(n10973), .out(n10973_0));
mux3 mux_5808 (.in({n12447_1, n12366_1/**/, n953}), .out(n10974), .config_in(config_chain[19419:19418]), .config_rst(config_rst)); 
buffer_wire buffer_10974 (.in(n10974), .out(n10974_0));
mux15 mux_5809 (.in({n13491_1, n13467_0/**/, n13450_0, n13436_0, n13431_0, n13424_0, n13419_0, n13392_1, n13386_1, n11115_1, n3999, n3991, n3899, n3891, n3883}), .out(n10975), .config_in(config_chain[19425:19420]), .config_rst(config_rst)); 
buffer_wire buffer_10975 (.in(n10975), .out(n10975_0));
mux3 mux_5810 (.in({n12387_0, n12386_0, n957}), .out(n10976), .config_in(config_chain[19427:19426]), .config_rst(config_rst)); 
buffer_wire buffer_10976 (.in(n10976), .out(n10976_0));
mux15 mux_5811 (.in({n12713_1/**/, n12691_0, n12686_0, n12665_0, n12660_0, n12652_0, n12637_0, n12618_1, n12609_1, n11053_1, n1061, n1053, n965, n957, n949}), .out(n10977), .config_in(config_chain[19433:19428]), .config_rst(config_rst)); 
buffer_wire buffer_10977 (.in(n10977), .out(n10977_0));
mux3 mux_5812 (.in({n12407_0, n12406_0, n957}), .out(n10978), .config_in(config_chain[19435:19434]), .config_rst(config_rst)); 
buffer_wire buffer_10978 (.in(n10978), .out(n10978_0));
mux15 mux_5813 (.in({n12969_1, n12948_0, n12933_0, n12927_0, n12922_0/**/, n12901_0, n12896_0, n12874_1, n12865_0, n11073_1, n2039, n2031, n1943, n1935, n1927}), .out(n10979), .config_in(config_chain[19441:19436]), .config_rst(config_rst)); 
buffer_wire buffer_10979 (.in(n10979), .out(n10979_0));
mux3 mux_5814 (.in({n12429_0, n12428_0/**/, n957}), .out(n10980), .config_in(config_chain[19443:19442]), .config_rst(config_rst)); 
buffer_wire buffer_10980 (.in(n10980), .out(n10980_0));
mux15 mux_5815 (.in({n13227_1, n13204_0/**/, n13199_0, n13187_0, n13170_0, n13158_0, n13153_0, n13134_1, n13128_1, n11095_1, n3021, n3013, n3005, n2913, n2905}), .out(n10981), .config_in(config_chain[19449:19444]), .config_rst(config_rst)); 
buffer_wire buffer_10981 (.in(n10981), .out(n10981_0));
mux3 mux_5816 (.in({n12449_1, n12368_1, n957}), .out(n10982), .config_in(config_chain[19451:19450]), .config_rst(config_rst)); 
buffer_wire buffer_10982 (.in(n10982), .out(n10982_0));
mux15 mux_5817 (.in({n13489_1, n13458_0, n13453_0, n13444_0, n13439_0/**/, n13427_0, n13410_0, n13394_1, n13388_1, n11117_1, n3999, n3991, n3983, n3891, n3883}), .out(n10983), .config_in(config_chain[19457:19452]), .config_rst(config_rst)); 
buffer_wire buffer_10983 (.in(n10983), .out(n10983_0));
mux3 mux_5818 (.in({n12389_0/**/, n12388_0, n957}), .out(n10984), .config_in(config_chain[19459:19458]), .config_rst(config_rst)); 
buffer_wire buffer_10984 (.in(n10984), .out(n10984_0));
mux15 mux_5819 (.in({n12711_1, n12685_0, n12680_0, n12674_0, n12659_0, n12651_0, n12646_0, n12620_1, n12611_1, n11055_1, n1061, n1053, n965, n957, n949}), .out(n10985), .config_in(config_chain[19465:19460]), .config_rst(config_rst)); 
buffer_wire buffer_10985 (.in(n10985), .out(n10985_0));
mux3 mux_5820 (.in({n12409_0, n12408_0/**/, n961}), .out(n10986), .config_in(config_chain[19467:19466]), .config_rst(config_rst)); 
buffer_wire buffer_10986 (.in(n10986), .out(n10986_0));
mux15 mux_5821 (.in({n12967_1, n12947_0, n12942_0, n12921_0, n12916_0, n12910_0, n12895_0, n12876_1, n12867_1, n11075_1, n2039, n2031, n1943, n1935, n1927/**/}), .out(n10987), .config_in(config_chain[19473:19468]), .config_rst(config_rst)); 
buffer_wire buffer_10987 (.in(n10987), .out(n10987_0));
mux3 mux_5822 (.in({n12431_0, n12430_0/**/, n961}), .out(n10988), .config_in(config_chain[19475:19474]), .config_rst(config_rst)); 
buffer_wire buffer_10988 (.in(n10988), .out(n10988_0));
mux14 mux_5823 (.in({n13225_1, n13207_0, n13190_0, n13178_0, n13173_0, n13166_0, n13161_0, n13136_1, n11097_1, n3021, n3013, n3005, n2917/**/, n2905}), .out(n10989), .config_in(config_chain[19481:19476]), .config_rst(config_rst)); 
buffer_wire buffer_10989 (.in(n10989), .out(n10989_0));
mux3 mux_5824 (.in({n12451_1, n12370_1/**/, n961}), .out(n10990), .config_in(config_chain[19483:19482]), .config_rst(config_rst)); 
buffer_wire buffer_10990 (.in(n10990), .out(n10990_0));
mux14 mux_5825 (.in({n13487_1, n13466_0, n13461_0, n13447_0, n13430_0, n13418_0, n13413_0, n13396_1/**/, n11119_1, n3999, n3991, n3983, n3895, n3883}), .out(n10991), .config_in(config_chain[19489:19484]), .config_rst(config_rst)); 
buffer_wire buffer_10991 (.in(n10991), .out(n10991_0));
mux3 mux_5826 (.in({n12391_0, n12390_0, n961}), .out(n10992), .config_in(config_chain[19491:19490]), .config_rst(config_rst)); 
buffer_wire buffer_10992 (.in(n10992), .out(n10992_0));
mux15 mux_5827 (.in({n12709_1, n12694_0, n12679_0, n12673_0, n12668_0, n12645_0, n12640_0, n12622_1, n12613_1, n11057_1, n1061, n1053, n965, n957, n949}), .out(n10993), .config_in(config_chain[19497:19492]), .config_rst(config_rst)); 
buffer_wire buffer_10993 (.in(n10993), .out(n10993_0));
mux3 mux_5828 (.in({n12411_0, n12410_0, n961}), .out(n10994), .config_in(config_chain[19499:19498]), .config_rst(config_rst)); 
buffer_wire buffer_10994 (.in(n10994), .out(n10994_0));
mux15 mux_5829 (.in({n12965_1, n12941_0, n12936_0, n12930_0/**/, n12915_0, n12909_0, n12904_0, n12878_1, n12869_1, n11077_1, n2039, n2031, n1943, n1935, n1927}), .out(n10995), .config_in(config_chain[19505:19500]), .config_rst(config_rst)); 
buffer_wire buffer_10995 (.in(n10995), .out(n10995_0));
mux3 mux_5830 (.in({n12433_0, n12432_0/**/, n965}), .out(n10996), .config_in(config_chain[19507:19506]), .config_rst(config_rst)); 
buffer_wire buffer_10996 (.in(n10996), .out(n10996_0));
mux14 mux_5831 (.in({n13223_1, n13198_0, n13193_0, n13186_0, n13181_0/**/, n13169_0, n13152_0, n13138_1, n11099_1, n3021, n3013, n3005, n2917, n2909}), .out(n10997), .config_in(config_chain[19513:19508]), .config_rst(config_rst)); 
buffer_wire buffer_10997 (.in(n10997), .out(n10997_0));
mux3 mux_5832 (.in({n12453_1, n12372_1/**/, n965}), .out(n10998), .config_in(config_chain[19515:19514]), .config_rst(config_rst)); 
buffer_wire buffer_10998 (.in(n10998), .out(n10998_0));
mux14 mux_5833 (.in({n13485_1, n13469_0, n13452_0, n13438_0, n13433_0, n13426_0, n13421_0, n13398_1, n11121_1, n3999, n3991, n3983/**/, n3895, n3887}), .out(n10999), .config_in(config_chain[19521:19516]), .config_rst(config_rst)); 
buffer_wire buffer_10999 (.in(n10999), .out(n10999_0));
mux3 mux_5834 (.in({n12393_0, n12392_0, n965}), .out(n11000), .config_in(config_chain[19523:19522]), .config_rst(config_rst)); 
buffer_wire buffer_11000 (.in(n11000), .out(n11000_0));
mux15 mux_5835 (.in({n12707_1, n12693_0, n12688_0, n12667_0, n12662_0, n12654_0, n12639_0, n12624_1, n12615_1, n11059_1/**/, n1065, n1057, n1049, n961, n953}), .out(n11001), .config_in(config_chain[19529:19524]), .config_rst(config_rst)); 
buffer_wire buffer_11001 (.in(n11001), .out(n11001_0));
mux3 mux_5836 (.in({n12413_0, n12412_0/**/, n965}), .out(n11002), .config_in(config_chain[19531:19530]), .config_rst(config_rst)); 
buffer_wire buffer_11002 (.in(n11002), .out(n11002_0));
mux15 mux_5837 (.in({n12963_1, n12950_0, n12935_0, n12929_0, n12924_0, n12903_0, n12898_0, n12880_1, n12871_1, n11079_1, n2043, n2035, n2027, n1939, n1931}), .out(n11003), .config_in(config_chain[19537:19532]), .config_rst(config_rst)); 
buffer_wire buffer_11003 (.in(n11003), .out(n11003_0));
mux3 mux_5838 (.in({n12435_0, n12434_0, n965}), .out(n11004), .config_in(config_chain[19539:19538]), .config_rst(config_rst)); 
buffer_wire buffer_11004 (.in(n11004), .out(n11004_0));
mux13 mux_5839 (.in({n13221_1, n13206_0, n13201_0/**/, n13189_0, n13172_0, n13160_0, n13155_0, n13140_1, n11101_1, n3013, n3005, n2917, n2909}), .out(n11005), .config_in(config_chain[19545:19540]), .config_rst(config_rst)); 
buffer_wire buffer_11005 (.in(n11005), .out(n11005_0));
mux3 mux_5840 (.in({n12455_1, n12374_1/**/, n1049}), .out(n11006), .config_in(config_chain[19547:19546]), .config_rst(config_rst)); 
buffer_wire buffer_11006 (.in(n11006), .out(n11006_0));
mux13 mux_5841 (.in({n13483_1/**/, n13460_0, n13455_0, n13446_0, n13441_0, n13429_0, n13412_0, n13400_1, n11123_1, n3991, n3983, n3895, n3887}), .out(n11007), .config_in(config_chain[19553:19548]), .config_rst(config_rst)); 
buffer_wire buffer_11007 (.in(n11007), .out(n11007_0));
mux3 mux_5842 (.in({n12395_0, n12394_0, n1049}), .out(n11008), .config_in(config_chain[19555:19554]), .config_rst(config_rst)); 
buffer_wire buffer_11008 (.in(n11008), .out(n11008_0));
mux15 mux_5843 (.in({n12705_1, n12687_0, n12682_0, n12661_0, n12656_0, n12653_0, n12648_0/**/, n12626_1, n12604_1, n11061_1, n1065, n1057, n1049, n961, n953}), .out(n11009), .config_in(config_chain[19561:19556]), .config_rst(config_rst)); 
buffer_wire buffer_11009 (.in(n11009), .out(n11009_0));
mux3 mux_5844 (.in({n12415_0/**/, n12414_0, n1049}), .out(n11010), .config_in(config_chain[19563:19562]), .config_rst(config_rst)); 
buffer_wire buffer_11010 (.in(n11010), .out(n11010_0));
mux15 mux_5845 (.in({n12961_1, n12949_0, n12944_0, n12923_0, n12918_0, n12897_0, n12892_0, n12882_1, n12860_1, n11081_1, n2043, n2035, n2027, n1939, n1931}), .out(n11011), .config_in(config_chain[19569:19564]), .config_rst(config_rst)); 
buffer_wire buffer_11011 (.in(n11011), .out(n11011_0));
mux3 mux_5846 (.in({n12437_0, n12436_0/**/, n1049}), .out(n11012), .config_in(config_chain[19571:19570]), .config_rst(config_rst)); 
buffer_wire buffer_11012 (.in(n11012), .out(n11012_0));
mux13 mux_5847 (.in({n13219_1, n13209_0, n13192_0, n13180_0/**/, n13175_0, n13168_0, n13163_0, n13142_1, n11103_1, n3017, n3005, n2917, n2909}), .out(n11013), .config_in(config_chain[19577:19572]), .config_rst(config_rst)); 
buffer_wire buffer_11013 (.in(n11013), .out(n11013_0));
mux3 mux_5848 (.in({n12457_1, n12376_1/**/, n1049}), .out(n11014), .config_in(config_chain[19579:19578]), .config_rst(config_rst)); 
buffer_wire buffer_11014 (.in(n11014), .out(n11014_0));
mux13 mux_5849 (.in({n13481_1, n13468_0, n13463_0, n13449_0, n13432_0, n13420_0, n13415_0, n13402_1, n11125_1, n3995, n3983/**/, n3895, n3887}), .out(n11015), .config_in(config_chain[19585:19580]), .config_rst(config_rst)); 
buffer_wire buffer_11015 (.in(n11015), .out(n11015_0));
mux3 mux_5850 (.in({n12397_0, n12396_0, n1053}), .out(n11016), .config_in(config_chain[19587:19586]), .config_rst(config_rst)); 
buffer_wire buffer_11016 (.in(n11016), .out(n11016_0));
mux15 mux_5851 (.in({n12703_1, n12681_0, n12676_0, n12675_0, n12670_0, n12647_0, n12642_0, n12628_1/**/, n12606_1, n11063_1, n1065, n1057, n1049, n961, n953}), .out(n11017), .config_in(config_chain[19593:19588]), .config_rst(config_rst)); 
buffer_wire buffer_11017 (.in(n11017), .out(n11017_0));
mux3 mux_5852 (.in({n12417_0, n12416_0, n1053/**/}), .out(n11018), .config_in(config_chain[19595:19594]), .config_rst(config_rst)); 
buffer_wire buffer_11018 (.in(n11018), .out(n11018_0));
mux15 mux_5853 (.in({n12959_1, n12943_0, n12938_0, n12917_0, n12912_0/**/, n12911_0, n12906_0, n12884_1, n12862_1, n11083_1, n2043, n2035, n2027, n1939, n1931}), .out(n11019), .config_in(config_chain[19601:19596]), .config_rst(config_rst)); 
buffer_wire buffer_11019 (.in(n11019), .out(n11019_0));
mux3 mux_5854 (.in({n12439_0, n12438_0/**/, n1053}), .out(n11020), .config_in(config_chain[19603:19602]), .config_rst(config_rst)); 
buffer_wire buffer_11020 (.in(n11020), .out(n11020_0));
mux13 mux_5855 (.in({n13217_1, n13200_0, n13195_0, n13188_0/**/, n13183_0, n13154_0, n13144_1, n13121_0, n11105_1, n3017, n3009, n2917, n2909}), .out(n11021), .config_in(config_chain[19609:19604]), .config_rst(config_rst)); 
buffer_wire buffer_11021 (.in(n11021), .out(n11021_0));
mux3 mux_5856 (.in({n12459_1, n12378_1/**/, n1053}), .out(n11022), .config_in(config_chain[19611:19610]), .config_rst(config_rst)); 
buffer_wire buffer_11022 (.in(n11022), .out(n11022_0));
mux13 mux_5857 (.in({n13479_1, n13471_1, n13454_0/**/, n13440_0, n13435_0, n13428_0, n13423_0, n13404_1, n11127_1, n3995, n3987, n3895, n3887}), .out(n11023), .config_in(config_chain[19617:19612]), .config_rst(config_rst)); 
buffer_wire buffer_11023 (.in(n11023), .out(n11023_0));
mux3 mux_5858 (.in({n12399_0/**/, n12398_0, n1053}), .out(n11024), .config_in(config_chain[19619:19618]), .config_rst(config_rst)); 
buffer_wire buffer_11024 (.in(n11024), .out(n11024_0));
mux15 mux_5859 (.in({n12701_1, n12695_0, n12690_0, n12669_0, n12664_0, n12641_0, n12636_0, n12630_1, n12608_1, n11065_1, n1065, n1057, n1049, n961, n953}), .out(n11025), .config_in(config_chain[19625:19620]), .config_rst(config_rst)); 
buffer_wire buffer_11025 (.in(n11025), .out(n11025_0));
mux3 mux_5860 (.in({n12419_0, n12418_0/**/, n1057}), .out(n11026), .config_in(config_chain[19627:19626]), .config_rst(config_rst)); 
buffer_wire buffer_11026 (.in(n11026), .out(n11026_0));
mux15 mux_5861 (.in({n12957_1, n12937_0, n12932_0, n12931_0, n12926_0, n12905_0, n12900_0, n12886_1, n12864_1, n11085_1/**/, n2043, n2035, n2027, n1939, n1931}), .out(n11027), .config_in(config_chain[19633:19628]), .config_rst(config_rst)); 
buffer_wire buffer_11027 (.in(n11027), .out(n11027_0));
mux3 mux_5862 (.in({n12441_0, n12440_0/**/, n1057}), .out(n11028), .config_in(config_chain[19635:19634]), .config_rst(config_rst)); 
buffer_wire buffer_11028 (.in(n11028), .out(n11028_0));
mux13 mux_5863 (.in({n13215_1, n13208_0/**/, n13203_0, n13174_0, n13162_0, n13157_0, n13146_1, n13123_0, n11107_1, n3017, n3009, n2921, n2909}), .out(n11029), .config_in(config_chain[19641:19636]), .config_rst(config_rst)); 
buffer_wire buffer_11029 (.in(n11029), .out(n11029_0));
mux3 mux_5864 (.in({n12461_1, n12380_1, n1057}), .out(n11030), .config_in(config_chain[19643:19642]), .config_rst(config_rst)); 
buffer_wire buffer_11030 (.in(n11030), .out(n11030_0));
mux13 mux_5865 (.in({n13477_1, n13462_0, n13457_0, n13448_0, n13443_0, n13414_0, n13406_1, n13383_0, n11129_1/**/, n3995, n3987, n3899, n3887}), .out(n11031), .config_in(config_chain[19649:19644]), .config_rst(config_rst)); 
buffer_wire buffer_11031 (.in(n11031), .out(n11031_0));
mux3 mux_5866 (.in({n12401_0, n12400_0, n1057}), .out(n11032), .config_in(config_chain[19651:19650]), .config_rst(config_rst)); 
buffer_wire buffer_11032 (.in(n11032), .out(n11032_0));
mux15 mux_5867 (.in({n12699_1, n12689_0, n12684_0, n12663_0, n12658_0, n12655_0, n12650_0, n12632_1, n12610_1, n11067_1, n1065, n1057, n1049, n961/**/, n953}), .out(n11033), .config_in(config_chain[19657:19652]), .config_rst(config_rst)); 
buffer_wire buffer_11033 (.in(n11033), .out(n11033_0));
mux3 mux_5868 (.in({n12421_0, n12420_0, n1057}), .out(n11034), .config_in(config_chain[19659:19658]), .config_rst(config_rst)); 
buffer_wire buffer_11034 (.in(n11034), .out(n11034_0));
mux15 mux_5869 (.in({n12955_1, n12951_0, n12946_0, n12925_0, n12920_0, n12899_0, n12894_0, n12888_1, n12866_1, n11087_1, n2043, n2035, n2027, n1939, n1931}), .out(n11035), .config_in(config_chain[19665:19660]), .config_rst(config_rst)); 
buffer_wire buffer_11035 (.in(n11035), .out(n11035_0));
mux3 mux_5870 (.in({n12351_0, n12350_1, n1061}), .out(n11036), .config_in(config_chain[19667:19666]), .config_rst(config_rst)); 
buffer_wire buffer_11036 (.in(n11036), .out(n11036_0));
mux13 mux_5871 (.in({n13213_1, n13194_0, n13182_0, n13177_0, n13165_0, n13148_1, n13125_0, n13120_1, n11109_1, n3017, n3009, n2921/**/, n2913}), .out(n11037), .config_in(config_chain[19673:19668]), .config_rst(config_rst)); 
buffer_wire buffer_11037 (.in(n11037), .out(n11037_0));
mux3 mux_5872 (.in({n12353_1/**/, n12352_1, n1061}), .out(n11038), .config_in(config_chain[19675:19674]), .config_rst(config_rst)); 
buffer_wire buffer_11038 (.in(n11038), .out(n11038_0));
mux13 mux_5873 (.in({n13475_1, n13470_0, n13465_0, n13434_0, n13422_0, n13417_0, n13408_1, n13385_0, n11131_1, n3995, n3987/**/, n3899, n3891}), .out(n11039), .config_in(config_chain[19681:19676]), .config_rst(config_rst)); 
buffer_wire buffer_11039 (.in(n11039), .out(n11039_0));
mux3 mux_5874 (.in({n12355_1/**/, n12354_1, n1061}), .out(n11040), .config_in(config_chain[19683:19682]), .config_rst(config_rst)); 
buffer_wire buffer_11040 (.in(n11040), .out(n11040_0));
mux13 mux_5875 (.in({n13739_1, n13726_0, n13721_0, n13712_0, n13707_0, n13676_0, n13670_1, n13647_0, n11153_1, n4973, n4965, n4877, n4869}), .out(n11041), .config_in(config_chain[19689:19684]), .config_rst(config_rst)); 
buffer_wire buffer_11041 (.in(n11041), .out(n11041_0));
mux3 mux_5876 (.in({n12357_1, n12356_1, n1061}), .out(n11042), .config_in(config_chain[19691:19690]), .config_rst(config_rst)); 
buffer_wire buffer_11042 (.in(n11042), .out(n11042_0));
mux13 mux_5877 (.in({n14005_1, n14001_1, n13984_0, n13970_0, n13965_0, n13956_0, n13951_0, n13934_1, n11175_0, n5951, n5943, n5855, n5847}), .out(n11043), .config_in(config_chain[19697:19692]), .config_rst(config_rst)); 
buffer_wire buffer_11043 (.in(n11043), .out(n11043_0));
mux3 mux_5878 (.in({n12359_1, n12358_1, n1061}), .out(n11044), .config_in(config_chain[19699:19698]), .config_rst(config_rst)); 
buffer_wire buffer_11044 (.in(n11044), .out(n11044_0));
mux13 mux_5879 (.in({n14271_1, n14250_0, n14245_1, n14236_0, n14231_0, n14217_0/**/, n14200_1, n14198_1, n11197_0, n6929, n6921, n6833, n6825}), .out(n11045), .config_in(config_chain[19705:19700]), .config_rst(config_rst)); 
buffer_wire buffer_11045 (.in(n11045), .out(n11045_0));
mux3 mux_5880 (.in({n12361_1, n12360_1, n1065}), .out(n11046), .config_in(config_chain[19707:19706]), .config_rst(config_rst)); 
buffer_wire buffer_11046 (.in(n11046), .out(n11046_0));
mux13 mux_5881 (.in({n14535_1, n14525_0, n14492_0, n14487_1, n14478_0, n14473_0, n14462_1, n14432_1, n11219_0/**/, n7907, n7899, n7811, n7803}), .out(n11047), .config_in(config_chain[19713:19708]), .config_rst(config_rst)); 
buffer_wire buffer_11047 (.in(n11047), .out(n11047_0));
mux16 mux_5882 (.in({n12715_1, n12682_0, n12679_0, n12673_0, n12656_0, n12648_0, n12645_0, n12632_1, n12613_1, n12604_1, n10960_0, n2039, n2031, n1943, n1935, n1927/**/}), .out(n11048), .config_in(config_chain[19719:19714]), .config_rst(config_rst)); 
buffer_wire buffer_11048 (.in(n11048), .out(n11048_0));
mux15 mux_5883 (.in({n13737_1, n13734_0, n13729_0, n13698_0, n13693_0, n13684_0, n13679_0, n13649_0, n13644_1, n11133_1, n4973, n4965, n4877, n4869, n4861}), .out(n11049), .config_in(config_chain[19725:19720]), .config_rst(config_rst)); 
buffer_wire buffer_11049 (.in(n11049), .out(n11049_0));
mux16 mux_5884 (.in({n12697_1, n12693_0, n12676_0, n12670_0, n12667_0, n12642_0, n12639_0/**/, n12630_1, n12615_1, n12606_1, n10968_0, n2039, n2031, n1943, n1935, n1927}), .out(n11050), .config_in(config_chain[19731:19726]), .config_rst(config_rst)); 
buffer_wire buffer_11050 (.in(n11050), .out(n11050_0));
mux15 mux_5885 (.in({n13757_1, n13720_0, n13715_0, n13706_0, n13701_0, n13687_0, n13652_1, n13651_0, n13646_1, n11135_1, n4977/**/, n4965, n4877, n4869, n4861}), .out(n11051), .config_in(config_chain[19737:19732]), .config_rst(config_rst)); 
buffer_wire buffer_11051 (.in(n11051), .out(n11051_0));
mux15 mux_5886 (.in({n12699_1, n12690_0, n12687_0, n12664_0, n12661_0, n12653_0, n12636_0, n12628_1, n12608_1, n10976_0, n2039, n2031, n1943, n1935, n1927/**/}), .out(n11052), .config_in(config_chain[19743:19738]), .config_rst(config_rst)); 
buffer_wire buffer_11052 (.in(n11052), .out(n11052_0));
mux15 mux_5887 (.in({n13755_1, n13728_0, n13723_0, n13709_0, n13692_0/**/, n13678_0, n13673_0, n13654_1, n13648_1, n11137_1, n4977, n4969, n4877, n4869, n4861}), .out(n11053), .config_in(config_chain[19749:19744]), .config_rst(config_rst)); 
buffer_wire buffer_11053 (.in(n11053), .out(n11053_0));
mux15 mux_5888 (.in({n12701_1, n12684_0, n12681_0, n12675_0, n12658_0, n12650_0, n12647_0, n12626_1, n12610_1, n10984_0/**/, n2039, n2031, n1943, n1935, n1927}), .out(n11054), .config_in(config_chain[19755:19750]), .config_rst(config_rst)); 
buffer_wire buffer_11054 (.in(n11054), .out(n11054_0));
mux15 mux_5889 (.in({n13753_1, n13731_0, n13714_0/**/, n13700_0, n13695_0, n13686_0, n13681_0, n13656_1, n13650_1, n11139_1, n4977, n4969, n4961, n4869, n4861}), .out(n11055), .config_in(config_chain[19761:19756]), .config_rst(config_rst)); 
buffer_wire buffer_11055 (.in(n11055), .out(n11055_0));
mux15 mux_5890 (.in({n12703_1, n12695_0, n12678_0, n12672_0, n12669_0, n12644_0/**/, n12641_0, n12624_1, n12612_1, n10992_0, n2039, n2031, n1943, n1935, n1927}), .out(n11056), .config_in(config_chain[19767:19762]), .config_rst(config_rst)); 
buffer_wire buffer_11056 (.in(n11056), .out(n11056_0));
mux14 mux_5891 (.in({n13751_1, n13722_0, n13717_0, n13708_0, n13703_0, n13689_0, n13672_0, n13658_1, n11141_1, n4977, n4969, n4961, n4873, n4861}), .out(n11057), .config_in(config_chain[19773:19768]), .config_rst(config_rst)); 
buffer_wire buffer_11057 (.in(n11057), .out(n11057_0));
mux15 mux_5892 (.in({n12705_1, n12692_0, n12689_0, n12666_0/**/, n12663_0, n12655_0, n12638_0, n12622_1, n12614_1, n11000_0, n2043, n2035, n2027, n1939, n1931}), .out(n11058), .config_in(config_chain[19779:19774]), .config_rst(config_rst)); 
buffer_wire buffer_11058 (.in(n11058), .out(n11058_0));
mux14 mux_5893 (.in({n13749_1, n13730_0, n13725_0, n13711_0, n13694_0, n13680_0, n13675_0, n13660_1/**/, n11143_1, n4977, n4969, n4961, n4873, n4865}), .out(n11059), .config_in(config_chain[19785:19780]), .config_rst(config_rst)); 
buffer_wire buffer_11059 (.in(n11059), .out(n11059_0));
mux15 mux_5894 (.in({n12707_1, n12686_0, n12683_0, n12660_0, n12657_0/**/, n12652_0, n12649_0, n12620_1, n12605_0, n11008_0, n2043, n2035, n2027, n1939, n1931}), .out(n11060), .config_in(config_chain[19791:19786]), .config_rst(config_rst)); 
buffer_wire buffer_11060 (.in(n11060), .out(n11060_0));
mux13 mux_5895 (.in({n13747_1, n13733_0, n13716_0, n13702_0, n13697_0, n13688_0, n13683_0, n13662_1/**/, n11145_1, n4969, n4961, n4873, n4865}), .out(n11061), .config_in(config_chain[19797:19792]), .config_rst(config_rst)); 
buffer_wire buffer_11061 (.in(n11061), .out(n11061_0));
mux15 mux_5896 (.in({n12709_1, n12680_0, n12677_0, n12674_0/**/, n12671_0, n12646_0, n12643_0, n12618_1, n12607_0, n11016_0, n2043, n2035, n2027, n1939, n1931}), .out(n11062), .config_in(config_chain[19803:19798]), .config_rst(config_rst)); 
buffer_wire buffer_11062 (.in(n11062), .out(n11062_0));
mux13 mux_5897 (.in({n13745_1, n13724_0, n13719_0, n13710_0, n13705_0, n13691_0, n13674_0, n13664_1, n11147_1, n4973/**/, n4961, n4873, n4865}), .out(n11063), .config_in(config_chain[19809:19804]), .config_rst(config_rst)); 
buffer_wire buffer_11063 (.in(n11063), .out(n11063_0));
mux15 mux_5898 (.in({n12711_1, n12694_0, n12691_0, n12668_0, n12665_0, n12640_0, n12637_0, n12616_1, n12609_1, n11024_0, n2043, n2035/**/, n2027, n1939, n1931}), .out(n11064), .config_in(config_chain[19815:19810]), .config_rst(config_rst)); 
buffer_wire buffer_11064 (.in(n11064), .out(n11064_0));
mux13 mux_5899 (.in({n13743_1, n13732_0, n13727_0, n13713_1, n13696_0, n13682_0, n13677_0, n13666_1, n11149_1, n4973, n4965, n4873, n4865}), .out(n11065), .config_in(config_chain[19821:19816]), .config_rst(config_rst)); 
buffer_wire buffer_11065 (.in(n11065), .out(n11065_0));
mux15 mux_5900 (.in({n12713_1, n12688_0, n12685_0/**/, n12662_0, n12659_0, n12654_0, n12651_0, n12634_1, n12611_1, n11032_0, n2043, n2035, n2027, n1939, n1931}), .out(n11066), .config_in(config_chain[19827:19822]), .config_rst(config_rst)); 
buffer_wire buffer_11066 (.in(n11066), .out(n11066_0));
mux13 mux_5901 (.in({n13741_1, n13735_1, n13718_0, n13704_0, n13699_0, n13690_0, n13685_0/**/, n13668_1, n11151_1, n4973, n4965, n4877, n4865}), .out(n11067), .config_in(config_chain[19833:19828]), .config_rst(config_rst)); 
buffer_wire buffer_11067 (.in(n11067), .out(n11067_0));
mux16 mux_5902 (.in({n12971_1, n12944_0, n12941_0, n12918_0, n12915_0, n12909_0, n12892_0, n12888_1, n12869_1, n12860_1, n10962_0, n3017/**/, n3009, n2921, n2913, n2905}), .out(n11068), .config_in(config_chain[19839:19834]), .config_rst(config_rst)); 
buffer_wire buffer_11068 (.in(n11068), .out(n11068_0));
mux15 mux_5903 (.in({n14003_1/**/, n13992_0, n13987_0, n13978_0, n13973_0, n13942_0, n13937_0, n13913_0, n13910_1, n11155_0, n5951, n5943, n5855, n5847, n5839}), .out(n11069), .config_in(config_chain[19845:19840]), .config_rst(config_rst)); 
buffer_wire buffer_11069 (.in(n11069), .out(n11069_0));
mux16 mux_5904 (.in({n12953_1, n12938_0, n12935_0/**/, n12929_0, n12912_0, n12906_0, n12903_0, n12886_1, n12871_1, n12862_1, n10970_0, n3017, n3009, n2921, n2913, n2905}), .out(n11070), .config_in(config_chain[19851:19846]), .config_rst(config_rst)); 
buffer_wire buffer_11070 (.in(n11070), .out(n11070_0));
mux15 mux_5905 (.in({n14023_1, n14000_0, n13995_0, n13964_0, n13959_0/**/, n13950_0, n13945_0, n13916_1, n13915_0, n11157_0, n5955, n5943, n5855, n5847, n5839}), .out(n11071), .config_in(config_chain[19857:19852]), .config_rst(config_rst)); 
buffer_wire buffer_11071 (.in(n11071), .out(n11071_0));
mux15 mux_5906 (.in({n12955_1, n12949_0, n12932_0, n12926_0, n12923_0, n12900_0, n12897_0/**/, n12884_1, n12864_1, n10978_0, n3017, n3009, n2921, n2913, n2905}), .out(n11072), .config_in(config_chain[19863:19858]), .config_rst(config_rst)); 
buffer_wire buffer_11072 (.in(n11072), .out(n11072_0));
mux15 mux_5907 (.in({n14021_1, n13986_0, n13981_0, n13972_0, n13967_0/**/, n13953_0, n13936_0, n13918_1, n13912_1, n11159_0, n5955, n5947, n5855, n5847, n5839}), .out(n11073), .config_in(config_chain[19869:19864]), .config_rst(config_rst)); 
buffer_wire buffer_11073 (.in(n11073), .out(n11073_0));
mux15 mux_5908 (.in({n12957_1, n12946_0, n12943_0, n12920_0, n12917_0, n12911_0, n12894_0, n12882_1, n12866_1, n10986_0, n3017, n3009, n2921, n2913/**/, n2905}), .out(n11074), .config_in(config_chain[19875:19870]), .config_rst(config_rst)); 
buffer_wire buffer_11074 (.in(n11074), .out(n11074_0));
mux15 mux_5909 (.in({n14019_1, n13994_0, n13989_0, n13975_0, n13958_0, n13944_0, n13939_0, n13920_1, n13914_1, n11161_0, n5955, n5947, n5939/**/, n5847, n5839}), .out(n11075), .config_in(config_chain[19881:19876]), .config_rst(config_rst)); 
buffer_wire buffer_11075 (.in(n11075), .out(n11075_0));
mux15 mux_5910 (.in({n12959_1, n12940_0, n12937_0, n12931_0, n12914_0, n12908_0, n12905_0, n12880_1/**/, n12868_1, n10994_0, n3017, n3009, n2921, n2913, n2905}), .out(n11076), .config_in(config_chain[19887:19882]), .config_rst(config_rst)); 
buffer_wire buffer_11076 (.in(n11076), .out(n11076_0));
mux14 mux_5911 (.in({n14017_1, n13997_0, n13980_0, n13966_0, n13961_0, n13952_0, n13947_0, n13922_1, n11163_0, n5955, n5947/**/, n5939, n5851, n5839}), .out(n11077), .config_in(config_chain[19893:19888]), .config_rst(config_rst)); 
buffer_wire buffer_11077 (.in(n11077), .out(n11077_0));
mux15 mux_5912 (.in({n12961_1, n12951_0, n12934_0, n12928_0, n12925_0, n12902_0, n12899_0, n12878_1, n12870_1, n11002_0/**/, n3021, n3013, n3005, n2917, n2909}), .out(n11078), .config_in(config_chain[19899:19894]), .config_rst(config_rst)); 
buffer_wire buffer_11078 (.in(n11078), .out(n11078_0));
mux14 mux_5913 (.in({n14015_1, n13988_0, n13983_0, n13974_0, n13969_0, n13955_0, n13938_0, n13924_1, n11165_0, n5955, n5947, n5939/**/, n5851, n5843}), .out(n11079), .config_in(config_chain[19905:19900]), .config_rst(config_rst)); 
buffer_wire buffer_11079 (.in(n11079), .out(n11079_0));
mux15 mux_5914 (.in({n12963_1, n12948_0/**/, n12945_0, n12922_0, n12919_0, n12896_0, n12893_0, n12876_1, n12861_0, n11010_0, n3021, n3013, n3005, n2917, n2909}), .out(n11080), .config_in(config_chain[19911:19906]), .config_rst(config_rst)); 
buffer_wire buffer_11080 (.in(n11080), .out(n11080_0));
mux13 mux_5915 (.in({n14013_1, n13996_0, n13991_0, n13977_0, n13960_0/**/, n13946_0, n13941_0, n13926_1, n11167_0, n5947, n5939, n5851, n5843}), .out(n11081), .config_in(config_chain[19917:19912]), .config_rst(config_rst)); 
buffer_wire buffer_11081 (.in(n11081), .out(n11081_0));
mux15 mux_5916 (.in({n12965_1, n12942_0, n12939_0/**/, n12916_0, n12913_0, n12910_0, n12907_0, n12874_1, n12863_0, n11018_0, n3021, n3013, n3005, n2917, n2909}), .out(n11082), .config_in(config_chain[19923:19918]), .config_rst(config_rst)); 
buffer_wire buffer_11082 (.in(n11082), .out(n11082_0));
mux13 mux_5917 (.in({n14011_1, n13999_0, n13982_0, n13968_0, n13963_0, n13954_0, n13949_0, n13928_1, n11169_0, n5951, n5939/**/, n5851, n5843}), .out(n11083), .config_in(config_chain[19929:19924]), .config_rst(config_rst)); 
buffer_wire buffer_11083 (.in(n11083), .out(n11083_0));
mux15 mux_5918 (.in({n12967_1, n12936_0, n12933_0, n12930_0, n12927_0, n12904_0, n12901_0, n12872_1, n12865_0, n11026_0/**/, n3021, n3013, n3005, n2917, n2909}), .out(n11084), .config_in(config_chain[19935:19930]), .config_rst(config_rst)); 
buffer_wire buffer_11084 (.in(n11084), .out(n11084_0));
mux13 mux_5919 (.in({n14009_1, n13990_0, n13985_0, n13976_0, n13971_0/**/, n13957_1, n13940_0, n13930_1, n11171_0, n5951, n5943, n5851, n5843}), .out(n11085), .config_in(config_chain[19941:19936]), .config_rst(config_rst)); 
buffer_wire buffer_11085 (.in(n11085), .out(n11085_0));
mux15 mux_5920 (.in({n12969_1, n12950_0, n12947_0, n12924_0, n12921_0/**/, n12898_0, n12895_0, n12890_1, n12867_1, n11034_0, n3021, n3013, n3005, n2917, n2909}), .out(n11086), .config_in(config_chain[19947:19942]), .config_rst(config_rst)); 
buffer_wire buffer_11086 (.in(n11086), .out(n11086_0));
mux13 mux_5921 (.in({n14007_1/**/, n13998_0, n13993_0, n13979_1, n13962_0, n13948_0, n13943_0, n13932_1, n11173_0, n5951, n5943, n5855, n5843}), .out(n11087), .config_in(config_chain[19953:19948]), .config_rst(config_rst)); 
buffer_wire buffer_11087 (.in(n11087), .out(n11087_0));
mux15 mux_5922 (.in({n13231_1, n13203_0, n13196_0, n13184_0, n13157_0, n13150_0, n13148_1, n13126_1, n13123_0, n10956_0/**/, n3995, n3987, n3899, n3891, n3883}), .out(n11088), .config_in(config_chain[19959:19954]), .config_rst(config_rst)); 
buffer_wire buffer_11088 (.in(n11088), .out(n11088_0));
mux15 mux_5923 (.in({n14269_1, n14267_1, n14258_0, n14253_0, n14239_0, n14222_0, n14208_0, n14203_0/**/, n14176_1, n11177_0, n6929, n6921, n6833, n6825, n6817}), .out(n11089), .config_in(config_chain[19965:19960]), .config_rst(config_rst)); 
buffer_wire buffer_11089 (.in(n11089), .out(n11089_0));
mux15 mux_5924 (.in({n13211_1, n13204_0, n13177_0, n13170_0, n13165_0, n13158_0, n13146_1/**/, n13128_1, n13125_0, n10964_0, n3999, n3987, n3899, n3891, n3883}), .out(n11090), .config_in(config_chain[19971:19966]), .config_rst(config_rst)); 
buffer_wire buffer_11090 (.in(n11090), .out(n11090_0));
mux15 mux_5925 (.in({n14289_1, n14261_0, n14244_0, n14230_0, n14225_0, n14216_0, n14211_0, n14180_1, n14179_0, n11179_0, n6933, n6921, n6833, n6825, n6817}), .out(n11091), .config_in(config_chain[19977:19972]), .config_rst(config_rst)); 
buffer_wire buffer_11091 (.in(n11091), .out(n11091_0));
mux15 mux_5926 (.in({n13213_1, n13197_0, n13190_0, n13185_0, n13178_0, n13166_0, n13151_0, n13144_1/**/, n13127_1, n10972_0, n3999, n3991, n3899, n3891, n3883}), .out(n11092), .config_in(config_chain[19983:19978]), .config_rst(config_rst)); 
buffer_wire buffer_11092 (.in(n11092), .out(n11092_0));
mux15 mux_5927 (.in({n14287_1, n14266_0, n14252_0, n14247_0, n14238_0, n14233_0/**/, n14219_0, n14202_0, n14182_1, n11181_0, n6933, n6925, n6833, n6825, n6817}), .out(n11093), .config_in(config_chain[19989:19984]), .config_rst(config_rst)); 
buffer_wire buffer_11093 (.in(n11093), .out(n11093_0));
mux15 mux_5928 (.in({n13215_1, n13205_0, n13198_0, n13186_0/**/, n13171_0, n13159_0, n13152_0, n13142_1, n13129_1, n10980_0, n3999, n3991, n3983, n3891, n3883}), .out(n11094), .config_in(config_chain[19995:19990]), .config_rst(config_rst)); 
buffer_wire buffer_11094 (.in(n11094), .out(n11094_0));
mux15 mux_5929 (.in({n14285_1, n14260_0/**/, n14255_0, n14241_0, n14224_0, n14210_0, n14205_0, n14184_1, n14178_1, n11183_0, n6933, n6925, n6917, n6825, n6817}), .out(n11095), .config_in(config_chain[20001:19996]), .config_rst(config_rst)); 
buffer_wire buffer_11095 (.in(n11095), .out(n11095_0));
mux14 mux_5930 (.in({n13217_1, n13206_0, n13191_0, n13179_0, n13172_0, n13167_0, n13160_0, n13140_1, n10988_0, n3999, n3991, n3983/**/, n3895, n3883}), .out(n11096), .config_in(config_chain[20007:20002]), .config_rst(config_rst)); 
buffer_wire buffer_11096 (.in(n11096), .out(n11096_0));
mux14 mux_5931 (.in({n14283_1, n14263_0, n14246_0, n14232_0, n14227_0, n14218_0, n14213_0, n14186_1, n11185_0, n6933/**/, n6925, n6917, n6829, n6817}), .out(n11097), .config_in(config_chain[20013:20008]), .config_rst(config_rst)); 
buffer_wire buffer_11097 (.in(n11097), .out(n11097_0));
mux14 mux_5932 (.in({n13219_1, n13199_0, n13192_0/**/, n13187_0, n13180_0, n13168_0, n13153_0, n13138_1, n10996_0, n3999, n3991, n3983, n3895, n3887}), .out(n11098), .config_in(config_chain[20019:20014]), .config_rst(config_rst)); 
buffer_wire buffer_11098 (.in(n11098), .out(n11098_0));
mux14 mux_5933 (.in({n14281_1, n14254_0, n14249_0, n14240_0, n14235_0, n14221_0, n14204_0, n14188_1, n11187_0, n6933, n6925, n6917, n6829, n6821/**/}), .out(n11099), .config_in(config_chain[20025:20020]), .config_rst(config_rst)); 
buffer_wire buffer_11099 (.in(n11099), .out(n11099_0));
mux13 mux_5934 (.in({n13221_1, n13207_0, n13200_0, n13188_0, n13173_0, n13161_0, n13154_0, n13136_1, n11004_0, n3991, n3983, n3895, n3887/**/}), .out(n11100), .config_in(config_chain[20031:20026]), .config_rst(config_rst)); 
buffer_wire buffer_11100 (.in(n11100), .out(n11100_0));
mux13 mux_5935 (.in({n14279_1, n14262_0, n14257_0, n14243_0/**/, n14226_0, n14212_0, n14207_0, n14190_1, n11189_0, n6925, n6917, n6829, n6821}), .out(n11101), .config_in(config_chain[20037:20032]), .config_rst(config_rst)); 
buffer_wire buffer_11101 (.in(n11101), .out(n11101_0));
mux13 mux_5936 (.in({n13223_1/**/, n13208_0, n13193_0, n13181_0, n13174_0, n13169_0, n13162_0, n13134_1, n11012_0, n3995, n3983, n3895, n3887}), .out(n11102), .config_in(config_chain[20043:20038]), .config_rst(config_rst)); 
buffer_wire buffer_11102 (.in(n11102), .out(n11102_0));
mux13 mux_5937 (.in({n14277_1, n14265_0, n14248_0, n14234_0, n14229_0, n14220_0, n14215_0, n14192_1, n11191_0, n6929, n6917/**/, n6829, n6821}), .out(n11103), .config_in(config_chain[20049:20044]), .config_rst(config_rst)); 
buffer_wire buffer_11103 (.in(n11103), .out(n11103_0));
mux13 mux_5938 (.in({n13225_1, n13201_0, n13194_0, n13189_0, n13182_0, n13155_0, n13132_1, n13120_1, n11020_0/**/, n3995, n3987, n3895, n3887}), .out(n11104), .config_in(config_chain[20055:20050]), .config_rst(config_rst)); 
buffer_wire buffer_11104 (.in(n11104), .out(n11104_0));
mux13 mux_5939 (.in({n14275_1, n14256_0, n14251_0, n14242_0, n14237_0, n14206_0, n14201_1, n14194_1, n11193_0, n6929, n6921, n6829/**/, n6821}), .out(n11105), .config_in(config_chain[20061:20056]), .config_rst(config_rst)); 
buffer_wire buffer_11105 (.in(n11105), .out(n11105_0));
mux13 mux_5940 (.in({n13227_1, n13209_0, n13202_0, n13175_0, n13163_0, n13156_0, n13130_1, n13122_1, n11028_0/**/, n3995, n3987, n3899, n3887}), .out(n11106), .config_in(config_chain[20067:20062]), .config_rst(config_rst)); 
buffer_wire buffer_11106 (.in(n11106), .out(n11106_0));
mux13 mux_5941 (.in({n14273_1, n14264_0, n14259_0, n14228_0, n14223_1, n14214_0/**/, n14209_0, n14196_1, n11195_0, n6929, n6921, n6833, n6821}), .out(n11107), .config_in(config_chain[20073:20068]), .config_rst(config_rst)); 
buffer_wire buffer_11107 (.in(n11107), .out(n11107_0));
mux13 mux_5942 (.in({n13229_1, n13195_0, n13183_0, n13176_0, n13164_0, n13124_1, n13121_0, n13118_1, n11036_0, n3995, n3987/**/, n3899, n3891}), .out(n11108), .config_in(config_chain[20079:20074]), .config_rst(config_rst)); 
buffer_wire buffer_11108 (.in(n11108), .out(n11108_0));
mux3 mux_5943 (.in({n14695_1, n14694_1, n8885}), .out(n11109), .config_in(config_chain[20081:20080]), .config_rst(config_rst)); 
buffer_wire buffer_11109 (.in(n11109), .out(n11109_0));
mux15 mux_5944 (.in({n13493_1, n13457_0, n13450_0, n13443_0, n13436_0, n13424_0, n13408_1, n13386_1/**/, n13383_0, n10958_1, n4973, n4965, n4877, n4869, n4861}), .out(n11110), .config_in(config_chain[20087:20082]), .config_rst(config_rst)); 
buffer_wire buffer_11110 (.in(n11110), .out(n11110_0));
mux15 mux_5945 (.in({n14533_1, n14516_0, n14511_0, n14509_1, n14500_0, n14495_0, n14481_0, n14464_1, n14442_1, n11199_0/**/, n7907, n7899, n7811, n7803, n7795}), .out(n11111), .config_in(config_chain[20093:20088]), .config_rst(config_rst)); 
buffer_wire buffer_11111 (.in(n11111), .out(n11111_0));
mux15 mux_5946 (.in({n13473_1, n13465_0, n13458_0, n13444_0, n13417_0, n13410_0/**/, n13406_1, n13388_1, n13385_0, n10966_1, n4977, n4965, n4877, n4869, n4861}), .out(n11112), .config_in(config_chain[20099:20094]), .config_rst(config_rst)); 
buffer_wire buffer_11112 (.in(n11112), .out(n11112_0));
mux15 mux_5947 (.in({n14553_1, n14531_1, n14524_0/**/, n14519_0, n14503_0, n14486_0, n14472_0, n14467_0, n14444_1, n11201_0, n7911, n7899, n7811, n7803, n7795}), .out(n11113), .config_in(config_chain[20105:20100]), .config_rst(config_rst)); 
buffer_wire buffer_11113 (.in(n11113), .out(n11113_0));
mux15 mux_5948 (.in({n13475_1, n13466_0, n13451_0, n13437_0, n13430_0/**/, n13425_0, n13418_0, n13404_1, n13387_0, n10974_1, n4977, n4969, n4877, n4869, n4861}), .out(n11114), .config_in(config_chain[20111:20106]), .config_rst(config_rst)); 
buffer_wire buffer_11114 (.in(n11114), .out(n11114_0));
mux15 mux_5949 (.in({n14551_1, n14527_0, n14510_0, n14508_0, n14494_0, n14489_0, n14480_0, n14475_0, n14446_1, n11203_0, n7911, n7903/**/, n7811, n7803, n7795}), .out(n11115), .config_in(config_chain[20117:20112]), .config_rst(config_rst)); 
buffer_wire buffer_11115 (.in(n11115), .out(n11115_0));
mux15 mux_5950 (.in({n13477_1, n13459_0, n13452_0, n13445_0, n13438_0, n13426_0, n13411_0/**/, n13402_1, n13389_1, n10982_1, n4977, n4969, n4961, n4869, n4861}), .out(n11116), .config_in(config_chain[20123:20118]), .config_rst(config_rst)); 
buffer_wire buffer_11116 (.in(n11116), .out(n11116_0));
mux15 mux_5951 (.in({n14549_1, n14530_0, n14518_0, n14513_0, n14502_0, n14497_0/**/, n14483_0, n14466_0, n14448_1, n11205_0, n7911, n7903, n7895, n7803, n7795}), .out(n11117), .config_in(config_chain[20129:20124]), .config_rst(config_rst)); 
buffer_wire buffer_11117 (.in(n11117), .out(n11117_0));
mux14 mux_5952 (.in({n13479_1, n13467_0, n13460_0, n13446_0, n13431_0, n13419_0, n13412_0, n13400_1, n10990_1, n4977, n4969/**/, n4961, n4873, n4861}), .out(n11118), .config_in(config_chain[20135:20130]), .config_rst(config_rst)); 
buffer_wire buffer_11118 (.in(n11118), .out(n11118_0));
mux14 mux_5953 (.in({n14547_1, n14526_0, n14521_0, n14505_0/**/, n14488_0, n14474_0, n14469_0, n14450_1, n11207_0, n7911, n7903, n7895, n7807, n7795}), .out(n11119), .config_in(config_chain[20141:20136]), .config_rst(config_rst)); 
buffer_wire buffer_11119 (.in(n11119), .out(n11119_0));
mux14 mux_5954 (.in({n13481_1, n13468_0, n13453_0, n13439_0, n13432_0, n13427_0, n13420_0, n13398_1, n10998_1/**/, n4977, n4969, n4961, n4873, n4865}), .out(n11120), .config_in(config_chain[20147:20142]), .config_rst(config_rst)); 
buffer_wire buffer_11120 (.in(n11120), .out(n11120_0));
mux14 mux_5955 (.in({n14545_1, n14529_0, n14512_0, n14496_0, n14491_0, n14482_0, n14477_0, n14452_1, n11209_0, n7911, n7903/**/, n7895, n7807, n7799}), .out(n11121), .config_in(config_chain[20153:20148]), .config_rst(config_rst)); 
buffer_wire buffer_11121 (.in(n11121), .out(n11121_0));
mux13 mux_5956 (.in({n13483_1, n13461_0, n13454_0, n13447_0, n13440_0, n13428_0, n13413_0, n13396_1/**/, n11006_1, n4969, n4961, n4873, n4865}), .out(n11122), .config_in(config_chain[20159:20154]), .config_rst(config_rst)); 
buffer_wire buffer_11122 (.in(n11122), .out(n11122_0));
mux13 mux_5957 (.in({n14543_1, n14520_0, n14515_0, n14504_0, n14499_0, n14485_0, n14468_0/**/, n14454_1, n11211_0, n7903, n7895, n7807, n7799}), .out(n11123), .config_in(config_chain[20165:20160]), .config_rst(config_rst)); 
buffer_wire buffer_11123 (.in(n11123), .out(n11123_0));
mux13 mux_5958 (.in({n13485_1, n13469_0, n13462_0, n13448_0, n13433_0/**/, n13421_0, n13414_0, n13394_1, n11014_1, n4973, n4961, n4873, n4865}), .out(n11124), .config_in(config_chain[20171:20166]), .config_rst(config_rst)); 
buffer_wire buffer_11124 (.in(n11124), .out(n11124_0));
mux13 mux_5959 (.in({n14541_1/**/, n14528_0, n14523_0, n14507_0, n14490_0, n14476_0, n14471_0, n14456_1, n11213_0, n7907, n7895, n7807, n7799}), .out(n11125), .config_in(config_chain[20177:20172]), .config_rst(config_rst)); 
buffer_wire buffer_11125 (.in(n11125), .out(n11125_0));
mux13 mux_5960 (.in({n13487_1, n13470_0, n13455_0, n13441_0, n13434_0, n13429_0, n13422_0, n13392_1/**/, n11022_1, n4973, n4965, n4873, n4865}), .out(n11126), .config_in(config_chain[20183:20178]), .config_rst(config_rst)); 
buffer_wire buffer_11126 (.in(n11126), .out(n11126_0));
mux13 mux_5961 (.in({n14539_1, n14514_0, n14498_0, n14493_0, n14484_0, n14479_0, n14458_1, n14433_1, n11215_0/**/, n7907, n7899, n7807, n7799}), .out(n11127), .config_in(config_chain[20189:20184]), .config_rst(config_rst)); 
buffer_wire buffer_11127 (.in(n11127), .out(n11127_0));
mux13 mux_5962 (.in({n13489_1, n13463_0, n13456_0, n13449_0, n13442_0, n13415_0, n13390_1/**/, n13382_1, n11030_1, n4973, n4965, n4877, n4865}), .out(n11128), .config_in(config_chain[20195:20190]), .config_rst(config_rst)); 
buffer_wire buffer_11128 (.in(n11128), .out(n11128_0));
mux13 mux_5963 (.in({n14537_1, n14522_0, n14517_0, n14506_0, n14501_0, n14470_0, n14465_1, n14460_1, n11217_0, n7907/**/, n7899, n7811, n7799}), .out(n11129), .config_in(config_chain[20201:20196]), .config_rst(config_rst)); 
buffer_wire buffer_11129 (.in(n11129), .out(n11129_0));
mux13 mux_5964 (.in({n13491_1, n13471_1, n13464_0, n13435_0/**/, n13423_0, n13416_0, n13384_1, n13380_1, n11038_1, n4973, n4965, n4877, n4869}), .out(n11130), .config_in(config_chain[20207:20202]), .config_rst(config_rst)); 
buffer_wire buffer_11130 (.in(n11130), .out(n11130_0));
mux3 mux_5965 (.in({n14697_1, n14696_1, n8885}), .out(n11131), .config_in(config_chain[20209:20208]), .config_rst(config_rst)); 
buffer_wire buffer_11131 (.in(n11131), .out(n11131_0));
mux15 mux_5966 (.in({n13757_1, n13735_1, n13728_0, n13699_0, n13692_0, n13685_0, n13678_0, n13670_1, n13648_1, n11048_1, n5951, n5943, n5855, n5847, n5839}), .out(n11132), .config_in(config_chain[20215:20210]), .config_rst(config_rst)); 
buffer_wire buffer_11132 (.in(n11132), .out(n11132_0));
mux4 mux_5967 (.in({n14795_1, n14706_1, n8889, n8773}), .out(n11133), .config_in(config_chain[20217:20216]), .config_rst(config_rst)); 
buffer_wire buffer_11133 (.in(n11133), .out(n11133_0));
mux15 mux_5968 (.in({n13737_1, n13721_0/**/, n13714_0, n13707_0, n13700_0, n13686_0, n13668_1, n13650_1, n13647_0, n11050_1, n5955, n5943, n5855, n5847, n5839}), .out(n11134), .config_in(config_chain[20223:20218]), .config_rst(config_rst)); 
buffer_wire buffer_11134 (.in(n11134), .out(n11134_0));
mux3 mux_5969 (.in({n14797_1, n14708_1/**/, n8777}), .out(n11135), .config_in(config_chain[20225:20224]), .config_rst(config_rst)); 
buffer_wire buffer_11135 (.in(n11135), .out(n11135_0));
mux15 mux_5970 (.in({n13739_1, n13729_0, n13722_0, n13708_0, n13693_0, n13679_0, n13672_0, n13666_1/**/, n13649_0, n11052_1, n5955, n5947, n5855, n5847, n5839}), .out(n11136), .config_in(config_chain[20231:20226]), .config_rst(config_rst)); 
buffer_wire buffer_11136 (.in(n11136), .out(n11136_0));
mux3 mux_5971 (.in({n14799_1, n14710_1/**/, n8781}), .out(n11137), .config_in(config_chain[20233:20232]), .config_rst(config_rst)); 
buffer_wire buffer_11137 (.in(n11137), .out(n11137_0));
mux15 mux_5972 (.in({n13741_1, n13730_0, n13715_0, n13701_0, n13694_0, n13687_0/**/, n13680_0, n13664_1, n13651_0, n11054_1, n5955, n5947, n5939, n5847, n5839}), .out(n11138), .config_in(config_chain[20239:20234]), .config_rst(config_rst)); 
buffer_wire buffer_11138 (.in(n11138), .out(n11138_0));
mux3 mux_5973 (.in({n14801_1, n14712_1, n8781}), .out(n11139), .config_in(config_chain[20241:20240]), .config_rst(config_rst)); 
buffer_wire buffer_11139 (.in(n11139), .out(n11139_0));
mux14 mux_5974 (.in({n13743_1, n13723_0, n13716_0, n13709_0, n13702_0, n13688_0, n13673_0/**/, n13662_1, n11056_1, n5955, n5947, n5939, n5851, n5839}), .out(n11140), .config_in(config_chain[20247:20242]), .config_rst(config_rst)); 
buffer_wire buffer_11140 (.in(n11140), .out(n11140_0));
mux3 mux_5975 (.in({n14803_1, n14714_1, n8785}), .out(n11141), .config_in(config_chain[20249:20248]), .config_rst(config_rst)); 
buffer_wire buffer_11141 (.in(n11141), .out(n11141_0));
mux14 mux_5976 (.in({n13745_1, n13731_0/**/, n13724_0, n13710_0, n13695_0, n13681_0, n13674_0, n13660_1, n11058_1, n5955, n5947, n5939, n5851, n5843}), .out(n11142), .config_in(config_chain[20255:20250]), .config_rst(config_rst)); 
buffer_wire buffer_11142 (.in(n11142), .out(n11142_0));
mux3 mux_5977 (.in({n14805_1, n14716_1, n8789}), .out(n11143), .config_in(config_chain[20257:20256]), .config_rst(config_rst)); 
buffer_wire buffer_11143 (.in(n11143), .out(n11143_0));
mux13 mux_5978 (.in({n13747_1, n13732_0, n13717_0, n13703_0, n13696_0, n13689_0, n13682_0/**/, n13658_1, n11060_1, n5947, n5939, n5851, n5843}), .out(n11144), .config_in(config_chain[20263:20258]), .config_rst(config_rst)); 
buffer_wire buffer_11144 (.in(n11144), .out(n11144_0));
mux3 mux_5979 (.in({n14807_1, n14718_1/**/, n8873}), .out(n11145), .config_in(config_chain[20265:20264]), .config_rst(config_rst)); 
buffer_wire buffer_11145 (.in(n11145), .out(n11145_0));
mux13 mux_5980 (.in({n13749_1, n13725_0, n13718_0, n13711_0, n13704_0, n13690_0, n13675_0, n13656_1, n11062_1/**/, n5951, n5939, n5851, n5843}), .out(n11146), .config_in(config_chain[20271:20266]), .config_rst(config_rst)); 
buffer_wire buffer_11146 (.in(n11146), .out(n11146_0));
mux3 mux_5981 (.in({n14809_1, n14720_1, n8877}), .out(n11147), .config_in(config_chain[20273:20272]), .config_rst(config_rst)); 
buffer_wire buffer_11147 (.in(n11147), .out(n11147_0));
mux13 mux_5982 (.in({n13751_1, n13733_0, n13726_0, n13712_0, n13697_0, n13683_0, n13676_0, n13654_1, n11064_1/**/, n5951, n5943, n5851, n5843}), .out(n11148), .config_in(config_chain[20279:20274]), .config_rst(config_rst)); 
buffer_wire buffer_11148 (.in(n11148), .out(n11148_0));
mux3 mux_5983 (.in({n14811_1, n14722_1/**/, n8877}), .out(n11149), .config_in(config_chain[20281:20280]), .config_rst(config_rst)); 
buffer_wire buffer_11149 (.in(n11149), .out(n11149_0));
mux13 mux_5984 (.in({n13753_1, n13734_0, n13719_0, n13705_0, n13698_0, n13691_0, n13684_0/**/, n13652_1, n11066_1, n5951, n5943, n5855, n5843}), .out(n11150), .config_in(config_chain[20287:20282]), .config_rst(config_rst)); 
buffer_wire buffer_11150 (.in(n11150), .out(n11150_0));
mux3 mux_5985 (.in({n14813_1, n14724_1/**/, n8881}), .out(n11151), .config_in(config_chain[20289:20288]), .config_rst(config_rst)); 
buffer_wire buffer_11151 (.in(n11151), .out(n11151_0));
mux13 mux_5986 (.in({n13755_1, n13727_0/**/, n13720_0, n13713_1, n13706_0, n13677_0, n13646_1, n13644_1, n11040_1, n5951, n5943, n5855, n5847}), .out(n11152), .config_in(config_chain[20295:20290]), .config_rst(config_rst)); 
buffer_wire buffer_11152 (.in(n11152), .out(n11152_0));
mux3 mux_5987 (.in({n14727_1, n14726_1, n8885}), .out(n11153), .config_in(config_chain[20297:20296]), .config_rst(config_rst)); 
buffer_wire buffer_11153 (.in(n11153), .out(n11153_0));
mux15 mux_5988 (.in({n14023_1, n13993_0, n13986_0, n13979_1, n13972_0, n13943_0, n13936_0, n13934_1, n13912_1, n11068_1, n6929/**/, n6921, n6833, n6825, n6817}), .out(n11154), .config_in(config_chain[20303:20298]), .config_rst(config_rst)); 
buffer_wire buffer_11154 (.in(n11154), .out(n11154_0));
mux4 mux_5989 (.in({n14729_0, n14728_0, n8889, n8773}), .out(n11155), .config_in(config_chain[20305:20304]), .config_rst(config_rst)); 
buffer_wire buffer_11155 (.in(n11155), .out(n11155_0));
mux15 mux_5990 (.in({n14003_1, n14001_1, n13994_0, n13965_0, n13958_0, n13951_0/**/, n13944_0, n13932_1, n13914_1, n11070_1, n6933, n6921, n6833, n6825, n6817}), .out(n11156), .config_in(config_chain[20311:20306]), .config_rst(config_rst)); 
buffer_wire buffer_11156 (.in(n11156), .out(n11156_0));
mux3 mux_5991 (.in({n14731_0/**/, n14730_0, n8777}), .out(n11157), .config_in(config_chain[20313:20312]), .config_rst(config_rst)); 
buffer_wire buffer_11157 (.in(n11157), .out(n11157_0));
mux15 mux_5992 (.in({n14005_1/**/, n13987_0, n13980_0, n13973_0, n13966_0, n13952_0, n13937_0, n13930_1, n13913_0, n11072_1, n6933, n6925, n6833, n6825, n6817}), .out(n11158), .config_in(config_chain[20319:20314]), .config_rst(config_rst)); 
buffer_wire buffer_11158 (.in(n11158), .out(n11158_0));
mux3 mux_5993 (.in({n14733_0, n14732_0, n8781}), .out(n11159), .config_in(config_chain[20321:20320]), .config_rst(config_rst)); 
buffer_wire buffer_11159 (.in(n11159), .out(n11159_0));
mux15 mux_5994 (.in({n14007_1/**/, n13995_0, n13988_0, n13974_0, n13959_0, n13945_0, n13938_0, n13928_1, n13915_0, n11074_1, n6933, n6925, n6917, n6825, n6817}), .out(n11160), .config_in(config_chain[20327:20322]), .config_rst(config_rst)); 
buffer_wire buffer_11160 (.in(n11160), .out(n11160_0));
mux3 mux_5995 (.in({n14735_0/**/, n14734_0, n8785}), .out(n11161), .config_in(config_chain[20329:20328]), .config_rst(config_rst)); 
buffer_wire buffer_11161 (.in(n11161), .out(n11161_0));
mux14 mux_5996 (.in({n14009_1, n13996_0, n13981_0, n13967_0, n13960_0, n13953_0, n13946_0, n13926_1, n11076_1, n6933, n6925, n6917/**/, n6829, n6817}), .out(n11162), .config_in(config_chain[20335:20330]), .config_rst(config_rst)); 
buffer_wire buffer_11162 (.in(n11162), .out(n11162_0));
mux3 mux_5997 (.in({n14737_0, n14736_0, n8785}), .out(n11163), .config_in(config_chain[20337:20336]), .config_rst(config_rst)); 
buffer_wire buffer_11163 (.in(n11163), .out(n11163_0));
mux14 mux_5998 (.in({n14011_1, n13989_0, n13982_0/**/, n13975_0, n13968_0, n13954_0, n13939_0, n13924_1, n11078_1, n6933, n6925, n6917, n6829, n6821}), .out(n11164), .config_in(config_chain[20343:20338]), .config_rst(config_rst)); 
buffer_wire buffer_11164 (.in(n11164), .out(n11164_0));
mux3 mux_5999 (.in({n14739_0, n14738_0, n8789}), .out(n11165), .config_in(config_chain[20345:20344]), .config_rst(config_rst)); 
buffer_wire buffer_11165 (.in(n11165), .out(n11165_0));
mux13 mux_6000 (.in({n14013_1, n13997_0, n13990_0, n13976_0, n13961_0, n13947_0, n13940_0, n13922_1, n11080_1, n6925, n6917/**/, n6829, n6821}), .out(n11166), .config_in(config_chain[20351:20346]), .config_rst(config_rst)); 
buffer_wire buffer_11166 (.in(n11166), .out(n11166_0));
mux3 mux_6001 (.in({n14741_0, n14740_0/**/, n8873}), .out(n11167), .config_in(config_chain[20353:20352]), .config_rst(config_rst)); 
buffer_wire buffer_11167 (.in(n11167), .out(n11167_0));
mux13 mux_6002 (.in({n14015_1, n13998_0, n13983_0, n13969_0, n13962_0, n13955_0, n13948_0, n13920_1, n11082_1, n6929, n6917, n6829, n6821/**/}), .out(n11168), .config_in(config_chain[20359:20354]), .config_rst(config_rst)); 
buffer_wire buffer_11168 (.in(n11168), .out(n11168_0));
mux3 mux_6003 (.in({n14743_0, n14742_0/**/, n8877}), .out(n11169), .config_in(config_chain[20361:20360]), .config_rst(config_rst)); 
buffer_wire buffer_11169 (.in(n11169), .out(n11169_0));
mux13 mux_6004 (.in({n14017_1, n13991_0, n13984_0, n13977_0, n13970_0, n13956_0, n13941_0, n13918_1, n11084_1/**/, n6929, n6921, n6829, n6821}), .out(n11170), .config_in(config_chain[20367:20362]), .config_rst(config_rst)); 
buffer_wire buffer_11170 (.in(n11170), .out(n11170_0));
mux3 mux_6005 (.in({n14745_0, n14744_0, n8881}), .out(n11171), .config_in(config_chain[20369:20368]), .config_rst(config_rst)); 
buffer_wire buffer_11171 (.in(n11171), .out(n11171_0));
mux13 mux_6006 (.in({n14019_1, n13999_0, n13992_0, n13978_0, n13963_0, n13949_0, n13942_0, n13916_1, n11086_1, n6929, n6921, n6833, n6821/**/}), .out(n11172), .config_in(config_chain[20375:20370]), .config_rst(config_rst)); 
buffer_wire buffer_11172 (.in(n11172), .out(n11172_0));
mux3 mux_6007 (.in({n14747_0/**/, n14746_0, n8881}), .out(n11173), .config_in(config_chain[20377:20376]), .config_rst(config_rst)); 
buffer_wire buffer_11173 (.in(n11173), .out(n11173_0));
mux13 mux_6008 (.in({n14021_1, n14000_0, n13985_0, n13971_0, n13964_0, n13957_1, n13950_0, n13910_1, n11042_1, n6929, n6921, n6833, n6825}), .out(n11174), .config_in(config_chain[20383:20378]), .config_rst(config_rst)); 
buffer_wire buffer_11174 (.in(n11174), .out(n11174_0));
mux3 mux_6009 (.in({n14749_1, n14748_0, n8885}), .out(n11175), .config_in(config_chain[20385:20384]), .config_rst(config_rst)); 
buffer_wire buffer_11175 (.in(n11175), .out(n11175_0));
mux15 mux_6010 (.in({n14289_1, n14266_0, n14259_0, n14252_0, n14238_0, n14223_1, n14209_0, n14202_0, n14198_1, n11088_1, n7907, n7899, n7811, n7803, n7795}), .out(n11176), .config_in(config_chain[20391:20386]), .config_rst(config_rst)); 
buffer_wire buffer_11176 (.in(n11176), .out(n11176_0));
mux4 mux_6011 (.in({n14751_0, n14750_0, n8889, n8773}), .out(n11177), .config_in(config_chain[20393:20392]), .config_rst(config_rst)); 
buffer_wire buffer_11177 (.in(n11177), .out(n11177_0));
mux15 mux_6012 (.in({n14269_1, n14260_0, n14245_1, n14231_0/**/, n14224_0, n14217_0, n14210_0, n14196_1, n14178_1, n11090_1, n7911, n7899, n7811, n7803, n7795}), .out(n11178), .config_in(config_chain[20399:20394]), .config_rst(config_rst)); 
buffer_wire buffer_11178 (.in(n11178), .out(n11178_0));
mux3 mux_6013 (.in({n14753_0, n14752_0, n8773}), .out(n11179), .config_in(config_chain[20401:20400]), .config_rst(config_rst)); 
buffer_wire buffer_11179 (.in(n11179), .out(n11179_0));
mux15 mux_6014 (.in({n14271_1, n14267_1, n14253_0, n14246_0, n14239_0, n14232_0, n14218_0, n14203_0, n14194_1, n11092_1, n7911, n7903, n7811, n7803, n7795}), .out(n11180), .config_in(config_chain[20407:20402]), .config_rst(config_rst)); 
buffer_wire buffer_11180 (.in(n11180), .out(n11180_0));
mux3 mux_6015 (.in({n14755_0, n14754_0, n8777}), .out(n11181), .config_in(config_chain[20409:20408]), .config_rst(config_rst)); 
buffer_wire buffer_11181 (.in(n11181), .out(n11181_0));
mux15 mux_6016 (.in({n14273_1, n14261_0, n14254_0, n14240_0, n14225_0, n14211_0, n14204_0, n14192_1, n14179_0, n11094_1, n7911/**/, n7903, n7895, n7803, n7795}), .out(n11182), .config_in(config_chain[20415:20410]), .config_rst(config_rst)); 
buffer_wire buffer_11182 (.in(n11182), .out(n11182_0));
mux3 mux_6017 (.in({n14757_0, n14756_0, n8781}), .out(n11183), .config_in(config_chain[20417:20416]), .config_rst(config_rst)); 
buffer_wire buffer_11183 (.in(n11183), .out(n11183_0));
mux14 mux_6018 (.in({n14275_1, n14262_0, n14247_0, n14233_0, n14226_0, n14219_0, n14212_0, n14190_1, n11096_1, n7911, n7903, n7895, n7807, n7795}), .out(n11184), .config_in(config_chain[20423:20418]), .config_rst(config_rst)); 
buffer_wire buffer_11184 (.in(n11184), .out(n11184_0));
mux3 mux_6019 (.in({n14759_0, n14758_0, n8785}), .out(n11185), .config_in(config_chain[20425:20424]), .config_rst(config_rst)); 
buffer_wire buffer_11185 (.in(n11185), .out(n11185_0));
mux14 mux_6020 (.in({n14277_1, n14255_0/**/, n14248_0, n14241_0, n14234_0, n14220_0, n14205_0, n14188_1, n11098_1, n7911, n7903, n7895, n7807, n7799}), .out(n11186), .config_in(config_chain[20431:20426]), .config_rst(config_rst)); 
buffer_wire buffer_11186 (.in(n11186), .out(n11186_0));
mux3 mux_6021 (.in({n14761_0, n14760_0, n8789}), .out(n11187), .config_in(config_chain[20433:20432]), .config_rst(config_rst)); 
buffer_wire buffer_11187 (.in(n11187), .out(n11187_0));
mux13 mux_6022 (.in({n14279_1, n14263_0, n14256_0, n14242_0, n14227_0, n14213_0/**/, n14206_0, n14186_1, n11100_1, n7903, n7895, n7807, n7799}), .out(n11188), .config_in(config_chain[20439:20434]), .config_rst(config_rst)); 
buffer_wire buffer_11188 (.in(n11188), .out(n11188_0));
mux3 mux_6023 (.in({n14763_0/**/, n14762_0, n8789}), .out(n11189), .config_in(config_chain[20441:20440]), .config_rst(config_rst)); 
buffer_wire buffer_11189 (.in(n11189), .out(n11189_0));
mux13 mux_6024 (.in({n14281_1, n14264_0, n14249_0, n14235_0, n14228_0, n14221_0, n14214_0, n14184_1, n11102_1, n7907, n7895, n7807/**/, n7799}), .out(n11190), .config_in(config_chain[20447:20442]), .config_rst(config_rst)); 
buffer_wire buffer_11190 (.in(n11190), .out(n11190_0));
mux3 mux_6025 (.in({n14765_0, n14764_0, n8873}), .out(n11191), .config_in(config_chain[20449:20448]), .config_rst(config_rst)); 
buffer_wire buffer_11191 (.in(n11191), .out(n11191_0));
mux13 mux_6026 (.in({n14283_1, n14257_0, n14250_0, n14243_0, n14236_0, n14207_0, n14200_1, n14182_1, n11104_1, n7907, n7899, n7807, n7799/**/}), .out(n11192), .config_in(config_chain[20455:20450]), .config_rst(config_rst)); 
buffer_wire buffer_11192 (.in(n11192), .out(n11192_0));
mux3 mux_6027 (.in({n14767_0, n14766_0, n8877}), .out(n11193), .config_in(config_chain[20457:20456]), .config_rst(config_rst)); 
buffer_wire buffer_11193 (.in(n11193), .out(n11193_0));
mux13 mux_6028 (.in({n14285_1, n14265_0, n14258_0, n14229_0, n14222_0, n14215_0, n14208_0, n14180_1, n11106_1/**/, n7907, n7899, n7811, n7799}), .out(n11194), .config_in(config_chain[20463:20458]), .config_rst(config_rst)); 
buffer_wire buffer_11194 (.in(n11194), .out(n11194_0));
mux3 mux_6029 (.in({n14769_0/**/, n14768_0, n8881}), .out(n11195), .config_in(config_chain[20465:20464]), .config_rst(config_rst)); 
buffer_wire buffer_11195 (.in(n11195), .out(n11195_0));
mux13 mux_6030 (.in({n14287_1, n14251_0, n14244_0, n14237_0, n14230_0, n14216_0, n14201_1, n14176_1, n11044_2, n7907, n7899, n7811, n7803}), .out(n11196), .config_in(config_chain[20471:20466]), .config_rst(config_rst)); 
buffer_wire buffer_11196 (.in(n11196), .out(n11196_0));
mux3 mux_6031 (.in({n14771_1, n14770_0, n8885}), .out(n11197), .config_in(config_chain[20473:20472]), .config_rst(config_rst)); 
buffer_wire buffer_11197 (.in(n11197), .out(n11197_0));
mux15 mux_6032 (.in({n14553_1, n14517_0, n14510_0, n14508_0, n14501_0, n14494_0, n14480_0, n14465_1, n14462_1, n11110_1, n8885, n8877, n8789, n8781, n8773}), .out(n11198), .config_in(config_chain[20479:20474]), .config_rst(config_rst)); 
buffer_wire buffer_11198 (.in(n11198), .out(n11198_0));
mux4 mux_6033 (.in({n14773_0, n14772_0/**/, n8889, n8773}), .out(n11199), .config_in(config_chain[20481:20480]), .config_rst(config_rst)); 
buffer_wire buffer_11199 (.in(n11199), .out(n11199_0));
mux15 mux_6034 (.in({n14533_1, n14530_0, n14525_0, n14518_0, n14502_0, n14487_1, n14473_0, n14466_0, n14460_1/**/, n11112_1, n8889, n8877, n8789, n8781, n8773}), .out(n11200), .config_in(config_chain[20487:20482]), .config_rst(config_rst)); 
buffer_wire buffer_11200 (.in(n11200), .out(n11200_0));
mux3 mux_6035 (.in({n14775_0, n14774_0, n8777}), .out(n11201), .config_in(config_chain[20489:20488]), .config_rst(config_rst)); 
buffer_wire buffer_11201 (.in(n11201), .out(n11201_0));
mux15 mux_6036 (.in({n14535_1, n14526_0, n14511_0, n14509_1, n14495_0, n14488_0, n14481_0, n14474_0, n14458_1/**/, n11114_1, n8889, n8881, n8789, n8781, n8773}), .out(n11202), .config_in(config_chain[20495:20490]), .config_rst(config_rst)); 
buffer_wire buffer_11202 (.in(n11202), .out(n11202_0));
mux3 mux_6037 (.in({n14777_0, n14776_0, n8777}), .out(n11203), .config_in(config_chain[20497:20496]), .config_rst(config_rst)); 
buffer_wire buffer_11203 (.in(n11203), .out(n11203_0));
mux15 mux_6038 (.in({n14537_1, n14531_1, n14519_0, n14512_0, n14503_0/**/, n14496_0, n14482_0, n14467_0, n14456_1, n11116_1, n8889, n8881, n8873, n8781, n8773}), .out(n11204), .config_in(config_chain[20503:20498]), .config_rst(config_rst)); 
buffer_wire buffer_11204 (.in(n11204), .out(n11204_0));
mux3 mux_6039 (.in({n14779_0, n14778_0, n8781}), .out(n11205), .config_in(config_chain[20505:20504]), .config_rst(config_rst)); 
buffer_wire buffer_11205 (.in(n11205), .out(n11205_0));
mux14 mux_6040 (.in({n14539_1, n14527_0, n14520_0/**/, n14504_0, n14489_0, n14475_0, n14468_0, n14454_1, n11118_1, n8889, n8881, n8873, n8785, n8773}), .out(n11206), .config_in(config_chain[20511:20506]), .config_rst(config_rst)); 
buffer_wire buffer_11206 (.in(n11206), .out(n11206_0));
mux3 mux_6041 (.in({n14781_0/**/, n14780_0, n8785}), .out(n11207), .config_in(config_chain[20513:20512]), .config_rst(config_rst)); 
buffer_wire buffer_11207 (.in(n11207), .out(n11207_0));
mux14 mux_6042 (.in({n14541_1, n14528_0, n14513_0, n14497_0, n14490_0, n14483_0, n14476_0, n14452_1, n11120_1, n8889, n8881, n8873, n8785, n8777}), .out(n11208), .config_in(config_chain[20519:20514]), .config_rst(config_rst)); 
buffer_wire buffer_11208 (.in(n11208), .out(n11208_0));
mux3 mux_6043 (.in({n14783_0, n14782_0, n8789}), .out(n11209), .config_in(config_chain[20521:20520]), .config_rst(config_rst)); 
buffer_wire buffer_11209 (.in(n11209), .out(n11209_0));
mux13 mux_6044 (.in({n14543_1, n14521_0, n14514_0, n14505_0, n14498_0, n14484_0, n14469_0, n14450_1/**/, n11122_1, n8881, n8873, n8785, n8777}), .out(n11210), .config_in(config_chain[20527:20522]), .config_rst(config_rst)); 
buffer_wire buffer_11210 (.in(n11210), .out(n11210_0));
mux3 mux_6045 (.in({n14785_0, n14784_0, n8873}), .out(n11211), .config_in(config_chain[20529:20528]), .config_rst(config_rst)); 
buffer_wire buffer_11211 (.in(n11211), .out(n11211_0));
mux13 mux_6046 (.in({n14545_1, n14529_0, n14522_0, n14506_0, n14491_0, n14477_0, n14470_0/**/, n14448_1, n11124_1, n8885, n8873, n8785, n8777}), .out(n11212), .config_in(config_chain[20535:20530]), .config_rst(config_rst)); 
buffer_wire buffer_11212 (.in(n11212), .out(n11212_0));
mux3 mux_6047 (.in({n14787_0, n14786_0, n8873}), .out(n11213), .config_in(config_chain[20537:20536]), .config_rst(config_rst)); 
buffer_wire buffer_11213 (.in(n11213), .out(n11213_0));
mux13 mux_6048 (.in({n14547_1, n14515_0, n14499_0, n14492_0, n14485_0, n14478_0, n14446_1, n14432_1, n11126_1, n8885, n8877, n8785, n8777}), .out(n11214), .config_in(config_chain[20543:20538]), .config_rst(config_rst)); 
buffer_wire buffer_11214 (.in(n11214), .out(n11214_0));
mux3 mux_6049 (.in({n14789_0, n14788_0, n8877/**/}), .out(n11215), .config_in(config_chain[20545:20544]), .config_rst(config_rst)); 
buffer_wire buffer_11215 (.in(n11215), .out(n11215_0));
mux13 mux_6050 (.in({n14549_1, n14523_0, n14516_0/**/, n14507_0, n14500_0, n14471_0, n14464_1, n14444_1, n11128_1, n8885, n8877, n8789, n8777}), .out(n11216), .config_in(config_chain[20551:20546]), .config_rst(config_rst)); 
buffer_wire buffer_11216 (.in(n11216), .out(n11216_0));
mux3 mux_6051 (.in({n14791_0, n14790_0, n8881}), .out(n11217), .config_in(config_chain[20553:20552]), .config_rst(config_rst)); 
buffer_wire buffer_11217 (.in(n11217), .out(n11217_0));
mux13 mux_6052 (.in({n14551_1, n14524_0, n14493_0, n14486_0, n14479_0, n14472_0, n14442_1, n14433_1, n11046_2, n8885, n8877, n8789, n8781}), .out(n11218), .config_in(config_chain[20559:20554]), .config_rst(config_rst)); 
buffer_wire buffer_11218 (.in(n11218), .out(n11218_0));
mux3 mux_6053 (.in({n14793_1, n14792_0/**/, n8889}), .out(n11219), .config_in(config_chain[20561:20560]), .config_rst(config_rst)); 
buffer_wire buffer_11219 (.in(n11219), .out(n11219_0));
mux4 mux_6054 (.in({n12423_0, n12422_0, n1163, n1047}), .out(n11220), .config_in(config_chain[20563:20562]), .config_rst(config_rst)); 
buffer_wire buffer_11220 (.in(n11220), .out(n11220_0));
mux15 mux_6055 (.in({n12973_0, n12964_0, n12959_0, n12947_0, n12918_0, n12913_0, n12869_0, n12864_1, n12860_1, n11333_1, n2137, n2129/**/, n2041, n2033, n2025}), .out(n11221), .config_in(config_chain[20569:20564]), .config_rst(config_rst)); 
buffer_wire buffer_11221 (.in(n11221), .out(n11221_0));
mux4 mux_6056 (.in({n12443_0, n12442_0, n1163, n1047}), .out(n11222), .config_in(config_chain[20571:20570]), .config_rst(config_rst)); 
buffer_wire buffer_11222 (.in(n11222), .out(n11222_0));
mux15 mux_6057 (.in({n13233_0, n13216_0, n13211_0, n13202_0, n13197_0, n13185_0, n13127_0, n13122_1, n13120_1, n11355_1, n3115, n3107, n3019/**/, n3011, n3003}), .out(n11223), .config_in(config_chain[20577:20572]), .config_rst(config_rst)); 
buffer_wire buffer_11223 (.in(n11223), .out(n11223_0));
mux4 mux_6058 (.in({n12463_0, n12382_1/**/, n1163, n1047}), .out(n11224), .config_in(config_chain[20579:20578]), .config_rst(config_rst)); 
buffer_wire buffer_11224 (.in(n11224), .out(n11224_0));
mux15 mux_6059 (.in({n13495_0, n13492_0, n13487_0, n13456_0, n13451_0, n13442_0, n13437_0, n13387_0, n13382_1, n11377_1, n4093, n4085/**/, n3997, n3989, n3981}), .out(n11225), .config_in(config_chain[20585:20580]), .config_rst(config_rst)); 
buffer_wire buffer_11225 (.in(n11225), .out(n11225_0));
mux4 mux_6060 (.in({n12403_0, n12402_0, n1163, n1047}), .out(n11226), .config_in(config_chain[20587:20586]), .config_rst(config_rst)); 
buffer_wire buffer_11226 (.in(n11226), .out(n11226_0));
mux16 mux_6061 (.in({n12717_0, n12709_0, n12704_0, n12683_0, n12678_0, n12672_0, n12657_0, n12654_1, n12612_1, n12605_0, n11313_1, n1159, n1151, n1063, n1055, n1047}), .out(n11227), .config_in(config_chain[20593:20588]), .config_rst(config_rst)); 
buffer_wire buffer_11227 (.in(n11227), .out(n11227_0));
mux3 mux_6062 (.in({n12425_0, n12424_0, n1047}), .out(n11228), .config_in(config_chain[20595:20594]), .config_rst(config_rst)); 
buffer_wire buffer_11228 (.in(n11228), .out(n11228_0));
mux15 mux_6063 (.in({n12993_0, n12967_0, n12938_0, n12933_0, n12926_0, n12921_0, n12892_1/**/, n12871_0, n12866_1, n11335_1, n2141, n2129, n2041, n2033, n2025}), .out(n11229), .config_in(config_chain[20601:20596]), .config_rst(config_rst)); 
buffer_wire buffer_11229 (.in(n11229), .out(n11229_0));
mux3 mux_6064 (.in({n12445_0, n12444_0, n1051}), .out(n11230), .config_in(config_chain[20603:20602]), .config_rst(config_rst)); 
buffer_wire buffer_11230 (.in(n11230), .out(n11230_0));
mux15 mux_6065 (.in({n13253_0, n13224_0, n13219_0, n13205_0, n13176_0, n13171_0, n13150_1/**/, n13129_0, n13124_1, n11357_1, n3119, n3107, n3019, n3011, n3003}), .out(n11231), .config_in(config_chain[20609:20604]), .config_rst(config_rst)); 
buffer_wire buffer_11231 (.in(n11231), .out(n11231_0));
mux3 mux_6066 (.in({n12465_0, n12384_1/**/, n1051}), .out(n11232), .config_in(config_chain[20611:20610]), .config_rst(config_rst)); 
buffer_wire buffer_11232 (.in(n11232), .out(n11232_0));
mux15 mux_6067 (.in({n13515_0, n13478_0, n13473_0, n13464_0, n13459_0, n13445_0, n13410_1, n13389_0, n13384_1, n11379_1, n4097, n4085, n3997, n3989, n3981}), .out(n11233), .config_in(config_chain[20617:20612]), .config_rst(config_rst)); 
buffer_wire buffer_11233 (.in(n11233), .out(n11233_0));
mux3 mux_6068 (.in({n12405_0, n12404_0/**/, n1051}), .out(n11234), .config_in(config_chain[20619:20618]), .config_rst(config_rst)); 
buffer_wire buffer_11234 (.in(n11234), .out(n11234_0));
mux16 mux_6069 (.in({n12735_0, n12703_0, n12698_0/**/, n12692_0, n12677_0, n12671_0, n12666_0, n12636_1, n12614_1, n12607_0, n11315_1, n1159, n1151, n1063, n1055, n1047}), .out(n11235), .config_in(config_chain[20625:20620]), .config_rst(config_rst)); 
buffer_wire buffer_11235 (.in(n11235), .out(n11235_0));
mux3 mux_6070 (.in({n12427_0, n12426_0, n1051/**/}), .out(n11236), .config_in(config_chain[20627:20626]), .config_rst(config_rst)); 
buffer_wire buffer_11236 (.in(n11236), .out(n11236_0));
mux15 mux_6071 (.in({n12991_0, n12958_0, n12953_0, n12946_0/**/, n12941_0, n12929_0, n12912_0, n12894_1, n12868_1, n11337_1, n2141, n2133, n2041, n2033, n2025}), .out(n11237), .config_in(config_chain[20633:20628]), .config_rst(config_rst)); 
buffer_wire buffer_11237 (.in(n11237), .out(n11237_0));
mux3 mux_6072 (.in({n12447_0, n12446_0/**/, n1051}), .out(n11238), .config_in(config_chain[20635:20634]), .config_rst(config_rst)); 
buffer_wire buffer_11238 (.in(n11238), .out(n11238_0));
mux15 mux_6073 (.in({n13251_0, n13227_0, n13210_0, n13196_0, n13191_0/**/, n13184_0, n13179_0, n13152_1, n13126_1, n11359_1, n3119, n3111, n3019, n3011, n3003}), .out(n11239), .config_in(config_chain[20641:20636]), .config_rst(config_rst)); 
buffer_wire buffer_11239 (.in(n11239), .out(n11239_0));
mux3 mux_6074 (.in({n12467_0, n12386_1, n1055}), .out(n11240), .config_in(config_chain[20643:20642]), .config_rst(config_rst)); 
buffer_wire buffer_11240 (.in(n11240), .out(n11240_0));
mux15 mux_6075 (.in({n13513_0, n13486_0, n13481_0, n13467_0, n13450_0, n13436_0, n13431_0, n13412_1, n13386_1, n11381_1/**/, n4097, n4089, n3997, n3989, n3981}), .out(n11241), .config_in(config_chain[20649:20644]), .config_rst(config_rst)); 
buffer_wire buffer_11241 (.in(n11241), .out(n11241_0));
mux3 mux_6076 (.in({n12407_0, n12406_0, n1055}), .out(n11242), .config_in(config_chain[20651:20650]), .config_rst(config_rst)); 
buffer_wire buffer_11242 (.in(n11242), .out(n11242_0));
mux15 mux_6077 (.in({n12733_0, n12712_0, n12697_0, n12691_0, n12686_0, n12665_0, n12660_0/**/, n12638_1, n12609_0, n11317_1, n1159, n1151, n1063, n1055, n1047}), .out(n11243), .config_in(config_chain[20657:20652]), .config_rst(config_rst)); 
buffer_wire buffer_11243 (.in(n11243), .out(n11243_0));
mux3 mux_6078 (.in({n12429_0, n12428_0/**/, n1055}), .out(n11244), .config_in(config_chain[20659:20658]), .config_rst(config_rst)); 
buffer_wire buffer_11244 (.in(n11244), .out(n11244_0));
mux15 mux_6079 (.in({n12989_0, n12966_0, n12961_0, n12949_0, n12932_0, n12920_0, n12915_0, n12896_1, n12870_1, n11339_1, n2141, n2133, n2125, n2033, n2025}), .out(n11245), .config_in(config_chain[20665:20660]), .config_rst(config_rst)); 
buffer_wire buffer_11245 (.in(n11245), .out(n11245_0));
mux3 mux_6080 (.in({n12449_0, n12448_0/**/, n1055}), .out(n11246), .config_in(config_chain[20667:20666]), .config_rst(config_rst)); 
buffer_wire buffer_11246 (.in(n11246), .out(n11246_0));
mux15 mux_6081 (.in({n13249_0, n13218_0/**/, n13213_0, n13204_0, n13199_0, n13187_0, n13170_0, n13154_1, n13128_1, n11361_1, n3119, n3111, n3103, n3011, n3003}), .out(n11247), .config_in(config_chain[20673:20668]), .config_rst(config_rst)); 
buffer_wire buffer_11247 (.in(n11247), .out(n11247_0));
mux3 mux_6082 (.in({n12469_0, n12388_1/**/, n1055}), .out(n11248), .config_in(config_chain[20675:20674]), .config_rst(config_rst)); 
buffer_wire buffer_11248 (.in(n11248), .out(n11248_0));
mux15 mux_6083 (.in({n13511_0, n13489_0, n13472_0, n13458_0, n13453_0, n13444_0, n13439_0, n13414_1, n13388_1, n11383_1, n4097, n4089, n4081/**/, n3989, n3981}), .out(n11249), .config_in(config_chain[20681:20676]), .config_rst(config_rst)); 
buffer_wire buffer_11249 (.in(n11249), .out(n11249_0));
mux3 mux_6084 (.in({n12409_0/**/, n12408_0, n1059}), .out(n11250), .config_in(config_chain[20683:20682]), .config_rst(config_rst)); 
buffer_wire buffer_11250 (.in(n11250), .out(n11250_0));
mux15 mux_6085 (.in({n12731_0/**/, n12711_0, n12706_0, n12685_0, n12680_0, n12674_0, n12659_0, n12640_1, n12611_0, n11319_1, n1159, n1151, n1063, n1055, n1047}), .out(n11251), .config_in(config_chain[20689:20684]), .config_rst(config_rst)); 
buffer_wire buffer_11251 (.in(n11251), .out(n11251_0));
mux3 mux_6086 (.in({n12431_0, n12430_0/**/, n1059}), .out(n11252), .config_in(config_chain[20691:20690]), .config_rst(config_rst)); 
buffer_wire buffer_11252 (.in(n11252), .out(n11252_0));
mux14 mux_6087 (.in({n12987_0, n12969_0, n12952_0, n12940_0, n12935_0, n12928_0/**/, n12923_0, n12898_1, n11341_1, n2141, n2133, n2125, n2037, n2025}), .out(n11253), .config_in(config_chain[20697:20692]), .config_rst(config_rst)); 
buffer_wire buffer_11253 (.in(n11253), .out(n11253_0));
mux3 mux_6088 (.in({n12451_0, n12450_0, n1059}), .out(n11254), .config_in(config_chain[20699:20698]), .config_rst(config_rst)); 
buffer_wire buffer_11254 (.in(n11254), .out(n11254_0));
mux14 mux_6089 (.in({n13247_0, n13226_0, n13221_0, n13207_0, n13190_0, n13178_0, n13173_0, n13156_1, n11363_1, n3119, n3111, n3103, n3015, n3003}), .out(n11255), .config_in(config_chain[20705:20700]), .config_rst(config_rst)); 
buffer_wire buffer_11255 (.in(n11255), .out(n11255_0));
mux3 mux_6090 (.in({n12471_0, n12390_1/**/, n1059}), .out(n11256), .config_in(config_chain[20707:20706]), .config_rst(config_rst)); 
buffer_wire buffer_11256 (.in(n11256), .out(n11256_0));
mux14 mux_6091 (.in({n13509_0, n13480_0, n13475_0, n13466_0/**/, n13461_0, n13447_0, n13430_0, n13416_1, n11385_1, n4097, n4089, n4081, n3993, n3981}), .out(n11257), .config_in(config_chain[20713:20708]), .config_rst(config_rst)); 
buffer_wire buffer_11257 (.in(n11257), .out(n11257_0));
mux3 mux_6092 (.in({n12411_0, n12410_0, n1059}), .out(n11258), .config_in(config_chain[20715:20714]), .config_rst(config_rst)); 
buffer_wire buffer_11258 (.in(n11258), .out(n11258_0));
mux15 mux_6093 (.in({n12729_0, n12705_0, n12700_0, n12694_0/**/, n12679_0, n12673_0, n12668_0, n12642_1, n12613_0, n11321_1, n1159, n1151, n1063, n1055, n1047}), .out(n11259), .config_in(config_chain[20721:20716]), .config_rst(config_rst)); 
buffer_wire buffer_11259 (.in(n11259), .out(n11259_0));
mux3 mux_6094 (.in({n12433_0, n12432_0/**/, n1063}), .out(n11260), .config_in(config_chain[20723:20722]), .config_rst(config_rst)); 
buffer_wire buffer_11260 (.in(n11260), .out(n11260_0));
mux14 mux_6095 (.in({n12985_0, n12960_0, n12955_0, n12948_0, n12943_0, n12931_0, n12914_0, n12900_1, n11343_1, n2141, n2133, n2125, n2037, n2029}), .out(n11261), .config_in(config_chain[20729:20724]), .config_rst(config_rst)); 
buffer_wire buffer_11261 (.in(n11261), .out(n11261_0));
mux3 mux_6096 (.in({n12453_0, n12452_0, n1063}), .out(n11262), .config_in(config_chain[20731:20730]), .config_rst(config_rst)); 
buffer_wire buffer_11262 (.in(n11262), .out(n11262_0));
mux14 mux_6097 (.in({n13245_0, n13229_0, n13212_0, n13198_0, n13193_0, n13186_0, n13181_0, n13158_1, n11365_1, n3119, n3111, n3103, n3015/**/, n3007}), .out(n11263), .config_in(config_chain[20737:20732]), .config_rst(config_rst)); 
buffer_wire buffer_11263 (.in(n11263), .out(n11263_0));
mux3 mux_6098 (.in({n12473_0, n12392_1, n1063/**/}), .out(n11264), .config_in(config_chain[20739:20738]), .config_rst(config_rst)); 
buffer_wire buffer_11264 (.in(n11264), .out(n11264_0));
mux14 mux_6099 (.in({n13507_0, n13488_0, n13483_0, n13469_0, n13452_0, n13438_0, n13433_0, n13418_1/**/, n11387_1, n4097, n4089, n4081, n3993, n3985}), .out(n11265), .config_in(config_chain[20745:20740]), .config_rst(config_rst)); 
buffer_wire buffer_11265 (.in(n11265), .out(n11265_0));
mux3 mux_6100 (.in({n12413_0, n12412_0, n1063}), .out(n11266), .config_in(config_chain[20747:20746]), .config_rst(config_rst)); 
buffer_wire buffer_11266 (.in(n11266), .out(n11266_0));
mux15 mux_6101 (.in({n12727_0, n12714_0, n12699_0, n12693_0, n12688_0/**/, n12667_0, n12662_0, n12644_1, n12615_0, n11323_1, n1163, n1155, n1147, n1059, n1051}), .out(n11267), .config_in(config_chain[20753:20748]), .config_rst(config_rst)); 
buffer_wire buffer_11267 (.in(n11267), .out(n11267_0));
mux3 mux_6102 (.in({n12435_0, n12434_0/**/, n1063}), .out(n11268), .config_in(config_chain[20755:20754]), .config_rst(config_rst)); 
buffer_wire buffer_11268 (.in(n11268), .out(n11268_0));
mux13 mux_6103 (.in({n12983_0, n12968_0, n12963_0, n12951_0, n12934_0, n12922_0/**/, n12917_0, n12902_1, n11345_1, n2133, n2125, n2037, n2029}), .out(n11269), .config_in(config_chain[20761:20756]), .config_rst(config_rst)); 
buffer_wire buffer_11269 (.in(n11269), .out(n11269_0));
mux3 mux_6104 (.in({n12455_0, n12454_0, n1147}), .out(n11270), .config_in(config_chain[20763:20762]), .config_rst(config_rst)); 
buffer_wire buffer_11270 (.in(n11270), .out(n11270_0));
mux13 mux_6105 (.in({n13243_0, n13220_0, n13215_0, n13206_0, n13201_0, n13189_0, n13172_0, n13160_1, n11367_1/**/, n3111, n3103, n3015, n3007}), .out(n11271), .config_in(config_chain[20769:20764]), .config_rst(config_rst)); 
buffer_wire buffer_11271 (.in(n11271), .out(n11271_0));
mux3 mux_6106 (.in({n12475_0, n12394_1, n1147}), .out(n11272), .config_in(config_chain[20771:20770]), .config_rst(config_rst)); 
buffer_wire buffer_11272 (.in(n11272), .out(n11272_0));
mux13 mux_6107 (.in({n13505_0, n13491_0, n13474_0, n13460_0, n13455_0, n13446_0, n13441_0, n13420_1, n11389_1, n4089, n4081, n3993, n3985/**/}), .out(n11273), .config_in(config_chain[20777:20772]), .config_rst(config_rst)); 
buffer_wire buffer_11273 (.in(n11273), .out(n11273_0));
mux3 mux_6108 (.in({n12415_0, n12414_0, n1147}), .out(n11274), .config_in(config_chain[20779:20778]), .config_rst(config_rst)); 
buffer_wire buffer_11274 (.in(n11274), .out(n11274_0));
mux15 mux_6109 (.in({n12725_0, n12713_0, n12708_0, n12687_0, n12682_0, n12661_0, n12656_0, n12646_1, n12604_1, n11325_1, n1163/**/, n1155, n1147, n1059, n1051}), .out(n11275), .config_in(config_chain[20785:20780]), .config_rst(config_rst)); 
buffer_wire buffer_11275 (.in(n11275), .out(n11275_0));
mux3 mux_6110 (.in({n12437_0, n12436_0, n1147}), .out(n11276), .config_in(config_chain[20787:20786]), .config_rst(config_rst)); 
buffer_wire buffer_11276 (.in(n11276), .out(n11276_0));
mux13 mux_6111 (.in({n12981_0/**/, n12971_0, n12954_0, n12942_0, n12937_0, n12930_0, n12925_0, n12904_1, n11347_1, n2137, n2125, n2037, n2029}), .out(n11277), .config_in(config_chain[20793:20788]), .config_rst(config_rst)); 
buffer_wire buffer_11277 (.in(n11277), .out(n11277_0));
mux3 mux_6112 (.in({n12457_0, n12456_0, n1147}), .out(n11278), .config_in(config_chain[20795:20794]), .config_rst(config_rst)); 
buffer_wire buffer_11278 (.in(n11278), .out(n11278_0));
mux13 mux_6113 (.in({n13241_0, n13228_0, n13223_0, n13209_0, n13192_0, n13180_0, n13175_0, n13162_1, n11369_1, n3115/**/, n3103, n3015, n3007}), .out(n11279), .config_in(config_chain[20801:20796]), .config_rst(config_rst)); 
buffer_wire buffer_11279 (.in(n11279), .out(n11279_0));
mux3 mux_6114 (.in({n12477_0, n12396_1, n1151}), .out(n11280), .config_in(config_chain[20803:20802]), .config_rst(config_rst)); 
buffer_wire buffer_11280 (.in(n11280), .out(n11280_0));
mux13 mux_6115 (.in({n13503_0, n13482_0, n13477_0, n13468_0, n13463_0, n13449_0, n13432_0, n13422_1, n11391_1, n4093, n4081, n3993, n3985/**/}), .out(n11281), .config_in(config_chain[20809:20804]), .config_rst(config_rst)); 
buffer_wire buffer_11281 (.in(n11281), .out(n11281_0));
mux3 mux_6116 (.in({n12417_0, n12416_0, n1151}), .out(n11282), .config_in(config_chain[20811:20810]), .config_rst(config_rst)); 
buffer_wire buffer_11282 (.in(n11282), .out(n11282_0));
mux15 mux_6117 (.in({n12723_0, n12707_0, n12702_0, n12681_0, n12676_0/**/, n12675_0, n12670_0, n12648_1, n12606_1, n11327_1, n1163, n1155, n1147, n1059, n1051}), .out(n11283), .config_in(config_chain[20817:20812]), .config_rst(config_rst)); 
buffer_wire buffer_11283 (.in(n11283), .out(n11283_0));
mux3 mux_6118 (.in({n12439_0, n12438_0/**/, n1151}), .out(n11284), .config_in(config_chain[20819:20818]), .config_rst(config_rst)); 
buffer_wire buffer_11284 (.in(n11284), .out(n11284_0));
mux13 mux_6119 (.in({n12979_0, n12962_0/**/, n12957_0, n12950_0, n12945_0, n12916_0, n12906_1, n12863_0, n11349_1, n2137, n2129, n2037, n2029}), .out(n11285), .config_in(config_chain[20825:20820]), .config_rst(config_rst)); 
buffer_wire buffer_11285 (.in(n11285), .out(n11285_0));
mux3 mux_6120 (.in({n12459_0, n12458_0/**/, n1151}), .out(n11286), .config_in(config_chain[20827:20826]), .config_rst(config_rst)); 
buffer_wire buffer_11286 (.in(n11286), .out(n11286_0));
mux13 mux_6121 (.in({n13239_0, n13231_0, n13214_0, n13200_0, n13195_0, n13188_0, n13183_0, n13164_1, n11371_1, n3115/**/, n3107, n3015, n3007}), .out(n11287), .config_in(config_chain[20833:20828]), .config_rst(config_rst)); 
buffer_wire buffer_11287 (.in(n11287), .out(n11287_0));
mux3 mux_6122 (.in({n12479_0/**/, n12398_1, n1151}), .out(n11288), .config_in(config_chain[20835:20834]), .config_rst(config_rst)); 
buffer_wire buffer_11288 (.in(n11288), .out(n11288_0));
mux13 mux_6123 (.in({n13501_0, n13490_0, n13485_0, n13471_0, n13454_0, n13440_0, n13435_0, n13424_1, n11393_1, n4093, n4085, n3993, n3985}), .out(n11289), .config_in(config_chain[20841:20836]), .config_rst(config_rst)); 
buffer_wire buffer_11289 (.in(n11289), .out(n11289_0));
mux3 mux_6124 (.in({n12419_0, n12418_0, n1155}), .out(n11290), .config_in(config_chain[20843:20842]), .config_rst(config_rst)); 
buffer_wire buffer_11290 (.in(n11290), .out(n11290_0));
mux15 mux_6125 (.in({n12721_0, n12701_0, n12696_0, n12695_0, n12690_0/**/, n12669_0, n12664_0, n12650_1, n12608_1, n11329_1, n1163, n1155, n1147, n1059, n1051}), .out(n11291), .config_in(config_chain[20849:20844]), .config_rst(config_rst)); 
buffer_wire buffer_11291 (.in(n11291), .out(n11291_0));
mux3 mux_6126 (.in({n12441_0, n12440_0/**/, n1155}), .out(n11292), .config_in(config_chain[20851:20850]), .config_rst(config_rst)); 
buffer_wire buffer_11292 (.in(n11292), .out(n11292_0));
mux13 mux_6127 (.in({n12977_0, n12970_0, n12965_0, n12936_0, n12924_0, n12919_0, n12908_1, n12865_0, n11351_1/**/, n2137, n2129, n2041, n2029}), .out(n11293), .config_in(config_chain[20857:20852]), .config_rst(config_rst)); 
buffer_wire buffer_11293 (.in(n11293), .out(n11293_0));
mux3 mux_6128 (.in({n12461_0, n12460_0, n1155}), .out(n11294), .config_in(config_chain[20859:20858]), .config_rst(config_rst)); 
buffer_wire buffer_11294 (.in(n11294), .out(n11294_0));
mux13 mux_6129 (.in({n13237_0, n13222_0, n13217_0/**/, n13208_0, n13203_0, n13174_0, n13166_1, n13123_0, n11373_1, n3115, n3107, n3019, n3007}), .out(n11295), .config_in(config_chain[20865:20860]), .config_rst(config_rst)); 
buffer_wire buffer_11295 (.in(n11295), .out(n11295_0));
mux3 mux_6130 (.in({n12481_0, n12400_1, n1155}), .out(n11296), .config_in(config_chain[20867:20866]), .config_rst(config_rst)); 
buffer_wire buffer_11296 (.in(n11296), .out(n11296_0));
mux13 mux_6131 (.in({n13499_0, n13493_0, n13476_0, n13462_0, n13457_0, n13448_0, n13443_0/**/, n13426_1, n11395_1, n4093, n4085, n3997, n3985}), .out(n11297), .config_in(config_chain[20873:20868]), .config_rst(config_rst)); 
buffer_wire buffer_11297 (.in(n11297), .out(n11297_0));
mux3 mux_6132 (.in({n12421_0, n12420_0, n1155}), .out(n11298), .config_in(config_chain[20875:20874]), .config_rst(config_rst)); 
buffer_wire buffer_11298 (.in(n11298), .out(n11298_0));
mux15 mux_6133 (.in({n12719_0, n12715_0, n12710_0, n12689_0, n12684_0, n12663_0, n12658_0, n12652_1, n12610_1, n11331_1, n1163, n1155, n1147, n1059, n1051}), .out(n11299), .config_in(config_chain[20881:20876]), .config_rst(config_rst)); 
buffer_wire buffer_11299 (.in(n11299), .out(n11299_0));
mux3 mux_6134 (.in({n12351_0, n12350_1, n1159}), .out(n11300), .config_in(config_chain[20883:20882]), .config_rst(config_rst)); 
buffer_wire buffer_11300 (.in(n11300), .out(n11300_0));
mux13 mux_6135 (.in({n12975_0, n12956_0, n12944_0, n12939_0, n12927_0, n12910_1, n12867_0, n12862_1, n11353_2, n2137, n2129, n2041/**/, n2033}), .out(n11301), .config_in(config_chain[20889:20884]), .config_rst(config_rst)); 
buffer_wire buffer_11301 (.in(n11301), .out(n11301_0));
mux3 mux_6136 (.in({n12353_0, n12352_1, n1159}), .out(n11302), .config_in(config_chain[20891:20890]), .config_rst(config_rst)); 
buffer_wire buffer_11302 (.in(n11302), .out(n11302_0));
mux13 mux_6137 (.in({n13235_0, n13230_0, n13225_0, n13194_0, n13182_0/**/, n13177_0, n13168_1, n13125_0, n11375_1, n3115, n3107, n3019, n3011}), .out(n11303), .config_in(config_chain[20897:20892]), .config_rst(config_rst)); 
buffer_wire buffer_11303 (.in(n11303), .out(n11303_0));
mux3 mux_6138 (.in({n12355_0, n12354_1, n1159}), .out(n11304), .config_in(config_chain[20899:20898]), .config_rst(config_rst)); 
buffer_wire buffer_11304 (.in(n11304), .out(n11304_0));
mux13 mux_6139 (.in({n13497_0, n13484_0, n13479_0, n13470_0/**/, n13465_0, n13434_0, n13428_1, n13385_0, n11397_1, n4093, n4085, n3997, n3989}), .out(n11305), .config_in(config_chain[20905:20900]), .config_rst(config_rst)); 
buffer_wire buffer_11305 (.in(n11305), .out(n11305_0));
mux3 mux_6140 (.in({n12357_0, n12356_1, n1159}), .out(n11306), .config_in(config_chain[20907:20906]), .config_rst(config_rst)); 
buffer_wire buffer_11306 (.in(n11306), .out(n11306_0));
mux13 mux_6141 (.in({n13761_0/**/, n13757_0, n13740_0, n13726_0, n13721_0, n13712_0, n13707_0, n13690_1, n11419_1, n5071, n5063, n4975, n4967}), .out(n11307), .config_in(config_chain[20913:20908]), .config_rst(config_rst)); 
buffer_wire buffer_11307 (.in(n11307), .out(n11307_0));
mux3 mux_6142 (.in({n12359_0, n12358_1, n1159}), .out(n11308), .config_in(config_chain[20915:20914]), .config_rst(config_rst)); 
buffer_wire buffer_11308 (.in(n11308), .out(n11308_0));
mux13 mux_6143 (.in({n14027_0, n14006_0, n14001_0, n13992_0, n13987_0, n13973_0, n13956_1, n13954_1/**/, n11441_0, n6049, n6041, n5953, n5945}), .out(n11309), .config_in(config_chain[20921:20916]), .config_rst(config_rst)); 
buffer_wire buffer_11309 (.in(n11309), .out(n11309_0));
mux3 mux_6144 (.in({n12361_0, n12360_1, n1163}), .out(n11310), .config_in(config_chain[20923:20922]), .config_rst(config_rst)); 
buffer_wire buffer_11310 (.in(n11310), .out(n11310_0));
mux13 mux_6145 (.in({n14293_0, n14283_0, n14250_0, n14245_0, n14236_0, n14231_0, n14220_1, n14200_1, n11463_0/**/, n7027, n7019, n6931, n6923}), .out(n11311), .config_in(config_chain[20929:20924]), .config_rst(config_rst)); 
buffer_wire buffer_11311 (.in(n11311), .out(n11311_0));
mux16 mux_6146 (.in({n12735_0, n12708_0, n12705_0, n12682_0, n12679_0, n12673_0, n12656_0, n12652_1, n12613_0, n12604_1/**/, n11226_0, n2137, n2129, n2041, n2033, n2025}), .out(n11312), .config_in(config_chain[20935:20930]), .config_rst(config_rst)); 
buffer_wire buffer_11312 (.in(n11312), .out(n11312_0));
mux15 mux_6147 (.in({n13759_0, n13748_0, n13743_0, n13734_0, n13729_0, n13698_0, n13693_0, n13649_0, n13646_1, n11399_1, n5071, n5063/**/, n4975, n4967, n4959}), .out(n11313), .config_in(config_chain[20941:20936]), .config_rst(config_rst)); 
buffer_wire buffer_11313 (.in(n11313), .out(n11313_0));
mux16 mux_6148 (.in({n12717_0, n12702_0, n12699_0, n12693_0, n12676_0, n12670_0, n12667_0, n12650_1, n12615_0, n12606_1, n11234_0, n2137, n2129/**/, n2041, n2033, n2025}), .out(n11314), .config_in(config_chain[20947:20942]), .config_rst(config_rst)); 
buffer_wire buffer_11314 (.in(n11314), .out(n11314_0));
mux15 mux_6149 (.in({n13779_0, n13756_0, n13751_0, n13720_0, n13715_0, n13706_0, n13701_0, n13672_1, n13651_0, n11401_1, n5075, n5063, n4975, n4967, n4959}), .out(n11315), .config_in(config_chain[20953:20948]), .config_rst(config_rst)); 
buffer_wire buffer_11315 (.in(n11315), .out(n11315_0));
mux15 mux_6150 (.in({n12719_0, n12713_0, n12696_0, n12690_0, n12687_0, n12664_0/**/, n12661_0, n12648_1, n12608_1, n11242_0, n2137, n2129, n2041, n2033, n2025}), .out(n11316), .config_in(config_chain[20959:20954]), .config_rst(config_rst)); 
buffer_wire buffer_11316 (.in(n11316), .out(n11316_0));
mux15 mux_6151 (.in({n13777_0, n13742_0, n13737_0, n13728_0, n13723_0/**/, n13709_0, n13692_0, n13674_1, n13648_1, n11403_1, n5075, n5067, n4975, n4967, n4959}), .out(n11317), .config_in(config_chain[20965:20960]), .config_rst(config_rst)); 
buffer_wire buffer_11317 (.in(n11317), .out(n11317_0));
mux15 mux_6152 (.in({n12721_0, n12710_0, n12707_0, n12684_0, n12681_0, n12675_0, n12658_0, n12646_1, n12610_1, n11250_0, n2137/**/, n2129, n2041, n2033, n2025}), .out(n11318), .config_in(config_chain[20971:20966]), .config_rst(config_rst)); 
buffer_wire buffer_11318 (.in(n11318), .out(n11318_0));
mux15 mux_6153 (.in({n13775_0, n13750_0, n13745_0, n13731_0, n13714_0, n13700_0, n13695_0, n13676_1, n13650_1, n11405_1, n5075, n5067/**/, n5059, n4967, n4959}), .out(n11319), .config_in(config_chain[20977:20972]), .config_rst(config_rst)); 
buffer_wire buffer_11319 (.in(n11319), .out(n11319_0));
mux15 mux_6154 (.in({n12723_0, n12704_0, n12701_0, n12695_0, n12678_0, n12672_0/**/, n12669_0, n12644_1, n12612_1, n11258_0, n2137, n2129, n2041, n2033, n2025}), .out(n11320), .config_in(config_chain[20983:20978]), .config_rst(config_rst)); 
buffer_wire buffer_11320 (.in(n11320), .out(n11320_0));
mux14 mux_6155 (.in({n13773_0, n13753_0, n13736_0, n13722_0, n13717_0, n13708_0, n13703_0, n13678_1, n11407_1, n5075, n5067, n5059/**/, n4971, n4959}), .out(n11321), .config_in(config_chain[20989:20984]), .config_rst(config_rst)); 
buffer_wire buffer_11321 (.in(n11321), .out(n11321_0));
mux15 mux_6156 (.in({n12725_0, n12715_0/**/, n12698_0, n12692_0, n12689_0, n12666_0, n12663_0, n12642_1, n12614_1, n11266_0, n2141, n2133, n2125, n2037, n2029}), .out(n11322), .config_in(config_chain[20995:20990]), .config_rst(config_rst)); 
buffer_wire buffer_11322 (.in(n11322), .out(n11322_0));
mux14 mux_6157 (.in({n13771_0, n13744_0, n13739_0, n13730_0, n13725_0, n13711_0, n13694_0, n13680_1, n11409_1, n5075, n5067, n5059, n4971, n4963}), .out(n11323), .config_in(config_chain[21001:20996]), .config_rst(config_rst)); 
buffer_wire buffer_11323 (.in(n11323), .out(n11323_0));
mux15 mux_6158 (.in({n12727_0, n12712_0, n12709_0, n12686_0/**/, n12683_0, n12660_0, n12657_0, n12640_1, n12605_0, n11274_0, n2141, n2133, n2125, n2037, n2029}), .out(n11324), .config_in(config_chain[21007:21002]), .config_rst(config_rst)); 
buffer_wire buffer_11324 (.in(n11324), .out(n11324_0));
mux13 mux_6159 (.in({n13769_0, n13752_0, n13747_0, n13733_0, n13716_0, n13702_0, n13697_0/**/, n13682_1, n11411_1, n5067, n5059, n4971, n4963}), .out(n11325), .config_in(config_chain[21013:21008]), .config_rst(config_rst)); 
buffer_wire buffer_11325 (.in(n11325), .out(n11325_0));
mux15 mux_6160 (.in({n12729_0, n12706_0, n12703_0, n12680_0/**/, n12677_0, n12674_0, n12671_0, n12638_1, n12607_0, n11282_0, n2141, n2133, n2125, n2037, n2029}), .out(n11326), .config_in(config_chain[21019:21014]), .config_rst(config_rst)); 
buffer_wire buffer_11326 (.in(n11326), .out(n11326_0));
mux13 mux_6161 (.in({n13767_0, n13755_0, n13738_0, n13724_0, n13719_0, n13710_0, n13705_0, n13684_1, n11413_1, n5071/**/, n5059, n4971, n4963}), .out(n11327), .config_in(config_chain[21025:21020]), .config_rst(config_rst)); 
buffer_wire buffer_11327 (.in(n11327), .out(n11327_0));
mux15 mux_6162 (.in({n12731_0, n12700_0, n12697_0/**/, n12694_0, n12691_0, n12668_0, n12665_0, n12636_1, n12609_0, n11290_0, n2141, n2133, n2125, n2037, n2029}), .out(n11328), .config_in(config_chain[21031:21026]), .config_rst(config_rst)); 
buffer_wire buffer_11328 (.in(n11328), .out(n11328_0));
mux13 mux_6163 (.in({n13765_0, n13746_0, n13741_0, n13732_0, n13727_0, n13713_0, n13696_0, n13686_1, n11415_1/**/, n5071, n5063, n4971, n4963}), .out(n11329), .config_in(config_chain[21037:21032]), .config_rst(config_rst)); 
buffer_wire buffer_11329 (.in(n11329), .out(n11329_0));
mux15 mux_6164 (.in({n12733_0, n12714_0, n12711_0, n12688_0, n12685_0, n12662_0, n12659_0, n12654_1, n12611_0, n11298_0, n2141, n2133/**/, n2125, n2037, n2029}), .out(n11330), .config_in(config_chain[21043:21038]), .config_rst(config_rst)); 
buffer_wire buffer_11330 (.in(n11330), .out(n11330_0));
mux13 mux_6165 (.in({n13763_0, n13754_0, n13749_0, n13735_0, n13718_0, n13704_0, n13699_0, n13688_1/**/, n11417_1, n5071, n5063, n4975, n4963}), .out(n11331), .config_in(config_chain[21049:21044]), .config_rst(config_rst)); 
buffer_wire buffer_11331 (.in(n11331), .out(n11331_0));
mux15 mux_6166 (.in({n12993_0, n12965_0, n12958_0, n12946_0, n12919_0, n12912_0, n12910_1, n12868_1, n12865_0, n11220_0, n3115, n3107, n3019, n3011, n3003}), .out(n11332), .config_in(config_chain[21055:21050]), .config_rst(config_rst)); 
buffer_wire buffer_11332 (.in(n11332), .out(n11332_0));
mux15 mux_6167 (.in({n14025_0, n14023_0, n14014_0, n14009_0, n13995_0, n13978_0, n13964_0, n13959_0, n13912_1, n11421_0, n6049, n6041/**/, n5953, n5945, n5937}), .out(n11333), .config_in(config_chain[21061:21056]), .config_rst(config_rst)); 
buffer_wire buffer_11333 (.in(n11333), .out(n11333_0));
mux15 mux_6168 (.in({n12973_0, n12966_0, n12939_0, n12932_0, n12927_0, n12920_0/**/, n12908_1, n12870_1, n12867_0, n11228_0, n3119, n3107, n3019, n3011, n3003}), .out(n11334), .config_in(config_chain[21067:21062]), .config_rst(config_rst)); 
buffer_wire buffer_11334 (.in(n11334), .out(n11334_0));
mux15 mux_6169 (.in({n14045_0, n14017_0, n14000_0, n13986_0, n13981_0, n13972_0, n13967_0, n13936_1/**/, n13915_0, n11423_0, n6053, n6041, n5953, n5945, n5937}), .out(n11335), .config_in(config_chain[21073:21068]), .config_rst(config_rst)); 
buffer_wire buffer_11335 (.in(n11335), .out(n11335_0));
mux15 mux_6170 (.in({n12975_0, n12959_0, n12952_0, n12947_0, n12940_0/**/, n12928_0, n12913_0, n12906_1, n12869_0, n11236_0, n3119, n3111, n3019, n3011, n3003}), .out(n11336), .config_in(config_chain[21079:21074]), .config_rst(config_rst)); 
buffer_wire buffer_11336 (.in(n11336), .out(n11336_0));
mux15 mux_6171 (.in({n14043_0, n14022_0, n14008_0, n14003_0, n13994_0, n13989_0, n13975_0, n13958_0, n13938_1, n11425_0, n6053, n6045/**/, n5953, n5945, n5937}), .out(n11337), .config_in(config_chain[21085:21080]), .config_rst(config_rst)); 
buffer_wire buffer_11337 (.in(n11337), .out(n11337_0));
mux15 mux_6172 (.in({n12977_0, n12967_0, n12960_0, n12948_0, n12933_0/**/, n12921_0, n12914_0, n12904_1, n12871_0, n11244_0, n3119, n3111, n3103, n3011, n3003}), .out(n11338), .config_in(config_chain[21091:21086]), .config_rst(config_rst)); 
buffer_wire buffer_11338 (.in(n11338), .out(n11338_0));
mux15 mux_6173 (.in({n14041_0, n14016_0, n14011_0, n13997_0, n13980_0, n13966_0/**/, n13961_0, n13940_1, n13914_1, n11427_0, n6053, n6045, n6037, n5945, n5937}), .out(n11339), .config_in(config_chain[21097:21092]), .config_rst(config_rst)); 
buffer_wire buffer_11339 (.in(n11339), .out(n11339_0));
mux14 mux_6174 (.in({n12979_0/**/, n12968_0, n12953_0, n12941_0, n12934_0, n12929_0, n12922_0, n12902_1, n11252_0, n3119, n3111, n3103, n3015, n3003}), .out(n11340), .config_in(config_chain[21103:21098]), .config_rst(config_rst)); 
buffer_wire buffer_11340 (.in(n11340), .out(n11340_0));
mux14 mux_6175 (.in({n14039_0, n14019_0, n14002_0, n13988_0, n13983_0, n13974_0, n13969_0, n13942_1, n11429_0, n6053, n6045, n6037, n5949, n5937/**/}), .out(n11341), .config_in(config_chain[21109:21104]), .config_rst(config_rst)); 
buffer_wire buffer_11341 (.in(n11341), .out(n11341_0));
mux14 mux_6176 (.in({n12981_0, n12961_0, n12954_0, n12949_0, n12942_0/**/, n12930_0, n12915_0, n12900_1, n11260_0, n3119, n3111, n3103, n3015, n3007}), .out(n11342), .config_in(config_chain[21115:21110]), .config_rst(config_rst)); 
buffer_wire buffer_11342 (.in(n11342), .out(n11342_0));
mux14 mux_6177 (.in({n14037_0, n14010_0, n14005_0, n13996_0, n13991_0, n13977_0, n13960_0, n13944_1/**/, n11431_0, n6053, n6045, n6037, n5949, n5941}), .out(n11343), .config_in(config_chain[21121:21116]), .config_rst(config_rst)); 
buffer_wire buffer_11343 (.in(n11343), .out(n11343_0));
mux13 mux_6178 (.in({n12983_0, n12969_0, n12962_0, n12950_0, n12935_0, n12923_0, n12916_0, n12898_1, n11268_0/**/, n3111, n3103, n3015, n3007}), .out(n11344), .config_in(config_chain[21127:21122]), .config_rst(config_rst)); 
buffer_wire buffer_11344 (.in(n11344), .out(n11344_0));
mux13 mux_6179 (.in({n14035_0, n14018_0, n14013_0, n13999_0, n13982_0, n13968_0, n13963_0, n13946_1/**/, n11433_0, n6045, n6037, n5949, n5941}), .out(n11345), .config_in(config_chain[21133:21128]), .config_rst(config_rst)); 
buffer_wire buffer_11345 (.in(n11345), .out(n11345_0));
mux13 mux_6180 (.in({n12985_0, n12970_0, n12955_0, n12943_0/**/, n12936_0, n12931_0, n12924_0, n12896_1, n11276_0, n3115, n3103, n3015, n3007}), .out(n11346), .config_in(config_chain[21139:21134]), .config_rst(config_rst)); 
buffer_wire buffer_11346 (.in(n11346), .out(n11346_0));
mux13 mux_6181 (.in({n14033_0, n14021_0, n14004_0, n13990_0, n13985_0, n13976_0, n13971_0, n13948_1/**/, n11435_0, n6049, n6037, n5949, n5941}), .out(n11347), .config_in(config_chain[21145:21140]), .config_rst(config_rst)); 
buffer_wire buffer_11347 (.in(n11347), .out(n11347_0));
mux13 mux_6182 (.in({n12987_0, n12963_0, n12956_0, n12951_0, n12944_0, n12917_0, n12894_1, n12862_1, n11284_0/**/, n3115, n3107, n3015, n3007}), .out(n11348), .config_in(config_chain[21151:21146]), .config_rst(config_rst)); 
buffer_wire buffer_11348 (.in(n11348), .out(n11348_0));
mux13 mux_6183 (.in({n14031_0, n14012_0, n14007_0, n13998_0, n13993_0, n13962_0, n13957_0, n13950_1, n11437_0, n6049, n6041/**/, n5949, n5941}), .out(n11349), .config_in(config_chain[21157:21152]), .config_rst(config_rst)); 
buffer_wire buffer_11349 (.in(n11349), .out(n11349_0));
mux13 mux_6184 (.in({n12989_0, n12971_0, n12964_0, n12937_0, n12925_0/**/, n12918_0, n12892_1, n12864_1, n11292_0, n3115, n3107, n3019, n3007}), .out(n11350), .config_in(config_chain[21163:21158]), .config_rst(config_rst)); 
buffer_wire buffer_11350 (.in(n11350), .out(n11350_0));
mux13 mux_6185 (.in({n14029_0, n14020_0, n14015_0, n13984_0, n13979_0, n13970_0, n13965_0, n13952_1, n11439_0/**/, n6049, n6041, n5953, n5941}), .out(n11351), .config_in(config_chain[21169:21164]), .config_rst(config_rst)); 
buffer_wire buffer_11351 (.in(n11351), .out(n11351_0));
mux13 mux_6186 (.in({n12991_0/**/, n12957_0, n12945_0, n12938_0, n12926_0, n12866_1, n12863_0, n12860_1, n11300_0, n3115, n3107, n3019, n3011}), .out(n11352), .config_in(config_chain[21175:21170]), .config_rst(config_rst)); 
buffer_wire buffer_11352 (.in(n11352), .out(n11352_0));
mux3 mux_6187 (.in({n14695_0, n14694_1, n8983}), .out(n11353), .config_in(config_chain[21177:21176]), .config_rst(config_rst)); 
buffer_wire buffer_11353 (.in(n11353), .out(n11353_0));
mux15 mux_6188 (.in({n13253_0, n13217_0, n13210_0, n13203_0, n13196_0/**/, n13184_0, n13168_1, n13126_1, n13123_0, n11222_0, n4093, n4085, n3997, n3989, n3981}), .out(n11354), .config_in(config_chain[21183:21178]), .config_rst(config_rst)); 
buffer_wire buffer_11354 (.in(n11354), .out(n11354_0));
mux15 mux_6189 (.in({n14291_0, n14274_0, n14269_0, n14267_0, n14258_0/**/, n14253_0, n14239_0, n14222_1, n14178_1, n11443_0, n7027, n7019, n6931, n6923, n6915}), .out(n11355), .config_in(config_chain[21189:21184]), .config_rst(config_rst)); 
buffer_wire buffer_11355 (.in(n11355), .out(n11355_0));
mux15 mux_6190 (.in({n13233_0, n13225_0/**/, n13218_0, n13204_0, n13177_0, n13170_0, n13166_1, n13128_1, n13125_0, n11230_0, n4097, n4085, n3997, n3989, n3981}), .out(n11356), .config_in(config_chain[21195:21190]), .config_rst(config_rst)); 
buffer_wire buffer_11356 (.in(n11356), .out(n11356_0));
mux15 mux_6191 (.in({n14311_0, n14289_0, n14282_0, n14277_0, n14261_0, n14244_0, n14230_0, n14225_0, n14202_1, n11445_0/**/, n7031, n7019, n6931, n6923, n6915}), .out(n11357), .config_in(config_chain[21201:21196]), .config_rst(config_rst)); 
buffer_wire buffer_11357 (.in(n11357), .out(n11357_0));
mux15 mux_6192 (.in({n13235_0, n13226_0/**/, n13211_0, n13197_0, n13190_0, n13185_0, n13178_0, n13164_1, n13127_0, n11238_0, n4097, n4089, n3997, n3989, n3981}), .out(n11358), .config_in(config_chain[21207:21202]), .config_rst(config_rst)); 
buffer_wire buffer_11358 (.in(n11358), .out(n11358_0));
mux15 mux_6193 (.in({n14309_0, n14285_0, n14268_0, n14266_0/**/, n14252_0, n14247_0, n14238_0, n14233_0, n14204_1, n11447_0, n7031, n7023, n6931, n6923, n6915}), .out(n11359), .config_in(config_chain[21213:21208]), .config_rst(config_rst)); 
buffer_wire buffer_11359 (.in(n11359), .out(n11359_0));
mux15 mux_6194 (.in({n13237_0, n13219_0, n13212_0, n13205_0, n13198_0, n13186_0, n13171_0/**/, n13162_1, n13129_0, n11246_0, n4097, n4089, n4081, n3989, n3981}), .out(n11360), .config_in(config_chain[21219:21214]), .config_rst(config_rst)); 
buffer_wire buffer_11360 (.in(n11360), .out(n11360_0));
mux15 mux_6195 (.in({n14307_0, n14288_0, n14276_0, n14271_0, n14260_0, n14255_0, n14241_0, n14224_0, n14206_1, n11449_0, n7031, n7023/**/, n7015, n6923, n6915}), .out(n11361), .config_in(config_chain[21225:21220]), .config_rst(config_rst)); 
buffer_wire buffer_11361 (.in(n11361), .out(n11361_0));
mux14 mux_6196 (.in({n13239_0, n13227_0, n13220_0, n13206_0, n13191_0/**/, n13179_0, n13172_0, n13160_1, n11254_0, n4097, n4089, n4081, n3993, n3981}), .out(n11362), .config_in(config_chain[21231:21226]), .config_rst(config_rst)); 
buffer_wire buffer_11362 (.in(n11362), .out(n11362_0));
mux14 mux_6197 (.in({n14305_0, n14284_0, n14279_0, n14263_0, n14246_0, n14232_0, n14227_0, n14208_1, n11451_0/**/, n7031, n7023, n7015, n6927, n6915}), .out(n11363), .config_in(config_chain[21237:21232]), .config_rst(config_rst)); 
buffer_wire buffer_11363 (.in(n11363), .out(n11363_0));
mux14 mux_6198 (.in({n13241_0, n13228_0, n13213_0, n13199_0, n13192_0, n13187_0, n13180_0, n13158_1, n11262_0, n4097, n4089/**/, n4081, n3993, n3985}), .out(n11364), .config_in(config_chain[21243:21238]), .config_rst(config_rst)); 
buffer_wire buffer_11364 (.in(n11364), .out(n11364_0));
mux14 mux_6199 (.in({n14303_0, n14287_0, n14270_0, n14254_0, n14249_0, n14240_0, n14235_0, n14210_1, n11453_0, n7031, n7023, n7015, n6927, n6919}), .out(n11365), .config_in(config_chain[21249:21244]), .config_rst(config_rst)); 
buffer_wire buffer_11365 (.in(n11365), .out(n11365_0));
mux13 mux_6200 (.in({n13243_0, n13221_0, n13214_0, n13207_0, n13200_0, n13188_0, n13173_0/**/, n13156_1, n11270_0, n4089, n4081, n3993, n3985}), .out(n11366), .config_in(config_chain[21255:21250]), .config_rst(config_rst)); 
buffer_wire buffer_11366 (.in(n11366), .out(n11366_0));
mux13 mux_6201 (.in({n14301_0, n14278_0, n14273_0, n14262_0, n14257_0, n14243_0, n14226_0, n14212_1, n11455_0, n7023, n7015, n6927, n6919/**/}), .out(n11367), .config_in(config_chain[21261:21256]), .config_rst(config_rst)); 
buffer_wire buffer_11367 (.in(n11367), .out(n11367_0));
mux13 mux_6202 (.in({n13245_0, n13229_0, n13222_0, n13208_0, n13193_0, n13181_0, n13174_0, n13154_1/**/, n11278_0, n4093, n4081, n3993, n3985}), .out(n11368), .config_in(config_chain[21267:21262]), .config_rst(config_rst)); 
buffer_wire buffer_11368 (.in(n11368), .out(n11368_0));
mux13 mux_6203 (.in({n14299_0, n14286_0, n14281_0, n14265_0, n14248_0, n14234_0, n14229_0, n14214_1/**/, n11457_0, n7027, n7015, n6927, n6919}), .out(n11369), .config_in(config_chain[21273:21268]), .config_rst(config_rst)); 
buffer_wire buffer_11369 (.in(n11369), .out(n11369_0));
mux13 mux_6204 (.in({n13247_0, n13230_0, n13215_0, n13201_0, n13194_0, n13189_0, n13182_0, n13152_1/**/, n11286_0, n4093, n4085, n3993, n3985}), .out(n11370), .config_in(config_chain[21279:21274]), .config_rst(config_rst)); 
buffer_wire buffer_11370 (.in(n11370), .out(n11370_0));
mux13 mux_6205 (.in({n14297_0, n14272_0, n14256_0, n14251_0, n14242_0, n14237_0, n14216_1, n14201_0, n11459_0/**/, n7027, n7019, n6927, n6919}), .out(n11371), .config_in(config_chain[21285:21280]), .config_rst(config_rst)); 
buffer_wire buffer_11371 (.in(n11371), .out(n11371_0));
mux13 mux_6206 (.in({n13249_0, n13223_0, n13216_0, n13209_0, n13202_0, n13175_0, n13150_1/**/, n13122_1, n11294_0, n4093, n4085, n3997, n3985}), .out(n11372), .config_in(config_chain[21291:21286]), .config_rst(config_rst)); 
buffer_wire buffer_11372 (.in(n11372), .out(n11372_0));
mux13 mux_6207 (.in({n14295_0, n14280_0, n14275_0, n14264_0/**/, n14259_0, n14228_0, n14223_0, n14218_1, n11461_0, n7027, n7019, n6931, n6919}), .out(n11373), .config_in(config_chain[21297:21292]), .config_rst(config_rst)); 
buffer_wire buffer_11373 (.in(n11373), .out(n11373_0));
mux13 mux_6208 (.in({n13251_0, n13231_0, n13224_0, n13195_0, n13183_0, n13176_0, n13124_1, n13120_1, n11302_0, n4093, n4085/**/, n3997, n3989}), .out(n11374), .config_in(config_chain[21303:21298]), .config_rst(config_rst)); 
buffer_wire buffer_11374 (.in(n11374), .out(n11374_0));
mux3 mux_6209 (.in({n14697_0, n14696_1, n8983}), .out(n11375), .config_in(config_chain[21305:21304]), .config_rst(config_rst)); 
buffer_wire buffer_11375 (.in(n11375), .out(n11375_0));
mux15 mux_6210 (.in({n13515_0, n13493_0, n13486_0, n13457_0, n13450_0, n13443_0, n13436_0, n13428_1, n13386_1, n11224_1, n5071, n5063, n4975/**/, n4967, n4959}), .out(n11376), .config_in(config_chain[21311:21306]), .config_rst(config_rst)); 
buffer_wire buffer_11376 (.in(n11376), .out(n11376_0));
mux16 mux_6211 (.in({n14555_0, n14539_0, n14534_0/**/, n14530_0, n14526_0, n14511_0, n14501_0, n14496_0, n14484_1, n14433_0, n11465_0, n8005, n7997, n7909, n7901, n7893}), .out(n11377), .config_in(config_chain[21317:21312]), .config_rst(config_rst)); 
buffer_wire buffer_11377 (.in(n11377), .out(n11377_0));
mux15 mux_6212 (.in({n13495_0, n13479_0, n13472_0/**/, n13465_0, n13458_0, n13444_0, n13426_1, n13388_1, n13385_0, n11232_1, n5075, n5063, n4975, n4967, n4959}), .out(n11378), .config_in(config_chain[21323:21318]), .config_rst(config_rst)); 
buffer_wire buffer_11378 (.in(n11378), .out(n11378_0));
mux16 mux_6213 (.in({n14573_0, n14552_0, n14548_0, n14533_0, n14525_0, n14520_0, n14495_0, n14490_0, n14466_1, n14465_0, n11467_0/**/, n8005, n7997, n7909, n7901, n7893}), .out(n11379), .config_in(config_chain[21329:21324]), .config_rst(config_rst)); 
buffer_wire buffer_11379 (.in(n11379), .out(n11379_0));
mux15 mux_6214 (.in({n13497_0, n13487_0, n13480_0, n13466_0, n13451_0, n13437_0/**/, n13430_0, n13424_1, n13387_0, n11240_1, n5075, n5067, n4975, n4967, n4959}), .out(n11380), .config_in(config_chain[21335:21330]), .config_rst(config_rst)); 
buffer_wire buffer_11380 (.in(n11380), .out(n11380_0));
mux15 mux_6215 (.in({n14571_0, n14547_0, n14542_0, n14519_0, n14514_0, n14504_0, n14489_0, n14487_0, n14468_1, n11469_0, n8005/**/, n7997, n7909, n7901, n7893}), .out(n11381), .config_in(config_chain[21341:21336]), .config_rst(config_rst)); 
buffer_wire buffer_11381 (.in(n11381), .out(n11381_0));
mux15 mux_6216 (.in({n13499_0, n13488_0, n13473_0, n13459_0, n13452_0, n13445_0, n13438_0, n13422_1/**/, n13389_0, n11248_1, n5075, n5067, n5059, n4967, n4959}), .out(n11382), .config_in(config_chain[21347:21342]), .config_rst(config_rst)); 
buffer_wire buffer_11382 (.in(n11382), .out(n11382_0));
mux15 mux_6217 (.in({n14569_0, n14541_0, n14536_0/**/, n14528_0, n14513_0, n14509_0, n14503_0, n14498_0, n14470_1, n11471_0, n8005, n7997, n7909, n7901, n7893}), .out(n11383), .config_in(config_chain[21353:21348]), .config_rst(config_rst)); 
buffer_wire buffer_11383 (.in(n11383), .out(n11383_0));
mux14 mux_6218 (.in({n13501_0, n13481_0, n13474_0, n13467_0, n13460_0, n13446_0, n13431_0, n13420_1, n11256_1, n5075, n5067, n5059/**/, n4971, n4959}), .out(n11384), .config_in(config_chain[21359:21354]), .config_rst(config_rst)); 
buffer_wire buffer_11384 (.in(n11384), .out(n11384_0));
mux15 mux_6219 (.in({n14567_0, n14550_0/**/, n14535_0, n14531_0, n14527_0, n14522_0, n14497_0, n14492_0, n14472_1, n11473_0, n8005, n7997, n7909, n7901, n7893}), .out(n11385), .config_in(config_chain[21365:21360]), .config_rst(config_rst)); 
buffer_wire buffer_11385 (.in(n11385), .out(n11385_0));
mux14 mux_6220 (.in({n13503_0, n13489_0, n13482_0, n13468_0, n13453_0, n13439_0, n13432_0/**/, n13418_1, n11264_1, n5075, n5067, n5059, n4971, n4963}), .out(n11386), .config_in(config_chain[21371:21366]), .config_rst(config_rst)); 
buffer_wire buffer_11386 (.in(n11386), .out(n11386_0));
mux15 mux_6221 (.in({n14565_0/**/, n14553_0, n14549_0, n14544_0, n14521_0, n14516_0, n14506_0, n14491_0, n14474_1, n11475_0, n8009, n8001, n7993, n7905, n7897}), .out(n11387), .config_in(config_chain[21377:21372]), .config_rst(config_rst)); 
buffer_wire buffer_11387 (.in(n11387), .out(n11387_0));
mux13 mux_6222 (.in({n13505_0, n13490_0, n13475_0, n13461_0/**/, n13454_0, n13447_0, n13440_0, n13416_1, n11272_1, n5067, n5059, n4971, n4963}), .out(n11388), .config_in(config_chain[21383:21378]), .config_rst(config_rst)); 
buffer_wire buffer_11388 (.in(n11388), .out(n11388_0));
mux15 mux_6223 (.in({n14563_0/**/, n14543_0, n14538_0, n14515_0, n14510_0, n14505_0, n14500_0, n14476_1, n14432_1, n11477_0, n8009, n8001, n7993, n7905, n7897}), .out(n11389), .config_in(config_chain[21389:21384]), .config_rst(config_rst)); 
buffer_wire buffer_11389 (.in(n11389), .out(n11389_0));
mux13 mux_6224 (.in({n13507_0, n13483_0, n13476_0, n13469_0, n13462_0, n13448_0, n13433_0, n13414_1, n11280_1, n5071, n5059, n4971/**/, n4963}), .out(n11390), .config_in(config_chain[21395:21390]), .config_rst(config_rst)); 
buffer_wire buffer_11390 (.in(n11390), .out(n11390_0));
mux15 mux_6225 (.in({n14561_0, n14537_0/**/, n14532_0, n14529_0, n14524_0, n14499_0, n14494_0, n14478_1, n14464_1, n11479_0, n8009, n8001, n7993, n7905, n7897}), .out(n11391), .config_in(config_chain[21401:21396]), .config_rst(config_rst)); 
buffer_wire buffer_11391 (.in(n11391), .out(n11391_0));
mux13 mux_6226 (.in({n13509_0/**/, n13491_0, n13484_0, n13470_0, n13455_0, n13441_0, n13434_0, n13412_1, n11288_1, n5071, n5063, n4971, n4963}), .out(n11392), .config_in(config_chain[21407:21402]), .config_rst(config_rst)); 
buffer_wire buffer_11392 (.in(n11392), .out(n11392_0));
mux15 mux_6227 (.in({n14559_0, n14551_0, n14546_0, n14523_0, n14518_0/**/, n14493_0, n14488_0, n14486_1, n14480_1, n11481_0, n8009, n8001, n7993, n7905, n7897}), .out(n11393), .config_in(config_chain[21413:21408]), .config_rst(config_rst)); 
buffer_wire buffer_11393 (.in(n11393), .out(n11393_0));
mux13 mux_6228 (.in({n13511_0/**/, n13492_0, n13477_0, n13463_0, n13456_0, n13449_0, n13442_0, n13410_1, n11296_1, n5071, n5063, n4975, n4963}), .out(n11394), .config_in(config_chain[21419:21414]), .config_rst(config_rst)); 
buffer_wire buffer_11394 (.in(n11394), .out(n11394_0));
mux15 mux_6229 (.in({n14557_0, n14545_0, n14540_0, n14517_0, n14512_0/**/, n14508_0, n14507_0, n14502_0, n14482_1, n11483_0, n8009, n8001, n7993, n7905, n7897}), .out(n11395), .config_in(config_chain[21425:21420]), .config_rst(config_rst)); 
buffer_wire buffer_11395 (.in(n11395), .out(n11395_0));
mux13 mux_6230 (.in({n13513_0, n13485_0, n13478_0/**/, n13471_0, n13464_0, n13435_0, n13384_1, n13382_1, n11304_1, n5071, n5063, n4975, n4967}), .out(n11396), .config_in(config_chain[21431:21426]), .config_rst(config_rst)); 
buffer_wire buffer_11396 (.in(n11396), .out(n11396_0));
mux3 mux_6231 (.in({n14727_0, n14726_1, n8983}), .out(n11397), .config_in(config_chain[21433:21432]), .config_rst(config_rst)); 
buffer_wire buffer_11397 (.in(n11397), .out(n11397_0));
mux15 mux_6232 (.in({n13779_0, n13749_0, n13742_0, n13735_0, n13728_0, n13699_0, n13692_0, n13690_1, n13648_1, n11312_1, n6049, n6041, n5953, n5945, n5937/**/}), .out(n11398), .config_in(config_chain[21439:21434]), .config_rst(config_rst)); 
buffer_wire buffer_11398 (.in(n11398), .out(n11398_0));
mux4 mux_6233 (.in({n14815_0, n14728_1, n8987, n8871}), .out(n11399), .config_in(config_chain[21441:21440]), .config_rst(config_rst)); 
buffer_wire buffer_11399 (.in(n11399), .out(n11399_0));
mux15 mux_6234 (.in({n13759_0/**/, n13757_0, n13750_0, n13721_0, n13714_0, n13707_0, n13700_0, n13688_1, n13650_1, n11314_1, n6053, n6041, n5953, n5945, n5937}), .out(n11400), .config_in(config_chain[21447:21442]), .config_rst(config_rst)); 
buffer_wire buffer_11400 (.in(n11400), .out(n11400_0));
mux3 mux_6235 (.in({n14817_0, n14730_1, n8875}), .out(n11401), .config_in(config_chain[21449:21448]), .config_rst(config_rst)); 
buffer_wire buffer_11401 (.in(n11401), .out(n11401_0));
mux15 mux_6236 (.in({n13761_0, n13743_0, n13736_0, n13729_0, n13722_0, n13708_0, n13693_0/**/, n13686_1, n13649_0, n11316_1, n6053, n6045, n5953, n5945, n5937}), .out(n11402), .config_in(config_chain[21455:21450]), .config_rst(config_rst)); 
buffer_wire buffer_11402 (.in(n11402), .out(n11402_0));
mux3 mux_6237 (.in({n14819_0, n14732_1/**/, n8879}), .out(n11403), .config_in(config_chain[21457:21456]), .config_rst(config_rst)); 
buffer_wire buffer_11403 (.in(n11403), .out(n11403_0));
mux15 mux_6238 (.in({n13763_0, n13751_0, n13744_0/**/, n13730_0, n13715_0, n13701_0, n13694_0, n13684_1, n13651_0, n11318_1, n6053, n6045, n6037, n5945, n5937}), .out(n11404), .config_in(config_chain[21463:21458]), .config_rst(config_rst)); 
buffer_wire buffer_11404 (.in(n11404), .out(n11404_0));
mux3 mux_6239 (.in({n14821_0, n14734_1/**/, n8883}), .out(n11405), .config_in(config_chain[21465:21464]), .config_rst(config_rst)); 
buffer_wire buffer_11405 (.in(n11405), .out(n11405_0));
mux14 mux_6240 (.in({n13765_0, n13752_0, n13737_0, n13723_0, n13716_0, n13709_0, n13702_0, n13682_1, n11320_1/**/, n6053, n6045, n6037, n5949, n5937}), .out(n11406), .config_in(config_chain[21471:21466]), .config_rst(config_rst)); 
buffer_wire buffer_11406 (.in(n11406), .out(n11406_0));
mux3 mux_6241 (.in({n14823_0, n14736_1/**/, n8883}), .out(n11407), .config_in(config_chain[21473:21472]), .config_rst(config_rst)); 
buffer_wire buffer_11407 (.in(n11407), .out(n11407_0));
mux14 mux_6242 (.in({n13767_0/**/, n13745_0, n13738_0, n13731_0, n13724_0, n13710_0, n13695_0, n13680_1, n11322_1, n6053, n6045, n6037, n5949, n5941}), .out(n11408), .config_in(config_chain[21479:21474]), .config_rst(config_rst)); 
buffer_wire buffer_11408 (.in(n11408), .out(n11408_0));
mux3 mux_6243 (.in({n14825_0, n14738_1, n8887}), .out(n11409), .config_in(config_chain[21481:21480]), .config_rst(config_rst)); 
buffer_wire buffer_11409 (.in(n11409), .out(n11409_0));
mux13 mux_6244 (.in({n13769_0, n13753_0, n13746_0, n13732_0, n13717_0, n13703_0, n13696_0, n13678_1, n11324_1, n6045, n6037, n5949, n5941/**/}), .out(n11410), .config_in(config_chain[21487:21482]), .config_rst(config_rst)); 
buffer_wire buffer_11410 (.in(n11410), .out(n11410_0));
mux3 mux_6245 (.in({n14827_0, n14740_1, n8971}), .out(n11411), .config_in(config_chain[21489:21488]), .config_rst(config_rst)); 
buffer_wire buffer_11411 (.in(n11411), .out(n11411_0));
mux13 mux_6246 (.in({n13771_0, n13754_0, n13739_0, n13725_0, n13718_0, n13711_0, n13704_0, n13676_1, n11326_1, n6049/**/, n6037, n5949, n5941}), .out(n11412), .config_in(config_chain[21495:21490]), .config_rst(config_rst)); 
buffer_wire buffer_11412 (.in(n11412), .out(n11412_0));
mux3 mux_6247 (.in({n14829_0, n14742_1/**/, n8975}), .out(n11413), .config_in(config_chain[21497:21496]), .config_rst(config_rst)); 
buffer_wire buffer_11413 (.in(n11413), .out(n11413_0));
mux13 mux_6248 (.in({n13773_0, n13747_0, n13740_0, n13733_0, n13726_0, n13712_0, n13697_0, n13674_1, n11328_1, n6049/**/, n6041, n5949, n5941}), .out(n11414), .config_in(config_chain[21503:21498]), .config_rst(config_rst)); 
buffer_wire buffer_11414 (.in(n11414), .out(n11414_0));
mux3 mux_6249 (.in({n14831_0, n14744_1, n8979/**/}), .out(n11415), .config_in(config_chain[21505:21504]), .config_rst(config_rst)); 
buffer_wire buffer_11415 (.in(n11415), .out(n11415_0));
mux13 mux_6250 (.in({n13775_0, n13755_0, n13748_0, n13734_0, n13719_0, n13705_0, n13698_0, n13672_1, n11330_1, n6049, n6041/**/, n5953, n5941}), .out(n11416), .config_in(config_chain[21511:21506]), .config_rst(config_rst)); 
buffer_wire buffer_11416 (.in(n11416), .out(n11416_0));
mux3 mux_6251 (.in({n14833_0, n14746_1, n8979/**/}), .out(n11417), .config_in(config_chain[21513:21512]), .config_rst(config_rst)); 
buffer_wire buffer_11417 (.in(n11417), .out(n11417_0));
mux13 mux_6252 (.in({n13777_0, n13756_0, n13741_0, n13727_0/**/, n13720_0, n13713_0, n13706_0, n13646_1, n11306_1, n6049, n6041, n5953, n5945}), .out(n11418), .config_in(config_chain[21519:21514]), .config_rst(config_rst)); 
buffer_wire buffer_11418 (.in(n11418), .out(n11418_0));
mux3 mux_6253 (.in({n14749_0, n14748_1, n8983}), .out(n11419), .config_in(config_chain[21521:21520]), .config_rst(config_rst)); 
buffer_wire buffer_11419 (.in(n11419), .out(n11419_0));
mux15 mux_6254 (.in({n14045_0, n14022_0, n14015_0, n14008_0, n13994_0, n13979_0, n13965_0, n13958_0, n13954_1, n11332_1, n7027/**/, n7019, n6931, n6923, n6915}), .out(n11420), .config_in(config_chain[21527:21522]), .config_rst(config_rst)); 
buffer_wire buffer_11420 (.in(n11420), .out(n11420_0));
mux4 mux_6255 (.in({n14751_0, n14750_0, n8987, n8871}), .out(n11421), .config_in(config_chain[21529:21528]), .config_rst(config_rst)); 
buffer_wire buffer_11421 (.in(n11421), .out(n11421_0));
mux15 mux_6256 (.in({n14025_0, n14016_0/**/, n14001_0, n13987_0, n13980_0, n13973_0, n13966_0, n13952_1, n13914_1, n11334_1, n7031, n7019, n6931, n6923, n6915}), .out(n11422), .config_in(config_chain[21535:21530]), .config_rst(config_rst)); 
buffer_wire buffer_11422 (.in(n11422), .out(n11422_0));
mux3 mux_6257 (.in({n14753_0, n14752_0/**/, n8871}), .out(n11423), .config_in(config_chain[21537:21536]), .config_rst(config_rst)); 
buffer_wire buffer_11423 (.in(n11423), .out(n11423_0));
mux15 mux_6258 (.in({n14027_0, n14023_0, n14009_0, n14002_0, n13995_0, n13988_0, n13974_0, n13959_0, n13950_1/**/, n11336_1, n7031, n7023, n6931, n6923, n6915}), .out(n11424), .config_in(config_chain[21543:21538]), .config_rst(config_rst)); 
buffer_wire buffer_11424 (.in(n11424), .out(n11424_0));
mux3 mux_6259 (.in({n14755_0, n14754_0, n8875}), .out(n11425), .config_in(config_chain[21545:21544]), .config_rst(config_rst)); 
buffer_wire buffer_11425 (.in(n11425), .out(n11425_0));
mux15 mux_6260 (.in({n14029_0, n14017_0, n14010_0, n13996_0, n13981_0, n13967_0, n13960_0/**/, n13948_1, n13915_0, n11338_1, n7031, n7023, n7015, n6923, n6915}), .out(n11426), .config_in(config_chain[21551:21546]), .config_rst(config_rst)); 
buffer_wire buffer_11426 (.in(n11426), .out(n11426_0));
mux3 mux_6261 (.in({n14757_0, n14756_0, n8879/**/}), .out(n11427), .config_in(config_chain[21553:21552]), .config_rst(config_rst)); 
buffer_wire buffer_11427 (.in(n11427), .out(n11427_0));
mux14 mux_6262 (.in({n14031_0, n14018_0, n14003_0, n13989_0, n13982_0/**/, n13975_0, n13968_0, n13946_1, n11340_1, n7031, n7023, n7015, n6927, n6915}), .out(n11428), .config_in(config_chain[21559:21554]), .config_rst(config_rst)); 
buffer_wire buffer_11428 (.in(n11428), .out(n11428_0));
mux3 mux_6263 (.in({n14759_0, n14758_0, n8883}), .out(n11429), .config_in(config_chain[21561:21560]), .config_rst(config_rst)); 
buffer_wire buffer_11429 (.in(n11429), .out(n11429_0));
mux14 mux_6264 (.in({n14033_0, n14011_0, n14004_0, n13997_0, n13990_0, n13976_0, n13961_0, n13944_1, n11342_1, n7031/**/, n7023, n7015, n6927, n6919}), .out(n11430), .config_in(config_chain[21567:21562]), .config_rst(config_rst)); 
buffer_wire buffer_11430 (.in(n11430), .out(n11430_0));
mux3 mux_6265 (.in({n14761_0, n14760_0/**/, n8887}), .out(n11431), .config_in(config_chain[21569:21568]), .config_rst(config_rst)); 
buffer_wire buffer_11431 (.in(n11431), .out(n11431_0));
mux13 mux_6266 (.in({n14035_0, n14019_0, n14012_0, n13998_0, n13983_0, n13969_0, n13962_0, n13942_1, n11344_1/**/, n7023, n7015, n6927, n6919}), .out(n11432), .config_in(config_chain[21575:21570]), .config_rst(config_rst)); 
buffer_wire buffer_11432 (.in(n11432), .out(n11432_0));
mux3 mux_6267 (.in({n14763_0, n14762_0/**/, n8887}), .out(n11433), .config_in(config_chain[21577:21576]), .config_rst(config_rst)); 
buffer_wire buffer_11433 (.in(n11433), .out(n11433_0));
mux13 mux_6268 (.in({n14037_0, n14020_0, n14005_0, n13991_0, n13984_0, n13977_0, n13970_0, n13940_1, n11346_1, n7027, n7015, n6927, n6919/**/}), .out(n11434), .config_in(config_chain[21583:21578]), .config_rst(config_rst)); 
buffer_wire buffer_11434 (.in(n11434), .out(n11434_0));
mux3 mux_6269 (.in({n14765_0, n14764_0/**/, n8971}), .out(n11435), .config_in(config_chain[21585:21584]), .config_rst(config_rst)); 
buffer_wire buffer_11435 (.in(n11435), .out(n11435_0));
mux13 mux_6270 (.in({n14039_0, n14013_0, n14006_0, n13999_0, n13992_0, n13963_0, n13956_1, n13938_1, n11348_1/**/, n7027, n7019, n6927, n6919}), .out(n11436), .config_in(config_chain[21591:21586]), .config_rst(config_rst)); 
buffer_wire buffer_11436 (.in(n11436), .out(n11436_0));
mux3 mux_6271 (.in({n14767_0, n14766_0/**/, n8975}), .out(n11437), .config_in(config_chain[21593:21592]), .config_rst(config_rst)); 
buffer_wire buffer_11437 (.in(n11437), .out(n11437_0));
mux13 mux_6272 (.in({n14041_0, n14021_0, n14014_0, n13985_0/**/, n13978_0, n13971_0, n13964_0, n13936_1, n11350_1, n7027, n7019, n6931, n6919}), .out(n11438), .config_in(config_chain[21599:21594]), .config_rst(config_rst)); 
buffer_wire buffer_11438 (.in(n11438), .out(n11438_0));
mux3 mux_6273 (.in({n14769_0, n14768_0/**/, n8979}), .out(n11439), .config_in(config_chain[21601:21600]), .config_rst(config_rst)); 
buffer_wire buffer_11439 (.in(n11439), .out(n11439_0));
mux13 mux_6274 (.in({n14043_0, n14007_0/**/, n14000_0, n13993_0, n13986_0, n13972_0, n13957_0, n13912_1, n11308_1, n7027, n7019, n6931, n6923}), .out(n11440), .config_in(config_chain[21607:21602]), .config_rst(config_rst)); 
buffer_wire buffer_11440 (.in(n11440), .out(n11440_0));
mux3 mux_6275 (.in({n14771_0, n14770_0, n8983}), .out(n11441), .config_in(config_chain[21609:21608]), .config_rst(config_rst)); 
buffer_wire buffer_11441 (.in(n11441), .out(n11441_0));
mux15 mux_6276 (.in({n14311_0, n14275_0, n14268_0, n14266_0, n14259_0, n14252_0, n14238_0, n14223_0, n14220_1, n11354_1/**/, n8005, n7997, n7909, n7901, n7893}), .out(n11442), .config_in(config_chain[21615:21610]), .config_rst(config_rst)); 
buffer_wire buffer_11442 (.in(n11442), .out(n11442_0));
mux4 mux_6277 (.in({n14773_0, n14772_0, n8987, n8871}), .out(n11443), .config_in(config_chain[21617:21616]), .config_rst(config_rst)); 
buffer_wire buffer_11443 (.in(n11443), .out(n11443_0));
mux15 mux_6278 (.in({n14291_0, n14288_0, n14283_0, n14276_0, n14260_0, n14245_0, n14231_0, n14224_0, n14218_1, n11356_1, n8009, n7997, n7909, n7901, n7893}), .out(n11444), .config_in(config_chain[21623:21618]), .config_rst(config_rst)); 
buffer_wire buffer_11444 (.in(n11444), .out(n11444_0));
mux3 mux_6279 (.in({n14775_0, n14774_0/**/, n8875}), .out(n11445), .config_in(config_chain[21625:21624]), .config_rst(config_rst)); 
buffer_wire buffer_11445 (.in(n11445), .out(n11445_0));
mux15 mux_6280 (.in({n14293_0, n14284_0, n14269_0, n14267_0, n14253_0, n14246_0, n14239_0, n14232_0, n14216_1, n11358_1, n8009, n8001, n7909, n7901, n7893/**/}), .out(n11446), .config_in(config_chain[21631:21626]), .config_rst(config_rst)); 
buffer_wire buffer_11446 (.in(n11446), .out(n11446_0));
mux3 mux_6281 (.in({n14777_0, n14776_0, n8875}), .out(n11447), .config_in(config_chain[21633:21632]), .config_rst(config_rst)); 
buffer_wire buffer_11447 (.in(n11447), .out(n11447_0));
mux15 mux_6282 (.in({n14295_0, n14289_0, n14277_0, n14270_0, n14261_0, n14254_0, n14240_0, n14225_0, n14214_1/**/, n11360_1, n8009, n8001, n7993, n7901, n7893}), .out(n11448), .config_in(config_chain[21639:21634]), .config_rst(config_rst)); 
buffer_wire buffer_11448 (.in(n11448), .out(n11448_0));
mux3 mux_6283 (.in({n14779_0, n14778_0, n8879}), .out(n11449), .config_in(config_chain[21641:21640]), .config_rst(config_rst)); 
buffer_wire buffer_11449 (.in(n11449), .out(n11449_0));
mux14 mux_6284 (.in({n14297_0, n14285_0, n14278_0, n14262_0, n14247_0, n14233_0, n14226_0, n14212_1, n11362_1/**/, n8009, n8001, n7993, n7905, n7893}), .out(n11450), .config_in(config_chain[21647:21642]), .config_rst(config_rst)); 
buffer_wire buffer_11450 (.in(n11450), .out(n11450_0));
mux3 mux_6285 (.in({n14781_0, n14780_0/**/, n8883}), .out(n11451), .config_in(config_chain[21649:21648]), .config_rst(config_rst)); 
buffer_wire buffer_11451 (.in(n11451), .out(n11451_0));
mux14 mux_6286 (.in({n14299_0, n14286_0, n14271_0/**/, n14255_0, n14248_0, n14241_0, n14234_0, n14210_1, n11364_1, n8009, n8001, n7993, n7905, n7897}), .out(n11452), .config_in(config_chain[21655:21650]), .config_rst(config_rst)); 
buffer_wire buffer_11452 (.in(n11452), .out(n11452_0));
mux3 mux_6287 (.in({n14783_0, n14782_0, n8887}), .out(n11453), .config_in(config_chain[21657:21656]), .config_rst(config_rst)); 
buffer_wire buffer_11453 (.in(n11453), .out(n11453_0));
mux13 mux_6288 (.in({n14301_0, n14279_0, n14272_0, n14263_0, n14256_0, n14242_0, n14227_0, n14208_1, n11366_1, n8001/**/, n7993, n7905, n7897}), .out(n11454), .config_in(config_chain[21663:21658]), .config_rst(config_rst)); 
buffer_wire buffer_11454 (.in(n11454), .out(n11454_0));
mux3 mux_6289 (.in({n14785_0, n14784_0/**/, n8971}), .out(n11455), .config_in(config_chain[21665:21664]), .config_rst(config_rst)); 
buffer_wire buffer_11455 (.in(n11455), .out(n11455_0));
mux13 mux_6290 (.in({n14303_0, n14287_0, n14280_0, n14264_0, n14249_0, n14235_0, n14228_0, n14206_1, n11368_1, n8005, n7993, n7905, n7897}), .out(n11456), .config_in(config_chain[21671:21666]), .config_rst(config_rst)); 
buffer_wire buffer_11456 (.in(n11456), .out(n11456_0));
mux3 mux_6291 (.in({n14787_0, n14786_0, n8971}), .out(n11457), .config_in(config_chain[21673:21672]), .config_rst(config_rst)); 
buffer_wire buffer_11457 (.in(n11457), .out(n11457_0));
mux13 mux_6292 (.in({n14305_0, n14273_0, n14257_0, n14250_0, n14243_0, n14236_0, n14204_1, n14200_1, n11370_1, n8005, n7997, n7905, n7897}), .out(n11458), .config_in(config_chain[21679:21674]), .config_rst(config_rst)); 
buffer_wire buffer_11458 (.in(n11458), .out(n11458_0));
mux3 mux_6293 (.in({n14789_0, n14788_0/**/, n8975}), .out(n11459), .config_in(config_chain[21681:21680]), .config_rst(config_rst)); 
buffer_wire buffer_11459 (.in(n11459), .out(n11459_0));
mux13 mux_6294 (.in({n14307_0, n14281_0/**/, n14274_0, n14265_0, n14258_0, n14229_0, n14222_1, n14202_1, n11372_1, n8005, n7997, n7909, n7897}), .out(n11460), .config_in(config_chain[21687:21682]), .config_rst(config_rst)); 
buffer_wire buffer_11460 (.in(n11460), .out(n11460_0));
mux3 mux_6295 (.in({n14791_0, n14790_0, n8979/**/}), .out(n11461), .config_in(config_chain[21689:21688]), .config_rst(config_rst)); 
buffer_wire buffer_11461 (.in(n11461), .out(n11461_0));
mux13 mux_6296 (.in({n14309_0/**/, n14282_0, n14251_0, n14244_0, n14237_0, n14230_0, n14201_0, n14178_1, n11310_2, n8005, n7997, n7909, n7901}), .out(n11462), .config_in(config_chain[21695:21690]), .config_rst(config_rst)); 
buffer_wire buffer_11462 (.in(n11462), .out(n11462_0));
mux3 mux_6297 (.in({n14793_0, n14792_0/**/, n8987}), .out(n11463), .config_in(config_chain[21697:21696]), .config_rst(config_rst)); 
buffer_wire buffer_11463 (.in(n11463), .out(n11463_0));
mux16 mux_6298 (.in({n14573_0, n14538_0, n14535_0, n14531_0, n14527_0, n14510_0, n14500_0, n14497_0, n14482_1, n14432_1, n11376_1/**/, n8983, n8975, n8887, n8879, n8871}), .out(n11464), .config_in(config_chain[21703:21698]), .config_rst(config_rst)); 
buffer_wire buffer_11464 (.in(n11464), .out(n11464_0));
mux4 mux_6299 (.in({n14795_0, n14794_0, n8987, n8871}), .out(n11465), .config_in(config_chain[21705:21704]), .config_rst(config_rst)); 
buffer_wire buffer_11465 (.in(n11465), .out(n11465_0));
mux16 mux_6300 (.in({n14555_0, n14553_0, n14549_0, n14532_0, n14524_0, n14521_0, n14494_0, n14491_0, n14480_1, n14464_1, n11378_1, n8983, n8975, n8887, n8879/**/, n8871}), .out(n11466), .config_in(config_chain[21711:21706]), .config_rst(config_rst)); 
buffer_wire buffer_11466 (.in(n11466), .out(n11466_0));
mux3 mux_6301 (.in({n14797_0/**/, n14796_0, n8875}), .out(n11467), .config_in(config_chain[21713:21712]), .config_rst(config_rst)); 
buffer_wire buffer_11467 (.in(n11467), .out(n11467_0));
mux15 mux_6302 (.in({n14557_0, n14546_0, n14543_0, n14518_0, n14515_0, n14505_0, n14488_0, n14486_1, n14478_1, n11380_1, n8983, n8975, n8887, n8879, n8871}), .out(n11468), .config_in(config_chain[21719:21714]), .config_rst(config_rst)); 
buffer_wire buffer_11468 (.in(n11468), .out(n11468_0));
mux3 mux_6303 (.in({n14799_0, n14798_0, n8879}), .out(n11469), .config_in(config_chain[21721:21720]), .config_rst(config_rst)); 
buffer_wire buffer_11469 (.in(n11469), .out(n11469_0));
mux15 mux_6304 (.in({n14559_0, n14540_0, n14537_0, n14529_0, n14512_0/**/, n14508_0, n14502_0, n14499_0, n14476_1, n11382_1, n8983, n8975, n8887, n8879, n8871}), .out(n11470), .config_in(config_chain[21727:21722]), .config_rst(config_rst)); 
buffer_wire buffer_11470 (.in(n11470), .out(n11470_0));
mux3 mux_6305 (.in({n14801_0, n14800_0, n8879}), .out(n11471), .config_in(config_chain[21729:21728]), .config_rst(config_rst)); 
buffer_wire buffer_11471 (.in(n11471), .out(n11471_0));
mux15 mux_6306 (.in({n14561_0, n14551_0, n14534_0, n14530_0, n14526_0, n14523_0/**/, n14496_0, n14493_0, n14474_1, n11384_1, n8983, n8975, n8887, n8879, n8871}), .out(n11472), .config_in(config_chain[21735:21730]), .config_rst(config_rst)); 
buffer_wire buffer_11472 (.in(n11472), .out(n11472_0));
mux3 mux_6307 (.in({n14803_0, n14802_0, n8883}), .out(n11473), .config_in(config_chain[21737:21736]), .config_rst(config_rst)); 
buffer_wire buffer_11473 (.in(n11473), .out(n11473_0));
mux15 mux_6308 (.in({n14563_0, n14552_0, n14548_0/**/, n14545_0, n14520_0, n14517_0, n14507_0, n14490_0, n14472_1, n11386_1, n8987, n8979, n8971, n8883, n8875}), .out(n11474), .config_in(config_chain[21743:21738]), .config_rst(config_rst)); 
buffer_wire buffer_11474 (.in(n11474), .out(n11474_0));
mux3 mux_6309 (.in({n14805_0, n14804_0, n8887/**/}), .out(n11475), .config_in(config_chain[21745:21744]), .config_rst(config_rst)); 
buffer_wire buffer_11475 (.in(n11475), .out(n11475_0));
mux15 mux_6310 (.in({n14565_0, n14542_0, n14539_0, n14514_0, n14511_0, n14504_0, n14501_0, n14470_1, n14433_0, n11388_1, n8987/**/, n8979, n8971, n8883, n8875}), .out(n11476), .config_in(config_chain[21751:21746]), .config_rst(config_rst)); 
buffer_wire buffer_11476 (.in(n11476), .out(n11476_0));
mux3 mux_6311 (.in({n14807_0, n14806_0, n8971}), .out(n11477), .config_in(config_chain[21753:21752]), .config_rst(config_rst)); 
buffer_wire buffer_11477 (.in(n11477), .out(n11477_0));
mux15 mux_6312 (.in({n14567_0, n14536_0, n14533_0, n14528_0, n14525_0, n14498_0, n14495_0, n14468_1, n14465_0, n11390_1, n8987, n8979, n8971, n8883/**/, n8875}), .out(n11478), .config_in(config_chain[21759:21754]), .config_rst(config_rst)); 
buffer_wire buffer_11478 (.in(n11478), .out(n11478_0));
mux3 mux_6313 (.in({n14809_0, n14808_0, n8975}), .out(n11479), .config_in(config_chain[21761:21760]), .config_rst(config_rst)); 
buffer_wire buffer_11479 (.in(n11479), .out(n11479_0));
mux15 mux_6314 (.in({n14569_0, n14550_0, n14547_0, n14522_0/**/, n14519_0, n14492_0, n14489_0, n14487_0, n14466_1, n11392_1, n8987, n8979, n8971, n8883, n8875}), .out(n11480), .config_in(config_chain[21767:21762]), .config_rst(config_rst)); 
buffer_wire buffer_11480 (.in(n11480), .out(n11480_0));
mux3 mux_6315 (.in({n14811_0, n14810_0, n8975}), .out(n11481), .config_in(config_chain[21769:21768]), .config_rst(config_rst)); 
buffer_wire buffer_11481 (.in(n11481), .out(n11481_0));
mux15 mux_6316 (.in({n14571_0, n14544_0, n14541_0/**/, n14516_0, n14513_0, n14509_0, n14506_0, n14503_0, n14484_1, n11394_1, n8987, n8979, n8971, n8883, n8875}), .out(n11482), .config_in(config_chain[21775:21770]), .config_rst(config_rst)); 
buffer_wire buffer_11482 (.in(n11482), .out(n11482_0));
mux3 mux_6317 (.in({n14813_0, n14812_0, n8979}), .out(n11483), .config_in(config_chain[21777:21776]), .config_rst(config_rst)); 
buffer_wire buffer_11483 (.in(n11483), .out(n11483_0));
mux4 mux_6318 (.in({n12423_0, n12422_0, n1261, n1145}), .out(n11484), .config_in(config_chain[21779:21778]), .config_rst(config_rst)); 
buffer_wire buffer_11484 (.in(n11484), .out(n11484_0));
mux15 mux_6319 (.in({n12737_0, n12728_0, n12723_0, n12711_0, n12682_0, n12677_0, n12613_0, n12608_2, n12604_2, n11577_1, n1257, n1249, n1161, n1153, n1145}), .out(n11485), .config_in(config_chain[21785:21780]), .config_rst(config_rst)); 
buffer_wire buffer_11485 (.in(n11485), .out(n11485_0));
mux4 mux_6320 (.in({n12443_0, n12442_0, n1261, n1145}), .out(n11486), .config_in(config_chain[21787:21786]), .config_rst(config_rst)); 
buffer_wire buffer_11486 (.in(n11486), .out(n11486_0));
mux15 mux_6321 (.in({n12995_0, n12978_0, n12973_0, n12964_0, n12959_0, n12947_0, n12869_0, n12864_2, n12862_2, n11599_1/**/, n2235, n2227, n2139, n2131, n2123}), .out(n11487), .config_in(config_chain[21793:21788]), .config_rst(config_rst)); 
buffer_wire buffer_11487 (.in(n11487), .out(n11487_0));
mux4 mux_6322 (.in({n12463_0, n12462_0, n1261, n1145}), .out(n11488), .config_in(config_chain[21795:21794]), .config_rst(config_rst)); 
buffer_wire buffer_11488 (.in(n11488), .out(n11488_0));
mux15 mux_6323 (.in({n13255_0, n13252_0, n13247_0, n13216_0, n13211_0, n13202_0, n13197_0, n13127_0, n13122_2, n11621_1/**/, n3213, n3205, n3117, n3109, n3101}), .out(n11489), .config_in(config_chain[21801:21796]), .config_rst(config_rst)); 
buffer_wire buffer_11489 (.in(n11489), .out(n11489_0));
mux4 mux_6324 (.in({n12483_0, n12402_1, n1261, n1145}), .out(n11490), .config_in(config_chain[21803:21802]), .config_rst(config_rst)); 
buffer_wire buffer_11490 (.in(n11490), .out(n11490_0));
mux15 mux_6325 (.in({n13517_0, n13506_0, n13501_0, n13492_0, n13487_0, n13456_0, n13451_0, n13387_0, n13384_2, n11643_1/**/, n4191, n4183, n4095, n4087, n4079}), .out(n11491), .config_in(config_chain[21809:21804]), .config_rst(config_rst)); 
buffer_wire buffer_11491 (.in(n11491), .out(n11491_0));
mux3 mux_6326 (.in({n12425_0, n12424_0, n1145}), .out(n11492), .config_in(config_chain[21811:21810]), .config_rst(config_rst)); 
buffer_wire buffer_11492 (.in(n11492), .out(n11492_0));
mux15 mux_6327 (.in({n12757_0, n12731_0, n12702_0, n12697_0, n12690_0, n12685_0, n12656_1, n12615_0, n12610_2, n11579_1, n1261, n1249, n1161, n1153, n1145}), .out(n11493), .config_in(config_chain[21817:21812]), .config_rst(config_rst)); 
buffer_wire buffer_11493 (.in(n11493), .out(n11493_0));
mux3 mux_6328 (.in({n12445_0, n12444_0, n1149}), .out(n11494), .config_in(config_chain[21819:21818]), .config_rst(config_rst)); 
buffer_wire buffer_11494 (.in(n11494), .out(n11494_0));
mux15 mux_6329 (.in({n13015_0, n12986_0, n12981_0, n12967_0, n12938_0, n12933_0, n12912_1, n12871_0, n12866_2, n11601_1, n2239, n2227, n2139, n2131, n2123}), .out(n11495), .config_in(config_chain[21825:21820]), .config_rst(config_rst)); 
buffer_wire buffer_11495 (.in(n11495), .out(n11495_0));
mux3 mux_6330 (.in({n12465_0, n12464_0, n1149}), .out(n11496), .config_in(config_chain[21827:21826]), .config_rst(config_rst)); 
buffer_wire buffer_11496 (.in(n11496), .out(n11496_0));
mux15 mux_6331 (.in({n13275_0, n13238_0, n13233_0, n13224_0, n13219_0/**/, n13205_0, n13170_1, n13129_0, n13124_2, n11623_1, n3217, n3205, n3117, n3109, n3101}), .out(n11497), .config_in(config_chain[21833:21828]), .config_rst(config_rst)); 
buffer_wire buffer_11497 (.in(n11497), .out(n11497_0));
mux3 mux_6332 (.in({n12485_0, n12404_1, n1149}), .out(n11498), .config_in(config_chain[21835:21834]), .config_rst(config_rst)); 
buffer_wire buffer_11498 (.in(n11498), .out(n11498_0));
mux15 mux_6333 (.in({n13537_0, n13514_0, n13509_0, n13478_0, n13473_0, n13464_0, n13459_0, n13430_1/**/, n13389_0, n11645_1, n4195, n4183, n4095, n4087, n4079}), .out(n11499), .config_in(config_chain[21841:21836]), .config_rst(config_rst)); 
buffer_wire buffer_11499 (.in(n11499), .out(n11499_0));
mux3 mux_6334 (.in({n12427_0, n12426_0, n1149}), .out(n11500), .config_in(config_chain[21843:21842]), .config_rst(config_rst)); 
buffer_wire buffer_11500 (.in(n11500), .out(n11500_0));
mux15 mux_6335 (.in({n12755_0, n12722_0, n12717_0, n12710_0, n12705_0, n12693_0, n12676_0/**/, n12658_1, n12612_2, n11581_1, n1261, n1253, n1161, n1153, n1145}), .out(n11501), .config_in(config_chain[21849:21844]), .config_rst(config_rst)); 
buffer_wire buffer_11501 (.in(n11501), .out(n11501_0));
mux3 mux_6336 (.in({n12447_0, n12446_0, n1149}), .out(n11502), .config_in(config_chain[21851:21850]), .config_rst(config_rst)); 
buffer_wire buffer_11502 (.in(n11502), .out(n11502_0));
mux15 mux_6337 (.in({n13013_0, n12989_0, n12972_0, n12958_0, n12953_0, n12946_0, n12941_0, n12914_1, n12868_2, n11603_1, n2239, n2231, n2139/**/, n2131, n2123}), .out(n11503), .config_in(config_chain[21857:21852]), .config_rst(config_rst)); 
buffer_wire buffer_11503 (.in(n11503), .out(n11503_0));
mux3 mux_6338 (.in({n12467_0, n12466_0/**/, n1153}), .out(n11504), .config_in(config_chain[21859:21858]), .config_rst(config_rst)); 
buffer_wire buffer_11504 (.in(n11504), .out(n11504_0));
mux15 mux_6339 (.in({n13273_0, n13246_0, n13241_0, n13227_0, n13210_0, n13196_0, n13191_0, n13172_1, n13126_2, n11625_1, n3217, n3209, n3117/**/, n3109, n3101}), .out(n11505), .config_in(config_chain[21865:21860]), .config_rst(config_rst)); 
buffer_wire buffer_11505 (.in(n11505), .out(n11505_0));
mux3 mux_6340 (.in({n12487_0, n12406_1/**/, n1153}), .out(n11506), .config_in(config_chain[21867:21866]), .config_rst(config_rst)); 
buffer_wire buffer_11506 (.in(n11506), .out(n11506_0));
mux15 mux_6341 (.in({n13535_0, n13500_0, n13495_0, n13486_0, n13481_0, n13467_0/**/, n13450_0, n13432_1, n13386_2, n11647_1, n4195, n4187, n4095, n4087, n4079}), .out(n11507), .config_in(config_chain[21873:21868]), .config_rst(config_rst)); 
buffer_wire buffer_11507 (.in(n11507), .out(n11507_0));
mux3 mux_6342 (.in({n12429_0, n12428_0/**/, n1153}), .out(n11508), .config_in(config_chain[21875:21874]), .config_rst(config_rst)); 
buffer_wire buffer_11508 (.in(n11508), .out(n11508_0));
mux15 mux_6343 (.in({n12753_0, n12730_0, n12725_0, n12713_0, n12696_0, n12684_0, n12679_0, n12660_1, n12614_2, n11583_1/**/, n1261, n1253, n1245, n1153, n1145}), .out(n11509), .config_in(config_chain[21881:21876]), .config_rst(config_rst)); 
buffer_wire buffer_11509 (.in(n11509), .out(n11509_0));
mux3 mux_6344 (.in({n12449_0, n12448_0, n1153}), .out(n11510), .config_in(config_chain[21883:21882]), .config_rst(config_rst)); 
buffer_wire buffer_11510 (.in(n11510), .out(n11510_0));
mux15 mux_6345 (.in({n13011_0, n12980_0/**/, n12975_0, n12966_0, n12961_0, n12949_0, n12932_0, n12916_1, n12870_2, n11605_1, n2239, n2231, n2223, n2131, n2123}), .out(n11511), .config_in(config_chain[21889:21884]), .config_rst(config_rst)); 
buffer_wire buffer_11511 (.in(n11511), .out(n11511_0));
mux3 mux_6346 (.in({n12469_0, n12468_0, n1153}), .out(n11512), .config_in(config_chain[21891:21890]), .config_rst(config_rst)); 
buffer_wire buffer_11512 (.in(n11512), .out(n11512_0));
mux15 mux_6347 (.in({n13271_0, n13249_0, n13232_0/**/, n13218_0, n13213_0, n13204_0, n13199_0, n13174_1, n13128_2, n11627_1, n3217, n3209, n3201, n3109, n3101}), .out(n11513), .config_in(config_chain[21897:21892]), .config_rst(config_rst)); 
buffer_wire buffer_11513 (.in(n11513), .out(n11513_0));
mux3 mux_6348 (.in({n12489_0, n12408_1, n1157}), .out(n11514), .config_in(config_chain[21899:21898]), .config_rst(config_rst)); 
buffer_wire buffer_11514 (.in(n11514), .out(n11514_0));
mux15 mux_6349 (.in({n13533_0, n13508_0, n13503_0, n13489_0, n13472_0, n13458_0, n13453_0, n13434_1, n13388_2, n11649_1, n4195, n4187, n4179, n4087, n4079}), .out(n11515), .config_in(config_chain[21905:21900]), .config_rst(config_rst)); 
buffer_wire buffer_11515 (.in(n11515), .out(n11515_0));
mux3 mux_6350 (.in({n12431_0, n12430_0, n1157}), .out(n11516), .config_in(config_chain[21907:21906]), .config_rst(config_rst)); 
buffer_wire buffer_11516 (.in(n11516), .out(n11516_0));
mux14 mux_6351 (.in({n12751_0, n12733_0, n12716_0, n12704_0, n12699_0, n12692_0, n12687_0, n12662_1, n11585_1, n1261, n1253, n1245, n1157, n1145}), .out(n11517), .config_in(config_chain[21913:21908]), .config_rst(config_rst)); 
buffer_wire buffer_11517 (.in(n11517), .out(n11517_0));
mux3 mux_6352 (.in({n12451_0/**/, n12450_0, n1157}), .out(n11518), .config_in(config_chain[21915:21914]), .config_rst(config_rst)); 
buffer_wire buffer_11518 (.in(n11518), .out(n11518_0));
mux14 mux_6353 (.in({n13009_0, n12988_0, n12983_0, n12969_0, n12952_0, n12940_0, n12935_0, n12918_1, n11607_1, n2239, n2231, n2223, n2135, n2123}), .out(n11519), .config_in(config_chain[21921:21916]), .config_rst(config_rst)); 
buffer_wire buffer_11519 (.in(n11519), .out(n11519_0));
mux3 mux_6354 (.in({n12471_0, n12470_0/**/, n1157}), .out(n11520), .config_in(config_chain[21923:21922]), .config_rst(config_rst)); 
buffer_wire buffer_11520 (.in(n11520), .out(n11520_0));
mux14 mux_6355 (.in({n13269_0, n13240_0, n13235_0, n13226_0, n13221_0, n13207_0, n13190_0, n13176_1, n11629_1, n3217, n3209, n3201, n3113/**/, n3101}), .out(n11521), .config_in(config_chain[21929:21924]), .config_rst(config_rst)); 
buffer_wire buffer_11521 (.in(n11521), .out(n11521_0));
mux3 mux_6356 (.in({n12491_0, n12410_1, n1157}), .out(n11522), .config_in(config_chain[21931:21930]), .config_rst(config_rst)); 
buffer_wire buffer_11522 (.in(n11522), .out(n11522_0));
mux14 mux_6357 (.in({n13531_0, n13511_0, n13494_0, n13480_0, n13475_0, n13466_0/**/, n13461_0, n13436_1, n11651_1, n4195, n4187, n4179, n4091, n4079}), .out(n11523), .config_in(config_chain[21937:21932]), .config_rst(config_rst)); 
buffer_wire buffer_11523 (.in(n11523), .out(n11523_0));
mux3 mux_6358 (.in({n12433_0, n12432_0/**/, n1161}), .out(n11524), .config_in(config_chain[21939:21938]), .config_rst(config_rst)); 
buffer_wire buffer_11524 (.in(n11524), .out(n11524_0));
mux14 mux_6359 (.in({n12749_0/**/, n12724_0, n12719_0, n12712_0, n12707_0, n12695_0, n12678_0, n12664_1, n11587_1, n1261, n1253, n1245, n1157, n1149}), .out(n11525), .config_in(config_chain[21945:21940]), .config_rst(config_rst)); 
buffer_wire buffer_11525 (.in(n11525), .out(n11525_0));
mux3 mux_6360 (.in({n12453_0, n12452_0, n1161/**/}), .out(n11526), .config_in(config_chain[21947:21946]), .config_rst(config_rst)); 
buffer_wire buffer_11526 (.in(n11526), .out(n11526_0));
mux14 mux_6361 (.in({n13007_0, n12991_0, n12974_0, n12960_0, n12955_0, n12948_0, n12943_0, n12920_1/**/, n11609_1, n2239, n2231, n2223, n2135, n2127}), .out(n11527), .config_in(config_chain[21953:21948]), .config_rst(config_rst)); 
buffer_wire buffer_11527 (.in(n11527), .out(n11527_0));
mux3 mux_6362 (.in({n12473_0, n12472_0/**/, n1161}), .out(n11528), .config_in(config_chain[21955:21954]), .config_rst(config_rst)); 
buffer_wire buffer_11528 (.in(n11528), .out(n11528_0));
mux14 mux_6363 (.in({n13267_0, n13248_0, n13243_0, n13229_0, n13212_0, n13198_0, n13193_0, n13178_1, n11631_1, n3217, n3209, n3201, n3113, n3105/**/}), .out(n11529), .config_in(config_chain[21961:21956]), .config_rst(config_rst)); 
buffer_wire buffer_11529 (.in(n11529), .out(n11529_0));
mux3 mux_6364 (.in({n12493_0, n12412_1/**/, n1161}), .out(n11530), .config_in(config_chain[21963:21962]), .config_rst(config_rst)); 
buffer_wire buffer_11530 (.in(n11530), .out(n11530_0));
mux14 mux_6365 (.in({n13529_0, n13502_0, n13497_0, n13488_0, n13483_0, n13469_0, n13452_0, n13438_1/**/, n11653_1, n4195, n4187, n4179, n4091, n4083}), .out(n11531), .config_in(config_chain[21969:21964]), .config_rst(config_rst)); 
buffer_wire buffer_11531 (.in(n11531), .out(n11531_0));
mux3 mux_6366 (.in({n12435_0, n12434_0/**/, n1161}), .out(n11532), .config_in(config_chain[21971:21970]), .config_rst(config_rst)); 
buffer_wire buffer_11532 (.in(n11532), .out(n11532_0));
mux13 mux_6367 (.in({n12747_0, n12732_0, n12727_0, n12715_0, n12698_0, n12686_0, n12681_0, n12666_1, n11589_1, n1253, n1245, n1157, n1149}), .out(n11533), .config_in(config_chain[21977:21972]), .config_rst(config_rst)); 
buffer_wire buffer_11533 (.in(n11533), .out(n11533_0));
mux3 mux_6368 (.in({n12455_0, n12454_0, n1245}), .out(n11534), .config_in(config_chain[21979:21978]), .config_rst(config_rst)); 
buffer_wire buffer_11534 (.in(n11534), .out(n11534_0));
mux13 mux_6369 (.in({n13005_0, n12982_0, n12977_0, n12968_0, n12963_0, n12951_0, n12934_0, n12922_1/**/, n11611_1, n2231, n2223, n2135, n2127}), .out(n11535), .config_in(config_chain[21985:21980]), .config_rst(config_rst)); 
buffer_wire buffer_11535 (.in(n11535), .out(n11535_0));
mux3 mux_6370 (.in({n12475_0, n12474_0, n1245}), .out(n11536), .config_in(config_chain[21987:21986]), .config_rst(config_rst)); 
buffer_wire buffer_11536 (.in(n11536), .out(n11536_0));
mux13 mux_6371 (.in({n13265_0, n13251_0, n13234_0, n13220_0, n13215_0, n13206_0, n13201_0, n13180_1, n11633_1, n3209, n3201, n3113, n3105/**/}), .out(n11537), .config_in(config_chain[21993:21988]), .config_rst(config_rst)); 
buffer_wire buffer_11537 (.in(n11537), .out(n11537_0));
mux3 mux_6372 (.in({n12495_0, n12414_1/**/, n1245}), .out(n11538), .config_in(config_chain[21995:21994]), .config_rst(config_rst)); 
buffer_wire buffer_11538 (.in(n11538), .out(n11538_0));
mux13 mux_6373 (.in({n13527_0, n13510_0, n13505_0, n13491_0, n13474_0/**/, n13460_0, n13455_0, n13440_1, n11655_1, n4187, n4179, n4091, n4083}), .out(n11539), .config_in(config_chain[22001:21996]), .config_rst(config_rst)); 
buffer_wire buffer_11539 (.in(n11539), .out(n11539_0));
mux3 mux_6374 (.in({n12437_0, n12436_0, n1245/**/}), .out(n11540), .config_in(config_chain[22003:22002]), .config_rst(config_rst)); 
buffer_wire buffer_11540 (.in(n11540), .out(n11540_0));
mux13 mux_6375 (.in({n12745_0, n12735_0, n12718_0, n12706_0, n12701_0, n12694_0, n12689_0, n12668_1, n11591_1, n1257, n1245, n1157, n1149}), .out(n11541), .config_in(config_chain[22009:22004]), .config_rst(config_rst)); 
buffer_wire buffer_11541 (.in(n11541), .out(n11541_0));
mux3 mux_6376 (.in({n12457_0, n12456_0, n1245}), .out(n11542), .config_in(config_chain[22011:22010]), .config_rst(config_rst)); 
buffer_wire buffer_11542 (.in(n11542), .out(n11542_0));
mux13 mux_6377 (.in({n13003_0, n12990_0, n12985_0, n12971_0, n12954_0, n12942_0/**/, n12937_0, n12924_1, n11613_1, n2235, n2223, n2135, n2127}), .out(n11543), .config_in(config_chain[22017:22012]), .config_rst(config_rst)); 
buffer_wire buffer_11543 (.in(n11543), .out(n11543_0));
mux3 mux_6378 (.in({n12477_0, n12476_0, n1249}), .out(n11544), .config_in(config_chain[22019:22018]), .config_rst(config_rst)); 
buffer_wire buffer_11544 (.in(n11544), .out(n11544_0));
mux13 mux_6379 (.in({n13263_0, n13242_0, n13237_0/**/, n13228_0, n13223_0, n13209_0, n13192_0, n13182_1, n11635_1, n3213, n3201, n3113, n3105}), .out(n11545), .config_in(config_chain[22025:22020]), .config_rst(config_rst)); 
buffer_wire buffer_11545 (.in(n11545), .out(n11545_0));
mux3 mux_6380 (.in({n12497_0, n12416_1, n1249}), .out(n11546), .config_in(config_chain[22027:22026]), .config_rst(config_rst)); 
buffer_wire buffer_11546 (.in(n11546), .out(n11546_0));
mux13 mux_6381 (.in({n13525_0, n13513_0, n13496_0, n13482_0, n13477_0, n13468_0, n13463_0, n13442_1/**/, n11657_1, n4191, n4179, n4091, n4083}), .out(n11547), .config_in(config_chain[22033:22028]), .config_rst(config_rst)); 
buffer_wire buffer_11547 (.in(n11547), .out(n11547_0));
mux3 mux_6382 (.in({n12439_0, n12438_0/**/, n1249}), .out(n11548), .config_in(config_chain[22035:22034]), .config_rst(config_rst)); 
buffer_wire buffer_11548 (.in(n11548), .out(n11548_0));
mux13 mux_6383 (.in({n12743_0/**/, n12726_0, n12721_0, n12714_0, n12709_0, n12680_0, n12670_1, n12607_0, n11593_1, n1257, n1249, n1157, n1149}), .out(n11549), .config_in(config_chain[22041:22036]), .config_rst(config_rst)); 
buffer_wire buffer_11549 (.in(n11549), .out(n11549_0));
mux3 mux_6384 (.in({n12459_0, n12458_0, n1249}), .out(n11550), .config_in(config_chain[22043:22042]), .config_rst(config_rst)); 
buffer_wire buffer_11550 (.in(n11550), .out(n11550_0));
mux13 mux_6385 (.in({n13001_0, n12993_0, n12976_0, n12962_0, n12957_0, n12950_0, n12945_0, n12926_1, n11615_1, n2235, n2227, n2135, n2127}), .out(n11551), .config_in(config_chain[22049:22044]), .config_rst(config_rst)); 
buffer_wire buffer_11551 (.in(n11551), .out(n11551_0));
mux3 mux_6386 (.in({n12479_0, n12478_0, n1249}), .out(n11552), .config_in(config_chain[22051:22050]), .config_rst(config_rst)); 
buffer_wire buffer_11552 (.in(n11552), .out(n11552_0));
mux13 mux_6387 (.in({n13261_0, n13250_0, n13245_0, n13231_0, n13214_0, n13200_0, n13195_0, n13184_1, n11637_1, n3213, n3205, n3113, n3105}), .out(n11553), .config_in(config_chain[22057:22052]), .config_rst(config_rst)); 
buffer_wire buffer_11553 (.in(n11553), .out(n11553_0));
mux3 mux_6388 (.in({n12499_0, n12418_1/**/, n1253}), .out(n11554), .config_in(config_chain[22059:22058]), .config_rst(config_rst)); 
buffer_wire buffer_11554 (.in(n11554), .out(n11554_0));
mux13 mux_6389 (.in({n13523_0, n13504_0, n13499_0, n13490_0, n13485_0, n13471_0, n13454_0, n13444_1, n11659_1, n4191, n4183, n4091/**/, n4083}), .out(n11555), .config_in(config_chain[22065:22060]), .config_rst(config_rst)); 
buffer_wire buffer_11555 (.in(n11555), .out(n11555_0));
mux3 mux_6390 (.in({n12441_0, n12440_0/**/, n1253}), .out(n11556), .config_in(config_chain[22067:22066]), .config_rst(config_rst)); 
buffer_wire buffer_11556 (.in(n11556), .out(n11556_0));
mux13 mux_6391 (.in({n12741_0, n12734_0, n12729_0, n12700_0, n12688_0, n12683_0, n12672_1/**/, n12609_0, n11595_1, n1257, n1249, n1161, n1149}), .out(n11557), .config_in(config_chain[22073:22068]), .config_rst(config_rst)); 
buffer_wire buffer_11557 (.in(n11557), .out(n11557_0));
mux3 mux_6392 (.in({n12461_0, n12460_0, n1253/**/}), .out(n11558), .config_in(config_chain[22075:22074]), .config_rst(config_rst)); 
buffer_wire buffer_11558 (.in(n11558), .out(n11558_0));
mux13 mux_6393 (.in({n12999_0, n12984_0, n12979_0, n12970_0, n12965_0/**/, n12936_0, n12928_1, n12865_0, n11617_1, n2235, n2227, n2139, n2127}), .out(n11559), .config_in(config_chain[22081:22076]), .config_rst(config_rst)); 
buffer_wire buffer_11559 (.in(n11559), .out(n11559_0));
mux3 mux_6394 (.in({n12481_0, n12480_0/**/, n1253}), .out(n11560), .config_in(config_chain[22083:22082]), .config_rst(config_rst)); 
buffer_wire buffer_11560 (.in(n11560), .out(n11560_0));
mux13 mux_6395 (.in({n13259_0, n13253_0, n13236_0, n13222_0/**/, n13217_0, n13208_0, n13203_0, n13186_1, n11639_1, n3213, n3205, n3117, n3105}), .out(n11561), .config_in(config_chain[22089:22084]), .config_rst(config_rst)); 
buffer_wire buffer_11561 (.in(n11561), .out(n11561_0));
mux3 mux_6396 (.in({n12501_0, n12420_1/**/, n1253}), .out(n11562), .config_in(config_chain[22091:22090]), .config_rst(config_rst)); 
buffer_wire buffer_11562 (.in(n11562), .out(n11562_0));
mux13 mux_6397 (.in({n13521_0, n13512_0, n13507_0, n13493_0, n13476_0, n13462_0, n13457_0, n13446_1, n11661_1/**/, n4191, n4183, n4095, n4083}), .out(n11563), .config_in(config_chain[22097:22092]), .config_rst(config_rst)); 
buffer_wire buffer_11563 (.in(n11563), .out(n11563_0));
mux3 mux_6398 (.in({n12351_0, n12350_2, n1257}), .out(n11564), .config_in(config_chain[22099:22098]), .config_rst(config_rst)); 
buffer_wire buffer_11564 (.in(n11564), .out(n11564_0));
mux13 mux_6399 (.in({n12739_0, n12720_0, n12708_0, n12703_0, n12691_0, n12674_1, n12611_0, n12606_2, n11597_2, n1257, n1249, n1161, n1153}), .out(n11565), .config_in(config_chain[22105:22100]), .config_rst(config_rst)); 
buffer_wire buffer_11565 (.in(n11565), .out(n11565_0));
mux3 mux_6400 (.in({n12353_0, n12352_2, n1257}), .out(n11566), .config_in(config_chain[22107:22106]), .config_rst(config_rst)); 
buffer_wire buffer_11566 (.in(n11566), .out(n11566_0));
mux13 mux_6401 (.in({n12997_0, n12992_0, n12987_0, n12956_0, n12944_0, n12939_0, n12930_1, n12867_0, n11619_2, n2235, n2227, n2139, n2131/**/}), .out(n11567), .config_in(config_chain[22113:22108]), .config_rst(config_rst)); 
buffer_wire buffer_11567 (.in(n11567), .out(n11567_0));
mux3 mux_6402 (.in({n12355_0, n12354_2, n1257}), .out(n11568), .config_in(config_chain[22115:22114]), .config_rst(config_rst)); 
buffer_wire buffer_11568 (.in(n11568), .out(n11568_0));
mux13 mux_6403 (.in({n13257_0, n13244_0, n13239_0, n13230_0, n13225_0, n13194_0, n13188_1/**/, n13125_0, n11641_1, n3213, n3205, n3117, n3109}), .out(n11569), .config_in(config_chain[22121:22116]), .config_rst(config_rst)); 
buffer_wire buffer_11569 (.in(n11569), .out(n11569_0));
mux3 mux_6404 (.in({n12357_0, n12356_2, n1257/**/}), .out(n11570), .config_in(config_chain[22123:22122]), .config_rst(config_rst)); 
buffer_wire buffer_11570 (.in(n11570), .out(n11570_0));
mux13 mux_6405 (.in({n13519_0, n13515_0, n13498_0, n13484_0, n13479_0, n13470_0, n13465_0, n13448_1, n11663_1, n4191, n4183, n4095/**/, n4087}), .out(n11571), .config_in(config_chain[22129:22124]), .config_rst(config_rst)); 
buffer_wire buffer_11571 (.in(n11571), .out(n11571_0));
mux3 mux_6406 (.in({n12359_0, n12358_2, n1257}), .out(n11572), .config_in(config_chain[22131:22130]), .config_rst(config_rst)); 
buffer_wire buffer_11572 (.in(n11572), .out(n11572_0));
mux13 mux_6407 (.in({n13783_0, n13762_0, n13757_0, n13748_0, n13743_0, n13729_0, n13712_1, n13710_1/**/, n11685_1, n5169, n5161, n5073, n5065}), .out(n11573), .config_in(config_chain[22137:22132]), .config_rst(config_rst)); 
buffer_wire buffer_11573 (.in(n11573), .out(n11573_0));
mux3 mux_6408 (.in({n12361_0, n12360_2, n1261}), .out(n11574), .config_in(config_chain[22139:22138]), .config_rst(config_rst)); 
buffer_wire buffer_11574 (.in(n11574), .out(n11574_0));
mux13 mux_6409 (.in({n14049_0, n14039_0, n14006_0, n14001_0, n13992_0, n13987_0, n13976_1, n13956_1, n11707_0/**/, n6147, n6139, n6051, n6043}), .out(n11575), .config_in(config_chain[22145:22140]), .config_rst(config_rst)); 
buffer_wire buffer_11575 (.in(n11575), .out(n11575_0));
mux15 mux_6410 (.in({n12757_0, n12729_0, n12722_0, n12710_0/**/, n12683_0, n12676_0, n12674_1, n12612_2, n12609_0, n11484_0, n2235, n2227, n2139, n2131, n2123}), .out(n11576), .config_in(config_chain[22151:22146]), .config_rst(config_rst)); 
buffer_wire buffer_11576 (.in(n11576), .out(n11576_0));
mux15 mux_6411 (.in({n13781_0/**/, n13779_0, n13770_0, n13765_0, n13751_0, n13734_0, n13720_0, n13715_0, n13648_2, n11665_1, n5169, n5161, n5073, n5065, n5057}), .out(n11577), .config_in(config_chain[22157:22152]), .config_rst(config_rst)); 
buffer_wire buffer_11577 (.in(n11577), .out(n11577_0));
mux15 mux_6412 (.in({n12737_0, n12730_0/**/, n12703_0, n12696_0, n12691_0, n12684_0, n12672_1, n12614_2, n12611_0, n11492_0, n2239, n2227, n2139, n2131, n2123}), .out(n11578), .config_in(config_chain[22163:22158]), .config_rst(config_rst)); 
buffer_wire buffer_11578 (.in(n11578), .out(n11578_0));
mux15 mux_6413 (.in({n13801_0, n13773_0, n13756_0, n13742_0, n13737_0, n13728_0, n13723_0, n13692_1, n13651_0, n11667_1, n5173/**/, n5161, n5073, n5065, n5057}), .out(n11579), .config_in(config_chain[22169:22164]), .config_rst(config_rst)); 
buffer_wire buffer_11579 (.in(n11579), .out(n11579_0));
mux15 mux_6414 (.in({n12739_0, n12723_0, n12716_0, n12711_0, n12704_0, n12692_0, n12677_0, n12670_1, n12613_0, n11500_0, n2239, n2231, n2139, n2131/**/, n2123}), .out(n11580), .config_in(config_chain[22175:22170]), .config_rst(config_rst)); 
buffer_wire buffer_11580 (.in(n11580), .out(n11580_0));
mux15 mux_6415 (.in({n13799_0, n13778_0, n13764_0, n13759_0, n13750_0, n13745_0, n13731_0, n13714_0, n13694_1, n11669_1/**/, n5173, n5165, n5073, n5065, n5057}), .out(n11581), .config_in(config_chain[22181:22176]), .config_rst(config_rst)); 
buffer_wire buffer_11581 (.in(n11581), .out(n11581_0));
mux15 mux_6416 (.in({n12741_0, n12731_0, n12724_0, n12712_0, n12697_0, n12685_0, n12678_0, n12668_1, n12615_0, n11508_0, n2239, n2231, n2223, n2131/**/, n2123}), .out(n11582), .config_in(config_chain[22187:22182]), .config_rst(config_rst)); 
buffer_wire buffer_11582 (.in(n11582), .out(n11582_0));
mux15 mux_6417 (.in({n13797_0, n13772_0, n13767_0, n13753_0, n13736_0, n13722_0/**/, n13717_0, n13696_1, n13650_2, n11671_1, n5173, n5165, n5157, n5065, n5057}), .out(n11583), .config_in(config_chain[22193:22188]), .config_rst(config_rst)); 
buffer_wire buffer_11583 (.in(n11583), .out(n11583_0));
mux14 mux_6418 (.in({n12743_0, n12732_0/**/, n12717_0, n12705_0, n12698_0, n12693_0, n12686_0, n12666_1, n11516_0, n2239, n2231, n2223, n2135, n2123}), .out(n11584), .config_in(config_chain[22199:22194]), .config_rst(config_rst)); 
buffer_wire buffer_11584 (.in(n11584), .out(n11584_0));
mux14 mux_6419 (.in({n13795_0, n13775_0, n13758_0, n13744_0, n13739_0, n13730_0, n13725_0, n13698_1, n11673_1, n5173, n5165, n5157, n5069/**/, n5057}), .out(n11585), .config_in(config_chain[22205:22200]), .config_rst(config_rst)); 
buffer_wire buffer_11585 (.in(n11585), .out(n11585_0));
mux14 mux_6420 (.in({n12745_0, n12725_0, n12718_0, n12713_0, n12706_0, n12694_0, n12679_0, n12664_1, n11524_0/**/, n2239, n2231, n2223, n2135, n2127}), .out(n11586), .config_in(config_chain[22211:22206]), .config_rst(config_rst)); 
buffer_wire buffer_11586 (.in(n11586), .out(n11586_0));
mux14 mux_6421 (.in({n13793_0, n13766_0/**/, n13761_0, n13752_0, n13747_0, n13733_0, n13716_0, n13700_1, n11675_1, n5173, n5165, n5157, n5069, n5061}), .out(n11587), .config_in(config_chain[22217:22212]), .config_rst(config_rst)); 
buffer_wire buffer_11587 (.in(n11587), .out(n11587_0));
mux13 mux_6422 (.in({n12747_0, n12733_0, n12726_0, n12714_0, n12699_0, n12687_0, n12680_0, n12662_1, n11532_0/**/, n2231, n2223, n2135, n2127}), .out(n11588), .config_in(config_chain[22223:22218]), .config_rst(config_rst)); 
buffer_wire buffer_11588 (.in(n11588), .out(n11588_0));
mux13 mux_6423 (.in({n13791_0, n13774_0, n13769_0, n13755_0, n13738_0, n13724_0, n13719_0, n13702_1/**/, n11677_1, n5165, n5157, n5069, n5061}), .out(n11589), .config_in(config_chain[22229:22224]), .config_rst(config_rst)); 
buffer_wire buffer_11589 (.in(n11589), .out(n11589_0));
mux13 mux_6424 (.in({n12749_0, n12734_0, n12719_0, n12707_0, n12700_0/**/, n12695_0, n12688_0, n12660_1, n11540_0, n2235, n2223, n2135, n2127}), .out(n11590), .config_in(config_chain[22235:22230]), .config_rst(config_rst)); 
buffer_wire buffer_11590 (.in(n11590), .out(n11590_0));
mux13 mux_6425 (.in({n13789_0, n13777_0, n13760_0, n13746_0, n13741_0, n13732_0, n13727_0, n13704_1, n11679_1, n5169/**/, n5157, n5069, n5061}), .out(n11591), .config_in(config_chain[22241:22236]), .config_rst(config_rst)); 
buffer_wire buffer_11591 (.in(n11591), .out(n11591_0));
mux13 mux_6426 (.in({n12751_0, n12727_0, n12720_0, n12715_0, n12708_0, n12681_0, n12658_1, n12606_2, n11548_0, n2235/**/, n2227, n2135, n2127}), .out(n11592), .config_in(config_chain[22247:22242]), .config_rst(config_rst)); 
buffer_wire buffer_11592 (.in(n11592), .out(n11592_0));
mux13 mux_6427 (.in({n13787_0, n13768_0, n13763_0/**/, n13754_0, n13749_0, n13718_0, n13713_0, n13706_1, n11681_1, n5169, n5161, n5069, n5061}), .out(n11593), .config_in(config_chain[22253:22248]), .config_rst(config_rst)); 
buffer_wire buffer_11593 (.in(n11593), .out(n11593_0));
mux13 mux_6428 (.in({n12753_0, n12735_0, n12728_0, n12701_0, n12689_0, n12682_0, n12656_1, n12608_2, n11556_0/**/, n2235, n2227, n2139, n2127}), .out(n11594), .config_in(config_chain[22259:22254]), .config_rst(config_rst)); 
buffer_wire buffer_11594 (.in(n11594), .out(n11594_0));
mux13 mux_6429 (.in({n13785_0, n13776_0, n13771_0, n13740_0, n13735_0, n13726_0, n13721_0, n13708_1, n11683_1, n5169, n5161, n5073, n5061}), .out(n11595), .config_in(config_chain[22265:22260]), .config_rst(config_rst)); 
buffer_wire buffer_11595 (.in(n11595), .out(n11595_0));
mux13 mux_6430 (.in({n12755_0, n12721_0, n12709_0, n12702_0, n12690_0, n12610_2, n12607_0, n12604_2, n11564_0, n2235, n2227, n2139, n2131/**/}), .out(n11596), .config_in(config_chain[22271:22266]), .config_rst(config_rst)); 
buffer_wire buffer_11596 (.in(n11596), .out(n11596_0));
mux3 mux_6431 (.in({n14695_0/**/, n14694_2, n9081}), .out(n11597), .config_in(config_chain[22273:22272]), .config_rst(config_rst)); 
buffer_wire buffer_11597 (.in(n11597), .out(n11597_0));
mux15 mux_6432 (.in({n13015_0, n12979_0, n12972_0, n12965_0, n12958_0, n12946_0, n12930_1/**/, n12868_2, n12865_0, n11486_0, n3213, n3205, n3117, n3109, n3101}), .out(n11598), .config_in(config_chain[22279:22274]), .config_rst(config_rst)); 
buffer_wire buffer_11598 (.in(n11598), .out(n11598_0));
mux15 mux_6433 (.in({n14047_0, n14030_0, n14025_0, n14023_0, n14014_0, n14009_0, n13995_0, n13978_1, n13914_2, n11687_0, n6147, n6139, n6051, n6043, n6035/**/}), .out(n11599), .config_in(config_chain[22285:22280]), .config_rst(config_rst)); 
buffer_wire buffer_11599 (.in(n11599), .out(n11599_0));
mux15 mux_6434 (.in({n12995_0, n12987_0, n12980_0, n12966_0, n12939_0, n12932_0, n12928_1/**/, n12870_2, n12867_0, n11494_0, n3217, n3205, n3117, n3109, n3101}), .out(n11600), .config_in(config_chain[22291:22286]), .config_rst(config_rst)); 
buffer_wire buffer_11600 (.in(n11600), .out(n11600_0));
mux15 mux_6435 (.in({n14067_0, n14045_0, n14038_0, n14033_0, n14017_0, n14000_0, n13986_0, n13981_0, n13958_1, n11689_0, n6151, n6139, n6051/**/, n6043, n6035}), .out(n11601), .config_in(config_chain[22297:22292]), .config_rst(config_rst)); 
buffer_wire buffer_11601 (.in(n11601), .out(n11601_0));
mux15 mux_6436 (.in({n12997_0, n12988_0, n12973_0, n12959_0, n12952_0, n12947_0, n12940_0, n12926_1, n12869_0, n11502_0, n3217, n3209, n3117, n3109/**/, n3101}), .out(n11602), .config_in(config_chain[22303:22298]), .config_rst(config_rst)); 
buffer_wire buffer_11602 (.in(n11602), .out(n11602_0));
mux15 mux_6437 (.in({n14065_0, n14041_0, n14024_0, n14022_0/**/, n14008_0, n14003_0, n13994_0, n13989_0, n13960_1, n11691_0, n6151, n6143, n6051, n6043, n6035}), .out(n11603), .config_in(config_chain[22309:22304]), .config_rst(config_rst)); 
buffer_wire buffer_11603 (.in(n11603), .out(n11603_0));
mux15 mux_6438 (.in({n12999_0, n12981_0, n12974_0, n12967_0, n12960_0, n12948_0, n12933_0, n12924_1/**/, n12871_0, n11510_0, n3217, n3209, n3201, n3109, n3101}), .out(n11604), .config_in(config_chain[22315:22310]), .config_rst(config_rst)); 
buffer_wire buffer_11604 (.in(n11604), .out(n11604_0));
mux15 mux_6439 (.in({n14063_0, n14044_0, n14032_0/**/, n14027_0, n14016_0, n14011_0, n13997_0, n13980_0, n13962_1, n11693_0, n6151, n6143, n6135, n6043, n6035}), .out(n11605), .config_in(config_chain[22321:22316]), .config_rst(config_rst)); 
buffer_wire buffer_11605 (.in(n11605), .out(n11605_0));
mux14 mux_6440 (.in({n13001_0, n12989_0, n12982_0, n12968_0, n12953_0, n12941_0, n12934_0, n12922_1/**/, n11518_0, n3217, n3209, n3201, n3113, n3101}), .out(n11606), .config_in(config_chain[22327:22322]), .config_rst(config_rst)); 
buffer_wire buffer_11606 (.in(n11606), .out(n11606_0));
mux14 mux_6441 (.in({n14061_0, n14040_0, n14035_0, n14019_0, n14002_0, n13988_0, n13983_0, n13964_1, n11695_0, n6151, n6143, n6135, n6047/**/, n6035}), .out(n11607), .config_in(config_chain[22333:22328]), .config_rst(config_rst)); 
buffer_wire buffer_11607 (.in(n11607), .out(n11607_0));
mux14 mux_6442 (.in({n13003_0, n12990_0, n12975_0, n12961_0, n12954_0, n12949_0, n12942_0, n12920_1/**/, n11526_0, n3217, n3209, n3201, n3113, n3105}), .out(n11608), .config_in(config_chain[22339:22334]), .config_rst(config_rst)); 
buffer_wire buffer_11608 (.in(n11608), .out(n11608_0));
mux14 mux_6443 (.in({n14059_0, n14043_0, n14026_0, n14010_0, n14005_0, n13996_0, n13991_0, n13966_1, n11697_0, n6151/**/, n6143, n6135, n6047, n6039}), .out(n11609), .config_in(config_chain[22345:22340]), .config_rst(config_rst)); 
buffer_wire buffer_11609 (.in(n11609), .out(n11609_0));
mux13 mux_6444 (.in({n13005_0, n12983_0, n12976_0, n12969_0, n12962_0, n12950_0, n12935_0, n12918_1/**/, n11534_0, n3209, n3201, n3113, n3105}), .out(n11610), .config_in(config_chain[22351:22346]), .config_rst(config_rst)); 
buffer_wire buffer_11610 (.in(n11610), .out(n11610_0));
mux13 mux_6445 (.in({n14057_0, n14034_0, n14029_0/**/, n14018_0, n14013_0, n13999_0, n13982_0, n13968_1, n11699_0, n6143, n6135, n6047, n6039}), .out(n11611), .config_in(config_chain[22357:22352]), .config_rst(config_rst)); 
buffer_wire buffer_11611 (.in(n11611), .out(n11611_0));
mux13 mux_6446 (.in({n13007_0, n12991_0, n12984_0/**/, n12970_0, n12955_0, n12943_0, n12936_0, n12916_1, n11542_0, n3213, n3201, n3113, n3105}), .out(n11612), .config_in(config_chain[22363:22358]), .config_rst(config_rst)); 
buffer_wire buffer_11612 (.in(n11612), .out(n11612_0));
mux13 mux_6447 (.in({n14055_0, n14042_0, n14037_0, n14021_0, n14004_0, n13990_0, n13985_0, n13970_1, n11701_0, n6147, n6135, n6047, n6039}), .out(n11613), .config_in(config_chain[22369:22364]), .config_rst(config_rst)); 
buffer_wire buffer_11613 (.in(n11613), .out(n11613_0));
mux13 mux_6448 (.in({n13009_0, n12992_0, n12977_0, n12963_0, n12956_0, n12951_0, n12944_0, n12914_1, n11550_0, n3213, n3205/**/, n3113, n3105}), .out(n11614), .config_in(config_chain[22375:22370]), .config_rst(config_rst)); 
buffer_wire buffer_11614 (.in(n11614), .out(n11614_0));
mux13 mux_6449 (.in({n14053_0/**/, n14028_0, n14012_0, n14007_0, n13998_0, n13993_0, n13972_1, n13957_0, n11703_0, n6147, n6139, n6047, n6039}), .out(n11615), .config_in(config_chain[22381:22376]), .config_rst(config_rst)); 
buffer_wire buffer_11615 (.in(n11615), .out(n11615_0));
mux13 mux_6450 (.in({n13011_0, n12985_0, n12978_0, n12971_0, n12964_0, n12937_0, n12912_1, n12864_2, n11558_0, n3213, n3205, n3117, n3105/**/}), .out(n11616), .config_in(config_chain[22387:22382]), .config_rst(config_rst)); 
buffer_wire buffer_11616 (.in(n11616), .out(n11616_0));
mux13 mux_6451 (.in({n14051_0, n14036_0, n14031_0, n14020_0, n14015_0, n13984_0, n13979_0, n13974_1, n11705_0/**/, n6147, n6139, n6051, n6039}), .out(n11617), .config_in(config_chain[22393:22388]), .config_rst(config_rst)); 
buffer_wire buffer_11617 (.in(n11617), .out(n11617_0));
mux13 mux_6452 (.in({n13013_0, n12993_0, n12986_0, n12957_0, n12945_0/**/, n12938_0, n12866_2, n12862_2, n11566_0, n3213, n3205, n3117, n3109}), .out(n11618), .config_in(config_chain[22399:22394]), .config_rst(config_rst)); 
buffer_wire buffer_11618 (.in(n11618), .out(n11618_0));
mux3 mux_6453 (.in({n14697_0, n14696_2, n9081}), .out(n11619), .config_in(config_chain[22401:22400]), .config_rst(config_rst)); 
buffer_wire buffer_11619 (.in(n11619), .out(n11619_0));
mux15 mux_6454 (.in({n13275_0, n13253_0, n13246_0, n13217_0, n13210_0, n13203_0, n13196_0, n13188_1, n13126_2, n11488_0, n4191, n4183, n4095, n4087, n4079}), .out(n11620), .config_in(config_chain[22407:22402]), .config_rst(config_rst)); 
buffer_wire buffer_11620 (.in(n11620), .out(n11620_0));
mux16 mux_6455 (.in({n14313_0, n14297_0, n14292_0, n14288_0, n14284_0, n14269_0, n14259_0, n14254_0, n14242_1, n14201_0, n11709_0, n7125, n7117/**/, n7029, n7021, n7013}), .out(n11621), .config_in(config_chain[22413:22408]), .config_rst(config_rst)); 
buffer_wire buffer_11621 (.in(n11621), .out(n11621_0));
mux15 mux_6456 (.in({n13255_0, n13239_0/**/, n13232_0, n13225_0, n13218_0, n13204_0, n13186_1, n13128_2, n13125_0, n11496_0, n4195, n4183, n4095, n4087, n4079}), .out(n11622), .config_in(config_chain[22419:22414]), .config_rst(config_rst)); 
buffer_wire buffer_11622 (.in(n11622), .out(n11622_0));
mux16 mux_6457 (.in({n14331_0, n14310_0, n14306_0, n14291_0, n14283_0, n14278_0, n14253_0, n14248_0/**/, n14224_1, n14223_0, n11711_0, n7125, n7117, n7029, n7021, n7013}), .out(n11623), .config_in(config_chain[22425:22420]), .config_rst(config_rst)); 
buffer_wire buffer_11623 (.in(n11623), .out(n11623_0));
mux15 mux_6458 (.in({n13257_0, n13247_0, n13240_0, n13226_0, n13211_0, n13197_0, n13190_0, n13184_1, n13127_0, n11504_0, n4195, n4187/**/, n4095, n4087, n4079}), .out(n11624), .config_in(config_chain[22431:22426]), .config_rst(config_rst)); 
buffer_wire buffer_11624 (.in(n11624), .out(n11624_0));
mux15 mux_6459 (.in({n14329_0, n14305_0, n14300_0/**/, n14277_0, n14272_0, n14262_0, n14247_0, n14245_0, n14226_1, n11713_0, n7125, n7117, n7029, n7021, n7013}), .out(n11625), .config_in(config_chain[22437:22432]), .config_rst(config_rst)); 
buffer_wire buffer_11625 (.in(n11625), .out(n11625_0));
mux15 mux_6460 (.in({n13259_0, n13248_0/**/, n13233_0, n13219_0, n13212_0, n13205_0, n13198_0, n13182_1, n13129_0, n11512_0, n4195, n4187, n4179, n4087, n4079}), .out(n11626), .config_in(config_chain[22443:22438]), .config_rst(config_rst)); 
buffer_wire buffer_11626 (.in(n11626), .out(n11626_0));
mux15 mux_6461 (.in({n14327_0, n14299_0, n14294_0, n14286_0, n14271_0, n14267_0, n14261_0, n14256_0, n14228_1, n11715_0, n7125, n7117/**/, n7029, n7021, n7013}), .out(n11627), .config_in(config_chain[22449:22444]), .config_rst(config_rst)); 
buffer_wire buffer_11627 (.in(n11627), .out(n11627_0));
mux14 mux_6462 (.in({n13261_0, n13241_0, n13234_0, n13227_0, n13220_0/**/, n13206_0, n13191_0, n13180_1, n11520_0, n4195, n4187, n4179, n4091, n4079}), .out(n11628), .config_in(config_chain[22455:22450]), .config_rst(config_rst)); 
buffer_wire buffer_11628 (.in(n11628), .out(n11628_0));
mux15 mux_6463 (.in({n14325_0, n14308_0, n14293_0, n14289_0, n14285_0/**/, n14280_0, n14255_0, n14250_0, n14230_1, n11717_0, n7125, n7117, n7029, n7021, n7013}), .out(n11629), .config_in(config_chain[22461:22456]), .config_rst(config_rst)); 
buffer_wire buffer_11629 (.in(n11629), .out(n11629_0));
mux14 mux_6464 (.in({n13263_0, n13249_0, n13242_0, n13228_0, n13213_0, n13199_0, n13192_0, n13178_1, n11528_0/**/, n4195, n4187, n4179, n4091, n4083}), .out(n11630), .config_in(config_chain[22467:22462]), .config_rst(config_rst)); 
buffer_wire buffer_11630 (.in(n11630), .out(n11630_0));
mux15 mux_6465 (.in({n14323_0, n14311_0/**/, n14307_0, n14302_0, n14279_0, n14274_0, n14264_0, n14249_0, n14232_1, n11719_0, n7129, n7121, n7113, n7025, n7017}), .out(n11631), .config_in(config_chain[22473:22468]), .config_rst(config_rst)); 
buffer_wire buffer_11631 (.in(n11631), .out(n11631_0));
mux13 mux_6466 (.in({n13265_0, n13250_0, n13235_0, n13221_0, n13214_0/**/, n13207_0, n13200_0, n13176_1, n11536_0, n4187, n4179, n4091, n4083}), .out(n11632), .config_in(config_chain[22479:22474]), .config_rst(config_rst)); 
buffer_wire buffer_11632 (.in(n11632), .out(n11632_0));
mux15 mux_6467 (.in({n14321_0, n14301_0, n14296_0/**/, n14273_0, n14268_0, n14263_0, n14258_0, n14234_1, n14200_1, n11721_0, n7129, n7121, n7113, n7025, n7017}), .out(n11633), .config_in(config_chain[22485:22480]), .config_rst(config_rst)); 
buffer_wire buffer_11633 (.in(n11633), .out(n11633_0));
mux13 mux_6468 (.in({n13267_0, n13243_0, n13236_0/**/, n13229_0, n13222_0, n13208_0, n13193_0, n13174_1, n11544_0, n4191, n4179, n4091, n4083}), .out(n11634), .config_in(config_chain[22491:22486]), .config_rst(config_rst)); 
buffer_wire buffer_11634 (.in(n11634), .out(n11634_0));
mux15 mux_6469 (.in({n14319_0, n14295_0, n14290_0, n14287_0, n14282_0/**/, n14257_0, n14252_0, n14236_1, n14222_1, n11723_0, n7129, n7121, n7113, n7025, n7017}), .out(n11635), .config_in(config_chain[22497:22492]), .config_rst(config_rst)); 
buffer_wire buffer_11635 (.in(n11635), .out(n11635_0));
mux13 mux_6470 (.in({n13269_0, n13251_0, n13244_0, n13230_0, n13215_0, n13201_0/**/, n13194_0, n13172_1, n11552_0, n4191, n4183, n4091, n4083}), .out(n11636), .config_in(config_chain[22503:22498]), .config_rst(config_rst)); 
buffer_wire buffer_11636 (.in(n11636), .out(n11636_0));
mux15 mux_6471 (.in({n14317_0, n14309_0, n14304_0, n14281_0, n14276_0, n14251_0, n14246_0/**/, n14244_1, n14238_1, n11725_0, n7129, n7121, n7113, n7025, n7017}), .out(n11637), .config_in(config_chain[22509:22504]), .config_rst(config_rst)); 
buffer_wire buffer_11637 (.in(n11637), .out(n11637_0));
mux13 mux_6472 (.in({n13271_0/**/, n13252_0, n13237_0, n13223_0, n13216_0, n13209_0, n13202_0, n13170_1, n11560_0, n4191, n4183, n4095, n4083}), .out(n11638), .config_in(config_chain[22515:22510]), .config_rst(config_rst)); 
buffer_wire buffer_11638 (.in(n11638), .out(n11638_0));
mux15 mux_6473 (.in({n14315_0/**/, n14303_0, n14298_0, n14275_0, n14270_0, n14266_0, n14265_0, n14260_0, n14240_1, n11727_0, n7129, n7121, n7113, n7025, n7017}), .out(n11639), .config_in(config_chain[22521:22516]), .config_rst(config_rst)); 
buffer_wire buffer_11639 (.in(n11639), .out(n11639_0));
mux13 mux_6474 (.in({n13273_0/**/, n13245_0, n13238_0, n13231_0, n13224_0, n13195_0, n13124_2, n13122_2, n11568_0, n4191, n4183, n4095, n4087}), .out(n11640), .config_in(config_chain[22527:22522]), .config_rst(config_rst)); 
buffer_wire buffer_11640 (.in(n11640), .out(n11640_0));
mux3 mux_6475 (.in({n14727_0, n14726_1, n9081}), .out(n11641), .config_in(config_chain[22529:22528]), .config_rst(config_rst)); 
buffer_wire buffer_11641 (.in(n11641), .out(n11641_0));
mux15 mux_6476 (.in({n13537_0, n13507_0, n13500_0, n13493_0, n13486_0, n13457_0, n13450_0, n13448_1/**/, n13386_2, n11490_1, n5169, n5161, n5073, n5065, n5057}), .out(n11642), .config_in(config_chain[22535:22530]), .config_rst(config_rst)); 
buffer_wire buffer_11642 (.in(n11642), .out(n11642_0));
mux16 mux_6477 (.in({n14575_0, n14567_0, n14562_0, n14539_0, n14534_0, n14530_0, n14526_0, n14511_0, n14506_1, n14433_0, n11729_0, n8103/**/, n8095, n8007, n7999, n7991}), .out(n11643), .config_in(config_chain[22541:22536]), .config_rst(config_rst)); 
buffer_wire buffer_11643 (.in(n11643), .out(n11643_0));
mux15 mux_6478 (.in({n13517_0/**/, n13515_0, n13508_0, n13479_0, n13472_0, n13465_0, n13458_0, n13446_1, n13388_2, n11498_1, n5173, n5161, n5073, n5065, n5057}), .out(n11644), .config_in(config_chain[22547:22542]), .config_rst(config_rst)); 
buffer_wire buffer_11644 (.in(n11644), .out(n11644_0));
mux16 mux_6479 (.in({n14593_0, n14561_0, n14556_0/**/, n14552_0, n14548_0, n14533_0, n14525_0, n14520_0, n14488_1, n14465_0, n11731_0, n8103, n8095, n8007, n7999, n7991}), .out(n11645), .config_in(config_chain[22553:22548]), .config_rst(config_rst)); 
buffer_wire buffer_11645 (.in(n11645), .out(n11645_0));
mux15 mux_6480 (.in({n13519_0, n13501_0, n13494_0/**/, n13487_0, n13480_0, n13466_0, n13451_0, n13444_1, n13387_0, n11506_1, n5173, n5165, n5073, n5065, n5057}), .out(n11646), .config_in(config_chain[22559:22554]), .config_rst(config_rst)); 
buffer_wire buffer_11646 (.in(n11646), .out(n11646_0));
mux15 mux_6481 (.in({n14591_0, n14570_0/**/, n14555_0, n14547_0, n14542_0, n14519_0, n14514_0, n14490_1, n14487_0, n11733_0, n8103, n8095, n8007, n7999, n7991}), .out(n11647), .config_in(config_chain[22565:22560]), .config_rst(config_rst)); 
buffer_wire buffer_11647 (.in(n11647), .out(n11647_0));
mux15 mux_6482 (.in({n13521_0, n13509_0, n13502_0, n13488_0, n13473_0, n13459_0/**/, n13452_0, n13442_1, n13389_0, n11514_1, n5173, n5165, n5157, n5065, n5057}), .out(n11648), .config_in(config_chain[22571:22566]), .config_rst(config_rst)); 
buffer_wire buffer_11648 (.in(n11648), .out(n11648_0));
mux15 mux_6483 (.in({n14589_0, n14569_0, n14564_0, n14541_0, n14536_0, n14528_0, n14513_0, n14509_0, n14492_1, n11735_0, n8103, n8095, n8007, n7999, n7991}), .out(n11649), .config_in(config_chain[22577:22572]), .config_rst(config_rst)); 
buffer_wire buffer_11649 (.in(n11649), .out(n11649_0));
mux14 mux_6484 (.in({n13523_0, n13510_0, n13495_0, n13481_0, n13474_0, n13467_0, n13460_0, n13440_1, n11522_1, n5173, n5165/**/, n5157, n5069, n5057}), .out(n11650), .config_in(config_chain[22583:22578]), .config_rst(config_rst)); 
buffer_wire buffer_11650 (.in(n11650), .out(n11650_0));
mux15 mux_6485 (.in({n14587_0, n14563_0, n14558_0, n14550_0, n14535_0, n14531_0, n14527_0, n14522_0, n14494_1, n11737_0/**/, n8103, n8095, n8007, n7999, n7991}), .out(n11651), .config_in(config_chain[22589:22584]), .config_rst(config_rst)); 
buffer_wire buffer_11651 (.in(n11651), .out(n11651_0));
mux14 mux_6486 (.in({n13525_0, n13503_0, n13496_0, n13489_0, n13482_0, n13468_0, n13453_0, n13438_1, n11530_1/**/, n5173, n5165, n5157, n5069, n5061}), .out(n11652), .config_in(config_chain[22595:22590]), .config_rst(config_rst)); 
buffer_wire buffer_11652 (.in(n11652), .out(n11652_0));
mux15 mux_6487 (.in({n14585_0, n14572_0, n14557_0, n14553_0, n14549_0, n14544_0, n14521_0, n14516_0, n14496_1, n11739_0, n8107, n8099, n8091, n8003/**/, n7995}), .out(n11653), .config_in(config_chain[22601:22596]), .config_rst(config_rst)); 
buffer_wire buffer_11653 (.in(n11653), .out(n11653_0));
mux13 mux_6488 (.in({n13527_0, n13511_0, n13504_0, n13490_0, n13475_0, n13461_0, n13454_0, n13436_1, n11538_1/**/, n5165, n5157, n5069, n5061}), .out(n11654), .config_in(config_chain[22607:22602]), .config_rst(config_rst)); 
buffer_wire buffer_11654 (.in(n11654), .out(n11654_0));
mux15 mux_6489 (.in({n14583_0, n14571_0, n14566_0, n14543_0, n14538_0, n14515_0, n14510_0, n14498_1, n14432_2, n11741_0, n8107, n8099, n8091/**/, n8003, n7995}), .out(n11655), .config_in(config_chain[22613:22608]), .config_rst(config_rst)); 
buffer_wire buffer_11655 (.in(n11655), .out(n11655_0));
mux13 mux_6490 (.in({n13529_0, n13512_0, n13497_0, n13483_0, n13476_0/**/, n13469_0, n13462_0, n13434_1, n11546_1, n5169, n5157, n5069, n5061}), .out(n11656), .config_in(config_chain[22619:22614]), .config_rst(config_rst)); 
buffer_wire buffer_11656 (.in(n11656), .out(n11656_0));
mux15 mux_6491 (.in({n14581_0, n14565_0, n14560_0, n14537_0, n14532_0, n14529_0, n14524_0, n14500_1, n14464_1/**/, n11743_0, n8107, n8099, n8091, n8003, n7995}), .out(n11657), .config_in(config_chain[22625:22620]), .config_rst(config_rst)); 
buffer_wire buffer_11657 (.in(n11657), .out(n11657_0));
mux13 mux_6492 (.in({n13531_0, n13505_0, n13498_0, n13491_0, n13484_0, n13470_0, n13455_0, n13432_1, n11554_1/**/, n5169, n5161, n5069, n5061}), .out(n11658), .config_in(config_chain[22631:22626]), .config_rst(config_rst)); 
buffer_wire buffer_11658 (.in(n11658), .out(n11658_0));
mux15 mux_6493 (.in({n14579_0, n14559_0, n14554_0, n14551_0, n14546_0/**/, n14523_0, n14518_0, n14502_1, n14486_1, n11745_0, n8107, n8099, n8091, n8003, n7995}), .out(n11659), .config_in(config_chain[22637:22632]), .config_rst(config_rst)); 
buffer_wire buffer_11659 (.in(n11659), .out(n11659_0));
mux13 mux_6494 (.in({n13533_0, n13513_0, n13506_0, n13492_0, n13477_0, n13463_0/**/, n13456_0, n13430_1, n11562_1, n5169, n5161, n5073, n5061}), .out(n11660), .config_in(config_chain[22643:22638]), .config_rst(config_rst)); 
buffer_wire buffer_11660 (.in(n11660), .out(n11660_0));
mux15 mux_6495 (.in({n14577_0, n14573_0, n14568_0, n14545_0, n14540_0, n14517_0, n14512_0, n14508_1, n14504_1, n11747_0, n8107, n8099, n8091/**/, n8003, n7995}), .out(n11661), .config_in(config_chain[22649:22644]), .config_rst(config_rst)); 
buffer_wire buffer_11661 (.in(n11661), .out(n11661_0));
mux13 mux_6496 (.in({n13535_0, n13514_0, n13499_0, n13485_0, n13478_0, n13471_0, n13464_0, n13384_2, n11570_1/**/, n5169, n5161, n5073, n5065}), .out(n11662), .config_in(config_chain[22655:22650]), .config_rst(config_rst)); 
buffer_wire buffer_11662 (.in(n11662), .out(n11662_0));
mux3 mux_6497 (.in({n14749_0, n14748_1, n9081}), .out(n11663), .config_in(config_chain[22657:22656]), .config_rst(config_rst)); 
buffer_wire buffer_11663 (.in(n11663), .out(n11663_0));
mux15 mux_6498 (.in({n13801_0, n13778_0/**/, n13771_0, n13764_0, n13750_0, n13735_0, n13721_0, n13714_0, n13710_1, n11576_1, n6147, n6139, n6051, n6043, n6035}), .out(n11664), .config_in(config_chain[22663:22658]), .config_rst(config_rst)); 
buffer_wire buffer_11664 (.in(n11664), .out(n11664_0));
mux4 mux_6499 (.in({n14835_0, n14750_1, n9085, n8969/**/}), .out(n11665), .config_in(config_chain[22665:22664]), .config_rst(config_rst)); 
buffer_wire buffer_11665 (.in(n11665), .out(n11665_0));
mux15 mux_6500 (.in({n13781_0, n13772_0, n13757_0, n13743_0, n13736_0, n13729_0, n13722_0, n13708_1, n13650_2, n11578_1, n6151, n6139/**/, n6051, n6043, n6035}), .out(n11666), .config_in(config_chain[22671:22666]), .config_rst(config_rst)); 
buffer_wire buffer_11666 (.in(n11666), .out(n11666_0));
mux3 mux_6501 (.in({n14837_0, n14752_1, n8969}), .out(n11667), .config_in(config_chain[22673:22672]), .config_rst(config_rst)); 
buffer_wire buffer_11667 (.in(n11667), .out(n11667_0));
mux15 mux_6502 (.in({n13783_0, n13779_0, n13765_0, n13758_0, n13751_0, n13744_0, n13730_0, n13715_0, n13706_1, n11580_1, n6151, n6143, n6051, n6043/**/, n6035}), .out(n11668), .config_in(config_chain[22679:22674]), .config_rst(config_rst)); 
buffer_wire buffer_11668 (.in(n11668), .out(n11668_0));
mux3 mux_6503 (.in({n14839_0, n14754_1/**/, n8973}), .out(n11669), .config_in(config_chain[22681:22680]), .config_rst(config_rst)); 
buffer_wire buffer_11669 (.in(n11669), .out(n11669_0));
mux15 mux_6504 (.in({n13785_0, n13773_0, n13766_0, n13752_0, n13737_0, n13723_0, n13716_0, n13704_1, n13651_0, n11582_1/**/, n6151, n6143, n6135, n6043, n6035}), .out(n11670), .config_in(config_chain[22687:22682]), .config_rst(config_rst)); 
buffer_wire buffer_11670 (.in(n11670), .out(n11670_0));
mux3 mux_6505 (.in({n14841_0/**/, n14756_1, n8977}), .out(n11671), .config_in(config_chain[22689:22688]), .config_rst(config_rst)); 
buffer_wire buffer_11671 (.in(n11671), .out(n11671_0));
mux14 mux_6506 (.in({n13787_0, n13774_0, n13759_0, n13745_0, n13738_0, n13731_0, n13724_0, n13702_1, n11584_1, n6151, n6143, n6135, n6047, n6035/**/}), .out(n11672), .config_in(config_chain[22695:22690]), .config_rst(config_rst)); 
buffer_wire buffer_11672 (.in(n11672), .out(n11672_0));
mux3 mux_6507 (.in({n14843_0, n14758_1, n8981/**/}), .out(n11673), .config_in(config_chain[22697:22696]), .config_rst(config_rst)); 
buffer_wire buffer_11673 (.in(n11673), .out(n11673_0));
mux14 mux_6508 (.in({n13789_0, n13767_0, n13760_0, n13753_0, n13746_0, n13732_0, n13717_0, n13700_1, n11586_1/**/, n6151, n6143, n6135, n6047, n6039}), .out(n11674), .config_in(config_chain[22703:22698]), .config_rst(config_rst)); 
buffer_wire buffer_11674 (.in(n11674), .out(n11674_0));
mux3 mux_6509 (.in({n14845_0/**/, n14760_1, n8985}), .out(n11675), .config_in(config_chain[22705:22704]), .config_rst(config_rst)); 
buffer_wire buffer_11675 (.in(n11675), .out(n11675_0));
mux13 mux_6510 (.in({n13791_0, n13775_0, n13768_0, n13754_0, n13739_0, n13725_0, n13718_0, n13698_1, n11588_1/**/, n6143, n6135, n6047, n6039}), .out(n11676), .config_in(config_chain[22711:22706]), .config_rst(config_rst)); 
buffer_wire buffer_11676 (.in(n11676), .out(n11676_0));
mux3 mux_6511 (.in({n14847_0, n14762_1/**/, n8985}), .out(n11677), .config_in(config_chain[22713:22712]), .config_rst(config_rst)); 
buffer_wire buffer_11677 (.in(n11677), .out(n11677_0));
mux13 mux_6512 (.in({n13793_0, n13776_0, n13761_0, n13747_0/**/, n13740_0, n13733_0, n13726_0, n13696_1, n11590_1, n6147, n6135, n6047, n6039}), .out(n11678), .config_in(config_chain[22719:22714]), .config_rst(config_rst)); 
buffer_wire buffer_11678 (.in(n11678), .out(n11678_0));
mux3 mux_6513 (.in({n14849_0/**/, n14764_1, n9069}), .out(n11679), .config_in(config_chain[22721:22720]), .config_rst(config_rst)); 
buffer_wire buffer_11679 (.in(n11679), .out(n11679_0));
mux13 mux_6514 (.in({n13795_0, n13769_0, n13762_0, n13755_0, n13748_0, n13719_0, n13712_1, n13694_1, n11592_1, n6147, n6139, n6047, n6039/**/}), .out(n11680), .config_in(config_chain[22727:22722]), .config_rst(config_rst)); 
buffer_wire buffer_11680 (.in(n11680), .out(n11680_0));
mux3 mux_6515 (.in({n14851_0, n14766_1, n9073}), .out(n11681), .config_in(config_chain[22729:22728]), .config_rst(config_rst)); 
buffer_wire buffer_11681 (.in(n11681), .out(n11681_0));
mux13 mux_6516 (.in({n13797_0, n13777_0, n13770_0, n13741_0, n13734_0, n13727_0, n13720_0, n13692_1, n11594_1/**/, n6147, n6139, n6051, n6039}), .out(n11682), .config_in(config_chain[22735:22730]), .config_rst(config_rst)); 
buffer_wire buffer_11682 (.in(n11682), .out(n11682_0));
mux3 mux_6517 (.in({n14853_0/**/, n14768_1, n9077}), .out(n11683), .config_in(config_chain[22737:22736]), .config_rst(config_rst)); 
buffer_wire buffer_11683 (.in(n11683), .out(n11683_0));
mux13 mux_6518 (.in({n13799_0, n13763_0, n13756_0, n13749_0, n13742_0, n13728_0, n13713_0, n13648_2, n11572_1, n6147, n6139/**/, n6051, n6043}), .out(n11684), .config_in(config_chain[22743:22738]), .config_rst(config_rst)); 
buffer_wire buffer_11684 (.in(n11684), .out(n11684_0));
mux3 mux_6519 (.in({n14771_0, n14770_1, n9081}), .out(n11685), .config_in(config_chain[22745:22744]), .config_rst(config_rst)); 
buffer_wire buffer_11685 (.in(n11685), .out(n11685_0));
mux15 mux_6520 (.in({n14067_0, n14031_0, n14024_0, n14022_0, n14015_0, n14008_0, n13994_0, n13979_0, n13976_1/**/, n11598_1, n7125, n7117, n7029, n7021, n7013}), .out(n11686), .config_in(config_chain[22751:22746]), .config_rst(config_rst)); 
buffer_wire buffer_11686 (.in(n11686), .out(n11686_0));
mux4 mux_6521 (.in({n14773_0, n14772_0, n9085, n8969/**/}), .out(n11687), .config_in(config_chain[22753:22752]), .config_rst(config_rst)); 
buffer_wire buffer_11687 (.in(n11687), .out(n11687_0));
mux15 mux_6522 (.in({n14047_0, n14044_0, n14039_0, n14032_0, n14016_0, n14001_0, n13987_0, n13980_0, n13974_1, n11600_1, n7129/**/, n7117, n7029, n7021, n7013}), .out(n11688), .config_in(config_chain[22759:22754]), .config_rst(config_rst)); 
buffer_wire buffer_11688 (.in(n11688), .out(n11688_0));
mux3 mux_6523 (.in({n14775_0, n14774_0, n8973}), .out(n11689), .config_in(config_chain[22761:22760]), .config_rst(config_rst)); 
buffer_wire buffer_11689 (.in(n11689), .out(n11689_0));
mux15 mux_6524 (.in({n14049_0, n14040_0, n14025_0, n14023_0, n14009_0, n14002_0, n13995_0, n13988_0, n13972_1, n11602_1, n7129, n7121, n7029/**/, n7021, n7013}), .out(n11690), .config_in(config_chain[22767:22762]), .config_rst(config_rst)); 
buffer_wire buffer_11690 (.in(n11690), .out(n11690_0));
mux3 mux_6525 (.in({n14777_0, n14776_0, n8973/**/}), .out(n11691), .config_in(config_chain[22769:22768]), .config_rst(config_rst)); 
buffer_wire buffer_11691 (.in(n11691), .out(n11691_0));
mux15 mux_6526 (.in({n14051_0, n14045_0, n14033_0, n14026_0, n14017_0/**/, n14010_0, n13996_0, n13981_0, n13970_1, n11604_1, n7129, n7121, n7113, n7021, n7013}), .out(n11692), .config_in(config_chain[22775:22770]), .config_rst(config_rst)); 
buffer_wire buffer_11692 (.in(n11692), .out(n11692_0));
mux3 mux_6527 (.in({n14779_0, n14778_0/**/, n8977}), .out(n11693), .config_in(config_chain[22777:22776]), .config_rst(config_rst)); 
buffer_wire buffer_11693 (.in(n11693), .out(n11693_0));
mux14 mux_6528 (.in({n14053_0, n14041_0, n14034_0, n14018_0, n14003_0, n13989_0, n13982_0/**/, n13968_1, n11606_1, n7129, n7121, n7113, n7025, n7013}), .out(n11694), .config_in(config_chain[22783:22778]), .config_rst(config_rst)); 
buffer_wire buffer_11694 (.in(n11694), .out(n11694_0));
mux3 mux_6529 (.in({n14781_0, n14780_0, n8981}), .out(n11695), .config_in(config_chain[22785:22784]), .config_rst(config_rst)); 
buffer_wire buffer_11695 (.in(n11695), .out(n11695_0));
mux14 mux_6530 (.in({n14055_0, n14042_0, n14027_0, n14011_0, n14004_0, n13997_0, n13990_0, n13966_1, n11608_1, n7129, n7121, n7113, n7025/**/, n7017}), .out(n11696), .config_in(config_chain[22791:22786]), .config_rst(config_rst)); 
buffer_wire buffer_11696 (.in(n11696), .out(n11696_0));
mux3 mux_6531 (.in({n14783_0, n14782_0, n8985}), .out(n11697), .config_in(config_chain[22793:22792]), .config_rst(config_rst)); 
buffer_wire buffer_11697 (.in(n11697), .out(n11697_0));
mux13 mux_6532 (.in({n14057_0, n14035_0, n14028_0, n14019_0, n14012_0, n13998_0, n13983_0, n13964_1, n11610_1/**/, n7121, n7113, n7025, n7017}), .out(n11698), .config_in(config_chain[22799:22794]), .config_rst(config_rst)); 
buffer_wire buffer_11698 (.in(n11698), .out(n11698_0));
mux3 mux_6533 (.in({n14785_0, n14784_0/**/, n9069}), .out(n11699), .config_in(config_chain[22801:22800]), .config_rst(config_rst)); 
buffer_wire buffer_11699 (.in(n11699), .out(n11699_0));
mux13 mux_6534 (.in({n14059_0, n14043_0, n14036_0, n14020_0, n14005_0/**/, n13991_0, n13984_0, n13962_1, n11612_1, n7125, n7113, n7025, n7017}), .out(n11700), .config_in(config_chain[22807:22802]), .config_rst(config_rst)); 
buffer_wire buffer_11700 (.in(n11700), .out(n11700_0));
mux3 mux_6535 (.in({n14787_0, n14786_0, n9069}), .out(n11701), .config_in(config_chain[22809:22808]), .config_rst(config_rst)); 
buffer_wire buffer_11701 (.in(n11701), .out(n11701_0));
mux13 mux_6536 (.in({n14061_0, n14029_0, n14013_0, n14006_0, n13999_0/**/, n13992_0, n13960_1, n13956_1, n11614_1, n7125, n7117, n7025, n7017}), .out(n11702), .config_in(config_chain[22815:22810]), .config_rst(config_rst)); 
buffer_wire buffer_11702 (.in(n11702), .out(n11702_0));
mux3 mux_6537 (.in({n14789_0, n14788_0/**/, n9073}), .out(n11703), .config_in(config_chain[22817:22816]), .config_rst(config_rst)); 
buffer_wire buffer_11703 (.in(n11703), .out(n11703_0));
mux13 mux_6538 (.in({n14063_0, n14037_0, n14030_0, n14021_0, n14014_0, n13985_0, n13978_1, n13958_1, n11616_1, n7125, n7117, n7029, n7017}), .out(n11704), .config_in(config_chain[22823:22818]), .config_rst(config_rst)); 
buffer_wire buffer_11704 (.in(n11704), .out(n11704_0));
mux3 mux_6539 (.in({n14791_0, n14790_0/**/, n9077}), .out(n11705), .config_in(config_chain[22825:22824]), .config_rst(config_rst)); 
buffer_wire buffer_11705 (.in(n11705), .out(n11705_0));
mux13 mux_6540 (.in({n14065_0, n14038_0/**/, n14007_0, n14000_0, n13993_0, n13986_0, n13957_0, n13914_2, n11574_1, n7125, n7117, n7029, n7021}), .out(n11706), .config_in(config_chain[22831:22826]), .config_rst(config_rst)); 
buffer_wire buffer_11706 (.in(n11706), .out(n11706_0));
mux3 mux_6541 (.in({n14793_0, n14792_0/**/, n9085}), .out(n11707), .config_in(config_chain[22833:22832]), .config_rst(config_rst)); 
buffer_wire buffer_11707 (.in(n11707), .out(n11707_0));
mux16 mux_6542 (.in({n14331_0, n14296_0, n14293_0, n14289_0, n14285_0, n14268_0, n14258_0, n14255_0, n14240_1, n14200_1, n11620_1, n8103, n8095, n8007, n7999/**/, n7991}), .out(n11708), .config_in(config_chain[22839:22834]), .config_rst(config_rst)); 
buffer_wire buffer_11708 (.in(n11708), .out(n11708_0));
mux4 mux_6543 (.in({n14795_0, n14794_0, n9085, n8969}), .out(n11709), .config_in(config_chain[22841:22840]), .config_rst(config_rst)); 
buffer_wire buffer_11709 (.in(n11709), .out(n11709_0));
mux16 mux_6544 (.in({n14313_0, n14311_0, n14307_0, n14290_0, n14282_0, n14279_0, n14252_0, n14249_0, n14238_1, n14222_1, n11622_1, n8103, n8095, n8007, n7999, n7991}), .out(n11710), .config_in(config_chain[22847:22842]), .config_rst(config_rst)); 
buffer_wire buffer_11710 (.in(n11710), .out(n11710_0));
mux3 mux_6545 (.in({n14797_0, n14796_0, n8973}), .out(n11711), .config_in(config_chain[22849:22848]), .config_rst(config_rst)); 
buffer_wire buffer_11711 (.in(n11711), .out(n11711_0));
mux15 mux_6546 (.in({n14315_0, n14304_0/**/, n14301_0, n14276_0, n14273_0, n14263_0, n14246_0, n14244_1, n14236_1, n11624_1, n8103, n8095, n8007, n7999, n7991}), .out(n11712), .config_in(config_chain[22855:22850]), .config_rst(config_rst)); 
buffer_wire buffer_11712 (.in(n11712), .out(n11712_0));
mux3 mux_6547 (.in({n14799_0/**/, n14798_0, n8977}), .out(n11713), .config_in(config_chain[22857:22856]), .config_rst(config_rst)); 
buffer_wire buffer_11713 (.in(n11713), .out(n11713_0));
mux15 mux_6548 (.in({n14317_0, n14298_0, n14295_0/**/, n14287_0, n14270_0, n14266_0, n14260_0, n14257_0, n14234_1, n11626_1, n8103, n8095, n8007, n7999, n7991}), .out(n11714), .config_in(config_chain[22863:22858]), .config_rst(config_rst)); 
buffer_wire buffer_11714 (.in(n11714), .out(n11714_0));
mux3 mux_6549 (.in({n14801_0, n14800_0, n8977}), .out(n11715), .config_in(config_chain[22865:22864]), .config_rst(config_rst)); 
buffer_wire buffer_11715 (.in(n11715), .out(n11715_0));
mux15 mux_6550 (.in({n14319_0, n14309_0, n14292_0, n14288_0, n14284_0, n14281_0, n14254_0, n14251_0, n14232_1, n11628_1, n8103, n8095, n8007, n7999, n7991}), .out(n11716), .config_in(config_chain[22871:22866]), .config_rst(config_rst)); 
buffer_wire buffer_11716 (.in(n11716), .out(n11716_0));
mux3 mux_6551 (.in({n14803_0, n14802_0, n8981}), .out(n11717), .config_in(config_chain[22873:22872]), .config_rst(config_rst)); 
buffer_wire buffer_11717 (.in(n11717), .out(n11717_0));
mux15 mux_6552 (.in({n14321_0, n14310_0, n14306_0, n14303_0, n14278_0, n14275_0, n14265_0, n14248_0, n14230_1, n11630_1, n8107, n8099, n8091, n8003, n7995}), .out(n11718), .config_in(config_chain[22879:22874]), .config_rst(config_rst)); 
buffer_wire buffer_11718 (.in(n11718), .out(n11718_0));
mux3 mux_6553 (.in({n14805_0, n14804_0/**/, n8985}), .out(n11719), .config_in(config_chain[22881:22880]), .config_rst(config_rst)); 
buffer_wire buffer_11719 (.in(n11719), .out(n11719_0));
mux15 mux_6554 (.in({n14323_0, n14300_0, n14297_0, n14272_0, n14269_0, n14262_0, n14259_0, n14228_1, n14201_0, n11632_1, n8107, n8099, n8091, n8003, n7995}), .out(n11720), .config_in(config_chain[22887:22882]), .config_rst(config_rst)); 
buffer_wire buffer_11720 (.in(n11720), .out(n11720_0));
mux3 mux_6555 (.in({n14807_0, n14806_0, n9069}), .out(n11721), .config_in(config_chain[22889:22888]), .config_rst(config_rst)); 
buffer_wire buffer_11721 (.in(n11721), .out(n11721_0));
mux15 mux_6556 (.in({n14325_0, n14294_0, n14291_0, n14286_0, n14283_0/**/, n14256_0, n14253_0, n14226_1, n14223_0, n11634_1, n8107, n8099, n8091, n8003, n7995}), .out(n11722), .config_in(config_chain[22895:22890]), .config_rst(config_rst)); 
buffer_wire buffer_11722 (.in(n11722), .out(n11722_0));
mux3 mux_6557 (.in({n14809_0, n14808_0, n9073/**/}), .out(n11723), .config_in(config_chain[22897:22896]), .config_rst(config_rst)); 
buffer_wire buffer_11723 (.in(n11723), .out(n11723_0));
mux15 mux_6558 (.in({n14327_0, n14308_0, n14305_0, n14280_0, n14277_0, n14250_0, n14247_0, n14245_0, n14224_1, n11636_1, n8107, n8099, n8091/**/, n8003, n7995}), .out(n11724), .config_in(config_chain[22903:22898]), .config_rst(config_rst)); 
buffer_wire buffer_11724 (.in(n11724), .out(n11724_0));
mux3 mux_6559 (.in({n14811_0, n14810_0, n9073}), .out(n11725), .config_in(config_chain[22905:22904]), .config_rst(config_rst)); 
buffer_wire buffer_11725 (.in(n11725), .out(n11725_0));
mux15 mux_6560 (.in({n14329_0, n14302_0, n14299_0/**/, n14274_0, n14271_0, n14267_0, n14264_0, n14261_0, n14242_1, n11638_1, n8107, n8099, n8091, n8003, n7995}), .out(n11726), .config_in(config_chain[22911:22906]), .config_rst(config_rst)); 
buffer_wire buffer_11726 (.in(n11726), .out(n11726_0));
mux3 mux_6561 (.in({n14813_0, n14812_0, n9077}), .out(n11727), .config_in(config_chain[22913:22912]), .config_rst(config_rst)); 
buffer_wire buffer_11727 (.in(n11727), .out(n11727_0));
mux16 mux_6562 (.in({n14593_0, n14566_0, n14563_0, n14538_0, n14535_0, n14531_0, n14527_0, n14510_0, n14504_1, n14432_2, n11642_1, n9081, n9073, n8985, n8977, n8969}), .out(n11728), .config_in(config_chain[22919:22914]), .config_rst(config_rst)); 
buffer_wire buffer_11728 (.in(n11728), .out(n11728_0));
mux4 mux_6563 (.in({n14815_0, n14814_0/**/, n9085, n8969}), .out(n11729), .config_in(config_chain[22921:22920]), .config_rst(config_rst)); 
buffer_wire buffer_11729 (.in(n11729), .out(n11729_0));
mux16 mux_6564 (.in({n14575_0, n14560_0, n14557_0, n14553_0, n14549_0, n14532_0, n14524_0/**/, n14521_0, n14502_1, n14464_1, n11644_1, n9081, n9073, n8985, n8977, n8969}), .out(n11730), .config_in(config_chain[22927:22922]), .config_rst(config_rst)); 
buffer_wire buffer_11730 (.in(n11730), .out(n11730_0));
mux3 mux_6565 (.in({n14817_0, n14816_0, n8973}), .out(n11731), .config_in(config_chain[22929:22928]), .config_rst(config_rst)); 
buffer_wire buffer_11731 (.in(n11731), .out(n11731_0));
mux15 mux_6566 (.in({n14577_0, n14571_0, n14554_0/**/, n14546_0, n14543_0, n14518_0, n14515_0, n14500_1, n14486_1, n11646_1, n9081, n9073, n8985, n8977, n8969}), .out(n11732), .config_in(config_chain[22935:22930]), .config_rst(config_rst)); 
buffer_wire buffer_11732 (.in(n11732), .out(n11732_0));
mux3 mux_6567 (.in({n14819_0, n14818_0, n8977}), .out(n11733), .config_in(config_chain[22937:22936]), .config_rst(config_rst)); 
buffer_wire buffer_11733 (.in(n11733), .out(n11733_0));
mux15 mux_6568 (.in({n14579_0, n14568_0, n14565_0, n14540_0, n14537_0/**/, n14529_0, n14512_0, n14508_1, n14498_1, n11648_1, n9081, n9073, n8985, n8977, n8969}), .out(n11734), .config_in(config_chain[22943:22938]), .config_rst(config_rst)); 
buffer_wire buffer_11734 (.in(n11734), .out(n11734_0));
mux3 mux_6569 (.in({n14821_0, n14820_0, n8981}), .out(n11735), .config_in(config_chain[22945:22944]), .config_rst(config_rst)); 
buffer_wire buffer_11735 (.in(n11735), .out(n11735_0));
mux15 mux_6570 (.in({n14581_0, n14562_0, n14559_0, n14551_0, n14534_0, n14530_0, n14526_0, n14523_0, n14496_1/**/, n11650_1, n9081, n9073, n8985, n8977, n8969}), .out(n11736), .config_in(config_chain[22951:22946]), .config_rst(config_rst)); 
buffer_wire buffer_11736 (.in(n11736), .out(n11736_0));
mux3 mux_6571 (.in({n14823_0/**/, n14822_0, n8981}), .out(n11737), .config_in(config_chain[22953:22952]), .config_rst(config_rst)); 
buffer_wire buffer_11737 (.in(n11737), .out(n11737_0));
mux15 mux_6572 (.in({n14583_0, n14573_0, n14556_0, n14552_0, n14548_0, n14545_0, n14520_0, n14517_0, n14494_1, n11652_1/**/, n9085, n9077, n9069, n8981, n8973}), .out(n11738), .config_in(config_chain[22959:22954]), .config_rst(config_rst)); 
buffer_wire buffer_11738 (.in(n11738), .out(n11738_0));
mux3 mux_6573 (.in({n14825_0, n14824_0, n8985}), .out(n11739), .config_in(config_chain[22961:22960]), .config_rst(config_rst)); 
buffer_wire buffer_11739 (.in(n11739), .out(n11739_0));
mux15 mux_6574 (.in({n14585_0/**/, n14570_0, n14567_0, n14542_0, n14539_0, n14514_0, n14511_0, n14492_1, n14433_0, n11654_1, n9085, n9077, n9069, n8981, n8973}), .out(n11740), .config_in(config_chain[22967:22962]), .config_rst(config_rst)); 
buffer_wire buffer_11740 (.in(n11740), .out(n11740_0));
mux3 mux_6575 (.in({n14827_0, n14826_0, n9069}), .out(n11741), .config_in(config_chain[22969:22968]), .config_rst(config_rst)); 
buffer_wire buffer_11741 (.in(n11741), .out(n11741_0));
mux15 mux_6576 (.in({n14587_0, n14564_0/**/, n14561_0, n14536_0, n14533_0, n14528_0, n14525_0, n14490_1, n14465_0, n11656_1, n9085, n9077, n9069, n8981, n8973}), .out(n11742), .config_in(config_chain[22975:22970]), .config_rst(config_rst)); 
buffer_wire buffer_11742 (.in(n11742), .out(n11742_0));
mux3 mux_6577 (.in({n14829_0, n14828_0, n9073}), .out(n11743), .config_in(config_chain[22977:22976]), .config_rst(config_rst)); 
buffer_wire buffer_11743 (.in(n11743), .out(n11743_0));
mux15 mux_6578 (.in({n14589_0, n14558_0, n14555_0, n14550_0, n14547_0, n14522_0, n14519_0, n14488_1, n14487_0, n11658_1/**/, n9085, n9077, n9069, n8981, n8973}), .out(n11744), .config_in(config_chain[22983:22978]), .config_rst(config_rst)); 
buffer_wire buffer_11744 (.in(n11744), .out(n11744_0));
mux3 mux_6579 (.in({n14831_0, n14830_0, n9077}), .out(n11745), .config_in(config_chain[22985:22984]), .config_rst(config_rst)); 
buffer_wire buffer_11745 (.in(n11745), .out(n11745_0));
mux15 mux_6580 (.in({n14591_0/**/, n14572_0, n14569_0, n14544_0, n14541_0, n14516_0, n14513_0, n14509_0, n14506_1, n11660_1, n9085, n9077, n9069, n8981, n8973}), .out(n11746), .config_in(config_chain[22991:22986]), .config_rst(config_rst)); 
buffer_wire buffer_11746 (.in(n11746), .out(n11746_0));
mux3 mux_6581 (.in({n14833_0, n14832_0, n9077}), .out(n11747), .config_in(config_chain[22993:22992]), .config_rst(config_rst)); 
buffer_wire buffer_11747 (.in(n11747), .out(n11747_0));
mux4 mux_6582 (.in({n12503_0, n12422_1/**/, n1359, n1243}), .out(n11748), .config_in(config_chain[22995:22994]), .config_rst(config_rst)); 
buffer_wire buffer_11748 (.in(n11748), .out(n11748_0));
mux15 mux_6583 (.in({n13539_0, n13537_0, n13528_0, n13523_0, n13509_0, n13492_0, n13478_0, n13473_0, n13386_2, n11907_1, n4289, n4281, n4193, n4185, n4177}), .out(n11749), .config_in(config_chain[23001:22996]), .config_rst(config_rst)); 
buffer_wire buffer_11749 (.in(n11749), .out(n11749_0));
mux4 mux_6584 (.in({n12443_0, n12442_0/**/, n1359, n1243}), .out(n11750), .config_in(config_chain[23003:23002]), .config_rst(config_rst)); 
buffer_wire buffer_11750 (.in(n11750), .out(n11750_0));
mux15 mux_6585 (.in({n12759_0, n12742_0/**/, n12737_0, n12728_0, n12723_0, n12711_0, n12613_0, n12608_2, n12606_2, n11841_1, n1355, n1347, n1259, n1251, n1243}), .out(n11751), .config_in(config_chain[23009:23004]), .config_rst(config_rst)); 
buffer_wire buffer_11751 (.in(n11751), .out(n11751_0));
mux4 mux_6586 (.in({n12463_0, n12462_0, n1359, n1243}), .out(n11752), .config_in(config_chain[23011:23010]), .config_rst(config_rst)); 
buffer_wire buffer_11752 (.in(n11752), .out(n11752_0));
mux15 mux_6587 (.in({n13017_0, n13014_0, n13009_0, n12978_0, n12973_0/**/, n12964_0, n12959_0, n12869_0, n12864_2, n11863_1, n2333, n2325, n2237, n2229, n2221}), .out(n11753), .config_in(config_chain[23017:23012]), .config_rst(config_rst)); 
buffer_wire buffer_11753 (.in(n11753), .out(n11753_0));
mux4 mux_6588 (.in({n12483_0, n12482_0, n1359, n1243}), .out(n11754), .config_in(config_chain[23019:23018]), .config_rst(config_rst)); 
buffer_wire buffer_11754 (.in(n11754), .out(n11754_0));
mux15 mux_6589 (.in({n13277_0, n13266_0, n13261_0, n13252_0, n13247_0, n13216_0, n13211_0, n13127_0, n13124_2, n11885_1, n3311, n3303/**/, n3215, n3207, n3199}), .out(n11755), .config_in(config_chain[23025:23020]), .config_rst(config_rst)); 
buffer_wire buffer_11755 (.in(n11755), .out(n11755_0));
mux3 mux_6590 (.in({n12505_0, n12424_1, n1243}), .out(n11756), .config_in(config_chain[23027:23026]), .config_rst(config_rst)); 
buffer_wire buffer_11756 (.in(n11756), .out(n11756_0));
mux15 mux_6591 (.in({n13559_0, n13531_0, n13514_0, n13500_0, n13495_0, n13486_0, n13481_0, n13450_1, n13389_0, n11909_1, n4293, n4281, n4193, n4185, n4177}), .out(n11757), .config_in(config_chain[23033:23028]), .config_rst(config_rst)); 
buffer_wire buffer_11757 (.in(n11757), .out(n11757_0));
mux3 mux_6592 (.in({n12445_0, n12444_0, n1247}), .out(n11758), .config_in(config_chain[23035:23034]), .config_rst(config_rst)); 
buffer_wire buffer_11758 (.in(n11758), .out(n11758_0));
mux15 mux_6593 (.in({n12779_0, n12750_0/**/, n12745_0, n12731_0, n12702_0, n12697_0, n12676_1, n12615_0, n12610_2, n11843_1, n1359, n1347, n1259, n1251, n1243}), .out(n11759), .config_in(config_chain[23041:23036]), .config_rst(config_rst)); 
buffer_wire buffer_11759 (.in(n11759), .out(n11759_0));
mux3 mux_6594 (.in({n12465_0, n12464_0, n1247}), .out(n11760), .config_in(config_chain[23043:23042]), .config_rst(config_rst)); 
buffer_wire buffer_11760 (.in(n11760), .out(n11760_0));
mux15 mux_6595 (.in({n13037_0, n13000_0, n12995_0, n12986_0, n12981_0, n12967_0, n12932_1, n12871_0, n12866_2, n11865_1, n2337, n2325, n2237, n2229, n2221}), .out(n11761), .config_in(config_chain[23049:23044]), .config_rst(config_rst)); 
buffer_wire buffer_11761 (.in(n11761), .out(n11761_0));
mux3 mux_6596 (.in({n12485_0, n12484_0, n1247}), .out(n11762), .config_in(config_chain[23051:23050]), .config_rst(config_rst)); 
buffer_wire buffer_11762 (.in(n11762), .out(n11762_0));
mux15 mux_6597 (.in({n13297_0, n13274_0, n13269_0, n13238_0/**/, n13233_0, n13224_0, n13219_0, n13190_1, n13129_0, n11887_1, n3315, n3303, n3215, n3207, n3199}), .out(n11763), .config_in(config_chain[23057:23052]), .config_rst(config_rst)); 
buffer_wire buffer_11763 (.in(n11763), .out(n11763_0));
mux3 mux_6598 (.in({n12507_0, n12426_1/**/, n1247}), .out(n11764), .config_in(config_chain[23059:23058]), .config_rst(config_rst)); 
buffer_wire buffer_11764 (.in(n11764), .out(n11764_0));
mux15 mux_6599 (.in({n13557_0, n13536_0, n13522_0/**/, n13517_0, n13508_0, n13503_0, n13489_0, n13472_0, n13452_1, n11911_1, n4293, n4285, n4193, n4185, n4177}), .out(n11765), .config_in(config_chain[23065:23060]), .config_rst(config_rst)); 
buffer_wire buffer_11765 (.in(n11765), .out(n11765_0));
mux3 mux_6600 (.in({n12447_0/**/, n12446_0, n1247}), .out(n11766), .config_in(config_chain[23067:23066]), .config_rst(config_rst)); 
buffer_wire buffer_11766 (.in(n11766), .out(n11766_0));
mux15 mux_6601 (.in({n12777_0/**/, n12753_0, n12736_0, n12722_0, n12717_0, n12710_0, n12705_0, n12678_1, n12612_2, n11845_1, n1359, n1351, n1259, n1251, n1243}), .out(n11767), .config_in(config_chain[23073:23068]), .config_rst(config_rst)); 
buffer_wire buffer_11767 (.in(n11767), .out(n11767_0));
mux3 mux_6602 (.in({n12467_0, n12466_0, n1251}), .out(n11768), .config_in(config_chain[23075:23074]), .config_rst(config_rst)); 
buffer_wire buffer_11768 (.in(n11768), .out(n11768_0));
mux15 mux_6603 (.in({n13035_0, n13008_0, n13003_0, n12989_0/**/, n12972_0, n12958_0, n12953_0, n12934_1, n12868_2, n11867_1, n2337, n2329, n2237, n2229, n2221}), .out(n11769), .config_in(config_chain[23081:23076]), .config_rst(config_rst)); 
buffer_wire buffer_11769 (.in(n11769), .out(n11769_0));
mux3 mux_6604 (.in({n12487_0, n12486_0/**/, n1251}), .out(n11770), .config_in(config_chain[23083:23082]), .config_rst(config_rst)); 
buffer_wire buffer_11770 (.in(n11770), .out(n11770_0));
mux15 mux_6605 (.in({n13295_0, n13260_0, n13255_0, n13246_0, n13241_0, n13227_0, n13210_0, n13192_1, n13126_2, n11889_1, n3315, n3307, n3215/**/, n3207, n3199}), .out(n11771), .config_in(config_chain[23089:23084]), .config_rst(config_rst)); 
buffer_wire buffer_11771 (.in(n11771), .out(n11771_0));
mux3 mux_6606 (.in({n12509_0, n12428_1/**/, n1251}), .out(n11772), .config_in(config_chain[23091:23090]), .config_rst(config_rst)); 
buffer_wire buffer_11772 (.in(n11772), .out(n11772_0));
mux15 mux_6607 (.in({n13555_0, n13530_0, n13525_0, n13511_0, n13494_0, n13480_0, n13475_0, n13454_1, n13388_2, n11913_1/**/, n4293, n4285, n4277, n4185, n4177}), .out(n11773), .config_in(config_chain[23097:23092]), .config_rst(config_rst)); 
buffer_wire buffer_11773 (.in(n11773), .out(n11773_0));
mux3 mux_6608 (.in({n12449_0, n12448_0, n1251/**/}), .out(n11774), .config_in(config_chain[23099:23098]), .config_rst(config_rst)); 
buffer_wire buffer_11774 (.in(n11774), .out(n11774_0));
mux15 mux_6609 (.in({n12775_0, n12744_0, n12739_0, n12730_0, n12725_0, n12713_0, n12696_0, n12680_1, n12614_2, n11847_1, n1359, n1351, n1343, n1251, n1243}), .out(n11775), .config_in(config_chain[23105:23100]), .config_rst(config_rst)); 
buffer_wire buffer_11775 (.in(n11775), .out(n11775_0));
mux3 mux_6610 (.in({n12469_0, n12468_0, n1251/**/}), .out(n11776), .config_in(config_chain[23107:23106]), .config_rst(config_rst)); 
buffer_wire buffer_11776 (.in(n11776), .out(n11776_0));
mux15 mux_6611 (.in({n13033_0, n13011_0, n12994_0, n12980_0, n12975_0/**/, n12966_0, n12961_0, n12936_1, n12870_2, n11869_1, n2337, n2329, n2321, n2229, n2221}), .out(n11777), .config_in(config_chain[23113:23108]), .config_rst(config_rst)); 
buffer_wire buffer_11777 (.in(n11777), .out(n11777_0));
mux3 mux_6612 (.in({n12489_0, n12488_0, n1255}), .out(n11778), .config_in(config_chain[23115:23114]), .config_rst(config_rst)); 
buffer_wire buffer_11778 (.in(n11778), .out(n11778_0));
mux15 mux_6613 (.in({n13293_0, n13268_0, n13263_0, n13249_0, n13232_0, n13218_0, n13213_0, n13194_1, n13128_2, n11891_1/**/, n3315, n3307, n3299, n3207, n3199}), .out(n11779), .config_in(config_chain[23121:23116]), .config_rst(config_rst)); 
buffer_wire buffer_11779 (.in(n11779), .out(n11779_0));
mux3 mux_6614 (.in({n12511_0, n12430_1/**/, n1255}), .out(n11780), .config_in(config_chain[23123:23122]), .config_rst(config_rst)); 
buffer_wire buffer_11780 (.in(n11780), .out(n11780_0));
mux14 mux_6615 (.in({n13553_0, n13533_0, n13516_0, n13502_0, n13497_0, n13488_0, n13483_0, n13456_1, n11915_1, n4293, n4285, n4277, n4189, n4177}), .out(n11781), .config_in(config_chain[23129:23124]), .config_rst(config_rst)); 
buffer_wire buffer_11781 (.in(n11781), .out(n11781_0));
mux3 mux_6616 (.in({n12451_0, n12450_0, n1255}), .out(n11782), .config_in(config_chain[23131:23130]), .config_rst(config_rst)); 
buffer_wire buffer_11782 (.in(n11782), .out(n11782_0));
mux14 mux_6617 (.in({n12773_0, n12752_0, n12747_0, n12733_0, n12716_0, n12704_0, n12699_0, n12682_1, n11849_1, n1359, n1351, n1343, n1255, n1243}), .out(n11783), .config_in(config_chain[23137:23132]), .config_rst(config_rst)); 
buffer_wire buffer_11783 (.in(n11783), .out(n11783_0));
mux3 mux_6618 (.in({n12471_0, n12470_0, n1255}), .out(n11784), .config_in(config_chain[23139:23138]), .config_rst(config_rst)); 
buffer_wire buffer_11784 (.in(n11784), .out(n11784_0));
mux14 mux_6619 (.in({n13031_0, n13002_0, n12997_0, n12988_0, n12983_0, n12969_0, n12952_0, n12938_1, n11871_1, n2337, n2329, n2321, n2233, n2221}), .out(n11785), .config_in(config_chain[23145:23140]), .config_rst(config_rst)); 
buffer_wire buffer_11785 (.in(n11785), .out(n11785_0));
mux3 mux_6620 (.in({n12491_0, n12490_0, n1255}), .out(n11786), .config_in(config_chain[23147:23146]), .config_rst(config_rst)); 
buffer_wire buffer_11786 (.in(n11786), .out(n11786_0));
mux14 mux_6621 (.in({n13291_0, n13271_0, n13254_0/**/, n13240_0, n13235_0, n13226_0, n13221_0, n13196_1, n11893_1, n3315, n3307, n3299, n3211, n3199}), .out(n11787), .config_in(config_chain[23153:23148]), .config_rst(config_rst)); 
buffer_wire buffer_11787 (.in(n11787), .out(n11787_0));
mux3 mux_6622 (.in({n12513_0, n12432_1/**/, n1259}), .out(n11788), .config_in(config_chain[23155:23154]), .config_rst(config_rst)); 
buffer_wire buffer_11788 (.in(n11788), .out(n11788_0));
mux14 mux_6623 (.in({n13551_0, n13524_0, n13519_0, n13510_0, n13505_0, n13491_0, n13474_0, n13458_1, n11917_1, n4293/**/, n4285, n4277, n4189, n4181}), .out(n11789), .config_in(config_chain[23161:23156]), .config_rst(config_rst)); 
buffer_wire buffer_11789 (.in(n11789), .out(n11789_0));
mux3 mux_6624 (.in({n12453_0, n12452_0, n1259}), .out(n11790), .config_in(config_chain[23163:23162]), .config_rst(config_rst)); 
buffer_wire buffer_11790 (.in(n11790), .out(n11790_0));
mux14 mux_6625 (.in({n12771_0, n12755_0, n12738_0, n12724_0, n12719_0, n12712_0, n12707_0, n12684_1, n11851_1, n1359, n1351, n1343, n1255/**/, n1247}), .out(n11791), .config_in(config_chain[23169:23164]), .config_rst(config_rst)); 
buffer_wire buffer_11791 (.in(n11791), .out(n11791_0));
mux3 mux_6626 (.in({n12473_0, n12472_0, n1259}), .out(n11792), .config_in(config_chain[23171:23170]), .config_rst(config_rst)); 
buffer_wire buffer_11792 (.in(n11792), .out(n11792_0));
mux14 mux_6627 (.in({n13029_0, n13010_0, n13005_0, n12991_0, n12974_0, n12960_0, n12955_0, n12940_1, n11873_1/**/, n2337, n2329, n2321, n2233, n2225}), .out(n11793), .config_in(config_chain[23177:23172]), .config_rst(config_rst)); 
buffer_wire buffer_11793 (.in(n11793), .out(n11793_0));
mux3 mux_6628 (.in({n12493_0, n12492_0/**/, n1259}), .out(n11794), .config_in(config_chain[23179:23178]), .config_rst(config_rst)); 
buffer_wire buffer_11794 (.in(n11794), .out(n11794_0));
mux14 mux_6629 (.in({n13289_0, n13262_0/**/, n13257_0, n13248_0, n13243_0, n13229_0, n13212_0, n13198_1, n11895_1, n3315, n3307, n3299, n3211, n3203}), .out(n11795), .config_in(config_chain[23185:23180]), .config_rst(config_rst)); 
buffer_wire buffer_11795 (.in(n11795), .out(n11795_0));
mux3 mux_6630 (.in({n12515_0, n12434_1/**/, n1259}), .out(n11796), .config_in(config_chain[23187:23186]), .config_rst(config_rst)); 
buffer_wire buffer_11796 (.in(n11796), .out(n11796_0));
mux13 mux_6631 (.in({n13549_0, n13532_0, n13527_0, n13513_0, n13496_0, n13482_0/**/, n13477_0, n13460_1, n11919_1, n4285, n4277, n4189, n4181}), .out(n11797), .config_in(config_chain[23193:23188]), .config_rst(config_rst)); 
buffer_wire buffer_11797 (.in(n11797), .out(n11797_0));
mux3 mux_6632 (.in({n12455_0, n12454_0, n1343}), .out(n11798), .config_in(config_chain[23195:23194]), .config_rst(config_rst)); 
buffer_wire buffer_11798 (.in(n11798), .out(n11798_0));
mux13 mux_6633 (.in({n12769_0, n12746_0, n12741_0, n12732_0, n12727_0, n12715_0, n12698_0, n12686_1, n11853_1, n1351, n1343, n1255, n1247}), .out(n11799), .config_in(config_chain[23201:23196]), .config_rst(config_rst)); 
buffer_wire buffer_11799 (.in(n11799), .out(n11799_0));
mux3 mux_6634 (.in({n12475_0, n12474_0, n1343}), .out(n11800), .config_in(config_chain[23203:23202]), .config_rst(config_rst)); 
buffer_wire buffer_11800 (.in(n11800), .out(n11800_0));
mux13 mux_6635 (.in({n13027_0, n13013_0, n12996_0/**/, n12982_0, n12977_0, n12968_0, n12963_0, n12942_1, n11875_1, n2329, n2321, n2233, n2225}), .out(n11801), .config_in(config_chain[23209:23204]), .config_rst(config_rst)); 
buffer_wire buffer_11801 (.in(n11801), .out(n11801_0));
mux3 mux_6636 (.in({n12495_0, n12494_0, n1343}), .out(n11802), .config_in(config_chain[23211:23210]), .config_rst(config_rst)); 
buffer_wire buffer_11802 (.in(n11802), .out(n11802_0));
mux13 mux_6637 (.in({n13287_0/**/, n13270_0, n13265_0, n13251_0, n13234_0, n13220_0, n13215_0, n13200_1, n11897_1, n3307, n3299, n3211, n3203}), .out(n11803), .config_in(config_chain[23217:23212]), .config_rst(config_rst)); 
buffer_wire buffer_11803 (.in(n11803), .out(n11803_0));
mux3 mux_6638 (.in({n12517_0/**/, n12436_1, n1343}), .out(n11804), .config_in(config_chain[23219:23218]), .config_rst(config_rst)); 
buffer_wire buffer_11804 (.in(n11804), .out(n11804_0));
mux13 mux_6639 (.in({n13547_0/**/, n13535_0, n13518_0, n13504_0, n13499_0, n13490_0, n13485_0, n13462_1, n11921_1, n4289, n4277, n4189, n4181}), .out(n11805), .config_in(config_chain[23225:23220]), .config_rst(config_rst)); 
buffer_wire buffer_11805 (.in(n11805), .out(n11805_0));
mux3 mux_6640 (.in({n12457_0, n12456_0, n1343}), .out(n11806), .config_in(config_chain[23227:23226]), .config_rst(config_rst)); 
buffer_wire buffer_11806 (.in(n11806), .out(n11806_0));
mux13 mux_6641 (.in({n12767_0, n12754_0, n12749_0, n12735_0, n12718_0, n12706_0, n12701_0, n12688_1, n11855_1, n1355, n1343, n1255, n1247}), .out(n11807), .config_in(config_chain[23233:23228]), .config_rst(config_rst)); 
buffer_wire buffer_11807 (.in(n11807), .out(n11807_0));
mux3 mux_6642 (.in({n12477_0, n12476_0, n1347}), .out(n11808), .config_in(config_chain[23235:23234]), .config_rst(config_rst)); 
buffer_wire buffer_11808 (.in(n11808), .out(n11808_0));
mux13 mux_6643 (.in({n13025_0/**/, n13004_0, n12999_0, n12990_0, n12985_0, n12971_0, n12954_0, n12944_1, n11877_1, n2333, n2321, n2233, n2225}), .out(n11809), .config_in(config_chain[23241:23236]), .config_rst(config_rst)); 
buffer_wire buffer_11809 (.in(n11809), .out(n11809_0));
mux3 mux_6644 (.in({n12497_0, n12496_0, n1347}), .out(n11810), .config_in(config_chain[23243:23242]), .config_rst(config_rst)); 
buffer_wire buffer_11810 (.in(n11810), .out(n11810_0));
mux13 mux_6645 (.in({n13285_0, n13273_0, n13256_0, n13242_0, n13237_0, n13228_0, n13223_0, n13202_1/**/, n11899_1, n3311, n3299, n3211, n3203}), .out(n11811), .config_in(config_chain[23249:23244]), .config_rst(config_rst)); 
buffer_wire buffer_11811 (.in(n11811), .out(n11811_0));
mux3 mux_6646 (.in({n12519_0, n12438_1/**/, n1347}), .out(n11812), .config_in(config_chain[23251:23250]), .config_rst(config_rst)); 
buffer_wire buffer_11812 (.in(n11812), .out(n11812_0));
mux13 mux_6647 (.in({n13545_0, n13526_0, n13521_0/**/, n13512_0, n13507_0, n13476_0, n13471_0, n13464_1, n11923_1, n4289, n4281, n4189, n4181}), .out(n11813), .config_in(config_chain[23257:23252]), .config_rst(config_rst)); 
buffer_wire buffer_11813 (.in(n11813), .out(n11813_0));
mux3 mux_6648 (.in({n12459_0, n12458_0, n1347}), .out(n11814), .config_in(config_chain[23259:23258]), .config_rst(config_rst)); 
buffer_wire buffer_11814 (.in(n11814), .out(n11814_0));
mux13 mux_6649 (.in({n12765_0, n12757_0, n12740_0, n12726_0, n12721_0, n12714_0/**/, n12709_0, n12690_1, n11857_1, n1355, n1347, n1255, n1247}), .out(n11815), .config_in(config_chain[23265:23260]), .config_rst(config_rst)); 
buffer_wire buffer_11815 (.in(n11815), .out(n11815_0));
mux3 mux_6650 (.in({n12479_0, n12478_0, n1347}), .out(n11816), .config_in(config_chain[23267:23266]), .config_rst(config_rst)); 
buffer_wire buffer_11816 (.in(n11816), .out(n11816_0));
mux13 mux_6651 (.in({n13023_0, n13012_0/**/, n13007_0, n12993_0, n12976_0, n12962_0, n12957_0, n12946_1, n11879_1, n2333, n2325, n2233, n2225}), .out(n11817), .config_in(config_chain[23273:23268]), .config_rst(config_rst)); 
buffer_wire buffer_11817 (.in(n11817), .out(n11817_0));
mux3 mux_6652 (.in({n12499_0, n12498_0, n1351}), .out(n11818), .config_in(config_chain[23275:23274]), .config_rst(config_rst)); 
buffer_wire buffer_11818 (.in(n11818), .out(n11818_0));
mux13 mux_6653 (.in({n13283_0/**/, n13264_0, n13259_0, n13250_0, n13245_0, n13231_0, n13214_0, n13204_1, n11901_1, n3311, n3303, n3211, n3203}), .out(n11819), .config_in(config_chain[23281:23276]), .config_rst(config_rst)); 
buffer_wire buffer_11819 (.in(n11819), .out(n11819_0));
mux3 mux_6654 (.in({n12521_0, n12440_1/**/, n1351}), .out(n11820), .config_in(config_chain[23283:23282]), .config_rst(config_rst)); 
buffer_wire buffer_11820 (.in(n11820), .out(n11820_0));
mux13 mux_6655 (.in({n13543_0, n13534_0, n13529_0/**/, n13498_0, n13493_0, n13484_0, n13479_0, n13466_1, n11925_1, n4289, n4281, n4193, n4181}), .out(n11821), .config_in(config_chain[23289:23284]), .config_rst(config_rst)); 
buffer_wire buffer_11821 (.in(n11821), .out(n11821_0));
mux3 mux_6656 (.in({n12461_0, n12460_0, n1351}), .out(n11822), .config_in(config_chain[23291:23290]), .config_rst(config_rst)); 
buffer_wire buffer_11822 (.in(n11822), .out(n11822_0));
mux13 mux_6657 (.in({n12763_0, n12748_0, n12743_0, n12734_0, n12729_0, n12700_0, n12692_1/**/, n12609_0, n11859_1, n1355, n1347, n1259, n1247}), .out(n11823), .config_in(config_chain[23297:23292]), .config_rst(config_rst)); 
buffer_wire buffer_11823 (.in(n11823), .out(n11823_0));
mux3 mux_6658 (.in({n12481_0/**/, n12480_0, n1351}), .out(n11824), .config_in(config_chain[23299:23298]), .config_rst(config_rst)); 
buffer_wire buffer_11824 (.in(n11824), .out(n11824_0));
mux13 mux_6659 (.in({n13021_0, n13015_0, n12998_0, n12984_0, n12979_0, n12970_0, n12965_0, n12948_1, n11881_1, n2333, n2325, n2237, n2225}), .out(n11825), .config_in(config_chain[23305:23300]), .config_rst(config_rst)); 
buffer_wire buffer_11825 (.in(n11825), .out(n11825_0));
mux3 mux_6660 (.in({n12501_0, n12500_0, n1351}), .out(n11826), .config_in(config_chain[23307:23306]), .config_rst(config_rst)); 
buffer_wire buffer_11826 (.in(n11826), .out(n11826_0));
mux13 mux_6661 (.in({n13281_0/**/, n13272_0, n13267_0, n13253_0, n13236_0, n13222_0, n13217_0, n13206_1, n11903_1, n3311, n3303, n3215, n3203}), .out(n11827), .config_in(config_chain[23313:23308]), .config_rst(config_rst)); 
buffer_wire buffer_11827 (.in(n11827), .out(n11827_0));
mux3 mux_6662 (.in({n12523_0, n12350_2, n1355}), .out(n11828), .config_in(config_chain[23315:23314]), .config_rst(config_rst)); 
buffer_wire buffer_11828 (.in(n11828), .out(n11828_0));
mux3 mux_6663 (.in({n14695_0, n14694_2, n9179}), .out(n11829), .config_in(config_chain[23317:23316]), .config_rst(config_rst)); 
buffer_wire buffer_11829 (.in(n11829), .out(n11829_0));
mux3 mux_6664 (.in({n12353_0, n12352_2, n1355}), .out(n11830), .config_in(config_chain[23319:23318]), .config_rst(config_rst)); 
buffer_wire buffer_11830 (.in(n11830), .out(n11830_0));
mux13 mux_6665 (.in({n12761_0, n12756_0, n12751_0, n12720_0, n12708_0, n12703_0, n12694_1, n12611_0, n11861_2, n1355, n1347, n1259, n1251/**/}), .out(n11831), .config_in(config_chain[23325:23320]), .config_rst(config_rst)); 
buffer_wire buffer_11831 (.in(n11831), .out(n11831_0));
mux3 mux_6666 (.in({n12355_0, n12354_2, n1355}), .out(n11832), .config_in(config_chain[23327:23326]), .config_rst(config_rst)); 
buffer_wire buffer_11832 (.in(n11832), .out(n11832_0));
mux13 mux_6667 (.in({n13019_0, n13006_0, n13001_0, n12992_0, n12987_0, n12956_0, n12950_1, n12867_0, n11883_2, n2333, n2325/**/, n2237, n2229}), .out(n11833), .config_in(config_chain[23333:23328]), .config_rst(config_rst)); 
buffer_wire buffer_11833 (.in(n11833), .out(n11833_0));
mux3 mux_6668 (.in({n12357_0, n12356_2, n1355}), .out(n11834), .config_in(config_chain[23335:23334]), .config_rst(config_rst)); 
buffer_wire buffer_11834 (.in(n11834), .out(n11834_0));
mux13 mux_6669 (.in({n13279_0, n13275_0, n13258_0, n13244_0, n13239_0, n13230_0, n13225_0, n13208_1, n11905_1, n3311, n3303, n3215, n3207}), .out(n11835), .config_in(config_chain[23341:23336]), .config_rst(config_rst)); 
buffer_wire buffer_11835 (.in(n11835), .out(n11835_0));
mux3 mux_6670 (.in({n12359_0, n12358_2, n1355}), .out(n11836), .config_in(config_chain[23343:23342]), .config_rst(config_rst)); 
buffer_wire buffer_11836 (.in(n11836), .out(n11836_0));
mux13 mux_6671 (.in({n13541_0, n13520_0, n13515_0, n13506_0, n13501_0, n13487_0, n13470_1, n13468_1, n11927_1, n4289, n4281, n4193, n4185}), .out(n11837), .config_in(config_chain[23349:23344]), .config_rst(config_rst)); 
buffer_wire buffer_11837 (.in(n11837), .out(n11837_0));
mux3 mux_6672 (.in({n12361_0, n12360_2, n1359}), .out(n11838), .config_in(config_chain[23351:23350]), .config_rst(config_rst)); 
buffer_wire buffer_11838 (.in(n11838), .out(n11838_0));
mux13 mux_6673 (.in({n13805_0, n13795_0, n13762_0, n13757_0, n13748_0, n13743_0, n13732_1, n13712_1, n11949_1/**/, n5267, n5259, n5171, n5163}), .out(n11839), .config_in(config_chain[23357:23352]), .config_rst(config_rst)); 
buffer_wire buffer_11839 (.in(n11839), .out(n11839_0));
mux15 mux_6674 (.in({n12779_0, n12743_0, n12736_0/**/, n12729_0, n12722_0, n12710_0, n12694_1, n12612_2, n12609_0, n11750_0, n2333, n2325, n2237, n2229, n2221}), .out(n11840), .config_in(config_chain[23363:23358]), .config_rst(config_rst)); 
buffer_wire buffer_11840 (.in(n11840), .out(n11840_0));
mux15 mux_6675 (.in({n13803_0, n13786_0, n13781_0, n13779_0, n13770_0, n13765_0, n13751_0/**/, n13734_1, n13650_2, n11929_1, n5267, n5259, n5171, n5163, n5155}), .out(n11841), .config_in(config_chain[23369:23364]), .config_rst(config_rst)); 
buffer_wire buffer_11841 (.in(n11841), .out(n11841_0));
mux15 mux_6676 (.in({n12759_0, n12751_0, n12744_0, n12730_0, n12703_0, n12696_0/**/, n12692_1, n12614_2, n12611_0, n11758_0, n2337, n2325, n2237, n2229, n2221}), .out(n11842), .config_in(config_chain[23375:23370]), .config_rst(config_rst)); 
buffer_wire buffer_11842 (.in(n11842), .out(n11842_0));
mux15 mux_6677 (.in({n13823_0, n13801_0, n13794_0, n13789_0, n13773_0, n13756_0, n13742_0, n13737_0, n13714_1, n11931_1, n5271, n5259/**/, n5171, n5163, n5155}), .out(n11843), .config_in(config_chain[23381:23376]), .config_rst(config_rst)); 
buffer_wire buffer_11843 (.in(n11843), .out(n11843_0));
mux15 mux_6678 (.in({n12761_0, n12752_0, n12737_0/**/, n12723_0, n12716_0, n12711_0, n12704_0, n12690_1, n12613_0, n11766_0, n2337, n2329, n2237, n2229, n2221}), .out(n11844), .config_in(config_chain[23387:23382]), .config_rst(config_rst)); 
buffer_wire buffer_11844 (.in(n11844), .out(n11844_0));
mux15 mux_6679 (.in({n13821_0, n13797_0, n13780_0, n13778_0, n13764_0, n13759_0, n13750_0, n13745_0, n13716_1, n11933_1, n5271, n5263, n5171, n5163, n5155}), .out(n11845), .config_in(config_chain[23393:23388]), .config_rst(config_rst)); 
buffer_wire buffer_11845 (.in(n11845), .out(n11845_0));
mux15 mux_6680 (.in({n12763_0, n12745_0, n12738_0, n12731_0, n12724_0, n12712_0, n12697_0, n12688_1, n12615_0, n11774_0/**/, n2337, n2329, n2321, n2229, n2221}), .out(n11846), .config_in(config_chain[23399:23394]), .config_rst(config_rst)); 
buffer_wire buffer_11846 (.in(n11846), .out(n11846_0));
mux15 mux_6681 (.in({n13819_0, n13800_0, n13788_0, n13783_0, n13772_0, n13767_0, n13753_0/**/, n13736_0, n13718_1, n11935_1, n5271, n5263, n5255, n5163, n5155}), .out(n11847), .config_in(config_chain[23405:23400]), .config_rst(config_rst)); 
buffer_wire buffer_11847 (.in(n11847), .out(n11847_0));
mux14 mux_6682 (.in({n12765_0, n12753_0, n12746_0, n12732_0, n12717_0, n12705_0, n12698_0, n12686_1, n11782_0, n2337, n2329/**/, n2321, n2233, n2221}), .out(n11848), .config_in(config_chain[23411:23406]), .config_rst(config_rst)); 
buffer_wire buffer_11848 (.in(n11848), .out(n11848_0));
mux14 mux_6683 (.in({n13817_0, n13796_0/**/, n13791_0, n13775_0, n13758_0, n13744_0, n13739_0, n13720_1, n11937_1, n5271, n5263, n5255, n5167, n5155}), .out(n11849), .config_in(config_chain[23417:23412]), .config_rst(config_rst)); 
buffer_wire buffer_11849 (.in(n11849), .out(n11849_0));
mux14 mux_6684 (.in({n12767_0, n12754_0, n12739_0, n12725_0, n12718_0, n12713_0, n12706_0, n12684_1/**/, n11790_0, n2337, n2329, n2321, n2233, n2225}), .out(n11850), .config_in(config_chain[23423:23418]), .config_rst(config_rst)); 
buffer_wire buffer_11850 (.in(n11850), .out(n11850_0));
mux14 mux_6685 (.in({n13815_0, n13799_0, n13782_0, n13766_0, n13761_0, n13752_0, n13747_0, n13722_1, n11939_1, n5271, n5263, n5255, n5167, n5159}), .out(n11851), .config_in(config_chain[23429:23424]), .config_rst(config_rst)); 
buffer_wire buffer_11851 (.in(n11851), .out(n11851_0));
mux13 mux_6686 (.in({n12769_0, n12747_0, n12740_0/**/, n12733_0, n12726_0, n12714_0, n12699_0, n12682_1, n11798_0, n2329, n2321, n2233, n2225}), .out(n11852), .config_in(config_chain[23435:23430]), .config_rst(config_rst)); 
buffer_wire buffer_11852 (.in(n11852), .out(n11852_0));
mux13 mux_6687 (.in({n13813_0, n13790_0, n13785_0, n13774_0, n13769_0, n13755_0, n13738_0, n13724_1/**/, n11941_1, n5263, n5255, n5167, n5159}), .out(n11853), .config_in(config_chain[23441:23436]), .config_rst(config_rst)); 
buffer_wire buffer_11853 (.in(n11853), .out(n11853_0));
mux13 mux_6688 (.in({n12771_0, n12755_0, n12748_0, n12734_0, n12719_0, n12707_0, n12700_0, n12680_1, n11806_0, n2333, n2321, n2233, n2225/**/}), .out(n11854), .config_in(config_chain[23447:23442]), .config_rst(config_rst)); 
buffer_wire buffer_11854 (.in(n11854), .out(n11854_0));
mux13 mux_6689 (.in({n13811_0, n13798_0, n13793_0, n13777_0, n13760_0, n13746_0/**/, n13741_0, n13726_1, n11943_1, n5267, n5255, n5167, n5159}), .out(n11855), .config_in(config_chain[23453:23448]), .config_rst(config_rst)); 
buffer_wire buffer_11855 (.in(n11855), .out(n11855_0));
mux13 mux_6690 (.in({n12773_0/**/, n12756_0, n12741_0, n12727_0, n12720_0, n12715_0, n12708_0, n12678_1, n11814_0, n2333, n2325, n2233, n2225}), .out(n11856), .config_in(config_chain[23459:23454]), .config_rst(config_rst)); 
buffer_wire buffer_11856 (.in(n11856), .out(n11856_0));
mux13 mux_6691 (.in({n13809_0, n13784_0, n13768_0, n13763_0, n13754_0, n13749_0, n13728_1, n13713_0, n11945_1/**/, n5267, n5259, n5167, n5159}), .out(n11857), .config_in(config_chain[23465:23460]), .config_rst(config_rst)); 
buffer_wire buffer_11857 (.in(n11857), .out(n11857_0));
mux13 mux_6692 (.in({n12775_0, n12749_0, n12742_0, n12735_0, n12728_0, n12701_0, n12676_1, n12608_2, n11822_0, n2333, n2325, n2237, n2225/**/}), .out(n11858), .config_in(config_chain[23471:23466]), .config_rst(config_rst)); 
buffer_wire buffer_11858 (.in(n11858), .out(n11858_0));
mux13 mux_6693 (.in({n13807_0, n13792_0, n13787_0, n13776_0, n13771_0, n13740_0, n13735_0, n13730_1, n11947_1/**/, n5267, n5259, n5171, n5159}), .out(n11859), .config_in(config_chain[23477:23472]), .config_rst(config_rst)); 
buffer_wire buffer_11859 (.in(n11859), .out(n11859_0));
mux13 mux_6694 (.in({n12777_0, n12757_0, n12750_0, n12721_0, n12709_0, n12702_0, n12610_2, n12606_2, n11830_0, n2333, n2325/**/, n2237, n2229}), .out(n11860), .config_in(config_chain[23483:23478]), .config_rst(config_rst)); 
buffer_wire buffer_11860 (.in(n11860), .out(n11860_0));
mux3 mux_6695 (.in({n14697_0, n14696_2, n9179}), .out(n11861), .config_in(config_chain[23485:23484]), .config_rst(config_rst)); 
buffer_wire buffer_11861 (.in(n11861), .out(n11861_0));
mux15 mux_6696 (.in({n13037_0, n13015_0, n13008_0/**/, n12979_0, n12972_0, n12965_0, n12958_0, n12950_1, n12868_2, n11752_0, n3311, n3303, n3215, n3207, n3199}), .out(n11862), .config_in(config_chain[23491:23486]), .config_rst(config_rst)); 
buffer_wire buffer_11862 (.in(n11862), .out(n11862_0));
mux16 mux_6697 (.in({n14069_0, n14053_0, n14048_0, n14044_0, n14040_0, n14025_0, n14015_0, n14010_0, n13998_1/**/, n13957_0, n11951_0, n6245, n6237, n6149, n6141, n6133}), .out(n11863), .config_in(config_chain[23497:23492]), .config_rst(config_rst)); 
buffer_wire buffer_11863 (.in(n11863), .out(n11863_0));
mux15 mux_6698 (.in({n13017_0, n13001_0, n12994_0/**/, n12987_0, n12980_0, n12966_0, n12948_1, n12870_2, n12867_0, n11760_0, n3315, n3303, n3215, n3207, n3199}), .out(n11864), .config_in(config_chain[23503:23498]), .config_rst(config_rst)); 
buffer_wire buffer_11864 (.in(n11864), .out(n11864_0));
mux16 mux_6699 (.in({n14087_0, n14066_0, n14062_0, n14047_0, n14039_0, n14034_0, n14009_0, n14004_0, n13980_1, n13979_0, n11953_0, n6245, n6237, n6149/**/, n6141, n6133}), .out(n11865), .config_in(config_chain[23509:23504]), .config_rst(config_rst)); 
buffer_wire buffer_11865 (.in(n11865), .out(n11865_0));
mux15 mux_6700 (.in({n13019_0, n13009_0, n13002_0, n12988_0, n12973_0, n12959_0, n12952_0, n12946_1, n12869_0, n11768_0, n3315/**/, n3307, n3215, n3207, n3199}), .out(n11866), .config_in(config_chain[23515:23510]), .config_rst(config_rst)); 
buffer_wire buffer_11866 (.in(n11866), .out(n11866_0));
mux15 mux_6701 (.in({n14085_0, n14061_0, n14056_0/**/, n14033_0, n14028_0, n14018_0, n14003_0, n14001_0, n13982_1, n11955_0, n6245, n6237, n6149, n6141, n6133}), .out(n11867), .config_in(config_chain[23521:23516]), .config_rst(config_rst)); 
buffer_wire buffer_11867 (.in(n11867), .out(n11867_0));
mux15 mux_6702 (.in({n13021_0, n13010_0, n12995_0, n12981_0, n12974_0, n12967_0, n12960_0, n12944_1, n12871_0, n11776_0/**/, n3315, n3307, n3299, n3207, n3199}), .out(n11868), .config_in(config_chain[23527:23522]), .config_rst(config_rst)); 
buffer_wire buffer_11868 (.in(n11868), .out(n11868_0));
mux15 mux_6703 (.in({n14083_0, n14055_0, n14050_0, n14042_0, n14027_0, n14023_0, n14017_0, n14012_0/**/, n13984_1, n11957_0, n6245, n6237, n6149, n6141, n6133}), .out(n11869), .config_in(config_chain[23533:23528]), .config_rst(config_rst)); 
buffer_wire buffer_11869 (.in(n11869), .out(n11869_0));
mux14 mux_6704 (.in({n13023_0, n13003_0, n12996_0, n12989_0, n12982_0, n12968_0/**/, n12953_0, n12942_1, n11784_0, n3315, n3307, n3299, n3211, n3199}), .out(n11870), .config_in(config_chain[23539:23534]), .config_rst(config_rst)); 
buffer_wire buffer_11870 (.in(n11870), .out(n11870_0));
mux15 mux_6705 (.in({n14081_0, n14064_0, n14049_0, n14045_0, n14041_0/**/, n14036_0, n14011_0, n14006_0, n13986_1, n11959_0, n6245, n6237, n6149, n6141, n6133}), .out(n11871), .config_in(config_chain[23545:23540]), .config_rst(config_rst)); 
buffer_wire buffer_11871 (.in(n11871), .out(n11871_0));
mux14 mux_6706 (.in({n13025_0, n13011_0, n13004_0, n12990_0, n12975_0, n12961_0, n12954_0, n12940_1, n11792_0, n3315, n3307/**/, n3299, n3211, n3203}), .out(n11872), .config_in(config_chain[23551:23546]), .config_rst(config_rst)); 
buffer_wire buffer_11872 (.in(n11872), .out(n11872_0));
mux15 mux_6707 (.in({n14079_0, n14067_0, n14063_0, n14058_0, n14035_0, n14030_0, n14020_0, n14005_0, n13988_1, n11961_0, n6249, n6241, n6233, n6145, n6137/**/}), .out(n11873), .config_in(config_chain[23557:23552]), .config_rst(config_rst)); 
buffer_wire buffer_11873 (.in(n11873), .out(n11873_0));
mux13 mux_6708 (.in({n13027_0, n13012_0/**/, n12997_0, n12983_0, n12976_0, n12969_0, n12962_0, n12938_1, n11800_0, n3307, n3299, n3211, n3203}), .out(n11874), .config_in(config_chain[23563:23558]), .config_rst(config_rst)); 
buffer_wire buffer_11874 (.in(n11874), .out(n11874_0));
mux15 mux_6709 (.in({n14077_0, n14057_0, n14052_0, n14029_0/**/, n14024_0, n14019_0, n14014_0, n13990_1, n13956_1, n11963_0, n6249, n6241, n6233, n6145, n6137}), .out(n11875), .config_in(config_chain[23569:23564]), .config_rst(config_rst)); 
buffer_wire buffer_11875 (.in(n11875), .out(n11875_0));
mux13 mux_6710 (.in({n13029_0, n13005_0, n12998_0/**/, n12991_0, n12984_0, n12970_0, n12955_0, n12936_1, n11808_0, n3311, n3299, n3211, n3203}), .out(n11876), .config_in(config_chain[23575:23570]), .config_rst(config_rst)); 
buffer_wire buffer_11876 (.in(n11876), .out(n11876_0));
mux15 mux_6711 (.in({n14075_0, n14051_0, n14046_0, n14043_0, n14038_0, n14013_0, n14008_0, n13992_1/**/, n13978_1, n11965_0, n6249, n6241, n6233, n6145, n6137}), .out(n11877), .config_in(config_chain[23581:23576]), .config_rst(config_rst)); 
buffer_wire buffer_11877 (.in(n11877), .out(n11877_0));
mux13 mux_6712 (.in({n13031_0, n13013_0, n13006_0/**/, n12992_0, n12977_0, n12963_0, n12956_0, n12934_1, n11816_0, n3311, n3303, n3211, n3203}), .out(n11878), .config_in(config_chain[23587:23582]), .config_rst(config_rst)); 
buffer_wire buffer_11878 (.in(n11878), .out(n11878_0));
mux15 mux_6713 (.in({n14073_0, n14065_0/**/, n14060_0, n14037_0, n14032_0, n14007_0, n14002_0, n14000_1, n13994_1, n11967_0, n6249, n6241, n6233, n6145, n6137}), .out(n11879), .config_in(config_chain[23593:23588]), .config_rst(config_rst)); 
buffer_wire buffer_11879 (.in(n11879), .out(n11879_0));
mux13 mux_6714 (.in({n13033_0, n13014_0, n12999_0, n12985_0, n12978_0, n12971_0, n12964_0, n12932_1/**/, n11824_0, n3311, n3303, n3215, n3203}), .out(n11880), .config_in(config_chain[23599:23594]), .config_rst(config_rst)); 
buffer_wire buffer_11880 (.in(n11880), .out(n11880_0));
mux15 mux_6715 (.in({n14071_0, n14059_0, n14054_0, n14031_0, n14026_0, n14022_0, n14021_0, n14016_0, n13996_1, n11969_0, n6249, n6241, n6233, n6145, n6137}), .out(n11881), .config_in(config_chain[23605:23600]), .config_rst(config_rst)); 
buffer_wire buffer_11881 (.in(n11881), .out(n11881_0));
mux13 mux_6716 (.in({n13035_0, n13007_0, n13000_0, n12993_0, n12986_0, n12957_0, n12866_2, n12864_2, n11832_0, n3311, n3303/**/, n3215, n3207}), .out(n11882), .config_in(config_chain[23611:23606]), .config_rst(config_rst)); 
buffer_wire buffer_11882 (.in(n11882), .out(n11882_0));
mux3 mux_6717 (.in({n14727_0, n14726_2/**/, n9179}), .out(n11883), .config_in(config_chain[23613:23612]), .config_rst(config_rst)); 
buffer_wire buffer_11883 (.in(n11883), .out(n11883_0));
mux15 mux_6718 (.in({n13297_0, n13267_0, n13260_0, n13253_0, n13246_0, n13217_0, n13210_0, n13208_1, n13126_2, n11754_0, n4289/**/, n4281, n4193, n4185, n4177}), .out(n11884), .config_in(config_chain[23619:23614]), .config_rst(config_rst)); 
buffer_wire buffer_11884 (.in(n11884), .out(n11884_0));
mux16 mux_6719 (.in({n14333_0, n14325_0, n14320_0, n14297_0, n14292_0, n14288_0, n14284_0, n14269_0, n14264_1, n14201_0, n11971_0, n7223, n7215, n7127, n7119/**/, n7111}), .out(n11885), .config_in(config_chain[23625:23620]), .config_rst(config_rst)); 
buffer_wire buffer_11885 (.in(n11885), .out(n11885_0));
mux15 mux_6720 (.in({n13277_0, n13275_0/**/, n13268_0, n13239_0, n13232_0, n13225_0, n13218_0, n13206_1, n13128_2, n11762_0, n4293, n4281, n4193, n4185, n4177}), .out(n11886), .config_in(config_chain[23631:23626]), .config_rst(config_rst)); 
buffer_wire buffer_11886 (.in(n11886), .out(n11886_0));
mux16 mux_6721 (.in({n14351_0, n14319_0, n14314_0, n14310_0, n14306_0/**/, n14291_0, n14283_0, n14278_0, n14246_1, n14223_0, n11973_0, n7223, n7215, n7127, n7119, n7111}), .out(n11887), .config_in(config_chain[23637:23632]), .config_rst(config_rst)); 
buffer_wire buffer_11887 (.in(n11887), .out(n11887_0));
mux15 mux_6722 (.in({n13279_0/**/, n13261_0, n13254_0, n13247_0, n13240_0, n13226_0, n13211_0, n13204_1, n13127_0, n11770_0, n4293, n4285, n4193, n4185, n4177}), .out(n11888), .config_in(config_chain[23643:23638]), .config_rst(config_rst)); 
buffer_wire buffer_11888 (.in(n11888), .out(n11888_0));
mux15 mux_6723 (.in({n14349_0, n14328_0, n14313_0, n14305_0, n14300_0, n14277_0, n14272_0, n14248_1, n14245_0, n11975_0, n7223/**/, n7215, n7127, n7119, n7111}), .out(n11889), .config_in(config_chain[23649:23644]), .config_rst(config_rst)); 
buffer_wire buffer_11889 (.in(n11889), .out(n11889_0));
mux15 mux_6724 (.in({n13281_0, n13269_0, n13262_0/**/, n13248_0, n13233_0, n13219_0, n13212_0, n13202_1, n13129_0, n11778_0, n4293, n4285, n4277, n4185, n4177}), .out(n11890), .config_in(config_chain[23655:23650]), .config_rst(config_rst)); 
buffer_wire buffer_11890 (.in(n11890), .out(n11890_0));
mux15 mux_6725 (.in({n14347_0, n14327_0, n14322_0, n14299_0, n14294_0, n14286_0, n14271_0, n14267_0, n14250_1/**/, n11977_0, n7223, n7215, n7127, n7119, n7111}), .out(n11891), .config_in(config_chain[23661:23656]), .config_rst(config_rst)); 
buffer_wire buffer_11891 (.in(n11891), .out(n11891_0));
mux14 mux_6726 (.in({n13283_0, n13270_0, n13255_0, n13241_0, n13234_0, n13227_0, n13220_0, n13200_1, n11786_0, n4293, n4285/**/, n4277, n4189, n4177}), .out(n11892), .config_in(config_chain[23667:23662]), .config_rst(config_rst)); 
buffer_wire buffer_11892 (.in(n11892), .out(n11892_0));
mux15 mux_6727 (.in({n14345_0, n14321_0, n14316_0, n14308_0/**/, n14293_0, n14289_0, n14285_0, n14280_0, n14252_1, n11979_0, n7223, n7215, n7127, n7119, n7111}), .out(n11893), .config_in(config_chain[23673:23668]), .config_rst(config_rst)); 
buffer_wire buffer_11893 (.in(n11893), .out(n11893_0));
mux14 mux_6728 (.in({n13285_0, n13263_0, n13256_0, n13249_0, n13242_0, n13228_0/**/, n13213_0, n13198_1, n11794_0, n4293, n4285, n4277, n4189, n4181}), .out(n11894), .config_in(config_chain[23679:23674]), .config_rst(config_rst)); 
buffer_wire buffer_11894 (.in(n11894), .out(n11894_0));
mux15 mux_6729 (.in({n14343_0, n14330_0, n14315_0, n14311_0, n14307_0, n14302_0, n14279_0, n14274_0/**/, n14254_1, n11981_0, n7227, n7219, n7211, n7123, n7115}), .out(n11895), .config_in(config_chain[23685:23680]), .config_rst(config_rst)); 
buffer_wire buffer_11895 (.in(n11895), .out(n11895_0));
mux13 mux_6730 (.in({n13287_0, n13271_0, n13264_0/**/, n13250_0, n13235_0, n13221_0, n13214_0, n13196_1, n11802_0, n4285, n4277, n4189, n4181}), .out(n11896), .config_in(config_chain[23691:23686]), .config_rst(config_rst)); 
buffer_wire buffer_11896 (.in(n11896), .out(n11896_0));
mux15 mux_6731 (.in({n14341_0, n14329_0, n14324_0, n14301_0, n14296_0, n14273_0, n14268_0, n14256_1, n14200_2, n11983_0/**/, n7227, n7219, n7211, n7123, n7115}), .out(n11897), .config_in(config_chain[23697:23692]), .config_rst(config_rst)); 
buffer_wire buffer_11897 (.in(n11897), .out(n11897_0));
mux13 mux_6732 (.in({n13289_0, n13272_0, n13257_0, n13243_0, n13236_0, n13229_0, n13222_0, n13194_1, n11810_0, n4289/**/, n4277, n4189, n4181}), .out(n11898), .config_in(config_chain[23703:23698]), .config_rst(config_rst)); 
buffer_wire buffer_11898 (.in(n11898), .out(n11898_0));
mux15 mux_6733 (.in({n14339_0, n14323_0, n14318_0, n14295_0, n14290_0, n14287_0, n14282_0, n14258_1, n14222_1, n11985_0, n7227, n7219, n7211, n7123, n7115}), .out(n11899), .config_in(config_chain[23709:23704]), .config_rst(config_rst)); 
buffer_wire buffer_11899 (.in(n11899), .out(n11899_0));
mux13 mux_6734 (.in({n13291_0, n13265_0, n13258_0/**/, n13251_0, n13244_0, n13230_0, n13215_0, n13192_1, n11818_0, n4289, n4281, n4189, n4181}), .out(n11900), .config_in(config_chain[23715:23710]), .config_rst(config_rst)); 
buffer_wire buffer_11900 (.in(n11900), .out(n11900_0));
mux15 mux_6735 (.in({n14337_0, n14317_0, n14312_0, n14309_0, n14304_0, n14281_0, n14276_0, n14260_1, n14244_1/**/, n11987_0, n7227, n7219, n7211, n7123, n7115}), .out(n11901), .config_in(config_chain[23721:23716]), .config_rst(config_rst)); 
buffer_wire buffer_11901 (.in(n11901), .out(n11901_0));
mux13 mux_6736 (.in({n13293_0, n13273_0, n13266_0, n13252_0/**/, n13237_0, n13223_0, n13216_0, n13190_1, n11826_0, n4289, n4281, n4193, n4181}), .out(n11902), .config_in(config_chain[23727:23722]), .config_rst(config_rst)); 
buffer_wire buffer_11902 (.in(n11902), .out(n11902_0));
mux15 mux_6737 (.in({n14335_0, n14331_0/**/, n14326_0, n14303_0, n14298_0, n14275_0, n14270_0, n14266_1, n14262_1, n11989_0, n7227, n7219, n7211, n7123, n7115}), .out(n11903), .config_in(config_chain[23733:23728]), .config_rst(config_rst)); 
buffer_wire buffer_11903 (.in(n11903), .out(n11903_0));
mux13 mux_6738 (.in({n13295_0, n13274_0, n13259_0, n13245_0, n13238_0, n13231_0, n13224_0, n13124_2, n11834_0, n4289, n4281, n4193/**/, n4185}), .out(n11904), .config_in(config_chain[23739:23734]), .config_rst(config_rst)); 
buffer_wire buffer_11904 (.in(n11904), .out(n11904_0));
mux3 mux_6739 (.in({n14749_0, n14748_1, n9179}), .out(n11905), .config_in(config_chain[23741:23740]), .config_rst(config_rst)); 
buffer_wire buffer_11905 (.in(n11905), .out(n11905_0));
mux15 mux_6740 (.in({n13559_0, n13536_0, n13529_0, n13522_0, n13508_0, n13493_0, n13479_0, n13472_0, n13468_1, n11748_1/**/, n5267, n5259, n5171, n5163, n5155}), .out(n11906), .config_in(config_chain[23747:23742]), .config_rst(config_rst)); 
buffer_wire buffer_11906 (.in(n11906), .out(n11906_0));
mux16 mux_6741 (.in({n14595_0, n14587_0, n14582_0, n14561_0, n14556_0, n14548_0, n14533_0, n14530_1, n14528_1, n14433_0, n11991_0, n8201/**/, n8193, n8105, n8097, n8089}), .out(n11907), .config_in(config_chain[23753:23748]), .config_rst(config_rst)); 
buffer_wire buffer_11907 (.in(n11907), .out(n11907_0));
mux15 mux_6742 (.in({n13539_0, n13530_0, n13515_0, n13501_0, n13494_0, n13487_0, n13480_0, n13466_1/**/, n13388_2, n11756_1, n5271, n5259, n5171, n5163, n5155}), .out(n11908), .config_in(config_chain[23759:23754]), .config_rst(config_rst)); 
buffer_wire buffer_11908 (.in(n11908), .out(n11908_0));
mux16 mux_6743 (.in({n14613_0, n14581_0, n14576_0, n14570_0, n14555_0, n14552_0, n14547_0, n14542_0, n14510_1, n14465_0, n11993_0, n8201, n8193, n8105/**/, n8097, n8089}), .out(n11909), .config_in(config_chain[23765:23760]), .config_rst(config_rst)); 
buffer_wire buffer_11909 (.in(n11909), .out(n11909_0));
mux15 mux_6744 (.in({n13541_0, n13537_0, n13523_0, n13516_0, n13509_0, n13502_0, n13488_0, n13473_0, n13464_1, n11764_1/**/, n5271, n5263, n5171, n5163, n5155}), .out(n11910), .config_in(config_chain[23771:23766]), .config_rst(config_rst)); 
buffer_wire buffer_11910 (.in(n11910), .out(n11910_0));
mux15 mux_6745 (.in({n14611_0, n14590_0, n14575_0, n14569_0, n14564_0, n14541_0, n14536_0, n14512_1/**/, n14487_0, n11995_0, n8201, n8193, n8105, n8097, n8089}), .out(n11911), .config_in(config_chain[23777:23772]), .config_rst(config_rst)); 
buffer_wire buffer_11911 (.in(n11911), .out(n11911_0));
mux15 mux_6746 (.in({n13543_0, n13531_0, n13524_0, n13510_0, n13495_0, n13481_0, n13474_0, n13462_1, n13389_0, n11772_1/**/, n5271, n5263, n5255, n5163, n5155}), .out(n11912), .config_in(config_chain[23783:23778]), .config_rst(config_rst)); 
buffer_wire buffer_11912 (.in(n11912), .out(n11912_0));
mux15 mux_6747 (.in({n14609_0, n14589_0, n14584_0/**/, n14563_0, n14558_0, n14550_0, n14535_0, n14514_1, n14509_0, n11997_0, n8201, n8193, n8105, n8097, n8089}), .out(n11913), .config_in(config_chain[23789:23784]), .config_rst(config_rst)); 
buffer_wire buffer_11913 (.in(n11913), .out(n11913_0));
mux14 mux_6748 (.in({n13545_0, n13532_0, n13517_0, n13503_0, n13496_0, n13489_0, n13482_0, n13460_1, n11780_1/**/, n5271, n5263, n5255, n5167, n5155}), .out(n11914), .config_in(config_chain[23795:23790]), .config_rst(config_rst)); 
buffer_wire buffer_11914 (.in(n11914), .out(n11914_0));
mux15 mux_6749 (.in({n14607_0, n14583_0, n14578_0, n14572_0/**/, n14557_0, n14549_0, n14544_0, n14531_0, n14516_1, n11999_0, n8201, n8193, n8105, n8097, n8089}), .out(n11915), .config_in(config_chain[23801:23796]), .config_rst(config_rst)); 
buffer_wire buffer_11915 (.in(n11915), .out(n11915_0));
mux14 mux_6750 (.in({n13547_0, n13525_0, n13518_0, n13511_0, n13504_0, n13490_0, n13475_0, n13458_1, n11788_1, n5271, n5263/**/, n5255, n5167, n5159}), .out(n11916), .config_in(config_chain[23807:23802]), .config_rst(config_rst)); 
buffer_wire buffer_11916 (.in(n11916), .out(n11916_0));
mux15 mux_6751 (.in({n14605_0, n14592_0, n14577_0, n14571_0, n14566_0/**/, n14553_0, n14543_0, n14538_0, n14518_1, n12001_0, n8205, n8197, n8189, n8101, n8093}), .out(n11917), .config_in(config_chain[23813:23808]), .config_rst(config_rst)); 
buffer_wire buffer_11917 (.in(n11917), .out(n11917_0));
mux13 mux_6752 (.in({n13549_0, n13533_0, n13526_0, n13512_0, n13497_0, n13483_0, n13476_0, n13456_1, n11796_1/**/, n5263, n5255, n5167, n5159}), .out(n11918), .config_in(config_chain[23819:23814]), .config_rst(config_rst)); 
buffer_wire buffer_11918 (.in(n11918), .out(n11918_0));
mux15 mux_6753 (.in({n14603_0, n14591_0, n14586_0, n14565_0, n14560_0, n14537_0, n14532_0/**/, n14520_1, n14432_2, n12003_0, n8205, n8197, n8189, n8101, n8093}), .out(n11919), .config_in(config_chain[23825:23820]), .config_rst(config_rst)); 
buffer_wire buffer_11919 (.in(n11919), .out(n11919_0));
mux13 mux_6754 (.in({n13551_0, n13534_0, n13519_0, n13505_0, n13498_0, n13491_0, n13484_0, n13454_1, n11804_1, n5267, n5255, n5167/**/, n5159}), .out(n11920), .config_in(config_chain[23831:23826]), .config_rst(config_rst)); 
buffer_wire buffer_11920 (.in(n11920), .out(n11920_0));
mux15 mux_6755 (.in({n14601_0, n14585_0, n14580_0, n14559_0, n14554_0, n14551_0, n14546_0, n14522_1/**/, n14464_2, n12005_0, n8205, n8197, n8189, n8101, n8093}), .out(n11921), .config_in(config_chain[23837:23832]), .config_rst(config_rst)); 
buffer_wire buffer_11921 (.in(n11921), .out(n11921_0));
mux13 mux_6756 (.in({n13553_0, n13527_0, n13520_0, n13513_0, n13506_0, n13477_0, n13470_1, n13452_1, n11812_1/**/, n5267, n5259, n5167, n5159}), .out(n11922), .config_in(config_chain[23843:23838]), .config_rst(config_rst)); 
buffer_wire buffer_11922 (.in(n11922), .out(n11922_0));
mux15 mux_6757 (.in({n14599_0, n14579_0, n14574_0, n14573_0, n14568_0, n14545_0, n14540_0, n14524_1, n14486_1, n12007_0, n8205, n8197, n8189, n8101, n8093/**/}), .out(n11923), .config_in(config_chain[23849:23844]), .config_rst(config_rst)); 
buffer_wire buffer_11923 (.in(n11923), .out(n11923_0));
mux13 mux_6758 (.in({n13555_0, n13535_0, n13528_0, n13499_0, n13492_0, n13485_0, n13478_0, n13450_1, n11820_1/**/, n5267, n5259, n5171, n5159}), .out(n11924), .config_in(config_chain[23855:23850]), .config_rst(config_rst)); 
buffer_wire buffer_11924 (.in(n11924), .out(n11924_0));
mux15 mux_6759 (.in({n14597_0, n14593_0, n14588_0, n14567_0, n14562_0, n14539_0, n14534_0, n14526_1, n14508_1, n12009_0/**/, n8205, n8197, n8189, n8101, n8093}), .out(n11925), .config_in(config_chain[23861:23856]), .config_rst(config_rst)); 
buffer_wire buffer_11925 (.in(n11925), .out(n11925_0));
mux13 mux_6760 (.in({n13557_0, n13521_0, n13514_0, n13507_0, n13500_0, n13486_0, n13471_0, n13386_2, n11836_1, n5267, n5259, n5171/**/, n5163}), .out(n11926), .config_in(config_chain[23867:23862]), .config_rst(config_rst)); 
buffer_wire buffer_11926 (.in(n11926), .out(n11926_0));
mux3 mux_6761 (.in({n14771_0, n14770_1/**/, n9179}), .out(n11927), .config_in(config_chain[23869:23868]), .config_rst(config_rst)); 
buffer_wire buffer_11927 (.in(n11927), .out(n11927_0));
mux15 mux_6762 (.in({n13823_0, n13787_0, n13780_0/**/, n13778_0, n13771_0, n13764_0, n13750_0, n13735_0, n13732_1, n11840_1, n6245, n6237, n6149, n6141, n6133}), .out(n11928), .config_in(config_chain[23875:23870]), .config_rst(config_rst)); 
buffer_wire buffer_11928 (.in(n11928), .out(n11928_0));
mux4 mux_6763 (.in({n14855_0, n14772_1, n9183, n9067/**/}), .out(n11929), .config_in(config_chain[23877:23876]), .config_rst(config_rst)); 
buffer_wire buffer_11929 (.in(n11929), .out(n11929_0));
mux15 mux_6764 (.in({n13803_0, n13800_0, n13795_0, n13788_0, n13772_0, n13757_0, n13743_0, n13736_0/**/, n13730_1, n11842_1, n6249, n6237, n6149, n6141, n6133}), .out(n11930), .config_in(config_chain[23883:23878]), .config_rst(config_rst)); 
buffer_wire buffer_11930 (.in(n11930), .out(n11930_0));
mux3 mux_6765 (.in({n14857_0, n14774_1/**/, n9071}), .out(n11931), .config_in(config_chain[23885:23884]), .config_rst(config_rst)); 
buffer_wire buffer_11931 (.in(n11931), .out(n11931_0));
mux15 mux_6766 (.in({n13805_0, n13796_0, n13781_0, n13779_0, n13765_0, n13758_0, n13751_0, n13744_0, n13728_1, n11844_1, n6249, n6241, n6149, n6141, n6133}), .out(n11932), .config_in(config_chain[23891:23886]), .config_rst(config_rst)); 
buffer_wire buffer_11932 (.in(n11932), .out(n11932_0));
mux3 mux_6767 (.in({n14859_0, n14776_1, n9071}), .out(n11933), .config_in(config_chain[23893:23892]), .config_rst(config_rst)); 
buffer_wire buffer_11933 (.in(n11933), .out(n11933_0));
mux15 mux_6768 (.in({n13807_0, n13801_0, n13789_0/**/, n13782_0, n13773_0, n13766_0, n13752_0, n13737_0, n13726_1, n11846_1, n6249, n6241, n6233, n6141, n6133}), .out(n11934), .config_in(config_chain[23899:23894]), .config_rst(config_rst)); 
buffer_wire buffer_11934 (.in(n11934), .out(n11934_0));
mux3 mux_6769 (.in({n14861_0, n14778_1/**/, n9075}), .out(n11935), .config_in(config_chain[23901:23900]), .config_rst(config_rst)); 
buffer_wire buffer_11935 (.in(n11935), .out(n11935_0));
mux14 mux_6770 (.in({n13809_0, n13797_0, n13790_0, n13774_0, n13759_0, n13745_0, n13738_0, n13724_1, n11848_1/**/, n6249, n6241, n6233, n6145, n6133}), .out(n11936), .config_in(config_chain[23907:23902]), .config_rst(config_rst)); 
buffer_wire buffer_11936 (.in(n11936), .out(n11936_0));
mux3 mux_6771 (.in({n14863_0/**/, n14780_1, n9079}), .out(n11937), .config_in(config_chain[23909:23908]), .config_rst(config_rst)); 
buffer_wire buffer_11937 (.in(n11937), .out(n11937_0));
mux14 mux_6772 (.in({n13811_0, n13798_0, n13783_0, n13767_0, n13760_0, n13753_0, n13746_0, n13722_1, n11850_1/**/, n6249, n6241, n6233, n6145, n6137}), .out(n11938), .config_in(config_chain[23915:23910]), .config_rst(config_rst)); 
buffer_wire buffer_11938 (.in(n11938), .out(n11938_0));
mux3 mux_6773 (.in({n14865_0, n14782_1, n9083}), .out(n11939), .config_in(config_chain[23917:23916]), .config_rst(config_rst)); 
buffer_wire buffer_11939 (.in(n11939), .out(n11939_0));
mux13 mux_6774 (.in({n13813_0, n13791_0, n13784_0/**/, n13775_0, n13768_0, n13754_0, n13739_0, n13720_1, n11852_1, n6241, n6233, n6145, n6137}), .out(n11940), .config_in(config_chain[23923:23918]), .config_rst(config_rst)); 
buffer_wire buffer_11940 (.in(n11940), .out(n11940_0));
mux3 mux_6775 (.in({n14867_0, n14784_1, n9167}), .out(n11941), .config_in(config_chain[23925:23924]), .config_rst(config_rst)); 
buffer_wire buffer_11941 (.in(n11941), .out(n11941_0));
mux13 mux_6776 (.in({n13815_0, n13799_0, n13792_0, n13776_0, n13761_0, n13747_0, n13740_0, n13718_1, n11854_1, n6245, n6233, n6145, n6137}), .out(n11942), .config_in(config_chain[23931:23926]), .config_rst(config_rst)); 
buffer_wire buffer_11942 (.in(n11942), .out(n11942_0));
mux3 mux_6777 (.in({n14869_0, n14786_1/**/, n9167}), .out(n11943), .config_in(config_chain[23933:23932]), .config_rst(config_rst)); 
buffer_wire buffer_11943 (.in(n11943), .out(n11943_0));
mux13 mux_6778 (.in({n13817_0, n13785_0, n13769_0, n13762_0, n13755_0, n13748_0, n13716_1, n13712_1, n11856_1, n6245, n6237, n6145, n6137}), .out(n11944), .config_in(config_chain[23939:23934]), .config_rst(config_rst)); 
buffer_wire buffer_11944 (.in(n11944), .out(n11944_0));
mux3 mux_6779 (.in({n14871_0, n14788_1/**/, n9171}), .out(n11945), .config_in(config_chain[23941:23940]), .config_rst(config_rst)); 
buffer_wire buffer_11945 (.in(n11945), .out(n11945_0));
mux13 mux_6780 (.in({n13819_0, n13793_0, n13786_0, n13777_0, n13770_0, n13741_0, n13734_1, n13714_1, n11858_1, n6245, n6237, n6149, n6137}), .out(n11946), .config_in(config_chain[23947:23942]), .config_rst(config_rst)); 
buffer_wire buffer_11946 (.in(n11946), .out(n11946_0));
mux3 mux_6781 (.in({n14873_0, n14790_1/**/, n9175}), .out(n11947), .config_in(config_chain[23949:23948]), .config_rst(config_rst)); 
buffer_wire buffer_11947 (.in(n11947), .out(n11947_0));
mux13 mux_6782 (.in({n13821_0, n13794_0, n13763_0, n13756_0, n13749_0, n13742_0/**/, n13713_0, n13650_2, n11838_1, n6245, n6237, n6149, n6141}), .out(n11948), .config_in(config_chain[23955:23950]), .config_rst(config_rst)); 
buffer_wire buffer_11948 (.in(n11948), .out(n11948_0));
mux3 mux_6783 (.in({n14793_0, n14792_1/**/, n9183}), .out(n11949), .config_in(config_chain[23957:23956]), .config_rst(config_rst)); 
buffer_wire buffer_11949 (.in(n11949), .out(n11949_0));
mux16 mux_6784 (.in({n14087_0, n14052_0/**/, n14049_0, n14045_0, n14041_0, n14024_0, n14014_0, n14011_0, n13996_1, n13956_1, n11862_1, n7223, n7215, n7127, n7119, n7111}), .out(n11950), .config_in(config_chain[23963:23958]), .config_rst(config_rst)); 
buffer_wire buffer_11950 (.in(n11950), .out(n11950_0));
mux4 mux_6785 (.in({n14795_0, n14794_0, n9183, n9067}), .out(n11951), .config_in(config_chain[23965:23964]), .config_rst(config_rst)); 
buffer_wire buffer_11951 (.in(n11951), .out(n11951_0));
mux16 mux_6786 (.in({n14069_0, n14067_0, n14063_0, n14046_0, n14038_0, n14035_0, n14008_0/**/, n14005_0, n13994_1, n13978_1, n11864_1, n7223, n7215, n7127, n7119, n7111}), .out(n11952), .config_in(config_chain[23971:23966]), .config_rst(config_rst)); 
buffer_wire buffer_11952 (.in(n11952), .out(n11952_0));
mux3 mux_6787 (.in({n14797_0, n14796_0/**/, n9071}), .out(n11953), .config_in(config_chain[23973:23972]), .config_rst(config_rst)); 
buffer_wire buffer_11953 (.in(n11953), .out(n11953_0));
mux15 mux_6788 (.in({n14071_0, n14060_0, n14057_0, n14032_0, n14029_0, n14019_0, n14002_0, n14000_1, n13992_1, n11866_1, n7223, n7215, n7127, n7119, n7111}), .out(n11954), .config_in(config_chain[23979:23974]), .config_rst(config_rst)); 
buffer_wire buffer_11954 (.in(n11954), .out(n11954_0));
mux3 mux_6789 (.in({n14799_0, n14798_0/**/, n9075}), .out(n11955), .config_in(config_chain[23981:23980]), .config_rst(config_rst)); 
buffer_wire buffer_11955 (.in(n11955), .out(n11955_0));
mux15 mux_6790 (.in({n14073_0, n14054_0/**/, n14051_0, n14043_0, n14026_0, n14022_0, n14016_0, n14013_0, n13990_1, n11868_1, n7223, n7215, n7127, n7119, n7111}), .out(n11956), .config_in(config_chain[23987:23982]), .config_rst(config_rst)); 
buffer_wire buffer_11956 (.in(n11956), .out(n11956_0));
mux3 mux_6791 (.in({n14801_0, n14800_0, n9075}), .out(n11957), .config_in(config_chain[23989:23988]), .config_rst(config_rst)); 
buffer_wire buffer_11957 (.in(n11957), .out(n11957_0));
mux15 mux_6792 (.in({n14075_0, n14065_0, n14048_0, n14044_0, n14040_0, n14037_0/**/, n14010_0, n14007_0, n13988_1, n11870_1, n7223, n7215, n7127, n7119, n7111}), .out(n11958), .config_in(config_chain[23995:23990]), .config_rst(config_rst)); 
buffer_wire buffer_11958 (.in(n11958), .out(n11958_0));
mux3 mux_6793 (.in({n14803_0, n14802_0, n9079}), .out(n11959), .config_in(config_chain[23997:23996]), .config_rst(config_rst)); 
buffer_wire buffer_11959 (.in(n11959), .out(n11959_0));
mux15 mux_6794 (.in({n14077_0, n14066_0, n14062_0, n14059_0, n14034_0, n14031_0, n14021_0, n14004_0, n13986_1/**/, n11872_1, n7227, n7219, n7211, n7123, n7115}), .out(n11960), .config_in(config_chain[24003:23998]), .config_rst(config_rst)); 
buffer_wire buffer_11960 (.in(n11960), .out(n11960_0));
mux3 mux_6795 (.in({n14805_0, n14804_0, n9083}), .out(n11961), .config_in(config_chain[24005:24004]), .config_rst(config_rst)); 
buffer_wire buffer_11961 (.in(n11961), .out(n11961_0));
mux15 mux_6796 (.in({n14079_0, n14056_0, n14053_0, n14028_0, n14025_0, n14018_0, n14015_0, n13984_1/**/, n13957_0, n11874_1, n7227, n7219, n7211, n7123, n7115}), .out(n11962), .config_in(config_chain[24011:24006]), .config_rst(config_rst)); 
buffer_wire buffer_11962 (.in(n11962), .out(n11962_0));
mux3 mux_6797 (.in({n14807_0, n14806_0, n9167}), .out(n11963), .config_in(config_chain[24013:24012]), .config_rst(config_rst)); 
buffer_wire buffer_11963 (.in(n11963), .out(n11963_0));
mux15 mux_6798 (.in({n14081_0, n14050_0, n14047_0, n14042_0, n14039_0, n14012_0, n14009_0/**/, n13982_1, n13979_0, n11876_1, n7227, n7219, n7211, n7123, n7115}), .out(n11964), .config_in(config_chain[24019:24014]), .config_rst(config_rst)); 
buffer_wire buffer_11964 (.in(n11964), .out(n11964_0));
mux3 mux_6799 (.in({n14809_0, n14808_0, n9171}), .out(n11965), .config_in(config_chain[24021:24020]), .config_rst(config_rst)); 
buffer_wire buffer_11965 (.in(n11965), .out(n11965_0));
mux15 mux_6800 (.in({n14083_0, n14064_0, n14061_0, n14036_0, n14033_0, n14006_0, n14003_0, n14001_0, n13980_1, n11878_1, n7227, n7219, n7211, n7123, n7115}), .out(n11966), .config_in(config_chain[24027:24022]), .config_rst(config_rst)); 
buffer_wire buffer_11966 (.in(n11966), .out(n11966_0));
mux3 mux_6801 (.in({n14811_0, n14810_0, n9171}), .out(n11967), .config_in(config_chain[24029:24028]), .config_rst(config_rst)); 
buffer_wire buffer_11967 (.in(n11967), .out(n11967_0));
mux15 mux_6802 (.in({n14085_0, n14058_0, n14055_0, n14030_0, n14027_0, n14023_0, n14020_0, n14017_0, n13998_1/**/, n11880_1, n7227, n7219, n7211, n7123, n7115}), .out(n11968), .config_in(config_chain[24035:24030]), .config_rst(config_rst)); 
buffer_wire buffer_11968 (.in(n11968), .out(n11968_0));
mux3 mux_6803 (.in({n14813_0, n14812_0/**/, n9175}), .out(n11969), .config_in(config_chain[24037:24036]), .config_rst(config_rst)); 
buffer_wire buffer_11969 (.in(n11969), .out(n11969_0));
mux16 mux_6804 (.in({n14351_0, n14324_0, n14321_0, n14296_0, n14293_0, n14289_0, n14285_0, n14268_0/**/, n14262_1, n14200_2, n11884_1, n8201, n8193, n8105, n8097, n8089}), .out(n11970), .config_in(config_chain[24043:24038]), .config_rst(config_rst)); 
buffer_wire buffer_11970 (.in(n11970), .out(n11970_0));
mux4 mux_6805 (.in({n14815_0, n14814_0, n9183, n9067}), .out(n11971), .config_in(config_chain[24045:24044]), .config_rst(config_rst)); 
buffer_wire buffer_11971 (.in(n11971), .out(n11971_0));
mux16 mux_6806 (.in({n14333_0, n14318_0, n14315_0, n14311_0, n14307_0, n14290_0, n14282_0, n14279_0, n14260_1, n14222_1, n11886_1, n8201, n8193, n8105, n8097, n8089}), .out(n11972), .config_in(config_chain[24051:24046]), .config_rst(config_rst)); 
buffer_wire buffer_11972 (.in(n11972), .out(n11972_0));
mux3 mux_6807 (.in({n14817_0, n14816_0, n9071}), .out(n11973), .config_in(config_chain[24053:24052]), .config_rst(config_rst)); 
buffer_wire buffer_11973 (.in(n11973), .out(n11973_0));
mux15 mux_6808 (.in({n14335_0, n14329_0, n14312_0, n14304_0, n14301_0, n14276_0, n14273_0, n14258_1/**/, n14244_1, n11888_1, n8201, n8193, n8105, n8097, n8089}), .out(n11974), .config_in(config_chain[24059:24054]), .config_rst(config_rst)); 
buffer_wire buffer_11974 (.in(n11974), .out(n11974_0));
mux3 mux_6809 (.in({n14819_0, n14818_0, n9075}), .out(n11975), .config_in(config_chain[24061:24060]), .config_rst(config_rst)); 
buffer_wire buffer_11975 (.in(n11975), .out(n11975_0));
mux15 mux_6810 (.in({n14337_0/**/, n14326_0, n14323_0, n14298_0, n14295_0, n14287_0, n14270_0, n14266_1, n14256_1, n11890_1, n8201, n8193, n8105, n8097, n8089}), .out(n11976), .config_in(config_chain[24067:24062]), .config_rst(config_rst)); 
buffer_wire buffer_11976 (.in(n11976), .out(n11976_0));
mux3 mux_6811 (.in({n14821_0, n14820_0, n9079}), .out(n11977), .config_in(config_chain[24069:24068]), .config_rst(config_rst)); 
buffer_wire buffer_11977 (.in(n11977), .out(n11977_0));
mux15 mux_6812 (.in({n14339_0/**/, n14320_0, n14317_0, n14309_0, n14292_0, n14288_0, n14284_0, n14281_0, n14254_1, n11892_1, n8201, n8193, n8105, n8097, n8089}), .out(n11978), .config_in(config_chain[24075:24070]), .config_rst(config_rst)); 
buffer_wire buffer_11978 (.in(n11978), .out(n11978_0));
mux3 mux_6813 (.in({n14823_0, n14822_0, n9079}), .out(n11979), .config_in(config_chain[24077:24076]), .config_rst(config_rst)); 
buffer_wire buffer_11979 (.in(n11979), .out(n11979_0));
mux15 mux_6814 (.in({n14341_0, n14331_0, n14314_0, n14310_0, n14306_0, n14303_0, n14278_0, n14275_0, n14252_1, n11894_1, n8205, n8197, n8189, n8101, n8093/**/}), .out(n11980), .config_in(config_chain[24083:24078]), .config_rst(config_rst)); 
buffer_wire buffer_11980 (.in(n11980), .out(n11980_0));
mux3 mux_6815 (.in({n14825_0, n14824_0, n9083/**/}), .out(n11981), .config_in(config_chain[24085:24084]), .config_rst(config_rst)); 
buffer_wire buffer_11981 (.in(n11981), .out(n11981_0));
mux15 mux_6816 (.in({n14343_0, n14328_0, n14325_0, n14300_0, n14297_0, n14272_0, n14269_0, n14250_1/**/, n14201_0, n11896_1, n8205, n8197, n8189, n8101, n8093}), .out(n11982), .config_in(config_chain[24091:24086]), .config_rst(config_rst)); 
buffer_wire buffer_11982 (.in(n11982), .out(n11982_0));
mux3 mux_6817 (.in({n14827_0/**/, n14826_0, n9167}), .out(n11983), .config_in(config_chain[24093:24092]), .config_rst(config_rst)); 
buffer_wire buffer_11983 (.in(n11983), .out(n11983_0));
mux15 mux_6818 (.in({n14345_0, n14322_0, n14319_0, n14294_0, n14291_0, n14286_0, n14283_0, n14248_1, n14223_0, n11898_1/**/, n8205, n8197, n8189, n8101, n8093}), .out(n11984), .config_in(config_chain[24099:24094]), .config_rst(config_rst)); 
buffer_wire buffer_11984 (.in(n11984), .out(n11984_0));
mux3 mux_6819 (.in({n14829_0, n14828_0, n9171}), .out(n11985), .config_in(config_chain[24101:24100]), .config_rst(config_rst)); 
buffer_wire buffer_11985 (.in(n11985), .out(n11985_0));
mux15 mux_6820 (.in({n14347_0, n14316_0, n14313_0, n14308_0, n14305_0, n14280_0, n14277_0, n14246_1, n14245_0, n11900_1, n8205, n8197/**/, n8189, n8101, n8093}), .out(n11986), .config_in(config_chain[24107:24102]), .config_rst(config_rst)); 
buffer_wire buffer_11986 (.in(n11986), .out(n11986_0));
mux3 mux_6821 (.in({n14831_0, n14830_0, n9175}), .out(n11987), .config_in(config_chain[24109:24108]), .config_rst(config_rst)); 
buffer_wire buffer_11987 (.in(n11987), .out(n11987_0));
mux15 mux_6822 (.in({n14349_0, n14330_0, n14327_0, n14302_0, n14299_0, n14274_0, n14271_0, n14267_0, n14264_1, n11902_1, n8205, n8197, n8189, n8101, n8093}), .out(n11988), .config_in(config_chain[24115:24110]), .config_rst(config_rst)); 
buffer_wire buffer_11988 (.in(n11988), .out(n11988_0));
mux3 mux_6823 (.in({n14833_0, n14832_0, n9175}), .out(n11989), .config_in(config_chain[24117:24116]), .config_rst(config_rst)); 
buffer_wire buffer_11989 (.in(n11989), .out(n11989_0));
mux16 mux_6824 (.in({n14613_0, n14586_0, n14583_0, n14560_0, n14557_0, n14549_0, n14532_0, n14531_0, n14526_1, n14432_2, n11906_1, n9179, n9171, n9083, n9075, n9067}), .out(n11990), .config_in(config_chain[24123:24118]), .config_rst(config_rst)); 
buffer_wire buffer_11990 (.in(n11990), .out(n11990_0));
mux4 mux_6825 (.in({n14835_0, n14834_0, n9183, n9067}), .out(n11991), .config_in(config_chain[24125:24124]), .config_rst(config_rst)); 
buffer_wire buffer_11991 (.in(n11991), .out(n11991_0));
mux16 mux_6826 (.in({n14595_0, n14580_0, n14577_0, n14571_0, n14554_0/**/, n14553_0, n14546_0, n14543_0, n14524_1, n14464_2, n11908_1, n9179, n9171, n9083, n9075, n9067}), .out(n11992), .config_in(config_chain[24131:24126]), .config_rst(config_rst)); 
buffer_wire buffer_11992 (.in(n11992), .out(n11992_0));
mux3 mux_6827 (.in({n14837_0, n14836_0, n9067}), .out(n11993), .config_in(config_chain[24133:24132]), .config_rst(config_rst)); 
buffer_wire buffer_11993 (.in(n11993), .out(n11993_0));
mux15 mux_6828 (.in({n14597_0, n14591_0, n14574_0, n14568_0, n14565_0, n14540_0, n14537_0, n14522_1/**/, n14486_1, n11910_1, n9179, n9171, n9083, n9075, n9067}), .out(n11994), .config_in(config_chain[24139:24134]), .config_rst(config_rst)); 
buffer_wire buffer_11994 (.in(n11994), .out(n11994_0));
mux3 mux_6829 (.in({n14839_0, n14838_0/**/, n9071}), .out(n11995), .config_in(config_chain[24141:24140]), .config_rst(config_rst)); 
buffer_wire buffer_11995 (.in(n11995), .out(n11995_0));
mux15 mux_6830 (.in({n14599_0, n14588_0, n14585_0, n14562_0, n14559_0, n14551_0, n14534_0, n14520_1, n14508_1, n11912_1/**/, n9179, n9171, n9083, n9075, n9067}), .out(n11996), .config_in(config_chain[24147:24142]), .config_rst(config_rst)); 
buffer_wire buffer_11996 (.in(n11996), .out(n11996_0));
mux3 mux_6831 (.in({n14841_0, n14840_0, n9075}), .out(n11997), .config_in(config_chain[24149:24148]), .config_rst(config_rst)); 
buffer_wire buffer_11997 (.in(n11997), .out(n11997_0));
mux15 mux_6832 (.in({n14601_0, n14582_0, n14579_0, n14573_0, n14556_0, n14548_0, n14545_0, n14530_1, n14518_1, n11914_1/**/, n9179, n9171, n9083, n9075, n9067}), .out(n11998), .config_in(config_chain[24155:24150]), .config_rst(config_rst)); 
buffer_wire buffer_11998 (.in(n11998), .out(n11998_0));
mux3 mux_6833 (.in({n14843_0, n14842_0/**/, n9079}), .out(n11999), .config_in(config_chain[24157:24156]), .config_rst(config_rst)); 
buffer_wire buffer_11999 (.in(n11999), .out(n11999_0));
mux15 mux_6834 (.in({n14603_0/**/, n14593_0, n14576_0, n14570_0, n14567_0, n14552_0, n14542_0, n14539_0, n14516_1, n11916_1, n9183, n9175, n9167, n9079, n9071}), .out(n12000), .config_in(config_chain[24163:24158]), .config_rst(config_rst)); 
buffer_wire buffer_12000 (.in(n12000), .out(n12000_0));
mux3 mux_6835 (.in({n14845_0, n14844_0, n9083}), .out(n12001), .config_in(config_chain[24165:24164]), .config_rst(config_rst)); 
buffer_wire buffer_12001 (.in(n12001), .out(n12001_0));
mux15 mux_6836 (.in({n14605_0, n14590_0, n14587_0, n14564_0, n14561_0, n14536_0, n14533_0, n14514_1, n14433_0, n11918_1/**/, n9183, n9175, n9167, n9079, n9071}), .out(n12002), .config_in(config_chain[24171:24166]), .config_rst(config_rst)); 
buffer_wire buffer_12002 (.in(n12002), .out(n12002_0));
mux3 mux_6837 (.in({n14847_0, n14846_0, n9083}), .out(n12003), .config_in(config_chain[24173:24172]), .config_rst(config_rst)); 
buffer_wire buffer_12003 (.in(n12003), .out(n12003_0));
mux15 mux_6838 (.in({n14607_0, n14584_0, n14581_0, n14558_0, n14555_0, n14550_0, n14547_0, n14512_1, n14465_0, n11920_1, n9183, n9175, n9167, n9079, n9071}), .out(n12004), .config_in(config_chain[24179:24174]), .config_rst(config_rst)); 
buffer_wire buffer_12004 (.in(n12004), .out(n12004_0));
mux3 mux_6839 (.in({n14849_0, n14848_0, n9167}), .out(n12005), .config_in(config_chain[24181:24180]), .config_rst(config_rst)); 
buffer_wire buffer_12005 (.in(n12005), .out(n12005_0));
mux15 mux_6840 (.in({n14609_0, n14578_0, n14575_0, n14572_0, n14569_0/**/, n14544_0, n14541_0, n14510_1, n14487_0, n11922_1, n9183, n9175, n9167, n9079, n9071}), .out(n12006), .config_in(config_chain[24187:24182]), .config_rst(config_rst)); 
buffer_wire buffer_12006 (.in(n12006), .out(n12006_0));
mux3 mux_6841 (.in({n14851_0, n14850_0, n9171}), .out(n12007), .config_in(config_chain[24189:24188]), .config_rst(config_rst)); 
buffer_wire buffer_12007 (.in(n12007), .out(n12007_0));
mux15 mux_6842 (.in({n14611_0, n14592_0, n14589_0/**/, n14566_0, n14563_0, n14538_0, n14535_0, n14528_1, n14509_0, n11924_1, n9183, n9175, n9167, n9079, n9071}), .out(n12008), .config_in(config_chain[24195:24190]), .config_rst(config_rst)); 
buffer_wire buffer_12008 (.in(n12008), .out(n12008_0));
mux3 mux_6843 (.in({n14853_0/**/, n14852_0, n9175}), .out(n12009), .config_in(config_chain[24197:24196]), .config_rst(config_rst)); 
buffer_wire buffer_12009 (.in(n12009), .out(n12009_0));
mux3 mux_6844 (.in({n12358_2, n1399, n1341}), .out(n12010), .config_in(config_chain[24199:24198]), .config_rst(config_rst)); 
buffer_wire buffer_12010 (.in(n12010), .out(n12010_0));
mux12 mux_6845 (.in({n13280_0, n13264_0, n13248_0, n13210_1, n13126_2, n12147_1, n3361/**/, n3352, n3346, n3313, n3305, n3297}), .out(n12011), .config_in(config_chain[24205:24200]), .config_rst(config_rst)); 
buffer_wire buffer_12011 (.in(n12011), .out(n12011_0));
mux3 mux_6846 (.in({n12356_2, n1399, n1341}), .out(n12012), .config_in(config_chain[24207:24206]), .config_rst(config_rst)); 
buffer_wire buffer_12012 (.in(n12012), .out(n12012_0));
mux12 mux_6847 (.in({n13558_0, n13538_0, n13520_0, n13504_0, n13488_1, n12169_1, n4339, n4330, n4324, n4291, n4283/**/, n4275}), .out(n12013), .config_in(config_chain[24213:24208]), .config_rst(config_rst)); 
buffer_wire buffer_12013 (.in(n12013), .out(n12013_0));
mux3 mux_6848 (.in({n12354_2, n1399, n1341}), .out(n12014), .config_in(config_chain[24215:24214]), .config_rst(config_rst)); 
buffer_wire buffer_12014 (.in(n12014), .out(n12014_0));
mux12 mux_6849 (.in({n12774_0/**/, n12736_0, n12720_0, n12706_1, n12612_2, n12103_1, n1405, n1396, n1390, n1357, n1349, n1341}), .out(n12015), .config_in(config_chain[24221:24216]), .config_rst(config_rst)); 
buffer_wire buffer_12015 (.in(n12015), .out(n12015_0));
mux3 mux_6850 (.in({n12352_2, n1399, n1341}), .out(n12016), .config_in(config_chain[24223:24222]), .config_rst(config_rst)); 
buffer_wire buffer_12016 (.in(n12016), .out(n12016_0));
mux12 mux_6851 (.in({n13026_0, n13010_0, n12972_0/**/, n12956_1, n12868_2, n12125_1, n2383, n2374, n2368, n2335, n2327, n2319}), .out(n12017), .config_in(config_chain[24229:24224]), .config_rst(config_rst)); 
buffer_wire buffer_12017 (.in(n12017), .out(n12017_0));
mux3 mux_6852 (.in({n12522_0, n1402, n1341}), .out(n12018), .config_in(config_chain[24231:24230]), .config_rst(config_rst)); 
buffer_wire buffer_12018 (.in(n12018), .out(n12018_0));
mux12 mux_6853 (.in({n13286_0, n13270_0, n13232_0, n13216_1, n13128_2, n12149_1, n3361, n3355, n3346, n3313, n3305, n3297/**/}), .out(n12019), .config_in(config_chain[24237:24232]), .config_rst(config_rst)); 
buffer_wire buffer_12019 (.in(n12019), .out(n12019_0));
mux3 mux_6854 (.in({n12500_0, n1402, n1345}), .out(n12020), .config_in(config_chain[24239:24238]), .config_rst(config_rst)); 
buffer_wire buffer_12020 (.in(n12020), .out(n12020_0));
mux12 mux_6855 (.in({n13544_0, n13526_0, n13510_0, n13472_1, n13388_2, n12171_1, n4339, n4333, n4324, n4291, n4283, n4275/**/}), .out(n12021), .config_in(config_chain[24245:24240]), .config_rst(config_rst)); 
buffer_wire buffer_12021 (.in(n12021), .out(n12021_0));
mux3 mux_6856 (.in({n12480_0, n1402, n1345}), .out(n12022), .config_in(config_chain[24247:24246]), .config_rst(config_rst)); 
buffer_wire buffer_12022 (.in(n12022), .out(n12022_0));
mux12 mux_6857 (.in({n12758_0, n12742_0, n12726_0, n12712_1, n12614_2, n12105_1/**/, n1405, n1399, n1390, n1357, n1349, n1341}), .out(n12023), .config_in(config_chain[24253:24248]), .config_rst(config_rst)); 
buffer_wire buffer_12023 (.in(n12023), .out(n12023_0));
mux3 mux_6858 (.in({n12460_1/**/, n1402, n1345}), .out(n12024), .config_in(config_chain[24255:24254]), .config_rst(config_rst)); 
buffer_wire buffer_12024 (.in(n12024), .out(n12024_0));
mux12 mux_6859 (.in({n13032_0, n12994_0, n12978_0, n12962_1, n12870_2, n12127_1, n2383, n2377, n2368, n2335/**/, n2327, n2319}), .out(n12025), .config_in(config_chain[24261:24256]), .config_rst(config_rst)); 
buffer_wire buffer_12025 (.in(n12025), .out(n12025_0));
mux3 mux_6860 (.in({n12520_0/**/, n1402, n1345}), .out(n12026), .config_in(config_chain[24263:24262]), .config_rst(config_rst)); 
buffer_wire buffer_12026 (.in(n12026), .out(n12026_0));
mux11 mux_6861 (.in({n13292_0, n13254_0, n13238_0, n13222_1, n12151_1, n3361/**/, n3355, n3349, n3313, n3305, n3297}), .out(n12027), .config_in(config_chain[24269:24264]), .config_rst(config_rst)); 
buffer_wire buffer_12027 (.in(n12027), .out(n12027_0));
mux3 mux_6862 (.in({n12498_0/**/, n1405, n1345}), .out(n12028), .config_in(config_chain[24271:24270]), .config_rst(config_rst)); 
buffer_wire buffer_12028 (.in(n12028), .out(n12028_0));
mux11 mux_6863 (.in({n13550_0, n13532_0, n13494_0/**/, n13478_1, n12173_1, n4339, n4333, n4327, n4291, n4283, n4275}), .out(n12029), .config_in(config_chain[24277:24272]), .config_rst(config_rst)); 
buffer_wire buffer_12029 (.in(n12029), .out(n12029_0));
mux3 mux_6864 (.in({n12478_0/**/, n1405, n1349}), .out(n12030), .config_in(config_chain[24279:24278]), .config_rst(config_rst)); 
buffer_wire buffer_12030 (.in(n12030), .out(n12030_0));
mux11 mux_6865 (.in({n12764_0/**/, n12748_0, n12732_0, n12696_1, n12107_1, n1405, n1399, n1393, n1357, n1349, n1341}), .out(n12031), .config_in(config_chain[24285:24280]), .config_rst(config_rst)); 
buffer_wire buffer_12031 (.in(n12031), .out(n12031_0));
mux3 mux_6866 (.in({n12458_1, n1405, n1349}), .out(n12032), .config_in(config_chain[24287:24286]), .config_rst(config_rst)); 
buffer_wire buffer_12032 (.in(n12032), .out(n12032_0));
mux11 mux_6867 (.in({n13016_0, n13000_0, n12984_0/**/, n12968_1, n12129_1, n2383, n2377, n2371, n2335, n2327, n2319}), .out(n12033), .config_in(config_chain[24293:24288]), .config_rst(config_rst)); 
buffer_wire buffer_12033 (.in(n12033), .out(n12033_0));
mux3 mux_6868 (.in({n12518_0/**/, n1405, n1349}), .out(n12034), .config_in(config_chain[24295:24294]), .config_rst(config_rst)); 
buffer_wire buffer_12034 (.in(n12034), .out(n12034_0));
mux11 mux_6869 (.in({n13276_0, n13260_0, n13244_0, n13228_1, n12153_1, n3361/**/, n3355, n3349, n3343, n3305, n3297}), .out(n12035), .config_in(config_chain[24301:24296]), .config_rst(config_rst)); 
buffer_wire buffer_12035 (.in(n12035), .out(n12035_0));
mux3 mux_6870 (.in({n12496_0, n1405, n1349}), .out(n12036), .config_in(config_chain[24303:24302]), .config_rst(config_rst)); 
buffer_wire buffer_12036 (.in(n12036), .out(n12036_0));
mux11 mux_6871 (.in({n13556_0/**/, n13516_0, n13500_0, n13484_1, n12175_1, n4339, n4333, n4327, n4321, n4283, n4275}), .out(n12037), .config_in(config_chain[24309:24304]), .config_rst(config_rst)); 
buffer_wire buffer_12037 (.in(n12037), .out(n12037_0));
mux3 mux_6872 (.in({n12476_0, n1408, n1349}), .out(n12038), .config_in(config_chain[24311:24310]), .config_rst(config_rst)); 
buffer_wire buffer_12038 (.in(n12038), .out(n12038_0));
mux11 mux_6873 (.in({n12770_0, n12754_0, n12716_0, n12702_1, n12109_1, n1405, n1399, n1393, n1387, n1349, n1341}), .out(n12039), .config_in(config_chain[24317:24312]), .config_rst(config_rst)); 
buffer_wire buffer_12039 (.in(n12039), .out(n12039_0));
mux3 mux_6874 (.in({n12456_1, n1408, n1353}), .out(n12040), .config_in(config_chain[24319:24318]), .config_rst(config_rst)); 
buffer_wire buffer_12040 (.in(n12040), .out(n12040_0));
mux11 mux_6875 (.in({n13022_0, n13006_0, n12990_0, n12952_1, n12131_1, n2383, n2377, n2371, n2365, n2327, n2319}), .out(n12041), .config_in(config_chain[24325:24320]), .config_rst(config_rst)); 
buffer_wire buffer_12041 (.in(n12041), .out(n12041_0));
mux3 mux_6876 (.in({n12516_0/**/, n1408, n1353}), .out(n12042), .config_in(config_chain[24327:24326]), .config_rst(config_rst)); 
buffer_wire buffer_12042 (.in(n12042), .out(n12042_0));
mux11 mux_6877 (.in({n13282_0, n13266_0, n13250_0, n13212_1, n12155_1, n3361/**/, n3355, n3349, n3343, n3309, n3297}), .out(n12043), .config_in(config_chain[24333:24328]), .config_rst(config_rst)); 
buffer_wire buffer_12043 (.in(n12043), .out(n12043_0));
mux3 mux_6878 (.in({n12494_0, n1408, n1353}), .out(n12044), .config_in(config_chain[24335:24334]), .config_rst(config_rst)); 
buffer_wire buffer_12044 (.in(n12044), .out(n12044_0));
mux11 mux_6879 (.in({n13540_0, n13522_0, n13506_0, n13490_1/**/, n12177_1, n4339, n4333, n4327, n4321, n4287, n4275}), .out(n12045), .config_in(config_chain[24341:24336]), .config_rst(config_rst)); 
buffer_wire buffer_12045 (.in(n12045), .out(n12045_0));
mux3 mux_6880 (.in({n12474_0, n1408, n1353}), .out(n12046), .config_in(config_chain[24343:24342]), .config_rst(config_rst)); 
buffer_wire buffer_12046 (.in(n12046), .out(n12046_0));
mux11 mux_6881 (.in({n12776_0, n12738_0/**/, n12722_0, n12708_1, n12111_1, n1405, n1399, n1393, n1387, n1353, n1341}), .out(n12047), .config_in(config_chain[24349:24344]), .config_rst(config_rst)); 
buffer_wire buffer_12047 (.in(n12047), .out(n12047_0));
mux2 mux_6882 (.in({n12454_1/**/, n1353}), .out(n12048), .config_in(config_chain[24350:24350]), .config_rst(config_rst)); 
buffer_wire buffer_12048 (.in(n12048), .out(n12048_0));
mux11 mux_6883 (.in({n13028_0, n13012_0, n12974_0, n12958_1, n12133_1, n2383, n2377, n2371, n2365, n2331, n2319}), .out(n12049), .config_in(config_chain[24356:24351]), .config_rst(config_rst)); 
buffer_wire buffer_12049 (.in(n12049), .out(n12049_0));
mux2 mux_6884 (.in({n12514_0, n1357}), .out(n12050), .config_in(config_chain[24357:24357]), .config_rst(config_rst)); 
buffer_wire buffer_12050 (.in(n12050), .out(n12050_0));
mux11 mux_6885 (.in({n13288_0, n13272_0/**/, n13234_0, n13218_1, n12157_1, n3364, n3355, n3349, n3343, n3309, n3301}), .out(n12051), .config_in(config_chain[24363:24358]), .config_rst(config_rst)); 
buffer_wire buffer_12051 (.in(n12051), .out(n12051_0));
mux2 mux_6886 (.in({n12492_0/**/, n1357}), .out(n12052), .config_in(config_chain[24364:24364]), .config_rst(config_rst)); 
buffer_wire buffer_12052 (.in(n12052), .out(n12052_0));
mux11 mux_6887 (.in({n13546_0/**/, n13528_0, n13512_0, n13474_1, n12179_1, n4342, n4333, n4327, n4321, n4287, n4279}), .out(n12053), .config_in(config_chain[24370:24365]), .config_rst(config_rst)); 
buffer_wire buffer_12053 (.in(n12053), .out(n12053_0));
mux2 mux_6888 (.in({n12472_0/**/, n1357}), .out(n12054), .config_in(config_chain[24371:24371]), .config_rst(config_rst)); 
buffer_wire buffer_12054 (.in(n12054), .out(n12054_0));
mux11 mux_6889 (.in({n12760_0, n12744_0, n12728_0, n12714_1, n12113_1, n1408, n1399, n1393, n1387, n1353, n1345}), .out(n12055), .config_in(config_chain[24377:24372]), .config_rst(config_rst)); 
buffer_wire buffer_12055 (.in(n12055), .out(n12055_0));
mux2 mux_6890 (.in({n12452_1, n1357}), .out(n12056), .config_in(config_chain[24378:24378]), .config_rst(config_rst)); 
buffer_wire buffer_12056 (.in(n12056), .out(n12056_0));
mux11 mux_6891 (.in({n13034_0, n12996_0, n12980_0, n12964_1, n12135_1, n2386, n2377, n2371, n2365, n2331, n2323}), .out(n12057), .config_in(config_chain[24384:24379]), .config_rst(config_rst)); 
buffer_wire buffer_12057 (.in(n12057), .out(n12057_0));
mux2 mux_6892 (.in({n12512_0/**/, n1357}), .out(n12058), .config_in(config_chain[24385:24385]), .config_rst(config_rst)); 
buffer_wire buffer_12058 (.in(n12058), .out(n12058_0));
mux11 mux_6893 (.in({n13294_0, n13256_0, n13240_0/**/, n13224_1, n12159_1, n3364, n3358, n3349, n3343, n3309, n3301}), .out(n12059), .config_in(config_chain[24391:24386]), .config_rst(config_rst)); 
buffer_wire buffer_12059 (.in(n12059), .out(n12059_0));
mux2 mux_6894 (.in({n12490_0/**/, n1387}), .out(n12060), .config_in(config_chain[24392:24392]), .config_rst(config_rst)); 
buffer_wire buffer_12060 (.in(n12060), .out(n12060_0));
mux11 mux_6895 (.in({n13552_0/**/, n13534_0, n13496_0, n13480_1, n12181_1, n4342, n4336, n4327, n4321, n4287, n4279}), .out(n12061), .config_in(config_chain[24398:24393]), .config_rst(config_rst)); 
buffer_wire buffer_12061 (.in(n12061), .out(n12061_0));
mux2 mux_6896 (.in({n12470_0, n1387}), .out(n12062), .config_in(config_chain[24399:24399]), .config_rst(config_rst)); 
buffer_wire buffer_12062 (.in(n12062), .out(n12062_0));
mux11 mux_6897 (.in({n12766_0, n12750_0, n12734_0, n12698_1, n12115_1, n1408, n1402, n1393, n1387, n1353, n1345}), .out(n12063), .config_in(config_chain[24405:24400]), .config_rst(config_rst)); 
buffer_wire buffer_12063 (.in(n12063), .out(n12063_0));
mux2 mux_6898 (.in({n12450_1/**/, n1387}), .out(n12064), .config_in(config_chain[24406:24406]), .config_rst(config_rst)); 
buffer_wire buffer_12064 (.in(n12064), .out(n12064_0));
mux11 mux_6899 (.in({n13018_0, n13002_0/**/, n12986_0, n12970_1, n12137_1, n2386, n2380, n2371, n2365, n2331, n2323}), .out(n12065), .config_in(config_chain[24412:24407]), .config_rst(config_rst)); 
buffer_wire buffer_12065 (.in(n12065), .out(n12065_0));
mux2 mux_6900 (.in({n12510_0/**/, n1387}), .out(n12066), .config_in(config_chain[24413:24413]), .config_rst(config_rst)); 
buffer_wire buffer_12066 (.in(n12066), .out(n12066_0));
mux11 mux_6901 (.in({n13278_0, n13262_0/**/, n13246_0, n13230_1, n12161_1, n3364, n3358, n3352, n3343, n3309, n3301}), .out(n12067), .config_in(config_chain[24419:24414]), .config_rst(config_rst)); 
buffer_wire buffer_12067 (.in(n12067), .out(n12067_0));
mux2 mux_6902 (.in({n12488_0/**/, n1387}), .out(n12068), .config_in(config_chain[24420:24420]), .config_rst(config_rst)); 
buffer_wire buffer_12068 (.in(n12068), .out(n12068_0));
mux11 mux_6903 (.in({n13518_0, n13502_0/**/, n13486_1, n13470_1, n12183_1, n4342, n4336, n4330, n4321, n4287, n4279}), .out(n12069), .config_in(config_chain[24426:24421]), .config_rst(config_rst)); 
buffer_wire buffer_12069 (.in(n12069), .out(n12069_0));
mux2 mux_6904 (.in({n12468_0, n1390}), .out(n12070), .config_in(config_chain[24427:24427]), .config_rst(config_rst)); 
buffer_wire buffer_12070 (.in(n12070), .out(n12070_0));
mux11 mux_6905 (.in({n12772_0, n12756_0, n12718_0, n12704_1, n12117_1, n1408, n1402, n1396, n1387, n1353, n1345}), .out(n12071), .config_in(config_chain[24433:24428]), .config_rst(config_rst)); 
buffer_wire buffer_12071 (.in(n12071), .out(n12071_0));
mux2 mux_6906 (.in({n12448_1, n1390}), .out(n12072), .config_in(config_chain[24434:24434]), .config_rst(config_rst)); 
buffer_wire buffer_12072 (.in(n12072), .out(n12072_0));
mux11 mux_6907 (.in({n13024_0, n13008_0, n12992_0, n12954_1, n12139_1, n2386, n2380, n2374, n2365, n2331, n2323}), .out(n12073), .config_in(config_chain[24440:24435]), .config_rst(config_rst)); 
buffer_wire buffer_12073 (.in(n12073), .out(n12073_0));
mux2 mux_6908 (.in({n12508_0, n1390}), .out(n12074), .config_in(config_chain[24441:24441]), .config_rst(config_rst)); 
buffer_wire buffer_12074 (.in(n12074), .out(n12074_0));
mux11 mux_6909 (.in({n13284_0, n13268_0, n13252_0, n13214_1, n12163_1, n3364, n3358, n3352, n3346, n3309/**/, n3301}), .out(n12075), .config_in(config_chain[24447:24442]), .config_rst(config_rst)); 
buffer_wire buffer_12075 (.in(n12075), .out(n12075_0));
mux2 mux_6910 (.in({n12486_0, n1390}), .out(n12076), .config_in(config_chain[24448:24448]), .config_rst(config_rst)); 
buffer_wire buffer_12076 (.in(n12076), .out(n12076_0));
mux11 mux_6911 (.in({n13542_0/**/, n13524_0, n13508_0, n13492_1, n12185_1, n4342, n4336, n4330, n4324, n4287, n4279}), .out(n12077), .config_in(config_chain[24454:24449]), .config_rst(config_rst)); 
buffer_wire buffer_12077 (.in(n12077), .out(n12077_0));
mux2 mux_6912 (.in({n12466_0, n1390}), .out(n12078), .config_in(config_chain[24455:24455]), .config_rst(config_rst)); 
buffer_wire buffer_12078 (.in(n12078), .out(n12078_0));
mux11 mux_6913 (.in({n12778_0, n12740_0, n12724_0, n12710_1, n12119_1, n1408, n1402, n1396, n1390, n1353, n1345}), .out(n12079), .config_in(config_chain[24461:24456]), .config_rst(config_rst)); 
buffer_wire buffer_12079 (.in(n12079), .out(n12079_0));
mux2 mux_6914 (.in({n12446_1, n1393}), .out(n12080), .config_in(config_chain[24462:24462]), .config_rst(config_rst)); 
buffer_wire buffer_12080 (.in(n12080), .out(n12080_0));
mux11 mux_6915 (.in({n13030_0, n13014_0/**/, n12976_0, n12960_1, n12141_1, n2386, n2380, n2374, n2368, n2331, n2323}), .out(n12081), .config_in(config_chain[24468:24463]), .config_rst(config_rst)); 
buffer_wire buffer_12081 (.in(n12081), .out(n12081_0));
mux2 mux_6916 (.in({n12506_0/**/, n1393}), .out(n12082), .config_in(config_chain[24469:24469]), .config_rst(config_rst)); 
buffer_wire buffer_12082 (.in(n12082), .out(n12082_0));
mux11 mux_6917 (.in({n13290_0, n13274_0/**/, n13236_0, n13220_1, n12165_1, n3364, n3358, n3352, n3346, n3313, n3301}), .out(n12083), .config_in(config_chain[24475:24470]), .config_rst(config_rst)); 
buffer_wire buffer_12083 (.in(n12083), .out(n12083_0));
mux2 mux_6918 (.in({n12484_0/**/, n1393}), .out(n12084), .config_in(config_chain[24476:24476]), .config_rst(config_rst)); 
buffer_wire buffer_12084 (.in(n12084), .out(n12084_0));
mux11 mux_6919 (.in({n13548_0, n13530_0, n13514_0, n13476_1, n12187_1, n4342, n4336, n4330, n4324, n4291, n4279/**/}), .out(n12085), .config_in(config_chain[24482:24477]), .config_rst(config_rst)); 
buffer_wire buffer_12085 (.in(n12085), .out(n12085_0));
mux2 mux_6920 (.in({n12464_0, n1393}), .out(n12086), .config_in(config_chain[24483:24483]), .config_rst(config_rst)); 
buffer_wire buffer_12086 (.in(n12086), .out(n12086_0));
mux11 mux_6921 (.in({n12762_0, n12746_0, n12730_0, n12608_2, n12121_1, n1408, n1402, n1396, n1390, n1357, n1345}), .out(n12087), .config_in(config_chain[24489:24484]), .config_rst(config_rst)); 
buffer_wire buffer_12087 (.in(n12087), .out(n12087_0));
mux2 mux_6922 (.in({n12444_1/**/, n1393}), .out(n12088), .config_in(config_chain[24490:24490]), .config_rst(config_rst)); 
buffer_wire buffer_12088 (.in(n12088), .out(n12088_0));
mux11 mux_6923 (.in({n13036_0, n12998_0, n12982_0, n12966_1, n12143_1, n2386, n2380, n2374, n2368, n2335, n2323}), .out(n12089), .config_in(config_chain[24496:24491]), .config_rst(config_rst)); 
buffer_wire buffer_12089 (.in(n12089), .out(n12089_0));
mux2 mux_6924 (.in({n12504_0/**/, n1396}), .out(n12090), .config_in(config_chain[24497:24497]), .config_rst(config_rst)); 
buffer_wire buffer_12090 (.in(n12090), .out(n12090_0));
mux2 mux_6925 (.in({n14832_0/**/, n9220}), .out(n12091), .config_in(config_chain[24498:24498]), .config_rst(config_rst)); 
buffer_wire buffer_12091 (.in(n12091), .out(n12091_0));
mux2 mux_6926 (.in({n12482_0/**/, n1396}), .out(n12092), .config_in(config_chain[24499:24499]), .config_rst(config_rst)); 
buffer_wire buffer_12092 (.in(n12092), .out(n12092_0));
mux2 mux_6927 (.in({n14694_2, n9220}), .out(n12093), .config_in(config_chain[24500:24500]), .config_rst(config_rst)); 
buffer_wire buffer_12093 (.in(n12093), .out(n12093_0));
mux2 mux_6928 (.in({n12462_0/**/, n1396}), .out(n12094), .config_in(config_chain[24501:24501]), .config_rst(config_rst)); 
buffer_wire buffer_12094 (.in(n12094), .out(n12094_0));
mux10 mux_6929 (.in({n12768_0, n12752_0, n12700_1, n12610_2, n12123_2, n1402, n1396, n1390, n1357, n1349}), .out(n12095), .config_in(config_chain[24507:24502]), .config_rst(config_rst)); 
buffer_wire buffer_12095 (.in(n12095), .out(n12095_0));
mux2 mux_6930 (.in({n12442_1, n1396}), .out(n12096), .config_in(config_chain[24508:24508]), .config_rst(config_rst)); 
buffer_wire buffer_12096 (.in(n12096), .out(n12096_0));
mux10 mux_6931 (.in({n13020_0, n13004_0, n12988_0, n12866_2, n12145_2, n2380, n2374, n2368, n2335, n2327}), .out(n12097), .config_in(config_chain[24514:24509]), .config_rst(config_rst)); 
buffer_wire buffer_12097 (.in(n12097), .out(n12097_0));
mux2 mux_6932 (.in({n12502_0/**/, n1396}), .out(n12098), .config_in(config_chain[24515:24515]), .config_rst(config_rst)); 
buffer_wire buffer_12098 (.in(n12098), .out(n12098_0));
mux10 mux_6933 (.in({n13296_0, n13258_0, n13242_0, n13226_1, n12167_1, n3358, n3352, n3346, n3313, n3305}), .out(n12099), .config_in(config_chain[24521:24516]), .config_rst(config_rst)); 
buffer_wire buffer_12099 (.in(n12099), .out(n12099_0));
mux2 mux_6934 (.in({n12360_2, n1399}), .out(n12100), .config_in(config_chain[24522:24522]), .config_rst(config_rst)); 
buffer_wire buffer_12100 (.in(n12100), .out(n12100_0));
mux10 mux_6935 (.in({n13554_0, n13536_0, n13498_0/**/, n13482_1, n12189_1, n4336, n4330, n4324, n4291, n4283}), .out(n12101), .config_in(config_chain[24528:24523]), .config_rst(config_rst)); 
buffer_wire buffer_12101 (.in(n12101), .out(n12101_0));
mux12 mux_6936 (.in({n12774_0, n12736_0/**/, n12720_0, n12706_1, n12612_2, n12014_0, n2383, n2374, n2368, n2335, n2327, n2319}), .out(n12102), .config_in(config_chain[24534:24529]), .config_rst(config_rst)); 
buffer_wire buffer_12102 (.in(n12102), .out(n12102_0));
mux13 mux_6937 (.in({n13790_0/**/, n13780_0, n13750_1, n13740_1, n13712_1, n12191_1, n5320, n5314, n5308, n5302, n5269, n5261, n5253}), .out(n12103), .config_in(config_chain[24540:24535]), .config_rst(config_rst)); 
buffer_wire buffer_12103 (.in(n12103), .out(n12103_0));
mux12 mux_6938 (.in({n12758_0/**/, n12742_0, n12726_0, n12712_1, n12614_2, n12022_0, n2383, n2377, n2368, n2335, n2327, n2319}), .out(n12104), .config_in(config_chain[24546:24541]), .config_rst(config_rst)); 
buffer_wire buffer_12104 (.in(n12104), .out(n12104_0));
mux13 mux_6939 (.in({n13812_0, n13802_0, n13772_0/**/, n13762_0, n13734_1, n12193_1, n5320, n5314, n5308, n5302, n5269, n5261, n5253}), .out(n12105), .config_in(config_chain[24552:24547]), .config_rst(config_rst)); 
buffer_wire buffer_12105 (.in(n12105), .out(n12105_0));
mux11 mux_6940 (.in({n12764_0, n12748_0, n12732_0, n12696_1, n12030_0/**/, n2383, n2377, n2371, n2335, n2327, n2319}), .out(n12106), .config_in(config_chain[24558:24553]), .config_rst(config_rst)); 
buffer_wire buffer_12106 (.in(n12106), .out(n12106_0));
mux13 mux_6941 (.in({n13796_0, n13786_0, n13756_1, n13746_1/**/, n13736_1, n12195_1, n5320, n5314, n5308, n5302, n5269, n5261, n5253}), .out(n12107), .config_in(config_chain[24564:24559]), .config_rst(config_rst)); 
buffer_wire buffer_12107 (.in(n12107), .out(n12107_0));
mux11 mux_6942 (.in({n12770_0, n12754_0, n12716_0, n12702_1/**/, n12038_0, n2383, n2377, n2371, n2365, n2327, n2319}), .out(n12108), .config_in(config_chain[24570:24565]), .config_rst(config_rst)); 
buffer_wire buffer_12108 (.in(n12108), .out(n12108_0));
mux13 mux_6943 (.in({n13818_0, n13808_0, n13778_0, n13768_0, n13758_0, n12197_1/**/, n5320, n5314, n5308, n5302, n5269, n5261, n5253}), .out(n12109), .config_in(config_chain[24576:24571]), .config_rst(config_rst)); 
buffer_wire buffer_12109 (.in(n12109), .out(n12109_0));
mux11 mux_6944 (.in({n12776_0/**/, n12738_0, n12722_0, n12708_1, n12046_0, n2383, n2377, n2371, n2365, n2331, n2319}), .out(n12110), .config_in(config_chain[24582:24577]), .config_rst(config_rst)); 
buffer_wire buffer_12110 (.in(n12110), .out(n12110_0));
mux13 mux_6945 (.in({n13800_0/**/, n13792_0, n13782_0, n13752_1, n13742_1, n12199_1, n5320, n5314, n5308, n5302, n5269, n5261, n5253}), .out(n12111), .config_in(config_chain[24588:24583]), .config_rst(config_rst)); 
buffer_wire buffer_12111 (.in(n12111), .out(n12111_0));
mux11 mux_6946 (.in({n12760_0, n12744_0, n12728_0, n12714_1, n12054_0/**/, n2386, n2377, n2371, n2365, n2331, n2323}), .out(n12112), .config_in(config_chain[24594:24589]), .config_rst(config_rst)); 
buffer_wire buffer_12112 (.in(n12112), .out(n12112_0));
mux12 mux_6947 (.in({n13822_0, n13814_0, n13804_0, n13774_0, n13764_0, n12201_1, n5317, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12113), .config_in(config_chain[24600:24595]), .config_rst(config_rst)); 
buffer_wire buffer_12113 (.in(n12113), .out(n12113_0));
mux11 mux_6948 (.in({n12766_0, n12750_0, n12734_0, n12698_1, n12062_0, n2386, n2380, n2371, n2365, n2331/**/, n2323}), .out(n12114), .config_in(config_chain[24606:24601]), .config_rst(config_rst)); 
buffer_wire buffer_12114 (.in(n12114), .out(n12114_0));
mux11 mux_6949 (.in({n13798_0, n13788_0, n13748_1, n13738_1, n12203_1, n5317, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12115), .config_in(config_chain[24612:24607]), .config_rst(config_rst)); 
buffer_wire buffer_12115 (.in(n12115), .out(n12115_0));
mux11 mux_6950 (.in({n12772_0, n12756_0, n12718_0, n12704_1/**/, n12070_0, n2386, n2380, n2374, n2365, n2331, n2323}), .out(n12116), .config_in(config_chain[24618:24613]), .config_rst(config_rst)); 
buffer_wire buffer_12116 (.in(n12116), .out(n12116_0));
mux11 mux_6951 (.in({n13820_0, n13810_0, n13770_0, n13760_0, n12205_1, n5317, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12117), .config_in(config_chain[24624:24619]), .config_rst(config_rst)); 
buffer_wire buffer_12117 (.in(n12117), .out(n12117_0));
mux11 mux_6952 (.in({n12778_0/**/, n12740_0, n12724_0, n12710_1, n12078_0, n2386, n2380, n2374, n2368, n2331, n2323}), .out(n12118), .config_in(config_chain[24630:24625]), .config_rst(config_rst)); 
buffer_wire buffer_12118 (.in(n12118), .out(n12118_0));
mux11 mux_6953 (.in({n13794_0, n13784_0, n13754_1, n13744_1, n12207_1, n5317, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12119), .config_in(config_chain[24636:24631]), .config_rst(config_rst)); 
buffer_wire buffer_12119 (.in(n12119), .out(n12119_0));
mux11 mux_6954 (.in({n12762_0/**/, n12746_0, n12730_0, n12608_2, n12086_0, n2386, n2380, n2374, n2368, n2335, n2323}), .out(n12120), .config_in(config_chain[24642:24637]), .config_rst(config_rst)); 
buffer_wire buffer_12120 (.in(n12120), .out(n12120_0));
mux11 mux_6955 (.in({n13816_0, n13806_0, n13776_0, n13766_0, n12209_1, n5317, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12121), .config_in(config_chain[24648:24643]), .config_rst(config_rst)); 
buffer_wire buffer_12121 (.in(n12121), .out(n12121_0));
mux10 mux_6956 (.in({n12768_0, n12752_0, n12700_1, n12610_2, n12094_0/**/, n2380, n2374, n2368, n2335, n2327}), .out(n12122), .config_in(config_chain[24654:24649]), .config_rst(config_rst)); 
buffer_wire buffer_12122 (.in(n12122), .out(n12122_0));
mux2 mux_6957 (.in({n14696_2, n9220}), .out(n12123), .config_in(config_chain[24655:24655]), .config_rst(config_rst)); 
buffer_wire buffer_12123 (.in(n12123), .out(n12123_0));
mux12 mux_6958 (.in({n13026_0/**/, n13010_0, n12972_0, n12956_1, n12868_2, n12016_0, n3361, n3352, n3346, n3313, n3305, n3297}), .out(n12124), .config_in(config_chain[24661:24656]), .config_rst(config_rst)); 
buffer_wire buffer_12124 (.in(n12124), .out(n12124_0));
mux13 mux_6959 (.in({n14082_0, n14072_0, n14034_0/**/, n14024_0, n13956_2, n12211_0, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12125), .config_in(config_chain[24667:24662]), .config_rst(config_rst)); 
buffer_wire buffer_12125 (.in(n12125), .out(n12125_0));
mux12 mux_6960 (.in({n13032_0, n12994_0, n12978_0, n12962_1, n12870_2, n12024_0, n3361/**/, n3355, n3346, n3313, n3305, n3297}), .out(n12126), .config_in(config_chain[24673:24668]), .config_rst(config_rst)); 
buffer_wire buffer_12126 (.in(n12126), .out(n12126_0));
mux13 mux_6961 (.in({n14056_0, n14046_0, n14016_1, n14006_1, n13978_1, n12213_0, n6298, n6292, n6286, n6280, n6247, n6239/**/, n6231}), .out(n12127), .config_in(config_chain[24679:24674]), .config_rst(config_rst)); 
buffer_wire buffer_12127 (.in(n12127), .out(n12127_0));
mux11 mux_6962 (.in({n13016_0, n13000_0, n12984_0, n12968_1, n12032_0, n3361/**/, n3355, n3349, n3313, n3305, n3297}), .out(n12128), .config_in(config_chain[24685:24680]), .config_rst(config_rst)); 
buffer_wire buffer_12128 (.in(n12128), .out(n12128_0));
mux13 mux_6963 (.in({n14078_0/**/, n14068_0, n14040_0, n14030_0, n14000_1, n12215_0, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12129), .config_in(config_chain[24691:24686]), .config_rst(config_rst)); 
buffer_wire buffer_12129 (.in(n12129), .out(n12129_0));
mux11 mux_6964 (.in({n13022_0, n13006_0, n12990_0, n12952_1, n12040_0, n3361/**/, n3355, n3349, n3343, n3305, n3297}), .out(n12130), .config_in(config_chain[24697:24692]), .config_rst(config_rst)); 
buffer_wire buffer_12130 (.in(n12130), .out(n12130_0));
mux13 mux_6965 (.in({n14062_0, n14052_0, n14022_1, n14012_1, n14002_1/**/, n12217_0, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12131), .config_in(config_chain[24703:24698]), .config_rst(config_rst)); 
buffer_wire buffer_12131 (.in(n12131), .out(n12131_0));
mux11 mux_6966 (.in({n13028_0, n13012_0, n12974_0, n12958_1, n12048_0, n3361/**/, n3355, n3349, n3343, n3309, n3297}), .out(n12132), .config_in(config_chain[24709:24704]), .config_rst(config_rst)); 
buffer_wire buffer_12132 (.in(n12132), .out(n12132_0));
mux13 mux_6967 (.in({n14084_0, n14074_0, n14044_0, n14036_0/**/, n14026_0, n12219_0, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12133), .config_in(config_chain[24715:24710]), .config_rst(config_rst)); 
buffer_wire buffer_12133 (.in(n12133), .out(n12133_0));
mux11 mux_6968 (.in({n13034_0/**/, n12996_0, n12980_0, n12964_1, n12056_0, n3364, n3355, n3349, n3343, n3309, n3301}), .out(n12134), .config_in(config_chain[24721:24716]), .config_rst(config_rst)); 
buffer_wire buffer_12134 (.in(n12134), .out(n12134_0));
mux12 mux_6969 (.in({n14066_0/**/, n14058_0, n14048_0, n14018_1, n14008_1, n12221_0, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12135), .config_in(config_chain[24727:24722]), .config_rst(config_rst)); 
buffer_wire buffer_12135 (.in(n12135), .out(n12135_0));
mux11 mux_6970 (.in({n13018_0, n13002_0/**/, n12986_0, n12970_1, n12064_0, n3364, n3358, n3349, n3343, n3309, n3301}), .out(n12136), .config_in(config_chain[24733:24728]), .config_rst(config_rst)); 
buffer_wire buffer_12136 (.in(n12136), .out(n12136_0));
mux11 mux_6971 (.in({n14080_0, n14070_0/**/, n14042_0, n14032_0, n12223_0, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12137), .config_in(config_chain[24739:24734]), .config_rst(config_rst)); 
buffer_wire buffer_12137 (.in(n12137), .out(n12137_0));
mux11 mux_6972 (.in({n13024_0/**/, n13008_0, n12992_0, n12954_1, n12072_0, n3364, n3358, n3352, n3343, n3309, n3301}), .out(n12138), .config_in(config_chain[24745:24740]), .config_rst(config_rst)); 
buffer_wire buffer_12138 (.in(n12138), .out(n12138_0));
mux11 mux_6973 (.in({n14064_0, n14054_0, n14014_1, n14004_1, n12225_0, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12139), .config_in(config_chain[24751:24746]), .config_rst(config_rst)); 
buffer_wire buffer_12139 (.in(n12139), .out(n12139_0));
mux11 mux_6974 (.in({n13030_0, n13014_0, n12976_0, n12960_1/**/, n12080_0, n3364, n3358, n3352, n3346, n3309, n3301}), .out(n12140), .config_in(config_chain[24757:24752]), .config_rst(config_rst)); 
buffer_wire buffer_12140 (.in(n12140), .out(n12140_0));
mux11 mux_6975 (.in({n14086_0, n14076_0, n14038_0, n14028_0/**/, n12227_0, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12141), .config_in(config_chain[24763:24758]), .config_rst(config_rst)); 
buffer_wire buffer_12141 (.in(n12141), .out(n12141_0));
mux11 mux_6976 (.in({n13036_0, n12998_0, n12982_0, n12966_1, n12088_0/**/, n3364, n3358, n3352, n3346, n3313, n3301}), .out(n12142), .config_in(config_chain[24769:24764]), .config_rst(config_rst)); 
buffer_wire buffer_12142 (.in(n12142), .out(n12142_0));
mux11 mux_6977 (.in({n14060_0, n14050_0, n14020_1, n14010_1, n12229_0, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12143), .config_in(config_chain[24775:24770]), .config_rst(config_rst)); 
buffer_wire buffer_12143 (.in(n12143), .out(n12143_0));
mux10 mux_6978 (.in({n13020_0, n13004_0, n12988_0/**/, n12866_2, n12096_0, n3358, n3352, n3346, n3313, n3305}), .out(n12144), .config_in(config_chain[24781:24776]), .config_rst(config_rst)); 
buffer_wire buffer_12144 (.in(n12144), .out(n12144_0));
mux2 mux_6979 (.in({n14726_2, n9220}), .out(n12145), .config_in(config_chain[24782:24782]), .config_rst(config_rst)); 
buffer_wire buffer_12145 (.in(n12145), .out(n12145_0));
mux12 mux_6980 (.in({n13280_0/**/, n13264_0, n13248_0, n13210_1, n13126_2, n12010_0, n4339, n4330, n4324, n4291, n4283, n4275}), .out(n12146), .config_in(config_chain[24788:24783]), .config_rst(config_rst)); 
buffer_wire buffer_12146 (.in(n12146), .out(n12146_0));
mux13 mux_6981 (.in({n14326_0, n14316_0, n14278_1, n14268_1, n14200_2, n12231_0/**/, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12147), .config_in(config_chain[24794:24789]), .config_rst(config_rst)); 
buffer_wire buffer_12147 (.in(n12147), .out(n12147_0));
mux12 mux_6982 (.in({n13286_0, n13270_0/**/, n13232_0, n13216_1, n13128_2, n12018_0, n4339, n4333, n4324, n4291, n4283, n4275}), .out(n12148), .config_in(config_chain[24800:24795]), .config_rst(config_rst)); 
buffer_wire buffer_12148 (.in(n12148), .out(n12148_0));
mux13 mux_6983 (.in({n14346_0, n14336_0, n14300_0, n14290_0/**/, n14222_2, n12233_0, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12149), .config_in(config_chain[24806:24801]), .config_rst(config_rst)); 
buffer_wire buffer_12149 (.in(n12149), .out(n12149_0));
mux11 mux_6984 (.in({n13292_0, n13254_0, n13238_0, n13222_1, n12026_0/**/, n4339, n4333, n4327, n4291, n4283, n4275}), .out(n12150), .config_in(config_chain[24812:24807]), .config_rst(config_rst)); 
buffer_wire buffer_12150 (.in(n12150), .out(n12150_0));
mux13 mux_6985 (.in({n14322_0, n14312_0, n14284_1, n14274_1, n14244_1, n12235_0, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12151), .config_in(config_chain[24818:24813]), .config_rst(config_rst)); 
buffer_wire buffer_12151 (.in(n12151), .out(n12151_0));
mux11 mux_6986 (.in({n13276_0, n13260_0, n13244_0, n13228_1, n12034_0/**/, n4339, n4333, n4327, n4321, n4283, n4275}), .out(n12152), .config_in(config_chain[24824:24819]), .config_rst(config_rst)); 
buffer_wire buffer_12152 (.in(n12152), .out(n12152_0));
mux13 mux_6987 (.in({n14342_0/**/, n14332_0, n14306_0, n14296_0, n14266_1, n12237_0, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12153), .config_in(config_chain[24830:24825]), .config_rst(config_rst)); 
buffer_wire buffer_12153 (.in(n12153), .out(n12153_0));
mux11 mux_6988 (.in({n13282_0/**/, n13266_0, n13250_0, n13212_1, n12042_0, n4339, n4333, n4327, n4321, n4287, n4275}), .out(n12154), .config_in(config_chain[24836:24831]), .config_rst(config_rst)); 
buffer_wire buffer_12154 (.in(n12154), .out(n12154_0));
mux13 mux_6989 (.in({n14328_0/**/, n14318_0, n14288_1, n14280_1, n14270_1, n12239_0, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12155), .config_in(config_chain[24842:24837]), .config_rst(config_rst)); 
buffer_wire buffer_12155 (.in(n12155), .out(n12155_0));
mux11 mux_6990 (.in({n13288_0, n13272_0/**/, n13234_0, n13218_1, n12050_0, n4342, n4333, n4327, n4321, n4287, n4279}), .out(n12156), .config_in(config_chain[24848:24843]), .config_rst(config_rst)); 
buffer_wire buffer_12156 (.in(n12156), .out(n12156_0));
mux12 mux_6991 (.in({n14348_0, n14338_0, n14310_0, n14302_0/**/, n14292_0, n12241_0, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12157), .config_in(config_chain[24854:24849]), .config_rst(config_rst)); 
buffer_wire buffer_12157 (.in(n12157), .out(n12157_0));
mux11 mux_6992 (.in({n13294_0, n13256_0, n13240_0, n13224_1, n12058_0, n4342, n4336, n4327, n4321, n4287, n4279/**/}), .out(n12158), .config_in(config_chain[24860:24855]), .config_rst(config_rst)); 
buffer_wire buffer_12158 (.in(n12158), .out(n12158_0));
mux11 mux_6993 (.in({n14324_0, n14314_0/**/, n14286_1, n14276_1, n12243_0, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12159), .config_in(config_chain[24866:24861]), .config_rst(config_rst)); 
buffer_wire buffer_12159 (.in(n12159), .out(n12159_0));
mux11 mux_6994 (.in({n13278_0, n13262_0, n13246_0, n13230_1/**/, n12066_0, n4342, n4336, n4330, n4321, n4287, n4279}), .out(n12160), .config_in(config_chain[24872:24867]), .config_rst(config_rst)); 
buffer_wire buffer_12160 (.in(n12160), .out(n12160_0));
mux11 mux_6995 (.in({n14344_0, n14334_0, n14308_0, n14298_0, n12245_0, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12161), .config_in(config_chain[24878:24873]), .config_rst(config_rst)); 
buffer_wire buffer_12161 (.in(n12161), .out(n12161_0));
mux11 mux_6996 (.in({n13284_0/**/, n13268_0, n13252_0, n13214_1, n12074_0, n4342, n4336, n4330, n4324, n4287, n4279}), .out(n12162), .config_in(config_chain[24884:24879]), .config_rst(config_rst)); 
buffer_wire buffer_12162 (.in(n12162), .out(n12162_0));
mux11 mux_6997 (.in({n14330_0, n14320_0/**/, n14282_1, n14272_1, n12247_0, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12163), .config_in(config_chain[24890:24885]), .config_rst(config_rst)); 
buffer_wire buffer_12163 (.in(n12163), .out(n12163_0));
mux11 mux_6998 (.in({n13290_0, n13274_0, n13236_0, n13220_1, n12082_0/**/, n4342, n4336, n4330, n4324, n4291, n4279}), .out(n12164), .config_in(config_chain[24896:24891]), .config_rst(config_rst)); 
buffer_wire buffer_12164 (.in(n12164), .out(n12164_0));
mux11 mux_6999 (.in({n14350_0, n14340_0, n14304_0, n14294_0, n12249_0/**/, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12165), .config_in(config_chain[24902:24897]), .config_rst(config_rst)); 
buffer_wire buffer_12165 (.in(n12165), .out(n12165_0));
mux10 mux_7000 (.in({n13296_0, n13258_0, n13242_0, n13226_1/**/, n12098_0, n4336, n4330, n4324, n4291, n4283}), .out(n12166), .config_in(config_chain[24908:24903]), .config_rst(config_rst)); 
buffer_wire buffer_12166 (.in(n12166), .out(n12166_0));
mux2 mux_7001 (.in({n14748_2/**/, n9220}), .out(n12167), .config_in(config_chain[24909:24909]), .config_rst(config_rst)); 
buffer_wire buffer_12167 (.in(n12167), .out(n12167_0));
mux12 mux_7002 (.in({n13558_0, n13538_0, n13520_0/**/, n13504_0, n13488_1, n12012_1, n5317, n5308, n5302, n5269, n5261, n5253}), .out(n12168), .config_in(config_chain[24915:24910]), .config_rst(config_rst)); 
buffer_wire buffer_12168 (.in(n12168), .out(n12168_0));
mux13 mux_7003 (.in({n14604_0, n14594_0/**/, n14568_0, n14558_0, n14432_2, n12251_0, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12169), .config_in(config_chain[24921:24916]), .config_rst(config_rst)); 
buffer_wire buffer_12169 (.in(n12169), .out(n12169_0));
mux12 mux_7004 (.in({n13544_0, n13526_0/**/, n13510_0, n13472_1, n13388_2, n12020_1, n5317, n5311, n5302, n5269, n5261, n5253}), .out(n12170), .config_in(config_chain[24927:24922]), .config_rst(config_rst)); 
buffer_wire buffer_12170 (.in(n12170), .out(n12170_0));
mux13 mux_7005 (.in({n14588_0, n14578_0, n14542_1, n14532_1, n14464_2, n12253_0/**/, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12171), .config_in(config_chain[24933:24928]), .config_rst(config_rst)); 
buffer_wire buffer_12171 (.in(n12171), .out(n12171_0));
mux11 mux_7006 (.in({n13550_0, n13532_0, n13494_0, n13478_1, n12028_1, n5317, n5311/**/, n5305, n5269, n5261, n5253}), .out(n12172), .config_in(config_chain[24939:24934]), .config_rst(config_rst)); 
buffer_wire buffer_12172 (.in(n12172), .out(n12172_0));
mux13 mux_7007 (.in({n14610_0, n14600_0, n14564_0, n14554_0, n14486_2, n12255_0, n8254, n8248, n8242, n8236, n8203, n8195, n8187/**/}), .out(n12173), .config_in(config_chain[24945:24940]), .config_rst(config_rst)); 
buffer_wire buffer_12173 (.in(n12173), .out(n12173_0));
mux11 mux_7008 (.in({n13556_0, n13516_0/**/, n13500_0, n13484_1, n12036_1, n5317, n5311, n5305, n5299, n5261, n5253}), .out(n12174), .config_in(config_chain[24951:24946]), .config_rst(config_rst)); 
buffer_wire buffer_12174 (.in(n12174), .out(n12174_0));
mux13 mux_7009 (.in({n14584_0, n14574_0/**/, n14548_1, n14538_1, n14508_1, n12257_0, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12175), .config_in(config_chain[24957:24952]), .config_rst(config_rst)); 
buffer_wire buffer_12175 (.in(n12175), .out(n12175_0));
mux11 mux_7010 (.in({n13540_0, n13522_0, n13506_0, n13490_1, n12044_1, n5317, n5311/**/, n5305, n5299, n5265, n5253}), .out(n12176), .config_in(config_chain[24963:24958]), .config_rst(config_rst)); 
buffer_wire buffer_12176 (.in(n12176), .out(n12176_0));
mux13 mux_7011 (.in({n14606_0, n14596_0/**/, n14570_0, n14560_0, n14530_1, n12259_0, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12177), .config_in(config_chain[24969:24964]), .config_rst(config_rst)); 
buffer_wire buffer_12177 (.in(n12177), .out(n12177_0));
mux11 mux_7012 (.in({n13546_0, n13528_0, n13512_0, n13474_1, n12052_1, n5320, n5311/**/, n5305, n5299, n5265, n5257}), .out(n12178), .config_in(config_chain[24975:24970]), .config_rst(config_rst)); 
buffer_wire buffer_12178 (.in(n12178), .out(n12178_0));
mux12 mux_7013 (.in({n14590_0, n14580_0/**/, n14552_1, n14544_1, n14534_1, n12261_0, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12179), .config_in(config_chain[24981:24976]), .config_rst(config_rst)); 
buffer_wire buffer_12179 (.in(n12179), .out(n12179_0));
mux11 mux_7014 (.in({n13552_0, n13534_0, n13496_0, n13480_1/**/, n12060_1, n5320, n5314, n5305, n5299, n5265, n5257}), .out(n12180), .config_in(config_chain[24987:24982]), .config_rst(config_rst)); 
buffer_wire buffer_12180 (.in(n12180), .out(n12180_0));
mux11 mux_7015 (.in({n14612_0/**/, n14602_0, n14566_0, n14556_0, n12263_0, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12181), .config_in(config_chain[24993:24988]), .config_rst(config_rst)); 
buffer_wire buffer_12181 (.in(n12181), .out(n12181_0));
mux11 mux_7016 (.in({n13518_0, n13502_0, n13486_1, n13470_1, n12068_1, n5320, n5314, n5308, n5299, n5265, n5257}), .out(n12182), .config_in(config_chain[24999:24994]), .config_rst(config_rst)); 
buffer_wire buffer_12182 (.in(n12182), .out(n12182_0));
mux11 mux_7017 (.in({n14586_0, n14576_0, n14550_1, n14540_1, n12265_0, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12183), .config_in(config_chain[25005:25000]), .config_rst(config_rst)); 
buffer_wire buffer_12183 (.in(n12183), .out(n12183_0));
mux11 mux_7018 (.in({n13542_0/**/, n13524_0, n13508_0, n13492_1, n12076_1, n5320, n5314, n5308, n5302, n5265, n5257}), .out(n12184), .config_in(config_chain[25011:25006]), .config_rst(config_rst)); 
buffer_wire buffer_12184 (.in(n12184), .out(n12184_0));
mux11 mux_7019 (.in({n14608_0, n14598_0/**/, n14572_0, n14562_0, n12267_0, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12185), .config_in(config_chain[25017:25012]), .config_rst(config_rst)); 
buffer_wire buffer_12185 (.in(n12185), .out(n12185_0));
mux11 mux_7020 (.in({n13548_0/**/, n13530_0, n13514_0, n13476_1, n12084_1, n5320, n5314, n5308, n5302, n5269, n5257}), .out(n12186), .config_in(config_chain[25023:25018]), .config_rst(config_rst)); 
buffer_wire buffer_12186 (.in(n12186), .out(n12186_0));
mux11 mux_7021 (.in({n14592_0, n14582_0/**/, n14546_1, n14536_1, n12269_0, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12187), .config_in(config_chain[25029:25024]), .config_rst(config_rst)); 
buffer_wire buffer_12187 (.in(n12187), .out(n12187_0));
mux10 mux_7022 (.in({n13554_0, n13536_0, n13498_0, n13482_1/**/, n12100_1, n5314, n5308, n5302, n5269, n5261}), .out(n12188), .config_in(config_chain[25035:25030]), .config_rst(config_rst)); 
buffer_wire buffer_12188 (.in(n12188), .out(n12188_0));
mux2 mux_7023 (.in({n14770_1, n9223}), .out(n12189), .config_in(config_chain[25036:25036]), .config_rst(config_rst)); 
buffer_wire buffer_12189 (.in(n12189), .out(n12189_0));
mux13 mux_7024 (.in({n13790_0, n13780_0, n13750_1, n13740_1, n13712_1, n12102_1/**/, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12190), .config_in(config_chain[25042:25037]), .config_rst(config_rst)); 
buffer_wire buffer_12190 (.in(n12190), .out(n12190_0));
mux3 mux_7025 (.in({n14854_0/**/, n9223, n9165}), .out(n12191), .config_in(config_chain[25044:25043]), .config_rst(config_rst)); 
buffer_wire buffer_12191 (.in(n12191), .out(n12191_0));
mux13 mux_7026 (.in({n13812_0, n13802_0/**/, n13772_0, n13762_0, n13734_1, n12104_1, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12192), .config_in(config_chain[25050:25045]), .config_rst(config_rst)); 
buffer_wire buffer_12192 (.in(n12192), .out(n12192_0));
mux3 mux_7027 (.in({n14856_0/**/, n9226, n9169}), .out(n12193), .config_in(config_chain[25052:25051]), .config_rst(config_rst)); 
buffer_wire buffer_12193 (.in(n12193), .out(n12193_0));
mux13 mux_7028 (.in({n13796_0, n13786_0/**/, n13756_1, n13746_1, n13736_1, n12106_1, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12194), .config_in(config_chain[25058:25053]), .config_rst(config_rst)); 
buffer_wire buffer_12194 (.in(n12194), .out(n12194_0));
mux3 mux_7029 (.in({n14858_0/**/, n9229, n9173}), .out(n12195), .config_in(config_chain[25060:25059]), .config_rst(config_rst)); 
buffer_wire buffer_12195 (.in(n12195), .out(n12195_0));
mux13 mux_7030 (.in({n13818_0/**/, n13808_0, n13778_0, n13768_0, n13758_0, n12108_1, n6298, n6292, n6286, n6280, n6247, n6239, n6231}), .out(n12196), .config_in(config_chain[25066:25061]), .config_rst(config_rst)); 
buffer_wire buffer_12196 (.in(n12196), .out(n12196_0));
mux3 mux_7031 (.in({n14860_0/**/, n9232, n9173}), .out(n12197), .config_in(config_chain[25068:25067]), .config_rst(config_rst)); 
buffer_wire buffer_12197 (.in(n12197), .out(n12197_0));
mux13 mux_7032 (.in({n13800_0, n13792_0, n13782_0, n13752_1, n13742_1, n12110_1, n6298, n6292, n6286, n6280, n6247/**/, n6239, n6231}), .out(n12198), .config_in(config_chain[25074:25069]), .config_rst(config_rst)); 
buffer_wire buffer_12198 (.in(n12198), .out(n12198_0));
mux3 mux_7033 (.in({n14862_0, n9232, n9177}), .out(n12199), .config_in(config_chain[25076:25075]), .config_rst(config_rst)); 
buffer_wire buffer_12199 (.in(n12199), .out(n12199_0));
mux12 mux_7034 (.in({n13822_0, n13814_0/**/, n13804_0, n13774_0, n13764_0, n12112_1, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12200), .config_in(config_chain[25082:25077]), .config_rst(config_rst)); 
buffer_wire buffer_12200 (.in(n12200), .out(n12200_0));
mux2 mux_7035 (.in({n14864_0/**/, n9181}), .out(n12201), .config_in(config_chain[25083:25083]), .config_rst(config_rst)); 
buffer_wire buffer_12201 (.in(n12201), .out(n12201_0));
mux11 mux_7036 (.in({n13798_0, n13788_0/**/, n13748_1, n13738_1, n12114_1, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12202), .config_in(config_chain[25089:25084]), .config_rst(config_rst)); 
buffer_wire buffer_12202 (.in(n12202), .out(n12202_0));
mux2 mux_7037 (.in({n14866_0/**/, n9211}), .out(n12203), .config_in(config_chain[25090:25090]), .config_rst(config_rst)); 
buffer_wire buffer_12203 (.in(n12203), .out(n12203_0));
mux11 mux_7038 (.in({n13820_0, n13810_0, n13770_0, n13760_0, n12116_1, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12204), .config_in(config_chain[25096:25091]), .config_rst(config_rst)); 
buffer_wire buffer_12204 (.in(n12204), .out(n12204_0));
mux2 mux_7039 (.in({n14868_0/**/, n9214}), .out(n12205), .config_in(config_chain[25097:25097]), .config_rst(config_rst)); 
buffer_wire buffer_12205 (.in(n12205), .out(n12205_0));
mux11 mux_7040 (.in({n13794_0, n13784_0, n13754_1, n13744_1, n12118_1, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12206), .config_in(config_chain[25103:25098]), .config_rst(config_rst)); 
buffer_wire buffer_12206 (.in(n12206), .out(n12206_0));
mux2 mux_7041 (.in({n14870_0/**/, n9214}), .out(n12207), .config_in(config_chain[25104:25104]), .config_rst(config_rst)); 
buffer_wire buffer_12207 (.in(n12207), .out(n12207_0));
mux11 mux_7042 (.in({n13816_0, n13806_0/**/, n13776_0, n13766_0, n12120_1, n6295, n6289, n6283, n6277, n6243, n6235}), .out(n12208), .config_in(config_chain[25110:25105]), .config_rst(config_rst)); 
buffer_wire buffer_12208 (.in(n12208), .out(n12208_0));
mux2 mux_7043 (.in({n14872_0/**/, n9217}), .out(n12209), .config_in(config_chain[25111:25111]), .config_rst(config_rst)); 
buffer_wire buffer_12209 (.in(n12209), .out(n12209_0));
mux13 mux_7044 (.in({n14082_0, n14072_0, n14034_0, n14024_0, n13956_2, n12124_1, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12210), .config_in(config_chain[25117:25112]), .config_rst(config_rst)); 
buffer_wire buffer_12210 (.in(n12210), .out(n12210_0));
mux3 mux_7045 (.in({n14794_1, n9223, n9165}), .out(n12211), .config_in(config_chain[25119:25118]), .config_rst(config_rst)); 
buffer_wire buffer_12211 (.in(n12211), .out(n12211_0));
mux13 mux_7046 (.in({n14056_0, n14046_0, n14016_1, n14006_1, n13978_1, n12126_1/**/, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12212), .config_in(config_chain[25125:25120]), .config_rst(config_rst)); 
buffer_wire buffer_12212 (.in(n12212), .out(n12212_0));
mux3 mux_7047 (.in({n14796_1, n9226, n9169}), .out(n12213), .config_in(config_chain[25127:25126]), .config_rst(config_rst)); 
buffer_wire buffer_12213 (.in(n12213), .out(n12213_0));
mux13 mux_7048 (.in({n14078_0, n14068_0, n14040_0, n14030_0, n14000_1, n12128_1/**/, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12214), .config_in(config_chain[25133:25128]), .config_rst(config_rst)); 
buffer_wire buffer_12214 (.in(n12214), .out(n12214_0));
mux3 mux_7049 (.in({n14798_1/**/, n9229, n9173}), .out(n12215), .config_in(config_chain[25135:25134]), .config_rst(config_rst)); 
buffer_wire buffer_12215 (.in(n12215), .out(n12215_0));
mux13 mux_7050 (.in({n14062_0/**/, n14052_0, n14022_1, n14012_1, n14002_1, n12130_1, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12216), .config_in(config_chain[25141:25136]), .config_rst(config_rst)); 
buffer_wire buffer_12216 (.in(n12216), .out(n12216_0));
mux3 mux_7051 (.in({n14800_1, n9232, n9177}), .out(n12217), .config_in(config_chain[25143:25142]), .config_rst(config_rst)); 
buffer_wire buffer_12217 (.in(n12217), .out(n12217_0));
mux13 mux_7052 (.in({n14084_0, n14074_0, n14044_0, n14036_0, n14026_0, n12132_1/**/, n7276, n7270, n7264, n7258, n7225, n7217, n7209}), .out(n12218), .config_in(config_chain[25149:25144]), .config_rst(config_rst)); 
buffer_wire buffer_12218 (.in(n12218), .out(n12218_0));
mux2 mux_7053 (.in({n14802_1, n9177}), .out(n12219), .config_in(config_chain[25150:25150]), .config_rst(config_rst)); 
buffer_wire buffer_12219 (.in(n12219), .out(n12219_0));
mux12 mux_7054 (.in({n14066_0, n14058_0, n14048_0, n14018_1, n14008_1, n12134_1, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12220), .config_in(config_chain[25156:25151]), .config_rst(config_rst)); 
buffer_wire buffer_12220 (.in(n12220), .out(n12220_0));
mux2 mux_7055 (.in({n14804_1/**/, n9181}), .out(n12221), .config_in(config_chain[25157:25157]), .config_rst(config_rst)); 
buffer_wire buffer_12221 (.in(n12221), .out(n12221_0));
mux11 mux_7056 (.in({n14080_0, n14070_0, n14042_0, n14032_0, n12136_1/**/, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12222), .config_in(config_chain[25163:25158]), .config_rst(config_rst)); 
buffer_wire buffer_12222 (.in(n12222), .out(n12222_0));
mux2 mux_7057 (.in({n14806_1, n9211}), .out(n12223), .config_in(config_chain[25164:25164]), .config_rst(config_rst)); 
buffer_wire buffer_12223 (.in(n12223), .out(n12223_0));
mux11 mux_7058 (.in({n14064_0, n14054_0, n14014_1, n14004_1, n12138_1/**/, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12224), .config_in(config_chain[25170:25165]), .config_rst(config_rst)); 
buffer_wire buffer_12224 (.in(n12224), .out(n12224_0));
mux2 mux_7059 (.in({n14808_1, n9214}), .out(n12225), .config_in(config_chain[25171:25171]), .config_rst(config_rst)); 
buffer_wire buffer_12225 (.in(n12225), .out(n12225_0));
mux11 mux_7060 (.in({n14086_0, n14076_0, n14038_0/**/, n14028_0, n12140_1, n7273, n7267, n7261, n7255, n7221, n7213}), .out(n12226), .config_in(config_chain[25177:25172]), .config_rst(config_rst)); 
buffer_wire buffer_12226 (.in(n12226), .out(n12226_0));
mux2 mux_7061 (.in({n14810_1, n9217}), .out(n12227), .config_in(config_chain[25178:25178]), .config_rst(config_rst)); 
buffer_wire buffer_12227 (.in(n12227), .out(n12227_0));
mux11 mux_7062 (.in({n14060_0, n14050_0, n14020_1, n14010_1, n12142_1, n7273, n7267, n7261, n7255, n7221/**/, n7213}), .out(n12228), .config_in(config_chain[25184:25179]), .config_rst(config_rst)); 
buffer_wire buffer_12228 (.in(n12228), .out(n12228_0));
mux2 mux_7063 (.in({n14812_1, n9217}), .out(n12229), .config_in(config_chain[25185:25185]), .config_rst(config_rst)); 
buffer_wire buffer_12229 (.in(n12229), .out(n12229_0));
mux13 mux_7064 (.in({n14326_0, n14316_0, n14278_1, n14268_1, n14200_2, n12146_1/**/, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12230), .config_in(config_chain[25191:25186]), .config_rst(config_rst)); 
buffer_wire buffer_12230 (.in(n12230), .out(n12230_0));
mux3 mux_7065 (.in({n14792_1/**/, n9223, n9165}), .out(n12231), .config_in(config_chain[25193:25192]), .config_rst(config_rst)); 
buffer_wire buffer_12231 (.in(n12231), .out(n12231_0));
mux13 mux_7066 (.in({n14346_0, n14336_0, n14300_0, n14290_0, n14222_2, n12148_1, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12232), .config_in(config_chain[25199:25194]), .config_rst(config_rst)); 
buffer_wire buffer_12232 (.in(n12232), .out(n12232_0));
mux3 mux_7067 (.in({n14814_0, n9226, n9165}), .out(n12233), .config_in(config_chain[25201:25200]), .config_rst(config_rst)); 
buffer_wire buffer_12233 (.in(n12233), .out(n12233_0));
mux13 mux_7068 (.in({n14322_0, n14312_0, n14284_1, n14274_1, n14244_1, n12150_1, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12234), .config_in(config_chain[25207:25202]), .config_rst(config_rst)); 
buffer_wire buffer_12234 (.in(n12234), .out(n12234_0));
mux3 mux_7069 (.in({n14816_0/**/, n9226, n9169}), .out(n12235), .config_in(config_chain[25209:25208]), .config_rst(config_rst)); 
buffer_wire buffer_12235 (.in(n12235), .out(n12235_0));
mux13 mux_7070 (.in({n14342_0, n14332_0, n14306_0, n14296_0, n14266_1, n12152_1, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12236), .config_in(config_chain[25215:25210]), .config_rst(config_rst)); 
buffer_wire buffer_12236 (.in(n12236), .out(n12236_0));
mux3 mux_7071 (.in({n14818_0/**/, n9229, n9173}), .out(n12237), .config_in(config_chain[25217:25216]), .config_rst(config_rst)); 
buffer_wire buffer_12237 (.in(n12237), .out(n12237_0));
mux13 mux_7072 (.in({n14328_0, n14318_0, n14288_1, n14280_1, n14270_1, n12154_1, n8254, n8248, n8242, n8236, n8203, n8195, n8187}), .out(n12238), .config_in(config_chain[25223:25218]), .config_rst(config_rst)); 
buffer_wire buffer_12238 (.in(n12238), .out(n12238_0));
mux3 mux_7073 (.in({n14820_0/**/, n9232, n9177}), .out(n12239), .config_in(config_chain[25225:25224]), .config_rst(config_rst)); 
buffer_wire buffer_12239 (.in(n12239), .out(n12239_0));
mux12 mux_7074 (.in({n14348_0, n14338_0, n14310_0/**/, n14302_0, n14292_0, n12156_1, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12240), .config_in(config_chain[25231:25226]), .config_rst(config_rst)); 
buffer_wire buffer_12240 (.in(n12240), .out(n12240_0));
mux2 mux_7075 (.in({n14822_0, n9181}), .out(n12241), .config_in(config_chain[25232:25232]), .config_rst(config_rst)); 
buffer_wire buffer_12241 (.in(n12241), .out(n12241_0));
mux11 mux_7076 (.in({n14324_0, n14314_0, n14286_1, n14276_1, n12158_1, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12242), .config_in(config_chain[25238:25233]), .config_rst(config_rst)); 
buffer_wire buffer_12242 (.in(n12242), .out(n12242_0));
mux2 mux_7077 (.in({n14824_0, n9181}), .out(n12243), .config_in(config_chain[25239:25239]), .config_rst(config_rst)); 
buffer_wire buffer_12243 (.in(n12243), .out(n12243_0));
mux11 mux_7078 (.in({n14344_0, n14334_0, n14308_0, n14298_0, n12160_1, n8251, n8245, n8239, n8233, n8199/**/, n8191}), .out(n12244), .config_in(config_chain[25245:25240]), .config_rst(config_rst)); 
buffer_wire buffer_12244 (.in(n12244), .out(n12244_0));
mux2 mux_7079 (.in({n14826_0, n9211}), .out(n12245), .config_in(config_chain[25246:25246]), .config_rst(config_rst)); 
buffer_wire buffer_12245 (.in(n12245), .out(n12245_0));
mux11 mux_7080 (.in({n14330_0, n14320_0, n14282_1, n14272_1, n12162_1, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12246), .config_in(config_chain[25252:25247]), .config_rst(config_rst)); 
buffer_wire buffer_12246 (.in(n12246), .out(n12246_0));
mux2 mux_7081 (.in({n14828_0/**/, n9214}), .out(n12247), .config_in(config_chain[25253:25253]), .config_rst(config_rst)); 
buffer_wire buffer_12247 (.in(n12247), .out(n12247_0));
mux11 mux_7082 (.in({n14350_0, n14340_0, n14304_0, n14294_0, n12164_1, n8251, n8245, n8239, n8233, n8199, n8191}), .out(n12248), .config_in(config_chain[25259:25254]), .config_rst(config_rst)); 
buffer_wire buffer_12248 (.in(n12248), .out(n12248_0));
mux2 mux_7083 (.in({n14830_0/**/, n9217}), .out(n12249), .config_in(config_chain[25260:25260]), .config_rst(config_rst)); 
buffer_wire buffer_12249 (.in(n12249), .out(n12249_0));
mux13 mux_7084 (.in({n14604_0, n14594_0, n14568_0, n14558_0, n14432_2, n12168_1, n9232, n9226, n9220, n9214, n9181, n9173, n9165}), .out(n12250), .config_in(config_chain[25266:25261]), .config_rst(config_rst)); 
buffer_wire buffer_12250 (.in(n12250), .out(n12250_0));
mux3 mux_7085 (.in({n14834_0, n9223, n9165}), .out(n12251), .config_in(config_chain[25268:25267]), .config_rst(config_rst)); 
buffer_wire buffer_12251 (.in(n12251), .out(n12251_0));
mux13 mux_7086 (.in({n14588_0, n14578_0, n14542_1, n14532_1, n14464_2, n12170_1, n9232, n9226, n9220, n9214, n9181, n9173, n9165}), .out(n12252), .config_in(config_chain[25274:25269]), .config_rst(config_rst)); 
buffer_wire buffer_12252 (.in(n12252), .out(n12252_0));
mux3 mux_7087 (.in({n14836_0/**/, n9226, n9169}), .out(n12253), .config_in(config_chain[25276:25275]), .config_rst(config_rst)); 
buffer_wire buffer_12253 (.in(n12253), .out(n12253_0));
mux13 mux_7088 (.in({n14610_0, n14600_0, n14564_0, n14554_0, n14486_2, n12172_1, n9232, n9226, n9220, n9214, n9181, n9173, n9165}), .out(n12254), .config_in(config_chain[25282:25277]), .config_rst(config_rst)); 
buffer_wire buffer_12254 (.in(n12254), .out(n12254_0));
mux3 mux_7089 (.in({n14838_0, n9229, n9169}), .out(n12255), .config_in(config_chain[25284:25283]), .config_rst(config_rst)); 
buffer_wire buffer_12255 (.in(n12255), .out(n12255_0));
mux13 mux_7090 (.in({n14584_0, n14574_0, n14548_1, n14538_1, n14508_1/**/, n12174_1, n9232, n9226, n9220, n9214, n9181, n9173, n9165}), .out(n12256), .config_in(config_chain[25290:25285]), .config_rst(config_rst)); 
buffer_wire buffer_12256 (.in(n12256), .out(n12256_0));
mux3 mux_7091 (.in({n14840_0, n9229, n9173}), .out(n12257), .config_in(config_chain[25292:25291]), .config_rst(config_rst)); 
buffer_wire buffer_12257 (.in(n12257), .out(n12257_0));
mux13 mux_7092 (.in({n14606_0, n14596_0, n14570_0, n14560_0, n14530_1, n12176_1, n9232, n9226, n9220, n9214, n9181, n9173, n9165}), .out(n12258), .config_in(config_chain[25298:25293]), .config_rst(config_rst)); 
buffer_wire buffer_12258 (.in(n12258), .out(n12258_0));
mux3 mux_7093 (.in({n14842_0, n9232, n9177}), .out(n12259), .config_in(config_chain[25300:25299]), .config_rst(config_rst)); 
buffer_wire buffer_12259 (.in(n12259), .out(n12259_0));
mux12 mux_7094 (.in({n14590_0/**/, n14580_0, n14552_1, n14544_1, n14534_1, n12178_1, n9229, n9223, n9217, n9211, n9177, n9169}), .out(n12260), .config_in(config_chain[25306:25301]), .config_rst(config_rst)); 
buffer_wire buffer_12260 (.in(n12260), .out(n12260_0));
mux2 mux_7095 (.in({n14844_0, n9181}), .out(n12261), .config_in(config_chain[25307:25307]), .config_rst(config_rst)); 
buffer_wire buffer_12261 (.in(n12261), .out(n12261_0));
mux11 mux_7096 (.in({n14612_0, n14602_0, n14566_0, n14556_0, n12180_1, n9229, n9223, n9217, n9211, n9177, n9169}), .out(n12262), .config_in(config_chain[25313:25308]), .config_rst(config_rst)); 
buffer_wire buffer_12262 (.in(n12262), .out(n12262_0));
mux2 mux_7097 (.in({n14846_0/**/, n9211}), .out(n12263), .config_in(config_chain[25314:25314]), .config_rst(config_rst)); 
buffer_wire buffer_12263 (.in(n12263), .out(n12263_0));
mux11 mux_7098 (.in({n14586_0/**/, n14576_0, n14550_1, n14540_1, n12182_1, n9229, n9223, n9217, n9211, n9177, n9169}), .out(n12264), .config_in(config_chain[25320:25315]), .config_rst(config_rst)); 
buffer_wire buffer_12264 (.in(n12264), .out(n12264_0));
mux2 mux_7099 (.in({n14848_0, n9211}), .out(n12265), .config_in(config_chain[25321:25321]), .config_rst(config_rst)); 
buffer_wire buffer_12265 (.in(n12265), .out(n12265_0));
mux11 mux_7100 (.in({n14608_0, n14598_0, n14572_0, n14562_0, n12184_1, n9229, n9223, n9217, n9211, n9177, n9169}), .out(n12266), .config_in(config_chain[25327:25322]), .config_rst(config_rst)); 
buffer_wire buffer_12266 (.in(n12266), .out(n12266_0));
mux2 mux_7101 (.in({n14850_0/**/, n9214}), .out(n12267), .config_in(config_chain[25328:25328]), .config_rst(config_rst)); 
buffer_wire buffer_12267 (.in(n12267), .out(n12267_0));
mux11 mux_7102 (.in({n14592_0, n14582_0/**/, n14546_1, n14536_1, n12186_1, n9229, n9223, n9217, n9211, n9177, n9169}), .out(n12268), .config_in(config_chain[25334:25329]), .config_rst(config_rst)); 
buffer_wire buffer_12268 (.in(n12268), .out(n12268_0));
mux2 mux_7103 (.in({n14852_0, n9217}), .out(n12269), .config_in(config_chain[25335:25335]), .config_rst(config_rst)); 
buffer_wire buffer_12269 (.in(n12269), .out(n12269_0));
mux3 mux_7104 (.in({n9669_0, n564, n25}), .out(n12270), .config_in(config_chain[25337:25336]), .config_rst(config_rst)); 
buffer_wire buffer_12270 (.in(n12270), .out(n12270_0));
mux13 mux_7105 (.in({n12423_1, n10775_1, n10755_0, n10735_1, n10715_0, n10695_1, n870, n862, n854, n187, n181, n175, n169}), .out(n12271), .config_in(config_chain[25343:25338]), .config_rst(config_rst)); 
buffer_wire buffer_12271 (.in(n12271), .out(n12271_0));
mux3 mux_7106 (.in({n9671_0/**/, n564, n25}), .out(n12272), .config_in(config_chain[25345:25344]), .config_rst(config_rst)); 
buffer_wire buffer_12272 (.in(n12272), .out(n12272_0));
mux13 mux_7107 (.in({n12363_1, n10001_2, n9981_0, n9961_0, n9941_0, n9921_0, n576, n568, n560, n43, n37, n31, n25}), .out(n12273), .config_in(config_chain[25351:25346]), .config_rst(config_rst)); 
buffer_wire buffer_12273 (.in(n12273), .out(n12273_0));
mux3 mux_7108 (.in({n9673_0, n564, n25}), .out(n12274), .config_in(config_chain[25353:25352]), .config_rst(config_rst)); 
buffer_wire buffer_12274 (.in(n12274), .out(n12274_0));
mux13 mux_7109 (.in({n12383_1, n10257_1, n10237_1, n10217_0, n10197_1, n10177_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12275), .config_in(config_chain[25359:25354]), .config_rst(config_rst)); 
buffer_wire buffer_12275 (.in(n12275), .out(n12275_0));
mux3 mux_7110 (.in({n9675_1, n564, n25}), .out(n12276), .config_in(config_chain[25361:25360]), .config_rst(config_rst)); 
buffer_wire buffer_12276 (.in(n12276), .out(n12276_0));
mux13 mux_7111 (.in({n12403_1, n10515_1, n10495_0, n10475_0, n10455_0, n10435_0, n772/**/, n764, n756, n139, n133, n127, n121}), .out(n12277), .config_in(config_chain[25367:25362]), .config_rst(config_rst)); 
buffer_wire buffer_12277 (.in(n12277), .out(n12277_0));
mux3 mux_7112 (.in({n9677_0, n568, n25}), .out(n12278), .config_in(config_chain[25369:25368]), .config_rst(config_rst)); 
buffer_wire buffer_12278 (.in(n12278), .out(n12278_0));
mux13 mux_7113 (.in({n12425_1, n10777_1, n10757_0, n10737_0, n10717_0/**/, n10697_0, n870, n862, n854, n187, n181, n175, n169}), .out(n12279), .config_in(config_chain[25375:25370]), .config_rst(config_rst)); 
buffer_wire buffer_12279 (.in(n12279), .out(n12279_0));
mux3 mux_7114 (.in({n9679_0, n568, n28}), .out(n12280), .config_in(config_chain[25377:25376]), .config_rst(config_rst)); 
buffer_wire buffer_12280 (.in(n12280), .out(n12280_0));
mux13 mux_7115 (.in({n12365_1/**/, n10003_2, n9983_0, n9963_1, n9943_0, n9923_1, n576, n568, n560, n43, n37, n31, n25}), .out(n12281), .config_in(config_chain[25383:25378]), .config_rst(config_rst)); 
buffer_wire buffer_12281 (.in(n12281), .out(n12281_0));
mux3 mux_7116 (.in({n9681_0/**/, n568, n28}), .out(n12282), .config_in(config_chain[25385:25384]), .config_rst(config_rst)); 
buffer_wire buffer_12282 (.in(n12282), .out(n12282_0));
mux13 mux_7117 (.in({n12385_1, n10259_2, n10239_0, n10219_0, n10199_0, n10179_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12283), .config_in(config_chain[25391:25386]), .config_rst(config_rst)); 
buffer_wire buffer_12283 (.in(n12283), .out(n12283_0));
mux3 mux_7118 (.in({n9683_1, n568, n28}), .out(n12284), .config_in(config_chain[25393:25392]), .config_rst(config_rst)); 
buffer_wire buffer_12284 (.in(n12284), .out(n12284_0));
mux13 mux_7119 (.in({n12405_1, n10517_1, n10497_1, n10477_0/**/, n10457_1, n10437_0, n772, n764, n756, n139, n133, n127, n121}), .out(n12285), .config_in(config_chain[25399:25394]), .config_rst(config_rst)); 
buffer_wire buffer_12285 (.in(n12285), .out(n12285_0));
mux3 mux_7120 (.in({n9685_0/**/, n568, n28}), .out(n12286), .config_in(config_chain[25401:25400]), .config_rst(config_rst)); 
buffer_wire buffer_12286 (.in(n12286), .out(n12286_0));
mux13 mux_7121 (.in({n12427_1, n10779_1, n10759_1, n10739_0, n10719_1, n10699_0, n870, n862/**/, n854, n187, n181, n175, n169}), .out(n12287), .config_in(config_chain[25407:25402]), .config_rst(config_rst)); 
buffer_wire buffer_12287 (.in(n12287), .out(n12287_0));
mux3 mux_7122 (.in({n9687_0, n572, n28}), .out(n12288), .config_in(config_chain[25409:25408]), .config_rst(config_rst)); 
buffer_wire buffer_12288 (.in(n12288), .out(n12288_0));
mux13 mux_7123 (.in({n12367_1/**/, n10005_2, n9985_0, n9965_0, n9945_0, n9925_0, n576, n568, n560, n43, n37, n31, n25}), .out(n12289), .config_in(config_chain[25415:25410]), .config_rst(config_rst)); 
buffer_wire buffer_12289 (.in(n12289), .out(n12289_0));
mux3 mux_7124 (.in({n9689_0, n572, n31}), .out(n12290), .config_in(config_chain[25417:25416]), .config_rst(config_rst)); 
buffer_wire buffer_12290 (.in(n12290), .out(n12290_0));
mux13 mux_7125 (.in({n12387_1, n10261_2, n10241_0, n10221_1, n10201_0, n10181_1, n674, n666, n658, n91, n85, n79, n73}), .out(n12291), .config_in(config_chain[25423:25418]), .config_rst(config_rst)); 
buffer_wire buffer_12291 (.in(n12291), .out(n12291_0));
mux3 mux_7126 (.in({n9691_1, n572, n31}), .out(n12292), .config_in(config_chain[25425:25424]), .config_rst(config_rst)); 
buffer_wire buffer_12292 (.in(n12292), .out(n12292_0));
mux13 mux_7127 (.in({n12407_1, n10519_2, n10499_0/**/, n10479_0, n10459_0, n10439_0, n772, n764, n756, n139, n133, n127, n121}), .out(n12293), .config_in(config_chain[25431:25426]), .config_rst(config_rst)); 
buffer_wire buffer_12293 (.in(n12293), .out(n12293_0));
mux3 mux_7128 (.in({n9693_0, n572, n31}), .out(n12294), .config_in(config_chain[25433:25432]), .config_rst(config_rst)); 
buffer_wire buffer_12294 (.in(n12294), .out(n12294_0));
mux13 mux_7129 (.in({n12429_1, n10781_2, n10761_0, n10741_0, n10721_0, n10701_0, n870/**/, n862, n854, n187, n181, n175, n169}), .out(n12295), .config_in(config_chain[25439:25434]), .config_rst(config_rst)); 
buffer_wire buffer_12295 (.in(n12295), .out(n12295_0));
mux3 mux_7130 (.in({n9695_0, n572, n31}), .out(n12296), .config_in(config_chain[25441:25440]), .config_rst(config_rst)); 
buffer_wire buffer_12296 (.in(n12296), .out(n12296_0));
mux13 mux_7131 (.in({n12369_1/**/, n10007_2, n9987_1, n9967_0, n9947_1, n9927_0, n576, n568, n560, n43, n37, n31, n25}), .out(n12297), .config_in(config_chain[25447:25442]), .config_rst(config_rst)); 
buffer_wire buffer_12297 (.in(n12297), .out(n12297_0));
mux3 mux_7132 (.in({n9697_0/**/, n576, n31}), .out(n12298), .config_in(config_chain[25449:25448]), .config_rst(config_rst)); 
buffer_wire buffer_12298 (.in(n12298), .out(n12298_0));
mux13 mux_7133 (.in({n12389_1, n10263_2, n10243_0, n10223_0, n10203_0, n10183_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12299), .config_in(config_chain[25455:25450]), .config_rst(config_rst)); 
buffer_wire buffer_12299 (.in(n12299), .out(n12299_0));
mux3 mux_7134 (.in({n9699_1, n576, n34}), .out(n12300), .config_in(config_chain[25457:25456]), .config_rst(config_rst)); 
buffer_wire buffer_12300 (.in(n12300), .out(n12300_0));
mux13 mux_7135 (.in({n12409_1, n10521_2, n10501_0, n10481_1, n10461_0, n10441_1, n772, n764, n756, n139, n133, n127, n121}), .out(n12301), .config_in(config_chain[25463:25458]), .config_rst(config_rst)); 
buffer_wire buffer_12301 (.in(n12301), .out(n12301_0));
mux3 mux_7136 (.in({n9701_0/**/, n576, n34}), .out(n12302), .config_in(config_chain[25465:25464]), .config_rst(config_rst)); 
buffer_wire buffer_12302 (.in(n12302), .out(n12302_0));
mux13 mux_7137 (.in({n12431_1/**/, n10783_2, n10763_0, n10743_1, n10723_0, n10703_1, n870, n862, n854, n187, n181, n175, n169}), .out(n12303), .config_in(config_chain[25471:25466]), .config_rst(config_rst)); 
buffer_wire buffer_12303 (.in(n12303), .out(n12303_0));
mux3 mux_7138 (.in({n9703_0, n576, n34}), .out(n12304), .config_in(config_chain[25473:25472]), .config_rst(config_rst)); 
buffer_wire buffer_12304 (.in(n12304), .out(n12304_0));
mux13 mux_7139 (.in({n12371_1, n10009_2, n9989_0, n9969_0, n9949_0, n9929_0, n576, n568, n560, n43, n37, n31, n25}), .out(n12305), .config_in(config_chain[25479:25474]), .config_rst(config_rst)); 
buffer_wire buffer_12305 (.in(n12305), .out(n12305_0));
mux3 mux_7140 (.in({n9705_0/**/, n576, n34}), .out(n12306), .config_in(config_chain[25481:25480]), .config_rst(config_rst)); 
buffer_wire buffer_12306 (.in(n12306), .out(n12306_0));
mux13 mux_7141 (.in({n12391_1, n10265_2, n10245_1, n10225_0, n10205_1, n10185_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12307), .config_in(config_chain[25487:25482]), .config_rst(config_rst)); 
buffer_wire buffer_12307 (.in(n12307), .out(n12307_0));
mux2 mux_7142 (.in({n9707_1, n34}), .out(n12308), .config_in(config_chain[25488:25488]), .config_rst(config_rst)); 
buffer_wire buffer_12308 (.in(n12308), .out(n12308_0));
mux13 mux_7143 (.in({n12411_1, n10523_2, n10503_0, n10483_0, n10463_0, n10443_0/**/, n772, n764, n756, n139, n133, n127, n121}), .out(n12309), .config_in(config_chain[25494:25489]), .config_rst(config_rst)); 
buffer_wire buffer_12309 (.in(n12309), .out(n12309_0));
mux2 mux_7144 (.in({n9709_0/**/, n37}), .out(n12310), .config_in(config_chain[25495:25495]), .config_rst(config_rst)); 
buffer_wire buffer_12310 (.in(n12310), .out(n12310_0));
mux12 mux_7145 (.in({n12433_1, n10785_2, n10765_0, n10745_0, n10725_0, n10705_0, n866, n858/**/, n190, n184, n178, n172}), .out(n12311), .config_in(config_chain[25501:25496]), .config_rst(config_rst)); 
buffer_wire buffer_12311 (.in(n12311), .out(n12311_0));
mux2 mux_7146 (.in({n9711_0, n37}), .out(n12312), .config_in(config_chain[25502:25502]), .config_rst(config_rst)); 
buffer_wire buffer_12312 (.in(n12312), .out(n12312_0));
mux12 mux_7147 (.in({n12373_1/**/, n10011_2, n9991_0, n9971_1, n9951_0, n9931_1, n572, n564, n46, n40, n34, n28}), .out(n12313), .config_in(config_chain[25508:25503]), .config_rst(config_rst)); 
buffer_wire buffer_12313 (.in(n12313), .out(n12313_0));
mux2 mux_7148 (.in({n9713_0, n37}), .out(n12314), .config_in(config_chain[25509:25509]), .config_rst(config_rst)); 
buffer_wire buffer_12314 (.in(n12314), .out(n12314_0));
mux12 mux_7149 (.in({n12393_1, n10267_2, n10247_0, n10227_0, n10207_0, n10187_0, n670, n662, n94, n88, n82, n76}), .out(n12315), .config_in(config_chain[25515:25510]), .config_rst(config_rst)); 
buffer_wire buffer_12315 (.in(n12315), .out(n12315_0));
mux2 mux_7150 (.in({n9715_1, n37}), .out(n12316), .config_in(config_chain[25516:25516]), .config_rst(config_rst)); 
buffer_wire buffer_12316 (.in(n12316), .out(n12316_0));
mux12 mux_7151 (.in({n12413_1, n10525_2, n10505_1, n10485_0, n10465_1, n10445_0, n768, n760, n142, n136, n130, n124}), .out(n12317), .config_in(config_chain[25522:25517]), .config_rst(config_rst)); 
buffer_wire buffer_12317 (.in(n12317), .out(n12317_0));
mux2 mux_7152 (.in({n9717_0/**/, n37}), .out(n12318), .config_in(config_chain[25523:25523]), .config_rst(config_rst)); 
buffer_wire buffer_12318 (.in(n12318), .out(n12318_0));
mux11 mux_7153 (.in({n12435_1, n10767_1, n10747_0, n10727_1, n10707_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12319), .config_in(config_chain[25529:25524]), .config_rst(config_rst)); 
buffer_wire buffer_12319 (.in(n12319), .out(n12319_0));
mux2 mux_7154 (.in({n9719_0, n40}), .out(n12320), .config_in(config_chain[25530:25530]), .config_rst(config_rst)); 
buffer_wire buffer_12320 (.in(n12320), .out(n12320_0));
mux11 mux_7155 (.in({n12375_1, n9993_0, n9973_0, n9953_0, n9933_0/**/, n572, n564, n46, n40, n34, n28}), .out(n12321), .config_in(config_chain[25536:25531]), .config_rst(config_rst)); 
buffer_wire buffer_12321 (.in(n12321), .out(n12321_0));
mux2 mux_7156 (.in({n9721_0/**/, n40}), .out(n12322), .config_in(config_chain[25537:25537]), .config_rst(config_rst)); 
buffer_wire buffer_12322 (.in(n12322), .out(n12322_0));
mux11 mux_7157 (.in({n12395_1, n10249_0/**/, n10229_1, n10209_0, n10189_1, n670, n662, n94, n88, n82, n76}), .out(n12323), .config_in(config_chain[25543:25538]), .config_rst(config_rst)); 
buffer_wire buffer_12323 (.in(n12323), .out(n12323_0));
mux2 mux_7158 (.in({n9723_1/**/, n40}), .out(n12324), .config_in(config_chain[25544:25544]), .config_rst(config_rst)); 
buffer_wire buffer_12324 (.in(n12324), .out(n12324_0));
mux11 mux_7159 (.in({n12415_1, n10507_0, n10487_0, n10467_0/**/, n10447_0, n768, n760, n142, n136, n130, n124}), .out(n12325), .config_in(config_chain[25550:25545]), .config_rst(config_rst)); 
buffer_wire buffer_12325 (.in(n12325), .out(n12325_0));
mux2 mux_7160 (.in({n9725_0, n40}), .out(n12326), .config_in(config_chain[25551:25551]), .config_rst(config_rst)); 
buffer_wire buffer_12326 (.in(n12326), .out(n12326_0));
mux11 mux_7161 (.in({n12437_1, n10769_0, n10749_0, n10729_0, n10709_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12327), .config_in(config_chain[25557:25552]), .config_rst(config_rst)); 
buffer_wire buffer_12327 (.in(n12327), .out(n12327_0));
mux2 mux_7162 (.in({n9727_0, n40}), .out(n12328), .config_in(config_chain[25558:25558]), .config_rst(config_rst)); 
buffer_wire buffer_12328 (.in(n12328), .out(n12328_0));
mux11 mux_7163 (.in({n12377_1/**/, n9995_1, n9975_0, n9955_1, n9935_0, n572, n564, n46, n40, n34, n28}), .out(n12329), .config_in(config_chain[25564:25559]), .config_rst(config_rst)); 
buffer_wire buffer_12329 (.in(n12329), .out(n12329_0));
mux2 mux_7164 (.in({n9729_0, n43}), .out(n12330), .config_in(config_chain[25565:25565]), .config_rst(config_rst)); 
buffer_wire buffer_12330 (.in(n12330), .out(n12330_0));
mux11 mux_7165 (.in({n12397_1, n10251_0, n10231_0, n10211_0, n10191_0, n670, n662, n94, n88, n82, n76}), .out(n12331), .config_in(config_chain[25571:25566]), .config_rst(config_rst)); 
buffer_wire buffer_12331 (.in(n12331), .out(n12331_0));
mux2 mux_7166 (.in({n9731_1, n43}), .out(n12332), .config_in(config_chain[25572:25572]), .config_rst(config_rst)); 
buffer_wire buffer_12332 (.in(n12332), .out(n12332_0));
mux11 mux_7167 (.in({n12417_1, n10509_0, n10489_1, n10469_0, n10449_1, n768, n760, n142, n136, n130, n124}), .out(n12333), .config_in(config_chain[25578:25573]), .config_rst(config_rst)); 
buffer_wire buffer_12333 (.in(n12333), .out(n12333_0));
mux2 mux_7168 (.in({n9733_0/**/, n43}), .out(n12334), .config_in(config_chain[25579:25579]), .config_rst(config_rst)); 
buffer_wire buffer_12334 (.in(n12334), .out(n12334_0));
mux11 mux_7169 (.in({n12439_1, n10771_0, n10751_1, n10731_0, n10711_1, n866, n858, n190, n184/**/, n178, n172}), .out(n12335), .config_in(config_chain[25585:25580]), .config_rst(config_rst)); 
buffer_wire buffer_12335 (.in(n12335), .out(n12335_0));
mux2 mux_7170 (.in({n9735_0, n43}), .out(n12336), .config_in(config_chain[25586:25586]), .config_rst(config_rst)); 
buffer_wire buffer_12336 (.in(n12336), .out(n12336_0));
mux11 mux_7171 (.in({n12379_1, n9997_0, n9977_0, n9957_0, n9937_0, n572, n564, n46, n40, n34, n28}), .out(n12337), .config_in(config_chain[25592:25587]), .config_rst(config_rst)); 
buffer_wire buffer_12337 (.in(n12337), .out(n12337_0));
mux2 mux_7172 (.in({n9737_0, n43}), .out(n12338), .config_in(config_chain[25593:25593]), .config_rst(config_rst)); 
buffer_wire buffer_12338 (.in(n12338), .out(n12338_0));
mux11 mux_7173 (.in({n12399_1, n10253_1, n10233_0, n10213_1, n10193_0, n670, n662, n94, n88, n82, n76}), .out(n12339), .config_in(config_chain[25599:25594]), .config_rst(config_rst)); 
buffer_wire buffer_12339 (.in(n12339), .out(n12339_0));
mux2 mux_7174 (.in({n9739_1, n46}), .out(n12340), .config_in(config_chain[25600:25600]), .config_rst(config_rst)); 
buffer_wire buffer_12340 (.in(n12340), .out(n12340_0));
mux11 mux_7175 (.in({n12419_1, n10511_0, n10491_0, n10471_0, n10451_0/**/, n768, n760, n142, n136, n130, n124}), .out(n12341), .config_in(config_chain[25606:25601]), .config_rst(config_rst)); 
buffer_wire buffer_12341 (.in(n12341), .out(n12341_0));
mux2 mux_7176 (.in({n9741_0, n46}), .out(n12342), .config_in(config_chain[25607:25607]), .config_rst(config_rst)); 
buffer_wire buffer_12342 (.in(n12342), .out(n12342_0));
mux11 mux_7177 (.in({n12441_1, n10773_0, n10753_0, n10733_0, n10713_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12343), .config_in(config_chain[25613:25608]), .config_rst(config_rst)); 
buffer_wire buffer_12343 (.in(n12343), .out(n12343_0));
mux2 mux_7178 (.in({n9743_0, n46}), .out(n12344), .config_in(config_chain[25614:25614]), .config_rst(config_rst)); 
buffer_wire buffer_12344 (.in(n12344), .out(n12344_0));
mux11 mux_7179 (.in({n12381_1/**/, n9999_0, n9979_1, n9959_0, n9939_1, n572, n564, n46, n40, n34, n28}), .out(n12345), .config_in(config_chain[25620:25615]), .config_rst(config_rst)); 
buffer_wire buffer_12345 (.in(n12345), .out(n12345_0));
mux2 mux_7180 (.in({n9745_0, n46}), .out(n12346), .config_in(config_chain[25621:25621]), .config_rst(config_rst)); 
buffer_wire buffer_12346 (.in(n12346), .out(n12346_0));
mux11 mux_7181 (.in({n12401_1, n10255_0, n10235_0, n10215_0, n10195_0, n670, n662, n94, n88, n82, n76}), .out(n12347), .config_in(config_chain[25627:25622]), .config_rst(config_rst)); 
buffer_wire buffer_12347 (.in(n12347), .out(n12347_0));
mux2 mux_7182 (.in({n9747_2, n46}), .out(n12348), .config_in(config_chain[25628:25628]), .config_rst(config_rst)); 
buffer_wire buffer_12348 (.in(n12348), .out(n12348_0));
mux11 mux_7183 (.in({n12421_1, n10513_1, n10493_0, n10473_1/**/, n10453_0, n768, n760, n142, n136, n130, n124}), .out(n12349), .config_in(config_chain[25634:25629]), .config_rst(config_rst)); 
buffer_wire buffer_12349 (.in(n12349), .out(n12349_0));
mux2 mux_7184 (.in({n9749_2, n560}), .out(n12350), .config_in(config_chain[25635:25635]), .config_rst(config_rst)); 
buffer_wire buffer_12350 (.in(n12350), .out(n12350_0));
mux10 mux_7185 (.in({n12523_0, n11835_0, n11813_1, n11791_0/**/, n11769_0, n1254, n1246, n379, n373, n367}), .out(n12351), .config_in(config_chain[25641:25636]), .config_rst(config_rst)); 
buffer_wire buffer_12351 (.in(n12351), .out(n12351_0));
mux2 mux_7186 (.in({n9751_2, n560}), .out(n12352), .config_in(config_chain[25642:25642]), .config_rst(config_rst)); 
buffer_wire buffer_12352 (.in(n12352), .out(n12352_0));
mux2 mux_7187 (.in({n12017_0/**/, n1344}), .out(n12353), .config_in(config_chain[25643:25643]), .config_rst(config_rst)); 
buffer_wire buffer_12353 (.in(n12353), .out(n12353_0));
mux2 mux_7188 (.in({n9753_2, n560}), .out(n12354), .config_in(config_chain[25644:25644]), .config_rst(config_rst)); 
buffer_wire buffer_12354 (.in(n12354), .out(n12354_0));
mux2 mux_7189 (.in({n12015_0/**/, n1344}), .out(n12355), .config_in(config_chain[25645:25645]), .config_rst(config_rst)); 
buffer_wire buffer_12355 (.in(n12355), .out(n12355_0));
mux2 mux_7190 (.in({n9755_2, n560}), .out(n12356), .config_in(config_chain[25646:25646]), .config_rst(config_rst)); 
buffer_wire buffer_12356 (.in(n12356), .out(n12356_0));
mux2 mux_7191 (.in({n12013_1, n1344}), .out(n12357), .config_in(config_chain[25647:25647]), .config_rst(config_rst)); 
buffer_wire buffer_12357 (.in(n12357), .out(n12357_0));
mux2 mux_7192 (.in({n9757_2, n560}), .out(n12358), .config_in(config_chain[25648:25648]), .config_rst(config_rst)); 
buffer_wire buffer_12358 (.in(n12358), .out(n12358_0));
mux2 mux_7193 (.in({n12011_0/**/, n1344}), .out(n12359), .config_in(config_chain[25649:25649]), .config_rst(config_rst)); 
buffer_wire buffer_12359 (.in(n12359), .out(n12359_0));
mux2 mux_7194 (.in({n9667_1, n564}), .out(n12360), .config_in(config_chain[25650:25650]), .config_rst(config_rst)); 
buffer_wire buffer_12360 (.in(n12360), .out(n12360_0));
mux2 mux_7195 (.in({n12101_1, n1348}), .out(n12361), .config_in(config_chain[25651:25651]), .config_rst(config_rst)); 
buffer_wire buffer_12361 (.in(n12361), .out(n12361_0));
mux13 mux_7196 (.in({n12272_0, n10001_2, n9981_0, n9961_0, n9941_0, n9921_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12362), .config_in(config_chain[25657:25652]), .config_rst(config_rst)); 
buffer_wire buffer_12362 (.in(n12362), .out(n12362_0));
mux13 mux_7197 (.in({n12443_1, n11037_0, n11017_0, n10997_0, n10977_0, n10957_0, n968/**/, n960, n952, n235, n229, n223, n217}), .out(n12363), .config_in(config_chain[25663:25658]), .config_rst(config_rst)); 
buffer_wire buffer_12363 (.in(n12363), .out(n12363_0));
mux13 mux_7198 (.in({n12280_0, n10003_2, n9983_0, n9963_1/**/, n9943_0, n9923_1, n674, n666, n658, n91, n85, n79, n73}), .out(n12364), .config_in(config_chain[25669:25664]), .config_rst(config_rst)); 
buffer_wire buffer_12364 (.in(n12364), .out(n12364_0));
mux13 mux_7199 (.in({n12445_1, n11039_1, n11019_0, n10999_1, n10979_0, n10959_1, n968, n960, n952, n235/**/, n229, n223, n217}), .out(n12365), .config_in(config_chain[25675:25670]), .config_rst(config_rst)); 
buffer_wire buffer_12365 (.in(n12365), .out(n12365_0));
mux13 mux_7200 (.in({n12288_0, n10005_2, n9985_0, n9965_0, n9945_0/**/, n9925_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12366), .config_in(config_chain[25681:25676]), .config_rst(config_rst)); 
buffer_wire buffer_12366 (.in(n12366), .out(n12366_0));
mux13 mux_7201 (.in({n12447_1, n11041_1, n11021_0, n11001_0, n10981_0, n10961_0, n968, n960, n952, n235/**/, n229, n223, n217}), .out(n12367), .config_in(config_chain[25687:25682]), .config_rst(config_rst)); 
buffer_wire buffer_12367 (.in(n12367), .out(n12367_0));
mux13 mux_7202 (.in({n12296_0, n10007_2, n9987_1/**/, n9967_0, n9947_1, n9927_0, n674, n666, n658, n91, n85, n79, n73}), .out(n12368), .config_in(config_chain[25693:25688]), .config_rst(config_rst)); 
buffer_wire buffer_12368 (.in(n12368), .out(n12368_0));
mux13 mux_7203 (.in({n12449_1, n11043_1, n11023_1, n11003_0, n10983_1, n10963_0, n968, n960, n952, n235, n229/**/, n223, n217}), .out(n12369), .config_in(config_chain[25699:25694]), .config_rst(config_rst)); 
buffer_wire buffer_12369 (.in(n12369), .out(n12369_0));
mux13 mux_7204 (.in({n12304_0, n10009_2, n9989_0, n9969_0, n9949_0, n9929_0/**/, n674, n666, n658, n91, n85, n79, n73}), .out(n12370), .config_in(config_chain[25705:25700]), .config_rst(config_rst)); 
buffer_wire buffer_12370 (.in(n12370), .out(n12370_0));
mux13 mux_7205 (.in({n12451_1, n11045_2, n11025_0, n11005_0, n10985_0, n10965_0, n968, n960, n952, n235, n229/**/, n223, n217}), .out(n12371), .config_in(config_chain[25711:25706]), .config_rst(config_rst)); 
buffer_wire buffer_12371 (.in(n12371), .out(n12371_0));
mux12 mux_7206 (.in({n12312_0, n10011_2, n9991_0, n9971_1, n9951_0, n9931_1/**/, n670, n662, n94, n88, n82, n76}), .out(n12372), .config_in(config_chain[25717:25712]), .config_rst(config_rst)); 
buffer_wire buffer_12372 (.in(n12372), .out(n12372_0));
mux12 mux_7207 (.in({n12453_1, n11047_2, n11027_0, n11007_1, n10987_0, n10967_1, n964, n956, n238, n232, n226/**/, n220}), .out(n12373), .config_in(config_chain[25723:25718]), .config_rst(config_rst)); 
buffer_wire buffer_12373 (.in(n12373), .out(n12373_0));
mux11 mux_7208 (.in({n12320_0, n9993_0, n9973_0, n9953_0/**/, n9933_0, n670, n662, n94, n88, n82, n76}), .out(n12374), .config_in(config_chain[25729:25724]), .config_rst(config_rst)); 
buffer_wire buffer_12374 (.in(n12374), .out(n12374_0));
mux11 mux_7209 (.in({n12455_1, n11029_0, n11009_0, n10989_0, n10969_0, n964, n956, n238, n232/**/, n226, n220}), .out(n12375), .config_in(config_chain[25735:25730]), .config_rst(config_rst)); 
buffer_wire buffer_12375 (.in(n12375), .out(n12375_0));
mux11 mux_7210 (.in({n12328_0, n9995_1, n9975_0, n9955_1, n9935_0/**/, n670, n662, n94, n88, n82, n76}), .out(n12376), .config_in(config_chain[25741:25736]), .config_rst(config_rst)); 
buffer_wire buffer_12376 (.in(n12376), .out(n12376_0));
mux11 mux_7211 (.in({n12457_1, n11031_1, n11011_0, n10991_1, n10971_0, n964, n956, n238, n232/**/, n226, n220}), .out(n12377), .config_in(config_chain[25747:25742]), .config_rst(config_rst)); 
buffer_wire buffer_12377 (.in(n12377), .out(n12377_0));
mux11 mux_7212 (.in({n12336_0, n9997_0, n9977_0, n9957_0/**/, n9937_0, n670, n662, n94, n88, n82, n76}), .out(n12378), .config_in(config_chain[25753:25748]), .config_rst(config_rst)); 
buffer_wire buffer_12378 (.in(n12378), .out(n12378_0));
mux11 mux_7213 (.in({n12459_1, n11033_0, n11013_0, n10993_0, n10973_0, n964, n956, n238, n232, n226/**/, n220}), .out(n12379), .config_in(config_chain[25759:25754]), .config_rst(config_rst)); 
buffer_wire buffer_12379 (.in(n12379), .out(n12379_0));
mux11 mux_7214 (.in({n12344_0, n9999_0, n9979_1, n9959_0/**/, n9939_1, n670, n662, n94, n88, n82, n76}), .out(n12380), .config_in(config_chain[25765:25760]), .config_rst(config_rst)); 
buffer_wire buffer_12380 (.in(n12380), .out(n12380_0));
mux11 mux_7215 (.in({n12461_1, n11035_0, n11015_1, n10995_0, n10975_1, n964, n956, n238/**/, n232, n226, n220}), .out(n12381), .config_in(config_chain[25771:25766]), .config_rst(config_rst)); 
buffer_wire buffer_12381 (.in(n12381), .out(n12381_0));
mux13 mux_7216 (.in({n12274_0, n10257_1, n10237_1, n10217_0, n10197_1, n10177_0/**/, n772, n764, n756, n139, n133, n127, n121}), .out(n12382), .config_in(config_chain[25777:25772]), .config_rst(config_rst)); 
buffer_wire buffer_12382 (.in(n12382), .out(n12382_0));
mux13 mux_7217 (.in({n12463_0, n11301_0, n11281_1/**/, n11261_0, n11241_1, n11221_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12383), .config_in(config_chain[25783:25778]), .config_rst(config_rst)); 
buffer_wire buffer_12383 (.in(n12383), .out(n12383_0));
mux13 mux_7218 (.in({n12282_0, n10259_2, n10239_0/**/, n10219_0, n10199_0, n10179_0, n772, n764, n756, n139, n133, n127, n121}), .out(n12384), .config_in(config_chain[25789:25784]), .config_rst(config_rst)); 
buffer_wire buffer_12384 (.in(n12384), .out(n12384_0));
mux13 mux_7219 (.in({n12465_0, n11303_0, n11283_0, n11263_0/**/, n11243_0, n11223_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12385), .config_in(config_chain[25795:25790]), .config_rst(config_rst)); 
buffer_wire buffer_12385 (.in(n12385), .out(n12385_0));
mux13 mux_7220 (.in({n12290_0, n10261_2, n10241_0, n10221_1, n10201_0/**/, n10181_1, n772, n764, n756, n139, n133, n127, n121}), .out(n12386), .config_in(config_chain[25801:25796]), .config_rst(config_rst)); 
buffer_wire buffer_12386 (.in(n12386), .out(n12386_0));
mux13 mux_7221 (.in({n12467_0, n11305_1, n11285_0, n11265_1, n11245_0, n11225_1, n1066/**/, n1058, n1050, n283, n277, n271, n265}), .out(n12387), .config_in(config_chain[25807:25802]), .config_rst(config_rst)); 
buffer_wire buffer_12387 (.in(n12387), .out(n12387_0));
mux13 mux_7222 (.in({n12298_0, n10263_2, n10243_0, n10223_0, n10203_0, n10183_0/**/, n772, n764, n756, n139, n133, n127, n121}), .out(n12388), .config_in(config_chain[25813:25808]), .config_rst(config_rst)); 
buffer_wire buffer_12388 (.in(n12388), .out(n12388_0));
mux13 mux_7223 (.in({n12469_0, n11307_1, n11287_0, n11267_0/**/, n11247_0, n11227_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12389), .config_in(config_chain[25819:25814]), .config_rst(config_rst)); 
buffer_wire buffer_12389 (.in(n12389), .out(n12389_0));
mux13 mux_7224 (.in({n12306_0/**/, n10265_2, n10245_1, n10225_0, n10205_1, n10185_0, n772, n764, n756, n139, n133, n127, n121}), .out(n12390), .config_in(config_chain[25825:25820]), .config_rst(config_rst)); 
buffer_wire buffer_12390 (.in(n12390), .out(n12390_0));
mux13 mux_7225 (.in({n12471_0, n11309_1, n11289_1, n11269_0, n11249_1, n11229_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12391), .config_in(config_chain[25831:25826]), .config_rst(config_rst)); 
buffer_wire buffer_12391 (.in(n12391), .out(n12391_0));
mux12 mux_7226 (.in({n12314_0, n10267_2, n10247_0, n10227_0, n10207_0/**/, n10187_0, n768, n760, n142, n136, n130, n124}), .out(n12392), .config_in(config_chain[25837:25832]), .config_rst(config_rst)); 
buffer_wire buffer_12392 (.in(n12392), .out(n12392_0));
mux12 mux_7227 (.in({n12473_0, n11311_2, n11291_0, n11271_0, n11251_0/**/, n11231_0, n1062, n1054, n286, n280, n274, n268}), .out(n12393), .config_in(config_chain[25843:25838]), .config_rst(config_rst)); 
buffer_wire buffer_12393 (.in(n12393), .out(n12393_0));
mux11 mux_7228 (.in({n12322_0, n10249_0/**/, n10229_1, n10209_0, n10189_1, n768, n760, n142, n136, n130, n124}), .out(n12394), .config_in(config_chain[25849:25844]), .config_rst(config_rst)); 
buffer_wire buffer_12394 (.in(n12394), .out(n12394_0));
mux11 mux_7229 (.in({n12475_0/**/, n11293_0, n11273_1, n11253_0, n11233_1, n1062, n1054, n286, n280, n274, n268}), .out(n12395), .config_in(config_chain[25855:25850]), .config_rst(config_rst)); 
buffer_wire buffer_12395 (.in(n12395), .out(n12395_0));
mux11 mux_7230 (.in({n12330_0, n10251_0, n10231_0, n10211_0, n10191_0/**/, n768, n760, n142, n136, n130, n124}), .out(n12396), .config_in(config_chain[25861:25856]), .config_rst(config_rst)); 
buffer_wire buffer_12396 (.in(n12396), .out(n12396_0));
mux11 mux_7231 (.in({n12477_0, n11295_0, n11275_0, n11255_0, n11235_0, n1062, n1054, n286, n280, n274, n268}), .out(n12397), .config_in(config_chain[25867:25862]), .config_rst(config_rst)); 
buffer_wire buffer_12397 (.in(n12397), .out(n12397_0));
mux11 mux_7232 (.in({n12338_0, n10253_1/**/, n10233_0, n10213_1, n10193_0, n768, n760, n142, n136, n130, n124}), .out(n12398), .config_in(config_chain[25873:25868]), .config_rst(config_rst)); 
buffer_wire buffer_12398 (.in(n12398), .out(n12398_0));
mux11 mux_7233 (.in({n12479_0, n11297_1, n11277_0/**/, n11257_1, n11237_0, n1062, n1054, n286, n280, n274, n268}), .out(n12399), .config_in(config_chain[25879:25874]), .config_rst(config_rst)); 
buffer_wire buffer_12399 (.in(n12399), .out(n12399_0));
mux11 mux_7234 (.in({n12346_0, n10255_0/**/, n10235_0, n10215_0, n10195_0, n768, n760, n142, n136, n130, n124}), .out(n12400), .config_in(config_chain[25885:25880]), .config_rst(config_rst)); 
buffer_wire buffer_12400 (.in(n12400), .out(n12400_0));
mux11 mux_7235 (.in({n12481_0, n11299_0, n11279_0, n11259_0, n11239_0/**/, n1062, n1054, n286, n280, n274, n268}), .out(n12401), .config_in(config_chain[25891:25886]), .config_rst(config_rst)); 
buffer_wire buffer_12401 (.in(n12401), .out(n12401_0));
mux13 mux_7236 (.in({n12276_0, n10515_1, n10495_0, n10475_0, n10455_0, n10435_0/**/, n870, n862, n854, n187, n181, n175, n169}), .out(n12402), .config_in(config_chain[25897:25892]), .config_rst(config_rst)); 
buffer_wire buffer_12402 (.in(n12402), .out(n12402_0));
mux13 mux_7237 (.in({n12483_0, n11565_0, n11545_0, n11525_0, n11505_0, n11485_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12403), .config_in(config_chain[25903:25898]), .config_rst(config_rst)); 
buffer_wire buffer_12403 (.in(n12403), .out(n12403_0));
mux13 mux_7238 (.in({n12284_0, n10517_1, n10497_1, n10477_0, n10457_1, n10437_0/**/, n870, n862, n854, n187, n181, n175, n169}), .out(n12404), .config_in(config_chain[25909:25904]), .config_rst(config_rst)); 
buffer_wire buffer_12404 (.in(n12404), .out(n12404_0));
mux13 mux_7239 (.in({n12485_0, n11567_0/**/, n11547_1, n11527_0, n11507_1, n11487_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12405), .config_in(config_chain[25915:25910]), .config_rst(config_rst)); 
buffer_wire buffer_12405 (.in(n12405), .out(n12405_0));
mux13 mux_7240 (.in({n12292_0, n10519_2, n10499_0, n10479_0, n10459_0/**/, n10439_0, n870, n862, n854, n187, n181, n175, n169}), .out(n12406), .config_in(config_chain[25921:25916]), .config_rst(config_rst)); 
buffer_wire buffer_12406 (.in(n12406), .out(n12406_0));
mux13 mux_7241 (.in({n12487_0, n11569_0, n11549_0, n11529_0, n11509_0/**/, n11489_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12407), .config_in(config_chain[25927:25922]), .config_rst(config_rst)); 
buffer_wire buffer_12407 (.in(n12407), .out(n12407_0));
mux13 mux_7242 (.in({n12300_0, n10521_2, n10501_0, n10481_1, n10461_0, n10441_1/**/, n870, n862, n854, n187, n181, n175, n169}), .out(n12408), .config_in(config_chain[25933:25928]), .config_rst(config_rst)); 
buffer_wire buffer_12408 (.in(n12408), .out(n12408_0));
mux13 mux_7243 (.in({n12489_0, n11571_1, n11551_0, n11531_1, n11511_0, n11491_1, n1164/**/, n1156, n1148, n331, n325, n319, n313}), .out(n12409), .config_in(config_chain[25939:25934]), .config_rst(config_rst)); 
buffer_wire buffer_12409 (.in(n12409), .out(n12409_0));
mux13 mux_7244 (.in({n12308_0, n10523_2, n10503_0, n10483_0, n10463_0, n10443_0/**/, n870, n862, n854, n187, n181, n175, n169}), .out(n12410), .config_in(config_chain[25945:25940]), .config_rst(config_rst)); 
buffer_wire buffer_12410 (.in(n12410), .out(n12410_0));
mux13 mux_7245 (.in({n12491_0, n11573_1, n11553_0, n11533_0, n11513_0/**/, n11493_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12411), .config_in(config_chain[25951:25946]), .config_rst(config_rst)); 
buffer_wire buffer_12411 (.in(n12411), .out(n12411_0));
mux12 mux_7246 (.in({n12316_0, n10525_2, n10505_1, n10485_0, n10465_1, n10445_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12412), .config_in(config_chain[25957:25952]), .config_rst(config_rst)); 
buffer_wire buffer_12412 (.in(n12412), .out(n12412_0));
mux12 mux_7247 (.in({n12493_0, n11575_1, n11555_1, n11535_0, n11515_1, n11495_0, n1160, n1152, n334, n328, n322, n316}), .out(n12413), .config_in(config_chain[25963:25958]), .config_rst(config_rst)); 
buffer_wire buffer_12413 (.in(n12413), .out(n12413_0));
mux11 mux_7248 (.in({n12324_0, n10507_0, n10487_0, n10467_0, n10447_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12414), .config_in(config_chain[25969:25964]), .config_rst(config_rst)); 
buffer_wire buffer_12414 (.in(n12414), .out(n12414_0));
mux11 mux_7249 (.in({n12495_0/**/, n11557_0, n11537_0, n11517_0, n11497_0, n1160, n1152, n334, n328, n322, n316}), .out(n12415), .config_in(config_chain[25975:25970]), .config_rst(config_rst)); 
buffer_wire buffer_12415 (.in(n12415), .out(n12415_0));
mux11 mux_7250 (.in({n12332_0, n10509_0, n10489_1, n10469_0, n10449_1, n866, n858/**/, n190, n184, n178, n172}), .out(n12416), .config_in(config_chain[25981:25976]), .config_rst(config_rst)); 
buffer_wire buffer_12416 (.in(n12416), .out(n12416_0));
mux11 mux_7251 (.in({n12497_0, n11559_0, n11539_1, n11519_0, n11499_1/**/, n1160, n1152, n334, n328, n322, n316}), .out(n12417), .config_in(config_chain[25987:25982]), .config_rst(config_rst)); 
buffer_wire buffer_12417 (.in(n12417), .out(n12417_0));
mux11 mux_7252 (.in({n12340_0, n10511_0, n10491_0, n10471_0, n10451_0, n866, n858, n190, n184/**/, n178, n172}), .out(n12418), .config_in(config_chain[25993:25988]), .config_rst(config_rst)); 
buffer_wire buffer_12418 (.in(n12418), .out(n12418_0));
mux11 mux_7253 (.in({n12499_0, n11561_0, n11541_0, n11521_0/**/, n11501_0, n1160, n1152, n334, n328, n322, n316}), .out(n12419), .config_in(config_chain[25999:25994]), .config_rst(config_rst)); 
buffer_wire buffer_12419 (.in(n12419), .out(n12419_0));
mux11 mux_7254 (.in({n12348_0, n10513_1, n10493_0, n10473_1, n10453_0, n866, n858/**/, n190, n184, n178, n172}), .out(n12420), .config_in(config_chain[26005:26000]), .config_rst(config_rst)); 
buffer_wire buffer_12420 (.in(n12420), .out(n12420_0));
mux11 mux_7255 (.in({n12501_0, n11563_1, n11543_0/**/, n11523_1, n11503_0, n1160, n1152, n334, n328, n322, n316}), .out(n12421), .config_in(config_chain[26011:26006]), .config_rst(config_rst)); 
buffer_wire buffer_12421 (.in(n12421), .out(n12421_0));
mux13 mux_7256 (.in({n12270_1, n10775_1, n10755_0, n10735_1, n10715_0, n10695_1, n968, n960, n952, n235, n229/**/, n223, n217}), .out(n12422), .config_in(config_chain[26017:26012]), .config_rst(config_rst)); 
buffer_wire buffer_12422 (.in(n12422), .out(n12422_0));
mux12 mux_7257 (.in({n12503_0, n11837_1, n11815_0/**/, n11793_0, n11771_0, n11749_1, n1258, n1246, n379, n373, n367, n361}), .out(n12423), .config_in(config_chain[26023:26018]), .config_rst(config_rst)); 
buffer_wire buffer_12423 (.in(n12423), .out(n12423_0));
mux13 mux_7258 (.in({n12278_1, n10777_1, n10757_0, n10737_0, n10717_0, n10697_0/**/, n968, n960, n952, n235, n229, n223, n217}), .out(n12424), .config_in(config_chain[26029:26024]), .config_rst(config_rst)); 
buffer_wire buffer_12424 (.in(n12424), .out(n12424_0));
mux12 mux_7259 (.in({n12505_0, n11839_1, n11817_0, n11795_0, n11773_1, n11751_0/**/, n1258, n1250, n379, n373, n367, n361}), .out(n12425), .config_in(config_chain[26035:26030]), .config_rst(config_rst)); 
buffer_wire buffer_12425 (.in(n12425), .out(n12425_0));
mux13 mux_7260 (.in({n12286_1, n10779_1, n10759_1, n10739_0, n10719_1, n10699_0, n968, n960, n952, n235/**/, n229, n223, n217}), .out(n12426), .config_in(config_chain[26041:26036]), .config_rst(config_rst)); 
buffer_wire buffer_12426 (.in(n12426), .out(n12426_0));
mux11 mux_7261 (.in({n12507_0, n11819_0, n11797_1, n11775_0, n11753_0/**/, n1258, n1250, n382, n373, n367, n361}), .out(n12427), .config_in(config_chain[26047:26042]), .config_rst(config_rst)); 
buffer_wire buffer_12427 (.in(n12427), .out(n12427_0));
mux13 mux_7262 (.in({n12294_1, n10781_2, n10761_0, n10741_0, n10721_0, n10701_0, n968, n960, n952, n235/**/, n229, n223, n217}), .out(n12428), .config_in(config_chain[26053:26048]), .config_rst(config_rst)); 
buffer_wire buffer_12428 (.in(n12428), .out(n12428_0));
mux11 mux_7263 (.in({n12509_0, n11821_1, n11799_0, n11777_0, n11755_0, n1258/**/, n1250, n382, n376, n367, n361}), .out(n12429), .config_in(config_chain[26059:26054]), .config_rst(config_rst)); 
buffer_wire buffer_12429 (.in(n12429), .out(n12429_0));
mux13 mux_7264 (.in({n12302_1, n10783_2, n10763_0, n10743_1, n10723_0, n10703_1, n968, n960, n952, n235, n229/**/, n223, n217}), .out(n12430), .config_in(config_chain[26065:26060]), .config_rst(config_rst)); 
buffer_wire buffer_12430 (.in(n12430), .out(n12430_0));
mux11 mux_7265 (.in({n12511_0, n11823_0, n11801_0/**/, n11779_0, n11757_1, n1258, n1250, n382, n376, n370, n361}), .out(n12431), .config_in(config_chain[26071:26066]), .config_rst(config_rst)); 
buffer_wire buffer_12431 (.in(n12431), .out(n12431_0));
mux12 mux_7266 (.in({n12310_1, n10785_2, n10765_0, n10745_0, n10725_0, n10705_0, n964, n956, n238, n232, n226/**/, n220}), .out(n12432), .config_in(config_chain[26077:26072]), .config_rst(config_rst)); 
buffer_wire buffer_12432 (.in(n12432), .out(n12432_0));
mux11 mux_7267 (.in({n12513_0, n11825_0, n11803_0, n11781_1, n11759_0, n1262, n1250, n382, n376, n370, n364}), .out(n12433), .config_in(config_chain[26083:26078]), .config_rst(config_rst)); 
buffer_wire buffer_12433 (.in(n12433), .out(n12433_0));
mux11 mux_7268 (.in({n12318_1, n10767_1, n10747_0, n10727_1, n10707_0, n964, n956, n238, n232, n226/**/, n220}), .out(n12434), .config_in(config_chain[26089:26084]), .config_rst(config_rst)); 
buffer_wire buffer_12434 (.in(n12434), .out(n12434_0));
mux11 mux_7269 (.in({n12515_0, n11827_0, n11805_1, n11783_0, n11761_0, n1262, n1254/**/, n382, n376, n370, n364}), .out(n12435), .config_in(config_chain[26095:26090]), .config_rst(config_rst)); 
buffer_wire buffer_12435 (.in(n12435), .out(n12435_0));
mux11 mux_7270 (.in({n12326_1, n10769_0, n10749_0, n10729_0, n10709_0, n964, n956, n238/**/, n232, n226, n220}), .out(n12436), .config_in(config_chain[26101:26096]), .config_rst(config_rst)); 
buffer_wire buffer_12436 (.in(n12436), .out(n12436_0));
mux11 mux_7271 (.in({n12517_0/**/, n11829_2, n11807_0, n11785_0, n11763_0, n1262, n1254, n1246, n376, n370, n364}), .out(n12437), .config_in(config_chain[26107:26102]), .config_rst(config_rst)); 
buffer_wire buffer_12437 (.in(n12437), .out(n12437_0));
mux11 mux_7272 (.in({n12334_1, n10771_0, n10751_1, n10731_0, n10711_1, n964, n956, n238, n232/**/, n226, n220}), .out(n12438), .config_in(config_chain[26113:26108]), .config_rst(config_rst)); 
buffer_wire buffer_12438 (.in(n12438), .out(n12438_0));
mux11 mux_7273 (.in({n12519_0, n11831_0, n11809_0, n11787_0, n11765_1, n1262, n1254, n1246, n379, n370, n364}), .out(n12439), .config_in(config_chain[26119:26114]), .config_rst(config_rst)); 
buffer_wire buffer_12439 (.in(n12439), .out(n12439_0));
mux11 mux_7274 (.in({n12342_1, n10773_0, n10753_0, n10733_0, n10713_0, n964, n956, n238/**/, n232, n226, n220}), .out(n12440), .config_in(config_chain[26125:26120]), .config_rst(config_rst)); 
buffer_wire buffer_12440 (.in(n12440), .out(n12440_0));
mux11 mux_7275 (.in({n12521_0, n11833_0, n11811_0, n11789_1, n11767_0/**/, n1262, n1254, n1246, n379, n373, n364}), .out(n12441), .config_in(config_chain[26131:26126]), .config_rst(config_rst)); 
buffer_wire buffer_12441 (.in(n12441), .out(n12441_0));
mux13 mux_7276 (.in({n12362_1, n11037_0/**/, n11017_0, n10997_0, n10977_0, n10957_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12442), .config_in(config_chain[26137:26132]), .config_rst(config_rst)); 
buffer_wire buffer_12442 (.in(n12442), .out(n12442_0));
mux3 mux_7277 (.in({n12097_0, n1348, n409}), .out(n12443), .config_in(config_chain[26139:26138]), .config_rst(config_rst)); 
buffer_wire buffer_12443 (.in(n12443), .out(n12443_0));
mux13 mux_7278 (.in({n12364_1, n11039_1, n11019_0, n10999_1/**/, n10979_0, n10959_1, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12444), .config_in(config_chain[26145:26140]), .config_rst(config_rst)); 
buffer_wire buffer_12444 (.in(n12444), .out(n12444_0));
mux3 mux_7279 (.in({n12089_0, n1352, n412}), .out(n12445), .config_in(config_chain[26147:26146]), .config_rst(config_rst)); 
buffer_wire buffer_12445 (.in(n12445), .out(n12445_0));
mux13 mux_7280 (.in({n12366_1, n11041_1, n11021_0/**/, n11001_0, n10981_0, n10961_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12446), .config_in(config_chain[26153:26148]), .config_rst(config_rst)); 
buffer_wire buffer_12446 (.in(n12446), .out(n12446_0));
mux3 mux_7281 (.in({n12081_0/**/, n1356, n412}), .out(n12447), .config_in(config_chain[26155:26154]), .config_rst(config_rst)); 
buffer_wire buffer_12447 (.in(n12447), .out(n12447_0));
mux13 mux_7282 (.in({n12368_1/**/, n11043_1, n11023_1, n11003_0, n10983_1, n10963_0, n1066, n1058, n1050, n283, n277, n271, n265}), .out(n12448), .config_in(config_chain[26161:26156]), .config_rst(config_rst)); 
buffer_wire buffer_12448 (.in(n12448), .out(n12448_0));
mux3 mux_7283 (.in({n12073_0, n1356, n415}), .out(n12449), .config_in(config_chain[26163:26162]), .config_rst(config_rst)); 
buffer_wire buffer_12449 (.in(n12449), .out(n12449_0));
mux13 mux_7284 (.in({n12370_1, n11045_2, n11025_0, n11005_0, n10985_0, n10965_0, n1066, n1058/**/, n1050, n283, n277, n271, n265}), .out(n12450), .config_in(config_chain[26169:26164]), .config_rst(config_rst)); 
buffer_wire buffer_12450 (.in(n12450), .out(n12450_0));
mux3 mux_7285 (.in({n12065_0/**/, n1360, n418}), .out(n12451), .config_in(config_chain[26171:26170]), .config_rst(config_rst)); 
buffer_wire buffer_12451 (.in(n12451), .out(n12451_0));
mux12 mux_7286 (.in({n12372_1, n11047_2, n11027_0/**/, n11007_1, n10987_0, n10967_1, n1062, n1054, n286, n280, n274, n268}), .out(n12452), .config_in(config_chain[26177:26172]), .config_rst(config_rst)); 
buffer_wire buffer_12452 (.in(n12452), .out(n12452_0));
mux2 mux_7287 (.in({n12057_0, n421}), .out(n12453), .config_in(config_chain[26178:26178]), .config_rst(config_rst)); 
buffer_wire buffer_12453 (.in(n12453), .out(n12453_0));
mux11 mux_7288 (.in({n12374_1, n11029_0, n11009_0/**/, n10989_0, n10969_0, n1062, n1054, n286, n280, n274, n268}), .out(n12454), .config_in(config_chain[26184:26179]), .config_rst(config_rst)); 
buffer_wire buffer_12454 (.in(n12454), .out(n12454_0));
mux2 mux_7289 (.in({n12049_0, n424}), .out(n12455), .config_in(config_chain[26185:26185]), .config_rst(config_rst)); 
buffer_wire buffer_12455 (.in(n12455), .out(n12455_0));
mux11 mux_7290 (.in({n12376_1, n11031_1, n11011_0, n10991_1/**/, n10971_0, n1062, n1054, n286, n280, n274, n268}), .out(n12456), .config_in(config_chain[26191:26186]), .config_rst(config_rst)); 
buffer_wire buffer_12456 (.in(n12456), .out(n12456_0));
mux2 mux_7291 (.in({n12041_0, n424}), .out(n12457), .config_in(config_chain[26192:26192]), .config_rst(config_rst)); 
buffer_wire buffer_12457 (.in(n12457), .out(n12457_0));
mux11 mux_7292 (.in({n12378_1, n11033_0/**/, n11013_0, n10993_0, n10973_0, n1062, n1054, n286, n280, n274, n268}), .out(n12458), .config_in(config_chain[26198:26193]), .config_rst(config_rst)); 
buffer_wire buffer_12458 (.in(n12458), .out(n12458_0));
mux2 mux_7293 (.in({n12033_0, n427}), .out(n12459), .config_in(config_chain[26199:26199]), .config_rst(config_rst)); 
buffer_wire buffer_12459 (.in(n12459), .out(n12459_0));
mux11 mux_7294 (.in({n12380_1, n11035_0, n11015_1, n10995_0/**/, n10975_1, n1062, n1054, n286, n280, n274, n268}), .out(n12460), .config_in(config_chain[26205:26200]), .config_rst(config_rst)); 
buffer_wire buffer_12460 (.in(n12460), .out(n12460_0));
mux2 mux_7295 (.in({n12025_0, n430}), .out(n12461), .config_in(config_chain[26206:26206]), .config_rst(config_rst)); 
buffer_wire buffer_12461 (.in(n12461), .out(n12461_0));
mux13 mux_7296 (.in({n12382_1, n11301_0/**/, n11281_1, n11261_0, n11241_1, n11221_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12462), .config_in(config_chain[26212:26207]), .config_rst(config_rst)); 
buffer_wire buffer_12462 (.in(n12462), .out(n12462_0));
mux3 mux_7297 (.in({n12095_0, n1348, n409}), .out(n12463), .config_in(config_chain[26214:26213]), .config_rst(config_rst)); 
buffer_wire buffer_12463 (.in(n12463), .out(n12463_0));
mux13 mux_7298 (.in({n12384_1, n11303_0, n11283_0, n11263_0, n11243_0, n11223_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12464), .config_in(config_chain[26220:26215]), .config_rst(config_rst)); 
buffer_wire buffer_12464 (.in(n12464), .out(n12464_0));
mux3 mux_7299 (.in({n12087_0, n1352, n412}), .out(n12465), .config_in(config_chain[26222:26221]), .config_rst(config_rst)); 
buffer_wire buffer_12465 (.in(n12465), .out(n12465_0));
mux13 mux_7300 (.in({n12386_1/**/, n11305_1, n11285_0, n11265_1, n11245_0, n11225_1, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12466), .config_in(config_chain[26228:26223]), .config_rst(config_rst)); 
buffer_wire buffer_12466 (.in(n12466), .out(n12466_0));
mux3 mux_7301 (.in({n12079_0, n1356, n415}), .out(n12467), .config_in(config_chain[26230:26229]), .config_rst(config_rst)); 
buffer_wire buffer_12467 (.in(n12467), .out(n12467_0));
mux13 mux_7302 (.in({n12388_1, n11307_1, n11287_0/**/, n11267_0, n11247_0, n11227_0, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12468), .config_in(config_chain[26236:26231]), .config_rst(config_rst)); 
buffer_wire buffer_12468 (.in(n12468), .out(n12468_0));
mux3 mux_7303 (.in({n12071_0, n1360, n415}), .out(n12469), .config_in(config_chain[26238:26237]), .config_rst(config_rst)); 
buffer_wire buffer_12469 (.in(n12469), .out(n12469_0));
mux13 mux_7304 (.in({n12390_1, n11309_1, n11289_1, n11269_0, n11249_1, n11229_0/**/, n1164, n1156, n1148, n331, n325, n319, n313}), .out(n12470), .config_in(config_chain[26244:26239]), .config_rst(config_rst)); 
buffer_wire buffer_12470 (.in(n12470), .out(n12470_0));
mux3 mux_7305 (.in({n12063_0, n1360, n418}), .out(n12471), .config_in(config_chain[26246:26245]), .config_rst(config_rst)); 
buffer_wire buffer_12471 (.in(n12471), .out(n12471_0));
mux12 mux_7306 (.in({n12392_1, n11311_2, n11291_0/**/, n11271_0, n11251_0, n11231_0, n1160, n1152, n334, n328, n322, n316}), .out(n12472), .config_in(config_chain[26252:26247]), .config_rst(config_rst)); 
buffer_wire buffer_12472 (.in(n12472), .out(n12472_0));
mux2 mux_7307 (.in({n12055_0, n421}), .out(n12473), .config_in(config_chain[26253:26253]), .config_rst(config_rst)); 
buffer_wire buffer_12473 (.in(n12473), .out(n12473_0));
mux11 mux_7308 (.in({n12394_1, n11293_0, n11273_1, n11253_0/**/, n11233_1, n1160, n1152, n334, n328, n322, n316}), .out(n12474), .config_in(config_chain[26259:26254]), .config_rst(config_rst)); 
buffer_wire buffer_12474 (.in(n12474), .out(n12474_0));
mux2 mux_7309 (.in({n12047_0/**/, n424}), .out(n12475), .config_in(config_chain[26260:26260]), .config_rst(config_rst)); 
buffer_wire buffer_12475 (.in(n12475), .out(n12475_0));
mux11 mux_7310 (.in({n12396_1, n11295_0, n11275_0, n11255_0, n11235_0, n1160, n1152, n334, n328, n322, n316}), .out(n12476), .config_in(config_chain[26266:26261]), .config_rst(config_rst)); 
buffer_wire buffer_12476 (.in(n12476), .out(n12476_0));
mux2 mux_7311 (.in({n12039_0, n427}), .out(n12477), .config_in(config_chain[26267:26267]), .config_rst(config_rst)); 
buffer_wire buffer_12477 (.in(n12477), .out(n12477_0));
mux11 mux_7312 (.in({n12398_1/**/, n11297_1, n11277_0, n11257_1, n11237_0, n1160, n1152, n334, n328, n322, n316}), .out(n12478), .config_in(config_chain[26273:26268]), .config_rst(config_rst)); 
buffer_wire buffer_12478 (.in(n12478), .out(n12478_0));
mux2 mux_7313 (.in({n12031_0/**/, n427}), .out(n12479), .config_in(config_chain[26274:26274]), .config_rst(config_rst)); 
buffer_wire buffer_12479 (.in(n12479), .out(n12479_0));
mux11 mux_7314 (.in({n12400_1/**/, n11299_0, n11279_0, n11259_0, n11239_0, n1160, n1152, n334, n328, n322, n316}), .out(n12480), .config_in(config_chain[26280:26275]), .config_rst(config_rst)); 
buffer_wire buffer_12480 (.in(n12480), .out(n12480_0));
mux2 mux_7315 (.in({n12023_0/**/, n430}), .out(n12481), .config_in(config_chain[26281:26281]), .config_rst(config_rst)); 
buffer_wire buffer_12481 (.in(n12481), .out(n12481_0));
mux13 mux_7316 (.in({n12402_1, n11565_0, n11545_0/**/, n11525_0, n11505_0, n11485_0, n1262, n1254, n1246, n379, n373, n367, n361}), .out(n12482), .config_in(config_chain[26287:26282]), .config_rst(config_rst)); 
buffer_wire buffer_12482 (.in(n12482), .out(n12482_0));
mux3 mux_7317 (.in({n12093_2, n1348, n409}), .out(n12483), .config_in(config_chain[26289:26288]), .config_rst(config_rst)); 
buffer_wire buffer_12483 (.in(n12483), .out(n12483_0));
mux13 mux_7318 (.in({n12404_1, n11567_0, n11547_1, n11527_0, n11507_1, n11487_0/**/, n1262, n1254, n1246, n379, n373, n367, n361}), .out(n12484), .config_in(config_chain[26295:26290]), .config_rst(config_rst)); 
buffer_wire buffer_12484 (.in(n12484), .out(n12484_0));
mux3 mux_7319 (.in({n12085_1, n1352, n412}), .out(n12485), .config_in(config_chain[26297:26296]), .config_rst(config_rst)); 
buffer_wire buffer_12485 (.in(n12485), .out(n12485_0));
mux13 mux_7320 (.in({n12406_1, n11569_0, n11549_0, n11529_0, n11509_0, n11489_0, n1262/**/, n1254, n1246, n379, n373, n367, n361}), .out(n12486), .config_in(config_chain[26303:26298]), .config_rst(config_rst)); 
buffer_wire buffer_12486 (.in(n12486), .out(n12486_0));
mux3 mux_7321 (.in({n12077_1, n1356, n415}), .out(n12487), .config_in(config_chain[26305:26304]), .config_rst(config_rst)); 
buffer_wire buffer_12487 (.in(n12487), .out(n12487_0));
mux13 mux_7322 (.in({n12408_1, n11571_1, n11551_0, n11531_1/**/, n11511_0, n11491_1, n1262, n1254, n1246, n379, n373, n367, n361}), .out(n12488), .config_in(config_chain[26311:26306]), .config_rst(config_rst)); 
buffer_wire buffer_12488 (.in(n12488), .out(n12488_0));
mux3 mux_7323 (.in({n12069_1, n1360, n418}), .out(n12489), .config_in(config_chain[26313:26312]), .config_rst(config_rst)); 
buffer_wire buffer_12489 (.in(n12489), .out(n12489_0));
mux13 mux_7324 (.in({n12410_1, n11573_1, n11553_0, n11533_0, n11513_0, n11493_0, n1262, n1254, n1246/**/, n379, n373, n367, n361}), .out(n12490), .config_in(config_chain[26319:26314]), .config_rst(config_rst)); 
buffer_wire buffer_12490 (.in(n12490), .out(n12490_0));
mux2 mux_7325 (.in({n12061_1, n418}), .out(n12491), .config_in(config_chain[26320:26320]), .config_rst(config_rst)); 
buffer_wire buffer_12491 (.in(n12491), .out(n12491_0));
mux12 mux_7326 (.in({n12412_1/**/, n11575_1, n11555_1, n11535_0, n11515_1, n11495_0, n1258, n1250, n382, n376, n370, n364}), .out(n12492), .config_in(config_chain[26326:26321]), .config_rst(config_rst)); 
buffer_wire buffer_12492 (.in(n12492), .out(n12492_0));
mux2 mux_7327 (.in({n12053_1, n421}), .out(n12493), .config_in(config_chain[26327:26327]), .config_rst(config_rst)); 
buffer_wire buffer_12493 (.in(n12493), .out(n12493_0));
mux11 mux_7328 (.in({n12414_1, n11557_0/**/, n11537_0, n11517_0, n11497_0, n1258, n1250, n382, n376, n370, n364}), .out(n12494), .config_in(config_chain[26333:26328]), .config_rst(config_rst)); 
buffer_wire buffer_12494 (.in(n12494), .out(n12494_0));
mux2 mux_7329 (.in({n12045_1/**/, n424}), .out(n12495), .config_in(config_chain[26334:26334]), .config_rst(config_rst)); 
buffer_wire buffer_12495 (.in(n12495), .out(n12495_0));
mux11 mux_7330 (.in({n12416_1, n11559_0, n11539_1, n11519_0, n11499_1, n1258, n1250, n382, n376, n370, n364}), .out(n12496), .config_in(config_chain[26340:26335]), .config_rst(config_rst)); 
buffer_wire buffer_12496 (.in(n12496), .out(n12496_0));
mux2 mux_7331 (.in({n12037_1, n427}), .out(n12497), .config_in(config_chain[26341:26341]), .config_rst(config_rst)); 
buffer_wire buffer_12497 (.in(n12497), .out(n12497_0));
mux11 mux_7332 (.in({n12418_1/**/, n11561_0, n11541_0, n11521_0, n11501_0, n1258, n1250, n382, n376, n370, n364}), .out(n12498), .config_in(config_chain[26347:26342]), .config_rst(config_rst)); 
buffer_wire buffer_12498 (.in(n12498), .out(n12498_0));
mux2 mux_7333 (.in({n12029_1, n430}), .out(n12499), .config_in(config_chain[26348:26348]), .config_rst(config_rst)); 
buffer_wire buffer_12499 (.in(n12499), .out(n12499_0));
mux11 mux_7334 (.in({n12420_1, n11563_1, n11543_0, n11523_1, n11503_0, n1258, n1250, n382, n376, n370, n364}), .out(n12500), .config_in(config_chain[26354:26349]), .config_rst(config_rst)); 
buffer_wire buffer_12500 (.in(n12500), .out(n12500_0));
mux2 mux_7335 (.in({n12021_1, n430}), .out(n12501), .config_in(config_chain[26355:26355]), .config_rst(config_rst)); 
buffer_wire buffer_12501 (.in(n12501), .out(n12501_0));
mux12 mux_7336 (.in({n12422_1/**/, n11837_1, n11815_0, n11793_0, n11771_0, n11749_1, n1356, n1344, n427, n421, n415, n409}), .out(n12502), .config_in(config_chain[26361:26356]), .config_rst(config_rst)); 
buffer_wire buffer_12502 (.in(n12502), .out(n12502_0));
mux3 mux_7337 (.in({n12099_0, n1348, n409}), .out(n12503), .config_in(config_chain[26363:26362]), .config_rst(config_rst)); 
buffer_wire buffer_12503 (.in(n12503), .out(n12503_0));
mux12 mux_7338 (.in({n12424_1, n11839_1/**/, n11817_0, n11795_0, n11773_1, n11751_0, n1356, n1348, n427, n421, n415, n409}), .out(n12504), .config_in(config_chain[26369:26364]), .config_rst(config_rst)); 
buffer_wire buffer_12504 (.in(n12504), .out(n12504_0));
mux3 mux_7339 (.in({n12091_2, n1352, n409}), .out(n12505), .config_in(config_chain[26371:26370]), .config_rst(config_rst)); 
buffer_wire buffer_12505 (.in(n12505), .out(n12505_0));
mux11 mux_7340 (.in({n12426_1/**/, n11819_0, n11797_1, n11775_0, n11753_0, n1356, n1348, n430, n421, n415, n409}), .out(n12506), .config_in(config_chain[26377:26372]), .config_rst(config_rst)); 
buffer_wire buffer_12506 (.in(n12506), .out(n12506_0));
mux3 mux_7341 (.in({n12083_0, n1352, n412}), .out(n12507), .config_in(config_chain[26379:26378]), .config_rst(config_rst)); 
buffer_wire buffer_12507 (.in(n12507), .out(n12507_0));
mux11 mux_7342 (.in({n12428_1, n11821_1, n11799_0, n11777_0, n11755_0, n1356, n1348, n430, n424, n415, n409}), .out(n12508), .config_in(config_chain[26385:26380]), .config_rst(config_rst)); 
buffer_wire buffer_12508 (.in(n12508), .out(n12508_0));
mux3 mux_7343 (.in({n12075_0, n1356, n415}), .out(n12509), .config_in(config_chain[26387:26386]), .config_rst(config_rst)); 
buffer_wire buffer_12509 (.in(n12509), .out(n12509_0));
mux11 mux_7344 (.in({n12430_1/**/, n11823_0, n11801_0, n11779_0, n11757_1, n1356, n1348, n430, n424, n418, n409}), .out(n12510), .config_in(config_chain[26393:26388]), .config_rst(config_rst)); 
buffer_wire buffer_12510 (.in(n12510), .out(n12510_0));
mux3 mux_7345 (.in({n12067_0, n1360, n418}), .out(n12511), .config_in(config_chain[26395:26394]), .config_rst(config_rst)); 
buffer_wire buffer_12511 (.in(n12511), .out(n12511_0));
mux11 mux_7346 (.in({n12432_1, n11825_0, n11803_0, n11781_1, n11759_0/**/, n1360, n1348, n430, n424, n418, n412}), .out(n12512), .config_in(config_chain[26401:26396]), .config_rst(config_rst)); 
buffer_wire buffer_12512 (.in(n12512), .out(n12512_0));
mux2 mux_7347 (.in({n12059_0, n421}), .out(n12513), .config_in(config_chain[26402:26402]), .config_rst(config_rst)); 
buffer_wire buffer_12513 (.in(n12513), .out(n12513_0));
mux11 mux_7348 (.in({n12434_1, n11827_0, n11805_1, n11783_0, n11761_0, n1360, n1352, n430, n424, n418, n412}), .out(n12514), .config_in(config_chain[26408:26403]), .config_rst(config_rst)); 
buffer_wire buffer_12514 (.in(n12514), .out(n12514_0));
mux2 mux_7349 (.in({n12051_0, n421}), .out(n12515), .config_in(config_chain[26409:26409]), .config_rst(config_rst)); 
buffer_wire buffer_12515 (.in(n12515), .out(n12515_0));
mux11 mux_7350 (.in({n12436_1/**/, n11829_2, n11807_0, n11785_0, n11763_0, n1360, n1352, n1344, n424, n418, n412}), .out(n12516), .config_in(config_chain[26415:26410]), .config_rst(config_rst)); 
buffer_wire buffer_12516 (.in(n12516), .out(n12516_0));
mux2 mux_7351 (.in({n12043_0/**/, n424}), .out(n12517), .config_in(config_chain[26416:26416]), .config_rst(config_rst)); 
buffer_wire buffer_12517 (.in(n12517), .out(n12517_0));
mux11 mux_7352 (.in({n12438_1, n11831_0/**/, n11809_0, n11787_0, n11765_1, n1360, n1352, n1344, n427, n418, n412}), .out(n12518), .config_in(config_chain[26422:26417]), .config_rst(config_rst)); 
buffer_wire buffer_12518 (.in(n12518), .out(n12518_0));
mux2 mux_7353 (.in({n12035_0, n427}), .out(n12519), .config_in(config_chain[26423:26423]), .config_rst(config_rst)); 
buffer_wire buffer_12519 (.in(n12519), .out(n12519_0));
mux11 mux_7354 (.in({n12440_1/**/, n11833_0, n11811_0, n11789_1, n11767_0, n1360, n1352, n1344, n427, n421, n412}), .out(n12520), .config_in(config_chain[26429:26424]), .config_rst(config_rst)); 
buffer_wire buffer_12520 (.in(n12520), .out(n12520_0));
mux2 mux_7355 (.in({n12027_0, n430}), .out(n12521), .config_in(config_chain[26430:26430]), .config_rst(config_rst)); 
buffer_wire buffer_12521 (.in(n12521), .out(n12521_0));
mux10 mux_7356 (.in({n12350_2, n11835_0, n11813_1, n11791_0, n11769_0, n1352, n1344, n427, n421, n415}), .out(n12522), .config_in(config_chain[26436:26431]), .config_rst(config_rst)); 
buffer_wire buffer_12522 (.in(n12522), .out(n12522_0));
mux2 mux_7357 (.in({n12019_0, n1344}), .out(n12523), .config_in(config_chain[26437:26437]), .config_rst(config_rst)); 
buffer_wire buffer_12523 (.in(n12523), .out(n12523_0));
mux4 mux_7358 (.in({n9667_0, n9666_0, n1554, n558}), .out(n12524), .config_in(config_chain[26439:26438]), .config_rst(config_rst)); 
buffer_wire buffer_12524 (.in(n12524), .out(n12524_0));
mux16 mux_7359 (.in({n12657_1, n10543_1, n10523_2, n10514_0, n10501_0, n10488_0, n10473_0, n10462_0, n10447_0, n10442_0, n10436_0, n1746, n1738, n770, n762, n754}), .out(n12525), .config_in(config_chain[26445:26440]), .config_rst(config_rst)); 
buffer_wire buffer_12525 (.in(n12525), .out(n12525_0));
mux4 mux_7360 (.in({n9759_1/**/, n9668_0, n1554, n558}), .out(n12526), .config_in(config_chain[26447:26446]), .config_rst(config_rst)); 
buffer_wire buffer_12526 (.in(n12526), .out(n12526_0));
mux16 mux_7361 (.in({n12677_1, n10803_1, n10783_2, n10774_0, n10759_0, n10748_0, n10733_0, n10722_0, n10707_0/**/, n10704_0, n10694_0, n1844, n1836, n868, n860, n852}), .out(n12527), .config_in(config_chain[26453:26448]), .config_rst(config_rst)); 
buffer_wire buffer_12527 (.in(n12527), .out(n12527_0));
mux4 mux_7362 (.in({n9671_0, n9670_0, n1554, n558}), .out(n12528), .config_in(config_chain[26455:26454]), .config_rst(config_rst)); 
buffer_wire buffer_12528 (.in(n12528), .out(n12528_0));
mux16 mux_7363 (.in({n12617_1, n10029_1, n10009_2, n10000_0, n9985_0, n9974_0, n9959_0, n9946_0, n9932_0, n9931_0, n9920_0, n1550, n1542, n574, n566, n558}), .out(n12529), .config_in(config_chain[26461:26456]), .config_rst(config_rst)); 
buffer_wire buffer_12529 (.in(n12529), .out(n12529_0));
mux4 mux_7364 (.in({n9673_0/**/, n9672_0, n1554, n558}), .out(n12530), .config_in(config_chain[26463:26462]), .config_rst(config_rst)); 
buffer_wire buffer_12530 (.in(n12530), .out(n12530_0));
mux16 mux_7365 (.in({n12637_1, n10285_1, n10265_2, n10256_0, n10241_0, n10228_0, n10213_0, n10202_0, n10190_0, n10187_0, n10176_0, n1648, n1640, n672, n664, n656}), .out(n12531), .config_in(config_chain[26469:26464]), .config_rst(config_rst)); 
buffer_wire buffer_12531 (.in(n12531), .out(n12531_0));
mux3 mux_7366 (.in({n9675_0, n9674_0/**/, n558}), .out(n12532), .config_in(config_chain[26471:26470]), .config_rst(config_rst)); 
buffer_wire buffer_12532 (.in(n12532), .out(n12532_0));
mux16 mux_7367 (.in({n12659_1, n10541_1, n10525_2, n10516_0, n10503_0, n10492_0, n10477_0, n10464_0, n10450_0/**/, n10449_0, n10438_0, n1746, n1738, n770, n762, n754}), .out(n12533), .config_in(config_chain[26477:26472]), .config_rst(config_rst)); 
buffer_wire buffer_12533 (.in(n12533), .out(n12533_0));
mux3 mux_7368 (.in({n9761_1, n9676_0, n562}), .out(n12534), .config_in(config_chain[26479:26478]), .config_rst(config_rst)); 
buffer_wire buffer_12534 (.in(n12534), .out(n12534_0));
mux16 mux_7369 (.in({n12679_1, n10801_1, n10785_2, n10776_0, n10763_0, n10750_0, n10735_0, n10724_0, n10712_0, n10709_0/**/, n10698_0, n1844, n1836, n868, n860, n852}), .out(n12535), .config_in(config_chain[26485:26480]), .config_rst(config_rst)); 
buffer_wire buffer_12535 (.in(n12535), .out(n12535_0));
mux3 mux_7370 (.in({n9679_0, n9678_0/**/, n562}), .out(n12536), .config_in(config_chain[26487:26486]), .config_rst(config_rst)); 
buffer_wire buffer_12536 (.in(n12536), .out(n12536_0));
mux16 mux_7371 (.in({n12619_1, n10027_1, n10011_2, n10002_0, n9987_0, n9976_0/**/, n9961_0, n9950_0, n9940_0, n9935_0, n9922_0, n1550, n1542, n574, n566, n558}), .out(n12537), .config_in(config_chain[26493:26488]), .config_rst(config_rst)); 
buffer_wire buffer_12537 (.in(n12537), .out(n12537_0));
mux3 mux_7372 (.in({n9681_0, n9680_0, n562}), .out(n12538), .config_in(config_chain[26495:26494]), .config_rst(config_rst)); 
buffer_wire buffer_12538 (.in(n12538), .out(n12538_0));
mux16 mux_7373 (.in({n12639_1, n10283_1, n10267_2, n10258_0, n10243_0, n10232_0, n10217_0, n10204_0, n10198_0, n10189_0, n10178_0, n1648, n1640, n672, n664, n656}), .out(n12539), .config_in(config_chain[26501:26496]), .config_rst(config_rst)); 
buffer_wire buffer_12539 (.in(n12539), .out(n12539_0));
mux3 mux_7374 (.in({n9683_0, n9682_0, n562}), .out(n12540), .config_in(config_chain[26503:26502]), .config_rst(config_rst)); 
buffer_wire buffer_12540 (.in(n12540), .out(n12540_0));
mux15 mux_7375 (.in({n12661_1, n10539_1, n10518_0, n10505_0, n10494_0, n10479_0, n10468_0, n10458_0/**/, n10453_0, n10440_0, n1746, n1738, n770, n762, n754}), .out(n12541), .config_in(config_chain[26509:26504]), .config_rst(config_rst)); 
buffer_wire buffer_12541 (.in(n12541), .out(n12541_0));
mux3 mux_7376 (.in({n9763_1/**/, n9684_0, n562}), .out(n12542), .config_in(config_chain[26511:26510]), .config_rst(config_rst)); 
buffer_wire buffer_12542 (.in(n12542), .out(n12542_0));
mux15 mux_7377 (.in({n12681_1, n10799_1, n10778_0, n10765_0, n10754_0, n10739_0, n10726_0, n10720_0, n10711_0, n10700_0, n1844, n1836, n868, n860, n852}), .out(n12543), .config_in(config_chain[26517:26512]), .config_rst(config_rst)); 
buffer_wire buffer_12543 (.in(n12543), .out(n12543_0));
mux3 mux_7378 (.in({n9687_0, n9686_0, n566}), .out(n12544), .config_in(config_chain[26519:26518]), .config_rst(config_rst)); 
buffer_wire buffer_12544 (.in(n12544), .out(n12544_0));
mux15 mux_7379 (.in({n12621_1, n10025_1, n10004_0, n9991_0, n9978_0, n9963_0, n9952_0, n9948_0/**/, n9937_0, n9926_0, n1550, n1542, n574, n566, n558}), .out(n12545), .config_in(config_chain[26525:26520]), .config_rst(config_rst)); 
buffer_wire buffer_12545 (.in(n12545), .out(n12545_0));
mux3 mux_7380 (.in({n9689_0/**/, n9688_0, n566}), .out(n12546), .config_in(config_chain[26527:26526]), .config_rst(config_rst)); 
buffer_wire buffer_12546 (.in(n12546), .out(n12546_0));
mux15 mux_7381 (.in({n12641_1, n10281_1, n10260_0, n10245_0, n10234_0, n10219_0, n10208_0, n10206_0, n10193_0, n10180_0, n1648/**/, n1640, n672, n664, n656}), .out(n12547), .config_in(config_chain[26533:26528]), .config_rst(config_rst)); 
buffer_wire buffer_12547 (.in(n12547), .out(n12547_0));
mux3 mux_7382 (.in({n9691_0, n9690_0, n566}), .out(n12548), .config_in(config_chain[26535:26534]), .config_rst(config_rst)); 
buffer_wire buffer_12548 (.in(n12548), .out(n12548_0));
mux15 mux_7383 (.in({n12663_1, n10537_1, n10520_0, n10509_0, n10496_0, n10481_0, n10470_0, n10466_0, n10455_0, n10444_0/**/, n1746, n1738, n770, n762, n754}), .out(n12549), .config_in(config_chain[26541:26536]), .config_rst(config_rst)); 
buffer_wire buffer_12549 (.in(n12549), .out(n12549_0));
mux3 mux_7384 (.in({n9765_1, n9692_0, n566}), .out(n12550), .config_in(config_chain[26543:26542]), .config_rst(config_rst)); 
buffer_wire buffer_12550 (.in(n12550), .out(n12550_0));
mux15 mux_7385 (.in({n12683_1/**/, n10797_1, n10780_0, n10767_0, n10756_0, n10741_0, n10730_0, n10728_0, n10715_0, n10702_0, n1844, n1836, n868, n860, n852}), .out(n12551), .config_in(config_chain[26549:26544]), .config_rst(config_rst)); 
buffer_wire buffer_12551 (.in(n12551), .out(n12551_0));
mux3 mux_7386 (.in({n9695_0, n9694_0/**/, n566}), .out(n12552), .config_in(config_chain[26551:26550]), .config_rst(config_rst)); 
buffer_wire buffer_12552 (.in(n12552), .out(n12552_0));
mux15 mux_7387 (.in({n12623_1, n10023_1, n10006_0, n9993_0/**/, n9982_0, n9967_0, n9956_0, n9954_0, n9939_0, n9928_0, n1550, n1542, n574, n566, n558}), .out(n12553), .config_in(config_chain[26557:26552]), .config_rst(config_rst)); 
buffer_wire buffer_12553 (.in(n12553), .out(n12553_0));
mux3 mux_7388 (.in({n9697_0, n9696_0, n570}), .out(n12554), .config_in(config_chain[26559:26558]), .config_rst(config_rst)); 
buffer_wire buffer_12554 (.in(n12554), .out(n12554_0));
mux15 mux_7389 (.in({n12643_1, n10279_1, n10262_0, n10249_0, n10236_0, n10221_0, n10214_0, n10210_0, n10195_0, n10184_0, n1648, n1640, n672, n664, n656}), .out(n12555), .config_in(config_chain[26565:26560]), .config_rst(config_rst)); 
buffer_wire buffer_12555 (.in(n12555), .out(n12555_0));
mux3 mux_7390 (.in({n9699_0/**/, n9698_0, n570}), .out(n12556), .config_in(config_chain[26567:26566]), .config_rst(config_rst)); 
buffer_wire buffer_12556 (.in(n12556), .out(n12556_0));
mux15 mux_7391 (.in({n12665_1, n10535_1, n10522_0, n10511_0, n10500_0, n10485_0, n10474_0, n10472_0, n10457_0, n10446_0, n1746, n1738, n770, n762, n754}), .out(n12557), .config_in(config_chain[26573:26568]), .config_rst(config_rst)); 
buffer_wire buffer_12557 (.in(n12557), .out(n12557_0));
mux3 mux_7392 (.in({n9767_1/**/, n9700_0, n570}), .out(n12558), .config_in(config_chain[26575:26574]), .config_rst(config_rst)); 
buffer_wire buffer_12558 (.in(n12558), .out(n12558_0));
mux15 mux_7393 (.in({n12685_1, n10795_1, n10782_0, n10771_0/**/, n10758_0, n10743_0, n10736_0, n10732_0, n10717_0, n10706_0, n1844, n1836, n868, n860, n852}), .out(n12559), .config_in(config_chain[26581:26576]), .config_rst(config_rst)); 
buffer_wire buffer_12559 (.in(n12559), .out(n12559_0));
mux3 mux_7394 (.in({n9703_0, n9702_0, n570}), .out(n12560), .config_in(config_chain[26583:26582]), .config_rst(config_rst)); 
buffer_wire buffer_12560 (.in(n12560), .out(n12560_0));
mux15 mux_7395 (.in({n12625_1, n10021_1, n10008_0, n9995_0, n9984_0/**/, n9969_0, n9964_0, n9958_0, n9943_0, n9930_0, n1550, n1542, n574, n566, n558}), .out(n12561), .config_in(config_chain[26589:26584]), .config_rst(config_rst)); 
buffer_wire buffer_12561 (.in(n12561), .out(n12561_0));
mux3 mux_7396 (.in({n9705_0, n9704_0, n570}), .out(n12562), .config_in(config_chain[26591:26590]), .config_rst(config_rst)); 
buffer_wire buffer_12562 (.in(n12562), .out(n12562_0));
mux15 mux_7397 (.in({n12645_1, n10277_1, n10264_0, n10251_0, n10240_0, n10225_0, n10222_0, n10212_0, n10197_0, n10186_0, n1648, n1640, n672, n664, n656}), .out(n12563), .config_in(config_chain[26597:26592]), .config_rst(config_rst)); 
buffer_wire buffer_12563 (.in(n12563), .out(n12563_0));
mux3 mux_7398 (.in({n9707_0, n9706_0, n574}), .out(n12564), .config_in(config_chain[26599:26598]), .config_rst(config_rst)); 
buffer_wire buffer_12564 (.in(n12564), .out(n12564_0));
mux15 mux_7399 (.in({n12667_1, n10533_1, n10524_0, n10513_0, n10502_0, n10487_0, n10482_0, n10476_0, n10461_0, n10448_0, n1750, n1742, n1734, n766, n758}), .out(n12565), .config_in(config_chain[26605:26600]), .config_rst(config_rst)); 
buffer_wire buffer_12565 (.in(n12565), .out(n12565_0));
mux3 mux_7400 (.in({n9769_1/**/, n9708_0, n574}), .out(n12566), .config_in(config_chain[26607:26606]), .config_rst(config_rst)); 
buffer_wire buffer_12566 (.in(n12566), .out(n12566_0));
mux15 mux_7401 (.in({n12687_1, n10793_1, n10784_0, n10773_0, n10762_0, n10747_0, n10744_0, n10734_0, n10719_0, n10708_0, n1848, n1840, n1832, n864, n856/**/}), .out(n12567), .config_in(config_chain[26613:26608]), .config_rst(config_rst)); 
buffer_wire buffer_12567 (.in(n12567), .out(n12567_0));
mux3 mux_7402 (.in({n9711_0, n9710_0, n574}), .out(n12568), .config_in(config_chain[26615:26614]), .config_rst(config_rst)); 
buffer_wire buffer_12568 (.in(n12568), .out(n12568_0));
mux15 mux_7403 (.in({n12627_1/**/, n10019_1, n10010_0, n9999_0, n9986_0, n9972_0, n9971_0, n9960_0, n9945_0, n9934_0, n1554, n1546, n1538, n570, n562}), .out(n12569), .config_in(config_chain[26621:26616]), .config_rst(config_rst)); 
buffer_wire buffer_12569 (.in(n12569), .out(n12569_0));
mux3 mux_7404 (.in({n9713_0, n9712_0, n574}), .out(n12570), .config_in(config_chain[26623:26622]), .config_rst(config_rst)); 
buffer_wire buffer_12570 (.in(n12570), .out(n12570_0));
mux15 mux_7405 (.in({n12647_1, n10275_1, n10266_0, n10253_0, n10242_0/**/, n10230_0, n10227_0, n10216_0, n10201_0, n10188_0, n1652, n1644, n1636, n668, n660}), .out(n12571), .config_in(config_chain[26629:26624]), .config_rst(config_rst)); 
buffer_wire buffer_12571 (.in(n12571), .out(n12571_0));
mux3 mux_7406 (.in({n9715_0, n9714_0, n574}), .out(n12572), .config_in(config_chain[26631:26630]), .config_rst(config_rst)); 
buffer_wire buffer_12572 (.in(n12572), .out(n12572_0));
mux15 mux_7407 (.in({n12669_1, n10531_1, n10515_1, n10504_0, n10490_0, n10489_0, n10478_0, n10463_0, n10452_0, n10437_0, n1750/**/, n1742, n1734, n766, n758}), .out(n12573), .config_in(config_chain[26637:26632]), .config_rst(config_rst)); 
buffer_wire buffer_12573 (.in(n12573), .out(n12573_0));
mux3 mux_7408 (.in({n9771_1/**/, n9716_0, n1538}), .out(n12574), .config_in(config_chain[26639:26638]), .config_rst(config_rst)); 
buffer_wire buffer_12574 (.in(n12574), .out(n12574_0));
mux15 mux_7409 (.in({n12689_1, n10791_1, n10775_0, n10764_0, n10752_0, n10749_0, n10738_0, n10723_0, n10710_0, n10695_0, n1848/**/, n1840, n1832, n864, n856}), .out(n12575), .config_in(config_chain[26645:26640]), .config_rst(config_rst)); 
buffer_wire buffer_12575 (.in(n12575), .out(n12575_0));
mux3 mux_7410 (.in({n9719_0, n9718_0, n1538}), .out(n12576), .config_in(config_chain[26647:26646]), .config_rst(config_rst)); 
buffer_wire buffer_12576 (.in(n12576), .out(n12576_0));
mux15 mux_7411 (.in({n12629_1, n10017_1, n10001_1, n9990_0, n9980_0, n9975_0, n9962_0, n9947_0, n9936_0, n9921_0/**/, n1554, n1546, n1538, n570, n562}), .out(n12577), .config_in(config_chain[26653:26648]), .config_rst(config_rst)); 
buffer_wire buffer_12577 (.in(n12577), .out(n12577_0));
mux3 mux_7412 (.in({n9721_0, n9720_0, n1538}), .out(n12578), .config_in(config_chain[26655:26654]), .config_rst(config_rst)); 
buffer_wire buffer_12578 (.in(n12578), .out(n12578_0));
mux15 mux_7413 (.in({n12649_1, n10273_1, n10257_1, n10244_0, n10238_0, n10229_0, n10218_0, n10203_0, n10192_0, n10177_0, n1652, n1644, n1636, n668, n660}), .out(n12579), .config_in(config_chain[26661:26656]), .config_rst(config_rst)); 
buffer_wire buffer_12579 (.in(n12579), .out(n12579_0));
mux3 mux_7414 (.in({n9723_0, n9722_0/**/, n1538}), .out(n12580), .config_in(config_chain[26663:26662]), .config_rst(config_rst)); 
buffer_wire buffer_12580 (.in(n12580), .out(n12580_0));
mux15 mux_7415 (.in({n12671_1, n10529_1, n10517_1, n10508_0, n10498_0, n10493_0, n10480_0, n10465_0, n10454_0, n10439_0, n1750, n1742, n1734, n766, n758}), .out(n12581), .config_in(config_chain[26669:26664]), .config_rst(config_rst)); 
buffer_wire buffer_12581 (.in(n12581), .out(n12581_0));
mux3 mux_7416 (.in({n9773_1, n9724_0, n1538}), .out(n12582), .config_in(config_chain[26671:26670]), .config_rst(config_rst)); 
buffer_wire buffer_12582 (.in(n12582), .out(n12582_0));
mux15 mux_7417 (.in({n12691_1, n10789_1, n10777_1, n10766_0, n10760_0, n10751_0, n10740_0, n10725_0/**/, n10714_0, n10699_0, n1848, n1840, n1832, n864, n856}), .out(n12583), .config_in(config_chain[26677:26672]), .config_rst(config_rst)); 
buffer_wire buffer_12583 (.in(n12583), .out(n12583_0));
mux3 mux_7418 (.in({n9727_0, n9726_0, n1542}), .out(n12584), .config_in(config_chain[26679:26678]), .config_rst(config_rst)); 
buffer_wire buffer_12584 (.in(n12584), .out(n12584_0));
mux15 mux_7419 (.in({n12631_1, n10015_1, n10003_2, n9992_0, n9988_0, n9977_0, n9966_0, n9951_0, n9938_0, n9923_0, n1554, n1546, n1538, n570, n562}), .out(n12585), .config_in(config_chain[26685:26680]), .config_rst(config_rst)); 
buffer_wire buffer_12585 (.in(n12585), .out(n12585_0));
mux3 mux_7420 (.in({n9729_0, n9728_0, n1542}), .out(n12586), .config_in(config_chain[26687:26686]), .config_rst(config_rst)); 
buffer_wire buffer_12586 (.in(n12586), .out(n12586_0));
mux15 mux_7421 (.in({n12651_1, n10271_1, n10259_1, n10248_0, n10246_0, n10233_0, n10220_0, n10205_0/**/, n10194_0, n10179_0, n1652, n1644, n1636, n668, n660}), .out(n12587), .config_in(config_chain[26693:26688]), .config_rst(config_rst)); 
buffer_wire buffer_12587 (.in(n12587), .out(n12587_0));
mux3 mux_7422 (.in({n9731_0/**/, n9730_0, n1542}), .out(n12588), .config_in(config_chain[26695:26694]), .config_rst(config_rst)); 
buffer_wire buffer_12588 (.in(n12588), .out(n12588_0));
mux15 mux_7423 (.in({n12673_1, n10527_1, n10519_1, n10510_0, n10506_0, n10495_0/**/, n10484_0, n10469_0, n10456_0, n10441_0, n1750, n1742, n1734, n766, n758}), .out(n12589), .config_in(config_chain[26701:26696]), .config_rst(config_rst)); 
buffer_wire buffer_12589 (.in(n12589), .out(n12589_0));
mux3 mux_7424 (.in({n9775_1/**/, n9732_0, n1542}), .out(n12590), .config_in(config_chain[26703:26702]), .config_rst(config_rst)); 
buffer_wire buffer_12590 (.in(n12590), .out(n12590_0));
mux15 mux_7425 (.in({n12693_1, n10787_1, n10779_1, n10770_0, n10768_0, n10755_0, n10742_0, n10727_0, n10716_0, n10701_0, n1848, n1840, n1832/**/, n864, n856}), .out(n12591), .config_in(config_chain[26709:26704]), .config_rst(config_rst)); 
buffer_wire buffer_12591 (.in(n12591), .out(n12591_0));
mux3 mux_7426 (.in({n9735_0, n9734_0, n1542}), .out(n12592), .config_in(config_chain[26711:26710]), .config_rst(config_rst)); 
buffer_wire buffer_12592 (.in(n12592), .out(n12592_0));
mux15 mux_7427 (.in({n12633_1, n10013_1, n10005_2, n9996_0, n9994_0, n9979_0, n9968_0, n9953_0, n9942_0, n9927_0, n1554, n1546, n1538, n570, n562}), .out(n12593), .config_in(config_chain[26717:26712]), .config_rst(config_rst)); 
buffer_wire buffer_12593 (.in(n12593), .out(n12593_0));
mux3 mux_7428 (.in({n9737_0, n9736_0, n1546}), .out(n12594), .config_in(config_chain[26719:26718]), .config_rst(config_rst)); 
buffer_wire buffer_12594 (.in(n12594), .out(n12594_0));
mux15 mux_7429 (.in({n12653_1, n10269_1, n10261_2, n10254_0/**/, n10250_0, n10235_0, n10224_0, n10209_0, n10196_0, n10181_0, n1652, n1644, n1636, n668, n660}), .out(n12595), .config_in(config_chain[26725:26720]), .config_rst(config_rst)); 
buffer_wire buffer_12595 (.in(n12595), .out(n12595_0));
mux3 mux_7430 (.in({n9739_0, n9738_0, n1546}), .out(n12596), .config_in(config_chain[26727:26726]), .config_rst(config_rst)); 
buffer_wire buffer_12596 (.in(n12596), .out(n12596_0));
mux15 mux_7431 (.in({n12675_1, n10545_1, n10521_2, n10512_0, n10497_0, n10486_0, n10471_0, n10460_0, n10445_0, n10434_0, n1750, n1742, n1734, n766, n758}), .out(n12597), .config_in(config_chain[26733:26728]), .config_rst(config_rst)); 
buffer_wire buffer_12597 (.in(n12597), .out(n12597_0));
mux3 mux_7432 (.in({n9777_1/**/, n9740_0, n1546}), .out(n12598), .config_in(config_chain[26735:26734]), .config_rst(config_rst)); 
buffer_wire buffer_12598 (.in(n12598), .out(n12598_0));
mux15 mux_7433 (.in({n12695_1, n10805_1, n10781_1, n10772_0, n10757_0, n10746_0, n10731_0, n10718_0, n10703_0, n10696_0, n1848, n1840, n1832, n864, n856/**/}), .out(n12599), .config_in(config_chain[26741:26736]), .config_rst(config_rst)); 
buffer_wire buffer_12599 (.in(n12599), .out(n12599_0));
mux3 mux_7434 (.in({n9743_0, n9742_0, n1546}), .out(n12600), .config_in(config_chain[26743:26742]), .config_rst(config_rst)); 
buffer_wire buffer_12600 (.in(n12600), .out(n12600_0));
mux15 mux_7435 (.in({n12635_1, n10031_1, n10007_2, n9998_0, n9983_0, n9970_0, n9955_0, n9944_0, n9929_0, n9924_0, n1554, n1546, n1538, n570, n562}), .out(n12601), .config_in(config_chain[26749:26744]), .config_rst(config_rst)); 
buffer_wire buffer_12601 (.in(n12601), .out(n12601_0));
mux3 mux_7436 (.in({n9745_0, n9744_0, n1546}), .out(n12602), .config_in(config_chain[26751:26750]), .config_rst(config_rst)); 
buffer_wire buffer_12602 (.in(n12602), .out(n12602_0));
mux15 mux_7437 (.in({n12655_1, n10287_1, n10263_2, n10252_0, n10237_0, n10226_0, n10211_0, n10200_0, n10185_0, n10182_0, n1652, n1644, n1636, n668, n660}), .out(n12603), .config_in(config_chain[26757:26752]), .config_rst(config_rst)); 
buffer_wire buffer_12603 (.in(n12603), .out(n12603_0));
mux3 mux_7438 (.in({n9747_2, n9746_0/**/, n1550}), .out(n12604), .config_in(config_chain[26759:26758]), .config_rst(config_rst)); 
buffer_wire buffer_12604 (.in(n12604), .out(n12604_0));
mux13 mux_7439 (.in({n12757_0, n11597_2, n11570_0, n11567_0/**/, n11542_0, n11537_0, n11512_0, n11507_0, n11484_0, n2138, n2130, n1162, n1154}), .out(n12605), .config_in(config_chain[26765:26760]), .config_rst(config_rst)); 
buffer_wire buffer_12605 (.in(n12605), .out(n12605_0));
mux3 mux_7440 (.in({n9749_2, n9748_0, n1550}), .out(n12606), .config_in(config_chain[26767:26766]), .config_rst(config_rst)); 
buffer_wire buffer_12606 (.in(n12606), .out(n12606_0));
mux13 mux_7441 (.in({n12779_0, n11861_2, n11834_0, n11829_2, n11804_0, n11801_0, n11776_0, n11771_0, n11750_0/**/, n2236, n2228, n1260, n1252}), .out(n12607), .config_in(config_chain[26773:26768]), .config_rst(config_rst)); 
buffer_wire buffer_12607 (.in(n12607), .out(n12607_0));
mux3 mux_7442 (.in({n9751_2, n9750_0, n1550}), .out(n12608), .config_in(config_chain[26775:26774]), .config_rst(config_rst)); 
buffer_wire buffer_12608 (.in(n12608), .out(n12608_0));
mux3 mux_7443 (.in({n12123_2, n12094_0, n2334}), .out(n12609), .config_in(config_chain[26777:26776]), .config_rst(config_rst)); 
buffer_wire buffer_12609 (.in(n12609), .out(n12609_0));
mux3 mux_7444 (.in({n9753_2, n9752_0, n1550}), .out(n12610), .config_in(config_chain[26779:26778]), .config_rst(config_rst)); 
buffer_wire buffer_12610 (.in(n12610), .out(n12610_0));
mux3 mux_7445 (.in({n12097_0, n12096_0, n2334}), .out(n12611), .config_in(config_chain[26781:26780]), .config_rst(config_rst)); 
buffer_wire buffer_12611 (.in(n12611), .out(n12611_0));
mux3 mux_7446 (.in({n9755_2, n9754_0, n1550}), .out(n12612), .config_in(config_chain[26783:26782]), .config_rst(config_rst)); 
buffer_wire buffer_12612 (.in(n12612), .out(n12612_0));
mux3 mux_7447 (.in({n12099_0, n12098_0, n2334}), .out(n12613), .config_in(config_chain[26785:26784]), .config_rst(config_rst)); 
buffer_wire buffer_12613 (.in(n12613), .out(n12613_0));
mux3 mux_7448 (.in({n9757_2, n9756_0, n1554}), .out(n12614), .config_in(config_chain[26787:26786]), .config_rst(config_rst)); 
buffer_wire buffer_12614 (.in(n12614), .out(n12614_0));
mux3 mux_7449 (.in({n12101_0, n12100_0, n2338}), .out(n12615), .config_in(config_chain[26789:26788]), .config_rst(config_rst)); 
buffer_wire buffer_12615 (.in(n12615), .out(n12615_0));
mux16 mux_7450 (.in({n12528_0, n10015_1/**/, n10008_0, n10001_1, n9984_0, n9975_0, n9958_0, n9947_0, n9930_0, n9924_0, n9921_0, n1648, n1640, n672, n664, n656}), .out(n12616), .config_in(config_chain[26795:26790]), .config_rst(config_rst)); 
buffer_wire buffer_12616 (.in(n12616), .out(n12616_0));
mux16 mux_7451 (.in({n12697_1, n11065_1, n11045_1, n11036_0, n11021_0, n11010_0, n10995_0/**/, n10982_0, n10968_0, n10967_0, n10956_0, n1942, n1934, n966, n958, n950}), .out(n12617), .config_in(config_chain[26801:26796]), .config_rst(config_rst)); 
buffer_wire buffer_12617 (.in(n12617), .out(n12617_0));
mux16 mux_7452 (.in({n12536_0, n10017_1/**/, n10010_0, n10003_2, n9996_0, n9986_0, n9977_0, n9960_0, n9951_0, n9934_0, n9923_0, n1648, n1640, n672, n664, n656}), .out(n12618), .config_in(config_chain[26807:26802]), .config_rst(config_rst)); 
buffer_wire buffer_12618 (.in(n12618), .out(n12618_0));
mux16 mux_7453 (.in({n12699_1, n11063_1, n11047_2, n11038_0, n11023_0/**/, n11012_0, n10997_0, n10986_0, n10976_0, n10971_0, n10958_0, n1942, n1934, n966, n958, n950}), .out(n12619), .config_in(config_chain[26813:26808]), .config_rst(config_rst)); 
buffer_wire buffer_12619 (.in(n12619), .out(n12619_0));
mux15 mux_7454 (.in({n12544_0, n10019_1/**/, n10005_2, n9990_0, n9988_0, n9979_0, n9962_0, n9953_0, n9936_0, n9927_0, n1648, n1640, n672, n664, n656}), .out(n12620), .config_in(config_chain[26819:26814]), .config_rst(config_rst)); 
buffer_wire buffer_12620 (.in(n12620), .out(n12620_0));
mux15 mux_7455 (.in({n12701_1, n11061_1, n11040_0, n11027_0, n11014_0, n10999_0/**/, n10988_0, n10984_0, n10973_0, n10962_0, n1942, n1934, n966, n958, n950}), .out(n12621), .config_in(config_chain[26825:26820]), .config_rst(config_rst)); 
buffer_wire buffer_12621 (.in(n12621), .out(n12621_0));
mux15 mux_7456 (.in({n12552_0, n10021_1/**/, n10007_2, n9992_0, n9983_0, n9980_0, n9966_0, n9955_0, n9938_0, n9929_0, n1648, n1640, n672, n664, n656}), .out(n12622), .config_in(config_chain[26831:26826]), .config_rst(config_rst)); 
buffer_wire buffer_12622 (.in(n12622), .out(n12622_0));
mux15 mux_7457 (.in({n12703_1, n11059_1, n11042_0, n11029_0, n11018_0/**/, n11003_0, n10992_0, n10990_0, n10975_0, n10964_0, n1942, n1934, n966, n958, n950}), .out(n12623), .config_in(config_chain[26837:26832]), .config_rst(config_rst)); 
buffer_wire buffer_12623 (.in(n12623), .out(n12623_0));
mux15 mux_7458 (.in({n12560_0, n10023_1, n10009_2, n9994_0, n9985_0, n9972_0, n9968_0, n9959_0, n9942_0, n9931_0/**/, n1648, n1640, n672, n664, n656}), .out(n12624), .config_in(config_chain[26843:26838]), .config_rst(config_rst)); 
buffer_wire buffer_12624 (.in(n12624), .out(n12624_0));
mux15 mux_7459 (.in({n12705_1, n11057_1, n11044_0, n11031_0, n11020_0/**/, n11005_0, n11000_0, n10994_0, n10979_0, n10966_0, n1942, n1934, n966, n958, n950}), .out(n12625), .config_in(config_chain[26849:26844]), .config_rst(config_rst)); 
buffer_wire buffer_12625 (.in(n12625), .out(n12625_0));
mux15 mux_7460 (.in({n12568_0, n10025_1/**/, n10011_2, n9998_0, n9987_0, n9970_0, n9964_0, n9961_0, n9944_0, n9935_0, n1652, n1644, n1636, n668, n660}), .out(n12626), .config_in(config_chain[26855:26850]), .config_rst(config_rst)); 
buffer_wire buffer_12626 (.in(n12626), .out(n12626_0));
mux15 mux_7461 (.in({n12707_1, n11055_1, n11046_0, n11035_0, n11022_0, n11008_0, n11007_0, n10996_0, n10981_0, n10970_0, n1946, n1938, n1930, n962, n954/**/}), .out(n12627), .config_in(config_chain[26861:26856]), .config_rst(config_rst)); 
buffer_wire buffer_12627 (.in(n12627), .out(n12627_0));
mux15 mux_7462 (.in({n12576_0, n10027_1, n10000_0, n9991_0, n9974_0, n9963_0/**/, n9956_0, n9946_0, n9937_0, n9920_0, n1652, n1644, n1636, n668, n660}), .out(n12628), .config_in(config_chain[26867:26862]), .config_rst(config_rst)); 
buffer_wire buffer_12628 (.in(n12628), .out(n12628_0));
mux15 mux_7463 (.in({n12709_1, n11053_1, n11037_0, n11026_0, n11016_0, n11011_0, n10998_0, n10983_0, n10972_0, n10957_0/**/, n1946, n1938, n1930, n962, n954}), .out(n12629), .config_in(config_chain[26873:26868]), .config_rst(config_rst)); 
buffer_wire buffer_12629 (.in(n12629), .out(n12629_0));
mux15 mux_7464 (.in({n12584_0, n10029_1/**/, n10002_0, n9993_0, n9976_0, n9967_0, n9950_0, n9948_0, n9939_0, n9922_0, n1652, n1644, n1636, n668, n660}), .out(n12630), .config_in(config_chain[26879:26874]), .config_rst(config_rst)); 
buffer_wire buffer_12630 (.in(n12630), .out(n12630_0));
mux15 mux_7465 (.in({n12711_1, n11051_1, n11039_0, n11028_0, n11024_0, n11013_0, n11002_0, n10987_0, n10974_0, n10959_0, n1946/**/, n1938, n1930, n962, n954}), .out(n12631), .config_in(config_chain[26885:26880]), .config_rst(config_rst)); 
buffer_wire buffer_12631 (.in(n12631), .out(n12631_0));
mux15 mux_7466 (.in({n12592_0, n10031_1, n10004_0, n9995_0, n9978_0, n9969_0, n9952_0, n9943_0, n9940_0, n9926_0, n1652/**/, n1644, n1636, n668, n660}), .out(n12632), .config_in(config_chain[26891:26886]), .config_rst(config_rst)); 
buffer_wire buffer_12632 (.in(n12632), .out(n12632_0));
mux15 mux_7467 (.in({n12713_1, n11049_1, n11041_1, n11032_0, n11030_0, n11015_0, n11004_0, n10989_0, n10978_0, n10963_0, n1946, n1938, n1930, n962, n954/**/}), .out(n12633), .config_in(config_chain[26897:26892]), .config_rst(config_rst)); 
buffer_wire buffer_12633 (.in(n12633), .out(n12633_0));
mux15 mux_7468 (.in({n12600_0, n10013_1/**/, n10006_0, n9999_0, n9982_0, n9971_0, n9954_0, n9945_0, n9932_0, n9928_0, n1652, n1644, n1636, n668, n660}), .out(n12634), .config_in(config_chain[26903:26898]), .config_rst(config_rst)); 
buffer_wire buffer_12634 (.in(n12634), .out(n12634_0));
mux15 mux_7469 (.in({n12715_1, n11067_1, n11043_1, n11034_0, n11019_0, n11006_0, n10991_0, n10980_0/**/, n10965_0, n10960_0, n1946, n1938, n1930, n962, n954}), .out(n12635), .config_in(config_chain[26909:26904]), .config_rst(config_rst)); 
buffer_wire buffer_12635 (.in(n12635), .out(n12635_0));
mux16 mux_7470 (.in({n12530_0/**/, n10271_1, n10264_0, n10257_1, n10240_0, n10229_0, n10212_0, n10203_0, n10186_0, n10182_0, n10177_0, n1746, n1738, n770, n762, n754}), .out(n12636), .config_in(config_chain[26915:26910]), .config_rst(config_rst)); 
buffer_wire buffer_12636 (.in(n12636), .out(n12636_0));
mux16 mux_7471 (.in({n12717_0, n11329_1, n11309_1, n11300_0, n11285_0, n11272_0, n11257_0, n11246_0, n11234_0, n11231_0, n11220_0, n2040, n2032, n1064, n1056, n1048}), .out(n12637), .config_in(config_chain[26921:26916]), .config_rst(config_rst)); 
buffer_wire buffer_12637 (.in(n12637), .out(n12637_0));
mux16 mux_7472 (.in({n12538_0, n10273_1/**/, n10266_0, n10259_1, n10254_0, n10242_0, n10233_0, n10216_0, n10205_0, n10188_0, n10179_0, n1746, n1738, n770, n762, n754}), .out(n12638), .config_in(config_chain[26927:26922]), .config_rst(config_rst)); 
buffer_wire buffer_12638 (.in(n12638), .out(n12638_0));
mux16 mux_7473 (.in({n12719_0, n11327_1, n11311_1, n11302_0, n11287_0, n11276_0, n11261_0, n11248_0, n11242_0, n11233_0, n11222_0, n2040, n2032, n1064, n1056, n1048/**/}), .out(n12639), .config_in(config_chain[26933:26928]), .config_rst(config_rst)); 
buffer_wire buffer_12639 (.in(n12639), .out(n12639_0));
mux15 mux_7474 (.in({n12546_0/**/, n10275_1, n10261_2, n10246_0, n10244_0, n10235_0, n10218_0, n10209_0, n10192_0, n10181_0, n1746, n1738, n770, n762, n754}), .out(n12640), .config_in(config_chain[26939:26934]), .config_rst(config_rst)); 
buffer_wire buffer_12640 (.in(n12640), .out(n12640_0));
mux15 mux_7475 (.in({n12721_0, n11325_1, n11304_0, n11289_0, n11278_0, n11263_0, n11252_0, n11250_0/**/, n11237_0, n11224_0, n2040, n2032, n1064, n1056, n1048}), .out(n12641), .config_in(config_chain[26945:26940]), .config_rst(config_rst)); 
buffer_wire buffer_12641 (.in(n12641), .out(n12641_0));
mux15 mux_7476 (.in({n12554_0, n10277_1, n10263_2, n10248_0, n10238_0, n10237_0/**/, n10220_0, n10211_0, n10194_0, n10185_0, n1746, n1738, n770, n762, n754}), .out(n12642), .config_in(config_chain[26951:26946]), .config_rst(config_rst)); 
buffer_wire buffer_12642 (.in(n12642), .out(n12642_0));
mux15 mux_7477 (.in({n12723_0, n11323_1, n11306_0, n11293_0, n11280_0, n11265_0, n11258_0, n11254_0, n11239_0, n11228_0, n2040/**/, n2032, n1064, n1056, n1048}), .out(n12643), .config_in(config_chain[26957:26952]), .config_rst(config_rst)); 
buffer_wire buffer_12643 (.in(n12643), .out(n12643_0));
mux15 mux_7478 (.in({n12562_0, n10279_1, n10265_2, n10250_0, n10241_0, n10230_0, n10224_0/**/, n10213_0, n10196_0, n10187_0, n1746, n1738, n770, n762, n754}), .out(n12644), .config_in(config_chain[26963:26958]), .config_rst(config_rst)); 
buffer_wire buffer_12644 (.in(n12644), .out(n12644_0));
mux15 mux_7479 (.in({n12725_0, n11321_1, n11308_0, n11295_0, n11284_0/**/, n11269_0, n11266_0, n11256_0, n11241_0, n11230_0, n2040, n2032, n1064, n1056, n1048}), .out(n12645), .config_in(config_chain[26969:26964]), .config_rst(config_rst)); 
buffer_wire buffer_12645 (.in(n12645), .out(n12645_0));
mux15 mux_7480 (.in({n12570_0, n10281_1, n10267_2, n10252_0, n10243_0, n10226_0, n10222_0, n10217_0/**/, n10200_0, n10189_0, n1750, n1742, n1734, n766, n758}), .out(n12646), .config_in(config_chain[26975:26970]), .config_rst(config_rst)); 
buffer_wire buffer_12646 (.in(n12646), .out(n12646_0));
mux15 mux_7481 (.in({n12727_0, n11319_1, n11310_0, n11297_0, n11286_0/**/, n11274_0, n11271_0, n11260_0, n11245_0, n11232_0, n2044, n2036, n2028, n1060, n1052}), .out(n12647), .config_in(config_chain[26981:26976]), .config_rst(config_rst)); 
buffer_wire buffer_12647 (.in(n12647), .out(n12647_0));
mux15 mux_7482 (.in({n12578_0, n10283_1/**/, n10256_0, n10245_0, n10228_0, n10219_0, n10214_0, n10202_0, n10193_0, n10176_0, n1750, n1742, n1734, n766, n758}), .out(n12648), .config_in(config_chain[26987:26982]), .config_rst(config_rst)); 
buffer_wire buffer_12648 (.in(n12648), .out(n12648_0));
mux15 mux_7483 (.in({n12729_0, n11317_1, n11301_0, n11288_0, n11282_0, n11273_0, n11262_0, n11247_0, n11236_0/**/, n11221_0, n2044, n2036, n2028, n1060, n1052}), .out(n12649), .config_in(config_chain[26993:26988]), .config_rst(config_rst)); 
buffer_wire buffer_12649 (.in(n12649), .out(n12649_0));
mux15 mux_7484 (.in({n12586_0, n10285_1, n10258_0, n10249_0, n10232_0, n10221_0/**/, n10206_0, n10204_0, n10195_0, n10178_0, n1750, n1742, n1734, n766, n758}), .out(n12650), .config_in(config_chain[26999:26994]), .config_rst(config_rst)); 
buffer_wire buffer_12650 (.in(n12650), .out(n12650_0));
mux15 mux_7485 (.in({n12731_0, n11315_1, n11303_0, n11292_0/**/, n11290_0, n11277_0, n11264_0, n11249_0, n11238_0, n11223_0, n2044, n2036, n2028, n1060, n1052}), .out(n12651), .config_in(config_chain[27005:27000]), .config_rst(config_rst)); 
buffer_wire buffer_12651 (.in(n12651), .out(n12651_0));
mux15 mux_7486 (.in({n12594_0, n10287_1, n10260_0, n10251_0, n10234_0, n10225_0, n10208_0, n10198_0/**/, n10197_0, n10180_0, n1750, n1742, n1734, n766, n758}), .out(n12652), .config_in(config_chain[27011:27006]), .config_rst(config_rst)); 
buffer_wire buffer_12652 (.in(n12652), .out(n12652_0));
mux15 mux_7487 (.in({n12733_0, n11313_1, n11305_0, n11298_0, n11294_0, n11279_0, n11268_0, n11253_0, n11240_0, n11225_0/**/, n2044, n2036, n2028, n1060, n1052}), .out(n12653), .config_in(config_chain[27017:27012]), .config_rst(config_rst)); 
buffer_wire buffer_12653 (.in(n12653), .out(n12653_0));
mux15 mux_7488 (.in({n12602_0, n10269_1, n10262_0, n10253_0, n10236_0, n10227_0, n10210_0/**/, n10201_0, n10190_0, n10184_0, n1750, n1742, n1734, n766, n758}), .out(n12654), .config_in(config_chain[27023:27018]), .config_rst(config_rst)); 
buffer_wire buffer_12654 (.in(n12654), .out(n12654_0));
mux15 mux_7489 (.in({n12735_0, n11331_1, n11307_1, n11296_0, n11281_0, n11270_0, n11255_0, n11244_0, n11229_0, n11226_0, n2044/**/, n2036, n2028, n1060, n1052}), .out(n12655), .config_in(config_chain[27029:27024]), .config_rst(config_rst)); 
buffer_wire buffer_12655 (.in(n12655), .out(n12655_0));
mux16 mux_7490 (.in({n12524_0, n10529_1, n10522_0, n10515_1, n10500_0, n10489_0, n10472_0, n10463_0, n10446_0, n10437_0, n10434_0/**/, n1844, n1836, n868, n860, n852}), .out(n12656), .config_in(config_chain[27035:27030]), .config_rst(config_rst)); 
buffer_wire buffer_12656 (.in(n12656), .out(n12656_0));
mux15 mux_7491 (.in({n12737_0, n11595_1, n11572_0, n11569_0, n11544_0, n11539_0, n11514_0, n11511_0, n11492_0, n11486_0, n2138, n2130, n1162/**/, n1154, n1146}), .out(n12657), .config_in(config_chain[27041:27036]), .config_rst(config_rst)); 
buffer_wire buffer_12657 (.in(n12657), .out(n12657_0));
mux16 mux_7492 (.in({n12532_0, n10531_1, n10524_0, n10517_1, n10506_0, n10502_0, n10493_0, n10476_0, n10465_0/**/, n10448_0, n10439_0, n1844, n1836, n868, n860, n852}), .out(n12658), .config_in(config_chain[27047:27042]), .config_rst(config_rst)); 
buffer_wire buffer_12658 (.in(n12658), .out(n12658_0));
mux15 mux_7493 (.in({n12739_0, n11593_1/**/, n11574_0, n11571_0, n11546_0, n11543_0, n11518_0, n11513_0, n11500_0, n11488_0, n2142, n2130, n1162, n1154, n1146}), .out(n12659), .config_in(config_chain[27053:27048]), .config_rst(config_rst)); 
buffer_wire buffer_12659 (.in(n12659), .out(n12659_0));
mux15 mux_7494 (.in({n12540_0, n10533_1, n10519_1, n10504_0, n10498_0, n10495_0, n10478_0, n10469_0, n10452_0/**/, n10441_0, n1844, n1836, n868, n860, n852}), .out(n12660), .config_in(config_chain[27059:27054]), .config_rst(config_rst)); 
buffer_wire buffer_12660 (.in(n12660), .out(n12660_0));
mux15 mux_7495 (.in({n12741_0/**/, n11591_1, n11573_1, n11550_0, n11545_0, n11520_0, n11515_0, n11508_0, n11490_0, n11487_0, n2142, n2134, n1162, n1154, n1146}), .out(n12661), .config_in(config_chain[27065:27060]), .config_rst(config_rst)); 
buffer_wire buffer_12661 (.in(n12661), .out(n12661_0));
mux15 mux_7496 (.in({n12548_0, n10535_1, n10521_2, n10508_0/**/, n10497_0, n10490_0, n10480_0, n10471_0, n10454_0, n10445_0, n1844, n1836, n868, n860, n852}), .out(n12662), .config_in(config_chain[27071:27066]), .config_rst(config_rst)); 
buffer_wire buffer_12662 (.in(n12662), .out(n12662_0));
mux15 mux_7497 (.in({n12743_0, n11589_1, n11575_1/**/, n11552_0, n11547_0, n11522_0, n11519_0, n11516_0, n11494_0, n11489_0, n2142, n2134, n2126, n1154, n1146}), .out(n12663), .config_in(config_chain[27077:27072]), .config_rst(config_rst)); 
buffer_wire buffer_12663 (.in(n12663), .out(n12663_0));
mux15 mux_7498 (.in({n12556_0, n10537_1, n10523_2, n10510_0, n10501_0, n10484_0/**/, n10482_0, n10473_0, n10456_0, n10447_0, n1844, n1836, n868, n860, n852}), .out(n12664), .config_in(config_chain[27083:27078]), .config_rst(config_rst)); 
buffer_wire buffer_12664 (.in(n12664), .out(n12664_0));
mux14 mux_7499 (.in({n12745_0/**/, n11587_1, n11554_0, n11551_0, n11526_0, n11524_0, n11521_0, n11496_0, n11491_0, n2142, n2134, n2126, n1158, n1146}), .out(n12665), .config_in(config_chain[27089:27084]), .config_rst(config_rst)); 
buffer_wire buffer_12665 (.in(n12665), .out(n12665_0));
mux15 mux_7500 (.in({n12564_0, n10539_1, n10525_2, n10512_0, n10503_0, n10486_0, n10477_0, n10474_0, n10460_0, n10449_0, n1848, n1840/**/, n1832, n864, n856}), .out(n12666), .config_in(config_chain[27095:27090]), .config_rst(config_rst)); 
buffer_wire buffer_12666 (.in(n12666), .out(n12666_0));
mux14 mux_7501 (.in({n12747_0, n11585_1/**/, n11558_0, n11553_0, n11532_0, n11528_0, n11523_0, n11498_0, n11495_0, n2142, n2134, n2126, n1158, n1150}), .out(n12667), .config_in(config_chain[27101:27096]), .config_rst(config_rst)); 
buffer_wire buffer_12667 (.in(n12667), .out(n12667_0));
mux15 mux_7502 (.in({n12572_0, n10541_1, n10514_0, n10505_0, n10488_0, n10479_0, n10466_0, n10462_0, n10453_0, n10436_0, n1848, n1840, n1832, n864, n856/**/}), .out(n12668), .config_in(config_chain[27107:27102]), .config_rst(config_rst)); 
buffer_wire buffer_12668 (.in(n12668), .out(n12668_0));
mux13 mux_7503 (.in({n12749_0, n11583_1, n11560_0, n11555_0, n11540_0/**/, n11530_0, n11527_0, n11502_0, n11497_0, n2134, n2126, n1158, n1150}), .out(n12669), .config_in(config_chain[27113:27108]), .config_rst(config_rst)); 
buffer_wire buffer_12669 (.in(n12669), .out(n12669_0));
mux15 mux_7504 (.in({n12580_0, n10543_1, n10516_0, n10509_0/**/, n10492_0, n10481_0, n10464_0, n10458_0, n10455_0, n10438_0, n1848, n1840, n1832, n864, n856}), .out(n12670), .config_in(config_chain[27119:27114]), .config_rst(config_rst)); 
buffer_wire buffer_12670 (.in(n12670), .out(n12670_0));
mux13 mux_7505 (.in({n12751_0, n11581_1/**/, n11562_0, n11559_0, n11548_0, n11534_0, n11529_0, n11504_0, n11499_0, n2138, n2126, n1158, n1150}), .out(n12671), .config_in(config_chain[27125:27120]), .config_rst(config_rst)); 
buffer_wire buffer_12671 (.in(n12671), .out(n12671_0));
mux15 mux_7506 (.in({n12588_0, n10545_1, n10518_0, n10511_0, n10494_0, n10485_0, n10468_0, n10457_0, n10450_0, n10440_0, n1848, n1840, n1832, n864, n856/**/}), .out(n12672), .config_in(config_chain[27131:27126]), .config_rst(config_rst)); 
buffer_wire buffer_12672 (.in(n12672), .out(n12672_0));
mux13 mux_7507 (.in({n12753_0, n11579_1, n11566_0, n11561_0, n11556_0/**/, n11536_0, n11531_0, n11506_0, n11503_0, n2138, n2130, n1158, n1150}), .out(n12673), .config_in(config_chain[27137:27132]), .config_rst(config_rst)); 
buffer_wire buffer_12673 (.in(n12673), .out(n12673_0));
mux15 mux_7508 (.in({n12596_0, n10527_1, n10520_0, n10513_0, n10496_0, n10487_0, n10470_0, n10461_0, n10444_0, n10442_0, n1848, n1840, n1832/**/, n864, n856}), .out(n12674), .config_in(config_chain[27143:27138]), .config_rst(config_rst)); 
buffer_wire buffer_12674 (.in(n12674), .out(n12674_0));
mux13 mux_7509 (.in({n12755_0, n11577_1, n11568_0, n11564_0, n11563_0, n11538_0, n11535_0, n11510_0, n11505_0, n2138, n2130, n1162, n1150}), .out(n12675), .config_in(config_chain[27149:27144]), .config_rst(config_rst)); 
buffer_wire buffer_12675 (.in(n12675), .out(n12675_0));
mux16 mux_7510 (.in({n12526_1/**/, n10789_1, n10782_0, n10775_0, n10758_0, n10749_0, n10732_0, n10723_0, n10706_0, n10696_0, n10695_0, n1942, n1934, n966, n958, n950}), .out(n12676), .config_in(config_chain[27155:27150]), .config_rst(config_rst)); 
buffer_wire buffer_12676 (.in(n12676), .out(n12676_0));
mux15 mux_7511 (.in({n12759_0, n11859_1/**/, n11836_0, n11833_0, n11808_0, n11803_0, n11778_0, n11773_0, n11758_0, n11748_0, n2236, n2228, n1260, n1252, n1244}), .out(n12677), .config_in(config_chain[27161:27156]), .config_rst(config_rst)); 
buffer_wire buffer_12677 (.in(n12677), .out(n12677_0));
mux16 mux_7512 (.in({n12534_1, n10791_1, n10784_0, n10777_1, n10768_0/**/, n10762_0, n10751_0, n10734_0, n10725_0, n10708_0, n10699_0, n1942, n1934, n966, n958, n950}), .out(n12678), .config_in(config_chain[27167:27162]), .config_rst(config_rst)); 
buffer_wire buffer_12678 (.in(n12678), .out(n12678_0));
mux15 mux_7513 (.in({n12761_0, n11857_1, n11838_0, n11835_0, n11810_0, n11805_0, n11780_0, n11777_0, n11766_0/**/, n11752_0, n2240, n2228, n1260, n1252, n1244}), .out(n12679), .config_in(config_chain[27173:27168]), .config_rst(config_rst)); 
buffer_wire buffer_12679 (.in(n12679), .out(n12679_0));
mux15 mux_7514 (.in({n12542_1/**/, n10793_1, n10779_1, n10764_0, n10760_0, n10755_0, n10738_0, n10727_0, n10710_0, n10701_0, n1942, n1934, n966, n958, n950}), .out(n12680), .config_in(config_chain[27179:27174]), .config_rst(config_rst)); 
buffer_wire buffer_12680 (.in(n12680), .out(n12680_0));
mux15 mux_7515 (.in({n12763_0, n11855_1, n11837_0, n11812_0, n11809_0/**/, n11784_0, n11779_0, n11774_0, n11754_0, n11749_0, n2240, n2232, n1260, n1252, n1244}), .out(n12681), .config_in(config_chain[27185:27180]), .config_rst(config_rst)); 
buffer_wire buffer_12681 (.in(n12681), .out(n12681_0));
mux15 mux_7516 (.in({n12550_1, n10795_1, n10781_1, n10766_0, n10757_0, n10752_0, n10740_0, n10731_0, n10714_0, n10703_0, n1942, n1934, n966/**/, n958, n950}), .out(n12682), .config_in(config_chain[27191:27186]), .config_rst(config_rst)); 
buffer_wire buffer_12682 (.in(n12682), .out(n12682_0));
mux15 mux_7517 (.in({n12765_0, n11853_1, n11839_1, n11816_0, n11811_0, n11786_0, n11782_0, n11781_0, n11756_0, n11753_0, n2240/**/, n2232, n2224, n1252, n1244}), .out(n12683), .config_in(config_chain[27197:27192]), .config_rst(config_rst)); 
buffer_wire buffer_12683 (.in(n12683), .out(n12683_0));
mux15 mux_7518 (.in({n12558_1/**/, n10797_1, n10783_2, n10770_0, n10759_0, n10744_0, n10742_0, n10733_0, n10716_0, n10707_0, n1942, n1934, n966, n958, n950}), .out(n12684), .config_in(config_chain[27203:27198]), .config_rst(config_rst)); 
buffer_wire buffer_12684 (.in(n12684), .out(n12684_0));
mux14 mux_7519 (.in({n12767_0, n11851_1, n11818_0, n11813_0, n11790_0, n11788_0, n11785_0, n11760_0, n11755_0, n2240, n2232/**/, n2224, n1256, n1244}), .out(n12685), .config_in(config_chain[27209:27204]), .config_rst(config_rst)); 
buffer_wire buffer_12685 (.in(n12685), .out(n12685_0));
mux15 mux_7520 (.in({n12566_1, n10799_1, n10785_2, n10772_0, n10763_0, n10746_0, n10736_0, n10735_0, n10718_0, n10709_0, n1946, n1938, n1930, n962/**/, n954}), .out(n12686), .config_in(config_chain[27215:27210]), .config_rst(config_rst)); 
buffer_wire buffer_12686 (.in(n12686), .out(n12686_0));
mux14 mux_7521 (.in({n12769_0, n11849_1, n11820_0, n11817_0, n11798_0, n11792_0, n11787_0/**/, n11762_0, n11757_0, n2240, n2232, n2224, n1256, n1248}), .out(n12687), .config_in(config_chain[27221:27216]), .config_rst(config_rst)); 
buffer_wire buffer_12687 (.in(n12687), .out(n12687_0));
mux15 mux_7522 (.in({n12574_1, n10801_1, n10774_0, n10765_0, n10748_0, n10739_0, n10728_0, n10722_0, n10711_0, n10694_0, n1946, n1938, n1930, n962, n954/**/}), .out(n12688), .config_in(config_chain[27227:27222]), .config_rst(config_rst)); 
buffer_wire buffer_12688 (.in(n12688), .out(n12688_0));
mux13 mux_7523 (.in({n12771_0, n11847_1, n11824_0, n11819_0/**/, n11806_0, n11794_0, n11789_0, n11764_0, n11761_0, n2232, n2224, n1256, n1248}), .out(n12689), .config_in(config_chain[27233:27228]), .config_rst(config_rst)); 
buffer_wire buffer_12689 (.in(n12689), .out(n12689_0));
mux15 mux_7524 (.in({n12582_1, n10803_1, n10776_0, n10767_0, n10750_0, n10741_0, n10724_0, n10720_0, n10715_0, n10698_0, n1946, n1938, n1930/**/, n962, n954}), .out(n12690), .config_in(config_chain[27239:27234]), .config_rst(config_rst)); 
buffer_wire buffer_12690 (.in(n12690), .out(n12690_0));
mux13 mux_7525 (.in({n12773_0, n11845_1, n11826_0, n11821_0, n11814_0, n11796_0, n11793_0/**/, n11768_0, n11763_0, n2236, n2224, n1256, n1248}), .out(n12691), .config_in(config_chain[27245:27240]), .config_rst(config_rst)); 
buffer_wire buffer_12691 (.in(n12691), .out(n12691_0));
mux15 mux_7526 (.in({n12590_1/**/, n10805_1, n10778_0, n10771_0, n10754_0, n10743_0, n10726_0, n10717_0, n10712_0, n10700_0, n1946, n1938, n1930, n962, n954}), .out(n12692), .config_in(config_chain[27251:27246]), .config_rst(config_rst)); 
buffer_wire buffer_12692 (.in(n12692), .out(n12692_0));
mux13 mux_7527 (.in({n12775_0, n11843_1, n11828_0, n11825_0, n11822_0, n11800_0, n11795_0, n11770_0, n11765_0, n2236, n2228, n1256, n1248}), .out(n12693), .config_in(config_chain[27257:27252]), .config_rst(config_rst)); 
buffer_wire buffer_12693 (.in(n12693), .out(n12693_0));
mux15 mux_7528 (.in({n12598_1/**/, n10787_1, n10780_0, n10773_0, n10756_0, n10747_0, n10730_0, n10719_0, n10704_0, n10702_0, n1946, n1938, n1930, n962, n954}), .out(n12694), .config_in(config_chain[27263:27258]), .config_rst(config_rst)); 
buffer_wire buffer_12694 (.in(n12694), .out(n12694_0));
mux13 mux_7529 (.in({n12777_0, n11841_1/**/, n11832_0, n11830_0, n11827_0, n11802_0, n11797_0, n11772_0, n11769_0, n2236, n2228, n1260, n1248}), .out(n12695), .config_in(config_chain[27269:27264]), .config_rst(config_rst)); 
buffer_wire buffer_12695 (.in(n12695), .out(n12695_0));
mux16 mux_7530 (.in({n12616_1, n11051_1, n11044_0, n11037_0, n11020_0, n11011_0, n10994_0, n10983_0, n10966_0, n10960_0/**/, n10957_0, n2040, n2032, n1064, n1056, n1048}), .out(n12696), .config_in(config_chain[27275:27270]), .config_rst(config_rst)); 
buffer_wire buffer_12696 (.in(n12696), .out(n12696_0));
mux4 mux_7531 (.in({n12103_1/**/, n12014_0, n2338, n1342}), .out(n12697), .config_in(config_chain[27277:27276]), .config_rst(config_rst)); 
buffer_wire buffer_12697 (.in(n12697), .out(n12697_0));
mux16 mux_7532 (.in({n12618_1, n11053_1, n11046_0, n11039_0, n11032_0, n11022_0, n11013_0, n10996_0, n10987_0/**/, n10970_0, n10959_0, n2040, n2032, n1064, n1056, n1048}), .out(n12698), .config_in(config_chain[27283:27278]), .config_rst(config_rst)); 
buffer_wire buffer_12698 (.in(n12698), .out(n12698_0));
mux3 mux_7533 (.in({n12105_1, n12022_0, n1346}), .out(n12699), .config_in(config_chain[27285:27284]), .config_rst(config_rst)); 
buffer_wire buffer_12699 (.in(n12699), .out(n12699_0));
mux15 mux_7534 (.in({n12620_1, n11055_1, n11041_1, n11026_0, n11024_0, n11015_0, n10998_0, n10989_0, n10972_0, n10963_0, n2040, n2032, n1064, n1056, n1048/**/}), .out(n12700), .config_in(config_chain[27291:27286]), .config_rst(config_rst)); 
buffer_wire buffer_12700 (.in(n12700), .out(n12700_0));
mux3 mux_7535 (.in({n12107_1, n12030_0, n1350}), .out(n12701), .config_in(config_chain[27293:27292]), .config_rst(config_rst)); 
buffer_wire buffer_12701 (.in(n12701), .out(n12701_0));
mux15 mux_7536 (.in({n12622_1, n11057_1, n11043_1, n11028_0, n11019_0, n11016_0, n11002_0/**/, n10991_0, n10974_0, n10965_0, n2040, n2032, n1064, n1056, n1048}), .out(n12702), .config_in(config_chain[27299:27294]), .config_rst(config_rst)); 
buffer_wire buffer_12702 (.in(n12702), .out(n12702_0));
mux3 mux_7537 (.in({n12109_1/**/, n12038_0, n1350}), .out(n12703), .config_in(config_chain[27301:27300]), .config_rst(config_rst)); 
buffer_wire buffer_12703 (.in(n12703), .out(n12703_0));
mux15 mux_7538 (.in({n12624_1, n11059_1, n11045_1, n11030_0, n11021_0, n11008_0, n11004_0, n10995_0, n10978_0, n10967_0, n2040, n2032, n1064, n1056, n1048/**/}), .out(n12704), .config_in(config_chain[27307:27302]), .config_rst(config_rst)); 
buffer_wire buffer_12704 (.in(n12704), .out(n12704_0));
mux3 mux_7539 (.in({n12111_1, n12046_0, n1354}), .out(n12705), .config_in(config_chain[27309:27308]), .config_rst(config_rst)); 
buffer_wire buffer_12705 (.in(n12705), .out(n12705_0));
mux15 mux_7540 (.in({n12626_1, n11061_1, n11047_2, n11034_0, n11023_0, n11006_0, n11000_0, n10997_0, n10980_0/**/, n10971_0, n2044, n2036, n2028, n1060, n1052}), .out(n12706), .config_in(config_chain[27315:27310]), .config_rst(config_rst)); 
buffer_wire buffer_12706 (.in(n12706), .out(n12706_0));
mux3 mux_7541 (.in({n12113_1, n12054_0, n1358}), .out(n12707), .config_in(config_chain[27317:27316]), .config_rst(config_rst)); 
buffer_wire buffer_12707 (.in(n12707), .out(n12707_0));
mux15 mux_7542 (.in({n12628_1, n11063_1, n11036_0, n11027_0, n11010_0, n10999_0, n10992_0, n10982_0, n10973_0, n10956_0/**/, n2044, n2036, n2028, n1060, n1052}), .out(n12708), .config_in(config_chain[27323:27318]), .config_rst(config_rst)); 
buffer_wire buffer_12708 (.in(n12708), .out(n12708_0));
mux3 mux_7543 (.in({n12115_1, n12062_0, n2322}), .out(n12709), .config_in(config_chain[27325:27324]), .config_rst(config_rst)); 
buffer_wire buffer_12709 (.in(n12709), .out(n12709_0));
mux15 mux_7544 (.in({n12630_1/**/, n11065_1, n11038_0, n11029_0, n11012_0, n11003_0, n10986_0, n10984_0, n10975_0, n10958_0, n2044, n2036, n2028, n1060, n1052}), .out(n12710), .config_in(config_chain[27331:27326]), .config_rst(config_rst)); 
buffer_wire buffer_12710 (.in(n12710), .out(n12710_0));
mux3 mux_7545 (.in({n12117_1, n12070_0, n2326}), .out(n12711), .config_in(config_chain[27333:27332]), .config_rst(config_rst)); 
buffer_wire buffer_12711 (.in(n12711), .out(n12711_0));
mux15 mux_7546 (.in({n12632_1, n11067_1, n11040_0, n11031_0, n11014_0, n11005_0, n10988_0, n10979_0/**/, n10976_0, n10962_0, n2044, n2036, n2028, n1060, n1052}), .out(n12712), .config_in(config_chain[27339:27334]), .config_rst(config_rst)); 
buffer_wire buffer_12712 (.in(n12712), .out(n12712_0));
mux3 mux_7547 (.in({n12119_1/**/, n12078_0, n2326}), .out(n12713), .config_in(config_chain[27341:27340]), .config_rst(config_rst)); 
buffer_wire buffer_12713 (.in(n12713), .out(n12713_0));
mux15 mux_7548 (.in({n12634_1, n11049_1, n11042_0, n11035_0, n11018_0, n11007_0, n10990_0, n10981_0/**/, n10968_0, n10964_0, n2044, n2036, n2028, n1060, n1052}), .out(n12714), .config_in(config_chain[27347:27342]), .config_rst(config_rst)); 
buffer_wire buffer_12714 (.in(n12714), .out(n12714_0));
mux3 mux_7549 (.in({n12121_1/**/, n12086_0, n2330}), .out(n12715), .config_in(config_chain[27349:27348]), .config_rst(config_rst)); 
buffer_wire buffer_12715 (.in(n12715), .out(n12715_0));
mux16 mux_7550 (.in({n12636_1, n11315_1, n11308_0, n11301_0, n11284_0, n11273_0, n11256_0, n11247_0, n11230_0, n11226_0, n11221_0/**/, n2138, n2130, n1162, n1154, n1146}), .out(n12716), .config_in(config_chain[27355:27350]), .config_rst(config_rst)); 
buffer_wire buffer_12716 (.in(n12716), .out(n12716_0));
mux4 mux_7551 (.in({n12017_0, n12016_0, n2338, n1342}), .out(n12717), .config_in(config_chain[27357:27356]), .config_rst(config_rst)); 
buffer_wire buffer_12717 (.in(n12717), .out(n12717_0));
mux16 mux_7552 (.in({n12638_1, n11317_1, n11310_0, n11303_0, n11298_0, n11286_0, n11277_0, n11260_0, n11249_0, n11232_0, n11223_0, n2138, n2130, n1162, n1154, n1146}), .out(n12718), .config_in(config_chain[27363:27358]), .config_rst(config_rst)); 
buffer_wire buffer_12718 (.in(n12718), .out(n12718_0));
mux3 mux_7553 (.in({n12025_0, n12024_0, n1346}), .out(n12719), .config_in(config_chain[27365:27364]), .config_rst(config_rst)); 
buffer_wire buffer_12719 (.in(n12719), .out(n12719_0));
mux15 mux_7554 (.in({n12640_1/**/, n11319_1, n11305_0, n11290_0, n11288_0, n11279_0, n11262_0, n11253_0, n11236_0, n11225_0, n2138, n2130, n1162, n1154, n1146}), .out(n12720), .config_in(config_chain[27371:27366]), .config_rst(config_rst)); 
buffer_wire buffer_12720 (.in(n12720), .out(n12720_0));
mux3 mux_7555 (.in({n12033_0/**/, n12032_0, n1350}), .out(n12721), .config_in(config_chain[27373:27372]), .config_rst(config_rst)); 
buffer_wire buffer_12721 (.in(n12721), .out(n12721_0));
mux15 mux_7556 (.in({n12642_1, n11321_1/**/, n11307_1, n11292_0, n11282_0, n11281_0, n11264_0, n11255_0, n11238_0, n11229_0, n2138, n2130, n1162, n1154, n1146}), .out(n12722), .config_in(config_chain[27379:27374]), .config_rst(config_rst)); 
buffer_wire buffer_12722 (.in(n12722), .out(n12722_0));
mux3 mux_7557 (.in({n12041_0, n12040_0, n1354}), .out(n12723), .config_in(config_chain[27381:27380]), .config_rst(config_rst)); 
buffer_wire buffer_12723 (.in(n12723), .out(n12723_0));
mux15 mux_7558 (.in({n12644_1, n11323_1, n11309_1, n11294_0, n11285_0, n11274_0, n11268_0, n11257_0, n11240_0, n11231_0/**/, n2138, n2130, n1162, n1154, n1146}), .out(n12724), .config_in(config_chain[27387:27382]), .config_rst(config_rst)); 
buffer_wire buffer_12724 (.in(n12724), .out(n12724_0));
mux3 mux_7559 (.in({n12049_0, n12048_0, n1354}), .out(n12725), .config_in(config_chain[27389:27388]), .config_rst(config_rst)); 
buffer_wire buffer_12725 (.in(n12725), .out(n12725_0));
mux15 mux_7560 (.in({n12646_1/**/, n11325_1, n11311_1, n11296_0, n11287_0, n11270_0, n11266_0, n11261_0, n11244_0, n11233_0, n2142, n2134, n2126, n1158, n1150}), .out(n12726), .config_in(config_chain[27395:27390]), .config_rst(config_rst)); 
buffer_wire buffer_12726 (.in(n12726), .out(n12726_0));
mux3 mux_7561 (.in({n12057_0, n12056_0, n1358}), .out(n12727), .config_in(config_chain[27397:27396]), .config_rst(config_rst)); 
buffer_wire buffer_12727 (.in(n12727), .out(n12727_0));
mux15 mux_7562 (.in({n12648_1, n11327_1, n11300_0, n11289_0, n11272_0, n11263_0, n11258_0, n11246_0, n11237_0, n11220_0, n2142, n2134, n2126, n1158, n1150}), .out(n12728), .config_in(config_chain[27403:27398]), .config_rst(config_rst)); 
buffer_wire buffer_12728 (.in(n12728), .out(n12728_0));
mux3 mux_7563 (.in({n12065_0, n12064_0, n2322}), .out(n12729), .config_in(config_chain[27405:27404]), .config_rst(config_rst)); 
buffer_wire buffer_12729 (.in(n12729), .out(n12729_0));
mux15 mux_7564 (.in({n12650_1, n11329_1, n11302_0, n11293_0, n11276_0, n11265_0, n11250_0, n11248_0, n11239_0, n11222_0, n2142/**/, n2134, n2126, n1158, n1150}), .out(n12730), .config_in(config_chain[27411:27406]), .config_rst(config_rst)); 
buffer_wire buffer_12730 (.in(n12730), .out(n12730_0));
mux3 mux_7565 (.in({n12073_0, n12072_0, n2326/**/}), .out(n12731), .config_in(config_chain[27413:27412]), .config_rst(config_rst)); 
buffer_wire buffer_12731 (.in(n12731), .out(n12731_0));
mux15 mux_7566 (.in({n12652_1, n11331_1, n11304_0, n11295_0, n11278_0, n11269_0, n11252_0, n11242_0, n11241_0, n11224_0/**/, n2142, n2134, n2126, n1158, n1150}), .out(n12732), .config_in(config_chain[27419:27414]), .config_rst(config_rst)); 
buffer_wire buffer_12732 (.in(n12732), .out(n12732_0));
mux3 mux_7567 (.in({n12081_0, n12080_0, n2330}), .out(n12733), .config_in(config_chain[27421:27420]), .config_rst(config_rst)); 
buffer_wire buffer_12733 (.in(n12733), .out(n12733_0));
mux15 mux_7568 (.in({n12654_1, n11313_1, n11306_0, n11297_0, n11280_0, n11271_0, n11254_0, n11245_0, n11234_0/**/, n11228_0, n2142, n2134, n2126, n1158, n1150}), .out(n12734), .config_in(config_chain[27427:27422]), .config_rst(config_rst)); 
buffer_wire buffer_12734 (.in(n12734), .out(n12734_0));
mux3 mux_7569 (.in({n12089_0, n12088_0, n2330}), .out(n12735), .config_in(config_chain[27429:27428]), .config_rst(config_rst)); 
buffer_wire buffer_12735 (.in(n12735), .out(n12735_0));
mux15 mux_7570 (.in({n12656_1, n11579_1, n11573_1, n11568_0, n11545_0, n11538_0, n11515_0, n11510_0, n11487_0, n11484_0, n2236, n2228, n1260/**/, n1252, n1244}), .out(n12736), .config_in(config_chain[27435:27430]), .config_rst(config_rst)); 
buffer_wire buffer_12736 (.in(n12736), .out(n12736_0));
mux4 mux_7571 (.in({n12011_0, n12010_0, n2338/**/, n1342}), .out(n12737), .config_in(config_chain[27437:27436]), .config_rst(config_rst)); 
buffer_wire buffer_12737 (.in(n12737), .out(n12737_0));
mux15 mux_7572 (.in({n12658_1, n11581_1, n11575_1, n11570_0, n11564_0, n11547_0, n11542_0, n11519_0, n11512_0, n11489_0, n2240, n2228, n1260, n1252, n1244/**/}), .out(n12738), .config_in(config_chain[27443:27438]), .config_rst(config_rst)); 
buffer_wire buffer_12738 (.in(n12738), .out(n12738_0));
mux3 mux_7573 (.in({n12019_0/**/, n12018_0, n1342}), .out(n12739), .config_in(config_chain[27445:27444]), .config_rst(config_rst)); 
buffer_wire buffer_12739 (.in(n12739), .out(n12739_0));
mux15 mux_7574 (.in({n12660_1, n11583_1, n11572_0, n11556_0, n11551_0, n11544_0, n11521_0, n11514_0, n11491_0, n11486_0, n2240, n2232/**/, n1260, n1252, n1244}), .out(n12740), .config_in(config_chain[27451:27446]), .config_rst(config_rst)); 
buffer_wire buffer_12740 (.in(n12740), .out(n12740_0));
mux3 mux_7575 (.in({n12027_0/**/, n12026_0, n1346}), .out(n12741), .config_in(config_chain[27453:27452]), .config_rst(config_rst)); 
buffer_wire buffer_12741 (.in(n12741), .out(n12741_0));
mux15 mux_7576 (.in({n12662_1, n11585_1, n11574_0, n11553_0, n11548_0/**/, n11546_0, n11523_0, n11518_0, n11495_0, n11488_0, n2240, n2232, n2224, n1252, n1244}), .out(n12742), .config_in(config_chain[27459:27454]), .config_rst(config_rst)); 
buffer_wire buffer_12742 (.in(n12742), .out(n12742_0));
mux3 mux_7577 (.in({n12035_0/**/, n12034_0, n1350}), .out(n12743), .config_in(config_chain[27461:27460]), .config_rst(config_rst)); 
buffer_wire buffer_12743 (.in(n12743), .out(n12743_0));
mux14 mux_7578 (.in({n12664_1, n11587_1, n11555_0, n11550_0, n11540_0, n11527_0, n11520_0, n11497_0, n11490_0, n2240, n2232, n2224, n1256, n1244}), .out(n12744), .config_in(config_chain[27467:27462]), .config_rst(config_rst)); 
buffer_wire buffer_12744 (.in(n12744), .out(n12744_0));
mux3 mux_7579 (.in({n12043_0/**/, n12042_0, n1354}), .out(n12745), .config_in(config_chain[27469:27468]), .config_rst(config_rst)); 
buffer_wire buffer_12745 (.in(n12745), .out(n12745_0));
mux14 mux_7580 (.in({n12666_1, n11589_1, n11559_0/**/, n11552_0, n11532_0, n11529_0, n11522_0, n11499_0, n11494_0, n2240, n2232, n2224, n1256, n1248}), .out(n12746), .config_in(config_chain[27475:27470]), .config_rst(config_rst)); 
buffer_wire buffer_12746 (.in(n12746), .out(n12746_0));
mux3 mux_7581 (.in({n12051_0, n12050_0, n1358}), .out(n12747), .config_in(config_chain[27477:27476]), .config_rst(config_rst)); 
buffer_wire buffer_12747 (.in(n12747), .out(n12747_0));
mux13 mux_7582 (.in({n12668_1, n11591_1, n11561_0, n11554_0, n11531_0, n11526_0, n11524_0, n11503_0, n11496_0, n2232, n2224, n1256, n1248}), .out(n12748), .config_in(config_chain[27483:27478]), .config_rst(config_rst)); 
buffer_wire buffer_12748 (.in(n12748), .out(n12748_0));
mux3 mux_7583 (.in({n12059_0/**/, n12058_0, n1358}), .out(n12749), .config_in(config_chain[27485:27484]), .config_rst(config_rst)); 
buffer_wire buffer_12749 (.in(n12749), .out(n12749_0));
mux13 mux_7584 (.in({n12670_1, n11593_1, n11563_0, n11558_0, n11535_0, n11528_0, n11516_0, n11505_0, n11498_0, n2236, n2224, n1256/**/, n1248}), .out(n12750), .config_in(config_chain[27491:27486]), .config_rst(config_rst)); 
buffer_wire buffer_12750 (.in(n12750), .out(n12750_0));
mux3 mux_7585 (.in({n12067_0, n12066_0, n2322}), .out(n12751), .config_in(config_chain[27493:27492]), .config_rst(config_rst)); 
buffer_wire buffer_12751 (.in(n12751), .out(n12751_0));
mux13 mux_7586 (.in({n12672_1, n11595_1, n11567_0, n11560_0, n11537_0, n11530_0, n11508_0/**/, n11507_0, n11502_0, n2236, n2228, n1256, n1248}), .out(n12752), .config_in(config_chain[27499:27494]), .config_rst(config_rst)); 
buffer_wire buffer_12752 (.in(n12752), .out(n12752_0));
mux3 mux_7587 (.in({n12075_0, n12074_0, n2326}), .out(n12753), .config_in(config_chain[27501:27500]), .config_rst(config_rst)); 
buffer_wire buffer_12753 (.in(n12753), .out(n12753_0));
mux13 mux_7588 (.in({n12674_1, n11597_2, n11569_0, n11562_0, n11539_0, n11534_0, n11511_0, n11504_0, n11500_0, n2236, n2228, n1260, n1248}), .out(n12754), .config_in(config_chain[27507:27502]), .config_rst(config_rst)); 
buffer_wire buffer_12754 (.in(n12754), .out(n12754_0));
mux3 mux_7589 (.in({n12083_0, n12082_0, n2330}), .out(n12755), .config_in(config_chain[27509:27508]), .config_rst(config_rst)); 
buffer_wire buffer_12755 (.in(n12755), .out(n12755_0));
mux13 mux_7590 (.in({n12604_2, n11577_1, n11571_0, n11566_0, n11543_0, n11536_0, n11513_0, n11506_0, n11492_0, n2236, n2228, n1260, n1252}), .out(n12756), .config_in(config_chain[27515:27510]), .config_rst(config_rst)); 
buffer_wire buffer_12756 (.in(n12756), .out(n12756_0));
mux3 mux_7591 (.in({n12091_2, n12090_0, n2334}), .out(n12757), .config_in(config_chain[27517:27516]), .config_rst(config_rst)); 
buffer_wire buffer_12757 (.in(n12757), .out(n12757_0));
mux15 mux_7592 (.in({n12676_1/**/, n11843_1, n11837_0, n11832_0, n11809_0, n11802_0, n11779_0, n11772_0, n11750_0, n11749_0, n2334, n2326, n1358, n1350, n1342}), .out(n12758), .config_in(config_chain[27523:27518]), .config_rst(config_rst)); 
buffer_wire buffer_12758 (.in(n12758), .out(n12758_0));
mux4 mux_7593 (.in({n12013_0, n12012_0, n2338, n1342}), .out(n12759), .config_in(config_chain[27525:27524]), .config_rst(config_rst)); 
buffer_wire buffer_12759 (.in(n12759), .out(n12759_0));
mux15 mux_7594 (.in({n12678_1, n11845_1, n11839_1, n11834_0, n11830_0, n11811_0, n11804_0, n11781_0, n11776_0, n11753_0, n2338, n2326, n1358, n1350, n1342}), .out(n12760), .config_in(config_chain[27531:27526]), .config_rst(config_rst)); 
buffer_wire buffer_12760 (.in(n12760), .out(n12760_0));
mux3 mux_7595 (.in({n12021_0, n12020_0, n1346}), .out(n12761), .config_in(config_chain[27533:27532]), .config_rst(config_rst)); 
buffer_wire buffer_12761 (.in(n12761), .out(n12761_0));
mux15 mux_7596 (.in({n12680_1, n11847_1, n11836_0, n11822_0, n11813_0, n11808_0, n11785_0, n11778_0, n11755_0/**/, n11748_0, n2338, n2330, n1358, n1350, n1342}), .out(n12762), .config_in(config_chain[27539:27534]), .config_rst(config_rst)); 
buffer_wire buffer_12762 (.in(n12762), .out(n12762_0));
mux3 mux_7597 (.in({n12029_0, n12028_0, n1346}), .out(n12763), .config_in(config_chain[27541:27540]), .config_rst(config_rst)); 
buffer_wire buffer_12763 (.in(n12763), .out(n12763_0));
mux15 mux_7598 (.in({n12682_1, n11849_1/**/, n11838_0, n11817_0, n11814_0, n11810_0, n11787_0, n11780_0, n11757_0, n11752_0, n2338, n2330, n2322, n1350, n1342}), .out(n12764), .config_in(config_chain[27547:27542]), .config_rst(config_rst)); 
buffer_wire buffer_12764 (.in(n12764), .out(n12764_0));
mux3 mux_7599 (.in({n12037_0, n12036_0, n1350}), .out(n12765), .config_in(config_chain[27549:27548]), .config_rst(config_rst)); 
buffer_wire buffer_12765 (.in(n12765), .out(n12765_0));
mux14 mux_7600 (.in({n12684_1, n11851_1, n11819_0, n11812_0, n11806_0, n11789_0, n11784_0, n11761_0, n11754_0, n2338, n2330, n2322, n1354, n1342}), .out(n12766), .config_in(config_chain[27555:27550]), .config_rst(config_rst)); 
buffer_wire buffer_12766 (.in(n12766), .out(n12766_0));
mux3 mux_7601 (.in({n12045_0, n12044_0, n1354}), .out(n12767), .config_in(config_chain[27557:27556]), .config_rst(config_rst)); 
buffer_wire buffer_12767 (.in(n12767), .out(n12767_0));
mux14 mux_7602 (.in({n12686_1, n11853_1, n11821_0, n11816_0, n11798_0, n11793_0, n11786_0, n11763_0, n11756_0, n2338, n2330, n2322, n1354, n1346}), .out(n12768), .config_in(config_chain[27563:27558]), .config_rst(config_rst)); 
buffer_wire buffer_12768 (.in(n12768), .out(n12768_0));
mux3 mux_7603 (.in({n12053_0, n12052_0, n1358}), .out(n12769), .config_in(config_chain[27565:27564]), .config_rst(config_rst)); 
buffer_wire buffer_12769 (.in(n12769), .out(n12769_0));
mux13 mux_7604 (.in({n12688_1, n11855_1, n11825_0, n11818_0, n11795_0, n11790_0, n11788_0, n11765_0, n11760_0, n2330, n2322, n1354, n1346}), .out(n12770), .config_in(config_chain[27571:27566]), .config_rst(config_rst)); 
buffer_wire buffer_12770 (.in(n12770), .out(n12770_0));
mux3 mux_7605 (.in({n12061_0, n12060_0, n2322}), .out(n12771), .config_in(config_chain[27573:27572]), .config_rst(config_rst)); 
buffer_wire buffer_12771 (.in(n12771), .out(n12771_0));
mux13 mux_7606 (.in({n12690_1/**/, n11857_1, n11827_0, n11820_0, n11797_0, n11792_0, n11782_0, n11769_0, n11762_0, n2334, n2322, n1354, n1346}), .out(n12772), .config_in(config_chain[27579:27574]), .config_rst(config_rst)); 
buffer_wire buffer_12772 (.in(n12772), .out(n12772_0));
mux3 mux_7607 (.in({n12069_0, n12068_0/**/, n2322}), .out(n12773), .config_in(config_chain[27581:27580]), .config_rst(config_rst)); 
buffer_wire buffer_12773 (.in(n12773), .out(n12773_0));
mux13 mux_7608 (.in({n12692_1, n11859_1, n11829_2, n11824_0, n11801_0, n11794_0, n11774_0, n11771_0, n11764_0/**/, n2334, n2326, n1354, n1346}), .out(n12774), .config_in(config_chain[27587:27582]), .config_rst(config_rst)); 
buffer_wire buffer_12774 (.in(n12774), .out(n12774_0));
mux3 mux_7609 (.in({n12077_0, n12076_0, n2326}), .out(n12775), .config_in(config_chain[27589:27588]), .config_rst(config_rst)); 
buffer_wire buffer_12775 (.in(n12775), .out(n12775_0));
mux13 mux_7610 (.in({n12694_1, n11861_2, n11833_0/**/, n11826_0, n11803_0, n11796_0, n11773_0, n11768_0, n11766_0, n2334, n2326, n1358, n1346}), .out(n12776), .config_in(config_chain[27595:27590]), .config_rst(config_rst)); 
buffer_wire buffer_12776 (.in(n12776), .out(n12776_0));
mux3 mux_7611 (.in({n12085_0, n12084_0/**/, n2330}), .out(n12777), .config_in(config_chain[27597:27596]), .config_rst(config_rst)); 
buffer_wire buffer_12777 (.in(n12777), .out(n12777_0));
mux13 mux_7612 (.in({n12606_2, n11841_1, n11835_0, n11828_0, n11805_0, n11800_0, n11777_0, n11770_0, n11758_0, n2334/**/, n2326, n1358, n1350}), .out(n12778), .config_in(config_chain[27603:27598]), .config_rst(config_rst)); 
buffer_wire buffer_12778 (.in(n12778), .out(n12778_0));
mux3 mux_7613 (.in({n12093_2, n12092_0, n2334}), .out(n12779), .config_in(config_chain[27605:27604]), .config_rst(config_rst)); 
buffer_wire buffer_12779 (.in(n12779), .out(n12779_0));
mux4 mux_7614 (.in({n9667_0/**/, n9666_0, n2532, n1536}), .out(n12780), .config_in(config_chain[27607:27606]), .config_rst(config_rst)); 
buffer_wire buffer_12780 (.in(n12780), .out(n12780_0));
mux16 mux_7615 (.in({n12893_1, n10305_1, n10280_0, n10277_0, n10265_2, n10256_0, n10243_0, n10204_0, n10189_0, n10184_0, n10178_0, n2626/**/, n2618, n1650, n1642, n1634}), .out(n12781), .config_in(config_chain[27613:27608]), .config_rst(config_rst)); 
buffer_wire buffer_12781 (.in(n12781), .out(n12781_0));
mux4 mux_7616 (.in({n9759_0/**/, n9758_0, n2532, n1536}), .out(n12782), .config_in(config_chain[27615:27614]), .config_rst(config_rst)); 
buffer_wire buffer_12782 (.in(n12782), .out(n12782_0));
mux16 mux_7617 (.in({n12913_1, n10563_1, n10543_0, n10526_0, n10523_2, n10514_0, n10488_0, n10473_0, n10462_0, n10447_0, n10444_0, n2724, n2716, n1748, n1740, n1732/**/}), .out(n12783), .config_in(config_chain[27621:27616]), .config_rst(config_rst)); 
buffer_wire buffer_12783 (.in(n12783), .out(n12783_0));
mux4 mux_7618 (.in({n9779_1, n9670_0, n2532, n1536}), .out(n12784), .config_in(config_chain[27623:27622]), .config_rst(config_rst)); 
buffer_wire buffer_12784 (.in(n12784), .out(n12784_0));
mux16 mux_7619 (.in({n12933_1, n10823_1, n10792_0, n10789_0, n10783_1, n10774_0, n10759_0, n10748_0, n10733_0, n10706_0, n10694_0, n2822, n2814, n1846, n1838, n1830}), .out(n12785), .config_in(config_chain[27629:27624]), .config_rst(config_rst)); 
buffer_wire buffer_12785 (.in(n12785), .out(n12785_0));
mux4 mux_7620 (.in({n9673_0, n9672_0, n2532/**/, n1536}), .out(n12786), .config_in(config_chain[27631:27630]), .config_rst(config_rst)); 
buffer_wire buffer_12786 (.in(n12786), .out(n12786_0));
mux16 mux_7621 (.in({n12873_1, n10049_1, n10024_0, n10021_0, n10009_2, n10000_0, n9985_0, n9946_0, n9934_0, n9931_0, n9920_0, n2528, n2520, n1552, n1544, n1536}), .out(n12787), .config_in(config_chain[27637:27632]), .config_rst(config_rst)); 
buffer_wire buffer_12787 (.in(n12787), .out(n12787_0));
mux3 mux_7622 (.in({n9675_0/**/, n9674_0, n1536}), .out(n12788), .config_in(config_chain[27639:27638]), .config_rst(config_rst)); 
buffer_wire buffer_12788 (.in(n12788), .out(n12788_0));
mux16 mux_7623 (.in({n12895_1, n10303_1, n10274_0, n10271_0, n10267_2, n10258_0, n10245_0, n10234_0, n10219_0, n10192_0, n10180_0, n2626, n2618, n1650, n1642, n1634}), .out(n12789), .config_in(config_chain[27645:27640]), .config_rst(config_rst)); 
buffer_wire buffer_12789 (.in(n12789), .out(n12789_0));
mux3 mux_7624 (.in({n9761_0/**/, n9760_0, n1540}), .out(n12790), .config_in(config_chain[27647:27646]), .config_rst(config_rst)); 
buffer_wire buffer_12790 (.in(n12790), .out(n12790_0));
mux16 mux_7625 (.in({n12915_1, n10561_1, n10540_0, n10537_0, n10525_2, n10516_0, n10503_0, n10464_0, n10452_0, n10449_0, n10438_0, n2724, n2716, n1748, n1740, n1732/**/}), .out(n12791), .config_in(config_chain[27653:27648]), .config_rst(config_rst)); 
buffer_wire buffer_12791 (.in(n12791), .out(n12791_0));
mux3 mux_7626 (.in({n9781_1, n9678_0/**/, n1540}), .out(n12792), .config_in(config_chain[27655:27654]), .config_rst(config_rst)); 
buffer_wire buffer_12792 (.in(n12792), .out(n12792_0));
mux16 mux_7627 (.in({n12935_1, n10821_1/**/, n10803_0, n10786_0, n10785_2, n10776_0, n10750_0, n10735_0, n10724_0, n10714_0, n10709_0, n2822, n2814, n1846, n1838, n1830}), .out(n12793), .config_in(config_chain[27661:27656]), .config_rst(config_rst)); 
buffer_wire buffer_12793 (.in(n12793), .out(n12793_0));
mux3 mux_7628 (.in({n9681_0, n9680_0, n1540}), .out(n12794), .config_in(config_chain[27663:27662]), .config_rst(config_rst)); 
buffer_wire buffer_12794 (.in(n12794), .out(n12794_0));
mux16 mux_7629 (.in({n12875_1, n10047_1, n10018_0, n10015_0, n10011_2, n10002_0, n9987_0, n9976_0, n9961_0, n9942_0, n9922_0, n2528, n2520, n1552, n1544, n1536}), .out(n12795), .config_in(config_chain[27669:27664]), .config_rst(config_rst)); 
buffer_wire buffer_12795 (.in(n12795), .out(n12795_0));
mux3 mux_7630 (.in({n9683_0, n9682_0, n1540}), .out(n12796), .config_in(config_chain[27671:27670]), .config_rst(config_rst)); 
buffer_wire buffer_12796 (.in(n12796), .out(n12796_0));
mux15 mux_7631 (.in({n12897_1, n10301_1, n10285_0, n10268_0, n10260_0, n10236_0, n10221_0, n10210_0, n10200_0, n10195_0, n2626, n2618, n1650/**/, n1642, n1634}), .out(n12797), .config_in(config_chain[27677:27672]), .config_rst(config_rst)); 
buffer_wire buffer_12797 (.in(n12797), .out(n12797_0));
mux3 mux_7632 (.in({n9763_0, n9762_0, n1540}), .out(n12798), .config_in(config_chain[27679:27678]), .config_rst(config_rst)); 
buffer_wire buffer_12798 (.in(n12798), .out(n12798_0));
mux15 mux_7633 (.in({n12917_1, n10559_1, n10534_0, n10531_0, n10518_0, n10505_0, n10494_0, n10479_0, n10460_0, n10440_0, n2724, n2716, n1748/**/, n1740, n1732}), .out(n12799), .config_in(config_chain[27685:27680]), .config_rst(config_rst)); 
buffer_wire buffer_12799 (.in(n12799), .out(n12799_0));
mux3 mux_7634 (.in({n9783_1, n9686_0/**/, n1544}), .out(n12800), .config_in(config_chain[27687:27686]), .config_rst(config_rst)); 
buffer_wire buffer_12800 (.in(n12800), .out(n12800_0));
mux15 mux_7635 (.in({n12937_1, n10819_1, n10800_0, n10797_0, n10778_0, n10765_0, n10726_0, n10722_0, n10711_0, n10700_0, n2822, n2814, n1846, n1838, n1830/**/}), .out(n12801), .config_in(config_chain[27693:27688]), .config_rst(config_rst)); 
buffer_wire buffer_12801 (.in(n12801), .out(n12801_0));
mux3 mux_7636 (.in({n9689_0, n9688_0, n1544}), .out(n12802), .config_in(config_chain[27695:27694]), .config_rst(config_rst)); 
buffer_wire buffer_12802 (.in(n12802), .out(n12802_0));
mux15 mux_7637 (.in({n12877_1, n10045_1, n10029_0, n10012_0, n10004_0, n9978_0, n9963_0, n9952_0, n9950_0, n9937_0, n2528, n2520/**/, n1552, n1544, n1536}), .out(n12803), .config_in(config_chain[27701:27696]), .config_rst(config_rst)); 
buffer_wire buffer_12803 (.in(n12803), .out(n12803_0));
mux3 mux_7638 (.in({n9691_0, n9690_0, n1544}), .out(n12804), .config_in(config_chain[27703:27702]), .config_rst(config_rst)); 
buffer_wire buffer_12804 (.in(n12804), .out(n12804_0));
mux15 mux_7639 (.in({n12899_1, n10299_1, n10282_0, n10279_0, n10262_0, n10251_0, n10212_0, n10208_0, n10197_0, n10186_0, n2626, n2618, n1650, n1642, n1634}), .out(n12805), .config_in(config_chain[27709:27704]), .config_rst(config_rst)); 
buffer_wire buffer_12805 (.in(n12805), .out(n12805_0));
mux3 mux_7640 (.in({n9765_0/**/, n9764_0, n1544}), .out(n12806), .config_in(config_chain[27711:27710]), .config_rst(config_rst)); 
buffer_wire buffer_12806 (.in(n12806), .out(n12806_0));
mux15 mux_7641 (.in({n12919_1/**/, n10557_1, n10545_0, n10528_0, n10520_0, n10496_0, n10481_0, n10470_0, n10468_0, n10455_0, n2724, n2716, n1748, n1740, n1732}), .out(n12807), .config_in(config_chain[27717:27712]), .config_rst(config_rst)); 
buffer_wire buffer_12807 (.in(n12807), .out(n12807_0));
mux3 mux_7642 (.in({n9785_1, n9694_0, n1544}), .out(n12808), .config_in(config_chain[27719:27718]), .config_rst(config_rst)); 
buffer_wire buffer_12808 (.in(n12808), .out(n12808_0));
mux15 mux_7643 (.in({n12939_1, n10817_1, n10794_0, n10791_0, n10780_0, n10767_0, n10756_0, n10741_0, n10730_0, n10702_0, n2822/**/, n2814, n1846, n1838, n1830}), .out(n12809), .config_in(config_chain[27725:27720]), .config_rst(config_rst)); 
buffer_wire buffer_12809 (.in(n12809), .out(n12809_0));
mux3 mux_7644 (.in({n9697_0, n9696_0, n1548}), .out(n12810), .config_in(config_chain[27727:27726]), .config_rst(config_rst)); 
buffer_wire buffer_12810 (.in(n12810), .out(n12810_0));
mux15 mux_7645 (.in({n12879_1, n10043_1, n10026_0, n10023_0, n10006_0, n9993_0, n9958_0, n9954_0, n9939_0, n9928_0, n2528, n2520, n1552, n1544, n1536}), .out(n12811), .config_in(config_chain[27733:27728]), .config_rst(config_rst)); 
buffer_wire buffer_12811 (.in(n12811), .out(n12811_0));
mux3 mux_7646 (.in({n9699_0, n9698_0, n1548}), .out(n12812), .config_in(config_chain[27735:27734]), .config_rst(config_rst)); 
buffer_wire buffer_12812 (.in(n12812), .out(n12812_0));
mux15 mux_7647 (.in({n12901_1/**/, n10297_1, n10276_0, n10273_0, n10264_0, n10253_0, n10242_0, n10227_0, n10216_0, n10188_0, n2626, n2618, n1650, n1642, n1634}), .out(n12813), .config_in(config_chain[27741:27736]), .config_rst(config_rst)); 
buffer_wire buffer_12813 (.in(n12813), .out(n12813_0));
mux3 mux_7648 (.in({n9767_0/**/, n9766_0, n1548}), .out(n12814), .config_in(config_chain[27743:27742]), .config_rst(config_rst)); 
buffer_wire buffer_12814 (.in(n12814), .out(n12814_0));
mux15 mux_7649 (.in({n12921_1, n10555_1, n10542_0, n10539_0, n10522_0, n10511_0, n10476_0, n10472_0, n10457_0, n10446_0, n2724, n2716, n1748, n1740, n1732}), .out(n12815), .config_in(config_chain[27749:27744]), .config_rst(config_rst)); 
buffer_wire buffer_12815 (.in(n12815), .out(n12815_0));
mux3 mux_7650 (.in({n9787_1, n9702_0, n1548}), .out(n12816), .config_in(config_chain[27751:27750]), .config_rst(config_rst)); 
buffer_wire buffer_12816 (.in(n12816), .out(n12816_0));
mux15 mux_7651 (.in({n12941_1, n10815_1, n10805_0, n10788_0, n10782_0, n10758_0, n10743_0, n10738_0, n10732_0, n10717_0, n2822/**/, n2814, n1846, n1838, n1830}), .out(n12817), .config_in(config_chain[27757:27752]), .config_rst(config_rst)); 
buffer_wire buffer_12817 (.in(n12817), .out(n12817_0));
mux3 mux_7652 (.in({n9705_0, n9704_0, n1548}), .out(n12818), .config_in(config_chain[27759:27758]), .config_rst(config_rst)); 
buffer_wire buffer_12818 (.in(n12818), .out(n12818_0));
mux15 mux_7653 (.in({n12881_1, n10041_1, n10020_0, n10017_0, n10008_0, n9995_0, n9984_0, n9969_0/**/, n9966_0, n9930_0, n2528, n2520, n1552, n1544, n1536}), .out(n12819), .config_in(config_chain[27765:27760]), .config_rst(config_rst)); 
buffer_wire buffer_12819 (.in(n12819), .out(n12819_0));
mux3 mux_7654 (.in({n9707_0, n9706_0, n1552}), .out(n12820), .config_in(config_chain[27767:27766]), .config_rst(config_rst)); 
buffer_wire buffer_12820 (.in(n12820), .out(n12820_0));
mux15 mux_7655 (.in({n12903_1, n10295_1, n10287_0, n10270_0, n10266_0, n10244_0, n10229_0, n10224_0, n10218_0, n10203_0, n2630, n2622, n2614, n1646, n1638/**/}), .out(n12821), .config_in(config_chain[27773:27768]), .config_rst(config_rst)); 
buffer_wire buffer_12821 (.in(n12821), .out(n12821_0));
mux3 mux_7656 (.in({n9769_0/**/, n9768_0, n1552}), .out(n12822), .config_in(config_chain[27775:27774]), .config_rst(config_rst)); 
buffer_wire buffer_12822 (.in(n12822), .out(n12822_0));
mux15 mux_7657 (.in({n12923_1, n10553_1, n10536_0, n10533_0, n10524_0, n10513_0, n10502_0, n10487_0, n10484_0, n10448_0, n2728, n2720, n2712, n1744, n1736}), .out(n12823), .config_in(config_chain[27781:27776]), .config_rst(config_rst)); 
buffer_wire buffer_12823 (.in(n12823), .out(n12823_0));
mux3 mux_7658 (.in({n9789_1, n9710_0/**/, n1552}), .out(n12824), .config_in(config_chain[27783:27782]), .config_rst(config_rst)); 
buffer_wire buffer_12824 (.in(n12824), .out(n12824_0));
mux15 mux_7659 (.in({n12943_1, n10813_1, n10802_0, n10799_0, n10784_0, n10773_0, n10746_0, n10734_0, n10719_0, n10708_0, n2826, n2818, n2810, n1842/**/, n1834}), .out(n12825), .config_in(config_chain[27789:27784]), .config_rst(config_rst)); 
buffer_wire buffer_12825 (.in(n12825), .out(n12825_0));
mux3 mux_7660 (.in({n9713_0, n9712_0, n1552}), .out(n12826), .config_in(config_chain[27791:27790]), .config_rst(config_rst)); 
buffer_wire buffer_12826 (.in(n12826), .out(n12826_0));
mux15 mux_7661 (.in({n12883_1, n10039_1, n10031_0, n10014_0, n10010_0, n9986_0/**/, n9974_0, n9971_0, n9960_0, n9945_0, n2532, n2524, n2516, n1548, n1540}), .out(n12827), .config_in(config_chain[27797:27792]), .config_rst(config_rst)); 
buffer_wire buffer_12827 (.in(n12827), .out(n12827_0));
mux3 mux_7662 (.in({n9715_0, n9714_0, n1552}), .out(n12828), .config_in(config_chain[27799:27798]), .config_rst(config_rst)); 
buffer_wire buffer_12828 (.in(n12828), .out(n12828_0));
mux15 mux_7663 (.in({n12905_1, n10293_1, n10284_0, n10281_0, n10257_1, n10232_0, n10220_0, n10205_0, n10194_0, n10179_0/**/, n2630, n2622, n2614, n1646, n1638}), .out(n12829), .config_in(config_chain[27805:27800]), .config_rst(config_rst)); 
buffer_wire buffer_12829 (.in(n12829), .out(n12829_0));
mux3 mux_7664 (.in({n9771_0, n9770_0, n2516}), .out(n12830), .config_in(config_chain[27807:27806]), .config_rst(config_rst)); 
buffer_wire buffer_12830 (.in(n12830), .out(n12830_0));
mux15 mux_7665 (.in({n12925_1/**/, n10551_1, n10530_0, n10527_0, n10515_0, n10504_0, n10492_0, n10489_0, n10478_0, n10463_0, n2728, n2720, n2712, n1744, n1736}), .out(n12831), .config_in(config_chain[27813:27808]), .config_rst(config_rst)); 
buffer_wire buffer_12831 (.in(n12831), .out(n12831_0));
mux3 mux_7666 (.in({n9791_1, n9718_0/**/, n2516}), .out(n12832), .config_in(config_chain[27815:27814]), .config_rst(config_rst)); 
buffer_wire buffer_12832 (.in(n12832), .out(n12832_0));
mux15 mux_7667 (.in({n12945_1, n10811_1/**/, n10796_0, n10793_0, n10775_0, n10764_0, n10754_0, n10749_0, n10710_0, n10695_0, n2826, n2818, n2810, n1842, n1834}), .out(n12833), .config_in(config_chain[27821:27816]), .config_rst(config_rst)); 
buffer_wire buffer_12833 (.in(n12833), .out(n12833_0));
mux3 mux_7668 (.in({n9721_0, n9720_0/**/, n2516}), .out(n12834), .config_in(config_chain[27823:27822]), .config_rst(config_rst)); 
buffer_wire buffer_12834 (.in(n12834), .out(n12834_0));
mux15 mux_7669 (.in({n12885_1, n10037_1, n10028_0, n10025_0, n10001_1, n9982_0, n9962_0, n9947_0, n9936_0, n9921_0, n2532, n2524, n2516, n1548, n1540}), .out(n12835), .config_in(config_chain[27829:27824]), .config_rst(config_rst)); 
buffer_wire buffer_12835 (.in(n12835), .out(n12835_0));
mux3 mux_7670 (.in({n9723_0, n9722_0, n2516}), .out(n12836), .config_in(config_chain[27831:27830]), .config_rst(config_rst)); 
buffer_wire buffer_12836 (.in(n12836), .out(n12836_0));
mux15 mux_7671 (.in({n12907_1, n10291_1, n10278_0, n10275_0, n10259_1, n10250_0/**/, n10240_0, n10235_0, n10196_0, n10181_0, n2630, n2622, n2614, n1646, n1638}), .out(n12837), .config_in(config_chain[27837:27832]), .config_rst(config_rst)); 
buffer_wire buffer_12837 (.in(n12837), .out(n12837_0));
mux3 mux_7672 (.in({n9773_0, n9772_0, n2516}), .out(n12838), .config_in(config_chain[27839:27838]), .config_rst(config_rst)); 
buffer_wire buffer_12838 (.in(n12838), .out(n12838_0));
mux15 mux_7673 (.in({n12927_1, n10549_1, n10544_0, n10541_0, n10517_1, n10500_0/**/, n10480_0, n10465_0, n10454_0, n10439_0, n2728, n2720, n2712, n1744, n1736}), .out(n12839), .config_in(config_chain[27845:27840]), .config_rst(config_rst)); 
buffer_wire buffer_12839 (.in(n12839), .out(n12839_0));
mux3 mux_7674 (.in({n9793_1, n9726_0, n2520}), .out(n12840), .config_in(config_chain[27847:27846]), .config_rst(config_rst)); 
buffer_wire buffer_12840 (.in(n12840), .out(n12840_0));
mux15 mux_7675 (.in({n12947_1, n10809_1, n10790_0, n10787_0, n10777_0, n10766_0, n10762_0, n10751_0, n10740_0, n10725_0, n2826/**/, n2818, n2810, n1842, n1834}), .out(n12841), .config_in(config_chain[27853:27848]), .config_rst(config_rst)); 
buffer_wire buffer_12841 (.in(n12841), .out(n12841_0));
mux3 mux_7676 (.in({n9729_0, n9728_0, n2520/**/}), .out(n12842), .config_in(config_chain[27855:27854]), .config_rst(config_rst)); 
buffer_wire buffer_12842 (.in(n12842), .out(n12842_0));
mux15 mux_7677 (.in({n12887_1, n10035_1, n10022_0, n10019_0, n10003_1, n9992_0, n9990_0, n9977_0, n9938_0, n9923_0, n2532, n2524, n2516, n1548, n1540}), .out(n12843), .config_in(config_chain[27861:27856]), .config_rst(config_rst)); 
buffer_wire buffer_12843 (.in(n12843), .out(n12843_0));
mux3 mux_7678 (.in({n9731_0, n9730_0, n2520}), .out(n12844), .config_in(config_chain[27863:27862]), .config_rst(config_rst)); 
buffer_wire buffer_12844 (.in(n12844), .out(n12844_0));
mux15 mux_7679 (.in({n12909_1, n10289_1, n10272_0, n10269_0/**/, n10261_1, n10252_0, n10248_0, n10237_0, n10226_0, n10211_0, n2630, n2622, n2614, n1646, n1638}), .out(n12845), .config_in(config_chain[27869:27864]), .config_rst(config_rst)); 
buffer_wire buffer_12845 (.in(n12845), .out(n12845_0));
mux3 mux_7680 (.in({n9775_0/**/, n9774_0, n2520}), .out(n12846), .config_in(config_chain[27871:27870]), .config_rst(config_rst)); 
buffer_wire buffer_12846 (.in(n12846), .out(n12846_0));
mux15 mux_7681 (.in({n12929_1, n10547_1, n10538_0, n10535_0, n10519_1, n10510_0, n10508_0, n10495_0, n10456_0, n10441_0, n2728, n2720, n2712, n1744, n1736}), .out(n12847), .config_in(config_chain[27877:27872]), .config_rst(config_rst)); 
buffer_wire buffer_12847 (.in(n12847), .out(n12847_0));
mux3 mux_7682 (.in({n9795_1, n9734_0, n2520}), .out(n12848), .config_in(config_chain[27879:27878]), .config_rst(config_rst)); 
buffer_wire buffer_12848 (.in(n12848), .out(n12848_0));
mux15 mux_7683 (.in({n12949_1/**/, n10807_1, n10804_0, n10801_0, n10779_1, n10770_0, n10742_0, n10727_0, n10716_0, n10701_0, n2826, n2818, n2810, n1842, n1834}), .out(n12849), .config_in(config_chain[27885:27880]), .config_rst(config_rst)); 
buffer_wire buffer_12849 (.in(n12849), .out(n12849_0));
mux3 mux_7684 (.in({n9737_0, n9736_0, n2524}), .out(n12850), .config_in(config_chain[27887:27886]), .config_rst(config_rst)); 
buffer_wire buffer_12850 (.in(n12850), .out(n12850_0));
mux15 mux_7685 (.in({n12889_1, n10033_1, n10016_0, n10013_0, n10005_2, n9998_0, n9994_0, n9979_0, n9968_0, n9953_0, n2532, n2524, n2516, n1548, n1540}), .out(n12851), .config_in(config_chain[27893:27888]), .config_rst(config_rst)); 
buffer_wire buffer_12851 (.in(n12851), .out(n12851_0));
mux3 mux_7686 (.in({n9739_0, n9738_0, n2524}), .out(n12852), .config_in(config_chain[27895:27894]), .config_rst(config_rst)); 
buffer_wire buffer_12852 (.in(n12852), .out(n12852_0));
mux15 mux_7687 (.in({n12911_1, n10307_1, n10286_0, n10283_0, n10263_2, n10228_0, n10213_0, n10202_0, n10187_0, n10176_0, n2630, n2622, n2614, n1646, n1638/**/}), .out(n12853), .config_in(config_chain[27901:27896]), .config_rst(config_rst)); 
buffer_wire buffer_12853 (.in(n12853), .out(n12853_0));
mux3 mux_7688 (.in({n9777_0/**/, n9776_0, n2524}), .out(n12854), .config_in(config_chain[27903:27902]), .config_rst(config_rst)); 
buffer_wire buffer_12854 (.in(n12854), .out(n12854_0));
mux15 mux_7689 (.in({n12931_1, n10565_1, n10532_0, n10529_0, n10521_1, n10512_0, n10497_0, n10486_0, n10471_0, n10436_0, n2728, n2720/**/, n2712, n1744, n1736}), .out(n12855), .config_in(config_chain[27909:27904]), .config_rst(config_rst)); 
buffer_wire buffer_12855 (.in(n12855), .out(n12855_0));
mux3 mux_7690 (.in({n9797_1, n9742_0/**/, n2524}), .out(n12856), .config_in(config_chain[27911:27910]), .config_rst(config_rst)); 
buffer_wire buffer_12856 (.in(n12856), .out(n12856_0));
mux15 mux_7691 (.in({n12951_1, n10825_1, n10798_0/**/, n10795_0, n10781_1, n10772_0, n10757_0, n10718_0, n10703_0, n10698_0, n2826, n2818, n2810, n1842, n1834}), .out(n12857), .config_in(config_chain[27917:27912]), .config_rst(config_rst)); 
buffer_wire buffer_12857 (.in(n12857), .out(n12857_0));
mux3 mux_7692 (.in({n9745_0, n9744_0, n2524}), .out(n12858), .config_in(config_chain[27919:27918]), .config_rst(config_rst)); 
buffer_wire buffer_12858 (.in(n12858), .out(n12858_0));
mux15 mux_7693 (.in({n12891_1, n10051_1, n10030_0, n10027_0, n10007_2, n9970_0, n9955_0, n9944_0, n9929_0, n9926_0, n2532, n2524, n2516, n1548, n1540}), .out(n12859), .config_in(config_chain[27925:27920]), .config_rst(config_rst)); 
buffer_wire buffer_12859 (.in(n12859), .out(n12859_0));
mux3 mux_7694 (.in({n9747_1, n9746_0, n2528}), .out(n12860), .config_in(config_chain[27927:27926]), .config_rst(config_rst)); 
buffer_wire buffer_12860 (.in(n12860), .out(n12860_0));
mux13 mux_7695 (.in({n12993_0, n11353_2, n11317_0, n11306_0, n11303_0, n11278_0, n11273_0, n11248_0, n11220_0, n3018, n3010, n2042, n2034}), .out(n12861), .config_in(config_chain[27933:27928]), .config_rst(config_rst)); 
buffer_wire buffer_12861 (.in(n12861), .out(n12861_0));
mux3 mux_7696 (.in({n9749_2, n9748_0, n2528}), .out(n12862), .config_in(config_chain[27935:27934]), .config_rst(config_rst)); 
buffer_wire buffer_12862 (.in(n12862), .out(n12862_0));
mux13 mux_7697 (.in({n13015_0, n11619_2, n11597_2, n11590_0, n11570_0, n11537_0, n11512_0, n11507_0, n11486_0, n3116, n3108, n2140/**/, n2132}), .out(n12863), .config_in(config_chain[27941:27936]), .config_rst(config_rst)); 
buffer_wire buffer_12863 (.in(n12863), .out(n12863_0));
mux3 mux_7698 (.in({n9751_2, n9750_0, n2528}), .out(n12864), .config_in(config_chain[27943:27942]), .config_rst(config_rst)); 
buffer_wire buffer_12864 (.in(n12864), .out(n12864_0));
mux13 mux_7699 (.in({n13037_0, n11883_2, n11853_0, n11846_0, n11834_0, n11829_2, n11804_0/**/, n11771_0, n11752_0, n3214, n3206, n2238, n2230}), .out(n12865), .config_in(config_chain[27949:27944]), .config_rst(config_rst)); 
buffer_wire buffer_12865 (.in(n12865), .out(n12865_0));
mux3 mux_7700 (.in({n9753_2, n9752_0, n2528}), .out(n12866), .config_in(config_chain[27951:27950]), .config_rst(config_rst)); 
buffer_wire buffer_12866 (.in(n12866), .out(n12866_0));
mux3 mux_7701 (.in({n12145_2, n12096_0, n3312}), .out(n12867), .config_in(config_chain[27953:27952]), .config_rst(config_rst)); 
buffer_wire buffer_12867 (.in(n12867), .out(n12867_0));
mux3 mux_7702 (.in({n9755_2, n9754_0, n2528}), .out(n12868), .config_in(config_chain[27955:27954]), .config_rst(config_rst)); 
buffer_wire buffer_12868 (.in(n12868), .out(n12868_0));
mux3 mux_7703 (.in({n12099_0, n12098_0/**/, n3312}), .out(n12869), .config_in(config_chain[27957:27956]), .config_rst(config_rst)); 
buffer_wire buffer_12869 (.in(n12869), .out(n12869_0));
mux3 mux_7704 (.in({n9757_2, n9756_0, n2532}), .out(n12870), .config_in(config_chain[27959:27958]), .config_rst(config_rst)); 
buffer_wire buffer_12870 (.in(n12870), .out(n12870_0));
mux3 mux_7705 (.in({n12101_0/**/, n12100_0, n3316}), .out(n12871), .config_in(config_chain[27961:27960]), .config_rst(config_rst)); 
buffer_wire buffer_12871 (.in(n12871), .out(n12871_0));
mux16 mux_7706 (.in({n12786_0, n10035_1, n10025_0, n10020_0, n10008_0, n10001_1, n9984_0, n9947_0, n9930_0/**/, n9926_0, n9921_0, n2626, n2618, n1650, n1642, n1634}), .out(n12872), .config_in(config_chain[27967:27962]), .config_rst(config_rst)); 
buffer_wire buffer_12872 (.in(n12872), .out(n12872_0));
mux16 mux_7707 (.in({n12953_1, n11085_1, n11060_0, n11057_0, n11045_1, n11036_0, n11021_0, n10982_0, n10970_0, n10967_0, n10956_0/**/, n2920, n2912, n1944, n1936, n1928}), .out(n12873), .config_in(config_chain[27973:27968]), .config_rst(config_rst)); 
buffer_wire buffer_12873 (.in(n12873), .out(n12873_0));
mux16 mux_7708 (.in({n12794_0, n10037_1/**/, n10019_0, n10014_0, n10010_0, n10003_1, n9998_0, n9986_0, n9977_0, n9960_0, n9923_0, n2626, n2618, n1650, n1642, n1634}), .out(n12874), .config_in(config_chain[27979:27974]), .config_rst(config_rst)); 
buffer_wire buffer_12874 (.in(n12874), .out(n12874_0));
mux16 mux_7709 (.in({n12955_1, n11083_1/**/, n11054_0, n11051_0, n11047_1, n11038_0, n11023_0, n11012_0, n10997_0, n10978_0, n10958_0, n2920, n2912, n1944, n1936, n1928}), .out(n12875), .config_in(config_chain[27985:27980]), .config_rst(config_rst)); 
buffer_wire buffer_12875 (.in(n12875), .out(n12875_0));
mux15 mux_7710 (.in({n12802_0, n10039_1/**/, n10028_0, n10013_0, n10005_2, n9990_0, n9979_0, n9962_0, n9953_0, n9936_0, n2626, n2618, n1650, n1642, n1634}), .out(n12876), .config_in(config_chain[27991:27986]), .config_rst(config_rst)); 
buffer_wire buffer_12876 (.in(n12876), .out(n12876_0));
mux15 mux_7711 (.in({n12957_1, n11081_1, n11065_0, n11048_0/**/, n11040_0, n11014_0, n10999_0, n10988_0, n10986_0, n10973_0, n2920, n2912, n1944, n1936, n1928}), .out(n12877), .config_in(config_chain[27997:27992]), .config_rst(config_rst)); 
buffer_wire buffer_12877 (.in(n12877), .out(n12877_0));
mux15 mux_7712 (.in({n12810_0, n10041_1, n10027_0, n10022_0, n10007_2, n9992_0/**/, n9982_0, n9955_0, n9938_0, n9929_0, n2626, n2618, n1650, n1642, n1634}), .out(n12878), .config_in(config_chain[28003:27998]), .config_rst(config_rst)); 
buffer_wire buffer_12878 (.in(n12878), .out(n12878_0));
mux15 mux_7713 (.in({n12959_1, n11079_1, n11062_0, n11059_0, n11042_0, n11029_0/**/, n10994_0, n10990_0, n10975_0, n10964_0, n2920, n2912, n1944, n1936, n1928}), .out(n12879), .config_in(config_chain[28009:28004]), .config_rst(config_rst)); 
buffer_wire buffer_12879 (.in(n12879), .out(n12879_0));
mux15 mux_7714 (.in({n12818_0, n10043_1, n10021_0, n10016_0, n10009_2, n9994_0, n9985_0, n9974_0, n9968_0, n9931_0, n2626/**/, n2618, n1650, n1642, n1634}), .out(n12880), .config_in(config_chain[28015:28010]), .config_rst(config_rst)); 
buffer_wire buffer_12880 (.in(n12880), .out(n12880_0));
mux15 mux_7715 (.in({n12961_1, n11077_1, n11056_0, n11053_0, n11044_0, n11031_0, n11020_0, n11005_0, n11002_0, n10966_0, n2920, n2912, n1944, n1936, n1928}), .out(n12881), .config_in(config_chain[28021:28016]), .config_rst(config_rst)); 
buffer_wire buffer_12881 (.in(n12881), .out(n12881_0));
mux15 mux_7716 (.in({n12826_0, n10045_1, n10030_0, n10015_0, n10011_2, n9987_0, n9970_0, n9966_0, n9961_0, n9944_0, n2630, n2622, n2614, n1646, n1638}), .out(n12882), .config_in(config_chain[28027:28022]), .config_rst(config_rst)); 
buffer_wire buffer_12882 (.in(n12882), .out(n12882_0));
mux15 mux_7717 (.in({n12963_1, n11075_1, n11067_0, n11050_0, n11046_0, n11022_0, n11010_0, n11007_0, n10996_0, n10981_0, n2924, n2916, n2908, n1940, n1932}), .out(n12883), .config_in(config_chain[28033:28028]), .config_rst(config_rst)); 
buffer_wire buffer_12883 (.in(n12883), .out(n12883_0));
mux15 mux_7718 (.in({n12834_0, n10047_1, n10029_0, n10024_0, n10000_0, n9963_0/**/, n9958_0, n9946_0, n9937_0, n9920_0, n2630, n2622, n2614, n1646, n1638}), .out(n12884), .config_in(config_chain[28039:28034]), .config_rst(config_rst)); 
buffer_wire buffer_12884 (.in(n12884), .out(n12884_0));
mux15 mux_7719 (.in({n12965_1, n11073_1, n11064_0, n11061_0, n11037_0, n11018_0, n10998_0, n10983_0, n10972_0, n10957_0, n2924, n2916, n2908, n1940, n1932}), .out(n12885), .config_in(config_chain[28045:28040]), .config_rst(config_rst)); 
buffer_wire buffer_12885 (.in(n12885), .out(n12885_0));
mux15 mux_7720 (.in({n12842_0/**/, n10049_1, n10023_0, n10018_0, n10002_0, n9993_0, n9976_0, n9950_0, n9939_0, n9922_0, n2630, n2622, n2614, n1646, n1638}), .out(n12886), .config_in(config_chain[28051:28046]), .config_rst(config_rst)); 
buffer_wire buffer_12886 (.in(n12886), .out(n12886_0));
mux15 mux_7721 (.in({n12967_1, n11071_1, n11058_0, n11055_0, n11039_0, n11028_0, n11026_0/**/, n11013_0, n10974_0, n10959_0, n2924, n2916, n2908, n1940, n1932}), .out(n12887), .config_in(config_chain[28057:28052]), .config_rst(config_rst)); 
buffer_wire buffer_12887 (.in(n12887), .out(n12887_0));
mux15 mux_7722 (.in({n12850_0, n10051_1, n10017_0, n10012_0, n10004_0, n9995_0, n9978_0, n9969_0, n9952_0, n9942_0, n2630, n2622/**/, n2614, n1646, n1638}), .out(n12888), .config_in(config_chain[28063:28058]), .config_rst(config_rst)); 
buffer_wire buffer_12888 (.in(n12888), .out(n12888_0));
mux15 mux_7723 (.in({n12969_1, n11069_1, n11052_0, n11049_0, n11041_0, n11034_0, n11030_0, n11015_0, n11004_0, n10989_0/**/, n2924, n2916, n2908, n1940, n1932}), .out(n12889), .config_in(config_chain[28069:28064]), .config_rst(config_rst)); 
buffer_wire buffer_12889 (.in(n12889), .out(n12889_0));
mux15 mux_7724 (.in({n12858_0, n10033_1, n10031_0, n10026_0, n10006_0, n9971_0, n9954_0, n9945_0, n9934_0, n9928_0, n2630/**/, n2622, n2614, n1646, n1638}), .out(n12890), .config_in(config_chain[28075:28070]), .config_rst(config_rst)); 
buffer_wire buffer_12890 (.in(n12890), .out(n12890_0));
mux15 mux_7725 (.in({n12971_1, n11087_1, n11066_0, n11063_0/**/, n11043_1, n11006_0, n10991_0, n10980_0, n10965_0, n10962_0, n2924, n2916, n2908, n1940, n1932}), .out(n12891), .config_in(config_chain[28081:28076]), .config_rst(config_rst)); 
buffer_wire buffer_12891 (.in(n12891), .out(n12891_0));
mux16 mux_7726 (.in({n12780_0, n10291_1, n10281_0, n10276_0, n10264_0, n10257_1, n10242_0, n10205_0, n10188_0, n10179_0, n10176_0, n2724, n2716, n1748, n1740, n1732/**/}), .out(n12892), .config_in(config_chain[28087:28082]), .config_rst(config_rst)); 
buffer_wire buffer_12892 (.in(n12892), .out(n12892_0));
mux15 mux_7727 (.in({n12973_0, n11351_1, n11325_0, n11318_0, n11308_0, n11305_0, n11280_0, n11247_0, n11228_0, n11222_0, n3018, n3010, n2042, n2034, n2026}), .out(n12893), .config_in(config_chain[28093:28088]), .config_rst(config_rst)); 
buffer_wire buffer_12893 (.in(n12893), .out(n12893_0));
mux16 mux_7728 (.in({n12788_0, n10293_1/**/, n10275_0, n10270_0, n10266_0, n10259_1, n10248_0, n10244_0, n10235_0, n10218_0, n10181_0, n2724, n2716, n1748, n1740, n1732}), .out(n12894), .config_in(config_chain[28099:28094]), .config_rst(config_rst)); 
buffer_wire buffer_12894 (.in(n12894), .out(n12894_0));
mux15 mux_7729 (.in({n12975_0, n11349_1, n11326_0, n11310_0, n11307_0, n11279_0/**/, n11254_0, n11249_0, n11236_0, n11224_0, n3022, n3010, n2042, n2034, n2026}), .out(n12895), .config_in(config_chain[28105:28100]), .config_rst(config_rst)); 
buffer_wire buffer_12895 (.in(n12895), .out(n12895_0));
mux15 mux_7730 (.in({n12796_0, n10295_1, n10284_0, n10269_0, n10261_1, n10240_0, n10237_0, n10220_0, n10211_0/**/, n10194_0, n2724, n2716, n1748, n1740, n1732}), .out(n12896), .config_in(config_chain[28111:28106]), .config_rst(config_rst)); 
buffer_wire buffer_12896 (.in(n12896), .out(n12896_0));
mux15 mux_7731 (.in({n12977_0, n11347_1, n11319_0, n11312_0, n11309_1, n11286_0, n11281_0, n11256_0, n11244_0, n11223_0, n3022/**/, n3014, n2042, n2034, n2026}), .out(n12897), .config_in(config_chain[28117:28112]), .config_rst(config_rst)); 
buffer_wire buffer_12897 (.in(n12897), .out(n12897_0));
mux15 mux_7732 (.in({n12804_0, n10297_1, n10283_0, n10278_0, n10263_2, n10250_0, n10232_0, n10213_0/**/, n10196_0, n10187_0, n2724, n2716, n1748, n1740, n1732}), .out(n12898), .config_in(config_chain[28123:28118]), .config_rst(config_rst)); 
buffer_wire buffer_12898 (.in(n12898), .out(n12898_0));
mux15 mux_7733 (.in({n12979_0/**/, n11345_1, n11327_0, n11320_0, n11311_1, n11288_0, n11255_0, n11252_0, n11230_0, n11225_0, n3022, n3014, n3006, n2034, n2026}), .out(n12899), .config_in(config_chain[28129:28124]), .config_rst(config_rst)); 
buffer_wire buffer_12899 (.in(n12899), .out(n12899_0));
mux15 mux_7734 (.in({n12812_0, n10299_1, n10277_0, n10272_0, n10265_2, n10252_0, n10243_0, n10226_0/**/, n10224_0, n10189_0, n2724, n2716, n1748, n1740, n1732}), .out(n12900), .config_in(config_chain[28135:28130]), .config_rst(config_rst)); 
buffer_wire buffer_12900 (.in(n12900), .out(n12900_0));
mux14 mux_7735 (.in({n12981_0/**/, n11343_1, n11328_0, n11313_0, n11287_0, n11262_0, n11260_0, n11257_0, n11232_0, n3022, n3014, n3006, n2038, n2026}), .out(n12901), .config_in(config_chain[28141:28136]), .config_rst(config_rst)); 
buffer_wire buffer_12901 (.in(n12901), .out(n12901_0));
mux15 mux_7736 (.in({n12820_0, n10301_1, n10286_0, n10271_0, n10267_2, n10245_0, n10228_0, n10219_0, n10216_0, n10202_0, n2728/**/, n2720, n2712, n1744, n1736}), .out(n12902), .config_in(config_chain[28147:28142]), .config_rst(config_rst)); 
buffer_wire buffer_12902 (.in(n12902), .out(n12902_0));
mux14 mux_7737 (.in({n12983_0, n11341_1/**/, n11321_0, n11314_0, n11294_0, n11289_0, n11268_0, n11264_0, n11231_0, n3022, n3014, n3006, n2038, n2030}), .out(n12903), .config_in(config_chain[28153:28148]), .config_rst(config_rst)); 
buffer_wire buffer_12903 (.in(n12903), .out(n12903_0));
mux15 mux_7738 (.in({n12828_0, n10303_1, n10285_0, n10280_0, n10256_0, n10221_0, n10208_0, n10204_0, n10195_0/**/, n10178_0, n2728, n2720, n2712, n1744, n1736}), .out(n12904), .config_in(config_chain[28159:28154]), .config_rst(config_rst)); 
buffer_wire buffer_12904 (.in(n12904), .out(n12904_0));
mux13 mux_7739 (.in({n12985_0, n11339_1, n11329_0, n11322_0/**/, n11296_0, n11276_0, n11263_0, n11238_0, n11233_0, n3014, n3006, n2038, n2030}), .out(n12905), .config_in(config_chain[28165:28160]), .config_rst(config_rst)); 
buffer_wire buffer_12905 (.in(n12905), .out(n12905_0));
mux15 mux_7740 (.in({n12836_0, n10305_1, n10279_0, n10274_0, n10258_0, n10251_0, n10234_0, n10200_0, n10197_0, n10180_0, n2728, n2720/**/, n2712, n1744, n1736}), .out(n12906), .config_in(config_chain[28171:28166]), .config_rst(config_rst)); 
buffer_wire buffer_12906 (.in(n12906), .out(n12906_0));
mux13 mux_7741 (.in({n12987_0/**/, n11337_1, n11330_0, n11315_0, n11295_0, n11284_0, n11270_0, n11265_0, n11240_0, n3018, n3006, n2038, n2030}), .out(n12907), .config_in(config_chain[28177:28172]), .config_rst(config_rst)); 
buffer_wire buffer_12907 (.in(n12907), .out(n12907_0));
mux15 mux_7742 (.in({n12844_0, n10307_1, n10273_0, n10268_0, n10260_0, n10253_0, n10236_0, n10227_0, n10210_0, n10192_0, n2728, n2720, n2712, n1744, n1736/**/}), .out(n12908), .config_in(config_chain[28183:28178]), .config_rst(config_rst)); 
buffer_wire buffer_12908 (.in(n12908), .out(n12908_0));
mux13 mux_7743 (.in({n12989_0, n11335_1, n11323_0, n11316_0, n11302_0, n11297_0, n11292_0, n11272_0, n11239_0, n3018, n3010, n2038, n2030}), .out(n12909), .config_in(config_chain[28189:28184]), .config_rst(config_rst)); 
buffer_wire buffer_12909 (.in(n12909), .out(n12909_0));
mux15 mux_7744 (.in({n12852_0, n10289_1, n10287_0, n10282_0, n10262_0, n10229_0/**/, n10212_0, n10203_0, n10186_0, n10184_0, n2728, n2720, n2712, n1744, n1736}), .out(n12910), .config_in(config_chain[28195:28190]), .config_rst(config_rst)); 
buffer_wire buffer_12910 (.in(n12910), .out(n12910_0));
mux13 mux_7745 (.in({n12991_0, n11333_1, n11331_0/**/, n11324_0, n11304_0, n11300_0, n11271_0, n11246_0, n11241_0, n3018, n3010, n2042, n2030}), .out(n12911), .config_in(config_chain[28201:28196]), .config_rst(config_rst)); 
buffer_wire buffer_12911 (.in(n12911), .out(n12911_0));
mux16 mux_7746 (.in({n12782_0, n10549_1, n10542_0, n10527_0, n10522_0, n10515_0, n10489_0/**/, n10472_0, n10463_0, n10446_0, n10436_0, n2822, n2814, n1846, n1838, n1830}), .out(n12912), .config_in(config_chain[28207:28202]), .config_rst(config_rst)); 
buffer_wire buffer_12912 (.in(n12912), .out(n12912_0));
mux15 mux_7747 (.in({n12995_0, n11617_1, n11583_0, n11576_0, n11572_0, n11569_0, n11544_0, n11539_0, n11514_0, n11494_0, n3116, n3108, n2140, n2132, n2124}), .out(n12913), .config_in(config_chain[28213:28208]), .config_rst(config_rst)); 
buffer_wire buffer_12913 (.in(n12913), .out(n12913_0));
mux16 mux_7748 (.in({n12790_0, n10551_1, n10541_0, n10536_0, n10524_0, n10517_1, n10508_0/**/, n10502_0, n10465_0, n10448_0, n10439_0, n2822, n2814, n1846, n1838, n1830}), .out(n12914), .config_in(config_chain[28219:28214]), .config_rst(config_rst)); 
buffer_wire buffer_12914 (.in(n12914), .out(n12914_0));
mux15 mux_7749 (.in({n12997_0, n11615_1, n11591_0, n11584_0, n11574_0, n11571_0, n11546_0, n11513_0, n11502_0, n11488_0, n3120, n3108, n2140, n2132, n2124}), .out(n12915), .config_in(config_chain[28225:28220]), .config_rst(config_rst)); 
buffer_wire buffer_12915 (.in(n12915), .out(n12915_0));
mux15 mux_7750 (.in({n12798_0, n10553_1, n10535_0/**/, n10530_0, n10519_1, n10504_0, n10500_0, n10495_0, n10478_0, n10441_0, n2822, n2814, n1846, n1838, n1830}), .out(n12916), .config_in(config_chain[28231:28226]), .config_rst(config_rst)); 
buffer_wire buffer_12916 (.in(n12916), .out(n12916_0));
mux15 mux_7751 (.in({n12999_0, n11613_1, n11592_0, n11577_0, n11573_0, n11545_0, n11520_0, n11515_0, n11510_0, n11490_0, n3120, n3112, n2140, n2132, n2124}), .out(n12917), .config_in(config_chain[28237:28232]), .config_rst(config_rst)); 
buffer_wire buffer_12917 (.in(n12917), .out(n12917_0));
mux15 mux_7752 (.in({n12806_0, n10555_1, n10544_0, n10529_0, n10521_1, n10497_0, n10492_0, n10480_0, n10471_0, n10454_0, n2822/**/, n2814, n1846, n1838, n1830}), .out(n12918), .config_in(config_chain[28243:28238]), .config_rst(config_rst)); 
buffer_wire buffer_12918 (.in(n12918), .out(n12918_0));
mux15 mux_7753 (.in({n13001_0, n11611_1, n11585_0, n11578_0, n11575_1, n11552_0, n11547_0, n11522_0, n11518_0, n11489_0/**/, n3120, n3112, n3104, n2132, n2124}), .out(n12919), .config_in(config_chain[28249:28244]), .config_rst(config_rst)); 
buffer_wire buffer_12919 (.in(n12919), .out(n12919_0));
mux15 mux_7754 (.in({n12814_0/**/, n10557_1, n10543_0, n10538_0, n10523_2, n10510_0, n10484_0, n10473_0, n10456_0, n10447_0, n2822, n2814, n1846, n1838, n1830}), .out(n12920), .config_in(config_chain[28255:28250]), .config_rst(config_rst)); 
buffer_wire buffer_12920 (.in(n12920), .out(n12920_0));
mux14 mux_7755 (.in({n13003_0, n11609_1, n11593_0, n11586_0, n11554_0, n11526_0, n11521_0, n11496_0, n11491_0, n3120/**/, n3112, n3104, n2136, n2124}), .out(n12921), .config_in(config_chain[28261:28256]), .config_rst(config_rst)); 
buffer_wire buffer_12921 (.in(n12921), .out(n12921_0));
mux15 mux_7756 (.in({n12822_0/**/, n10559_1, n10537_0, n10532_0, n10525_2, n10512_0, n10503_0, n10486_0, n10476_0, n10449_0, n2826, n2818, n2810, n1842, n1834}), .out(n12922), .config_in(config_chain[28267:28262]), .config_rst(config_rst)); 
buffer_wire buffer_12922 (.in(n12922), .out(n12922_0));
mux14 mux_7757 (.in({n13005_0, n11607_1, n11594_0, n11579_0, n11553_0, n11534_0, n11528_0, n11523_0, n11498_0, n3120, n3112, n3104, n2136, n2128}), .out(n12923), .config_in(config_chain[28273:28268]), .config_rst(config_rst)); 
buffer_wire buffer_12923 (.in(n12923), .out(n12923_0));
mux15 mux_7758 (.in({n12830_0, n10561_1, n10531_0, n10526_0, n10514_0, n10505_0, n10488_0, n10479_0, n10468_0, n10462_0, n2826, n2818, n2810/**/, n1842, n1834}), .out(n12924), .config_in(config_chain[28279:28274]), .config_rst(config_rst)); 
buffer_wire buffer_12924 (.in(n12924), .out(n12924_0));
mux13 mux_7759 (.in({n13007_0, n11605_1, n11587_0, n11580_0, n11560_0, n11555_0, n11542_0, n11530_0, n11497_0, n3112, n3104/**/, n2136, n2128}), .out(n12925), .config_in(config_chain[28285:28280]), .config_rst(config_rst)); 
buffer_wire buffer_12925 (.in(n12925), .out(n12925_0));
mux15 mux_7760 (.in({n12838_0, n10563_1, n10545_0, n10540_0, n10516_0, n10481_0/**/, n10464_0, n10460_0, n10455_0, n10438_0, n2826, n2818, n2810, n1842, n1834}), .out(n12926), .config_in(config_chain[28291:28286]), .config_rst(config_rst)); 
buffer_wire buffer_12926 (.in(n12926), .out(n12926_0));
mux13 mux_7761 (.in({n13009_0, n11603_1, n11595_0, n11588_0, n11562_0, n11550_0, n11529_0/**/, n11504_0, n11499_0, n3116, n3104, n2136, n2128}), .out(n12927), .config_in(config_chain[28297:28292]), .config_rst(config_rst)); 
buffer_wire buffer_12927 (.in(n12927), .out(n12927_0));
mux15 mux_7762 (.in({n12846_0/**/, n10565_1, n10539_0, n10534_0, n10518_0, n10511_0, n10494_0, n10457_0, n10452_0, n10440_0, n2826, n2818, n2810, n1842, n1834}), .out(n12928), .config_in(config_chain[28303:28298]), .config_rst(config_rst)); 
buffer_wire buffer_12928 (.in(n12928), .out(n12928_0));
mux13 mux_7763 (.in({n13011_0, n11601_1, n11596_0, n11581_0, n11561_0, n11558_0, n11536_0, n11531_0, n11506_0, n3116, n3108, n2136, n2128}), .out(n12929), .config_in(config_chain[28309:28304]), .config_rst(config_rst)); 
buffer_wire buffer_12929 (.in(n12929), .out(n12929_0));
mux15 mux_7764 (.in({n12854_0/**/, n10547_1, n10533_0, n10528_0, n10520_0, n10513_0, n10496_0, n10487_0, n10470_0, n10444_0, n2826, n2818, n2810, n1842, n1834}), .out(n12930), .config_in(config_chain[28315:28310]), .config_rst(config_rst)); 
buffer_wire buffer_12930 (.in(n12930), .out(n12930_0));
mux13 mux_7765 (.in({n13013_0, n11599_1, n11589_0, n11582_0, n11568_0, n11566_0, n11563_0/**/, n11538_0, n11505_0, n3116, n3108, n2140, n2128}), .out(n12931), .config_in(config_chain[28321:28316]), .config_rst(config_rst)); 
buffer_wire buffer_12931 (.in(n12931), .out(n12931_0));
mux16 mux_7766 (.in({n12784_1, n10809_1, n10793_0, n10788_0, n10782_0, n10775_0, n10758_0, n10749_0, n10732_0, n10698_0, n10695_0/**/, n2920, n2912, n1944, n1936, n1928}), .out(n12932), .config_in(config_chain[28327:28322]), .config_rst(config_rst)); 
buffer_wire buffer_12932 (.in(n12932), .out(n12932_0));
mux15 mux_7767 (.in({n13017_0, n11881_1, n11861_2, n11854_0, n11836_0, n11803_0, n11778_0, n11773_0, n11760_0, n11748_0, n3214, n3206/**/, n2238, n2230, n2222}), .out(n12933), .config_in(config_chain[28333:28328]), .config_rst(config_rst)); 
buffer_wire buffer_12933 (.in(n12933), .out(n12933_0));
mux16 mux_7768 (.in({n12792_1/**/, n10811_1, n10802_0, n10787_0, n10784_0, n10777_0, n10770_0, n10751_0, n10734_0, n10725_0, n10708_0, n2920, n2912, n1944, n1936, n1928}), .out(n12934), .config_in(config_chain[28339:28334]), .config_rst(config_rst)); 
buffer_wire buffer_12934 (.in(n12934), .out(n12934_0));
mux15 mux_7769 (.in({n13019_0, n11879_1, n11847_0, n11840_0, n11838_0, n11835_0, n11810_0, n11805_0, n11780_0, n11768_0, n3218/**/, n3206, n2238, n2230, n2222}), .out(n12935), .config_in(config_chain[28345:28340]), .config_rst(config_rst)); 
buffer_wire buffer_12935 (.in(n12935), .out(n12935_0));
mux15 mux_7770 (.in({n12800_1, n10813_1, n10801_0, n10796_0, n10779_1, n10764_0, n10762_0, n10727_0, n10710_0, n10701_0/**/, n2920, n2912, n1944, n1936, n1928}), .out(n12936), .config_in(config_chain[28351:28346]), .config_rst(config_rst)); 
buffer_wire buffer_12936 (.in(n12936), .out(n12936_0));
mux15 mux_7771 (.in({n13021_0, n11877_1, n11855_0, n11848_0, n11837_0, n11812_0/**/, n11779_0, n11776_0, n11754_0, n11749_0, n3218, n3210, n2238, n2230, n2222}), .out(n12937), .config_in(config_chain[28357:28352]), .config_rst(config_rst)); 
buffer_wire buffer_12937 (.in(n12937), .out(n12937_0));
mux15 mux_7772 (.in({n12808_1, n10815_1, n10795_0, n10790_0/**/, n10781_1, n10766_0, n10757_0, n10754_0, n10740_0, n10703_0, n2920, n2912, n1944, n1936, n1928}), .out(n12938), .config_in(config_chain[28363:28358]), .config_rst(config_rst)); 
buffer_wire buffer_12938 (.in(n12938), .out(n12938_0));
mux15 mux_7773 (.in({n13023_0, n11875_1, n11856_0, n11841_0, n11839_0, n11811_0, n11786_0, n11784_0, n11781_0, n11756_0, n3218, n3210, n3202, n2230, n2222/**/}), .out(n12939), .config_in(config_chain[28369:28364]), .config_rst(config_rst)); 
buffer_wire buffer_12939 (.in(n12939), .out(n12939_0));
mux15 mux_7774 (.in({n12816_1, n10817_1, n10804_0, n10789_0, n10783_1, n10759_0, n10746_0, n10742_0, n10733_0, n10716_0, n2920/**/, n2912, n1944, n1936, n1928}), .out(n12940), .config_in(config_chain[28375:28370]), .config_rst(config_rst)); 
buffer_wire buffer_12940 (.in(n12940), .out(n12940_0));
mux14 mux_7775 (.in({n13025_0, n11873_1, n11849_0, n11842_0, n11818_0, n11813_0, n11792_0, n11788_0, n11755_0/**/, n3218, n3210, n3202, n2234, n2222}), .out(n12941), .config_in(config_chain[28381:28376]), .config_rst(config_rst)); 
buffer_wire buffer_12941 (.in(n12941), .out(n12941_0));
mux15 mux_7776 (.in({n12824_1, n10819_1, n10803_0, n10798_0, n10785_2, n10772_0, n10738_0, n10735_0, n10718_0, n10709_0, n2924, n2916, n2908, n1940, n1932/**/}), .out(n12942), .config_in(config_chain[28387:28382]), .config_rst(config_rst)); 
buffer_wire buffer_12942 (.in(n12942), .out(n12942_0));
mux14 mux_7777 (.in({n13027_0/**/, n11871_1, n11857_0, n11850_0, n11820_0, n11800_0, n11787_0, n11762_0, n11757_0, n3218, n3210, n3202, n2234, n2226}), .out(n12943), .config_in(config_chain[28393:28388]), .config_rst(config_rst)); 
buffer_wire buffer_12943 (.in(n12943), .out(n12943_0));
mux15 mux_7778 (.in({n12832_1, n10821_1, n10797_0, n10792_0, n10774_0, n10765_0, n10748_0, n10730_0, n10711_0, n10694_0, n2924, n2916/**/, n2908, n1940, n1932}), .out(n12944), .config_in(config_chain[28399:28394]), .config_rst(config_rst)); 
buffer_wire buffer_12944 (.in(n12944), .out(n12944_0));
mux13 mux_7779 (.in({n13029_0, n11869_1, n11858_0, n11843_0/**/, n11819_0, n11808_0, n11794_0, n11789_0, n11764_0, n3210, n3202, n2234, n2226}), .out(n12945), .config_in(config_chain[28405:28400]), .config_rst(config_rst)); 
buffer_wire buffer_12945 (.in(n12945), .out(n12945_0));
mux15 mux_7780 (.in({n12840_1, n10823_1, n10791_0/**/, n10786_0, n10776_0, n10767_0, n10750_0, n10741_0, n10724_0, n10722_0, n2924, n2916, n2908, n1940, n1932}), .out(n12946), .config_in(config_chain[28411:28406]), .config_rst(config_rst)); 
buffer_wire buffer_12946 (.in(n12946), .out(n12946_0));
mux13 mux_7781 (.in({n13031_0/**/, n11867_1, n11851_0, n11844_0, n11826_0, n11821_0, n11816_0, n11796_0, n11763_0, n3214, n3202, n2234, n2226}), .out(n12947), .config_in(config_chain[28417:28412]), .config_rst(config_rst)); 
buffer_wire buffer_12947 (.in(n12947), .out(n12947_0));
mux15 mux_7782 (.in({n12848_1, n10825_1, n10805_0, n10800_0, n10778_0, n10743_0, n10726_0, n10717_0, n10714_0, n10700_0, n2924/**/, n2916, n2908, n1940, n1932}), .out(n12948), .config_in(config_chain[28423:28418]), .config_rst(config_rst)); 
buffer_wire buffer_12948 (.in(n12948), .out(n12948_0));
mux13 mux_7783 (.in({n13033_0/**/, n11865_1, n11859_0, n11852_0, n11828_0, n11824_0, n11795_0, n11770_0, n11765_0, n3214, n3206, n2234, n2226}), .out(n12949), .config_in(config_chain[28429:28424]), .config_rst(config_rst)); 
buffer_wire buffer_12949 (.in(n12949), .out(n12949_0));
mux15 mux_7784 (.in({n12856_1, n10807_1, n10799_0, n10794_0, n10780_0, n10773_0/**/, n10756_0, n10719_0, n10706_0, n10702_0, n2924, n2916, n2908, n1940, n1932}), .out(n12950), .config_in(config_chain[28435:28430]), .config_rst(config_rst)); 
buffer_wire buffer_12950 (.in(n12950), .out(n12950_0));
mux13 mux_7785 (.in({n13035_0/**/, n11863_1, n11860_0, n11845_0, n11832_0, n11827_0, n11802_0, n11797_0, n11772_0, n3214, n3206, n2238, n2226}), .out(n12951), .config_in(config_chain[28441:28436]), .config_rst(config_rst)); 
buffer_wire buffer_12951 (.in(n12951), .out(n12951_0));
mux16 mux_7786 (.in({n12872_1, n11071_1, n11061_0, n11056_0, n11044_0, n11037_0, n11020_0, n10983_0, n10966_0, n10962_0, n10957_0, n3018, n3010, n2042, n2034, n2026}), .out(n12952), .config_in(config_chain[28447:28442]), .config_rst(config_rst)); 
buffer_wire buffer_12952 (.in(n12952), .out(n12952_0));
mux4 mux_7787 (.in({n12125_1, n12016_0, n3316, n2320}), .out(n12953), .config_in(config_chain[28449:28448]), .config_rst(config_rst)); 
buffer_wire buffer_12953 (.in(n12953), .out(n12953_0));
mux16 mux_7788 (.in({n12874_1/**/, n11073_1, n11055_0, n11050_0, n11046_0, n11039_0, n11034_0, n11022_0, n11013_0, n10996_0, n10959_0, n3018, n3010, n2042, n2034, n2026}), .out(n12954), .config_in(config_chain[28455:28450]), .config_rst(config_rst)); 
buffer_wire buffer_12954 (.in(n12954), .out(n12954_0));
mux3 mux_7789 (.in({n12127_1, n12024_0/**/, n2324}), .out(n12955), .config_in(config_chain[28457:28456]), .config_rst(config_rst)); 
buffer_wire buffer_12955 (.in(n12955), .out(n12955_0));
mux15 mux_7790 (.in({n12876_1, n11075_1, n11064_0, n11049_0, n11041_0, n11026_0/**/, n11015_0, n10998_0, n10989_0, n10972_0, n3018, n3010, n2042, n2034, n2026}), .out(n12956), .config_in(config_chain[28463:28458]), .config_rst(config_rst)); 
buffer_wire buffer_12956 (.in(n12956), .out(n12956_0));
mux3 mux_7791 (.in({n12129_1, n12032_0, n2328}), .out(n12957), .config_in(config_chain[28465:28464]), .config_rst(config_rst)); 
buffer_wire buffer_12957 (.in(n12957), .out(n12957_0));
mux15 mux_7792 (.in({n12878_1, n11077_1, n11063_0, n11058_0, n11043_1, n11028_0, n11018_0, n10991_0/**/, n10974_0, n10965_0, n3018, n3010, n2042, n2034, n2026}), .out(n12958), .config_in(config_chain[28471:28466]), .config_rst(config_rst)); 
buffer_wire buffer_12958 (.in(n12958), .out(n12958_0));
mux3 mux_7793 (.in({n12131_1, n12040_0, n2332}), .out(n12959), .config_in(config_chain[28473:28472]), .config_rst(config_rst)); 
buffer_wire buffer_12959 (.in(n12959), .out(n12959_0));
mux15 mux_7794 (.in({n12880_1, n11079_1, n11057_0, n11052_0, n11045_1, n11030_0, n11021_0, n11010_0, n11004_0, n10967_0, n3018/**/, n3010, n2042, n2034, n2026}), .out(n12960), .config_in(config_chain[28479:28474]), .config_rst(config_rst)); 
buffer_wire buffer_12960 (.in(n12960), .out(n12960_0));
mux3 mux_7795 (.in({n12133_1, n12048_0/**/, n2332}), .out(n12961), .config_in(config_chain[28481:28480]), .config_rst(config_rst)); 
buffer_wire buffer_12961 (.in(n12961), .out(n12961_0));
mux15 mux_7796 (.in({n12882_1, n11081_1, n11066_0, n11051_0, n11047_1, n11023_0, n11006_0, n11002_0, n10997_0, n10980_0, n3022, n3014, n3006, n2038, n2030/**/}), .out(n12962), .config_in(config_chain[28487:28482]), .config_rst(config_rst)); 
buffer_wire buffer_12962 (.in(n12962), .out(n12962_0));
mux3 mux_7797 (.in({n12135_1, n12056_0, n2336}), .out(n12963), .config_in(config_chain[28489:28488]), .config_rst(config_rst)); 
buffer_wire buffer_12963 (.in(n12963), .out(n12963_0));
mux15 mux_7798 (.in({n12884_1, n11083_1, n11065_0, n11060_0, n11036_0, n10999_0, n10994_0, n10982_0, n10973_0, n10956_0/**/, n3022, n3014, n3006, n2038, n2030}), .out(n12964), .config_in(config_chain[28495:28490]), .config_rst(config_rst)); 
buffer_wire buffer_12964 (.in(n12964), .out(n12964_0));
mux3 mux_7799 (.in({n12137_1, n12064_0/**/, n3300}), .out(n12965), .config_in(config_chain[28497:28496]), .config_rst(config_rst)); 
buffer_wire buffer_12965 (.in(n12965), .out(n12965_0));
mux15 mux_7800 (.in({n12886_1, n11085_1, n11059_0, n11054_0, n11038_0, n11029_0, n11012_0/**/, n10986_0, n10975_0, n10958_0, n3022, n3014, n3006, n2038, n2030}), .out(n12966), .config_in(config_chain[28503:28498]), .config_rst(config_rst)); 
buffer_wire buffer_12966 (.in(n12966), .out(n12966_0));
mux3 mux_7801 (.in({n12139_1, n12072_0, n3304}), .out(n12967), .config_in(config_chain[28505:28504]), .config_rst(config_rst)); 
buffer_wire buffer_12967 (.in(n12967), .out(n12967_0));
mux15 mux_7802 (.in({n12888_1, n11087_1, n11053_0, n11048_0, n11040_0, n11031_0, n11014_0, n11005_0, n10988_0, n10978_0, n3022, n3014/**/, n3006, n2038, n2030}), .out(n12968), .config_in(config_chain[28511:28506]), .config_rst(config_rst)); 
buffer_wire buffer_12968 (.in(n12968), .out(n12968_0));
mux3 mux_7803 (.in({n12141_1/**/, n12080_0, n3308}), .out(n12969), .config_in(config_chain[28513:28512]), .config_rst(config_rst)); 
buffer_wire buffer_12969 (.in(n12969), .out(n12969_0));
mux15 mux_7804 (.in({n12890_1, n11069_1, n11067_0, n11062_0, n11042_0, n11007_0, n10990_0/**/, n10981_0, n10970_0, n10964_0, n3022, n3014, n3006, n2038, n2030}), .out(n12970), .config_in(config_chain[28519:28514]), .config_rst(config_rst)); 
buffer_wire buffer_12970 (.in(n12970), .out(n12970_0));
mux3 mux_7805 (.in({n12143_1, n12088_0, n3308}), .out(n12971), .config_in(config_chain[28521:28520]), .config_rst(config_rst)); 
buffer_wire buffer_12971 (.in(n12971), .out(n12971_0));
mux15 mux_7806 (.in({n12892_1, n11335_1, n11324_0, n11319_0, n11309_1, n11304_0, n11281_0, n11246_0, n11223_0/**/, n11220_0, n3116, n3108, n2140, n2132, n2124}), .out(n12972), .config_in(config_chain[28527:28522]), .config_rst(config_rst)); 
buffer_wire buffer_12972 (.in(n12972), .out(n12972_0));
mux4 mux_7807 (.in({n12011_0, n12010_0, n3316/**/, n2320}), .out(n12973), .config_in(config_chain[28529:28528]), .config_rst(config_rst)); 
buffer_wire buffer_12973 (.in(n12973), .out(n12973_0));
mux15 mux_7808 (.in({n12894_1, n11337_1, n11327_0, n11311_1/**/, n11306_0, n11300_0, n11278_0, n11255_0, n11248_0, n11225_0, n3120, n3108, n2140, n2132, n2124}), .out(n12974), .config_in(config_chain[28535:28530]), .config_rst(config_rst)); 
buffer_wire buffer_12974 (.in(n12974), .out(n12974_0));
mux3 mux_7809 (.in({n12019_0, n12018_0, n2320/**/}), .out(n12975), .config_in(config_chain[28537:28536]), .config_rst(config_rst)); 
buffer_wire buffer_12975 (.in(n12975), .out(n12975_0));
mux15 mux_7810 (.in({n12896_1, n11339_1, n11318_0, n11313_0/**/, n11308_0, n11292_0, n11287_0, n11280_0, n11257_0, n11222_0, n3120, n3112, n2140, n2132, n2124}), .out(n12976), .config_in(config_chain[28543:28538]), .config_rst(config_rst)); 
buffer_wire buffer_12976 (.in(n12976), .out(n12976_0));
mux3 mux_7811 (.in({n12027_0, n12026_0/**/, n2324}), .out(n12977), .config_in(config_chain[28545:28544]), .config_rst(config_rst)); 
buffer_wire buffer_12977 (.in(n12977), .out(n12977_0));
mux15 mux_7812 (.in({n12898_1, n11341_1, n11326_0, n11321_0, n11310_0, n11289_0, n11284_0, n11254_0, n11231_0/**/, n11224_0, n3120, n3112, n3104, n2132, n2124}), .out(n12978), .config_in(config_chain[28551:28546]), .config_rst(config_rst)); 
buffer_wire buffer_12978 (.in(n12978), .out(n12978_0));
mux3 mux_7813 (.in({n12035_0/**/, n12034_0, n2328}), .out(n12979), .config_in(config_chain[28553:28552]), .config_rst(config_rst)); 
buffer_wire buffer_12979 (.in(n12979), .out(n12979_0));
mux14 mux_7814 (.in({n12900_1, n11343_1, n11329_0/**/, n11312_0, n11286_0, n11276_0, n11263_0, n11256_0, n11233_0, n3120, n3112, n3104, n2136, n2124}), .out(n12980), .config_in(config_chain[28559:28554]), .config_rst(config_rst)); 
buffer_wire buffer_12980 (.in(n12980), .out(n12980_0));
mux3 mux_7815 (.in({n12043_0/**/, n12042_0, n2332}), .out(n12981), .config_in(config_chain[28561:28560]), .config_rst(config_rst)); 
buffer_wire buffer_12981 (.in(n12981), .out(n12981_0));
mux14 mux_7816 (.in({n12902_1, n11345_1, n11320_0, n11315_0, n11295_0, n11288_0, n11268_0, n11265_0, n11230_0, n3120, n3112/**/, n3104, n2136, n2128}), .out(n12982), .config_in(config_chain[28567:28562]), .config_rst(config_rst)); 
buffer_wire buffer_12982 (.in(n12982), .out(n12982_0));
mux3 mux_7817 (.in({n12051_0, n12050_0, n2336}), .out(n12983), .config_in(config_chain[28569:28568]), .config_rst(config_rst)); 
buffer_wire buffer_12983 (.in(n12983), .out(n12983_0));
mux13 mux_7818 (.in({n12904_1, n11347_1, n11328_0, n11323_0, n11297_0, n11262_0, n11260_0/**/, n11239_0, n11232_0, n3112, n3104, n2136, n2128}), .out(n12984), .config_in(config_chain[28575:28570]), .config_rst(config_rst)); 
buffer_wire buffer_12984 (.in(n12984), .out(n12984_0));
mux3 mux_7819 (.in({n12059_0, n12058_0, n2336}), .out(n12985), .config_in(config_chain[28577:28576]), .config_rst(config_rst)); 
buffer_wire buffer_12985 (.in(n12985), .out(n12985_0));
mux13 mux_7820 (.in({n12906_1, n11349_1, n11331_0, n11314_0, n11294_0, n11271_0, n11264_0, n11252_0/**/, n11241_0, n3116, n3104, n2136, n2128}), .out(n12986), .config_in(config_chain[28583:28578]), .config_rst(config_rst)); 
buffer_wire buffer_12986 (.in(n12986), .out(n12986_0));
mux3 mux_7821 (.in({n12067_0/**/, n12066_0, n3300}), .out(n12987), .config_in(config_chain[28585:28584]), .config_rst(config_rst)); 
buffer_wire buffer_12987 (.in(n12987), .out(n12987_0));
mux13 mux_7822 (.in({n12908_1, n11351_1, n11322_0, n11317_0, n11303_0, n11296_0, n11273_0, n11244_0/**/, n11238_0, n3116, n3108, n2136, n2128}), .out(n12988), .config_in(config_chain[28591:28586]), .config_rst(config_rst)); 
buffer_wire buffer_12988 (.in(n12988), .out(n12988_0));
mux3 mux_7823 (.in({n12075_0/**/, n12074_0, n3304}), .out(n12989), .config_in(config_chain[28593:28592]), .config_rst(config_rst)); 
buffer_wire buffer_12989 (.in(n12989), .out(n12989_0));
mux13 mux_7824 (.in({n12910_1, n11353_2, n11330_0, n11325_0, n11305_0/**/, n11270_0, n11247_0, n11240_0, n11236_0, n3116, n3108, n2140, n2128}), .out(n12990), .config_in(config_chain[28599:28594]), .config_rst(config_rst)); 
buffer_wire buffer_12990 (.in(n12990), .out(n12990_0));
mux3 mux_7825 (.in({n12083_0, n12082_0/**/, n3308}), .out(n12991), .config_in(config_chain[28601:28600]), .config_rst(config_rst)); 
buffer_wire buffer_12991 (.in(n12991), .out(n12991_0));
mux13 mux_7826 (.in({n12860_1, n11333_1, n11316_0, n11307_0, n11302_0, n11279_0, n11272_0, n11249_0, n11228_0, n3116, n3108, n2140, n2132}), .out(n12992), .config_in(config_chain[28607:28602]), .config_rst(config_rst)); 
buffer_wire buffer_12992 (.in(n12992), .out(n12992_0));
mux3 mux_7827 (.in({n12091_2, n12090_0, n3312}), .out(n12993), .config_in(config_chain[28609:28608]), .config_rst(config_rst)); 
buffer_wire buffer_12993 (.in(n12993), .out(n12993_0));
mux15 mux_7828 (.in({n12912_1, n11601_1, n11582_0, n11577_0, n11573_0, n11568_0, n11545_0, n11538_0, n11515_0, n11486_0, n3214, n3206/**/, n2238, n2230, n2222}), .out(n12994), .config_in(config_chain[28615:28610]), .config_rst(config_rst)); 
buffer_wire buffer_12994 (.in(n12994), .out(n12994_0));
mux4 mux_7829 (.in({n12013_0/**/, n12012_0, n3316, n2320}), .out(n12995), .config_in(config_chain[28617:28616]), .config_rst(config_rst)); 
buffer_wire buffer_12995 (.in(n12995), .out(n12995_0));
mux15 mux_7830 (.in({n12914_1, n11603_1, n11590_0, n11585_0, n11575_1, n11570_0, n11566_0, n11547_0, n11512_0, n11489_0, n3218, n3206, n2238, n2230, n2222/**/}), .out(n12996), .config_in(config_chain[28623:28618]), .config_rst(config_rst)); 
buffer_wire buffer_12996 (.in(n12996), .out(n12996_0));
mux3 mux_7831 (.in({n12021_0, n12020_0, n2324}), .out(n12997), .config_in(config_chain[28625:28624]), .config_rst(config_rst)); 
buffer_wire buffer_12997 (.in(n12997), .out(n12997_0));
mux15 mux_7832 (.in({n12916_1/**/, n11605_1, n11593_0, n11576_0, n11572_0, n11558_0, n11544_0, n11521_0, n11514_0, n11491_0, n3218, n3210, n2238, n2230, n2222}), .out(n12998), .config_in(config_chain[28631:28626]), .config_rst(config_rst)); 
buffer_wire buffer_12998 (.in(n12998), .out(n12998_0));
mux3 mux_7833 (.in({n12029_0, n12028_0, n2324}), .out(n12999), .config_in(config_chain[28633:28632]), .config_rst(config_rst)); 
buffer_wire buffer_12999 (.in(n12999), .out(n12999_0));
mux15 mux_7834 (.in({n12918_1, n11607_1, n11584_0, n11579_0/**/, n11574_0, n11553_0, n11550_0, n11546_0, n11523_0, n11488_0, n3218, n3210, n3202, n2230, n2222}), .out(n13000), .config_in(config_chain[28639:28634]), .config_rst(config_rst)); 
buffer_wire buffer_13000 (.in(n13000), .out(n13000_0));
mux3 mux_7835 (.in({n12037_0, n12036_0, n2328}), .out(n13001), .config_in(config_chain[28641:28640]), .config_rst(config_rst)); 
buffer_wire buffer_13001 (.in(n13001), .out(n13001_0));
mux14 mux_7836 (.in({n12920_1, n11609_1, n11592_0, n11587_0, n11555_0, n11542_0, n11520_0, n11497_0, n11490_0, n3218, n3210, n3202, n2234, n2222/**/}), .out(n13002), .config_in(config_chain[28647:28642]), .config_rst(config_rst)); 
buffer_wire buffer_13002 (.in(n13002), .out(n13002_0));
mux3 mux_7837 (.in({n12045_0, n12044_0, n2332}), .out(n13003), .config_in(config_chain[28649:28648]), .config_rst(config_rst)); 
buffer_wire buffer_13003 (.in(n13003), .out(n13003_0));
mux14 mux_7838 (.in({n12922_1/**/, n11611_1, n11595_0, n11578_0, n11552_0, n11534_0, n11529_0, n11522_0, n11499_0, n3218, n3210, n3202, n2234, n2226}), .out(n13004), .config_in(config_chain[28655:28650]), .config_rst(config_rst)); 
buffer_wire buffer_13004 (.in(n13004), .out(n13004_0));
mux3 mux_7839 (.in({n12053_0, n12052_0, n2336}), .out(n13005), .config_in(config_chain[28657:28656]), .config_rst(config_rst)); 
buffer_wire buffer_13005 (.in(n13005), .out(n13005_0));
mux13 mux_7840 (.in({n12924_1, n11613_1, n11586_0, n11581_0, n11561_0, n11554_0, n11531_0, n11526_0/**/, n11496_0, n3210, n3202, n2234, n2226}), .out(n13006), .config_in(config_chain[28663:28658]), .config_rst(config_rst)); 
buffer_wire buffer_13006 (.in(n13006), .out(n13006_0));
mux3 mux_7841 (.in({n12061_0, n12060_0, n3300}), .out(n13007), .config_in(config_chain[28665:28664]), .config_rst(config_rst)); 
buffer_wire buffer_13007 (.in(n13007), .out(n13007_0));
mux13 mux_7842 (.in({n12926_1, n11615_1, n11594_0, n11589_0, n11563_0, n11528_0, n11518_0/**/, n11505_0, n11498_0, n3214, n3202, n2234, n2226}), .out(n13008), .config_in(config_chain[28671:28666]), .config_rst(config_rst)); 
buffer_wire buffer_13008 (.in(n13008), .out(n13008_0));
mux3 mux_7843 (.in({n12069_0, n12068_0, n3300}), .out(n13009), .config_in(config_chain[28673:28672]), .config_rst(config_rst)); 
buffer_wire buffer_13009 (.in(n13009), .out(n13009_0));
mux13 mux_7844 (.in({n12928_1, n11617_1, n11597_2, n11580_0, n11560_0, n11537_0/**/, n11530_0, n11510_0, n11507_0, n3214, n3206, n2234, n2226}), .out(n13010), .config_in(config_chain[28679:28674]), .config_rst(config_rst)); 
buffer_wire buffer_13010 (.in(n13010), .out(n13010_0));
mux3 mux_7845 (.in({n12077_0, n12076_0, n3304}), .out(n13011), .config_in(config_chain[28681:28680]), .config_rst(config_rst)); 
buffer_wire buffer_13011 (.in(n13011), .out(n13011_0));
mux13 mux_7846 (.in({n12930_1/**/, n11619_2, n11588_0, n11583_0, n11569_0, n11562_0, n11539_0, n11504_0, n11502_0, n3214, n3206, n2238, n2226}), .out(n13012), .config_in(config_chain[28687:28682]), .config_rst(config_rst)); 
buffer_wire buffer_13012 (.in(n13012), .out(n13012_0));
mux3 mux_7847 (.in({n12085_0/**/, n12084_0, n3308}), .out(n13013), .config_in(config_chain[28689:28688]), .config_rst(config_rst)); 
buffer_wire buffer_13013 (.in(n13013), .out(n13013_0));
mux13 mux_7848 (.in({n12862_2, n11599_1, n11596_0, n11591_0, n11571_0, n11536_0, n11513_0, n11506_0, n11494_0, n3214, n3206, n2238/**/, n2230}), .out(n13014), .config_in(config_chain[28695:28690]), .config_rst(config_rst)); 
buffer_wire buffer_13014 (.in(n13014), .out(n13014_0));
mux3 mux_7849 (.in({n12093_2, n12092_0, n3312}), .out(n13015), .config_in(config_chain[28697:28696]), .config_rst(config_rst)); 
buffer_wire buffer_13015 (.in(n13015), .out(n13015_0));
mux15 mux_7850 (.in({n12932_1/**/, n11865_1, n11860_0, n11855_0, n11837_0, n11802_0, n11779_0, n11772_0, n11752_0, n11749_0, n3312, n3304, n2336, n2328, n2320}), .out(n13016), .config_in(config_chain[28703:28698]), .config_rst(config_rst)); 
buffer_wire buffer_13016 (.in(n13016), .out(n13016_0));
mux4 mux_7851 (.in({n12103_0, n12102_0, n3316, n2320}), .out(n13017), .config_in(config_chain[28705:28704]), .config_rst(config_rst)); 
buffer_wire buffer_13017 (.in(n13017), .out(n13017_0));
mux15 mux_7852 (.in({n12934_1, n11867_1, n11846_0, n11841_0, n11839_0, n11834_0, n11832_0, n11811_0, n11804_0, n11781_0, n3316, n3304, n2336, n2328, n2320}), .out(n13018), .config_in(config_chain[28711:28706]), .config_rst(config_rst)); 
buffer_wire buffer_13018 (.in(n13018), .out(n13018_0));
mux3 mux_7853 (.in({n12105_0, n12104_0, n2324}), .out(n13019), .config_in(config_chain[28713:28712]), .config_rst(config_rst)); 
buffer_wire buffer_13019 (.in(n13019), .out(n13019_0));
mux15 mux_7854 (.in({n12936_1, n11869_1, n11854_0, n11849_0, n11836_0, n11824_0, n11813_0, n11778_0, n11755_0, n11748_0/**/, n3316, n3308, n2336, n2328, n2320}), .out(n13020), .config_in(config_chain[28719:28714]), .config_rst(config_rst)); 
buffer_wire buffer_13020 (.in(n13020), .out(n13020_0));
mux3 mux_7855 (.in({n12107_0, n12106_0, n2328}), .out(n13021), .config_in(config_chain[28721:28720]), .config_rst(config_rst)); 
buffer_wire buffer_13021 (.in(n13021), .out(n13021_0));
mux15 mux_7856 (.in({n12938_1, n11871_1, n11857_0/**/, n11840_0, n11838_0, n11816_0, n11810_0, n11787_0, n11780_0, n11757_0, n3316, n3308, n3300, n2328, n2320}), .out(n13022), .config_in(config_chain[28727:28722]), .config_rst(config_rst)); 
buffer_wire buffer_13022 (.in(n13022), .out(n13022_0));
mux3 mux_7857 (.in({n12109_0, n12108_0, n2328}), .out(n13023), .config_in(config_chain[28729:28728]), .config_rst(config_rst)); 
buffer_wire buffer_13023 (.in(n13023), .out(n13023_0));
mux14 mux_7858 (.in({n12940_1, n11873_1, n11848_0, n11843_0, n11819_0, n11812_0/**/, n11808_0, n11789_0, n11754_0, n3316, n3308, n3300, n2332, n2320}), .out(n13024), .config_in(config_chain[28735:28730]), .config_rst(config_rst)); 
buffer_wire buffer_13024 (.in(n13024), .out(n13024_0));
mux3 mux_7859 (.in({n12111_0/**/, n12110_0, n2332}), .out(n13025), .config_in(config_chain[28737:28736]), .config_rst(config_rst)); 
buffer_wire buffer_13025 (.in(n13025), .out(n13025_0));
mux14 mux_7860 (.in({n12942_1/**/, n11875_1, n11856_0, n11851_0, n11821_0, n11800_0, n11786_0, n11763_0, n11756_0, n3316, n3308, n3300, n2332, n2324}), .out(n13026), .config_in(config_chain[28743:28738]), .config_rst(config_rst)); 
buffer_wire buffer_13026 (.in(n13026), .out(n13026_0));
mux3 mux_7861 (.in({n12113_0/**/, n12112_0, n2336}), .out(n13027), .config_in(config_chain[28745:28744]), .config_rst(config_rst)); 
buffer_wire buffer_13027 (.in(n13027), .out(n13027_0));
mux13 mux_7862 (.in({n12944_1, n11877_1, n11859_0, n11842_0, n11818_0, n11795_0, n11792_0, n11788_0, n11765_0, n3308, n3300, n2332, n2324}), .out(n13028), .config_in(config_chain[28751:28746]), .config_rst(config_rst)); 
buffer_wire buffer_13028 (.in(n13028), .out(n13028_0));
mux3 mux_7863 (.in({n12115_0, n12114_0, n3300}), .out(n13029), .config_in(config_chain[28753:28752]), .config_rst(config_rst)); 
buffer_wire buffer_13029 (.in(n13029), .out(n13029_0));
mux13 mux_7864 (.in({n12946_1, n11879_1, n11850_0/**/, n11845_0, n11827_0, n11820_0, n11797_0, n11784_0, n11762_0, n3312, n3300, n2332, n2324}), .out(n13030), .config_in(config_chain[28759:28754]), .config_rst(config_rst)); 
buffer_wire buffer_13030 (.in(n13030), .out(n13030_0));
mux3 mux_7865 (.in({n12117_0/**/, n12116_0, n3304}), .out(n13031), .config_in(config_chain[28761:28760]), .config_rst(config_rst)); 
buffer_wire buffer_13031 (.in(n13031), .out(n13031_0));
mux13 mux_7866 (.in({n12948_1, n11881_1, n11858_0, n11853_0, n11829_2, n11794_0, n11776_0, n11771_0, n11764_0, n3312, n3304, n2332, n2324}), .out(n13032), .config_in(config_chain[28767:28762]), .config_rst(config_rst)); 
buffer_wire buffer_13032 (.in(n13032), .out(n13032_0));
mux3 mux_7867 (.in({n12119_0/**/, n12118_0, n3304}), .out(n13033), .config_in(config_chain[28769:28768]), .config_rst(config_rst)); 
buffer_wire buffer_13033 (.in(n13033), .out(n13033_0));
mux13 mux_7868 (.in({n12950_1, n11883_2, n11861_2, n11844_0, n11826_0, n11803_0/**/, n11796_0, n11773_0, n11768_0, n3312, n3304, n2336, n2324}), .out(n13034), .config_in(config_chain[28775:28770]), .config_rst(config_rst)); 
buffer_wire buffer_13034 (.in(n13034), .out(n13034_0));
mux3 mux_7869 (.in({n12121_0/**/, n12120_0, n3308}), .out(n13035), .config_in(config_chain[28777:28776]), .config_rst(config_rst)); 
buffer_wire buffer_13035 (.in(n13035), .out(n13035_0));
mux13 mux_7870 (.in({n12864_2, n11863_1/**/, n11852_0, n11847_0, n11835_0, n11828_0, n11805_0, n11770_0, n11760_0, n3312, n3304, n2336, n2328}), .out(n13036), .config_in(config_chain[28783:28778]), .config_rst(config_rst)); 
buffer_wire buffer_13036 (.in(n13036), .out(n13036_0));
mux3 mux_7871 (.in({n12123_2, n12122_0, n3312}), .out(n13037), .config_in(config_chain[28785:28784]), .config_rst(config_rst)); 
buffer_wire buffer_13037 (.in(n13037), .out(n13037_0));
mux4 mux_7872 (.in({n9667_0, n9666_0, n3510, n2514}), .out(n13038), .config_in(config_chain[28787:28786]), .config_rst(config_rst)); 
buffer_wire buffer_13038 (.in(n13038), .out(n13038_0));
mux16 mux_7873 (.in({n13131_1, n10069_1/**/, n10044_0, n10041_0, n10018_0, n10015_0, n10009_1, n10000_0, n9987_0, n9928_0, n9922_0, n3506, n3498, n2530, n2522, n2514}), .out(n13039), .config_in(config_chain[28793:28788]), .config_rst(config_rst)); 
buffer_wire buffer_13039 (.in(n13039), .out(n13039_0));
mux4 mux_7874 (.in({n9759_0/**/, n9758_0, n3510, n2514}), .out(n13040), .config_in(config_chain[28795:28794]), .config_rst(config_rst)); 
buffer_wire buffer_13040 (.in(n13040), .out(n13040_0));
mux16 mux_7875 (.in({n13151_1, n10325_1, n10305_0, n10288_0, n10280_0, n10277_0, n10265_1, n10256_0, n10204_0, n10189_0, n10186_0, n3604, n3596, n2628, n2620, n2612}), .out(n13041), .config_in(config_chain[28801:28796]), .config_rst(config_rst)); 
buffer_wire buffer_13041 (.in(n13041), .out(n13041_0));
mux4 mux_7876 (.in({n9779_0, n9778_0, n3510, n2514}), .out(n13042), .config_in(config_chain[28803:28802]), .config_rst(config_rst)); 
buffer_wire buffer_13042 (.in(n13042), .out(n13042_0));
mux16 mux_7877 (.in({n13171_1, n10583_1, n10552_0, n10549_0, n10543_0, n10526_0, n10523_1, n10514_0, n10488_0, n10473_0, n10446_0/**/, n3702, n3694, n2726, n2718, n2710}), .out(n13043), .config_in(config_chain[28809:28804]), .config_rst(config_rst)); 
buffer_wire buffer_13043 (.in(n13043), .out(n13043_0));
mux4 mux_7878 (.in({n9799_1, n9672_0, n3510/**/, n2514}), .out(n13044), .config_in(config_chain[28811:28810]), .config_rst(config_rst)); 
buffer_wire buffer_13044 (.in(n13044), .out(n13044_0));
mux16 mux_7879 (.in({n13191_1, n10843_1, n10818_0/**/, n10815_0, n10792_0, n10789_0, n10783_1, n10774_0, n10759_0, n10708_0, n10694_0, n3800, n3792, n2824, n2816, n2808}), .out(n13045), .config_in(config_chain[28817:28812]), .config_rst(config_rst)); 
buffer_wire buffer_13045 (.in(n13045), .out(n13045_0));
mux3 mux_7880 (.in({n9675_0, n9674_0, n2514}), .out(n13046), .config_in(config_chain[28819:28818]), .config_rst(config_rst)); 
buffer_wire buffer_13046 (.in(n13046), .out(n13046_0));
mux16 mux_7881 (.in({n13133_1, n10067_1, n10038_0, n10035_0, n10029_0, n10012_0, n10011_1, n10002_0, n9978_0/**/, n9963_0, n9936_0, n3506, n3498, n2530, n2522, n2514}), .out(n13047), .config_in(config_chain[28825:28820]), .config_rst(config_rst)); 
buffer_wire buffer_13047 (.in(n13047), .out(n13047_0));
mux3 mux_7882 (.in({n9761_0/**/, n9760_0, n2518}), .out(n13048), .config_in(config_chain[28827:28826]), .config_rst(config_rst)); 
buffer_wire buffer_13048 (.in(n13048), .out(n13048_0));
mux16 mux_7883 (.in({n13153_1, n10323_1, n10302_0, n10299_0, n10274_0, n10271_0, n10267_1, n10258_0, n10245_0, n10194_0, n10180_0, n3604, n3596, n2628/**/, n2620, n2612}), .out(n13049), .config_in(config_chain[28833:28828]), .config_rst(config_rst)); 
buffer_wire buffer_13049 (.in(n13049), .out(n13049_0));
mux3 mux_7884 (.in({n9781_0, n9780_0, n2518}), .out(n13050), .config_in(config_chain[28835:28834]), .config_rst(config_rst)); 
buffer_wire buffer_13050 (.in(n13050), .out(n13050_0));
mux16 mux_7885 (.in({n13173_1, n10581_1, n10563_0, n10546_0, n10540_0, n10537_0, n10525_1, n10516_0, n10464_0, n10454_0, n10449_0, n3702, n3694/**/, n2726, n2718, n2710}), .out(n13051), .config_in(config_chain[28841:28836]), .config_rst(config_rst)); 
buffer_wire buffer_13051 (.in(n13051), .out(n13051_0));
mux3 mux_7886 (.in({n9801_1/**/, n9680_0, n2518}), .out(n13052), .config_in(config_chain[28843:28842]), .config_rst(config_rst)); 
buffer_wire buffer_13052 (.in(n13052), .out(n13052_0));
mux16 mux_7887 (.in({n13193_1, n10841_1, n10812_0, n10809_0, n10803_0/**/, n10786_0, n10785_1, n10776_0, n10750_0, n10735_0, n10716_0, n3800, n3792, n2824, n2816, n2808}), .out(n13053), .config_in(config_chain[28849:28844]), .config_rst(config_rst)); 
buffer_wire buffer_13053 (.in(n13053), .out(n13053_0));
mux3 mux_7888 (.in({n9683_0, n9682_0/**/, n2518}), .out(n13054), .config_in(config_chain[28851:28850]), .config_rst(config_rst)); 
buffer_wire buffer_13054 (.in(n13054), .out(n13054_0));
mux15 mux_7889 (.in({n13135_1, n10065_1, n10049_0, n10032_0, n10026_0, n10023_0, n10004_0, n9954_0, n9944_0, n9939_0, n3506, n3498, n2530, n2522, n2514}), .out(n13055), .config_in(config_chain[28857:28852]), .config_rst(config_rst)); 
buffer_wire buffer_13055 (.in(n13055), .out(n13055_0));
mux3 mux_7890 (.in({n9763_0/**/, n9762_0, n2518}), .out(n13056), .config_in(config_chain[28859:28858]), .config_rst(config_rst)); 
buffer_wire buffer_13056 (.in(n13056), .out(n13056_0));
mux15 mux_7891 (.in({n13155_1/**/, n10321_1, n10296_0, n10293_0, n10285_0, n10268_0, n10260_0, n10236_0, n10221_0, n10202_0, n3604, n3596, n2628, n2620, n2612}), .out(n13057), .config_in(config_chain[28865:28860]), .config_rst(config_rst)); 
buffer_wire buffer_13057 (.in(n13057), .out(n13057_0));
mux3 mux_7892 (.in({n9783_0/**/, n9782_0, n2522}), .out(n13058), .config_in(config_chain[28867:28866]), .config_rst(config_rst)); 
buffer_wire buffer_13058 (.in(n13058), .out(n13058_0));
mux15 mux_7893 (.in({n13175_1, n10579_1, n10560_0, n10557_0, n10534_0, n10531_0, n10518_0, n10505_0, n10462_0/**/, n10440_0, n3702, n3694, n2726, n2718, n2710}), .out(n13059), .config_in(config_chain[28873:28868]), .config_rst(config_rst)); 
buffer_wire buffer_13059 (.in(n13059), .out(n13059_0));
mux3 mux_7894 (.in({n9803_1/**/, n9688_0, n2522}), .out(n13060), .config_in(config_chain[28875:28874]), .config_rst(config_rst)); 
buffer_wire buffer_13060 (.in(n13060), .out(n13060_0));
mux15 mux_7895 (.in({n13195_1/**/, n10839_1, n10823_0, n10806_0, n10800_0, n10797_0, n10778_0, n10726_0, n10724_0, n10711_0, n3800, n3792, n2824, n2816, n2808}), .out(n13061), .config_in(config_chain[28881:28876]), .config_rst(config_rst)); 
buffer_wire buffer_13061 (.in(n13061), .out(n13061_0));
mux3 mux_7896 (.in({n9691_0, n9690_0, n2522}), .out(n13062), .config_in(config_chain[28883:28882]), .config_rst(config_rst)); 
buffer_wire buffer_13062 (.in(n13062), .out(n13062_0));
mux15 mux_7897 (.in({n13137_1, n10063_1/**/, n10046_0, n10043_0, n10020_0, n10017_0, n10006_0, n9995_0, n9952_0, n9930_0, n3506, n3498, n2530, n2522, n2514}), .out(n13063), .config_in(config_chain[28889:28884]), .config_rst(config_rst)); 
buffer_wire buffer_13063 (.in(n13063), .out(n13063_0));
mux3 mux_7898 (.in({n9765_0, n9764_0, n2522}), .out(n13064), .config_in(config_chain[28891:28890]), .config_rst(config_rst)); 
buffer_wire buffer_13064 (.in(n13064), .out(n13064_0));
mux15 mux_7899 (.in({n13157_1, n10319_1, n10307_0, n10290_0/**/, n10282_0, n10279_0, n10262_0, n10212_0, n10210_0, n10197_0, n3604, n3596, n2628, n2620, n2612}), .out(n13065), .config_in(config_chain[28897:28892]), .config_rst(config_rst)); 
buffer_wire buffer_13065 (.in(n13065), .out(n13065_0));
mux3 mux_7900 (.in({n9785_0, n9784_0/**/, n2522}), .out(n13066), .config_in(config_chain[28899:28898]), .config_rst(config_rst)); 
buffer_wire buffer_13066 (.in(n13066), .out(n13066_0));
mux15 mux_7901 (.in({n13177_1, n10577_1, n10554_0, n10551_0, n10545_0, n10528_0, n10520_0, n10496_0, n10481_0, n10470_0, n3702, n3694, n2726, n2718, n2710}), .out(n13067), .config_in(config_chain[28905:28900]), .config_rst(config_rst)); 
buffer_wire buffer_13067 (.in(n13067), .out(n13067_0));
mux3 mux_7902 (.in({n9805_1, n9696_0, n2526}), .out(n13068), .config_in(config_chain[28907:28906]), .config_rst(config_rst)); 
buffer_wire buffer_13068 (.in(n13068), .out(n13068_0));
mux15 mux_7903 (.in({n13197_1, n10837_1, n10820_0, n10817_0, n10794_0, n10791_0, n10780_0, n10767_0, n10732_0, n10702_0, n3800, n3792/**/, n2824, n2816, n2808}), .out(n13069), .config_in(config_chain[28913:28908]), .config_rst(config_rst)); 
buffer_wire buffer_13069 (.in(n13069), .out(n13069_0));
mux3 mux_7904 (.in({n9699_0, n9698_0, n2526}), .out(n13070), .config_in(config_chain[28915:28914]), .config_rst(config_rst)); 
buffer_wire buffer_13070 (.in(n13070), .out(n13070_0));
mux15 mux_7905 (.in({n13139_1, n10061_1, n10040_0, n10037_0, n10031_0, n10014_0, n10008_0, n9986_0, n9971_0, n9960_0, n3506, n3498, n2530, n2522, n2514}), .out(n13071), .config_in(config_chain[28921:28916]), .config_rst(config_rst)); 
buffer_wire buffer_13071 (.in(n13071), .out(n13071_0));
mux3 mux_7906 (.in({n9767_0/**/, n9766_0, n2526}), .out(n13072), .config_in(config_chain[28923:28922]), .config_rst(config_rst)); 
buffer_wire buffer_13072 (.in(n13072), .out(n13072_0));
mux15 mux_7907 (.in({n13159_1, n10317_1, n10304_0, n10301_0, n10276_0, n10273_0, n10264_0, n10253_0, n10218_0, n10188_0, n3604, n3596, n2628, n2620, n2612}), .out(n13073), .config_in(config_chain[28929:28924]), .config_rst(config_rst)); 
buffer_wire buffer_13073 (.in(n13073), .out(n13073_0));
mux3 mux_7908 (.in({n9787_0, n9786_0/**/, n2526}), .out(n13074), .config_in(config_chain[28931:28930]), .config_rst(config_rst)); 
buffer_wire buffer_13074 (.in(n13074), .out(n13074_0));
mux15 mux_7909 (.in({n13179_1, n10575_1, n10565_0, n10548_0, n10542_0, n10539_0, n10522_0, n10478_0, n10472_0, n10457_0, n3702, n3694, n2726/**/, n2718, n2710}), .out(n13075), .config_in(config_chain[28937:28932]), .config_rst(config_rst)); 
buffer_wire buffer_13075 (.in(n13075), .out(n13075_0));
mux3 mux_7910 (.in({n9807_1, n9704_0, n2526}), .out(n13076), .config_in(config_chain[28939:28938]), .config_rst(config_rst)); 
buffer_wire buffer_13076 (.in(n13076), .out(n13076_0));
mux15 mux_7911 (.in({n13199_1, n10835_1, n10814_0, n10811_0, n10805_0, n10788_0, n10782_0, n10758_0, n10743_0, n10740_0, n3800, n3792/**/, n2824, n2816, n2808}), .out(n13077), .config_in(config_chain[28945:28940]), .config_rst(config_rst)); 
buffer_wire buffer_13077 (.in(n13077), .out(n13077_0));
mux3 mux_7912 (.in({n9707_0/**/, n9706_0, n2530}), .out(n13078), .config_in(config_chain[28947:28946]), .config_rst(config_rst)); 
buffer_wire buffer_13078 (.in(n13078), .out(n13078_0));
mux15 mux_7913 (.in({n13141_1, n10059_1, n10051_0/**/, n10034_0, n10028_0, n10025_0, n10010_0, n9968_0, n9962_0, n9947_0, n3510, n3502, n3494, n2526, n2518}), .out(n13079), .config_in(config_chain[28953:28948]), .config_rst(config_rst)); 
buffer_wire buffer_13079 (.in(n13079), .out(n13079_0));
mux3 mux_7914 (.in({n9769_0/**/, n9768_0, n2530}), .out(n13080), .config_in(config_chain[28955:28954]), .config_rst(config_rst)); 
buffer_wire buffer_13080 (.in(n13080), .out(n13080_0));
mux15 mux_7915 (.in({n13161_1, n10315_1, n10298_0, n10295_0, n10287_0, n10270_0, n10266_0, n10244_0, n10229_0, n10226_0, n3608, n3600/**/, n3592, n2624, n2616}), .out(n13081), .config_in(config_chain[28961:28956]), .config_rst(config_rst)); 
buffer_wire buffer_13081 (.in(n13081), .out(n13081_0));
mux3 mux_7916 (.in({n9789_0/**/, n9788_0, n2530}), .out(n13082), .config_in(config_chain[28963:28962]), .config_rst(config_rst)); 
buffer_wire buffer_13082 (.in(n13082), .out(n13082_0));
mux15 mux_7917 (.in({n13181_1, n10573_1/**/, n10562_0, n10559_0, n10536_0, n10533_0, n10524_0, n10513_0, n10486_0, n10448_0, n3706, n3698, n3690, n2722, n2714}), .out(n13083), .config_in(config_chain[28969:28964]), .config_rst(config_rst)); 
buffer_wire buffer_13083 (.in(n13083), .out(n13083_0));
mux3 mux_7918 (.in({n9809_1, n9712_0, n2530/**/}), .out(n13084), .config_in(config_chain[28971:28970]), .config_rst(config_rst)); 
buffer_wire buffer_13084 (.in(n13084), .out(n13084_0));
mux15 mux_7919 (.in({n13201_1, n10833_1, n10825_0, n10808_0, n10802_0, n10799_0, n10784_0, n10748_0, n10734_0, n10719_0, n3804, n3796, n3788, n2820/**/, n2812}), .out(n13085), .config_in(config_chain[28977:28972]), .config_rst(config_rst)); 
buffer_wire buffer_13085 (.in(n13085), .out(n13085_0));
mux3 mux_7920 (.in({n9715_0, n9714_0, n2530}), .out(n13086), .config_in(config_chain[28979:28978]), .config_rst(config_rst)); 
buffer_wire buffer_13086 (.in(n13086), .out(n13086_0));
mux15 mux_7921 (.in({n13143_1, n10057_1, n10048_0, n10045_0, n10022_0, n10019_0, n10001_1, n9976_0, n9938_0/**/, n9923_0, n3510, n3502, n3494, n2526, n2518}), .out(n13087), .config_in(config_chain[28985:28980]), .config_rst(config_rst)); 
buffer_wire buffer_13087 (.in(n13087), .out(n13087_0));
mux3 mux_7922 (.in({n9771_0/**/, n9770_0, n3494}), .out(n13088), .config_in(config_chain[28987:28986]), .config_rst(config_rst)); 
buffer_wire buffer_13088 (.in(n13088), .out(n13088_0));
mux15 mux_7923 (.in({n13163_1, n10313_1, n10292_0, n10289_0, n10284_0, n10281_0, n10257_0, n10234_0, n10220_0, n10205_0, n3608/**/, n3600, n3592, n2624, n2616}), .out(n13089), .config_in(config_chain[28993:28988]), .config_rst(config_rst)); 
buffer_wire buffer_13089 (.in(n13089), .out(n13089_0));
mux3 mux_7924 (.in({n9791_0, n9790_0, n3494/**/}), .out(n13090), .config_in(config_chain[28995:28994]), .config_rst(config_rst)); 
buffer_wire buffer_13090 (.in(n13090), .out(n13090_0));
mux15 mux_7925 (.in({n13183_1, n10571_1, n10556_0, n10553_0, n10530_0, n10527_0, n10515_0, n10504_0, n10494_0, n10489_0, n3706/**/, n3698, n3690, n2722, n2714}), .out(n13091), .config_in(config_chain[29001:28996]), .config_rst(config_rst)); 
buffer_wire buffer_13091 (.in(n13091), .out(n13091_0));
mux3 mux_7926 (.in({n9811_1, n9720_0, n3494/**/}), .out(n13092), .config_in(config_chain[29003:29002]), .config_rst(config_rst)); 
buffer_wire buffer_13092 (.in(n13092), .out(n13092_0));
mux15 mux_7927 (.in({n13203_1, n10831_1, n10822_0, n10819_0, n10796_0, n10793_0, n10775_0, n10756_0, n10710_0, n10695_0, n3804/**/, n3796, n3788, n2820, n2812}), .out(n13093), .config_in(config_chain[29009:29004]), .config_rst(config_rst)); 
buffer_wire buffer_13093 (.in(n13093), .out(n13093_0));
mux3 mux_7928 (.in({n9723_0, n9722_0, n3494}), .out(n13094), .config_in(config_chain[29011:29010]), .config_rst(config_rst)); 
buffer_wire buffer_13094 (.in(n13094), .out(n13094_0));
mux15 mux_7929 (.in({n13145_1, n10055_1, n10042_0, n10039_0, n10016_0, n10013_0, n10003_1, n9994_0, n9984_0/**/, n9979_0, n3510, n3502, n3494, n2526, n2518}), .out(n13095), .config_in(config_chain[29017:29012]), .config_rst(config_rst)); 
buffer_wire buffer_13095 (.in(n13095), .out(n13095_0));
mux3 mux_7930 (.in({n9773_0/**/, n9772_0, n3494}), .out(n13096), .config_in(config_chain[29019:29018]), .config_rst(config_rst)); 
buffer_wire buffer_13096 (.in(n13096), .out(n13096_0));
mux15 mux_7931 (.in({n13165_1, n10311_1, n10306_0, n10303_0, n10278_0, n10275_0, n10259_1, n10242_0/**/, n10196_0, n10181_0, n3608, n3600, n3592, n2624, n2616}), .out(n13097), .config_in(config_chain[29025:29020]), .config_rst(config_rst)); 
buffer_wire buffer_13097 (.in(n13097), .out(n13097_0));
mux3 mux_7932 (.in({n9793_0, n9792_0, n3498/**/}), .out(n13098), .config_in(config_chain[29027:29026]), .config_rst(config_rst)); 
buffer_wire buffer_13098 (.in(n13098), .out(n13098_0));
mux15 mux_7933 (.in({n13185_1, n10569_1, n10550_0, n10547_0, n10544_0/**/, n10541_0, n10517_0, n10502_0, n10480_0, n10465_0, n3706, n3698, n3690, n2722, n2714}), .out(n13099), .config_in(config_chain[29033:29028]), .config_rst(config_rst)); 
buffer_wire buffer_13099 (.in(n13099), .out(n13099_0));
mux3 mux_7934 (.in({n9813_1, n9728_0, n3498}), .out(n13100), .config_in(config_chain[29035:29034]), .config_rst(config_rst)); 
buffer_wire buffer_13100 (.in(n13100), .out(n13100_0));
mux15 mux_7935 (.in({n13205_1, n10829_1, n10816_0, n10813_0, n10790_0, n10787_0, n10777_0, n10766_0, n10764_0/**/, n10751_0, n3804, n3796, n3788, n2820, n2812}), .out(n13101), .config_in(config_chain[29041:29036]), .config_rst(config_rst)); 
buffer_wire buffer_13101 (.in(n13101), .out(n13101_0));
mux3 mux_7936 (.in({n9731_0, n9730_0, n3498}), .out(n13102), .config_in(config_chain[29043:29042]), .config_rst(config_rst)); 
buffer_wire buffer_13102 (.in(n13102), .out(n13102_0));
mux15 mux_7937 (.in({n13147_1, n10053_1, n10036_0, n10033_0, n10030_0, n10027_0, n10005_1, n9992_0/**/, n9970_0, n9955_0, n3510, n3502, n3494, n2526, n2518}), .out(n13103), .config_in(config_chain[29049:29044]), .config_rst(config_rst)); 
buffer_wire buffer_13103 (.in(n13103), .out(n13103_0));
mux3 mux_7938 (.in({n9775_0/**/, n9774_0, n3498}), .out(n13104), .config_in(config_chain[29051:29050]), .config_rst(config_rst)); 
buffer_wire buffer_13104 (.in(n13104), .out(n13104_0));
mux15 mux_7939 (.in({n13167_1, n10309_1, n10300_0, n10297_0, n10272_0, n10269_0, n10261_1, n10252_0, n10250_0, n10237_0, n3608, n3600, n3592/**/, n2624, n2616}), .out(n13105), .config_in(config_chain[29057:29052]), .config_rst(config_rst)); 
buffer_wire buffer_13105 (.in(n13105), .out(n13105_0));
mux3 mux_7940 (.in({n9795_0, n9794_0, n3498}), .out(n13106), .config_in(config_chain[29059:29058]), .config_rst(config_rst)); 
buffer_wire buffer_13106 (.in(n13106), .out(n13106_0));
mux15 mux_7941 (.in({n13187_1, n10567_1, n10564_0, n10561_0, n10538_0, n10535_0, n10519_1, n10510_0, n10456_0, n10441_0, n3706, n3698, n3690, n2722, n2714/**/}), .out(n13107), .config_in(config_chain[29065:29060]), .config_rst(config_rst)); 
buffer_wire buffer_13107 (.in(n13107), .out(n13107_0));
mux3 mux_7942 (.in({n9815_1, n9736_0, n3502}), .out(n13108), .config_in(config_chain[29067:29066]), .config_rst(config_rst)); 
buffer_wire buffer_13108 (.in(n13108), .out(n13108_0));
mux15 mux_7943 (.in({n13207_1, n10827_1/**/, n10810_0, n10807_0, n10804_0, n10801_0, n10779_0, n10772_0, n10742_0, n10727_0, n3804, n3796, n3788, n2820, n2812}), .out(n13109), .config_in(config_chain[29073:29068]), .config_rst(config_rst)); 
buffer_wire buffer_13109 (.in(n13109), .out(n13109_0));
mux3 mux_7944 (.in({n9739_0, n9738_0, n3502}), .out(n13110), .config_in(config_chain[29075:29074]), .config_rst(config_rst)); 
buffer_wire buffer_13110 (.in(n13110), .out(n13110_0));
mux15 mux_7945 (.in({n13149_1, n10071_1, n10050_0, n10047_0, n10024_0, n10021_0, n10007_1, n9946_0, n9931_0, n9920_0, n3510, n3502, n3494, n2526, n2518}), .out(n13111), .config_in(config_chain[29081:29076]), .config_rst(config_rst)); 
buffer_wire buffer_13111 (.in(n13111), .out(n13111_0));
mux3 mux_7946 (.in({n9777_0/**/, n9776_0, n3502}), .out(n13112), .config_in(config_chain[29083:29082]), .config_rst(config_rst)); 
buffer_wire buffer_13112 (.in(n13112), .out(n13112_0));
mux15 mux_7947 (.in({n13169_1, n10327_1, n10294_0, n10291_0, n10286_0, n10283_0, n10263_1, n10228_0/**/, n10213_0, n10178_0, n3608, n3600, n3592, n2624, n2616}), .out(n13113), .config_in(config_chain[29089:29084]), .config_rst(config_rst)); 
buffer_wire buffer_13113 (.in(n13113), .out(n13113_0));
mux3 mux_7948 (.in({n9797_0/**/, n9796_0, n3502}), .out(n13114), .config_in(config_chain[29091:29090]), .config_rst(config_rst)); 
buffer_wire buffer_13114 (.in(n13114), .out(n13114_0));
mux15 mux_7949 (.in({n13189_1, n10585_1, n10558_0, n10555_0, n10532_0, n10529_0, n10521_1, n10512_0, n10497_0, n10438_0/**/, n3706, n3698, n3690, n2722, n2714}), .out(n13115), .config_in(config_chain[29097:29092]), .config_rst(config_rst)); 
buffer_wire buffer_13115 (.in(n13115), .out(n13115_0));
mux3 mux_7950 (.in({n9817_1, n9744_0, n3502}), .out(n13116), .config_in(config_chain[29099:29098]), .config_rst(config_rst)); 
buffer_wire buffer_13116 (.in(n13116), .out(n13116_0));
mux15 mux_7951 (.in({n13209_1/**/, n10845_1, n10824_0, n10821_0, n10798_0, n10795_0, n10781_1, n10718_0, n10703_0, n10700_0, n3804, n3796, n3788, n2820, n2812}), .out(n13117), .config_in(config_chain[29105:29100]), .config_rst(config_rst)); 
buffer_wire buffer_13117 (.in(n13117), .out(n13117_0));
mux3 mux_7952 (.in({n9747_1, n9746_0, n3506}), .out(n13118), .config_in(config_chain[29107:29106]), .config_rst(config_rst)); 
buffer_wire buffer_13118 (.in(n13118), .out(n13118_0));
mux13 mux_7953 (.in({n13231_1, n11109_1, n11073_0, n11061_0, n11054_0, n11042_0, n11039_0/**/, n11014_0, n10956_0, n3898, n3890, n2922, n2914}), .out(n13119), .config_in(config_chain[29113:29108]), .config_rst(config_rst)); 
buffer_wire buffer_13119 (.in(n13119), .out(n13119_0));
mux3 mux_7954 (.in({n9749_1, n9748_0, n3506}), .out(n13120), .config_in(config_chain[29115:29114]), .config_rst(config_rst)); 
buffer_wire buffer_13120 (.in(n13120), .out(n13120_0));
mux13 mux_7955 (.in({n13253_0, n11375_1, n11353_1, n11346_0, n11317_0, n11306_0, n11273_0/**/, n11248_0, n11222_0, n3996, n3988, n3020, n3012}), .out(n13121), .config_in(config_chain[29121:29116]), .config_rst(config_rst)); 
buffer_wire buffer_13121 (.in(n13121), .out(n13121_0));
mux3 mux_7956 (.in({n9751_1, n9750_0, n3506}), .out(n13122), .config_in(config_chain[29123:29122]), .config_rst(config_rst)); 
buffer_wire buffer_13122 (.in(n13122), .out(n13122_0));
mux13 mux_7957 (.in({n13275_0, n11641_1, n11611_0, n11604_0, n11597_1, n11590_0, n11570_0, n11507_0, n11488_0, n4094, n4086, n3118, n3110}), .out(n13123), .config_in(config_chain[29129:29124]), .config_rst(config_rst)); 
buffer_wire buffer_13123 (.in(n13123), .out(n13123_0));
mux3 mux_7958 (.in({n9753_1, n9752_0, n3506}), .out(n13124), .config_in(config_chain[29131:29130]), .config_rst(config_rst)); 
buffer_wire buffer_13124 (.in(n13124), .out(n13124_0));
mux13 mux_7959 (.in({n13297_0, n11905_1, n11882_0, n11867_0, n11853_0, n11846_0, n11829_1, n11804_0, n11754_0, n4192, n4184, n3216, n3208}), .out(n13125), .config_in(config_chain[29137:29132]), .config_rst(config_rst)); 
buffer_wire buffer_13125 (.in(n13125), .out(n13125_0));
mux3 mux_7960 (.in({n9755_1, n9754_0, n3506}), .out(n13126), .config_in(config_chain[29139:29138]), .config_rst(config_rst)); 
buffer_wire buffer_13126 (.in(n13126), .out(n13126_0));
mux3 mux_7961 (.in({n12167_1/**/, n12098_0, n4290}), .out(n13127), .config_in(config_chain[29141:29140]), .config_rst(config_rst)); 
buffer_wire buffer_13127 (.in(n13127), .out(n13127_0));
mux3 mux_7962 (.in({n9757_1, n9756_0, n3510}), .out(n13128), .config_in(config_chain[29143:29142]), .config_rst(config_rst)); 
buffer_wire buffer_13128 (.in(n13128), .out(n13128_0));
mux3 mux_7963 (.in({n12101_0, n12100_0, n4294}), .out(n13129), .config_in(config_chain[29145:29144]), .config_rst(config_rst)); 
buffer_wire buffer_13129 (.in(n13129), .out(n13129_0));
mux16 mux_7964 (.in({n13038_0, n10055_1/**/, n10045_0, n10040_0, n10019_0, n10014_0, n10008_0, n10001_1, n9986_0, n9923_0, n9920_0, n3604, n3596, n2628, n2620, n2612}), .out(n13130), .config_in(config_chain[29151:29146]), .config_rst(config_rst)); 
buffer_wire buffer_13130 (.in(n13130), .out(n13130_0));
mux15 mux_7965 (.in({n13211_1, n11107_1, n11081_0, n11074_0, n11062_0, n11044_0, n11041_0, n10983_0, n10964_0, n10958_0/**/, n3898, n3890, n2922, n2914, n2906}), .out(n13131), .config_in(config_chain[29157:29152]), .config_rst(config_rst)); 
buffer_wire buffer_13131 (.in(n13131), .out(n13131_0));
mux16 mux_7966 (.in({n13046_0, n10057_1, n10039_0/**/, n10034_0, n10028_0, n10013_0, n10010_0, n10003_1, n9992_0, n9979_0, n9962_0, n3604, n3596, n2628, n2620, n2612}), .out(n13132), .config_in(config_chain[29163:29158]), .config_rst(config_rst)); 
buffer_wire buffer_13132 (.in(n13132), .out(n13132_0));
mux15 mux_7967 (.in({n13213_1, n11105_1, n11082_0, n11055_0, n11048_0, n11046_0, n11043_0, n11015_0/**/, n10990_0, n10972_0, n3902, n3890, n2922, n2914, n2906}), .out(n13133), .config_in(config_chain[29169:29164]), .config_rst(config_rst)); 
buffer_wire buffer_13133 (.in(n13133), .out(n13133_0));
mux15 mux_7968 (.in({n13054_0, n10059_1, n10048_0/**/, n10033_0, n10027_0, n10022_0, n10005_1, n9984_0, n9955_0, n9938_0, n3604, n3596, n2628, n2620, n2612}), .out(n13134), .config_in(config_chain[29175:29170]), .config_rst(config_rst)); 
buffer_wire buffer_13134 (.in(n13134), .out(n13134_0));
mux15 mux_7969 (.in({n13215_1, n11103_1, n11075_0, n11068_0, n11063_0, n11056_0, n11045_1, n11022_0, n10980_0/**/, n10959_0, n3902, n3894, n2922, n2914, n2906}), .out(n13135), .config_in(config_chain[29181:29176]), .config_rst(config_rst)); 
buffer_wire buffer_13135 (.in(n13135), .out(n13135_0));
mux15 mux_7970 (.in({n13062_0, n10061_1, n10047_0, n10042_0, n10021_0, n10016_0, n10007_1, n9994_0/**/, n9976_0, n9931_0, n3604, n3596, n2628, n2620, n2612}), .out(n13136), .config_in(config_chain[29187:29182]), .config_rst(config_rst)); 
buffer_wire buffer_13136 (.in(n13136), .out(n13136_0));
mux15 mux_7971 (.in({n13217_1, n11101_1, n11083_0, n11076_0, n11064_0, n11049_0, n11047_1, n10991_0, n10988_0, n10966_0, n3902, n3894/**/, n3886, n2914, n2906}), .out(n13137), .config_in(config_chain[29193:29188]), .config_rst(config_rst)); 
buffer_wire buffer_13137 (.in(n13137), .out(n13137_0));
mux15 mux_7972 (.in({n13070_0, n10063_1, n10041_0, n10036_0, n10030_0, n10015_0, n10009_1, n9987_0, n9970_0/**/, n9968_0, n3604, n3596, n2628, n2620, n2612}), .out(n13138), .config_in(config_chain[29199:29194]), .config_rst(config_rst)); 
buffer_wire buffer_13138 (.in(n13138), .out(n13138_0));
mux14 mux_7973 (.in({n13219_1, n11099_1, n11084_0, n11069_0, n11057_0, n11050_0, n11023_0, n10998_0, n10996_0, n3902, n3894, n3886, n2918/**/, n2906}), .out(n13139), .config_in(config_chain[29205:29200]), .config_rst(config_rst)); 
buffer_wire buffer_13139 (.in(n13139), .out(n13139_0));
mux15 mux_7974 (.in({n13078_0/**/, n10065_1, n10050_0, n10035_0, n10029_0, n10024_0, n10011_1, n9963_0, n9960_0, n9946_0, n3608, n3600, n3592, n2624, n2616}), .out(n13140), .config_in(config_chain[29211:29206]), .config_rst(config_rst)); 
buffer_wire buffer_13140 (.in(n13140), .out(n13140_0));
mux14 mux_7975 (.in({n13221_1, n11097_1, n11077_0/**/, n11070_0, n11065_0, n11058_0, n11030_0, n11004_0, n10967_0, n3902, n3894, n3886, n2918, n2910}), .out(n13141), .config_in(config_chain[29217:29212]), .config_rst(config_rst)); 
buffer_wire buffer_13141 (.in(n13141), .out(n13141_0));
mux15 mux_7976 (.in({n13086_0, n10067_1, n10049_0, n10044_0, n10023_0, n10018_0, n10000_0, n9952_0, n9939_0, n9922_0/**/, n3608, n3600, n3592, n2624, n2616}), .out(n13142), .config_in(config_chain[29223:29218]), .config_rst(config_rst)); 
buffer_wire buffer_13142 (.in(n13142), .out(n13142_0));
mux13 mux_7977 (.in({n13223_1, n11095_1, n11085_0, n11078_0, n11066_0, n11051_0, n11012_0, n10999_0, n10974_0, n3894, n3886, n2918, n2910}), .out(n13143), .config_in(config_chain[29229:29224]), .config_rst(config_rst)); 
buffer_wire buffer_13143 (.in(n13143), .out(n13143_0));
mux15 mux_7978 (.in({n13094_0, n10069_1, n10043_0, n10038_0, n10017_0, n10012_0, n10002_0, n9995_0, n9978_0, n9944_0, n3608, n3600/**/, n3592, n2624, n2616}), .out(n13144), .config_in(config_chain[29235:29230]), .config_rst(config_rst)); 
buffer_wire buffer_13144 (.in(n13144), .out(n13144_0));
mux13 mux_7979 (.in({n13225_1, n11093_1, n11086_0, n11071_0, n11059_0, n11052_0, n11031_0, n11020_0, n11006_0, n3898, n3886, n2918/**/, n2910}), .out(n13145), .config_in(config_chain[29241:29236]), .config_rst(config_rst)); 
buffer_wire buffer_13145 (.in(n13145), .out(n13145_0));
mux15 mux_7980 (.in({n13102_0, n10071_1, n10037_0, n10032_0, n10031_0, n10026_0, n10004_0, n9971_0, n9954_0, n9936_0, n3608, n3600/**/, n3592, n2624, n2616}), .out(n13146), .config_in(config_chain[29247:29242]), .config_rst(config_rst)); 
buffer_wire buffer_13146 (.in(n13146), .out(n13146_0));
mux13 mux_7981 (.in({n13227_1, n11091_1, n11079_0, n11072_0, n11067_0, n11060_0, n11038_0, n11028_0/**/, n10975_0, n3898, n3890, n2918, n2910}), .out(n13147), .config_in(config_chain[29253:29248]), .config_rst(config_rst)); 
buffer_wire buffer_13147 (.in(n13147), .out(n13147_0));
mux15 mux_7982 (.in({n13110_0, n10053_1, n10051_0, n10046_0/**/, n10025_0, n10020_0, n10006_0, n9947_0, n9930_0, n9928_0, n3608, n3600, n3592, n2624, n2616}), .out(n13148), .config_in(config_chain[29259:29254]), .config_rst(config_rst)); 
buffer_wire buffer_13148 (.in(n13148), .out(n13148_0));
mux13 mux_7983 (.in({n13229_1, n11089_1, n11087_0, n11080_0, n11053_0, n11040_0, n11036_0, n11007_0, n10982_0, n3898, n3890/**/, n2922, n2910}), .out(n13149), .config_in(config_chain[29265:29260]), .config_rst(config_rst)); 
buffer_wire buffer_13149 (.in(n13149), .out(n13149_0));
mux16 mux_7984 (.in({n13040_0/**/, n10311_1, n10304_0, n10289_0, n10281_0, n10276_0, n10264_0, n10257_0, n10205_0, n10188_0, n10178_0, n3702, n3694, n2726, n2718, n2710}), .out(n13150), .config_in(config_chain[29271:29266]), .config_rst(config_rst)); 
buffer_wire buffer_13150 (.in(n13150), .out(n13150_0));
mux15 mux_7985 (.in({n13233_0, n11373_1, n11339_0, n11332_0, n11325_0, n11318_0, n11308_0, n11305_0, n11280_0, n11230_0, n3996, n3988, n3020, n3012, n3004}), .out(n13151), .config_in(config_chain[29277:29272]), .config_rst(config_rst)); 
buffer_wire buffer_13151 (.in(n13151), .out(n13151_0));
mux16 mux_7986 (.in({n13048_0/**/, n10313_1, n10303_0, n10298_0, n10275_0, n10270_0, n10266_0, n10259_1, n10250_0, n10244_0, n10181_0, n3702, n3694, n2726, n2718, n2710}), .out(n13152), .config_in(config_chain[29283:29278]), .config_rst(config_rst)); 
buffer_wire buffer_13152 (.in(n13152), .out(n13152_0));
mux15 mux_7987 (.in({n13235_0/**/, n11371_1, n11347_0, n11340_0, n11326_0, n11310_0, n11307_0, n11249_0, n11238_0, n11224_0, n4000, n3988, n3020, n3012, n3004}), .out(n13153), .config_in(config_chain[29289:29284]), .config_rst(config_rst)); 
buffer_wire buffer_13153 (.in(n13153), .out(n13153_0));
mux15 mux_7988 (.in({n13056_0/**/, n10315_1, n10297_0, n10292_0, n10284_0, n10269_0, n10261_1, n10242_0, n10237_0, n10220_0, n3702, n3694, n2726, n2718, n2710}), .out(n13154), .config_in(config_chain[29295:29290]), .config_rst(config_rst)); 
buffer_wire buffer_13154 (.in(n13154), .out(n13154_0));
mux15 mux_7989 (.in({n13237_0, n11369_1, n11348_0, n11333_0/**/, n11319_0, n11312_0, n11309_0, n11281_0, n11256_0, n11246_0, n4000, n3992, n3020, n3012, n3004}), .out(n13155), .config_in(config_chain[29301:29296]), .config_rst(config_rst)); 
buffer_wire buffer_13155 (.in(n13155), .out(n13155_0));
mux15 mux_7990 (.in({n13064_0, n10317_1, n10306_0, n10291_0, n10283_0, n10278_0, n10263_1, n10234_0, n10213_0, n10196_0, n3702, n3694, n2726, n2718, n2710/**/}), .out(n13156), .config_in(config_chain[29307:29302]), .config_rst(config_rst)); 
buffer_wire buffer_13156 (.in(n13156), .out(n13156_0));
mux15 mux_7991 (.in({n13239_0, n11367_1, n11341_0/**/, n11334_0, n11327_0, n11320_0, n11311_1, n11288_0, n11254_0, n11225_0, n4000, n3992, n3984, n3012, n3004}), .out(n13157), .config_in(config_chain[29313:29308]), .config_rst(config_rst)); 
buffer_wire buffer_13157 (.in(n13157), .out(n13157_0));
mux15 mux_7992 (.in({n13072_0, n10319_1, n10305_0/**/, n10300_0, n10277_0, n10272_0, n10265_1, n10252_0, n10226_0, n10189_0, n3702, n3694, n2726, n2718, n2710}), .out(n13158), .config_in(config_chain[29319:29314]), .config_rst(config_rst)); 
buffer_wire buffer_13158 (.in(n13158), .out(n13158_0));
mux14 mux_7993 (.in({n13241_0, n11365_1, n11349_0, n11342_0, n11328_0, n11313_0, n11262_0, n11257_0, n11232_0, n4000/**/, n3992, n3984, n3016, n3004}), .out(n13159), .config_in(config_chain[29325:29320]), .config_rst(config_rst)); 
buffer_wire buffer_13159 (.in(n13159), .out(n13159_0));
mux15 mux_7994 (.in({n13080_0/**/, n10321_1, n10299_0, n10294_0, n10286_0, n10271_0, n10267_1, n10245_0, n10228_0, n10218_0, n3706, n3698, n3690, n2722, n2714}), .out(n13160), .config_in(config_chain[29331:29326]), .config_rst(config_rst)); 
buffer_wire buffer_13160 (.in(n13160), .out(n13160_0));
mux14 mux_7995 (.in({n13243_0, n11363_1, n11350_0, n11335_0, n11321_0/**/, n11314_0, n11289_0, n11270_0, n11264_0, n4000, n3992, n3984, n3016, n3008}), .out(n13161), .config_in(config_chain[29337:29332]), .config_rst(config_rst)); 
buffer_wire buffer_13161 (.in(n13161), .out(n13161_0));
mux15 mux_7996 (.in({n13088_0, n10323_1, n10293_0, n10288_0, n10285_0, n10280_0, n10256_0, n10221_0, n10210_0/**/, n10204_0, n3706, n3698, n3690, n2722, n2714}), .out(n13162), .config_in(config_chain[29343:29338]), .config_rst(config_rst)); 
buffer_wire buffer_13162 (.in(n13162), .out(n13162_0));
mux13 mux_7997 (.in({n13245_0, n11361_1, n11343_0, n11336_0, n11329_0, n11322_0, n11296_0, n11278_0, n11233_0, n3992, n3984, n3016/**/, n3008}), .out(n13163), .config_in(config_chain[29349:29344]), .config_rst(config_rst)); 
buffer_wire buffer_13163 (.in(n13163), .out(n13163_0));
mux15 mux_7998 (.in({n13096_0/**/, n10325_1, n10307_0, n10302_0, n10279_0, n10274_0, n10258_0, n10202_0, n10197_0, n10180_0, n3706, n3698, n3690, n2722, n2714}), .out(n13164), .config_in(config_chain[29355:29350]), .config_rst(config_rst)); 
buffer_wire buffer_13164 (.in(n13164), .out(n13164_0));
mux13 mux_7999 (.in({n13247_0, n11359_1, n11351_0, n11344_0/**/, n11330_0, n11315_0, n11286_0, n11265_0, n11240_0, n3996, n3984, n3016, n3008}), .out(n13165), .config_in(config_chain[29361:29356]), .config_rst(config_rst)); 
buffer_wire buffer_13165 (.in(n13165), .out(n13165_0));
mux15 mux_8000 (.in({n13104_0/**/, n10327_1, n10301_0, n10296_0, n10273_0, n10268_0, n10260_0, n10253_0, n10236_0, n10194_0, n3706, n3698, n3690, n2722, n2714}), .out(n13166), .config_in(config_chain[29367:29362]), .config_rst(config_rst)); 
buffer_wire buffer_13166 (.in(n13166), .out(n13166_0));
mux13 mux_8001 (.in({n13249_0, n11357_1, n11352_0, n11337_0, n11323_0, n11316_0, n11297_0, n11294_0, n11272_0, n3996, n3988/**/, n3016, n3008}), .out(n13167), .config_in(config_chain[29373:29368]), .config_rst(config_rst)); 
buffer_wire buffer_13167 (.in(n13167), .out(n13167_0));
mux15 mux_8002 (.in({n13112_0, n10309_1, n10295_0, n10290_0, n10287_0, n10282_0, n10262_0, n10229_0/**/, n10212_0, n10186_0, n3706, n3698, n3690, n2722, n2714}), .out(n13168), .config_in(config_chain[29379:29374]), .config_rst(config_rst)); 
buffer_wire buffer_13168 (.in(n13168), .out(n13168_0));
mux13 mux_8003 (.in({n13251_0, n11355_1, n11345_0, n11338_0, n11331_0, n11324_0, n11304_0, n11302_0, n11241_0, n3996, n3988, n3020/**/, n3008}), .out(n13169), .config_in(config_chain[29385:29380]), .config_rst(config_rst)); 
buffer_wire buffer_13169 (.in(n13169), .out(n13169_0));
mux16 mux_8004 (.in({n13042_0, n10569_1, n10553_0, n10548_0, n10542_0, n10527_0, n10522_0, n10515_0, n10489_0, n10472_0, n10438_0, n3800, n3792, n2824, n2816, n2808}), .out(n13170), .config_in(config_chain[29391:29386]), .config_rst(config_rst)); 
buffer_wire buffer_13170 (.in(n13170), .out(n13170_0));
mux15 mux_8005 (.in({n13255_0/**/, n11639_1, n11619_1, n11612_0, n11583_0, n11576_0, n11572_0, n11539_0, n11514_0, n11496_0, n4094, n4086, n3118, n3110, n3102}), .out(n13171), .config_in(config_chain[29397:29392]), .config_rst(config_rst)); 
buffer_wire buffer_13171 (.in(n13171), .out(n13171_0));
mux16 mux_8006 (.in({n13050_0, n10571_1, n10562_0, n10547_0, n10541_0, n10536_0, n10524_0, n10517_0/**/, n10510_0, n10465_0, n10448_0, n3800, n3792, n2824, n2816, n2808}), .out(n13172), .config_in(config_chain[29403:29398]), .config_rst(config_rst)); 
buffer_wire buffer_13172 (.in(n13172), .out(n13172_0));
mux15 mux_8007 (.in({n13257_0, n11637_1, n11605_0, n11598_0, n11591_0/**/, n11584_0, n11574_0, n11571_0, n11546_0, n11504_0, n4098, n4086, n3118, n3110, n3102}), .out(n13173), .config_in(config_chain[29409:29404]), .config_rst(config_rst)); 
buffer_wire buffer_13173 (.in(n13173), .out(n13173_0));
mux15 mux_8008 (.in({n13058_0, n10573_1, n10561_0, n10556_0, n10535_0, n10530_0, n10519_1, n10504_0, n10502_0, n10441_0, n3800/**/, n3792, n2824, n2816, n2808}), .out(n13174), .config_in(config_chain[29415:29410]), .config_rst(config_rst)); 
buffer_wire buffer_13174 (.in(n13174), .out(n13174_0));
mux15 mux_8009 (.in({n13259_0, n11635_1, n11613_0, n11606_0, n11592_0, n11577_0, n11573_0, n11515_0, n11512_0, n11490_0, n4098, n4090, n3118, n3110, n3102}), .out(n13175), .config_in(config_chain[29421:29416]), .config_rst(config_rst)); 
buffer_wire buffer_13175 (.in(n13175), .out(n13175_0));
mux15 mux_8010 (.in({n13066_0/**/, n10575_1, n10555_0, n10550_0, n10544_0, n10529_0, n10521_1, n10497_0, n10494_0, n10480_0, n3800, n3792, n2824, n2816, n2808}), .out(n13176), .config_in(config_chain[29427:29422]), .config_rst(config_rst)); 
buffer_wire buffer_13176 (.in(n13176), .out(n13176_0));
mux15 mux_8011 (.in({n13261_0, n11633_1, n11614_0, n11599_0, n11585_0, n11578_0/**/, n11575_0, n11547_0, n11522_0, n11520_0, n4098, n4090, n4082, n3110, n3102}), .out(n13177), .config_in(config_chain[29433:29428]), .config_rst(config_rst)); 
buffer_wire buffer_13177 (.in(n13177), .out(n13177_0));
mux15 mux_8012 (.in({n13074_0/**/, n10577_1, n10564_0, n10549_0, n10543_0, n10538_0, n10523_1, n10486_0, n10473_0, n10456_0, n3800, n3792, n2824, n2816, n2808}), .out(n13178), .config_in(config_chain[29439:29434]), .config_rst(config_rst)); 
buffer_wire buffer_13178 (.in(n13178), .out(n13178_0));
mux14 mux_8013 (.in({n13263_0, n11631_1, n11607_0, n11600_0, n11593_0, n11586_0, n11554_0, n11528_0, n11491_0/**/, n4098, n4090, n4082, n3114, n3102}), .out(n13179), .config_in(config_chain[29445:29440]), .config_rst(config_rst)); 
buffer_wire buffer_13179 (.in(n13179), .out(n13179_0));
mux15 mux_8014 (.in({n13082_0, n10579_1, n10563_0, n10558_0, n10537_0, n10532_0, n10525_1, n10512_0, n10478_0, n10449_0, n3804, n3796, n3788/**/, n2820, n2812}), .out(n13180), .config_in(config_chain[29451:29446]), .config_rst(config_rst)); 
buffer_wire buffer_13180 (.in(n13180), .out(n13180_0));
mux14 mux_8015 (.in({n13265_0, n11629_1, n11615_0, n11608_0, n11594_0, n11579_0, n11536_0, n11523_0, n11498_0, n4098, n4090, n4082/**/, n3114, n3106}), .out(n13181), .config_in(config_chain[29457:29452]), .config_rst(config_rst)); 
buffer_wire buffer_13181 (.in(n13181), .out(n13181_0));
mux15 mux_8016 (.in({n13090_0, n10581_1, n10557_0, n10552_0, n10531_0, n10526_0, n10514_0, n10505_0, n10488_0, n10470_0, n3804, n3796, n3788, n2820/**/, n2812}), .out(n13182), .config_in(config_chain[29463:29458]), .config_rst(config_rst)); 
buffer_wire buffer_13182 (.in(n13182), .out(n13182_0));
mux13 mux_8017 (.in({n13267_0, n11627_1, n11616_0, n11601_0, n11587_0, n11580_0, n11555_0/**/, n11544_0, n11530_0, n4090, n4082, n3114, n3106}), .out(n13183), .config_in(config_chain[29469:29464]), .config_rst(config_rst)); 
buffer_wire buffer_13183 (.in(n13183), .out(n13183_0));
mux15 mux_8018 (.in({n13098_0, n10583_1/**/, n10551_0, n10546_0, n10545_0, n10540_0, n10516_0, n10481_0, n10464_0, n10462_0, n3804, n3796, n3788, n2820, n2812}), .out(n13184), .config_in(config_chain[29475:29470]), .config_rst(config_rst)); 
buffer_wire buffer_13184 (.in(n13184), .out(n13184_0));
mux13 mux_8019 (.in({n13269_0, n11625_1, n11609_0, n11602_0, n11595_0, n11588_0, n11562_0, n11552_0, n11499_0, n4094, n4082, n3114/**/, n3106}), .out(n13185), .config_in(config_chain[29481:29476]), .config_rst(config_rst)); 
buffer_wire buffer_13185 (.in(n13185), .out(n13185_0));
mux15 mux_8020 (.in({n13106_0, n10585_1, n10565_0, n10560_0, n10539_0, n10534_0, n10518_0, n10457_0, n10454_0, n10440_0, n3804, n3796, n3788/**/, n2820, n2812}), .out(n13186), .config_in(config_chain[29487:29482]), .config_rst(config_rst)); 
buffer_wire buffer_13186 (.in(n13186), .out(n13186_0));
mux13 mux_8021 (.in({n13271_0, n11623_1, n11617_0, n11610_0, n11596_0, n11581_0, n11560_0, n11531_0/**/, n11506_0, n4094, n4086, n3114, n3106}), .out(n13187), .config_in(config_chain[29493:29488]), .config_rst(config_rst)); 
buffer_wire buffer_13187 (.in(n13187), .out(n13187_0));
mux15 mux_8022 (.in({n13114_0, n10567_1, n10559_0, n10554_0/**/, n10533_0, n10528_0, n10520_0, n10513_0, n10496_0, n10446_0, n3804, n3796, n3788, n2820, n2812}), .out(n13188), .config_in(config_chain[29499:29494]), .config_rst(config_rst)); 
buffer_wire buffer_13188 (.in(n13188), .out(n13188_0));
mux13 mux_8023 (.in({n13273_0/**/, n11621_1, n11618_0, n11603_0, n11589_0, n11582_0, n11568_0, n11563_0, n11538_0, n4094, n4086, n3118, n3106}), .out(n13189), .config_in(config_chain[29505:29500]), .config_rst(config_rst)); 
buffer_wire buffer_13189 (.in(n13189), .out(n13189_0));
mux16 mux_8024 (.in({n13044_1, n10829_1, n10819_0, n10814_0, n10793_0, n10788_0, n10782_0, n10775_0, n10758_0, n10700_0, n10695_0, n3898, n3890, n2922, n2914, n2906}), .out(n13190), .config_in(config_chain[29511:29506]), .config_rst(config_rst)); 
buffer_wire buffer_13190 (.in(n13190), .out(n13190_0));
mux15 mux_8025 (.in({n13277_0, n11903_1, n11875_0, n11868_0, n11861_1, n11854_0, n11836_0, n11773_0, n11762_0, n11748_0, n4192, n4184, n3216, n3208, n3200/**/}), .out(n13191), .config_in(config_chain[29517:29512]), .config_rst(config_rst)); 
buffer_wire buffer_13191 (.in(n13191), .out(n13191_0));
mux16 mux_8026 (.in({n13052_1, n10831_1, n10813_0, n10808_0, n10802_0, n10787_0, n10784_0, n10777_0, n10772_0, n10751_0, n10734_0, n3898, n3890/**/, n2922, n2914, n2906}), .out(n13192), .config_in(config_chain[29523:29518]), .config_rst(config_rst)); 
buffer_wire buffer_13192 (.in(n13192), .out(n13192_0));
mux15 mux_8027 (.in({n13279_0, n11901_1, n11883_1, n11876_0, n11847_0, n11840_0, n11838_0, n11805_0, n11780_0, n11770_0/**/, n4196, n4184, n3216, n3208, n3200}), .out(n13193), .config_in(config_chain[29529:29524]), .config_rst(config_rst)); 
buffer_wire buffer_13193 (.in(n13193), .out(n13193_0));
mux15 mux_8028 (.in({n13060_1, n10833_1/**/, n10822_0, n10807_0, n10801_0, n10796_0, n10779_0, n10764_0, n10727_0, n10710_0, n3898, n3890, n2922, n2914, n2906}), .out(n13194), .config_in(config_chain[29535:29530]), .config_rst(config_rst)); 
buffer_wire buffer_13194 (.in(n13194), .out(n13194_0));
mux15 mux_8029 (.in({n13281_0/**/, n11899_1, n11869_0, n11862_0, n11855_0, n11848_0, n11837_0, n11812_0, n11778_0, n11749_0, n4196, n4188, n3216, n3208, n3200}), .out(n13195), .config_in(config_chain[29541:29536]), .config_rst(config_rst)); 
buffer_wire buffer_13195 (.in(n13195), .out(n13195_0));
mux15 mux_8030 (.in({n13068_1, n10835_1, n10821_0, n10816_0, n10795_0, n10790_0, n10781_1, n10766_0, n10756_0, n10703_0, n3898, n3890, n2922/**/, n2914, n2906}), .out(n13196), .config_in(config_chain[29547:29542]), .config_rst(config_rst)); 
buffer_wire buffer_13196 (.in(n13196), .out(n13196_0));
mux15 mux_8031 (.in({n13283_0, n11897_1, n11877_0, n11870_0, n11856_0/**/, n11841_0, n11839_0, n11786_0, n11781_0, n11756_0, n4196, n4188, n4180, n3208, n3200}), .out(n13197), .config_in(config_chain[29553:29548]), .config_rst(config_rst)); 
buffer_wire buffer_13197 (.in(n13197), .out(n13197_0));
mux15 mux_8032 (.in({n13076_1, n10837_1/**/, n10815_0, n10810_0, n10804_0, n10789_0, n10783_1, n10759_0, n10748_0, n10742_0, n3898, n3890, n2922, n2914, n2906}), .out(n13198), .config_in(config_chain[29559:29554]), .config_rst(config_rst)); 
buffer_wire buffer_13198 (.in(n13198), .out(n13198_0));
mux14 mux_8033 (.in({n13285_0, n11895_1, n11878_0, n11863_0, n11849_0, n11842_0, n11813_0, n11794_0, n11788_0, n4196, n4188/**/, n4180, n3212, n3200}), .out(n13199), .config_in(config_chain[29565:29560]), .config_rst(config_rst)); 
buffer_wire buffer_13199 (.in(n13199), .out(n13199_0));
mux15 mux_8034 (.in({n13084_1, n10839_1, n10824_0, n10809_0, n10803_0, n10798_0/**/, n10785_1, n10740_0, n10735_0, n10718_0, n3902, n3894, n3886, n2918, n2910}), .out(n13200), .config_in(config_chain[29571:29566]), .config_rst(config_rst)); 
buffer_wire buffer_13200 (.in(n13200), .out(n13200_0));
mux14 mux_8035 (.in({n13287_0, n11893_1, n11871_0, n11864_0, n11857_0, n11850_0, n11820_0/**/, n11802_0, n11757_0, n4196, n4188, n4180, n3212, n3204}), .out(n13201), .config_in(config_chain[29577:29572]), .config_rst(config_rst)); 
buffer_wire buffer_13201 (.in(n13201), .out(n13201_0));
mux15 mux_8036 (.in({n13092_1/**/, n10841_1, n10823_0, n10818_0, n10797_0, n10792_0, n10774_0, n10732_0, n10711_0, n10694_0, n3902, n3894, n3886, n2918, n2910}), .out(n13202), .config_in(config_chain[29583:29578]), .config_rst(config_rst)); 
buffer_wire buffer_13202 (.in(n13202), .out(n13202_0));
mux13 mux_8037 (.in({n13289_0, n11891_1, n11879_0, n11872_0, n11858_0, n11843_0, n11810_0, n11789_0, n11764_0/**/, n4188, n4180, n3212, n3204}), .out(n13203), .config_in(config_chain[29589:29584]), .config_rst(config_rst)); 
buffer_wire buffer_13203 (.in(n13203), .out(n13203_0));
mux15 mux_8038 (.in({n13100_1, n10843_1, n10817_0, n10812_0, n10791_0, n10786_0, n10776_0, n10767_0, n10750_0, n10724_0, n3902/**/, n3894, n3886, n2918, n2910}), .out(n13204), .config_in(config_chain[29595:29590]), .config_rst(config_rst)); 
buffer_wire buffer_13204 (.in(n13204), .out(n13204_0));
mux13 mux_8039 (.in({n13291_0, n11889_1, n11880_0, n11865_0, n11851_0, n11844_0, n11821_0, n11818_0, n11796_0/**/, n4192, n4180, n3212, n3204}), .out(n13205), .config_in(config_chain[29601:29596]), .config_rst(config_rst)); 
buffer_wire buffer_13205 (.in(n13205), .out(n13205_0));
mux15 mux_8040 (.in({n13108_1, n10845_1, n10811_0, n10806_0, n10805_0, n10800_0, n10778_0, n10743_0, n10726_0, n10716_0, n3902, n3894, n3886, n2918, n2910}), .out(n13206), .config_in(config_chain[29607:29602]), .config_rst(config_rst)); 
buffer_wire buffer_13206 (.in(n13206), .out(n13206_0));
mux13 mux_8041 (.in({n13293_0/**/, n11887_1, n11873_0, n11866_0, n11859_0, n11852_0, n11828_0, n11826_0, n11765_0, n4192, n4184, n3212, n3204}), .out(n13207), .config_in(config_chain[29613:29608]), .config_rst(config_rst)); 
buffer_wire buffer_13207 (.in(n13207), .out(n13207_0));
mux15 mux_8042 (.in({n13116_1, n10827_1, n10825_0, n10820_0, n10799_0, n10794_0, n10780_0, n10719_0, n10708_0, n10702_0, n3902, n3894, n3886, n2918/**/, n2910}), .out(n13208), .config_in(config_chain[29619:29614]), .config_rst(config_rst)); 
buffer_wire buffer_13208 (.in(n13208), .out(n13208_0));
mux13 mux_8043 (.in({n13295_0, n11885_1/**/, n11881_0, n11874_0, n11860_0, n11845_0, n11834_0, n11797_0, n11772_0, n4192, n4184, n3216, n3204}), .out(n13209), .config_in(config_chain[29625:29620]), .config_rst(config_rst)); 
buffer_wire buffer_13209 (.in(n13209), .out(n13209_0));
mux15 mux_8044 (.in({n13130_1/**/, n11091_1, n11080_0, n11075_0, n11063_0, n11045_1, n11040_0, n10982_0, n10959_0, n10956_0, n3996, n3988, n3020, n3012, n3004}), .out(n13210), .config_in(config_chain[29631:29626]), .config_rst(config_rst)); 
buffer_wire buffer_13210 (.in(n13210), .out(n13210_0));
mux4 mux_8045 (.in({n12147_1, n12010_0, n4294, n3298}), .out(n13211), .config_in(config_chain[29633:29632]), .config_rst(config_rst)); 
buffer_wire buffer_13211 (.in(n13211), .out(n13211_0));
mux15 mux_8046 (.in({n13132_1/**/, n11093_1, n11083_0, n11054_0, n11049_0, n11047_1, n11042_0, n11036_0, n11014_0, n10991_0, n4000, n3988, n3020, n3012, n3004}), .out(n13212), .config_in(config_chain[29639:29634]), .config_rst(config_rst)); 
buffer_wire buffer_13212 (.in(n13212), .out(n13212_0));
mux3 mux_8047 (.in({n12149_1/**/, n12018_0, n3298}), .out(n13213), .config_in(config_chain[29641:29640]), .config_rst(config_rst)); 
buffer_wire buffer_13213 (.in(n13213), .out(n13213_0));
mux15 mux_8048 (.in({n13134_1, n11095_1, n11074_0, n11069_0, n11062_0, n11057_0, n11044_0, n11028_0, n11023_0, n10958_0, n4000, n3992/**/, n3020, n3012, n3004}), .out(n13214), .config_in(config_chain[29647:29642]), .config_rst(config_rst)); 
buffer_wire buffer_13214 (.in(n13214), .out(n13214_0));
mux3 mux_8049 (.in({n12151_1, n12026_0/**/, n3302}), .out(n13215), .config_in(config_chain[29649:29648]), .config_rst(config_rst)); 
buffer_wire buffer_13215 (.in(n13215), .out(n13215_0));
mux15 mux_8050 (.in({n13136_1, n11097_1, n11082_0, n11077_0, n11065_0, n11048_0, n11046_0, n11020_0/**/, n10990_0, n10967_0, n4000, n3992, n3984, n3012, n3004}), .out(n13216), .config_in(config_chain[29655:29650]), .config_rst(config_rst)); 
buffer_wire buffer_13216 (.in(n13216), .out(n13216_0));
mux3 mux_8051 (.in({n12153_1/**/, n12034_0, n3306}), .out(n13217), .config_in(config_chain[29657:29656]), .config_rst(config_rst)); 
buffer_wire buffer_13217 (.in(n13217), .out(n13217_0));
mux14 mux_8052 (.in({n13138_1, n11099_1, n11085_0, n11068_0, n11056_0, n11051_0, n11022_0, n11012_0, n10999_0, n4000, n3992/**/, n3984, n3016, n3004}), .out(n13218), .config_in(config_chain[29663:29658]), .config_rst(config_rst)); 
buffer_wire buffer_13218 (.in(n13218), .out(n13218_0));
mux3 mux_8053 (.in({n12155_1, n12042_0, n3310/**/}), .out(n13219), .config_in(config_chain[29665:29664]), .config_rst(config_rst)); 
buffer_wire buffer_13219 (.in(n13219), .out(n13219_0));
mux14 mux_8054 (.in({n13140_1, n11101_1, n11076_0, n11071_0, n11064_0, n11059_0, n11031_0, n11004_0, n10966_0, n4000, n3992, n3984, n3016/**/, n3008}), .out(n13220), .config_in(config_chain[29671:29666]), .config_rst(config_rst)); 
buffer_wire buffer_13220 (.in(n13220), .out(n13220_0));
mux3 mux_8055 (.in({n12157_1, n12050_0, n3314}), .out(n13221), .config_in(config_chain[29673:29672]), .config_rst(config_rst)); 
buffer_wire buffer_13221 (.in(n13221), .out(n13221_0));
mux13 mux_8056 (.in({n13142_1, n11103_1, n11084_0, n11079_0/**/, n11067_0, n11050_0, n10998_0, n10996_0, n10975_0, n3992, n3984, n3016, n3008}), .out(n13222), .config_in(config_chain[29679:29674]), .config_rst(config_rst)); 
buffer_wire buffer_13222 (.in(n13222), .out(n13222_0));
mux3 mux_8057 (.in({n12159_1/**/, n12058_0, n3314}), .out(n13223), .config_in(config_chain[29681:29680]), .config_rst(config_rst)); 
buffer_wire buffer_13223 (.in(n13223), .out(n13223_0));
mux13 mux_8058 (.in({n13144_1, n11105_1/**/, n11087_0, n11070_0, n11058_0, n11053_0, n11030_0, n11007_0, n10988_0, n3996, n3984, n3016, n3008}), .out(n13224), .config_in(config_chain[29687:29682]), .config_rst(config_rst)); 
buffer_wire buffer_13224 (.in(n13224), .out(n13224_0));
mux3 mux_8059 (.in({n12161_1, n12066_0/**/, n4278}), .out(n13225), .config_in(config_chain[29689:29688]), .config_rst(config_rst)); 
buffer_wire buffer_13225 (.in(n13225), .out(n13225_0));
mux13 mux_8060 (.in({n13146_1, n11107_1, n11078_0, n11073_0, n11066_0, n11061_0, n11039_0, n10980_0/**/, n10974_0, n3996, n3988, n3016, n3008}), .out(n13226), .config_in(config_chain[29695:29690]), .config_rst(config_rst)); 
buffer_wire buffer_13226 (.in(n13226), .out(n13226_0));
mux3 mux_8061 (.in({n12163_1, n12074_0, n4282}), .out(n13227), .config_in(config_chain[29697:29696]), .config_rst(config_rst)); 
buffer_wire buffer_13227 (.in(n13227), .out(n13227_0));
mux13 mux_8062 (.in({n13148_1, n11109_1, n11086_0, n11081_0, n11052_0, n11041_0, n11006_0, n10983_0, n10972_0, n3996, n3988/**/, n3020, n3008}), .out(n13228), .config_in(config_chain[29703:29698]), .config_rst(config_rst)); 
buffer_wire buffer_13228 (.in(n13228), .out(n13228_0));
mux3 mux_8063 (.in({n12165_1, n12082_0/**/, n4286}), .out(n13229), .config_in(config_chain[29705:29704]), .config_rst(config_rst)); 
buffer_wire buffer_13229 (.in(n13229), .out(n13229_0));
mux13 mux_8064 (.in({n13118_1, n11089_1, n11072_0, n11060_0, n11055_0, n11043_0, n11038_0, n11015_0/**/, n10964_0, n3996, n3988, n3020, n3012}), .out(n13230), .config_in(config_chain[29711:29706]), .config_rst(config_rst)); 
buffer_wire buffer_13230 (.in(n13230), .out(n13230_0));
mux3 mux_8065 (.in({n12091_1, n12090_0, n4290}), .out(n13231), .config_in(config_chain[29713:29712]), .config_rst(config_rst)); 
buffer_wire buffer_13231 (.in(n13231), .out(n13231_0));
mux15 mux_8066 (.in({n13150_1/**/, n11357_1, n11338_0, n11333_0, n11324_0, n11319_0, n11309_0, n11304_0, n11281_0, n11222_0, n4094, n4086, n3118, n3110, n3102}), .out(n13232), .config_in(config_chain[29719:29714]), .config_rst(config_rst)); 
buffer_wire buffer_13232 (.in(n13232), .out(n13232_0));
mux4 mux_8067 (.in({n12013_0, n12012_0, n4294, n3298}), .out(n13233), .config_in(config_chain[29721:29720]), .config_rst(config_rst)); 
buffer_wire buffer_13233 (.in(n13233), .out(n13233_0));
mux15 mux_8068 (.in({n13152_1, n11359_1, n11346_0, n11341_0, n11327_0, n11311_1/**/, n11306_0, n11302_0, n11248_0, n11225_0, n4098, n4086, n3118, n3110, n3102}), .out(n13234), .config_in(config_chain[29727:29722]), .config_rst(config_rst)); 
buffer_wire buffer_13234 (.in(n13234), .out(n13234_0));
mux3 mux_8069 (.in({n12021_0/**/, n12020_0, n3302}), .out(n13235), .config_in(config_chain[29729:29728]), .config_rst(config_rst)); 
buffer_wire buffer_13235 (.in(n13235), .out(n13235_0));
mux15 mux_8070 (.in({n13154_1, n11361_1, n11349_0, n11332_0, n11318_0, n11313_0/**/, n11308_0, n11294_0, n11280_0, n11257_0, n4098, n4090, n3118, n3110, n3102}), .out(n13236), .config_in(config_chain[29735:29730]), .config_rst(config_rst)); 
buffer_wire buffer_13236 (.in(n13236), .out(n13236_0));
mux3 mux_8071 (.in({n12029_0, n12028_0/**/, n3302}), .out(n13237), .config_in(config_chain[29737:29736]), .config_rst(config_rst)); 
buffer_wire buffer_13237 (.in(n13237), .out(n13237_0));
mux15 mux_8072 (.in({n13156_1, n11363_1, n11340_0, n11335_0, n11326_0, n11321_0, n11310_0, n11289_0, n11286_0, n11224_0, n4098/**/, n4090, n4082, n3110, n3102}), .out(n13238), .config_in(config_chain[29743:29738]), .config_rst(config_rst)); 
buffer_wire buffer_13238 (.in(n13238), .out(n13238_0));
mux3 mux_8073 (.in({n12037_0/**/, n12036_0, n3306}), .out(n13239), .config_in(config_chain[29745:29744]), .config_rst(config_rst)); 
buffer_wire buffer_13239 (.in(n13239), .out(n13239_0));
mux14 mux_8074 (.in({n13158_1, n11365_1, n11348_0, n11343_0, n11329_0, n11312_0, n11278_0, n11256_0, n11233_0, n4098, n4090, n4082/**/, n3114, n3102}), .out(n13240), .config_in(config_chain[29751:29746]), .config_rst(config_rst)); 
buffer_wire buffer_13240 (.in(n13240), .out(n13240_0));
mux3 mux_8075 (.in({n12045_0, n12044_0, n3310}), .out(n13241), .config_in(config_chain[29753:29752]), .config_rst(config_rst)); 
buffer_wire buffer_13241 (.in(n13241), .out(n13241_0));
mux14 mux_8076 (.in({n13160_1, n11367_1, n11351_0, n11334_0, n11320_0, n11315_0, n11288_0, n11270_0, n11265_0/**/, n4098, n4090, n4082, n3114, n3106}), .out(n13242), .config_in(config_chain[29759:29754]), .config_rst(config_rst)); 
buffer_wire buffer_13242 (.in(n13242), .out(n13242_0));
mux3 mux_8077 (.in({n12053_0/**/, n12052_0, n3314}), .out(n13243), .config_in(config_chain[29761:29760]), .config_rst(config_rst)); 
buffer_wire buffer_13243 (.in(n13243), .out(n13243_0));
mux13 mux_8078 (.in({n13162_1, n11369_1, n11342_0, n11337_0, n11328_0, n11323_0, n11297_0, n11262_0, n11232_0/**/, n4090, n4082, n3114, n3106}), .out(n13244), .config_in(config_chain[29767:29762]), .config_rst(config_rst)); 
buffer_wire buffer_13244 (.in(n13244), .out(n13244_0));
mux3 mux_8079 (.in({n12061_0, n12060_0/**/, n4278}), .out(n13245), .config_in(config_chain[29769:29768]), .config_rst(config_rst)); 
buffer_wire buffer_13245 (.in(n13245), .out(n13245_0));
mux13 mux_8080 (.in({n13164_1, n11371_1, n11350_0, n11345_0, n11331_0, n11314_0, n11264_0/**/, n11254_0, n11241_0, n4094, n4082, n3114, n3106}), .out(n13246), .config_in(config_chain[29775:29770]), .config_rst(config_rst)); 
buffer_wire buffer_13246 (.in(n13246), .out(n13246_0));
mux3 mux_8081 (.in({n12069_0, n12068_0, n4278}), .out(n13247), .config_in(config_chain[29777:29776]), .config_rst(config_rst)); 
buffer_wire buffer_13247 (.in(n13247), .out(n13247_0));
mux13 mux_8082 (.in({n13166_1, n11373_1, n11353_1, n11336_0, n11322_0, n11317_0, n11296_0, n11273_0, n11246_0, n4094, n4086, n3114/**/, n3106}), .out(n13248), .config_in(config_chain[29783:29778]), .config_rst(config_rst)); 
buffer_wire buffer_13248 (.in(n13248), .out(n13248_0));
mux3 mux_8083 (.in({n12077_0, n12076_0, n4282}), .out(n13249), .config_in(config_chain[29785:29784]), .config_rst(config_rst)); 
buffer_wire buffer_13249 (.in(n13249), .out(n13249_0));
mux13 mux_8084 (.in({n13168_1, n11375_1, n11344_0, n11339_0, n11330_0, n11325_0/**/, n11305_0, n11240_0, n11238_0, n4094, n4086, n3118, n3106}), .out(n13250), .config_in(config_chain[29791:29786]), .config_rst(config_rst)); 
buffer_wire buffer_13250 (.in(n13250), .out(n13250_0));
mux3 mux_8085 (.in({n12085_0, n12084_0, n4286}), .out(n13251), .config_in(config_chain[29793:29792]), .config_rst(config_rst)); 
buffer_wire buffer_13251 (.in(n13251), .out(n13251_0));
mux13 mux_8086 (.in({n13120_1, n11355_1, n11352_0, n11347_0, n11316_0, n11307_0, n11272_0, n11249_0/**/, n11230_0, n4094, n4086, n3118, n3110}), .out(n13252), .config_in(config_chain[29799:29794]), .config_rst(config_rst)); 
buffer_wire buffer_13252 (.in(n13252), .out(n13252_0));
mux3 mux_8087 (.in({n12093_1, n12092_0, n4290}), .out(n13253), .config_in(config_chain[29801:29800]), .config_rst(config_rst)); 
buffer_wire buffer_13253 (.in(n13253), .out(n13253_0));
mux15 mux_8088 (.in({n13170_1, n11623_1, n11618_0, n11613_0, n11582_0, n11577_0, n11573_0, n11538_0, n11515_0, n11488_0, n4192, n4184, n3216, n3208, n3200/**/}), .out(n13254), .config_in(config_chain[29807:29802]), .config_rst(config_rst)); 
buffer_wire buffer_13254 (.in(n13254), .out(n13254_0));
mux4 mux_8089 (.in({n12103_0, n12102_0, n4294, n3298/**/}), .out(n13255), .config_in(config_chain[29809:29808]), .config_rst(config_rst)); 
buffer_wire buffer_13255 (.in(n13255), .out(n13255_0));
mux15 mux_8090 (.in({n13172_1, n11625_1, n11604_0, n11599_0, n11590_0, n11585_0, n11575_0, n11570_0, n11568_0, n11547_0/**/, n4196, n4184, n3216, n3208, n3200}), .out(n13256), .config_in(config_chain[29815:29810]), .config_rst(config_rst)); 
buffer_wire buffer_13256 (.in(n13256), .out(n13256_0));
mux3 mux_8091 (.in({n12105_0, n12104_0, n3302}), .out(n13257), .config_in(config_chain[29817:29816]), .config_rst(config_rst)); 
buffer_wire buffer_13257 (.in(n13257), .out(n13257_0));
mux15 mux_8092 (.in({n13174_1, n11627_1, n11612_0, n11607_0, n11593_0, n11576_0, n11572_0, n11560_0, n11514_0, n11491_0, n4196/**/, n4188, n3216, n3208, n3200}), .out(n13258), .config_in(config_chain[29823:29818]), .config_rst(config_rst)); 
buffer_wire buffer_13258 (.in(n13258), .out(n13258_0));
mux3 mux_8093 (.in({n12107_0, n12106_0, n3306}), .out(n13259), .config_in(config_chain[29825:29824]), .config_rst(config_rst)); 
buffer_wire buffer_13259 (.in(n13259), .out(n13259_0));
mux15 mux_8094 (.in({n13176_1, n11629_1, n11615_0, n11598_0, n11584_0, n11579_0, n11574_0, n11552_0, n11546_0, n11523_0/**/, n4196, n4188, n4180, n3208, n3200}), .out(n13260), .config_in(config_chain[29831:29826]), .config_rst(config_rst)); 
buffer_wire buffer_13260 (.in(n13260), .out(n13260_0));
mux3 mux_8095 (.in({n12109_0, n12108_0, n3306}), .out(n13261), .config_in(config_chain[29833:29832]), .config_rst(config_rst)); 
buffer_wire buffer_13261 (.in(n13261), .out(n13261_0));
mux14 mux_8096 (.in({n13178_1, n11631_1, n11606_0, n11601_0, n11592_0, n11587_0, n11555_0, n11544_0, n11490_0, n4196, n4188, n4180, n3212, n3200/**/}), .out(n13262), .config_in(config_chain[29839:29834]), .config_rst(config_rst)); 
buffer_wire buffer_13262 (.in(n13262), .out(n13262_0));
mux3 mux_8097 (.in({n12111_0, n12110_0, n3310}), .out(n13263), .config_in(config_chain[29841:29840]), .config_rst(config_rst)); 
buffer_wire buffer_13263 (.in(n13263), .out(n13263_0));
mux14 mux_8098 (.in({n13180_1, n11633_1, n11614_0, n11609_0/**/, n11595_0, n11578_0, n11536_0, n11522_0, n11499_0, n4196, n4188, n4180, n3212, n3204}), .out(n13264), .config_in(config_chain[29847:29842]), .config_rst(config_rst)); 
buffer_wire buffer_13264 (.in(n13264), .out(n13264_0));
mux3 mux_8099 (.in({n12113_0/**/, n12112_0, n3314}), .out(n13265), .config_in(config_chain[29849:29848]), .config_rst(config_rst)); 
buffer_wire buffer_13265 (.in(n13265), .out(n13265_0));
mux13 mux_8100 (.in({n13182_1, n11635_1, n11617_0, n11600_0, n11586_0, n11581_0, n11554_0, n11531_0, n11528_0, n4188, n4180, n3212, n3204}), .out(n13266), .config_in(config_chain[29855:29850]), .config_rst(config_rst)); 
buffer_wire buffer_13266 (.in(n13266), .out(n13266_0));
mux3 mux_8101 (.in({n12115_0, n12114_0, n4278}), .out(n13267), .config_in(config_chain[29857:29856]), .config_rst(config_rst)); 
buffer_wire buffer_13267 (.in(n13267), .out(n13267_0));
mux13 mux_8102 (.in({n13184_1, n11637_1, n11608_0, n11603_0, n11594_0, n11589_0, n11563_0, n11520_0/**/, n11498_0, n4192, n4180, n3212, n3204}), .out(n13268), .config_in(config_chain[29863:29858]), .config_rst(config_rst)); 
buffer_wire buffer_13268 (.in(n13268), .out(n13268_0));
mux3 mux_8103 (.in({n12117_0, n12116_0/**/, n4282}), .out(n13269), .config_in(config_chain[29865:29864]), .config_rst(config_rst)); 
buffer_wire buffer_13269 (.in(n13269), .out(n13269_0));
mux13 mux_8104 (.in({n13186_1/**/, n11639_1, n11616_0, n11611_0, n11597_1, n11580_0, n11530_0, n11512_0, n11507_0, n4192, n4184, n3212, n3204}), .out(n13270), .config_in(config_chain[29871:29866]), .config_rst(config_rst)); 
buffer_wire buffer_13270 (.in(n13270), .out(n13270_0));
mux3 mux_8105 (.in({n12119_0/**/, n12118_0, n4282}), .out(n13271), .config_in(config_chain[29873:29872]), .config_rst(config_rst)); 
buffer_wire buffer_13271 (.in(n13271), .out(n13271_0));
mux13 mux_8106 (.in({n13188_1/**/, n11641_1, n11619_1, n11602_0, n11588_0, n11583_0, n11562_0, n11539_0, n11504_0, n4192, n4184, n3216, n3204}), .out(n13272), .config_in(config_chain[29879:29874]), .config_rst(config_rst)); 
buffer_wire buffer_13272 (.in(n13272), .out(n13272_0));
mux3 mux_8107 (.in({n12121_0/**/, n12120_0, n4286}), .out(n13273), .config_in(config_chain[29881:29880]), .config_rst(config_rst)); 
buffer_wire buffer_13273 (.in(n13273), .out(n13273_0));
mux13 mux_8108 (.in({n13122_2, n11621_1/**/, n11610_0, n11605_0, n11596_0, n11591_0, n11571_0, n11506_0, n11496_0, n4192, n4184, n3216, n3208}), .out(n13274), .config_in(config_chain[29887:29882]), .config_rst(config_rst)); 
buffer_wire buffer_13274 (.in(n13274), .out(n13274_0));
mux3 mux_8109 (.in({n12123_1, n12122_0/**/, n4290}), .out(n13275), .config_in(config_chain[29889:29888]), .config_rst(config_rst)); 
buffer_wire buffer_13275 (.in(n13275), .out(n13275_0));
mux15 mux_8110 (.in({n13190_1, n11887_1, n11874_0, n11869_0, n11860_0, n11855_0, n11837_0, n11772_0/**/, n11754_0, n11749_0, n4290, n4282, n3314, n3306, n3298}), .out(n13276), .config_in(config_chain[29895:29890]), .config_rst(config_rst)); 
buffer_wire buffer_13276 (.in(n13276), .out(n13276_0));
mux4 mux_8111 (.in({n12125_0, n12124_0, n4294, n3298}), .out(n13277), .config_in(config_chain[29897:29896]), .config_rst(config_rst)); 
buffer_wire buffer_13277 (.in(n13277), .out(n13277_0));
mux15 mux_8112 (.in({n13192_1, n11889_1, n11882_0, n11877_0/**/, n11846_0, n11841_0, n11839_0, n11834_0, n11804_0, n11781_0, n4294, n4282, n3314, n3306, n3298}), .out(n13278), .config_in(config_chain[29903:29898]), .config_rst(config_rst)); 
buffer_wire buffer_13278 (.in(n13278), .out(n13278_0));
mux3 mux_8113 (.in({n12127_0, n12126_0/**/, n3302}), .out(n13279), .config_in(config_chain[29905:29904]), .config_rst(config_rst)); 
buffer_wire buffer_13279 (.in(n13279), .out(n13279_0));
mux15 mux_8114 (.in({n13194_1, n11891_1, n11868_0, n11863_0, n11854_0, n11849_0, n11836_0, n11826_0, n11813_0, n11748_0/**/, n4294, n4286, n3314, n3306, n3298}), .out(n13280), .config_in(config_chain[29911:29906]), .config_rst(config_rst)); 
buffer_wire buffer_13280 (.in(n13280), .out(n13280_0));
mux3 mux_8115 (.in({n12129_0, n12128_0/**/, n3306}), .out(n13281), .config_in(config_chain[29913:29912]), .config_rst(config_rst)); 
buffer_wire buffer_13281 (.in(n13281), .out(n13281_0));
mux15 mux_8116 (.in({n13196_1, n11893_1, n11876_0, n11871_0, n11857_0, n11840_0, n11838_0, n11818_0, n11780_0, n11757_0, n4294/**/, n4286, n4278, n3306, n3298}), .out(n13282), .config_in(config_chain[29919:29914]), .config_rst(config_rst)); 
buffer_wire buffer_13282 (.in(n13282), .out(n13282_0));
mux3 mux_8117 (.in({n12131_0, n12130_0, n3310/**/}), .out(n13283), .config_in(config_chain[29921:29920]), .config_rst(config_rst)); 
buffer_wire buffer_13283 (.in(n13283), .out(n13283_0));
mux14 mux_8118 (.in({n13198_1, n11895_1, n11879_0/**/, n11862_0, n11848_0, n11843_0, n11812_0, n11810_0, n11789_0, n4294, n4286, n4278, n3310, n3298}), .out(n13284), .config_in(config_chain[29927:29922]), .config_rst(config_rst)); 
buffer_wire buffer_13284 (.in(n13284), .out(n13284_0));
mux3 mux_8119 (.in({n12133_0, n12132_0, n3310}), .out(n13285), .config_in(config_chain[29929:29928]), .config_rst(config_rst)); 
buffer_wire buffer_13285 (.in(n13285), .out(n13285_0));
mux14 mux_8120 (.in({n13200_1, n11897_1, n11870_0, n11865_0, n11856_0, n11851_0, n11821_0, n11802_0, n11756_0, n4294, n4286, n4278, n3310, n3302}), .out(n13286), .config_in(config_chain[29935:29930]), .config_rst(config_rst)); 
buffer_wire buffer_13286 (.in(n13286), .out(n13286_0));
mux3 mux_8121 (.in({n12135_0, n12134_0, n3314/**/}), .out(n13287), .config_in(config_chain[29937:29936]), .config_rst(config_rst)); 
buffer_wire buffer_13287 (.in(n13287), .out(n13287_0));
mux13 mux_8122 (.in({n13202_1/**/, n11899_1, n11878_0, n11873_0, n11859_0, n11842_0, n11794_0, n11788_0, n11765_0, n4286, n4278, n3310, n3302}), .out(n13288), .config_in(config_chain[29943:29938]), .config_rst(config_rst)); 
buffer_wire buffer_13288 (.in(n13288), .out(n13288_0));
mux3 mux_8123 (.in({n12137_0, n12136_0, n4278}), .out(n13289), .config_in(config_chain[29945:29944]), .config_rst(config_rst)); 
buffer_wire buffer_13289 (.in(n13289), .out(n13289_0));
mux13 mux_8124 (.in({n13204_1, n11901_1, n11881_0, n11864_0, n11850_0, n11845_0, n11820_0, n11797_0, n11786_0, n4290, n4278, n3310, n3302}), .out(n13290), .config_in(config_chain[29951:29946]), .config_rst(config_rst)); 
buffer_wire buffer_13290 (.in(n13290), .out(n13290_0));
mux3 mux_8125 (.in({n12139_0, n12138_0, n4282}), .out(n13291), .config_in(config_chain[29953:29952]), .config_rst(config_rst)); 
buffer_wire buffer_13291 (.in(n13291), .out(n13291_0));
mux13 mux_8126 (.in({n13206_1, n11903_1, n11872_0, n11867_0, n11858_0, n11853_0, n11829_1, n11778_0, n11764_0, n4290, n4282, n3310, n3302}), .out(n13292), .config_in(config_chain[29959:29954]), .config_rst(config_rst)); 
buffer_wire buffer_13292 (.in(n13292), .out(n13292_0));
mux3 mux_8127 (.in({n12141_0, n12140_0/**/, n4286}), .out(n13293), .config_in(config_chain[29961:29960]), .config_rst(config_rst)); 
buffer_wire buffer_13293 (.in(n13293), .out(n13293_0));
mux13 mux_8128 (.in({n13208_1, n11905_1, n11880_0, n11875_0, n11861_1, n11844_0, n11796_0/**/, n11773_0, n11770_0, n4290, n4282, n3314, n3302}), .out(n13294), .config_in(config_chain[29967:29962]), .config_rst(config_rst)); 
buffer_wire buffer_13294 (.in(n13294), .out(n13294_0));
mux3 mux_8129 (.in({n12143_0, n12142_0, n4286}), .out(n13295), .config_in(config_chain[29969:29968]), .config_rst(config_rst)); 
buffer_wire buffer_13295 (.in(n13295), .out(n13295_0));
mux13 mux_8130 (.in({n13124_2, n11885_1, n11883_1, n11866_0, n11852_0, n11847_0, n11828_0, n11805_0/**/, n11762_0, n4290, n4282, n3314, n3306}), .out(n13296), .config_in(config_chain[29975:29970]), .config_rst(config_rst)); 
buffer_wire buffer_13296 (.in(n13296), .out(n13296_0));
mux3 mux_8131 (.in({n12145_1, n12144_0, n4290}), .out(n13297), .config_in(config_chain[29977:29976]), .config_rst(config_rst)); 
buffer_wire buffer_13297 (.in(n13297), .out(n13297_0));
mux4 mux_8132 (.in({n9819_1, n9666_1, n4488, n3492}), .out(n13298), .config_in(config_chain[29979:29978]), .config_rst(config_rst)); 
buffer_wire buffer_13298 (.in(n13298), .out(n13298_0));
mux15 mux_8133 (.in({n13451_1, n10865_1, n10839_0, n10832_0, n10820_0, n10793_0, n10786_0, n10782_1, n10779_0, n10702_1, n4778, n4770, n3802, n3794, n3786}), .out(n13299), .config_in(config_chain[29985:29980]), .config_rst(config_rst)); 
buffer_wire buffer_13299 (.in(n13299), .out(n13299_0));
mux4 mux_8134 (.in({n9759_0/**/, n9758_0, n4488, n3492}), .out(n13300), .config_in(config_chain[29987:29986]), .config_rst(config_rst)); 
buffer_wire buffer_13300 (.in(n13300), .out(n13300_0));
mux16 mux_8135 (.in({n13391_1, n10089_1, n10069_0, n10052_0, n10044_0, n10041_0/**/, n10018_0, n10015_0, n10009_1, n10000_1, n9930_1, n4484, n4476, n3508, n3500, n3492}), .out(n13301), .config_in(config_chain[29993:29988]), .config_rst(config_rst)); 
buffer_wire buffer_13301 (.in(n13301), .out(n13301_0));
mux4 mux_8136 (.in({n9779_0, n9778_0, n4488, n3492}), .out(n13302), .config_in(config_chain[29995:29994]), .config_rst(config_rst)); 
buffer_wire buffer_13302 (.in(n13302), .out(n13302_0));
mux16 mux_8137 (.in({n13411_1, n10345_1, n10314_0, n10311_0, n10305_0, n10288_0, n10280_0, n10277_0, n10265_1, n10256_1, n10188_1, n4582, n4574, n3606, n3598, n3590/**/}), .out(n13303), .config_in(config_chain[30001:29996]), .config_rst(config_rst)); 
buffer_wire buffer_13303 (.in(n13303), .out(n13303_0));
mux4 mux_8138 (.in({n9799_0, n9798_0, n4488/**/, n3492}), .out(n13304), .config_in(config_chain[30003:30002]), .config_rst(config_rst)); 
buffer_wire buffer_13304 (.in(n13304), .out(n13304_0));
mux16 mux_8139 (.in({n13431_1, n10603_1, n10578_0, n10575_0, n10552_0, n10549_0, n10543_0, n10526_0, n10523_1, n10514_1, n10448_1, n4680, n4672, n3704, n3696, n3688}), .out(n13305), .config_in(config_chain[30009:30004]), .config_rst(config_rst)); 
buffer_wire buffer_13305 (.in(n13305), .out(n13305_0));
mux3 mux_8140 (.in({n9821_1/**/, n9674_1, n3492}), .out(n13306), .config_in(config_chain[30011:30010]), .config_rst(config_rst)); 
buffer_wire buffer_13306 (.in(n13306), .out(n13306_0));
mux15 mux_8141 (.in({n13453_1, n10863_1, n10840_0, n10813_0/**/, n10806_0, n10801_0, n10794_0, n10784_1, n10781_0, n10710_1, n4782, n4770, n3802, n3794, n3786}), .out(n13307), .config_in(config_chain[30017:30012]), .config_rst(config_rst)); 
buffer_wire buffer_13307 (.in(n13307), .out(n13307_0));
mux3 mux_8142 (.in({n9761_0, n9760_0, n3496}), .out(n13308), .config_in(config_chain[30019:30018]), .config_rst(config_rst)); 
buffer_wire buffer_13308 (.in(n13308), .out(n13308_0));
mux16 mux_8143 (.in({n13393_1, n10087_1/**/, n10066_0, n10063_0, n10038_0, n10035_0, n10029_0, n10012_0, n10011_1, n10002_1, n9938_1, n4484, n4476, n3508, n3500, n3492}), .out(n13309), .config_in(config_chain[30025:30020]), .config_rst(config_rst)); 
buffer_wire buffer_13309 (.in(n13309), .out(n13309_0));
mux3 mux_8144 (.in({n9781_0, n9780_0, n3496}), .out(n13310), .config_in(config_chain[30027:30026]), .config_rst(config_rst)); 
buffer_wire buffer_13310 (.in(n13310), .out(n13310_0));
mux16 mux_8145 (.in({n13413_1, n10343_1, n10325_0, n10308_0, n10302_0, n10299_0, n10274_0, n10271_0, n10267_1, n10258_1, n10196_1, n4582, n4574, n3606, n3598, n3590}), .out(n13311), .config_in(config_chain[30033:30028]), .config_rst(config_rst)); 
buffer_wire buffer_13311 (.in(n13311), .out(n13311_0));
mux3 mux_8146 (.in({n9801_0, n9800_0, n3496/**/}), .out(n13312), .config_in(config_chain[30035:30034]), .config_rst(config_rst)); 
buffer_wire buffer_13312 (.in(n13312), .out(n13312_0));
mux16 mux_8147 (.in({n13433_1/**/, n10601_1, n10572_0, n10569_0, n10563_0, n10546_0, n10540_0, n10537_0, n10525_1, n10516_1, n10456_1, n4680, n4672, n3704, n3696, n3688}), .out(n13313), .config_in(config_chain[30041:30036]), .config_rst(config_rst)); 
buffer_wire buffer_13313 (.in(n13313), .out(n13313_0));
mux3 mux_8148 (.in({n9823_1, n9682_1, n3496/**/}), .out(n13314), .config_in(config_chain[30043:30042]), .config_rst(config_rst)); 
buffer_wire buffer_13314 (.in(n13314), .out(n13314_0));
mux15 mux_8149 (.in({n13455_1, n10861_1, n10833_0, n10826_0, n10821_0, n10814_0, n10802_0/**/, n10787_0, n10783_1, n10718_1, n4782, n4774, n3802, n3794, n3786}), .out(n13315), .config_in(config_chain[30049:30044]), .config_rst(config_rst)); 
buffer_wire buffer_13315 (.in(n13315), .out(n13315_0));
mux3 mux_8150 (.in({n9763_0/**/, n9762_0, n3496}), .out(n13316), .config_in(config_chain[30051:30050]), .config_rst(config_rst)); 
buffer_wire buffer_13316 (.in(n13316), .out(n13316_0));
mux15 mux_8151 (.in({n13395_1, n10085_1, n10060_0, n10057_0, n10049_0, n10032_0, n10026_0, n10023_0, n10004_1, n9946_1, n4484, n4476, n3508/**/, n3500, n3492}), .out(n13317), .config_in(config_chain[30057:30052]), .config_rst(config_rst)); 
buffer_wire buffer_13317 (.in(n13317), .out(n13317_0));
mux3 mux_8152 (.in({n9783_0, n9782_0, n3500}), .out(n13318), .config_in(config_chain[30059:30058]), .config_rst(config_rst)); 
buffer_wire buffer_13318 (.in(n13318), .out(n13318_0));
mux15 mux_8153 (.in({n13415_1, n10341_1, n10322_0, n10319_0, n10296_0, n10293_0, n10285_0, n10268_0, n10260_1, n10204_1, n4582, n4574/**/, n3606, n3598, n3590}), .out(n13319), .config_in(config_chain[30065:30060]), .config_rst(config_rst)); 
buffer_wire buffer_13319 (.in(n13319), .out(n13319_0));
mux3 mux_8154 (.in({n9803_0, n9802_0/**/, n3500}), .out(n13320), .config_in(config_chain[30067:30066]), .config_rst(config_rst)); 
buffer_wire buffer_13320 (.in(n13320), .out(n13320_0));
mux15 mux_8155 (.in({n13435_1, n10599_1, n10583_0, n10566_0, n10560_0, n10557_0, n10534_0, n10531_0, n10518_1, n10464_1, n4680, n4672, n3704, n3696, n3688/**/}), .out(n13321), .config_in(config_chain[30073:30068]), .config_rst(config_rst)); 
buffer_wire buffer_13321 (.in(n13321), .out(n13321_0));
mux3 mux_8156 (.in({n9825_1/**/, n9690_1, n3500}), .out(n13322), .config_in(config_chain[30075:30074]), .config_rst(config_rst)); 
buffer_wire buffer_13322 (.in(n13322), .out(n13322_0));
mux15 mux_8157 (.in({n13457_1, n10859_1/**/, n10841_0, n10834_0, n10822_0, n10807_0, n10795_0, n10788_0, n10785_1, n10726_1, n4782, n4774, n4766, n3794, n3786}), .out(n13323), .config_in(config_chain[30081:30076]), .config_rst(config_rst)); 
buffer_wire buffer_13323 (.in(n13323), .out(n13323_0));
mux3 mux_8158 (.in({n9765_0, n9764_0, n3500}), .out(n13324), .config_in(config_chain[30083:30082]), .config_rst(config_rst)); 
buffer_wire buffer_13324 (.in(n13324), .out(n13324_0));
mux15 mux_8159 (.in({n13397_1, n10083_1, n10071_0, n10054_0, n10046_0, n10043_0, n10020_0, n10017_0, n10006_1, n9954_1, n4484, n4476, n3508, n3500, n3492}), .out(n13325), .config_in(config_chain[30089:30084]), .config_rst(config_rst)); 
buffer_wire buffer_13325 (.in(n13325), .out(n13325_0));
mux3 mux_8160 (.in({n9785_0, n9784_0, n3500}), .out(n13326), .config_in(config_chain[30091:30090]), .config_rst(config_rst)); 
buffer_wire buffer_13326 (.in(n13326), .out(n13326_0));
mux15 mux_8161 (.in({n13417_1, n10339_1, n10316_0, n10313_0, n10307_0, n10290_0, n10282_0, n10279_0, n10262_1, n10212_1, n4582, n4574/**/, n3606, n3598, n3590}), .out(n13327), .config_in(config_chain[30097:30092]), .config_rst(config_rst)); 
buffer_wire buffer_13327 (.in(n13327), .out(n13327_0));
mux3 mux_8162 (.in({n9805_0, n9804_0, n3504}), .out(n13328), .config_in(config_chain[30099:30098]), .config_rst(config_rst)); 
buffer_wire buffer_13328 (.in(n13328), .out(n13328_0));
mux15 mux_8163 (.in({n13437_1, n10597_1, n10580_0, n10577_0, n10554_0, n10551_0, n10545_0, n10528_0, n10520_1, n10472_1, n4680, n4672, n3704, n3696, n3688/**/}), .out(n13329), .config_in(config_chain[30105:30100]), .config_rst(config_rst)); 
buffer_wire buffer_13329 (.in(n13329), .out(n13329_0));
mux3 mux_8164 (.in({n9827_1, n9698_1, n3504}), .out(n13330), .config_in(config_chain[30107:30106]), .config_rst(config_rst)); 
buffer_wire buffer_13330 (.in(n13330), .out(n13330_0));
mux14 mux_8165 (.in({n13459_1, n10857_1, n10842_0, n10827_0, n10815_0, n10808_0, n10803_0, n10796_0, n10734_1, n4782, n4774/**/, n4766, n3798, n3786}), .out(n13331), .config_in(config_chain[30113:30108]), .config_rst(config_rst)); 
buffer_wire buffer_13331 (.in(n13331), .out(n13331_0));
mux3 mux_8166 (.in({n9767_0/**/, n9766_0, n3504}), .out(n13332), .config_in(config_chain[30115:30114]), .config_rst(config_rst)); 
buffer_wire buffer_13332 (.in(n13332), .out(n13332_0));
mux15 mux_8167 (.in({n13399_1, n10081_1, n10068_0, n10065_0, n10040_0, n10037_0, n10031_0, n10014_0, n10008_1, n9962_1, n4484, n4476, n3508, n3500, n3492}), .out(n13333), .config_in(config_chain[30121:30116]), .config_rst(config_rst)); 
buffer_wire buffer_13333 (.in(n13333), .out(n13333_0));
mux3 mux_8168 (.in({n9787_0, n9786_0, n3504}), .out(n13334), .config_in(config_chain[30123:30122]), .config_rst(config_rst)); 
buffer_wire buffer_13334 (.in(n13334), .out(n13334_0));
mux15 mux_8169 (.in({n13419_1, n10337_1, n10327_0, n10310_0, n10304_0/**/, n10301_0, n10276_0, n10273_0, n10264_1, n10220_1, n4582, n4574, n3606, n3598, n3590}), .out(n13335), .config_in(config_chain[30129:30124]), .config_rst(config_rst)); 
buffer_wire buffer_13335 (.in(n13335), .out(n13335_0));
mux3 mux_8170 (.in({n9807_0, n9806_0, n3504}), .out(n13336), .config_in(config_chain[30131:30130]), .config_rst(config_rst)); 
buffer_wire buffer_13336 (.in(n13336), .out(n13336_0));
mux15 mux_8171 (.in({n13439_1, n10595_1, n10574_0, n10571_0, n10565_0, n10548_0, n10542_0, n10539_0, n10522_1, n10480_1, n4680, n4672, n3704, n3696, n3688}), .out(n13337), .config_in(config_chain[30137:30132]), .config_rst(config_rst)); 
buffer_wire buffer_13337 (.in(n13337), .out(n13337_0));
mux3 mux_8172 (.in({n9829_1, n9706_1/**/, n3508}), .out(n13338), .config_in(config_chain[30139:30138]), .config_rst(config_rst)); 
buffer_wire buffer_13338 (.in(n13338), .out(n13338_0));
mux14 mux_8173 (.in({n13461_1, n10855_1/**/, n10835_0, n10828_0, n10823_0, n10816_0, n10804_0, n10789_0, n10742_1, n4782, n4774, n4766, n3798, n3790}), .out(n13339), .config_in(config_chain[30145:30140]), .config_rst(config_rst)); 
buffer_wire buffer_13339 (.in(n13339), .out(n13339_0));
mux3 mux_8174 (.in({n9769_0/**/, n9768_0, n3508}), .out(n13340), .config_in(config_chain[30147:30146]), .config_rst(config_rst)); 
buffer_wire buffer_13340 (.in(n13340), .out(n13340_0));
mux15 mux_8175 (.in({n13401_1, n10079_1, n10062_0, n10059_0, n10051_0, n10034_0, n10028_0, n10025_0, n10010_1, n9970_1, n4488, n4480/**/, n4472, n3504, n3496}), .out(n13341), .config_in(config_chain[30153:30148]), .config_rst(config_rst)); 
buffer_wire buffer_13341 (.in(n13341), .out(n13341_0));
mux3 mux_8176 (.in({n9789_0, n9788_0, n3508}), .out(n13342), .config_in(config_chain[30155:30154]), .config_rst(config_rst)); 
buffer_wire buffer_13342 (.in(n13342), .out(n13342_0));
mux15 mux_8177 (.in({n13421_1, n10335_1, n10324_0, n10321_0, n10298_0, n10295_0, n10287_0, n10270_0, n10266_1, n10228_1, n4586, n4578, n4570, n3602, n3594}), .out(n13343), .config_in(config_chain[30161:30156]), .config_rst(config_rst)); 
buffer_wire buffer_13343 (.in(n13343), .out(n13343_0));
mux3 mux_8178 (.in({n9809_0/**/, n9808_0, n3508}), .out(n13344), .config_in(config_chain[30163:30162]), .config_rst(config_rst)); 
buffer_wire buffer_13344 (.in(n13344), .out(n13344_0));
mux15 mux_8179 (.in({n13441_1, n10593_1, n10585_0, n10568_0, n10562_0, n10559_0/**/, n10536_0, n10533_0, n10524_1, n10488_1, n4684, n4676, n4668, n3700, n3692}), .out(n13345), .config_in(config_chain[30169:30164]), .config_rst(config_rst)); 
buffer_wire buffer_13345 (.in(n13345), .out(n13345_0));
mux3 mux_8180 (.in({n9831_1, n9714_1, n3508}), .out(n13346), .config_in(config_chain[30171:30170]), .config_rst(config_rst)); 
buffer_wire buffer_13346 (.in(n13346), .out(n13346_0));
mux13 mux_8181 (.in({n13463_1, n10853_1, n10843_0/**/, n10836_0, n10824_0, n10809_0, n10797_0, n10790_0, n10750_1, n4774, n4766, n3798, n3790}), .out(n13347), .config_in(config_chain[30177:30172]), .config_rst(config_rst)); 
buffer_wire buffer_13347 (.in(n13347), .out(n13347_0));
mux3 mux_8182 (.in({n9771_0, n9770_0/**/, n4472}), .out(n13348), .config_in(config_chain[30179:30178]), .config_rst(config_rst)); 
buffer_wire buffer_13348 (.in(n13348), .out(n13348_0));
mux15 mux_8183 (.in({n13403_1, n10077_1, n10056_0, n10053_0, n10048_0, n10045_0, n10022_0, n10019_0, n10001_0, n9978_1, n4488, n4480, n4472, n3504, n3496/**/}), .out(n13349), .config_in(config_chain[30185:30180]), .config_rst(config_rst)); 
buffer_wire buffer_13349 (.in(n13349), .out(n13349_0));
mux3 mux_8184 (.in({n9791_0, n9790_0, n4472}), .out(n13350), .config_in(config_chain[30187:30186]), .config_rst(config_rst)); 
buffer_wire buffer_13350 (.in(n13350), .out(n13350_0));
mux15 mux_8185 (.in({n13423_1, n10333_1, n10318_0, n10315_0, n10292_0, n10289_0/**/, n10284_0, n10281_0, n10257_0, n10236_1, n4586, n4578, n4570, n3602, n3594}), .out(n13351), .config_in(config_chain[30193:30188]), .config_rst(config_rst)); 
buffer_wire buffer_13351 (.in(n13351), .out(n13351_0));
mux3 mux_8186 (.in({n9811_0/**/, n9810_0, n4472}), .out(n13352), .config_in(config_chain[30195:30194]), .config_rst(config_rst)); 
buffer_wire buffer_13352 (.in(n13352), .out(n13352_0));
mux15 mux_8187 (.in({n13443_1, n10591_1, n10582_0, n10579_0, n10556_0, n10553_0, n10530_0, n10527_0, n10515_0, n10496_1, n4684, n4676, n4668, n3700, n3692}), .out(n13353), .config_in(config_chain[30201:30196]), .config_rst(config_rst)); 
buffer_wire buffer_13353 (.in(n13353), .out(n13353_0));
mux3 mux_8188 (.in({n9833_1, n9722_1, n4472}), .out(n13354), .config_in(config_chain[30203:30202]), .config_rst(config_rst)); 
buffer_wire buffer_13354 (.in(n13354), .out(n13354_0));
mux13 mux_8189 (.in({n13465_1, n10851_1, n10844_0, n10829_0, n10817_0/**/, n10810_0, n10805_0, n10798_0, n10758_1, n4778, n4766, n3798, n3790}), .out(n13355), .config_in(config_chain[30209:30204]), .config_rst(config_rst)); 
buffer_wire buffer_13355 (.in(n13355), .out(n13355_0));
mux3 mux_8190 (.in({n9773_0, n9772_0, n4472}), .out(n13356), .config_in(config_chain[30211:30210]), .config_rst(config_rst)); 
buffer_wire buffer_13356 (.in(n13356), .out(n13356_0));
mux15 mux_8191 (.in({n13405_1, n10075_1, n10070_0, n10067_0, n10042_0, n10039_0, n10016_0, n10013_0, n10003_1, n9986_1/**/, n4488, n4480, n4472, n3504, n3496}), .out(n13357), .config_in(config_chain[30217:30212]), .config_rst(config_rst)); 
buffer_wire buffer_13357 (.in(n13357), .out(n13357_0));
mux3 mux_8192 (.in({n9793_0, n9792_0, n4476}), .out(n13358), .config_in(config_chain[30219:30218]), .config_rst(config_rst)); 
buffer_wire buffer_13358 (.in(n13358), .out(n13358_0));
mux15 mux_8193 (.in({n13425_1, n10331_1, n10312_0, n10309_0, n10306_0, n10303_0, n10278_0, n10275_0, n10259_0, n10244_1, n4586, n4578/**/, n4570, n3602, n3594}), .out(n13359), .config_in(config_chain[30225:30220]), .config_rst(config_rst)); 
buffer_wire buffer_13359 (.in(n13359), .out(n13359_0));
mux3 mux_8194 (.in({n9813_0, n9812_0, n4476}), .out(n13360), .config_in(config_chain[30227:30226]), .config_rst(config_rst)); 
buffer_wire buffer_13360 (.in(n13360), .out(n13360_0));
mux15 mux_8195 (.in({n13445_1, n10589_1, n10576_0, n10573_0, n10550_0, n10547_0, n10544_0, n10541_0/**/, n10517_0, n10504_1, n4684, n4676, n4668, n3700, n3692}), .out(n13361), .config_in(config_chain[30233:30228]), .config_rst(config_rst)); 
buffer_wire buffer_13361 (.in(n13361), .out(n13361_0));
mux3 mux_8196 (.in({n9835_1, n9730_1, n4476/**/}), .out(n13362), .config_in(config_chain[30235:30234]), .config_rst(config_rst)); 
buffer_wire buffer_13362 (.in(n13362), .out(n13362_0));
mux13 mux_8197 (.in({n13467_1, n10849_1, n10837_0, n10830_0, n10825_0, n10818_0, n10791_0, n10776_1, n10766_1/**/, n4778, n4770, n3798, n3790}), .out(n13363), .config_in(config_chain[30241:30236]), .config_rst(config_rst)); 
buffer_wire buffer_13363 (.in(n13363), .out(n13363_0));
mux3 mux_8198 (.in({n9775_0/**/, n9774_0, n4476}), .out(n13364), .config_in(config_chain[30243:30242]), .config_rst(config_rst)); 
buffer_wire buffer_13364 (.in(n13364), .out(n13364_0));
mux15 mux_8199 (.in({n13407_1, n10073_1, n10064_0, n10061_0, n10036_0, n10033_0, n10030_0, n10027_0, n10005_1, n9994_1, n4488, n4480, n4472, n3504, n3496}), .out(n13365), .config_in(config_chain[30249:30244]), .config_rst(config_rst)); 
buffer_wire buffer_13365 (.in(n13365), .out(n13365_0));
mux3 mux_8200 (.in({n9795_0, n9794_0/**/, n4476}), .out(n13366), .config_in(config_chain[30251:30250]), .config_rst(config_rst)); 
buffer_wire buffer_13366 (.in(n13366), .out(n13366_0));
mux15 mux_8201 (.in({n13427_1, n10329_1, n10326_0, n10323_0, n10300_0, n10297_0, n10272_0, n10269_0, n10261_1, n10252_1, n4586, n4578, n4570, n3602, n3594}), .out(n13367), .config_in(config_chain[30257:30252]), .config_rst(config_rst)); 
buffer_wire buffer_13367 (.in(n13367), .out(n13367_0));
mux3 mux_8202 (.in({n9815_0, n9814_0, n4480}), .out(n13368), .config_in(config_chain[30259:30258]), .config_rst(config_rst)); 
buffer_wire buffer_13368 (.in(n13368), .out(n13368_0));
mux15 mux_8203 (.in({n13447_1, n10587_1, n10570_0, n10567_0, n10564_0, n10561_0, n10538_0, n10535_0, n10519_0, n10512_1, n4684, n4676, n4668, n3700, n3692}), .out(n13369), .config_in(config_chain[30265:30260]), .config_rst(config_rst)); 
buffer_wire buffer_13369 (.in(n13369), .out(n13369_0));
mux3 mux_8204 (.in({n9837_1, n9738_1, n4480/**/}), .out(n13370), .config_in(config_chain[30267:30266]), .config_rst(config_rst)); 
buffer_wire buffer_13370 (.in(n13370), .out(n13370_0));
mux13 mux_8205 (.in({n13469_1, n10847_1, n10845_0, n10838_0, n10811_0, n10799_0/**/, n10792_0, n10778_1, n10774_1, n4778, n4770, n3802, n3790}), .out(n13371), .config_in(config_chain[30273:30268]), .config_rst(config_rst)); 
buffer_wire buffer_13371 (.in(n13371), .out(n13371_0));
mux3 mux_8206 (.in({n9777_0, n9776_0, n4480}), .out(n13372), .config_in(config_chain[30275:30274]), .config_rst(config_rst)); 
buffer_wire buffer_13372 (.in(n13372), .out(n13372_0));
mux15 mux_8207 (.in({n13409_1, n10091_1, n10058_0, n10055_0, n10050_0, n10047_0, n10024_0, n10021_0, n10007_1, n9922_1, n4488, n4480, n4472, n3504, n3496/**/}), .out(n13373), .config_in(config_chain[30281:30276]), .config_rst(config_rst)); 
buffer_wire buffer_13373 (.in(n13373), .out(n13373_0));
mux3 mux_8208 (.in({n9797_0, n9796_0, n4480/**/}), .out(n13374), .config_in(config_chain[30283:30282]), .config_rst(config_rst)); 
buffer_wire buffer_13374 (.in(n13374), .out(n13374_0));
mux15 mux_8209 (.in({n13429_1, n10347_1, n10320_0/**/, n10317_0, n10294_0, n10291_0, n10286_0, n10283_0, n10263_1, n10180_1, n4586, n4578, n4570, n3602, n3594}), .out(n13375), .config_in(config_chain[30289:30284]), .config_rst(config_rst)); 
buffer_wire buffer_13375 (.in(n13375), .out(n13375_0));
mux3 mux_8210 (.in({n9817_0, n9816_0, n4480}), .out(n13376), .config_in(config_chain[30291:30290]), .config_rst(config_rst)); 
buffer_wire buffer_13376 (.in(n13376), .out(n13376_0));
mux15 mux_8211 (.in({n13449_1, n10605_1, n10584_0, n10581_0, n10558_0, n10555_0, n10532_0, n10529_0/**/, n10521_1, n10440_1, n4684, n4676, n4668, n3700, n3692}), .out(n13377), .config_in(config_chain[30297:30292]), .config_rst(config_rst)); 
buffer_wire buffer_13377 (.in(n13377), .out(n13377_0));
mux3 mux_8212 (.in({n9747_1, n9746_1, n4484}), .out(n13378), .config_in(config_chain[30299:30298]), .config_rst(config_rst)); 
buffer_wire buffer_13378 (.in(n13378), .out(n13378_0));
mux13 mux_8213 (.in({n13471_1, n10867_1, n10831_0, n10819_0, n10812_0, n10800_0, n10780_1, n10777_0, n10694_1, n4778, n4770, n3802, n3794}), .out(n13379), .config_in(config_chain[30305:30300]), .config_rst(config_rst)); 
buffer_wire buffer_13379 (.in(n13379), .out(n13379_0));
mux3 mux_8214 (.in({n9749_1, n9748_1, n4484}), .out(n13380), .config_in(config_chain[30307:30306]), .config_rst(config_rst)); 
buffer_wire buffer_13380 (.in(n13380), .out(n13380_0));
mux13 mux_8215 (.in({n13493_1, n11131_1, n11109_1, n11102_0, n11073_0, n11061_0, n11054_0, n11042_1, n10958_1/**/, n4876, n4868, n3900, n3892}), .out(n13381), .config_in(config_chain[30313:30308]), .config_rst(config_rst)); 
buffer_wire buffer_13381 (.in(n13381), .out(n13381_0));
mux3 mux_8216 (.in({n9751_1, n9750_1, n4484}), .out(n13382), .config_in(config_chain[30315:30314]), .config_rst(config_rst)); 
buffer_wire buffer_13382 (.in(n13382), .out(n13382_0));
mux13 mux_8217 (.in({n13515_0, n11397_1, n11367_0, n11360_0, n11353_1, n11346_0, n11317_0, n11306_1, n11224_1, n4974, n4966, n3998, n3990}), .out(n13383), .config_in(config_chain[30321:30316]), .config_rst(config_rst)); 
buffer_wire buffer_13383 (.in(n13383), .out(n13383_0));
mux3 mux_8218 (.in({n9753_1/**/, n9752_1, n4484}), .out(n13384), .config_in(config_chain[30323:30322]), .config_rst(config_rst)); 
buffer_wire buffer_13384 (.in(n13384), .out(n13384_0));
mux13 mux_8219 (.in({n13537_0, n11663_1, n11640_0, n11625_0, n11611_0, n11604_0, n11597_1/**/, n11590_0, n11490_1, n5072, n5064, n4096, n4088}), .out(n13385), .config_in(config_chain[30329:30324]), .config_rst(config_rst)); 
buffer_wire buffer_13385 (.in(n13385), .out(n13385_0));
mux3 mux_8220 (.in({n9755_1/**/, n9754_1, n4484}), .out(n13386), .config_in(config_chain[30331:30330]), .config_rst(config_rst)); 
buffer_wire buffer_13386 (.in(n13386), .out(n13386_0));
mux13 mux_8221 (.in({n13559_0, n11927_1, n11889_0, n11882_0, n11875_0, n11868_0, n11854_0, n11829_1, n11748_1, n5170, n5162, n4194, n4186}), .out(n13387), .config_in(config_chain[30337:30332]), .config_rst(config_rst)); 
buffer_wire buffer_13387 (.in(n13387), .out(n13387_0));
mux3 mux_8222 (.in({n9757_1, n9756_1, n4488}), .out(n13388), .config_in(config_chain[30339:30338]), .config_rst(config_rst)); 
buffer_wire buffer_13388 (.in(n13388), .out(n13388_0));
mux3 mux_8223 (.in({n12189_1, n12100_1, n5272}), .out(n13389), .config_in(config_chain[30341:30340]), .config_rst(config_rst)); 
buffer_wire buffer_13389 (.in(n13389), .out(n13389_0));
mux16 mux_8224 (.in({n13300_0/**/, n10075_1, n10068_0, n10053_0, n10045_0, n10040_0, n10019_0, n10014_0, n10008_1, n10001_0, n9922_1, n4582, n4574, n3606, n3598, n3590}), .out(n13390), .config_in(config_chain[30347:30342]), .config_rst(config_rst)); 
buffer_wire buffer_13390 (.in(n13390), .out(n13390_0));
mux15 mux_8225 (.in({n13473_1, n11129_1, n11095_0, n11088_0/**/, n11081_0, n11074_0, n11062_0, n11044_1, n11041_0, n10966_1, n4876, n4868, n3900, n3892, n3884}), .out(n13391), .config_in(config_chain[30353:30348]), .config_rst(config_rst)); 
buffer_wire buffer_13391 (.in(n13391), .out(n13391_0));
mux16 mux_8226 (.in({n13308_0, n10077_1, n10067_0, n10062_0, n10039_0, n10034_0, n10028_0, n10013_0, n10010_1, n10003_1, n9994_1/**/, n4582, n4574, n3606, n3598, n3590}), .out(n13392), .config_in(config_chain[30359:30354]), .config_rst(config_rst)); 
buffer_wire buffer_13392 (.in(n13392), .out(n13392_0));
mux15 mux_8227 (.in({n13475_1, n11127_1, n11103_0/**/, n11096_0, n11082_0, n11055_0, n11048_0, n11046_1, n11043_0, n10974_1, n4880, n4868, n3900, n3892, n3884}), .out(n13393), .config_in(config_chain[30365:30360]), .config_rst(config_rst)); 
buffer_wire buffer_13393 (.in(n13393), .out(n13393_0));
mux15 mux_8228 (.in({n13316_0, n10079_1, n10061_0, n10056_0, n10048_0, n10033_0, n10027_0, n10022_0, n10005_1, n9986_1, n4582, n4574, n3606/**/, n3598, n3590}), .out(n13394), .config_in(config_chain[30371:30366]), .config_rst(config_rst)); 
buffer_wire buffer_13394 (.in(n13394), .out(n13394_0));
mux15 mux_8229 (.in({n13477_1/**/, n11125_1, n11104_0, n11089_0, n11075_0, n11068_0, n11063_0, n11056_0, n11045_0, n10982_1, n4880, n4872, n3900, n3892, n3884}), .out(n13395), .config_in(config_chain[30377:30372]), .config_rst(config_rst)); 
buffer_wire buffer_13395 (.in(n13395), .out(n13395_0));
mux15 mux_8230 (.in({n13324_0, n10081_1, n10070_0, n10055_0, n10047_0, n10042_0, n10021_0, n10016_0, n10007_1, n9978_1, n4582, n4574, n3606, n3598, n3590/**/}), .out(n13396), .config_in(config_chain[30383:30378]), .config_rst(config_rst)); 
buffer_wire buffer_13396 (.in(n13396), .out(n13396_0));
mux15 mux_8231 (.in({n13479_1, n11123_1, n11097_0, n11090_0, n11083_0, n11076_0, n11064_0, n11049_0, n11047_1, n10990_1, n4880, n4872, n4864, n3892, n3884/**/}), .out(n13397), .config_in(config_chain[30389:30384]), .config_rst(config_rst)); 
buffer_wire buffer_13397 (.in(n13397), .out(n13397_0));
mux15 mux_8232 (.in({n13332_0, n10083_1, n10069_0/**/, n10064_0, n10041_0, n10036_0, n10030_0, n10015_0, n10009_1, n9970_1, n4582, n4574, n3606, n3598, n3590}), .out(n13398), .config_in(config_chain[30395:30390]), .config_rst(config_rst)); 
buffer_wire buffer_13398 (.in(n13398), .out(n13398_0));
mux14 mux_8233 (.in({n13481_1, n11121_1/**/, n11105_0, n11098_0, n11084_0, n11069_0, n11057_0, n11050_0, n10998_1, n4880, n4872, n4864, n3896, n3884}), .out(n13399), .config_in(config_chain[30401:30396]), .config_rst(config_rst)); 
buffer_wire buffer_13399 (.in(n13399), .out(n13399_0));
mux15 mux_8234 (.in({n13340_0/**/, n10085_1, n10063_0, n10058_0, n10050_0, n10035_0, n10029_0, n10024_0, n10011_1, n9962_1, n4586, n4578, n4570, n3602, n3594}), .out(n13400), .config_in(config_chain[30407:30402]), .config_rst(config_rst)); 
buffer_wire buffer_13400 (.in(n13400), .out(n13400_0));
mux14 mux_8235 (.in({n13483_1, n11119_1, n11106_0, n11091_0, n11077_0, n11070_0, n11065_0, n11058_0, n11006_1, n4880/**/, n4872, n4864, n3896, n3888}), .out(n13401), .config_in(config_chain[30413:30408]), .config_rst(config_rst)); 
buffer_wire buffer_13401 (.in(n13401), .out(n13401_0));
mux15 mux_8236 (.in({n13348_0/**/, n10087_1, n10057_0, n10052_0, n10049_0, n10044_0, n10023_0, n10018_0, n10000_1, n9954_1, n4586, n4578, n4570, n3602, n3594}), .out(n13402), .config_in(config_chain[30419:30414]), .config_rst(config_rst)); 
buffer_wire buffer_13402 (.in(n13402), .out(n13402_0));
mux13 mux_8237 (.in({n13485_1, n11117_1, n11099_0, n11092_0, n11085_0, n11078_0, n11066_0/**/, n11051_0, n11014_1, n4872, n4864, n3896, n3888}), .out(n13403), .config_in(config_chain[30425:30420]), .config_rst(config_rst)); 
buffer_wire buffer_13403 (.in(n13403), .out(n13403_0));
mux15 mux_8238 (.in({n13356_0, n10089_1, n10071_0, n10066_0, n10043_0, n10038_0, n10017_0, n10012_0, n10002_1, n9946_1/**/, n4586, n4578, n4570, n3602, n3594}), .out(n13404), .config_in(config_chain[30431:30426]), .config_rst(config_rst)); 
buffer_wire buffer_13404 (.in(n13404), .out(n13404_0));
mux13 mux_8239 (.in({n13487_1, n11115_1, n11107_0, n11100_0, n11086_0, n11071_0, n11059_0, n11052_0/**/, n11022_1, n4876, n4864, n3896, n3888}), .out(n13405), .config_in(config_chain[30437:30432]), .config_rst(config_rst)); 
buffer_wire buffer_13405 (.in(n13405), .out(n13405_0));
mux15 mux_8240 (.in({n13364_0/**/, n10091_1, n10065_0, n10060_0, n10037_0, n10032_0, n10031_0, n10026_0, n10004_1, n9938_1, n4586, n4578, n4570, n3602, n3594}), .out(n13406), .config_in(config_chain[30443:30438]), .config_rst(config_rst)); 
buffer_wire buffer_13406 (.in(n13406), .out(n13406_0));
mux13 mux_8241 (.in({n13489_1, n11113_1, n11108_0, n11093_0, n11079_0, n11072_0, n11067_0, n11060_0/**/, n11030_1, n4876, n4868, n3896, n3888}), .out(n13407), .config_in(config_chain[30449:30444]), .config_rst(config_rst)); 
buffer_wire buffer_13407 (.in(n13407), .out(n13407_0));
mux15 mux_8242 (.in({n13372_0, n10073_1, n10059_0, n10054_0, n10051_0, n10046_0, n10025_0, n10020_0, n10006_1, n9930_1, n4586/**/, n4578, n4570, n3602, n3594}), .out(n13408), .config_in(config_chain[30455:30450]), .config_rst(config_rst)); 
buffer_wire buffer_13408 (.in(n13408), .out(n13408_0));
mux13 mux_8243 (.in({n13491_1, n11111_1, n11101_0, n11094_0, n11087_0/**/, n11080_0, n11053_0, n11040_1, n11038_1, n4876, n4868, n3900, n3888}), .out(n13409), .config_in(config_chain[30461:30456]), .config_rst(config_rst)); 
buffer_wire buffer_13409 (.in(n13409), .out(n13409_0));
mux16 mux_8244 (.in({n13302_0, n10331_1, n10315_0, n10310_0, n10304_0, n10289_0, n10281_0, n10276_0, n10264_1, n10257_0, n10180_1, n4680, n4672, n3704, n3696, n3688/**/}), .out(n13410), .config_in(config_chain[30467:30462]), .config_rst(config_rst)); 
buffer_wire buffer_13410 (.in(n13410), .out(n13410_0));
mux15 mux_8245 (.in({n13495_0, n11395_1, n11375_1, n11368_0, n11339_0, n11332_0, n11325_0, n11318_0, n11308_1, n11232_1, n4974/**/, n4966, n3998, n3990, n3982}), .out(n13411), .config_in(config_chain[30473:30468]), .config_rst(config_rst)); 
buffer_wire buffer_13411 (.in(n13411), .out(n13411_0));
mux16 mux_8246 (.in({n13310_0, n10333_1, n10324_0, n10309_0, n10303_0, n10298_0, n10275_0, n10270_0, n10266_1, n10259_0, n10252_1, n4680, n4672, n3704, n3696, n3688/**/}), .out(n13412), .config_in(config_chain[30479:30474]), .config_rst(config_rst)); 
buffer_wire buffer_13412 (.in(n13412), .out(n13412_0));
mux15 mux_8247 (.in({n13497_0, n11393_1, n11361_0, n11354_0, n11347_0, n11340_0/**/, n11326_0, n11310_1, n11307_0, n11240_1, n4978, n4966, n3998, n3990, n3982}), .out(n13413), .config_in(config_chain[30485:30480]), .config_rst(config_rst)); 
buffer_wire buffer_13413 (.in(n13413), .out(n13413_0));
mux15 mux_8248 (.in({n13318_0, n10335_1, n10323_0, n10318_0, n10297_0, n10292_0, n10284_0/**/, n10269_0, n10261_1, n10244_1, n4680, n4672, n3704, n3696, n3688}), .out(n13414), .config_in(config_chain[30491:30486]), .config_rst(config_rst)); 
buffer_wire buffer_13414 (.in(n13414), .out(n13414_0));
mux15 mux_8249 (.in({n13499_0, n11391_1, n11369_0, n11362_0, n11348_0, n11333_0, n11319_0, n11312_0, n11309_0, n11248_1/**/, n4978, n4970, n3998, n3990, n3982}), .out(n13415), .config_in(config_chain[30497:30492]), .config_rst(config_rst)); 
buffer_wire buffer_13415 (.in(n13415), .out(n13415_0));
mux15 mux_8250 (.in({n13326_0, n10337_1, n10317_0, n10312_0, n10306_0, n10291_0, n10283_0, n10278_0, n10263_1, n10236_1/**/, n4680, n4672, n3704, n3696, n3688}), .out(n13416), .config_in(config_chain[30503:30498]), .config_rst(config_rst)); 
buffer_wire buffer_13416 (.in(n13416), .out(n13416_0));
mux15 mux_8251 (.in({n13501_0, n11389_1, n11370_0, n11355_0, n11341_0, n11334_0, n11327_0, n11320_0, n11311_0, n11256_1/**/, n4978, n4970, n4962, n3990, n3982}), .out(n13417), .config_in(config_chain[30509:30504]), .config_rst(config_rst)); 
buffer_wire buffer_13417 (.in(n13417), .out(n13417_0));
mux15 mux_8252 (.in({n13334_0, n10339_1/**/, n10326_0, n10311_0, n10305_0, n10300_0, n10277_0, n10272_0, n10265_1, n10228_1, n4680, n4672, n3704, n3696, n3688}), .out(n13418), .config_in(config_chain[30515:30510]), .config_rst(config_rst)); 
buffer_wire buffer_13418 (.in(n13418), .out(n13418_0));
mux14 mux_8253 (.in({n13503_0, n11387_1, n11363_0, n11356_0, n11349_0, n11342_0, n11328_0, n11313_0, n11264_1, n4978, n4970, n4962, n3994, n3982}), .out(n13419), .config_in(config_chain[30521:30516]), .config_rst(config_rst)); 
buffer_wire buffer_13419 (.in(n13419), .out(n13419_0));
mux15 mux_8254 (.in({n13342_0, n10341_1, n10325_0, n10320_0, n10299_0, n10294_0, n10286_0, n10271_0, n10267_1, n10220_1, n4684, n4676, n4668/**/, n3700, n3692}), .out(n13420), .config_in(config_chain[30527:30522]), .config_rst(config_rst)); 
buffer_wire buffer_13420 (.in(n13420), .out(n13420_0));
mux14 mux_8255 (.in({n13505_0, n11385_1, n11371_0, n11364_0, n11350_0/**/, n11335_0, n11321_0, n11314_0, n11272_1, n4978, n4970, n4962, n3994, n3986}), .out(n13421), .config_in(config_chain[30533:30528]), .config_rst(config_rst)); 
buffer_wire buffer_13421 (.in(n13421), .out(n13421_0));
mux15 mux_8256 (.in({n13350_0, n10343_1, n10319_0, n10314_0, n10293_0, n10288_0, n10285_0, n10280_0, n10256_1, n10212_1, n4684, n4676, n4668/**/, n3700, n3692}), .out(n13422), .config_in(config_chain[30539:30534]), .config_rst(config_rst)); 
buffer_wire buffer_13422 (.in(n13422), .out(n13422_0));
mux13 mux_8257 (.in({n13507_0, n11383_1/**/, n11372_0, n11357_0, n11343_0, n11336_0, n11329_0, n11322_0, n11280_1, n4970, n4962, n3994, n3986}), .out(n13423), .config_in(config_chain[30545:30540]), .config_rst(config_rst)); 
buffer_wire buffer_13423 (.in(n13423), .out(n13423_0));
mux15 mux_8258 (.in({n13358_0, n10345_1, n10313_0, n10308_0, n10307_0, n10302_0, n10279_0/**/, n10274_0, n10258_1, n10204_1, n4684, n4676, n4668, n3700, n3692}), .out(n13424), .config_in(config_chain[30551:30546]), .config_rst(config_rst)); 
buffer_wire buffer_13424 (.in(n13424), .out(n13424_0));
mux13 mux_8259 (.in({n13509_0/**/, n11381_1, n11365_0, n11358_0, n11351_0, n11344_0, n11330_0, n11315_0, n11288_1, n4974, n4962, n3994, n3986}), .out(n13425), .config_in(config_chain[30557:30552]), .config_rst(config_rst)); 
buffer_wire buffer_13425 (.in(n13425), .out(n13425_0));
mux15 mux_8260 (.in({n13366_0, n10347_1, n10327_0, n10322_0, n10301_0/**/, n10296_0, n10273_0, n10268_0, n10260_1, n10196_1, n4684, n4676, n4668, n3700, n3692}), .out(n13426), .config_in(config_chain[30563:30558]), .config_rst(config_rst)); 
buffer_wire buffer_13426 (.in(n13426), .out(n13426_0));
mux13 mux_8261 (.in({n13511_0, n11379_1, n11373_0, n11366_0, n11352_0, n11337_0, n11323_0, n11316_0, n11296_1, n4974, n4966, n3994, n3986}), .out(n13427), .config_in(config_chain[30569:30564]), .config_rst(config_rst)); 
buffer_wire buffer_13427 (.in(n13427), .out(n13427_0));
mux15 mux_8262 (.in({n13374_0, n10329_1, n10321_0, n10316_0, n10295_0, n10290_0, n10287_0, n10282_0, n10262_1, n10188_1, n4684/**/, n4676, n4668, n3700, n3692}), .out(n13428), .config_in(config_chain[30575:30570]), .config_rst(config_rst)); 
buffer_wire buffer_13428 (.in(n13428), .out(n13428_0));
mux13 mux_8263 (.in({n13513_0, n11377_1, n11374_0, n11359_0, n11345_0, n11338_0, n11331_0, n11324_0, n11304_1, n4974/**/, n4966, n3998, n3986}), .out(n13429), .config_in(config_chain[30581:30576]), .config_rst(config_rst)); 
buffer_wire buffer_13429 (.in(n13429), .out(n13429_0));
mux16 mux_8264 (.in({n13304_0, n10589_1/**/, n10579_0, n10574_0, n10553_0, n10548_0, n10542_0, n10527_0, n10522_1, n10515_0, n10440_1, n4778, n4770, n3802, n3794, n3786}), .out(n13430), .config_in(config_chain[30587:30582]), .config_rst(config_rst)); 
buffer_wire buffer_13430 (.in(n13430), .out(n13430_0));
mux15 mux_8265 (.in({n13517_0, n11661_1, n11633_0, n11626_0/**/, n11619_1, n11612_0, n11583_0, n11576_0, n11572_1, n11498_1, n5072, n5064, n4096, n4088, n4080}), .out(n13431), .config_in(config_chain[30593:30588]), .config_rst(config_rst)); 
buffer_wire buffer_13431 (.in(n13431), .out(n13431_0));
mux16 mux_8266 (.in({n13312_0, n10591_1, n10573_0, n10568_0, n10562_0, n10547_0, n10541_0/**/, n10536_0, n10524_1, n10517_0, n10512_1, n4778, n4770, n3802, n3794, n3786}), .out(n13432), .config_in(config_chain[30599:30594]), .config_rst(config_rst)); 
buffer_wire buffer_13432 (.in(n13432), .out(n13432_0));
mux15 mux_8267 (.in({n13519_0/**/, n11659_1, n11641_1, n11634_0, n11605_0, n11598_0, n11591_0, n11584_0, n11574_1, n11506_1, n5076, n5064, n4096, n4088, n4080}), .out(n13433), .config_in(config_chain[30605:30600]), .config_rst(config_rst)); 
buffer_wire buffer_13433 (.in(n13433), .out(n13433_0));
mux15 mux_8268 (.in({n13320_0, n10593_1, n10582_0, n10567_0/**/, n10561_0, n10556_0, n10535_0, n10530_0, n10519_0, n10504_1, n4778, n4770, n3802, n3794, n3786}), .out(n13434), .config_in(config_chain[30611:30606]), .config_rst(config_rst)); 
buffer_wire buffer_13434 (.in(n13434), .out(n13434_0));
mux15 mux_8269 (.in({n13521_0, n11657_1, n11627_0, n11620_0, n11613_0, n11606_0, n11592_0, n11577_0, n11573_0, n11514_1, n5076, n5068/**/, n4096, n4088, n4080}), .out(n13435), .config_in(config_chain[30617:30612]), .config_rst(config_rst)); 
buffer_wire buffer_13435 (.in(n13435), .out(n13435_0));
mux15 mux_8270 (.in({n13328_0, n10595_1, n10581_0, n10576_0, n10555_0, n10550_0, n10544_0, n10529_0, n10521_1, n10496_1, n4778, n4770, n3802, n3794, n3786}), .out(n13436), .config_in(config_chain[30623:30618]), .config_rst(config_rst)); 
buffer_wire buffer_13436 (.in(n13436), .out(n13436_0));
mux15 mux_8271 (.in({n13523_0, n11655_1, n11635_0, n11628_0, n11614_0, n11599_0, n11585_0, n11578_0, n11575_0, n11522_1, n5076/**/, n5068, n5060, n4088, n4080}), .out(n13437), .config_in(config_chain[30629:30624]), .config_rst(config_rst)); 
buffer_wire buffer_13437 (.in(n13437), .out(n13437_0));
mux15 mux_8272 (.in({n13336_0, n10597_1, n10575_0, n10570_0, n10564_0/**/, n10549_0, n10543_0, n10538_0, n10523_1, n10488_1, n4778, n4770, n3802, n3794, n3786}), .out(n13438), .config_in(config_chain[30635:30630]), .config_rst(config_rst)); 
buffer_wire buffer_13438 (.in(n13438), .out(n13438_0));
mux14 mux_8273 (.in({n13525_0, n11653_1, n11636_0, n11621_0, n11607_0, n11600_0, n11593_0, n11586_0, n11530_1, n5076, n5068/**/, n5060, n4092, n4080}), .out(n13439), .config_in(config_chain[30641:30636]), .config_rst(config_rst)); 
buffer_wire buffer_13439 (.in(n13439), .out(n13439_0));
mux15 mux_8274 (.in({n13344_0, n10599_1, n10584_0, n10569_0, n10563_0, n10558_0, n10537_0, n10532_0, n10525_1, n10480_1, n4782, n4774, n4766/**/, n3798, n3790}), .out(n13440), .config_in(config_chain[30647:30642]), .config_rst(config_rst)); 
buffer_wire buffer_13440 (.in(n13440), .out(n13440_0));
mux14 mux_8275 (.in({n13527_0, n11651_1, n11629_0, n11622_0, n11615_0, n11608_0, n11594_0, n11579_0, n11538_1, n5076, n5068, n5060, n4092, n4084/**/}), .out(n13441), .config_in(config_chain[30653:30648]), .config_rst(config_rst)); 
buffer_wire buffer_13441 (.in(n13441), .out(n13441_0));
mux15 mux_8276 (.in({n13352_0, n10601_1, n10583_0, n10578_0, n10557_0, n10552_0, n10531_0/**/, n10526_0, n10514_1, n10472_1, n4782, n4774, n4766, n3798, n3790}), .out(n13442), .config_in(config_chain[30659:30654]), .config_rst(config_rst)); 
buffer_wire buffer_13442 (.in(n13442), .out(n13442_0));
mux13 mux_8277 (.in({n13529_0, n11649_1, n11637_0, n11630_0, n11616_0, n11601_0, n11587_0, n11580_0, n11546_1, n5068, n5060, n4092, n4084/**/}), .out(n13443), .config_in(config_chain[30665:30660]), .config_rst(config_rst)); 
buffer_wire buffer_13443 (.in(n13443), .out(n13443_0));
mux15 mux_8278 (.in({n13360_0, n10603_1, n10577_0/**/, n10572_0, n10551_0, n10546_0, n10545_0, n10540_0, n10516_1, n10464_1, n4782, n4774, n4766, n3798, n3790}), .out(n13444), .config_in(config_chain[30671:30666]), .config_rst(config_rst)); 
buffer_wire buffer_13444 (.in(n13444), .out(n13444_0));
mux13 mux_8279 (.in({n13531_0, n11647_1, n11638_0, n11623_0, n11609_0, n11602_0, n11595_0, n11588_0/**/, n11554_1, n5072, n5060, n4092, n4084}), .out(n13445), .config_in(config_chain[30677:30672]), .config_rst(config_rst)); 
buffer_wire buffer_13445 (.in(n13445), .out(n13445_0));
mux15 mux_8280 (.in({n13368_0, n10605_1, n10571_0, n10566_0, n10565_0, n10560_0, n10539_0, n10534_0, n10518_1, n10456_1, n4782/**/, n4774, n4766, n3798, n3790}), .out(n13446), .config_in(config_chain[30683:30678]), .config_rst(config_rst)); 
buffer_wire buffer_13446 (.in(n13446), .out(n13446_0));
mux13 mux_8281 (.in({n13533_0, n11645_1, n11631_0, n11624_0, n11617_0, n11610_0, n11596_0, n11581_0, n11562_1/**/, n5072, n5064, n4092, n4084}), .out(n13447), .config_in(config_chain[30689:30684]), .config_rst(config_rst)); 
buffer_wire buffer_13447 (.in(n13447), .out(n13447_0));
mux15 mux_8282 (.in({n13376_0, n10587_1, n10585_0, n10580_0, n10559_0, n10554_0, n10533_0, n10528_0, n10520_1, n10448_1, n4782, n4774, n4766, n3798/**/, n3790}), .out(n13448), .config_in(config_chain[30695:30690]), .config_rst(config_rst)); 
buffer_wire buffer_13448 (.in(n13448), .out(n13448_0));
mux13 mux_8283 (.in({n13535_0, n11643_1/**/, n11639_0, n11632_0, n11618_0, n11603_0, n11589_0, n11582_0, n11570_1, n5072, n5064, n4096, n4084}), .out(n13449), .config_in(config_chain[30701:30696]), .config_rst(config_rst)); 
buffer_wire buffer_13449 (.in(n13449), .out(n13449_0));
mux15 mux_8284 (.in({n13298_1, n10849_1/**/, n10838_0, n10833_0, n10821_0, n10792_0, n10787_0, n10783_1, n10778_1, n10694_1, n4876, n4868, n3900, n3892, n3884}), .out(n13450), .config_in(config_chain[30707:30702]), .config_rst(config_rst)); 
buffer_wire buffer_13450 (.in(n13450), .out(n13450_0));
mux15 mux_8285 (.in({n13539_0, n11925_1, n11904_0, n11897_0, n11890_0, n11876_0, n11861_1, n11847_0, n11840_0/**/, n11756_1, n5170, n5162, n4194, n4186, n4178}), .out(n13451), .config_in(config_chain[30713:30708]), .config_rst(config_rst)); 
buffer_wire buffer_13451 (.in(n13451), .out(n13451_0));
mux15 mux_8286 (.in({n13306_1, n10851_1, n10841_0, n10812_0, n10807_0, n10800_0, n10795_0/**/, n10785_1, n10780_1, n10774_1, n4880, n4868, n3900, n3892, n3884}), .out(n13452), .config_in(config_chain[30719:30714]), .config_rst(config_rst)); 
buffer_wire buffer_13452 (.in(n13452), .out(n13452_0));
mux15 mux_8287 (.in({n13541_0, n11923_1/**/, n11898_0, n11883_1, n11869_0, n11862_0, n11855_0, n11848_0, n11838_1, n11764_1, n5174, n5162, n4194, n4186, n4178}), .out(n13453), .config_in(config_chain[30725:30720]), .config_rst(config_rst)); 
buffer_wire buffer_13453 (.in(n13453), .out(n13453_0));
mux15 mux_8288 (.in({n13314_1/**/, n10853_1, n10832_0, n10827_0, n10820_0, n10815_0, n10803_0, n10786_0, n10782_1, n10766_1, n4880, n4872, n3900, n3892, n3884}), .out(n13454), .config_in(config_chain[30731:30726]), .config_rst(config_rst)); 
buffer_wire buffer_13454 (.in(n13454), .out(n13454_0));
mux15 mux_8289 (.in({n13543_0, n11921_1, n11905_1, n11891_0, n11884_0, n11877_0, n11870_0, n11856_0, n11841_0, n11772_1/**/, n5174, n5166, n4194, n4186, n4178}), .out(n13455), .config_in(config_chain[30737:30732]), .config_rst(config_rst)); 
buffer_wire buffer_13455 (.in(n13455), .out(n13455_0));
mux15 mux_8290 (.in({n13322_1, n10855_1, n10840_0, n10835_0/**/, n10823_0, n10806_0, n10794_0, n10789_0, n10784_1, n10758_1, n4880, n4872, n4864, n3892, n3884}), .out(n13456), .config_in(config_chain[30743:30738]), .config_rst(config_rst)); 
buffer_wire buffer_13456 (.in(n13456), .out(n13456_0));
mux15 mux_8291 (.in({n13545_0, n11919_1, n11899_0, n11892_0, n11878_0/**/, n11863_0, n11849_0, n11842_0, n11839_0, n11780_1, n5174, n5166, n5158, n4186, n4178}), .out(n13457), .config_in(config_chain[30749:30744]), .config_rst(config_rst)); 
buffer_wire buffer_13457 (.in(n13457), .out(n13457_0));
mux14 mux_8292 (.in({n13330_1, n10857_1, n10843_0, n10826_0, n10814_0, n10809_0, n10802_0, n10797_0, n10750_1, n4880, n4872, n4864, n3896, n3884}), .out(n13458), .config_in(config_chain[30755:30750]), .config_rst(config_rst)); 
buffer_wire buffer_13458 (.in(n13458), .out(n13458_0));
mux14 mux_8293 (.in({n13547_0, n11917_1, n11900_0, n11885_0, n11871_0, n11864_0, n11857_0, n11850_0, n11788_1/**/, n5174, n5166, n5158, n4190, n4178}), .out(n13459), .config_in(config_chain[30761:30756]), .config_rst(config_rst)); 
buffer_wire buffer_13459 (.in(n13459), .out(n13459_0));
mux14 mux_8294 (.in({n13338_1/**/, n10859_1, n10834_0, n10829_0, n10822_0, n10817_0, n10805_0, n10788_0, n10742_1, n4880, n4872, n4864, n3896, n3888}), .out(n13460), .config_in(config_chain[30767:30762]), .config_rst(config_rst)); 
buffer_wire buffer_13460 (.in(n13460), .out(n13460_0));
mux14 mux_8295 (.in({n13549_0, n11915_1, n11893_0, n11886_0, n11879_0, n11872_0, n11858_0, n11843_0, n11796_1/**/, n5174, n5166, n5158, n4190, n4182}), .out(n13461), .config_in(config_chain[30773:30768]), .config_rst(config_rst)); 
buffer_wire buffer_13461 (.in(n13461), .out(n13461_0));
mux13 mux_8296 (.in({n13346_1, n10861_1, n10842_0, n10837_0, n10825_0, n10808_0, n10796_0/**/, n10791_0, n10734_1, n4872, n4864, n3896, n3888}), .out(n13462), .config_in(config_chain[30779:30774]), .config_rst(config_rst)); 
buffer_wire buffer_13462 (.in(n13462), .out(n13462_0));
mux13 mux_8297 (.in({n13551_0, n11913_1, n11901_0, n11894_0/**/, n11880_0, n11865_0, n11851_0, n11844_0, n11804_1, n5166, n5158, n4190, n4182}), .out(n13463), .config_in(config_chain[30785:30780]), .config_rst(config_rst)); 
buffer_wire buffer_13463 (.in(n13463), .out(n13463_0));
mux13 mux_8298 (.in({n13354_1, n10863_1, n10845_0, n10828_0, n10816_0, n10811_0, n10804_0, n10799_0, n10726_1/**/, n4876, n4864, n3896, n3888}), .out(n13464), .config_in(config_chain[30791:30786]), .config_rst(config_rst)); 
buffer_wire buffer_13464 (.in(n13464), .out(n13464_0));
mux13 mux_8299 (.in({n13553_0, n11911_1, n11902_0, n11887_0, n11873_0, n11866_0, n11859_0, n11852_0/**/, n11812_1, n5170, n5158, n4190, n4182}), .out(n13465), .config_in(config_chain[30797:30792]), .config_rst(config_rst)); 
buffer_wire buffer_13465 (.in(n13465), .out(n13465_0));
mux13 mux_8300 (.in({n13362_1/**/, n10865_1, n10836_0, n10831_0, n10824_0, n10819_0, n10790_0, n10777_0, n10718_1, n4876, n4868, n3896, n3888}), .out(n13466), .config_in(config_chain[30803:30798]), .config_rst(config_rst)); 
buffer_wire buffer_13466 (.in(n13466), .out(n13466_0));
mux13 mux_8301 (.in({n13555_0, n11909_1, n11895_0, n11888_0, n11881_0, n11874_0, n11845_0, n11828_1, n11820_1, n5170, n5162, n4190/**/, n4182}), .out(n13467), .config_in(config_chain[30809:30804]), .config_rst(config_rst)); 
buffer_wire buffer_13467 (.in(n13467), .out(n13467_0));
mux13 mux_8302 (.in({n13370_1/**/, n10867_1, n10844_0, n10839_0, n10810_0, n10798_0, n10793_0, n10779_0, n10710_1, n4876, n4868, n3900, n3888}), .out(n13468), .config_in(config_chain[30815:30810]), .config_rst(config_rst)); 
buffer_wire buffer_13468 (.in(n13468), .out(n13468_0));
mux13 mux_8303 (.in({n13557_0, n11907_1, n11903_0, n11896_0, n11867_0, n11860_0, n11853_0/**/, n11846_0, n11836_1, n5170, n5162, n4194, n4182}), .out(n13469), .config_in(config_chain[30821:30816]), .config_rst(config_rst)); 
buffer_wire buffer_13469 (.in(n13469), .out(n13469_0));
mux13 mux_8304 (.in({n13378_1, n10847_1, n10830_0, n10818_0, n10813_0, n10801_0/**/, n10781_0, n10776_1, n10702_1, n4876, n4868, n3900, n3892}), .out(n13470), .config_in(config_chain[30827:30822]), .config_rst(config_rst)); 
buffer_wire buffer_13470 (.in(n13470), .out(n13470_0));
mux3 mux_8305 (.in({n12091_1, n12090_1/**/, n5268}), .out(n13471), .config_in(config_chain[30829:30828]), .config_rst(config_rst)); 
buffer_wire buffer_13471 (.in(n13471), .out(n13471_0));
mux15 mux_8306 (.in({n13390_1, n11113_1, n11094_0, n11089_0, n11080_0, n11075_0, n11063_0, n11045_0, n11040_1, n10958_1, n4974, n4966, n3998, n3990, n3982/**/}), .out(n13472), .config_in(config_chain[30835:30830]), .config_rst(config_rst)); 
buffer_wire buffer_13472 (.in(n13472), .out(n13472_0));
mux4 mux_8307 (.in({n12169_1/**/, n12012_1, n5272, n4276}), .out(n13473), .config_in(config_chain[30837:30836]), .config_rst(config_rst)); 
buffer_wire buffer_13473 (.in(n13473), .out(n13473_0));
mux15 mux_8308 (.in({n13392_1, n11115_1/**/, n11102_0, n11097_0, n11083_0, n11054_0, n11049_0, n11047_1, n11042_1, n11038_1, n4978, n4966, n3998, n3990, n3982}), .out(n13474), .config_in(config_chain[30843:30838]), .config_rst(config_rst)); 
buffer_wire buffer_13474 (.in(n13474), .out(n13474_0));
mux3 mux_8309 (.in({n12171_1, n12020_1, n4280}), .out(n13475), .config_in(config_chain[30845:30844]), .config_rst(config_rst)); 
buffer_wire buffer_13475 (.in(n13475), .out(n13475_0));
mux15 mux_8310 (.in({n13394_1, n11117_1, n11105_0, n11088_0, n11074_0, n11069_0, n11062_0, n11057_0, n11044_1, n11030_1, n4978/**/, n4970, n3998, n3990, n3982}), .out(n13476), .config_in(config_chain[30851:30846]), .config_rst(config_rst)); 
buffer_wire buffer_13476 (.in(n13476), .out(n13476_0));
mux3 mux_8311 (.in({n12173_1/**/, n12028_1, n4280}), .out(n13477), .config_in(config_chain[30853:30852]), .config_rst(config_rst)); 
buffer_wire buffer_13477 (.in(n13477), .out(n13477_0));
mux15 mux_8312 (.in({n13396_1, n11119_1, n11096_0, n11091_0, n11082_0, n11077_0, n11065_0, n11048_0, n11046_1, n11022_1, n4978, n4970/**/, n4962, n3990, n3982}), .out(n13478), .config_in(config_chain[30859:30854]), .config_rst(config_rst)); 
buffer_wire buffer_13478 (.in(n13478), .out(n13478_0));
mux3 mux_8313 (.in({n12175_1, n12036_1, n4284}), .out(n13479), .config_in(config_chain[30861:30860]), .config_rst(config_rst)); 
buffer_wire buffer_13479 (.in(n13479), .out(n13479_0));
mux14 mux_8314 (.in({n13398_1, n11121_1, n11104_0, n11099_0, n11085_0, n11068_0, n11056_0, n11051_0/**/, n11014_1, n4978, n4970, n4962, n3994, n3982}), .out(n13480), .config_in(config_chain[30867:30862]), .config_rst(config_rst)); 
buffer_wire buffer_13480 (.in(n13480), .out(n13480_0));
mux3 mux_8315 (.in({n12177_1/**/, n12044_1, n4288}), .out(n13481), .config_in(config_chain[30869:30868]), .config_rst(config_rst)); 
buffer_wire buffer_13481 (.in(n13481), .out(n13481_0));
mux14 mux_8316 (.in({n13400_1, n11123_1, n11107_0, n11090_0, n11076_0, n11071_0, n11064_0, n11059_0, n11006_1, n4978, n4970, n4962, n3994, n3986/**/}), .out(n13482), .config_in(config_chain[30875:30870]), .config_rst(config_rst)); 
buffer_wire buffer_13482 (.in(n13482), .out(n13482_0));
mux3 mux_8317 (.in({n12179_1, n12052_1/**/, n4292}), .out(n13483), .config_in(config_chain[30877:30876]), .config_rst(config_rst)); 
buffer_wire buffer_13483 (.in(n13483), .out(n13483_0));
mux13 mux_8318 (.in({n13402_1, n11125_1, n11098_0, n11093_0, n11084_0/**/, n11079_0, n11067_0, n11050_0, n10998_1, n4970, n4962, n3994, n3986}), .out(n13484), .config_in(config_chain[30883:30878]), .config_rst(config_rst)); 
buffer_wire buffer_13484 (.in(n13484), .out(n13484_0));
mux3 mux_8319 (.in({n12181_1/**/, n12060_1, n5256}), .out(n13485), .config_in(config_chain[30885:30884]), .config_rst(config_rst)); 
buffer_wire buffer_13485 (.in(n13485), .out(n13485_0));
mux13 mux_8320 (.in({n13404_1, n11127_1, n11106_0/**/, n11101_0, n11087_0, n11070_0, n11058_0, n11053_0, n10990_1, n4974, n4962, n3994, n3986}), .out(n13486), .config_in(config_chain[30891:30886]), .config_rst(config_rst)); 
buffer_wire buffer_13486 (.in(n13486), .out(n13486_0));
mux3 mux_8321 (.in({n12183_1, n12068_1, n5256}), .out(n13487), .config_in(config_chain[30893:30892]), .config_rst(config_rst)); 
buffer_wire buffer_13487 (.in(n13487), .out(n13487_0));
mux13 mux_8322 (.in({n13406_1/**/, n11129_1, n11109_1, n11092_0, n11078_0, n11073_0, n11066_0, n11061_0, n10982_1, n4974, n4966, n3994, n3986}), .out(n13488), .config_in(config_chain[30899:30894]), .config_rst(config_rst)); 
buffer_wire buffer_13488 (.in(n13488), .out(n13488_0));
mux3 mux_8323 (.in({n12185_1, n12076_1, n5260}), .out(n13489), .config_in(config_chain[30901:30900]), .config_rst(config_rst)); 
buffer_wire buffer_13489 (.in(n13489), .out(n13489_0));
mux13 mux_8324 (.in({n13408_1, n11131_1, n11100_0, n11095_0, n11086_0, n11081_0, n11052_0, n11041_0, n10974_1, n4974, n4966, n3998, n3986/**/}), .out(n13490), .config_in(config_chain[30907:30902]), .config_rst(config_rst)); 
buffer_wire buffer_13490 (.in(n13490), .out(n13490_0));
mux3 mux_8325 (.in({n12187_1, n12084_1, n5264}), .out(n13491), .config_in(config_chain[30909:30908]), .config_rst(config_rst)); 
buffer_wire buffer_13491 (.in(n13491), .out(n13491_0));
mux13 mux_8326 (.in({n13380_1, n11111_1, n11108_0, n11103_0, n11072_0, n11060_0, n11055_0, n11043_0, n10966_1/**/, n4974, n4966, n3998, n3990}), .out(n13492), .config_in(config_chain[30915:30910]), .config_rst(config_rst)); 
buffer_wire buffer_13492 (.in(n13492), .out(n13492_0));
mux3 mux_8327 (.in({n12093_1, n12092_1, n5268}), .out(n13493), .config_in(config_chain[30917:30916]), .config_rst(config_rst)); 
buffer_wire buffer_13493 (.in(n13493), .out(n13493_0));
mux15 mux_8328 (.in({n13410_1/**/, n11379_1, n11374_0, n11369_0, n11338_0, n11333_0, n11324_0, n11319_0, n11309_0, n11224_1, n5072, n5064, n4096, n4088, n4080}), .out(n13494), .config_in(config_chain[30923:30918]), .config_rst(config_rst)); 
buffer_wire buffer_13494 (.in(n13494), .out(n13494_0));
mux4 mux_8329 (.in({n12103_0, n12102_0, n5272, n4276}), .out(n13495), .config_in(config_chain[30925:30924]), .config_rst(config_rst)); 
buffer_wire buffer_13495 (.in(n13495), .out(n13495_0));
mux15 mux_8330 (.in({n13412_1, n11381_1, n11360_0, n11355_0, n11346_0, n11341_0, n11327_0/**/, n11311_0, n11306_1, n11304_1, n5076, n5064, n4096, n4088, n4080}), .out(n13496), .config_in(config_chain[30931:30926]), .config_rst(config_rst)); 
buffer_wire buffer_13496 (.in(n13496), .out(n13496_0));
mux3 mux_8331 (.in({n12105_0, n12104_0, n4280}), .out(n13497), .config_in(config_chain[30933:30932]), .config_rst(config_rst)); 
buffer_wire buffer_13497 (.in(n13497), .out(n13497_0));
mux15 mux_8332 (.in({n13414_1, n11383_1, n11368_0, n11363_0, n11349_0/**/, n11332_0, n11318_0, n11313_0, n11308_1, n11296_1, n5076, n5068, n4096, n4088, n4080}), .out(n13498), .config_in(config_chain[30939:30934]), .config_rst(config_rst)); 
buffer_wire buffer_13498 (.in(n13498), .out(n13498_0));
mux3 mux_8333 (.in({n12107_0, n12106_0, n4284}), .out(n13499), .config_in(config_chain[30941:30940]), .config_rst(config_rst)); 
buffer_wire buffer_13499 (.in(n13499), .out(n13499_0));
mux15 mux_8334 (.in({n13416_1, n11385_1, n11371_0, n11354_0, n11340_0, n11335_0, n11326_0, n11321_0, n11310_1, n11288_1, n5076, n5068, n5060, n4088, n4080}), .out(n13500), .config_in(config_chain[30947:30942]), .config_rst(config_rst)); 
buffer_wire buffer_13500 (.in(n13500), .out(n13500_0));
mux3 mux_8335 (.in({n12109_0, n12108_0/**/, n4284}), .out(n13501), .config_in(config_chain[30949:30948]), .config_rst(config_rst)); 
buffer_wire buffer_13501 (.in(n13501), .out(n13501_0));
mux14 mux_8336 (.in({n13418_1, n11387_1, n11362_0, n11357_0, n11348_0, n11343_0/**/, n11329_0, n11312_0, n11280_1, n5076, n5068, n5060, n4092, n4080}), .out(n13502), .config_in(config_chain[30955:30950]), .config_rst(config_rst)); 
buffer_wire buffer_13502 (.in(n13502), .out(n13502_0));
mux3 mux_8337 (.in({n12111_0, n12110_0, n4288}), .out(n13503), .config_in(config_chain[30957:30956]), .config_rst(config_rst)); 
buffer_wire buffer_13503 (.in(n13503), .out(n13503_0));
mux14 mux_8338 (.in({n13420_1, n11389_1/**/, n11370_0, n11365_0, n11351_0, n11334_0, n11320_0, n11315_0, n11272_1, n5076, n5068, n5060, n4092, n4084}), .out(n13504), .config_in(config_chain[30963:30958]), .config_rst(config_rst)); 
buffer_wire buffer_13504 (.in(n13504), .out(n13504_0));
mux3 mux_8339 (.in({n12113_0, n12112_0, n4292}), .out(n13505), .config_in(config_chain[30965:30964]), .config_rst(config_rst)); 
buffer_wire buffer_13505 (.in(n13505), .out(n13505_0));
mux13 mux_8340 (.in({n13422_1, n11391_1, n11373_0, n11356_0, n11342_0, n11337_0/**/, n11328_0, n11323_0, n11264_1, n5068, n5060, n4092, n4084}), .out(n13506), .config_in(config_chain[30971:30966]), .config_rst(config_rst)); 
buffer_wire buffer_13506 (.in(n13506), .out(n13506_0));
mux3 mux_8341 (.in({n12115_0/**/, n12114_0, n5256}), .out(n13507), .config_in(config_chain[30973:30972]), .config_rst(config_rst)); 
buffer_wire buffer_13507 (.in(n13507), .out(n13507_0));
mux13 mux_8342 (.in({n13424_1/**/, n11393_1, n11364_0, n11359_0, n11350_0, n11345_0, n11331_0, n11314_0, n11256_1, n5072, n5060, n4092, n4084}), .out(n13508), .config_in(config_chain[30979:30974]), .config_rst(config_rst)); 
buffer_wire buffer_13508 (.in(n13508), .out(n13508_0));
mux3 mux_8343 (.in({n12117_0/**/, n12116_0, n5260}), .out(n13509), .config_in(config_chain[30981:30980]), .config_rst(config_rst)); 
buffer_wire buffer_13509 (.in(n13509), .out(n13509_0));
mux13 mux_8344 (.in({n13426_1, n11395_1, n11372_0, n11367_0, n11353_1, n11336_0, n11322_0, n11317_0, n11248_1, n5072, n5064, n4092, n4084}), .out(n13510), .config_in(config_chain[30987:30982]), .config_rst(config_rst)); 
buffer_wire buffer_13510 (.in(n13510), .out(n13510_0));
mux3 mux_8345 (.in({n12119_0, n12118_0/**/, n5260}), .out(n13511), .config_in(config_chain[30989:30988]), .config_rst(config_rst)); 
buffer_wire buffer_13511 (.in(n13511), .out(n13511_0));
mux13 mux_8346 (.in({n13428_1, n11397_1, n11375_1, n11358_0, n11344_0, n11339_0, n11330_0, n11325_0, n11240_1, n5072, n5064, n4096, n4084}), .out(n13512), .config_in(config_chain[30995:30990]), .config_rst(config_rst)); 
buffer_wire buffer_13512 (.in(n13512), .out(n13512_0));
mux3 mux_8347 (.in({n12121_0, n12120_0, n5264}), .out(n13513), .config_in(config_chain[30997:30996]), .config_rst(config_rst)); 
buffer_wire buffer_13513 (.in(n13513), .out(n13513_0));
mux13 mux_8348 (.in({n13382_1, n11377_1, n11366_0, n11361_0, n11352_0, n11347_0, n11316_0, n11307_0, n11232_1, n5072, n5064, n4096, n4088}), .out(n13514), .config_in(config_chain[31003:30998]), .config_rst(config_rst)); 
buffer_wire buffer_13514 (.in(n13514), .out(n13514_0));
mux3 mux_8349 (.in({n12123_1, n12122_0, n5268}), .out(n13515), .config_in(config_chain[31005:31004]), .config_rst(config_rst)); 
buffer_wire buffer_13515 (.in(n13515), .out(n13515_0));
mux15 mux_8350 (.in({n13430_1, n11645_1, n11632_0, n11627_0, n11618_0, n11613_0, n11582_0, n11577_0/**/, n11573_0, n11490_1, n5170, n5162, n4194, n4186, n4178}), .out(n13516), .config_in(config_chain[31011:31006]), .config_rst(config_rst)); 
buffer_wire buffer_13516 (.in(n13516), .out(n13516_0));
mux4 mux_8351 (.in({n12125_0, n12124_0, n5272/**/, n4276}), .out(n13517), .config_in(config_chain[31013:31012]), .config_rst(config_rst)); 
buffer_wire buffer_13517 (.in(n13517), .out(n13517_0));
mux15 mux_8352 (.in({n13432_1, n11647_1, n11640_0, n11635_0, n11604_0/**/, n11599_0, n11590_0, n11585_0, n11575_0, n11570_1, n5174, n5162, n4194, n4186, n4178}), .out(n13518), .config_in(config_chain[31019:31014]), .config_rst(config_rst)); 
buffer_wire buffer_13518 (.in(n13518), .out(n13518_0));
mux3 mux_8353 (.in({n12127_0, n12126_0/**/, n4280}), .out(n13519), .config_in(config_chain[31021:31020]), .config_rst(config_rst)); 
buffer_wire buffer_13519 (.in(n13519), .out(n13519_0));
mux15 mux_8354 (.in({n13434_1, n11649_1, n11626_0, n11621_0, n11612_0, n11607_0, n11593_0, n11576_0, n11572_1, n11562_1, n5174, n5166/**/, n4194, n4186, n4178}), .out(n13520), .config_in(config_chain[31027:31022]), .config_rst(config_rst)); 
buffer_wire buffer_13520 (.in(n13520), .out(n13520_0));
mux3 mux_8355 (.in({n12129_0, n12128_0/**/, n4284}), .out(n13521), .config_in(config_chain[31029:31028]), .config_rst(config_rst)); 
buffer_wire buffer_13521 (.in(n13521), .out(n13521_0));
mux15 mux_8356 (.in({n13436_1, n11651_1, n11634_0, n11629_0, n11615_0, n11598_0, n11584_0, n11579_0, n11574_1, n11554_1, n5174/**/, n5166, n5158, n4186, n4178}), .out(n13522), .config_in(config_chain[31035:31030]), .config_rst(config_rst)); 
buffer_wire buffer_13522 (.in(n13522), .out(n13522_0));
mux3 mux_8357 (.in({n12131_0, n12130_0, n4288}), .out(n13523), .config_in(config_chain[31037:31036]), .config_rst(config_rst)); 
buffer_wire buffer_13523 (.in(n13523), .out(n13523_0));
mux14 mux_8358 (.in({n13438_1, n11653_1, n11637_0, n11620_0, n11606_0, n11601_0, n11592_0, n11587_0, n11546_1, n5174, n5166, n5158, n4190, n4178}), .out(n13524), .config_in(config_chain[31043:31038]), .config_rst(config_rst)); 
buffer_wire buffer_13524 (.in(n13524), .out(n13524_0));
mux3 mux_8359 (.in({n12133_0/**/, n12132_0, n4288}), .out(n13525), .config_in(config_chain[31045:31044]), .config_rst(config_rst)); 
buffer_wire buffer_13525 (.in(n13525), .out(n13525_0));
mux14 mux_8360 (.in({n13440_1, n11655_1, n11628_0, n11623_0, n11614_0, n11609_0, n11595_0, n11578_0, n11538_1/**/, n5174, n5166, n5158, n4190, n4182}), .out(n13526), .config_in(config_chain[31051:31046]), .config_rst(config_rst)); 
buffer_wire buffer_13526 (.in(n13526), .out(n13526_0));
mux3 mux_8361 (.in({n12135_0/**/, n12134_0, n4292}), .out(n13527), .config_in(config_chain[31053:31052]), .config_rst(config_rst)); 
buffer_wire buffer_13527 (.in(n13527), .out(n13527_0));
mux13 mux_8362 (.in({n13442_1, n11657_1, n11636_0, n11631_0, n11617_0, n11600_0, n11586_0, n11581_0, n11530_1/**/, n5166, n5158, n4190, n4182}), .out(n13528), .config_in(config_chain[31059:31054]), .config_rst(config_rst)); 
buffer_wire buffer_13528 (.in(n13528), .out(n13528_0));
mux3 mux_8363 (.in({n12137_0/**/, n12136_0, n5256}), .out(n13529), .config_in(config_chain[31061:31060]), .config_rst(config_rst)); 
buffer_wire buffer_13529 (.in(n13529), .out(n13529_0));
mux13 mux_8364 (.in({n13444_1, n11659_1, n11639_0, n11622_0, n11608_0/**/, n11603_0, n11594_0, n11589_0, n11522_1, n5170, n5158, n4190, n4182}), .out(n13530), .config_in(config_chain[31067:31062]), .config_rst(config_rst)); 
buffer_wire buffer_13530 (.in(n13530), .out(n13530_0));
mux3 mux_8365 (.in({n12139_0, n12138_0, n5260}), .out(n13531), .config_in(config_chain[31069:31068]), .config_rst(config_rst)); 
buffer_wire buffer_13531 (.in(n13531), .out(n13531_0));
mux13 mux_8366 (.in({n13446_1, n11661_1, n11630_0, n11625_0, n11616_0, n11611_0, n11597_1, n11580_0/**/, n11514_1, n5170, n5162, n4190, n4182}), .out(n13532), .config_in(config_chain[31075:31070]), .config_rst(config_rst)); 
buffer_wire buffer_13532 (.in(n13532), .out(n13532_0));
mux3 mux_8367 (.in({n12141_0, n12140_0, n5264}), .out(n13533), .config_in(config_chain[31077:31076]), .config_rst(config_rst)); 
buffer_wire buffer_13533 (.in(n13533), .out(n13533_0));
mux13 mux_8368 (.in({n13448_1, n11663_1, n11638_0, n11633_0, n11619_1, n11602_0/**/, n11588_0, n11583_0, n11506_1, n5170, n5162, n4194, n4182}), .out(n13534), .config_in(config_chain[31083:31078]), .config_rst(config_rst)); 
buffer_wire buffer_13534 (.in(n13534), .out(n13534_0));
mux3 mux_8369 (.in({n12143_0, n12142_0, n5264}), .out(n13535), .config_in(config_chain[31085:31084]), .config_rst(config_rst)); 
buffer_wire buffer_13535 (.in(n13535), .out(n13535_0));
mux13 mux_8370 (.in({n13384_2, n11643_1, n11641_1, n11624_0, n11610_0, n11605_0, n11596_0, n11591_0, n11498_1, n5170, n5162, n4194, n4186}), .out(n13536), .config_in(config_chain[31091:31086]), .config_rst(config_rst)); 
buffer_wire buffer_13536 (.in(n13536), .out(n13536_0));
mux3 mux_8371 (.in({n12145_1, n12144_0, n5268}), .out(n13537), .config_in(config_chain[31093:31092]), .config_rst(config_rst)); 
buffer_wire buffer_13537 (.in(n13537), .out(n13537_0));
mux15 mux_8372 (.in({n13450_1/**/, n11909_1, n11905_1, n11896_0, n11891_0, n11877_0, n11860_0, n11846_0, n11841_0, n11748_1, n5268, n5260, n4292, n4284, n4276}), .out(n13538), .config_in(config_chain[31099:31094]), .config_rst(config_rst)); 
buffer_wire buffer_13538 (.in(n13538), .out(n13538_0));
mux4 mux_8373 (.in({n12147_0, n12146_0, n5272, n4276}), .out(n13539), .config_in(config_chain[31101:31100]), .config_rst(config_rst)); 
buffer_wire buffer_13539 (.in(n13539), .out(n13539_0));
mux15 mux_8374 (.in({n13452_1, n11911_1, n11899_0, n11882_0, n11868_0, n11863_0, n11854_0, n11849_0, n11839_0, n11836_1, n5272, n5260, n4292, n4284, n4276}), .out(n13540), .config_in(config_chain[31107:31102]), .config_rst(config_rst)); 
buffer_wire buffer_13540 (.in(n13540), .out(n13540_0));
mux3 mux_8375 (.in({n12149_0, n12148_0, n4276}), .out(n13541), .config_in(config_chain[31109:31108]), .config_rst(config_rst)); 
buffer_wire buffer_13541 (.in(n13541), .out(n13541_0));
mux15 mux_8376 (.in({n13454_1, n11913_1, n11904_0, n11890_0, n11885_0, n11876_0, n11871_0, n11857_0, n11840_0, n11820_1/**/, n5272, n5264, n4292, n4284, n4276}), .out(n13542), .config_in(config_chain[31115:31110]), .config_rst(config_rst)); 
buffer_wire buffer_13542 (.in(n13542), .out(n13542_0));
mux3 mux_8377 (.in({n12151_0, n12150_0, n4280}), .out(n13543), .config_in(config_chain[31117:31116]), .config_rst(config_rst)); 
buffer_wire buffer_13543 (.in(n13543), .out(n13543_0));
mux15 mux_8378 (.in({n13456_1, n11915_1/**/, n11898_0, n11893_0, n11879_0, n11862_0, n11848_0, n11843_0, n11838_1, n11812_1, n5272, n5264, n5256, n4284, n4276}), .out(n13544), .config_in(config_chain[31123:31118]), .config_rst(config_rst)); 
buffer_wire buffer_13544 (.in(n13544), .out(n13544_0));
mux3 mux_8379 (.in({n12153_0, n12152_0, n4284}), .out(n13545), .config_in(config_chain[31125:31124]), .config_rst(config_rst)); 
buffer_wire buffer_13545 (.in(n13545), .out(n13545_0));
mux14 mux_8380 (.in({n13458_1, n11917_1, n11901_0, n11884_0, n11870_0, n11865_0, n11856_0, n11851_0, n11804_1/**/, n5272, n5264, n5256, n4288, n4276}), .out(n13546), .config_in(config_chain[31131:31126]), .config_rst(config_rst)); 
buffer_wire buffer_13546 (.in(n13546), .out(n13546_0));
mux3 mux_8381 (.in({n12155_0/**/, n12154_0, n4288}), .out(n13547), .config_in(config_chain[31133:31132]), .config_rst(config_rst)); 
buffer_wire buffer_13547 (.in(n13547), .out(n13547_0));
mux14 mux_8382 (.in({n13460_1, n11919_1, n11892_0, n11887_0, n11878_0, n11873_0, n11859_0, n11842_0, n11796_1/**/, n5272, n5264, n5256, n4288, n4280}), .out(n13548), .config_in(config_chain[31139:31134]), .config_rst(config_rst)); 
buffer_wire buffer_13548 (.in(n13548), .out(n13548_0));
mux3 mux_8383 (.in({n12157_0, n12156_0, n4292}), .out(n13549), .config_in(config_chain[31141:31140]), .config_rst(config_rst)); 
buffer_wire buffer_13549 (.in(n13549), .out(n13549_0));
mux13 mux_8384 (.in({n13462_1, n11921_1, n11900_0, n11895_0, n11881_0, n11864_0, n11850_0, n11845_0, n11788_1, n5264, n5256, n4288, n4280}), .out(n13550), .config_in(config_chain[31147:31142]), .config_rst(config_rst)); 
buffer_wire buffer_13550 (.in(n13550), .out(n13550_0));
mux3 mux_8385 (.in({n12159_0, n12158_0, n4292}), .out(n13551), .config_in(config_chain[31149:31148]), .config_rst(config_rst)); 
buffer_wire buffer_13551 (.in(n13551), .out(n13551_0));
mux13 mux_8386 (.in({n13464_1, n11923_1, n11903_0/**/, n11886_0, n11872_0, n11867_0, n11858_0, n11853_0, n11780_1, n5268, n5256, n4288, n4280}), .out(n13552), .config_in(config_chain[31155:31150]), .config_rst(config_rst)); 
buffer_wire buffer_13552 (.in(n13552), .out(n13552_0));
mux3 mux_8387 (.in({n12161_0, n12160_0, n5256}), .out(n13553), .config_in(config_chain[31157:31156]), .config_rst(config_rst)); 
buffer_wire buffer_13553 (.in(n13553), .out(n13553_0));
mux13 mux_8388 (.in({n13466_1, n11925_1, n11894_0, n11889_0, n11880_0, n11875_0, n11844_0, n11829_1, n11772_1, n5268, n5260, n4288, n4280}), .out(n13554), .config_in(config_chain[31163:31158]), .config_rst(config_rst)); 
buffer_wire buffer_13554 (.in(n13554), .out(n13554_0));
mux3 mux_8389 (.in({n12163_0, n12162_0, n5260}), .out(n13555), .config_in(config_chain[31165:31164]), .config_rst(config_rst)); 
buffer_wire buffer_13555 (.in(n13555), .out(n13555_0));
mux13 mux_8390 (.in({n13468_1, n11927_1, n11902_0, n11897_0, n11866_0, n11861_1, n11852_0, n11847_0/**/, n11764_1, n5268, n5260, n4292, n4280}), .out(n13556), .config_in(config_chain[31171:31166]), .config_rst(config_rst)); 
buffer_wire buffer_13556 (.in(n13556), .out(n13556_0));
mux3 mux_8391 (.in({n12165_0, n12164_0, n5264}), .out(n13557), .config_in(config_chain[31173:31172]), .config_rst(config_rst)); 
buffer_wire buffer_13557 (.in(n13557), .out(n13557_0));
mux13 mux_8392 (.in({n13386_2, n11907_1, n11888_0, n11883_1, n11874_0, n11869_0, n11855_0, n11828_1, n11756_1, n5268, n5260, n4292, n4284}), .out(n13558), .config_in(config_chain[31179:31174]), .config_rst(config_rst)); 
buffer_wire buffer_13558 (.in(n13558), .out(n13558_0));
mux3 mux_8393 (.in({n12167_1, n12166_0, n5268}), .out(n13559), .config_in(config_chain[31181:31180]), .config_rst(config_rst)); 
buffer_wire buffer_13559 (.in(n13559), .out(n13559_0));
mux4 mux_8394 (.in({n9819_0, n9818_0, n5466, n4470}), .out(n13560), .config_in(config_chain[31183:31182]), .config_rst(config_rst)); 
buffer_wire buffer_13560 (.in(n13560), .out(n13560_0));
mux15 mux_8395 (.in({n13693_1, n10625_1/**/, n10599_0, n10592_0, n10580_0, n10553_0, n10546_0, n10528_1, n10522_1, n10519_0, n5658, n5650, n4682, n4674, n4666}), .out(n13561), .config_in(config_chain[31189:31184]), .config_rst(config_rst)); 
buffer_wire buffer_13561 (.in(n13561), .out(n13561_0));
mux4 mux_8396 (.in({n9839_1, n9758_1/**/, n5466, n4470}), .out(n13562), .config_in(config_chain[31191:31190]), .config_rst(config_rst)); 
buffer_wire buffer_13562 (.in(n13562), .out(n13562_0));
mux15 mux_8397 (.in({n13715_1/**/, n10887_1, n10853_0, n10846_0, n10839_0, n10832_0, n10820_0, n10788_1, n10782_1, n10779_0, n5756, n5748, n4780, n4772, n4764}), .out(n13563), .config_in(config_chain[31197:31192]), .config_rst(config_rst)); 
buffer_wire buffer_13563 (.in(n13563), .out(n13563_0));
mux4 mux_8398 (.in({n9779_0, n9778_0, n5466, n4470/**/}), .out(n13564), .config_in(config_chain[31199:31198]), .config_rst(config_rst)); 
buffer_wire buffer_13564 (.in(n13564), .out(n13564_0));
mux16 mux_8399 (.in({n13653_1, n10109_1, n10078_0, n10075_0, n10069_0, n10052_0, n10044_0, n10041_0, n10014_1, n10009_1, n10000_1, n5462, n5454, n4486, n4478, n4470/**/}), .out(n13565), .config_in(config_chain[31205:31200]), .config_rst(config_rst)); 
buffer_wire buffer_13565 (.in(n13565), .out(n13565_0));
mux4 mux_8400 (.in({n9799_0, n9798_0, n5466, n4470/**/}), .out(n13566), .config_in(config_chain[31207:31206]), .config_rst(config_rst)); 
buffer_wire buffer_13566 (.in(n13566), .out(n13566_0));
mux16 mux_8401 (.in({n13673_1, n10365_1, n10340_0, n10337_0, n10314_0, n10311_0, n10305_0, n10288_0, n10270_1, n10265_1, n10256_1, n5560, n5552, n4584, n4576, n4568}), .out(n13567), .config_in(config_chain[31213:31208]), .config_rst(config_rst)); 
buffer_wire buffer_13567 (.in(n13567), .out(n13567_0));
mux3 mux_8402 (.in({n9821_0, n9820_0/**/, n4470}), .out(n13568), .config_in(config_chain[31215:31214]), .config_rst(config_rst)); 
buffer_wire buffer_13568 (.in(n13568), .out(n13568_0));
mux15 mux_8403 (.in({n13695_1, n10623_1, n10600_0, n10573_0, n10566_0, n10561_0, n10554_0/**/, n10530_1, n10524_1, n10521_0, n5662, n5650, n4682, n4674, n4666}), .out(n13569), .config_in(config_chain[31221:31216]), .config_rst(config_rst)); 
buffer_wire buffer_13569 (.in(n13569), .out(n13569_0));
mux3 mux_8404 (.in({n9841_1, n9760_1, n4474/**/}), .out(n13570), .config_in(config_chain[31223:31222]), .config_rst(config_rst)); 
buffer_wire buffer_13570 (.in(n13570), .out(n13570_0));
mux15 mux_8405 (.in({n13717_1/**/, n10885_1, n10861_0, n10854_0, n10840_0, n10813_0, n10806_0, n10790_1, n10784_1, n10781_0, n5760, n5748, n4780, n4772, n4764}), .out(n13571), .config_in(config_chain[31229:31224]), .config_rst(config_rst)); 
buffer_wire buffer_13571 (.in(n13571), .out(n13571_0));
mux3 mux_8406 (.in({n9781_0/**/, n9780_0, n4474}), .out(n13572), .config_in(config_chain[31231:31230]), .config_rst(config_rst)); 
buffer_wire buffer_13572 (.in(n13572), .out(n13572_0));
mux16 mux_8407 (.in({n13655_1, n10107_1, n10089_0, n10072_0, n10066_0, n10063_0, n10038_0, n10035_0, n10016_1, n10011_1, n10002_1, n5462, n5454, n4486, n4478, n4470/**/}), .out(n13573), .config_in(config_chain[31237:31232]), .config_rst(config_rst)); 
buffer_wire buffer_13573 (.in(n13573), .out(n13573_0));
mux3 mux_8408 (.in({n9801_0, n9800_0, n4474/**/}), .out(n13574), .config_in(config_chain[31239:31238]), .config_rst(config_rst)); 
buffer_wire buffer_13574 (.in(n13574), .out(n13574_0));
mux16 mux_8409 (.in({n13675_1, n10363_1, n10334_0, n10331_0, n10325_0, n10308_0/**/, n10302_0, n10299_0, n10272_1, n10267_1, n10258_1, n5560, n5552, n4584, n4576, n4568}), .out(n13575), .config_in(config_chain[31245:31240]), .config_rst(config_rst)); 
buffer_wire buffer_13575 (.in(n13575), .out(n13575_0));
mux3 mux_8410 (.in({n9823_0/**/, n9822_0, n4474}), .out(n13576), .config_in(config_chain[31247:31246]), .config_rst(config_rst)); 
buffer_wire buffer_13576 (.in(n13576), .out(n13576_0));
mux15 mux_8411 (.in({n13697_1, n10621_1, n10593_0, n10586_0, n10581_0, n10574_0, n10562_0, n10547_0, n10532_1, n10523_1, n5662, n5654, n4682, n4674, n4666}), .out(n13577), .config_in(config_chain[31253:31248]), .config_rst(config_rst)); 
buffer_wire buffer_13577 (.in(n13577), .out(n13577_0));
mux3 mux_8412 (.in({n9843_1, n9762_1/**/, n4474}), .out(n13578), .config_in(config_chain[31255:31254]), .config_rst(config_rst)); 
buffer_wire buffer_13578 (.in(n13578), .out(n13578_0));
mux15 mux_8413 (.in({n13719_1, n10883_1, n10862_0, n10847_0, n10833_0, n10826_0, n10821_0, n10814_0, n10792_1, n10783_0, n5760, n5752, n4780, n4772, n4764}), .out(n13579), .config_in(config_chain[31261:31256]), .config_rst(config_rst)); 
buffer_wire buffer_13579 (.in(n13579), .out(n13579_0));
mux3 mux_8414 (.in({n9783_0, n9782_0, n4478}), .out(n13580), .config_in(config_chain[31263:31262]), .config_rst(config_rst)); 
buffer_wire buffer_13580 (.in(n13580), .out(n13580_0));
mux15 mux_8415 (.in({n13657_1, n10105_1, n10086_0, n10083_0, n10060_0, n10057_0, n10049_0, n10032_0, n10018_1, n10004_1, n5462, n5454, n4486, n4478, n4470}), .out(n13581), .config_in(config_chain[31269:31264]), .config_rst(config_rst)); 
buffer_wire buffer_13581 (.in(n13581), .out(n13581_0));
mux3 mux_8416 (.in({n9803_0, n9802_0, n4478}), .out(n13582), .config_in(config_chain[31271:31270]), .config_rst(config_rst)); 
buffer_wire buffer_13582 (.in(n13582), .out(n13582_0));
mux15 mux_8417 (.in({n13677_1, n10361_1, n10345_0, n10328_0, n10322_0, n10319_0, n10296_0, n10293_0, n10274_1/**/, n10260_1, n5560, n5552, n4584, n4576, n4568}), .out(n13583), .config_in(config_chain[31277:31272]), .config_rst(config_rst)); 
buffer_wire buffer_13583 (.in(n13583), .out(n13583_0));
mux3 mux_8418 (.in({n9825_0, n9824_0/**/, n4478}), .out(n13584), .config_in(config_chain[31279:31278]), .config_rst(config_rst)); 
buffer_wire buffer_13584 (.in(n13584), .out(n13584_0));
mux15 mux_8419 (.in({n13699_1, n10619_1, n10601_0, n10594_0, n10582_0, n10567_0, n10555_0, n10548_0, n10534_1, n10525_1, n5662/**/, n5654, n5646, n4674, n4666}), .out(n13585), .config_in(config_chain[31285:31280]), .config_rst(config_rst)); 
buffer_wire buffer_13585 (.in(n13585), .out(n13585_0));
mux3 mux_8420 (.in({n9845_1, n9764_1, n4478}), .out(n13586), .config_in(config_chain[31287:31286]), .config_rst(config_rst)); 
buffer_wire buffer_13586 (.in(n13586), .out(n13586_0));
mux15 mux_8421 (.in({n13721_1, n10881_1, n10855_0, n10848_0, n10841_0, n10834_0, n10822_0, n10807_0, n10794_1, n10785_1, n5760, n5752, n5744, n4772, n4764/**/}), .out(n13587), .config_in(config_chain[31293:31288]), .config_rst(config_rst)); 
buffer_wire buffer_13587 (.in(n13587), .out(n13587_0));
mux3 mux_8422 (.in({n9785_0, n9784_0/**/, n4478}), .out(n13588), .config_in(config_chain[31295:31294]), .config_rst(config_rst)); 
buffer_wire buffer_13588 (.in(n13588), .out(n13588_0));
mux15 mux_8423 (.in({n13659_1, n10103_1, n10080_0, n10077_0, n10071_0, n10054_0, n10046_0, n10043_0, n10020_1, n10006_1, n5462, n5454, n4486, n4478, n4470}), .out(n13589), .config_in(config_chain[31301:31296]), .config_rst(config_rst)); 
buffer_wire buffer_13589 (.in(n13589), .out(n13589_0));
mux3 mux_8424 (.in({n9805_0, n9804_0, n4482}), .out(n13590), .config_in(config_chain[31303:31302]), .config_rst(config_rst)); 
buffer_wire buffer_13590 (.in(n13590), .out(n13590_0));
mux15 mux_8425 (.in({n13679_1, n10359_1, n10342_0, n10339_0, n10316_0, n10313_0/**/, n10307_0, n10290_0, n10276_1, n10262_1, n5560, n5552, n4584, n4576, n4568}), .out(n13591), .config_in(config_chain[31309:31304]), .config_rst(config_rst)); 
buffer_wire buffer_13591 (.in(n13591), .out(n13591_0));
mux3 mux_8426 (.in({n9827_0, n9826_0/**/, n4482}), .out(n13592), .config_in(config_chain[31311:31310]), .config_rst(config_rst)); 
buffer_wire buffer_13592 (.in(n13592), .out(n13592_0));
mux14 mux_8427 (.in({n13701_1/**/, n10617_1, n10602_0, n10587_0, n10575_0, n10568_0, n10563_0, n10556_0, n10536_1, n5662, n5654, n5646, n4678, n4666}), .out(n13593), .config_in(config_chain[31317:31312]), .config_rst(config_rst)); 
buffer_wire buffer_13593 (.in(n13593), .out(n13593_0));
mux3 mux_8428 (.in({n9847_1, n9766_1, n4482}), .out(n13594), .config_in(config_chain[31319:31318]), .config_rst(config_rst)); 
buffer_wire buffer_13594 (.in(n13594), .out(n13594_0));
mux14 mux_8429 (.in({n13723_1, n10879_1, n10863_0, n10856_0, n10842_0, n10827_0, n10815_0, n10808_0, n10796_1, n5760/**/, n5752, n5744, n4776, n4764}), .out(n13595), .config_in(config_chain[31325:31320]), .config_rst(config_rst)); 
buffer_wire buffer_13595 (.in(n13595), .out(n13595_0));
mux3 mux_8430 (.in({n9787_0, n9786_0/**/, n4482}), .out(n13596), .config_in(config_chain[31327:31326]), .config_rst(config_rst)); 
buffer_wire buffer_13596 (.in(n13596), .out(n13596_0));
mux15 mux_8431 (.in({n13661_1, n10101_1, n10091_0, n10074_0, n10068_0, n10065_0, n10040_0, n10037_0, n10022_1/**/, n10008_1, n5462, n5454, n4486, n4478, n4470}), .out(n13597), .config_in(config_chain[31333:31328]), .config_rst(config_rst)); 
buffer_wire buffer_13597 (.in(n13597), .out(n13597_0));
mux3 mux_8432 (.in({n9807_0, n9806_0, n4482}), .out(n13598), .config_in(config_chain[31335:31334]), .config_rst(config_rst)); 
buffer_wire buffer_13598 (.in(n13598), .out(n13598_0));
mux15 mux_8433 (.in({n13681_1, n10357_1, n10336_0, n10333_0, n10327_0, n10310_0/**/, n10304_0, n10301_0, n10278_1, n10264_1, n5560, n5552, n4584, n4576, n4568}), .out(n13599), .config_in(config_chain[31341:31336]), .config_rst(config_rst)); 
buffer_wire buffer_13599 (.in(n13599), .out(n13599_0));
mux3 mux_8434 (.in({n9829_0, n9828_0/**/, n4486}), .out(n13600), .config_in(config_chain[31343:31342]), .config_rst(config_rst)); 
buffer_wire buffer_13600 (.in(n13600), .out(n13600_0));
mux14 mux_8435 (.in({n13703_1, n10615_1/**/, n10595_0, n10588_0, n10583_0, n10576_0, n10564_0, n10549_0, n10538_1, n5662, n5654, n5646, n4678, n4670}), .out(n13601), .config_in(config_chain[31349:31344]), .config_rst(config_rst)); 
buffer_wire buffer_13601 (.in(n13601), .out(n13601_0));
mux3 mux_8436 (.in({n9849_1, n9768_1, n4486}), .out(n13602), .config_in(config_chain[31351:31350]), .config_rst(config_rst)); 
buffer_wire buffer_13602 (.in(n13602), .out(n13602_0));
mux14 mux_8437 (.in({n13725_1, n10877_1, n10864_0/**/, n10849_0, n10835_0, n10828_0, n10823_0, n10816_0, n10798_1, n5760, n5752, n5744, n4776, n4768}), .out(n13603), .config_in(config_chain[31357:31352]), .config_rst(config_rst)); 
buffer_wire buffer_13603 (.in(n13603), .out(n13603_0));
mux3 mux_8438 (.in({n9789_0, n9788_0, n4486/**/}), .out(n13604), .config_in(config_chain[31359:31358]), .config_rst(config_rst)); 
buffer_wire buffer_13604 (.in(n13604), .out(n13604_0));
mux15 mux_8439 (.in({n13663_1, n10099_1, n10088_0, n10085_0, n10062_0, n10059_0/**/, n10051_0, n10034_0, n10024_1, n10010_1, n5466, n5458, n5450, n4482, n4474}), .out(n13605), .config_in(config_chain[31365:31360]), .config_rst(config_rst)); 
buffer_wire buffer_13605 (.in(n13605), .out(n13605_0));
mux3 mux_8440 (.in({n9809_0, n9808_0, n4486}), .out(n13606), .config_in(config_chain[31367:31366]), .config_rst(config_rst)); 
buffer_wire buffer_13606 (.in(n13606), .out(n13606_0));
mux15 mux_8441 (.in({n13683_1, n10355_1, n10347_0, n10330_0, n10324_0, n10321_0, n10298_0, n10295_0, n10280_1, n10266_1, n5564, n5556, n5548, n4580, n4572}), .out(n13607), .config_in(config_chain[31373:31368]), .config_rst(config_rst)); 
buffer_wire buffer_13607 (.in(n13607), .out(n13607_0));
mux3 mux_8442 (.in({n9831_0, n9830_0/**/, n4486}), .out(n13608), .config_in(config_chain[31375:31374]), .config_rst(config_rst)); 
buffer_wire buffer_13608 (.in(n13608), .out(n13608_0));
mux13 mux_8443 (.in({n13705_1, n10613_1, n10603_0, n10596_0, n10584_0, n10569_0, n10557_0, n10550_0, n10540_1, n5654/**/, n5646, n4678, n4670}), .out(n13609), .config_in(config_chain[31381:31376]), .config_rst(config_rst)); 
buffer_wire buffer_13609 (.in(n13609), .out(n13609_0));
mux3 mux_8444 (.in({n9851_1, n9770_1, n5450}), .out(n13610), .config_in(config_chain[31383:31382]), .config_rst(config_rst)); 
buffer_wire buffer_13610 (.in(n13610), .out(n13610_0));
mux13 mux_8445 (.in({n13727_1/**/, n10875_1, n10857_0, n10850_0, n10843_0, n10836_0, n10824_0, n10809_0, n10800_1, n5752, n5744, n4776, n4768}), .out(n13611), .config_in(config_chain[31389:31384]), .config_rst(config_rst)); 
buffer_wire buffer_13611 (.in(n13611), .out(n13611_0));
mux3 mux_8446 (.in({n9791_0/**/, n9790_0, n5450}), .out(n13612), .config_in(config_chain[31391:31390]), .config_rst(config_rst)); 
buffer_wire buffer_13612 (.in(n13612), .out(n13612_0));
mux15 mux_8447 (.in({n13665_1, n10097_1, n10082_0, n10079_0, n10056_0, n10053_0, n10048_0, n10045_0, n10026_1, n10001_0, n5466, n5458, n5450, n4482, n4474}), .out(n13613), .config_in(config_chain[31397:31392]), .config_rst(config_rst)); 
buffer_wire buffer_13613 (.in(n13613), .out(n13613_0));
mux3 mux_8448 (.in({n9811_0, n9810_0, n5450}), .out(n13614), .config_in(config_chain[31399:31398]), .config_rst(config_rst)); 
buffer_wire buffer_13614 (.in(n13614), .out(n13614_0));
mux15 mux_8449 (.in({n13685_1, n10353_1, n10344_0, n10341_0, n10318_0/**/, n10315_0, n10292_0, n10289_0, n10282_1, n10257_0, n5564, n5556, n5548, n4580, n4572}), .out(n13615), .config_in(config_chain[31405:31400]), .config_rst(config_rst)); 
buffer_wire buffer_13615 (.in(n13615), .out(n13615_0));
mux3 mux_8450 (.in({n9833_0, n9832_0/**/, n5450}), .out(n13616), .config_in(config_chain[31407:31406]), .config_rst(config_rst)); 
buffer_wire buffer_13616 (.in(n13616), .out(n13616_0));
mux13 mux_8451 (.in({n13707_1, n10611_1, n10604_0, n10589_0, n10577_0, n10570_0, n10565_0, n10558_0, n10542_1, n5658, n5646, n4678, n4670}), .out(n13617), .config_in(config_chain[31413:31408]), .config_rst(config_rst)); 
buffer_wire buffer_13617 (.in(n13617), .out(n13617_0));
mux3 mux_8452 (.in({n9853_1, n9772_1, n5450}), .out(n13618), .config_in(config_chain[31415:31414]), .config_rst(config_rst)); 
buffer_wire buffer_13618 (.in(n13618), .out(n13618_0));
mux13 mux_8453 (.in({n13729_1, n10873_1, n10865_0, n10858_0/**/, n10844_0, n10829_0, n10817_0, n10810_0, n10802_1, n5756, n5744, n4776, n4768}), .out(n13619), .config_in(config_chain[31421:31416]), .config_rst(config_rst)); 
buffer_wire buffer_13619 (.in(n13619), .out(n13619_0));
mux3 mux_8454 (.in({n9793_0, n9792_0, n5454}), .out(n13620), .config_in(config_chain[31423:31422]), .config_rst(config_rst)); 
buffer_wire buffer_13620 (.in(n13620), .out(n13620_0));
mux15 mux_8455 (.in({n13667_1, n10095_1, n10076_0, n10073_0, n10070_0, n10067_0, n10042_0, n10039_0/**/, n10028_1, n10003_0, n5466, n5458, n5450, n4482, n4474}), .out(n13621), .config_in(config_chain[31429:31424]), .config_rst(config_rst)); 
buffer_wire buffer_13621 (.in(n13621), .out(n13621_0));
mux3 mux_8456 (.in({n9813_0, n9812_0, n5454}), .out(n13622), .config_in(config_chain[31431:31430]), .config_rst(config_rst)); 
buffer_wire buffer_13622 (.in(n13622), .out(n13622_0));
mux15 mux_8457 (.in({n13687_1, n10351_1, n10338_0, n10335_0, n10312_0, n10309_0/**/, n10306_0, n10303_0, n10284_1, n10259_0, n5564, n5556, n5548, n4580, n4572}), .out(n13623), .config_in(config_chain[31437:31432]), .config_rst(config_rst)); 
buffer_wire buffer_13623 (.in(n13623), .out(n13623_0));
mux3 mux_8458 (.in({n9835_0, n9834_0/**/, n5454}), .out(n13624), .config_in(config_chain[31439:31438]), .config_rst(config_rst)); 
buffer_wire buffer_13624 (.in(n13624), .out(n13624_0));
mux13 mux_8459 (.in({n13709_1, n10609_1, n10597_0, n10590_0, n10585_0, n10578_0, n10551_0, n10544_1, n10516_1, n5658, n5650, n4678/**/, n4670}), .out(n13625), .config_in(config_chain[31445:31440]), .config_rst(config_rst)); 
buffer_wire buffer_13625 (.in(n13625), .out(n13625_0));
mux3 mux_8460 (.in({n9855_1, n9774_1/**/, n5454}), .out(n13626), .config_in(config_chain[31447:31446]), .config_rst(config_rst)); 
buffer_wire buffer_13626 (.in(n13626), .out(n13626_0));
mux13 mux_8461 (.in({n13731_1, n10871_1, n10866_0, n10851_0, n10837_0, n10830_0, n10825_0, n10818_0, n10804_1, n5756, n5748, n4776/**/, n4768}), .out(n13627), .config_in(config_chain[31453:31448]), .config_rst(config_rst)); 
buffer_wire buffer_13627 (.in(n13627), .out(n13627_0));
mux3 mux_8462 (.in({n9795_0, n9794_0, n5454}), .out(n13628), .config_in(config_chain[31455:31454]), .config_rst(config_rst)); 
buffer_wire buffer_13628 (.in(n13628), .out(n13628_0));
mux15 mux_8463 (.in({n13669_1, n10093_1, n10090_0/**/, n10087_0, n10064_0, n10061_0, n10036_0, n10033_0, n10030_1, n10005_1, n5466, n5458, n5450, n4482, n4474}), .out(n13629), .config_in(config_chain[31461:31456]), .config_rst(config_rst)); 
buffer_wire buffer_13629 (.in(n13629), .out(n13629_0));
mux3 mux_8464 (.in({n9815_0, n9814_0, n5458}), .out(n13630), .config_in(config_chain[31463:31462]), .config_rst(config_rst)); 
buffer_wire buffer_13630 (.in(n13630), .out(n13630_0));
mux15 mux_8465 (.in({n13689_1, n10349_1, n10332_0, n10329_0, n10326_0, n10323_0, n10300_0, n10297_0, n10286_1, n10261_0, n5564, n5556, n5548, n4580, n4572}), .out(n13631), .config_in(config_chain[31469:31464]), .config_rst(config_rst)); 
buffer_wire buffer_13631 (.in(n13631), .out(n13631_0));
mux3 mux_8466 (.in({n9837_0, n9836_0/**/, n5458}), .out(n13632), .config_in(config_chain[31471:31470]), .config_rst(config_rst)); 
buffer_wire buffer_13632 (.in(n13632), .out(n13632_0));
mux13 mux_8467 (.in({n13711_1/**/, n10607_1, n10605_0, n10598_0, n10571_0, n10559_0, n10552_0, n10518_1, n10514_1, n5658, n5650, n4682, n4670}), .out(n13633), .config_in(config_chain[31477:31472]), .config_rst(config_rst)); 
buffer_wire buffer_13633 (.in(n13633), .out(n13633_0));
mux3 mux_8468 (.in({n9857_1, n9776_1, n5458}), .out(n13634), .config_in(config_chain[31479:31478]), .config_rst(config_rst)); 
buffer_wire buffer_13634 (.in(n13634), .out(n13634_0));
mux13 mux_8469 (.in({n13733_1, n10869_1, n10859_0, n10852_0, n10845_0/**/, n10838_0, n10811_0, n10778_1, n10776_1, n5756, n5748, n4780, n4768}), .out(n13635), .config_in(config_chain[31485:31480]), .config_rst(config_rst)); 
buffer_wire buffer_13635 (.in(n13635), .out(n13635_0));
mux3 mux_8470 (.in({n9797_0, n9796_0, n5458}), .out(n13636), .config_in(config_chain[31487:31486]), .config_rst(config_rst)); 
buffer_wire buffer_13636 (.in(n13636), .out(n13636_0));
mux15 mux_8471 (.in({n13671_1, n10111_1, n10084_0, n10081_0, n10058_0, n10055_0, n10050_0, n10047_0, n10012_1, n10007_1, n5466/**/, n5458, n5450, n4482, n4474}), .out(n13637), .config_in(config_chain[31493:31488]), .config_rst(config_rst)); 
buffer_wire buffer_13637 (.in(n13637), .out(n13637_0));
mux3 mux_8472 (.in({n9817_0, n9816_0/**/, n5458}), .out(n13638), .config_in(config_chain[31495:31494]), .config_rst(config_rst)); 
buffer_wire buffer_13638 (.in(n13638), .out(n13638_0));
mux15 mux_8473 (.in({n13691_1, n10367_1, n10346_0, n10343_0, n10320_0, n10317_0, n10294_0, n10291_0, n10268_1/**/, n10263_1, n5564, n5556, n5548, n4580, n4572}), .out(n13639), .config_in(config_chain[31501:31496]), .config_rst(config_rst)); 
buffer_wire buffer_13639 (.in(n13639), .out(n13639_0));
mux3 mux_8474 (.in({n9747_0, n9746_1, n5462}), .out(n13640), .config_in(config_chain[31503:31502]), .config_rst(config_rst)); 
buffer_wire buffer_13640 (.in(n13640), .out(n13640_0));
mux13 mux_8475 (.in({n13713_1, n10627_1, n10591_0, n10579_0, n10572_0, n10560_0/**/, n10526_1, n10520_1, n10517_0, n5658, n5650, n4682, n4674}), .out(n13641), .config_in(config_chain[31509:31504]), .config_rst(config_rst)); 
buffer_wire buffer_13641 (.in(n13641), .out(n13641_0));
mux3 mux_8476 (.in({n9749_1, n9748_1, n5462}), .out(n13642), .config_in(config_chain[31511:31510]), .config_rst(config_rst)); 
buffer_wire buffer_13642 (.in(n13642), .out(n13642_0));
mux13 mux_8477 (.in({n13735_1, n10889_1, n10867_1, n10860_0, n10831_0, n10819_0, n10812_0, n10786_1, n10780_1, n5756, n5748, n4780, n4772}), .out(n13643), .config_in(config_chain[31517:31512]), .config_rst(config_rst)); 
buffer_wire buffer_13643 (.in(n13643), .out(n13643_0));
mux3 mux_8478 (.in({n9751_1, n9750_1, n5462}), .out(n13644), .config_in(config_chain[31519:31518]), .config_rst(config_rst)); 
buffer_wire buffer_13644 (.in(n13644), .out(n13644_0));
mux13 mux_8479 (.in({n13757_1, n11153_1, n11123_0, n11116_0, n11109_1, n11102_0, n11073_0, n11048_1, n11042_1, n5854, n5846, n4878, n4870}), .out(n13645), .config_in(config_chain[31525:31520]), .config_rst(config_rst)); 
buffer_wire buffer_13645 (.in(n13645), .out(n13645_0));
mux3 mux_8480 (.in({n9753_1, n9752_1, n5462}), .out(n13646), .config_in(config_chain[31527:31526]), .config_rst(config_rst)); 
buffer_wire buffer_13646 (.in(n13646), .out(n13646_0));
mux13 mux_8481 (.in({n13779_0, n11419_1, n11396_0, n11381_0, n11367_0, n11360_0, n11353_1, n11346_0, n11312_1, n5952, n5944, n4976, n4968}), .out(n13647), .config_in(config_chain[31533:31528]), .config_rst(config_rst)); 
buffer_wire buffer_13647 (.in(n13647), .out(n13647_0));
mux3 mux_8482 (.in({n9755_1, n9754_1, n5462}), .out(n13648), .config_in(config_chain[31535:31534]), .config_rst(config_rst)); 
buffer_wire buffer_13648 (.in(n13648), .out(n13648_0));
mux13 mux_8483 (.in({n13801_0, n11685_1, n11647_0, n11640_0, n11633_0, n11626_0, n11612_0, n11597_1, n11576_1/**/, n6050, n6042, n5074, n5066}), .out(n13649), .config_in(config_chain[31541:31536]), .config_rst(config_rst)); 
buffer_wire buffer_13649 (.in(n13649), .out(n13649_0));
mux3 mux_8484 (.in({n9757_1, n9756_1, n5466}), .out(n13650), .config_in(config_chain[31543:31542]), .config_rst(config_rst)); 
buffer_wire buffer_13650 (.in(n13650), .out(n13650_0));
mux13 mux_8485 (.in({n13823_0, n11949_1, n11920_0, n11889_0, n11882_0, n11875_0, n11868_0/**/, n11840_1, n11829_1, n6148, n6140, n5172, n5164}), .out(n13651), .config_in(config_chain[31549:31544]), .config_rst(config_rst)); 
buffer_wire buffer_13651 (.in(n13651), .out(n13651_0));
mux16 mux_8486 (.in({n13564_0, n10095_1, n10079_0, n10074_0, n10068_0, n10053_0/**/, n10045_0, n10040_0, n10012_1, n10008_1, n10001_0, n5560, n5552, n4584, n4576, n4568}), .out(n13652), .config_in(config_chain[31555:31550]), .config_rst(config_rst)); 
buffer_wire buffer_13652 (.in(n13652), .out(n13652_0));
mux15 mux_8487 (.in({n13737_1, n11151_1, n11131_1, n11124_0, n11095_0, n11088_0, n11081_0, n11074_0, n11050_1, n11044_1, n5854, n5846, n4878/**/, n4870, n4862}), .out(n13653), .config_in(config_chain[31561:31556]), .config_rst(config_rst)); 
buffer_wire buffer_13653 (.in(n13653), .out(n13653_0));
mux16 mux_8488 (.in({n13572_0, n10097_1, n10088_0, n10073_0, n10067_0, n10062_0, n10039_0, n10034_0, n10030_1/**/, n10010_1, n10003_0, n5560, n5552, n4584, n4576, n4568}), .out(n13654), .config_in(config_chain[31567:31562]), .config_rst(config_rst)); 
buffer_wire buffer_13654 (.in(n13654), .out(n13654_0));
mux15 mux_8489 (.in({n13739_1, n11149_1, n11117_0, n11110_0, n11103_0, n11096_0, n11082_0, n11052_1/**/, n11046_1, n11043_0, n5858, n5846, n4878, n4870, n4862}), .out(n13655), .config_in(config_chain[31573:31568]), .config_rst(config_rst)); 
buffer_wire buffer_13655 (.in(n13655), .out(n13655_0));
mux15 mux_8490 (.in({n13580_0, n10099_1, n10087_0, n10082_0, n10061_0, n10056_0, n10048_0, n10033_0/**/, n10028_1, n10005_1, n5560, n5552, n4584, n4576, n4568}), .out(n13656), .config_in(config_chain[31579:31574]), .config_rst(config_rst)); 
buffer_wire buffer_13656 (.in(n13656), .out(n13656_0));
mux15 mux_8491 (.in({n13741_1, n11147_1, n11125_0, n11118_0, n11104_0/**/, n11089_0, n11075_0, n11068_0, n11054_1, n11045_0, n5858, n5850, n4878, n4870, n4862}), .out(n13657), .config_in(config_chain[31585:31580]), .config_rst(config_rst)); 
buffer_wire buffer_13657 (.in(n13657), .out(n13657_0));
mux15 mux_8492 (.in({n13588_0, n10101_1, n10081_0, n10076_0/**/, n10070_0, n10055_0, n10047_0, n10042_0, n10026_1, n10007_1, n5560, n5552, n4584, n4576, n4568}), .out(n13658), .config_in(config_chain[31591:31586]), .config_rst(config_rst)); 
buffer_wire buffer_13658 (.in(n13658), .out(n13658_0));
mux15 mux_8493 (.in({n13743_1, n11145_1, n11126_0, n11111_0/**/, n11097_0, n11090_0, n11083_0, n11076_0, n11056_1, n11047_0, n5858, n5850, n5842, n4870, n4862}), .out(n13659), .config_in(config_chain[31597:31592]), .config_rst(config_rst)); 
buffer_wire buffer_13659 (.in(n13659), .out(n13659_0));
mux15 mux_8494 (.in({n13596_0, n10103_1, n10090_0, n10075_0, n10069_0, n10064_0, n10041_0, n10036_0, n10024_1, n10009_1, n5560, n5552, n4584/**/, n4576, n4568}), .out(n13660), .config_in(config_chain[31603:31598]), .config_rst(config_rst)); 
buffer_wire buffer_13660 (.in(n13660), .out(n13660_0));
mux14 mux_8495 (.in({n13745_1, n11143_1, n11119_0, n11112_0, n11105_0, n11098_0, n11084_0, n11069_0, n11058_1, n5858, n5850, n5842/**/, n4874, n4862}), .out(n13661), .config_in(config_chain[31609:31604]), .config_rst(config_rst)); 
buffer_wire buffer_13661 (.in(n13661), .out(n13661_0));
mux15 mux_8496 (.in({n13604_0, n10105_1, n10089_0, n10084_0, n10063_0, n10058_0, n10050_0, n10035_0/**/, n10022_1, n10011_1, n5564, n5556, n5548, n4580, n4572}), .out(n13662), .config_in(config_chain[31615:31610]), .config_rst(config_rst)); 
buffer_wire buffer_13662 (.in(n13662), .out(n13662_0));
mux14 mux_8497 (.in({n13747_1, n11141_1, n11127_0, n11120_0, n11106_0, n11091_0, n11077_0, n11070_0, n11060_1, n5858/**/, n5850, n5842, n4874, n4866}), .out(n13663), .config_in(config_chain[31621:31616]), .config_rst(config_rst)); 
buffer_wire buffer_13663 (.in(n13663), .out(n13663_0));
mux15 mux_8498 (.in({n13612_0/**/, n10107_1, n10083_0, n10078_0, n10057_0, n10052_0, n10049_0, n10044_0, n10020_1, n10000_1, n5564, n5556, n5548, n4580, n4572}), .out(n13664), .config_in(config_chain[31627:31622]), .config_rst(config_rst)); 
buffer_wire buffer_13664 (.in(n13664), .out(n13664_0));
mux13 mux_8499 (.in({n13749_1, n11139_1, n11128_0, n11113_0, n11099_0, n11092_0, n11085_0, n11078_0/**/, n11062_1, n5850, n5842, n4874, n4866}), .out(n13665), .config_in(config_chain[31633:31628]), .config_rst(config_rst)); 
buffer_wire buffer_13665 (.in(n13665), .out(n13665_0));
mux15 mux_8500 (.in({n13620_0, n10109_1, n10077_0, n10072_0, n10071_0, n10066_0, n10043_0, n10038_0, n10018_1, n10002_1, n5564, n5556, n5548, n4580/**/, n4572}), .out(n13666), .config_in(config_chain[31639:31634]), .config_rst(config_rst)); 
buffer_wire buffer_13666 (.in(n13666), .out(n13666_0));
mux13 mux_8501 (.in({n13751_1, n11137_1, n11121_0, n11114_0, n11107_0, n11100_0/**/, n11086_0, n11071_0, n11064_1, n5854, n5842, n4874, n4866}), .out(n13667), .config_in(config_chain[31645:31640]), .config_rst(config_rst)); 
buffer_wire buffer_13667 (.in(n13667), .out(n13667_0));
mux15 mux_8502 (.in({n13628_0, n10111_1, n10091_0, n10086_0, n10065_0, n10060_0, n10037_0, n10032_0, n10016_1, n10004_1, n5564/**/, n5556, n5548, n4580, n4572}), .out(n13668), .config_in(config_chain[31651:31646]), .config_rst(config_rst)); 
buffer_wire buffer_13668 (.in(n13668), .out(n13668_0));
mux13 mux_8503 (.in({n13753_1, n11135_1, n11129_0, n11122_0, n11108_0, n11093_0, n11079_0/**/, n11072_0, n11066_1, n5854, n5846, n4874, n4866}), .out(n13669), .config_in(config_chain[31657:31652]), .config_rst(config_rst)); 
buffer_wire buffer_13669 (.in(n13669), .out(n13669_0));
mux15 mux_8504 (.in({n13636_0, n10093_1, n10085_0, n10080_0, n10059_0/**/, n10054_0, n10051_0, n10046_0, n10014_1, n10006_1, n5564, n5556, n5548, n4580, n4572}), .out(n13670), .config_in(config_chain[31663:31658]), .config_rst(config_rst)); 
buffer_wire buffer_13670 (.in(n13670), .out(n13670_0));
mux13 mux_8505 (.in({n13755_1, n11133_1, n11130_0, n11115_0, n11101_0, n11094_0, n11087_0, n11080_0, n11040_1, n5854/**/, n5846, n4878, n4866}), .out(n13671), .config_in(config_chain[31669:31664]), .config_rst(config_rst)); 
buffer_wire buffer_13671 (.in(n13671), .out(n13671_0));
mux16 mux_8506 (.in({n13566_0, n10351_1, n10341_0, n10336_0, n10315_0, n10310_0/**/, n10304_0, n10289_0, n10268_1, n10264_1, n10257_0, n5658, n5650, n4682, n4674, n4666}), .out(n13672), .config_in(config_chain[31675:31670]), .config_rst(config_rst)); 
buffer_wire buffer_13672 (.in(n13672), .out(n13672_0));
mux15 mux_8507 (.in({n13759_0, n11417_1, n11389_0, n11382_0, n11375_1, n11368_0, n11339_0, n11332_0, n11314_1, n11308_1, n5952, n5944, n4976/**/, n4968, n4960}), .out(n13673), .config_in(config_chain[31681:31676]), .config_rst(config_rst)); 
buffer_wire buffer_13673 (.in(n13673), .out(n13673_0));
mux16 mux_8508 (.in({n13574_0, n10353_1, n10335_0, n10330_0, n10324_0, n10309_0, n10303_0/**/, n10298_0, n10286_1, n10266_1, n10259_0, n5658, n5650, n4682, n4674, n4666}), .out(n13674), .config_in(config_chain[31687:31682]), .config_rst(config_rst)); 
buffer_wire buffer_13674 (.in(n13674), .out(n13674_0));
mux15 mux_8509 (.in({n13761_0/**/, n11415_1, n11397_1, n11390_0, n11361_0, n11354_0, n11347_0, n11340_0, n11316_1, n11310_1, n5956, n5944, n4976, n4968, n4960}), .out(n13675), .config_in(config_chain[31693:31688]), .config_rst(config_rst)); 
buffer_wire buffer_13675 (.in(n13675), .out(n13675_0));
mux15 mux_8510 (.in({n13582_0, n10355_1, n10344_0, n10329_0, n10323_0, n10318_0, n10297_0/**/, n10292_0, n10284_1, n10261_0, n5658, n5650, n4682, n4674, n4666}), .out(n13676), .config_in(config_chain[31699:31694]), .config_rst(config_rst)); 
buffer_wire buffer_13676 (.in(n13676), .out(n13676_0));
mux15 mux_8511 (.in({n13763_0, n11413_1, n11383_0, n11376_0, n11369_0/**/, n11362_0, n11348_0, n11333_0, n11318_1, n11309_0, n5956, n5948, n4976, n4968, n4960}), .out(n13677), .config_in(config_chain[31705:31700]), .config_rst(config_rst)); 
buffer_wire buffer_13677 (.in(n13677), .out(n13677_0));
mux15 mux_8512 (.in({n13590_0, n10357_1, n10343_0, n10338_0/**/, n10317_0, n10312_0, n10306_0, n10291_0, n10282_1, n10263_1, n5658, n5650, n4682, n4674, n4666}), .out(n13678), .config_in(config_chain[31711:31706]), .config_rst(config_rst)); 
buffer_wire buffer_13678 (.in(n13678), .out(n13678_0));
mux15 mux_8513 (.in({n13765_0, n11411_1, n11391_0, n11384_0, n11370_0, n11355_0, n11341_0, n11334_0/**/, n11320_1, n11311_0, n5956, n5948, n5940, n4968, n4960}), .out(n13679), .config_in(config_chain[31717:31712]), .config_rst(config_rst)); 
buffer_wire buffer_13679 (.in(n13679), .out(n13679_0));
mux15 mux_8514 (.in({n13598_0, n10359_1, n10337_0/**/, n10332_0, n10326_0, n10311_0, n10305_0, n10300_0, n10280_1, n10265_1, n5658, n5650, n4682, n4674, n4666}), .out(n13680), .config_in(config_chain[31723:31718]), .config_rst(config_rst)); 
buffer_wire buffer_13680 (.in(n13680), .out(n13680_0));
mux14 mux_8515 (.in({n13767_0, n11409_1, n11392_0, n11377_0, n11363_0, n11356_0, n11349_0, n11342_0, n11322_1, n5956/**/, n5948, n5940, n4972, n4960}), .out(n13681), .config_in(config_chain[31729:31724]), .config_rst(config_rst)); 
buffer_wire buffer_13681 (.in(n13681), .out(n13681_0));
mux15 mux_8516 (.in({n13606_0, n10361_1, n10346_0, n10331_0, n10325_0, n10320_0, n10299_0, n10294_0/**/, n10278_1, n10267_1, n5662, n5654, n5646, n4678, n4670}), .out(n13682), .config_in(config_chain[31735:31730]), .config_rst(config_rst)); 
buffer_wire buffer_13682 (.in(n13682), .out(n13682_0));
mux14 mux_8517 (.in({n13769_0, n11407_1, n11385_0, n11378_0/**/, n11371_0, n11364_0, n11350_0, n11335_0, n11324_1, n5956, n5948, n5940, n4972, n4964}), .out(n13683), .config_in(config_chain[31741:31736]), .config_rst(config_rst)); 
buffer_wire buffer_13683 (.in(n13683), .out(n13683_0));
mux15 mux_8518 (.in({n13614_0, n10363_1, n10345_0, n10340_0, n10319_0, n10314_0, n10293_0, n10288_0, n10276_1, n10256_1, n5662, n5654, n5646, n4678/**/, n4670}), .out(n13684), .config_in(config_chain[31747:31742]), .config_rst(config_rst)); 
buffer_wire buffer_13684 (.in(n13684), .out(n13684_0));
mux13 mux_8519 (.in({n13771_0, n11405_1, n11393_0, n11386_0, n11372_0, n11357_0, n11343_0, n11336_0, n11326_1, n5948, n5940, n4972/**/, n4964}), .out(n13685), .config_in(config_chain[31753:31748]), .config_rst(config_rst)); 
buffer_wire buffer_13685 (.in(n13685), .out(n13685_0));
mux15 mux_8520 (.in({n13622_0, n10365_1, n10339_0, n10334_0, n10313_0, n10308_0, n10307_0, n10302_0/**/, n10274_1, n10258_1, n5662, n5654, n5646, n4678, n4670}), .out(n13686), .config_in(config_chain[31759:31754]), .config_rst(config_rst)); 
buffer_wire buffer_13686 (.in(n13686), .out(n13686_0));
mux13 mux_8521 (.in({n13773_0, n11403_1, n11394_0, n11379_0, n11365_0, n11358_0, n11351_0, n11344_0/**/, n11328_1, n5952, n5940, n4972, n4964}), .out(n13687), .config_in(config_chain[31765:31760]), .config_rst(config_rst)); 
buffer_wire buffer_13687 (.in(n13687), .out(n13687_0));
mux15 mux_8522 (.in({n13630_0, n10367_1, n10333_0, n10328_0, n10327_0, n10322_0, n10301_0, n10296_0, n10272_1, n10260_1, n5662, n5654, n5646, n4678/**/, n4670}), .out(n13688), .config_in(config_chain[31771:31766]), .config_rst(config_rst)); 
buffer_wire buffer_13688 (.in(n13688), .out(n13688_0));
mux13 mux_8523 (.in({n13775_0, n11401_1, n11387_0, n11380_0, n11373_0/**/, n11366_0, n11352_0, n11337_0, n11330_1, n5952, n5944, n4972, n4964}), .out(n13689), .config_in(config_chain[31777:31772]), .config_rst(config_rst)); 
buffer_wire buffer_13689 (.in(n13689), .out(n13689_0));
mux15 mux_8524 (.in({n13638_0, n10349_1, n10347_0, n10342_0, n10321_0, n10316_0, n10295_0/**/, n10290_0, n10270_1, n10262_1, n5662, n5654, n5646, n4678, n4670}), .out(n13690), .config_in(config_chain[31783:31778]), .config_rst(config_rst)); 
buffer_wire buffer_13690 (.in(n13690), .out(n13690_0));
mux13 mux_8525 (.in({n13777_0, n11399_1, n11395_0/**/, n11388_0, n11374_0, n11359_0, n11345_0, n11338_0, n11306_1, n5952, n5944, n4976, n4964}), .out(n13691), .config_in(config_chain[31789:31784]), .config_rst(config_rst)); 
buffer_wire buffer_13691 (.in(n13691), .out(n13691_0));
mux15 mux_8526 (.in({n13560_0, n10609_1, n10598_0, n10593_0/**/, n10581_0, n10552_0, n10547_0, n10526_1, n10523_1, n10518_1, n5756, n5748, n4780, n4772, n4764}), .out(n13692), .config_in(config_chain[31795:31790]), .config_rst(config_rst)); 
buffer_wire buffer_13692 (.in(n13692), .out(n13692_0));
mux15 mux_8527 (.in({n13781_0, n11683_1, n11662_0, n11655_0, n11648_0, n11634_0, n11619_1, n11605_0, n11598_0, n11578_1, n6050, n6042, n5074, n5066, n5058/**/}), .out(n13693), .config_in(config_chain[31801:31796]), .config_rst(config_rst)); 
buffer_wire buffer_13693 (.in(n13693), .out(n13693_0));
mux15 mux_8528 (.in({n13568_0, n10611_1, n10601_0, n10572_0, n10567_0, n10560_0, n10555_0/**/, n10525_1, n10520_1, n10514_1, n5760, n5748, n4780, n4772, n4764}), .out(n13694), .config_in(config_chain[31807:31802]), .config_rst(config_rst)); 
buffer_wire buffer_13694 (.in(n13694), .out(n13694_0));
mux15 mux_8529 (.in({n13783_0, n11681_1, n11656_0, n11641_1, n11627_0, n11620_0, n11613_0, n11606_0, n11580_1, n11574_1, n6054, n6042, n5074, n5066, n5058/**/}), .out(n13695), .config_in(config_chain[31813:31808]), .config_rst(config_rst)); 
buffer_wire buffer_13695 (.in(n13695), .out(n13695_0));
mux15 mux_8530 (.in({n13576_0, n10613_1, n10592_0, n10587_0, n10580_0, n10575_0, n10563_0, n10546_0, n10544_1, n10522_1, n5760, n5752, n4780, n4772, n4764/**/}), .out(n13696), .config_in(config_chain[31819:31814]), .config_rst(config_rst)); 
buffer_wire buffer_13696 (.in(n13696), .out(n13696_0));
mux15 mux_8531 (.in({n13785_0, n11679_1, n11663_1, n11649_0, n11642_0, n11635_0, n11628_0, n11614_0, n11599_0, n11582_1, n6054, n6046, n5074, n5066, n5058/**/}), .out(n13697), .config_in(config_chain[31825:31820]), .config_rst(config_rst)); 
buffer_wire buffer_13697 (.in(n13697), .out(n13697_0));
mux15 mux_8532 (.in({n13584_0, n10615_1, n10600_0, n10595_0, n10583_0, n10566_0, n10554_0, n10549_0, n10542_1, n10524_1, n5760, n5752, n5744, n4772, n4764/**/}), .out(n13698), .config_in(config_chain[31831:31826]), .config_rst(config_rst)); 
buffer_wire buffer_13698 (.in(n13698), .out(n13698_0));
mux15 mux_8533 (.in({n13787_0, n11677_1, n11657_0, n11650_0, n11636_0, n11621_0, n11607_0, n11600_0, n11584_1, n11575_0, n6054, n6046/**/, n6038, n5066, n5058}), .out(n13699), .config_in(config_chain[31837:31832]), .config_rst(config_rst)); 
buffer_wire buffer_13699 (.in(n13699), .out(n13699_0));
mux14 mux_8534 (.in({n13592_0/**/, n10617_1, n10603_0, n10586_0, n10574_0, n10569_0, n10562_0, n10557_0, n10540_1, n5760, n5752, n5744, n4776, n4764}), .out(n13700), .config_in(config_chain[31843:31838]), .config_rst(config_rst)); 
buffer_wire buffer_13700 (.in(n13700), .out(n13700_0));
mux14 mux_8535 (.in({n13789_0, n11675_1, n11658_0, n11643_0, n11629_0, n11622_0, n11615_0, n11608_0, n11586_1, n6054/**/, n6046, n6038, n5070, n5058}), .out(n13701), .config_in(config_chain[31849:31844]), .config_rst(config_rst)); 
buffer_wire buffer_13701 (.in(n13701), .out(n13701_0));
mux14 mux_8536 (.in({n13600_0/**/, n10619_1, n10594_0, n10589_0, n10582_0, n10577_0, n10565_0, n10548_0, n10538_1, n5760, n5752, n5744, n4776, n4768}), .out(n13702), .config_in(config_chain[31855:31850]), .config_rst(config_rst)); 
buffer_wire buffer_13702 (.in(n13702), .out(n13702_0));
mux14 mux_8537 (.in({n13791_0, n11673_1, n11651_0, n11644_0, n11637_0, n11630_0, n11616_0/**/, n11601_0, n11588_1, n6054, n6046, n6038, n5070, n5062}), .out(n13703), .config_in(config_chain[31861:31856]), .config_rst(config_rst)); 
buffer_wire buffer_13703 (.in(n13703), .out(n13703_0));
mux13 mux_8538 (.in({n13608_0, n10621_1, n10602_0, n10597_0, n10585_0, n10568_0, n10556_0, n10551_0, n10536_1/**/, n5752, n5744, n4776, n4768}), .out(n13704), .config_in(config_chain[31867:31862]), .config_rst(config_rst)); 
buffer_wire buffer_13704 (.in(n13704), .out(n13704_0));
mux13 mux_8539 (.in({n13793_0, n11671_1, n11659_0, n11652_0, n11638_0, n11623_0, n11609_0, n11602_0, n11590_1, n6046, n6038, n5070, n5062}), .out(n13705), .config_in(config_chain[31873:31868]), .config_rst(config_rst)); 
buffer_wire buffer_13705 (.in(n13705), .out(n13705_0));
mux13 mux_8540 (.in({n13616_0, n10623_1/**/, n10605_0, n10588_0, n10576_0, n10571_0, n10564_0, n10559_0, n10534_1, n5756, n5744, n4776, n4768}), .out(n13706), .config_in(config_chain[31879:31874]), .config_rst(config_rst)); 
buffer_wire buffer_13706 (.in(n13706), .out(n13706_0));
mux13 mux_8541 (.in({n13795_0, n11669_1, n11660_0/**/, n11645_0, n11631_0, n11624_0, n11617_0, n11610_0, n11592_1, n6050, n6038, n5070, n5062}), .out(n13707), .config_in(config_chain[31885:31880]), .config_rst(config_rst)); 
buffer_wire buffer_13707 (.in(n13707), .out(n13707_0));
mux13 mux_8542 (.in({n13624_0/**/, n10625_1, n10596_0, n10591_0, n10584_0, n10579_0, n10550_0, n10532_1, n10517_0, n5756, n5748, n4776, n4768}), .out(n13708), .config_in(config_chain[31891:31886]), .config_rst(config_rst)); 
buffer_wire buffer_13708 (.in(n13708), .out(n13708_0));
mux13 mux_8543 (.in({n13797_0, n11667_1, n11653_0, n11646_0, n11639_0, n11632_0, n11603_0, n11596_1, n11594_1/**/, n6050, n6042, n5070, n5062}), .out(n13709), .config_in(config_chain[31897:31892]), .config_rst(config_rst)); 
buffer_wire buffer_13709 (.in(n13709), .out(n13709_0));
mux13 mux_8544 (.in({n13632_0, n10627_1, n10604_0, n10599_0, n10570_0, n10558_0, n10553_0, n10530_1/**/, n10519_0, n5756, n5748, n4780, n4768}), .out(n13710), .config_in(config_chain[31903:31898]), .config_rst(config_rst)); 
buffer_wire buffer_13710 (.in(n13710), .out(n13710_0));
mux13 mux_8545 (.in({n13799_0, n11665_1/**/, n11661_0, n11654_0, n11625_0, n11618_0, n11611_0, n11604_0, n11572_1, n6050, n6042, n5074, n5062}), .out(n13711), .config_in(config_chain[31909:31904]), .config_rst(config_rst)); 
buffer_wire buffer_13711 (.in(n13711), .out(n13711_0));
mux13 mux_8546 (.in({n13640_0, n10607_1, n10590_0, n10578_0, n10573_0, n10561_0, n10528_1, n10521_0, n10516_1, n5756, n5748, n4780, n4772}), .out(n13712), .config_in(config_chain[31915:31910]), .config_rst(config_rst)); 
buffer_wire buffer_13712 (.in(n13712), .out(n13712_0));
mux3 mux_8547 (.in({n12091_1, n12090_1, n6246}), .out(n13713), .config_in(config_chain[31917:31916]), .config_rst(config_rst)); 
buffer_wire buffer_13713 (.in(n13713), .out(n13713_0));
mux15 mux_8548 (.in({n13562_1, n10871_1, n10852_0, n10847_0, n10838_0, n10833_0, n10821_0, n10786_1/**/, n10783_0, n10778_1, n5854, n5846, n4878, n4870, n4862}), .out(n13714), .config_in(config_chain[31923:31918]), .config_rst(config_rst)); 
buffer_wire buffer_13714 (.in(n13714), .out(n13714_0));
mux15 mux_8549 (.in({n13803_0, n11947_1/**/, n11913_0, n11906_0, n11904_0, n11897_0, n11890_0, n11876_0, n11861_1, n11842_1, n6148, n6140, n5172, n5164, n5156}), .out(n13715), .config_in(config_chain[31929:31924]), .config_rst(config_rst)); 
buffer_wire buffer_13715 (.in(n13715), .out(n13715_0));
mux15 mux_8550 (.in({n13570_1, n10873_1, n10860_0, n10855_0, n10841_0, n10812_0, n10807_0, n10785_1, n10780_1, n10776_1, n5858, n5846, n4878, n4870, n4862}), .out(n13716), .config_in(config_chain[31935:31930]), .config_rst(config_rst)); 
buffer_wire buffer_13716 (.in(n13716), .out(n13716_0));
mux15 mux_8551 (.in({n13805_0, n11945_1, n11926_0, n11921_0, n11914_0, n11898_0/**/, n11883_1, n11869_0, n11862_0, n11844_1, n6152, n6140, n5172, n5164, n5156}), .out(n13717), .config_in(config_chain[31941:31936]), .config_rst(config_rst)); 
buffer_wire buffer_13717 (.in(n13717), .out(n13717_0));
mux15 mux_8552 (.in({n13578_1, n10875_1, n10863_0, n10846_0, n10832_0/**/, n10827_0, n10820_0, n10815_0, n10804_1, n10782_1, n5858, n5850, n4878, n4870, n4862}), .out(n13718), .config_in(config_chain[31947:31942]), .config_rst(config_rst)); 
buffer_wire buffer_13718 (.in(n13718), .out(n13718_0));
mux15 mux_8553 (.in({n13807_0, n11943_1, n11922_0, n11907_0, n11905_1, n11891_0, n11884_0, n11877_0, n11870_0, n11846_1, n6152, n6144, n5172/**/, n5164, n5156}), .out(n13719), .config_in(config_chain[31953:31948]), .config_rst(config_rst)); 
buffer_wire buffer_13719 (.in(n13719), .out(n13719_0));
mux15 mux_8554 (.in({n13586_1, n10877_1, n10854_0, n10849_0, n10840_0, n10835_0/**/, n10823_0, n10806_0, n10802_1, n10784_1, n5858, n5850, n5842, n4870, n4862}), .out(n13720), .config_in(config_chain[31959:31954]), .config_rst(config_rst)); 
buffer_wire buffer_13720 (.in(n13720), .out(n13720_0));
mux15 mux_8555 (.in({n13809_0, n11941_1, n11927_1, n11915_0, n11908_0, n11899_0, n11892_0, n11878_0, n11863_0, n11848_1, n6152, n6144/**/, n6136, n5164, n5156}), .out(n13721), .config_in(config_chain[31965:31960]), .config_rst(config_rst)); 
buffer_wire buffer_13721 (.in(n13721), .out(n13721_0));
mux14 mux_8556 (.in({n13594_1, n10879_1, n10862_0/**/, n10857_0, n10843_0, n10826_0, n10814_0, n10809_0, n10800_1, n5858, n5850, n5842, n4874, n4862}), .out(n13722), .config_in(config_chain[31971:31966]), .config_rst(config_rst)); 
buffer_wire buffer_13722 (.in(n13722), .out(n13722_0));
mux14 mux_8557 (.in({n13811_0, n11939_1, n11923_0, n11916_0, n11900_0, n11885_0, n11871_0, n11864_0, n11850_1, n6152, n6144, n6136, n5168/**/, n5156}), .out(n13723), .config_in(config_chain[31977:31972]), .config_rst(config_rst)); 
buffer_wire buffer_13723 (.in(n13723), .out(n13723_0));
mux14 mux_8558 (.in({n13602_1, n10881_1, n10865_0, n10848_0, n10834_0, n10829_0, n10822_0, n10817_0, n10798_1, n5858, n5850, n5842/**/, n4874, n4866}), .out(n13724), .config_in(config_chain[31983:31978]), .config_rst(config_rst)); 
buffer_wire buffer_13724 (.in(n13724), .out(n13724_0));
mux14 mux_8559 (.in({n13813_0, n11937_1, n11924_0/**/, n11909_0, n11893_0, n11886_0, n11879_0, n11872_0, n11852_1, n6152, n6144, n6136, n5168, n5160}), .out(n13725), .config_in(config_chain[31989:31984]), .config_rst(config_rst)); 
buffer_wire buffer_13725 (.in(n13725), .out(n13725_0));
mux13 mux_8560 (.in({n13610_1, n10883_1, n10856_0, n10851_0, n10842_0, n10837_0, n10825_0, n10808_0/**/, n10796_1, n5850, n5842, n4874, n4866}), .out(n13726), .config_in(config_chain[31995:31990]), .config_rst(config_rst)); 
buffer_wire buffer_13726 (.in(n13726), .out(n13726_0));
mux13 mux_8561 (.in({n13815_0, n11935_1, n11917_0, n11910_0/**/, n11901_0, n11894_0, n11880_0, n11865_0, n11854_1, n6144, n6136, n5168, n5160}), .out(n13727), .config_in(config_chain[32001:31996]), .config_rst(config_rst)); 
buffer_wire buffer_13727 (.in(n13727), .out(n13727_0));
mux13 mux_8562 (.in({n13618_1, n10885_1, n10864_0, n10859_0/**/, n10845_0, n10828_0, n10816_0, n10811_0, n10794_1, n5854, n5842, n4874, n4866}), .out(n13728), .config_in(config_chain[32007:32002]), .config_rst(config_rst)); 
buffer_wire buffer_13728 (.in(n13728), .out(n13728_0));
mux13 mux_8563 (.in({n13817_0, n11933_1, n11925_0, n11918_0/**/, n11902_0, n11887_0, n11873_0, n11866_0, n11856_1, n6148, n6136, n5168, n5160}), .out(n13729), .config_in(config_chain[32013:32008]), .config_rst(config_rst)); 
buffer_wire buffer_13729 (.in(n13729), .out(n13729_0));
mux13 mux_8564 (.in({n13626_1, n10887_1, n10867_1, n10850_0, n10836_0, n10831_0, n10824_0, n10819_0, n10792_1, n5854, n5846, n4874, n4866}), .out(n13730), .config_in(config_chain[32019:32014]), .config_rst(config_rst)); 
buffer_wire buffer_13730 (.in(n13730), .out(n13730_0));
mux13 mux_8565 (.in({n13819_0, n11931_1, n11911_0, n11895_0, n11888_0, n11881_0, n11874_0, n11858_1, n11828_1, n6148/**/, n6140, n5168, n5160}), .out(n13731), .config_in(config_chain[32025:32020]), .config_rst(config_rst)); 
buffer_wire buffer_13731 (.in(n13731), .out(n13731_0));
mux13 mux_8566 (.in({n13634_1, n10889_1, n10858_0, n10853_0, n10844_0, n10839_0, n10810_0, n10790_1/**/, n10779_0, n5854, n5846, n4878, n4866}), .out(n13732), .config_in(config_chain[32031:32026]), .config_rst(config_rst)); 
buffer_wire buffer_13732 (.in(n13732), .out(n13732_0));
mux13 mux_8567 (.in({n13821_0, n11929_1/**/, n11919_0, n11912_0, n11903_0, n11896_0, n11867_0, n11860_1, n11838_1, n6148, n6140, n5172, n5160}), .out(n13733), .config_in(config_chain[32037:32032]), .config_rst(config_rst)); 
buffer_wire buffer_13733 (.in(n13733), .out(n13733_0));
mux13 mux_8568 (.in({n13642_1, n10869_1, n10866_0, n10861_0, n10830_0, n10818_0, n10813_0, n10788_1/**/, n10781_0, n5854, n5846, n4878, n4870}), .out(n13734), .config_in(config_chain[32043:32038]), .config_rst(config_rst)); 
buffer_wire buffer_13734 (.in(n13734), .out(n13734_0));
mux3 mux_8569 (.in({n12093_1, n12092_1, n6246}), .out(n13735), .config_in(config_chain[32045:32044]), .config_rst(config_rst)); 
buffer_wire buffer_13735 (.in(n13735), .out(n13735_0));
mux15 mux_8570 (.in({n13652_1, n11135_1, n11130_0, n11125_0, n11094_0/**/, n11089_0, n11080_0, n11075_0, n11048_1, n11045_0, n5952, n5944, n4976, n4968, n4960}), .out(n13736), .config_in(config_chain[32051:32046]), .config_rst(config_rst)); 
buffer_wire buffer_13736 (.in(n13736), .out(n13736_0));
mux4 mux_8571 (.in({n12191_1/**/, n12102_1, n6250, n5254}), .out(n13737), .config_in(config_chain[32053:32052]), .config_rst(config_rst)); 
buffer_wire buffer_13737 (.in(n13737), .out(n13737_0));
mux15 mux_8572 (.in({n13654_1, n11137_1, n11116_0, n11111_0, n11102_0, n11097_0, n11083_0, n11047_0, n11042_1, n11040_1/**/, n5956, n5944, n4976, n4968, n4960}), .out(n13738), .config_in(config_chain[32059:32054]), .config_rst(config_rst)); 
buffer_wire buffer_13738 (.in(n13738), .out(n13738_0));
mux3 mux_8573 (.in({n12193_1/**/, n12104_1, n5258}), .out(n13739), .config_in(config_chain[32061:32060]), .config_rst(config_rst)); 
buffer_wire buffer_13739 (.in(n13739), .out(n13739_0));
mux15 mux_8574 (.in({n13656_1, n11139_1, n11124_0, n11119_0, n11105_0, n11088_0/**/, n11074_0, n11069_0, n11066_1, n11044_1, n5956, n5948, n4976, n4968, n4960}), .out(n13740), .config_in(config_chain[32067:32062]), .config_rst(config_rst)); 
buffer_wire buffer_13740 (.in(n13740), .out(n13740_0));
mux3 mux_8575 (.in({n12195_1, n12106_1/**/, n5262}), .out(n13741), .config_in(config_chain[32069:32068]), .config_rst(config_rst)); 
buffer_wire buffer_13741 (.in(n13741), .out(n13741_0));
mux15 mux_8576 (.in({n13658_1, n11141_1, n11127_0, n11110_0, n11096_0/**/, n11091_0, n11082_0, n11077_0, n11064_1, n11046_1, n5956, n5948, n5940, n4968, n4960}), .out(n13742), .config_in(config_chain[32075:32070]), .config_rst(config_rst)); 
buffer_wire buffer_13742 (.in(n13742), .out(n13742_0));
mux3 mux_8577 (.in({n12197_1, n12108_1, n5262}), .out(n13743), .config_in(config_chain[32077:32076]), .config_rst(config_rst)); 
buffer_wire buffer_13743 (.in(n13743), .out(n13743_0));
mux14 mux_8578 (.in({n13660_1/**/, n11143_1, n11118_0, n11113_0, n11104_0, n11099_0, n11085_0, n11068_0, n11062_1, n5956, n5948, n5940, n4972, n4960}), .out(n13744), .config_in(config_chain[32083:32078]), .config_rst(config_rst)); 
buffer_wire buffer_13744 (.in(n13744), .out(n13744_0));
mux3 mux_8579 (.in({n12199_1, n12110_1/**/, n5266}), .out(n13745), .config_in(config_chain[32085:32084]), .config_rst(config_rst)); 
buffer_wire buffer_13745 (.in(n13745), .out(n13745_0));
mux14 mux_8580 (.in({n13662_1/**/, n11145_1, n11126_0, n11121_0, n11107_0, n11090_0, n11076_0, n11071_0, n11060_1, n5956, n5948, n5940, n4972, n4964}), .out(n13746), .config_in(config_chain[32091:32086]), .config_rst(config_rst)); 
buffer_wire buffer_13746 (.in(n13746), .out(n13746_0));
mux3 mux_8581 (.in({n12201_1/**/, n12112_1, n5270}), .out(n13747), .config_in(config_chain[32093:32092]), .config_rst(config_rst)); 
buffer_wire buffer_13747 (.in(n13747), .out(n13747_0));
mux13 mux_8582 (.in({n13664_1, n11147_1, n11129_0, n11112_0, n11098_0, n11093_0, n11084_0, n11079_0, n11058_1/**/, n5948, n5940, n4972, n4964}), .out(n13748), .config_in(config_chain[32099:32094]), .config_rst(config_rst)); 
buffer_wire buffer_13748 (.in(n13748), .out(n13748_0));
mux3 mux_8583 (.in({n12203_1, n12114_1/**/, n6234}), .out(n13749), .config_in(config_chain[32101:32100]), .config_rst(config_rst)); 
buffer_wire buffer_13749 (.in(n13749), .out(n13749_0));
mux13 mux_8584 (.in({n13666_1, n11149_1, n11120_0, n11115_0, n11106_0/**/, n11101_0, n11087_0, n11070_0, n11056_1, n5952, n5940, n4972, n4964}), .out(n13750), .config_in(config_chain[32107:32102]), .config_rst(config_rst)); 
buffer_wire buffer_13750 (.in(n13750), .out(n13750_0));
mux3 mux_8585 (.in({n12205_1, n12116_1, n6238/**/}), .out(n13751), .config_in(config_chain[32109:32108]), .config_rst(config_rst)); 
buffer_wire buffer_13751 (.in(n13751), .out(n13751_0));
mux13 mux_8586 (.in({n13668_1, n11151_1, n11128_0, n11123_0, n11109_1, n11092_0, n11078_0/**/, n11073_0, n11054_1, n5952, n5944, n4972, n4964}), .out(n13752), .config_in(config_chain[32115:32110]), .config_rst(config_rst)); 
buffer_wire buffer_13752 (.in(n13752), .out(n13752_0));
mux3 mux_8587 (.in({n12207_1/**/, n12118_1, n6238}), .out(n13753), .config_in(config_chain[32117:32116]), .config_rst(config_rst)); 
buffer_wire buffer_13753 (.in(n13753), .out(n13753_0));
mux13 mux_8588 (.in({n13670_1/**/, n11153_1, n11131_1, n11114_0, n11100_0, n11095_0, n11086_0, n11081_0, n11052_1, n5952, n5944, n4976, n4964}), .out(n13754), .config_in(config_chain[32123:32118]), .config_rst(config_rst)); 
buffer_wire buffer_13754 (.in(n13754), .out(n13754_0));
mux3 mux_8589 (.in({n12209_1, n12120_1/**/, n6242}), .out(n13755), .config_in(config_chain[32125:32124]), .config_rst(config_rst)); 
buffer_wire buffer_13755 (.in(n13755), .out(n13755_0));
mux13 mux_8590 (.in({n13644_1, n11133_1, n11122_0, n11117_0/**/, n11108_0, n11103_0, n11072_0, n11050_1, n11043_0, n5952, n5944, n4976, n4968}), .out(n13756), .config_in(config_chain[32131:32126]), .config_rst(config_rst)); 
buffer_wire buffer_13756 (.in(n13756), .out(n13756_0));
mux3 mux_8591 (.in({n12123_1, n12122_1, n6246}), .out(n13757), .config_in(config_chain[32133:32132]), .config_rst(config_rst)); 
buffer_wire buffer_13757 (.in(n13757), .out(n13757_0));
mux15 mux_8592 (.in({n13672_1/**/, n11401_1, n11388_0, n11383_0, n11374_0, n11369_0, n11338_0, n11333_0, n11312_1, n11309_0, n6050, n6042, n5074, n5066, n5058}), .out(n13758), .config_in(config_chain[32139:32134]), .config_rst(config_rst)); 
buffer_wire buffer_13758 (.in(n13758), .out(n13758_0));
mux4 mux_8593 (.in({n12125_0/**/, n12124_0, n6250, n5254}), .out(n13759), .config_in(config_chain[32141:32140]), .config_rst(config_rst)); 
buffer_wire buffer_13759 (.in(n13759), .out(n13759_0));
mux15 mux_8594 (.in({n13674_1, n11403_1/**/, n11396_0, n11391_0, n11360_0, n11355_0, n11346_0, n11341_0, n11311_0, n11306_1, n6054, n6042, n5074, n5066, n5058}), .out(n13760), .config_in(config_chain[32147:32142]), .config_rst(config_rst)); 
buffer_wire buffer_13760 (.in(n13760), .out(n13760_0));
mux3 mux_8595 (.in({n12127_0/**/, n12126_0, n5258}), .out(n13761), .config_in(config_chain[32149:32148]), .config_rst(config_rst)); 
buffer_wire buffer_13761 (.in(n13761), .out(n13761_0));
mux15 mux_8596 (.in({n13676_1, n11405_1, n11382_0, n11377_0, n11368_0, n11363_0, n11349_0, n11332_0, n11330_1/**/, n11308_1, n6054, n6046, n5074, n5066, n5058}), .out(n13762), .config_in(config_chain[32155:32150]), .config_rst(config_rst)); 
buffer_wire buffer_13762 (.in(n13762), .out(n13762_0));
mux3 mux_8597 (.in({n12129_0, n12128_0/**/, n5262}), .out(n13763), .config_in(config_chain[32157:32156]), .config_rst(config_rst)); 
buffer_wire buffer_13763 (.in(n13763), .out(n13763_0));
mux15 mux_8598 (.in({n13678_1, n11407_1, n11390_0/**/, n11385_0, n11371_0, n11354_0, n11340_0, n11335_0, n11328_1, n11310_1, n6054, n6046, n6038, n5066, n5058}), .out(n13764), .config_in(config_chain[32163:32158]), .config_rst(config_rst)); 
buffer_wire buffer_13764 (.in(n13764), .out(n13764_0));
mux3 mux_8599 (.in({n12131_0, n12130_0, n5266}), .out(n13765), .config_in(config_chain[32165:32164]), .config_rst(config_rst)); 
buffer_wire buffer_13765 (.in(n13765), .out(n13765_0));
mux14 mux_8600 (.in({n13680_1, n11409_1, n11393_0, n11376_0, n11362_0, n11357_0, n11348_0/**/, n11343_0, n11326_1, n6054, n6046, n6038, n5070, n5058}), .out(n13766), .config_in(config_chain[32171:32166]), .config_rst(config_rst)); 
buffer_wire buffer_13766 (.in(n13766), .out(n13766_0));
mux3 mux_8601 (.in({n12133_0, n12132_0/**/, n5266}), .out(n13767), .config_in(config_chain[32173:32172]), .config_rst(config_rst)); 
buffer_wire buffer_13767 (.in(n13767), .out(n13767_0));
mux14 mux_8602 (.in({n13682_1, n11411_1, n11384_0, n11379_0, n11370_0, n11365_0, n11351_0, n11334_0, n11324_1, n6054, n6046, n6038/**/, n5070, n5062}), .out(n13768), .config_in(config_chain[32179:32174]), .config_rst(config_rst)); 
buffer_wire buffer_13768 (.in(n13768), .out(n13768_0));
mux3 mux_8603 (.in({n12135_0, n12134_0, n5270}), .out(n13769), .config_in(config_chain[32181:32180]), .config_rst(config_rst)); 
buffer_wire buffer_13769 (.in(n13769), .out(n13769_0));
mux13 mux_8604 (.in({n13684_1, n11413_1, n11392_0, n11387_0, n11373_0, n11356_0, n11342_0/**/, n11337_0, n11322_1, n6046, n6038, n5070, n5062}), .out(n13770), .config_in(config_chain[32187:32182]), .config_rst(config_rst)); 
buffer_wire buffer_13770 (.in(n13770), .out(n13770_0));
mux3 mux_8605 (.in({n12137_0, n12136_0, n6234}), .out(n13771), .config_in(config_chain[32189:32188]), .config_rst(config_rst)); 
buffer_wire buffer_13771 (.in(n13771), .out(n13771_0));
mux13 mux_8606 (.in({n13686_1, n11415_1, n11395_0, n11378_0, n11364_0, n11359_0, n11350_0, n11345_0/**/, n11320_1, n6050, n6038, n5070, n5062}), .out(n13772), .config_in(config_chain[32195:32190]), .config_rst(config_rst)); 
buffer_wire buffer_13772 (.in(n13772), .out(n13772_0));
mux3 mux_8607 (.in({n12139_0, n12138_0/**/, n6238}), .out(n13773), .config_in(config_chain[32197:32196]), .config_rst(config_rst)); 
buffer_wire buffer_13773 (.in(n13773), .out(n13773_0));
mux13 mux_8608 (.in({n13688_1, n11417_1, n11386_0, n11381_0, n11372_0, n11367_0, n11353_1, n11336_0, n11318_1/**/, n6050, n6042, n5070, n5062}), .out(n13774), .config_in(config_chain[32203:32198]), .config_rst(config_rst)); 
buffer_wire buffer_13774 (.in(n13774), .out(n13774_0));
mux3 mux_8609 (.in({n12141_0, n12140_0, n6242}), .out(n13775), .config_in(config_chain[32205:32204]), .config_rst(config_rst)); 
buffer_wire buffer_13775 (.in(n13775), .out(n13775_0));
mux13 mux_8610 (.in({n13690_1, n11419_1, n11394_0, n11389_0, n11375_1, n11358_0, n11344_0, n11339_0, n11316_1, n6050, n6042/**/, n5074, n5062}), .out(n13776), .config_in(config_chain[32211:32206]), .config_rst(config_rst)); 
buffer_wire buffer_13776 (.in(n13776), .out(n13776_0));
mux3 mux_8611 (.in({n12143_0, n12142_0/**/, n6242}), .out(n13777), .config_in(config_chain[32213:32212]), .config_rst(config_rst)); 
buffer_wire buffer_13777 (.in(n13777), .out(n13777_0));
mux13 mux_8612 (.in({n13646_1, n11399_1, n11397_1, n11380_0, n11366_0, n11361_0, n11352_0, n11347_0, n11314_1, n6050/**/, n6042, n5074, n5066}), .out(n13778), .config_in(config_chain[32219:32214]), .config_rst(config_rst)); 
buffer_wire buffer_13778 (.in(n13778), .out(n13778_0));
mux3 mux_8613 (.in({n12145_1, n12144_0, n6246}), .out(n13779), .config_in(config_chain[32221:32220]), .config_rst(config_rst)); 
buffer_wire buffer_13779 (.in(n13779), .out(n13779_0));
mux15 mux_8614 (.in({n13692_1, n11667_1, n11663_1, n11654_0, n11649_0, n11635_0, n11618_0, n11604_0, n11599_0, n11576_1, n6148, n6140/**/, n5172, n5164, n5156}), .out(n13780), .config_in(config_chain[32227:32222]), .config_rst(config_rst)); 
buffer_wire buffer_13780 (.in(n13780), .out(n13780_0));
mux4 mux_8615 (.in({n12147_0, n12146_0, n6250/**/, n5254}), .out(n13781), .config_in(config_chain[32229:32228]), .config_rst(config_rst)); 
buffer_wire buffer_13781 (.in(n13781), .out(n13781_0));
mux15 mux_8616 (.in({n13694_1, n11669_1, n11657_0, n11640_0, n11626_0, n11621_0, n11612_0, n11607_0/**/, n11575_0, n11572_1, n6152, n6140, n5172, n5164, n5156}), .out(n13782), .config_in(config_chain[32235:32230]), .config_rst(config_rst)); 
buffer_wire buffer_13782 (.in(n13782), .out(n13782_0));
mux3 mux_8617 (.in({n12149_0, n12148_0, n5254}), .out(n13783), .config_in(config_chain[32237:32236]), .config_rst(config_rst)); 
buffer_wire buffer_13783 (.in(n13783), .out(n13783_0));
mux15 mux_8618 (.in({n13696_1, n11671_1, n11662_0, n11648_0, n11643_0, n11634_0, n11629_0/**/, n11615_0, n11598_0, n11594_1, n6152, n6144, n5172, n5164, n5156}), .out(n13784), .config_in(config_chain[32243:32238]), .config_rst(config_rst)); 
buffer_wire buffer_13784 (.in(n13784), .out(n13784_0));
mux3 mux_8619 (.in({n12151_0, n12150_0, n5258}), .out(n13785), .config_in(config_chain[32245:32244]), .config_rst(config_rst)); 
buffer_wire buffer_13785 (.in(n13785), .out(n13785_0));
mux15 mux_8620 (.in({n13698_1, n11673_1, n11656_0, n11651_0, n11637_0, n11620_0, n11606_0, n11601_0/**/, n11592_1, n11574_1, n6152, n6144, n6136, n5164, n5156}), .out(n13786), .config_in(config_chain[32251:32246]), .config_rst(config_rst)); 
buffer_wire buffer_13786 (.in(n13786), .out(n13786_0));
mux3 mux_8621 (.in({n12153_0, n12152_0, n5262}), .out(n13787), .config_in(config_chain[32253:32252]), .config_rst(config_rst)); 
buffer_wire buffer_13787 (.in(n13787), .out(n13787_0));
mux14 mux_8622 (.in({n13700_1, n11675_1, n11659_0, n11642_0, n11628_0, n11623_0, n11614_0, n11609_0, n11590_1, n6152/**/, n6144, n6136, n5168, n5156}), .out(n13788), .config_in(config_chain[32259:32254]), .config_rst(config_rst)); 
buffer_wire buffer_13788 (.in(n13788), .out(n13788_0));
mux3 mux_8623 (.in({n12155_0, n12154_0/**/, n5266}), .out(n13789), .config_in(config_chain[32261:32260]), .config_rst(config_rst)); 
buffer_wire buffer_13789 (.in(n13789), .out(n13789_0));
mux14 mux_8624 (.in({n13702_1/**/, n11677_1, n11650_0, n11645_0, n11636_0, n11631_0, n11617_0, n11600_0, n11588_1, n6152, n6144, n6136, n5168, n5160}), .out(n13790), .config_in(config_chain[32267:32262]), .config_rst(config_rst)); 
buffer_wire buffer_13790 (.in(n13790), .out(n13790_0));
mux3 mux_8625 (.in({n12157_0, n12156_0, n5270}), .out(n13791), .config_in(config_chain[32269:32268]), .config_rst(config_rst)); 
buffer_wire buffer_13791 (.in(n13791), .out(n13791_0));
mux13 mux_8626 (.in({n13704_1, n11679_1, n11658_0, n11653_0, n11639_0, n11622_0, n11608_0, n11603_0, n11586_1, n6144, n6136, n5168, n5160}), .out(n13792), .config_in(config_chain[32275:32270]), .config_rst(config_rst)); 
buffer_wire buffer_13792 (.in(n13792), .out(n13792_0));
mux3 mux_8627 (.in({n12159_0, n12158_0, n5270}), .out(n13793), .config_in(config_chain[32277:32276]), .config_rst(config_rst)); 
buffer_wire buffer_13793 (.in(n13793), .out(n13793_0));
mux13 mux_8628 (.in({n13706_1, n11681_1, n11661_0, n11644_0/**/, n11630_0, n11625_0, n11616_0, n11611_0, n11584_1, n6148, n6136, n5168, n5160}), .out(n13794), .config_in(config_chain[32283:32278]), .config_rst(config_rst)); 
buffer_wire buffer_13794 (.in(n13794), .out(n13794_0));
mux3 mux_8629 (.in({n12161_0, n12160_0, n6234}), .out(n13795), .config_in(config_chain[32285:32284]), .config_rst(config_rst)); 
buffer_wire buffer_13795 (.in(n13795), .out(n13795_0));
mux13 mux_8630 (.in({n13708_1, n11683_1, n11652_0, n11647_0, n11638_0, n11633_0, n11602_0, n11597_1, n11582_1/**/, n6148, n6140, n5168, n5160}), .out(n13796), .config_in(config_chain[32291:32286]), .config_rst(config_rst)); 
buffer_wire buffer_13796 (.in(n13796), .out(n13796_0));
mux3 mux_8631 (.in({n12163_0, n12162_0, n6238}), .out(n13797), .config_in(config_chain[32293:32292]), .config_rst(config_rst)); 
buffer_wire buffer_13797 (.in(n13797), .out(n13797_0));
mux13 mux_8632 (.in({n13710_1, n11685_1, n11660_0, n11655_0, n11624_0, n11619_1, n11610_0, n11605_0, n11580_1, n6148, n6140, n5172, n5160}), .out(n13798), .config_in(config_chain[32299:32294]), .config_rst(config_rst)); 
buffer_wire buffer_13798 (.in(n13798), .out(n13798_0));
mux3 mux_8633 (.in({n12165_0/**/, n12164_0, n6242}), .out(n13799), .config_in(config_chain[32301:32300]), .config_rst(config_rst)); 
buffer_wire buffer_13799 (.in(n13799), .out(n13799_0));
mux13 mux_8634 (.in({n13648_2, n11665_1, n11646_0, n11641_1, n11632_0, n11627_0/**/, n11613_0, n11596_1, n11578_1, n6148, n6140, n5172, n5164}), .out(n13800), .config_in(config_chain[32307:32302]), .config_rst(config_rst)); 
buffer_wire buffer_13800 (.in(n13800), .out(n13800_0));
mux3 mux_8635 (.in({n12167_1, n12166_0, n6246}), .out(n13801), .config_in(config_chain[32309:32308]), .config_rst(config_rst)); 
buffer_wire buffer_13801 (.in(n13801), .out(n13801_0));
mux15 mux_8636 (.in({n13714_1, n11931_1, n11912_0, n11907_0, n11905_1, n11896_0/**/, n11891_0, n11877_0, n11860_1, n11840_1, n6246, n6238, n5270, n5262, n5254}), .out(n13802), .config_in(config_chain[32315:32310]), .config_rst(config_rst)); 
buffer_wire buffer_13802 (.in(n13802), .out(n13802_0));
mux4 mux_8637 (.in({n12169_0, n12168_0, n6250, n5254}), .out(n13803), .config_in(config_chain[32317:32316]), .config_rst(config_rst)); 
buffer_wire buffer_13803 (.in(n13803), .out(n13803_0));
mux15 mux_8638 (.in({n13716_1, n11933_1, n11927_1, n11920_0, n11915_0, n11899_0, n11882_0, n11868_0, n11863_0, n11838_1, n6250, n6238, n5270, n5262, n5254}), .out(n13804), .config_in(config_chain[32323:32318]), .config_rst(config_rst)); 
buffer_wire buffer_13804 (.in(n13804), .out(n13804_0));
mux3 mux_8639 (.in({n12171_0/**/, n12170_0, n5258}), .out(n13805), .config_in(config_chain[32325:32324]), .config_rst(config_rst)); 
buffer_wire buffer_13805 (.in(n13805), .out(n13805_0));
mux15 mux_8640 (.in({n13718_1, n11935_1, n11923_0, n11906_0/**/, n11904_0, n11890_0, n11885_0, n11876_0, n11871_0, n11858_1, n6250, n6242, n5270, n5262, n5254}), .out(n13806), .config_in(config_chain[32331:32326]), .config_rst(config_rst)); 
buffer_wire buffer_13806 (.in(n13806), .out(n13806_0));
mux3 mux_8641 (.in({n12173_0, n12172_0, n5258}), .out(n13807), .config_in(config_chain[32333:32332]), .config_rst(config_rst)); 
buffer_wire buffer_13807 (.in(n13807), .out(n13807_0));
mux15 mux_8642 (.in({n13720_1, n11937_1, n11926_0, n11914_0, n11909_0, n11898_0, n11893_0, n11879_0, n11862_0, n11856_1, n6250, n6242, n6234, n5262, n5254}), .out(n13808), .config_in(config_chain[32339:32334]), .config_rst(config_rst)); 
buffer_wire buffer_13808 (.in(n13808), .out(n13808_0));
mux3 mux_8643 (.in({n12175_0, n12174_0, n5262}), .out(n13809), .config_in(config_chain[32341:32340]), .config_rst(config_rst)); 
buffer_wire buffer_13809 (.in(n13809), .out(n13809_0));
mux14 mux_8644 (.in({n13722_1, n11939_1, n11922_0, n11917_0, n11901_0, n11884_0, n11870_0, n11865_0, n11854_1, n6250, n6242, n6234, n5266, n5254}), .out(n13810), .config_in(config_chain[32347:32342]), .config_rst(config_rst)); 
buffer_wire buffer_13810 (.in(n13810), .out(n13810_0));
mux3 mux_8645 (.in({n12177_0, n12176_0/**/, n5266}), .out(n13811), .config_in(config_chain[32349:32348]), .config_rst(config_rst)); 
buffer_wire buffer_13811 (.in(n13811), .out(n13811_0));
mux14 mux_8646 (.in({n13724_1, n11941_1, n11925_0, n11908_0, n11892_0/**/, n11887_0, n11878_0, n11873_0, n11852_1, n6250, n6242, n6234, n5266, n5258}), .out(n13812), .config_in(config_chain[32355:32350]), .config_rst(config_rst)); 
buffer_wire buffer_13812 (.in(n13812), .out(n13812_0));
mux3 mux_8647 (.in({n12179_0, n12178_0, n5270}), .out(n13813), .config_in(config_chain[32357:32356]), .config_rst(config_rst)); 
buffer_wire buffer_13813 (.in(n13813), .out(n13813_0));
mux13 mux_8648 (.in({n13726_1, n11943_1, n11916_0, n11911_0, n11900_0, n11895_0/**/, n11881_0, n11864_0, n11850_1, n6242, n6234, n5266, n5258}), .out(n13814), .config_in(config_chain[32363:32358]), .config_rst(config_rst)); 
buffer_wire buffer_13814 (.in(n13814), .out(n13814_0));
mux3 mux_8649 (.in({n12181_0, n12180_0, n6234}), .out(n13815), .config_in(config_chain[32365:32364]), .config_rst(config_rst)); 
buffer_wire buffer_13815 (.in(n13815), .out(n13815_0));
mux13 mux_8650 (.in({n13728_1, n11945_1, n11924_0, n11919_0, n11903_0, n11886_0, n11872_0, n11867_0, n11848_1, n6246, n6234, n5266, n5258}), .out(n13816), .config_in(config_chain[32371:32366]), .config_rst(config_rst)); 
buffer_wire buffer_13816 (.in(n13816), .out(n13816_0));
mux3 mux_8651 (.in({n12183_0, n12182_0, n6234}), .out(n13817), .config_in(config_chain[32373:32372]), .config_rst(config_rst)); 
buffer_wire buffer_13817 (.in(n13817), .out(n13817_0));
mux13 mux_8652 (.in({n13730_1, n11947_1, n11910_0, n11894_0, n11889_0/**/, n11880_0, n11875_0, n11846_1, n11829_1, n6246, n6238, n5266, n5258}), .out(n13818), .config_in(config_chain[32379:32374]), .config_rst(config_rst)); 
buffer_wire buffer_13818 (.in(n13818), .out(n13818_0));
mux3 mux_8653 (.in({n12185_0, n12184_0, n6238}), .out(n13819), .config_in(config_chain[32381:32380]), .config_rst(config_rst)); 
buffer_wire buffer_13819 (.in(n13819), .out(n13819_0));
mux13 mux_8654 (.in({n13732_1, n11949_1, n11918_0, n11913_0, n11902_0, n11897_0, n11866_0, n11861_1, n11844_1, n6246, n6238, n5270, n5258}), .out(n13820), .config_in(config_chain[32387:32382]), .config_rst(config_rst)); 
buffer_wire buffer_13820 (.in(n13820), .out(n13820_0));
mux3 mux_8655 (.in({n12187_0, n12186_0, n6242}), .out(n13821), .config_in(config_chain[32389:32388]), .config_rst(config_rst)); 
buffer_wire buffer_13821 (.in(n13821), .out(n13821_0));
mux13 mux_8656 (.in({n13650_2, n11929_1, n11921_0/**/, n11888_0, n11883_1, n11874_0, n11869_0, n11842_1, n11828_1, n6246, n6238, n5270, n5262}), .out(n13822), .config_in(config_chain[32395:32390]), .config_rst(config_rst)); 
buffer_wire buffer_13822 (.in(n13822), .out(n13822_0));
mux3 mux_8657 (.in({n12189_1, n12188_0, n6250}), .out(n13823), .config_in(config_chain[32397:32396]), .config_rst(config_rst)); 
buffer_wire buffer_13823 (.in(n13823), .out(n13823_0));
mux4 mux_8658 (.in({n9819_0/**/, n9818_0, n6444, n5448}), .out(n13824), .config_in(config_chain[32399:32398]), .config_rst(config_rst)); 
buffer_wire buffer_13824 (.in(n13824), .out(n13824_0));
mux15 mux_8659 (.in({n13937_1, n10387_0, n10361_0, n10354_0, n10342_0, n10315_0, n10308_0, n10290_1/**/, n10264_1, n10261_0, n6538, n6530, n5562, n5554, n5546}), .out(n13825), .config_in(config_chain[32405:32400]), .config_rst(config_rst)); 
buffer_wire buffer_13825 (.in(n13825), .out(n13825_0));
mux4 mux_8660 (.in({n9839_0, n9838_0, n6444/**/, n5448}), .out(n13826), .config_in(config_chain[32407:32406]), .config_rst(config_rst)); 
buffer_wire buffer_13826 (.in(n13826), .out(n13826_0));
mux15 mux_8661 (.in({n13959_1, n10647_0, n10613_0, n10606_0, n10599_0, n10592_0, n10580_0, n10548_1, n10522_1, n10519_0, n6636, n6628, n5660, n5652, n5644}), .out(n13827), .config_in(config_chain[32413:32408]), .config_rst(config_rst)); 
buffer_wire buffer_13827 (.in(n13827), .out(n13827_0));
mux4 mux_8662 (.in({n9859_0, n9778_1/**/, n6444, n5448}), .out(n13828), .config_in(config_chain[32415:32414]), .config_rst(config_rst)); 
buffer_wire buffer_13828 (.in(n13828), .out(n13828_0));
mux15 mux_8663 (.in({n13981_1, n10909_0, n10889_0, n10882_0/**/, n10853_0, n10846_0, n10839_0, n10832_0, n10808_1, n10782_1, n6734, n6726, n5758, n5750, n5742}), .out(n13829), .config_in(config_chain[32421:32416]), .config_rst(config_rst)); 
buffer_wire buffer_13829 (.in(n13829), .out(n13829_0));
mux4 mux_8664 (.in({n9799_0/**/, n9798_0, n6444, n5448}), .out(n13830), .config_in(config_chain[32423:32422]), .config_rst(config_rst)); 
buffer_wire buffer_13830 (.in(n13830), .out(n13830_0));
mux16 mux_8665 (.in({n13917_1, n10129_0, n10104_0, n10101_0/**/, n10078_0, n10075_0, n10069_0, n10052_0, n10034_1, n10009_0, n10000_1, n6440, n6432, n5464, n5456, n5448}), .out(n13831), .config_in(config_chain[32429:32424]), .config_rst(config_rst)); 
buffer_wire buffer_13831 (.in(n13831), .out(n13831_0));
mux3 mux_8666 (.in({n9821_0, n9820_0/**/, n5448}), .out(n13832), .config_in(config_chain[32431:32430]), .config_rst(config_rst)); 
buffer_wire buffer_13832 (.in(n13832), .out(n13832_0));
mux15 mux_8667 (.in({n13939_1, n10385_0, n10362_0, n10335_0, n10328_0, n10323_0/**/, n10316_0, n10292_1, n10266_1, n10263_0, n6542, n6530, n5562, n5554, n5546}), .out(n13833), .config_in(config_chain[32437:32432]), .config_rst(config_rst)); 
buffer_wire buffer_13833 (.in(n13833), .out(n13833_0));
mux3 mux_8668 (.in({n9841_0, n9840_0/**/, n5452}), .out(n13834), .config_in(config_chain[32439:32438]), .config_rst(config_rst)); 
buffer_wire buffer_13834 (.in(n13834), .out(n13834_0));
mux15 mux_8669 (.in({n13961_1, n10645_0, n10621_0, n10614_0, n10600_0/**/, n10573_0, n10566_0, n10550_1, n10524_1, n10521_0, n6640, n6628, n5660, n5652, n5644}), .out(n13835), .config_in(config_chain[32445:32440]), .config_rst(config_rst)); 
buffer_wire buffer_13835 (.in(n13835), .out(n13835_0));
mux3 mux_8670 (.in({n9861_0, n9780_1, n5452}), .out(n13836), .config_in(config_chain[32447:32446]), .config_rst(config_rst)); 
buffer_wire buffer_13836 (.in(n13836), .out(n13836_0));
mux15 mux_8671 (.in({n13983_1, n10907_0, n10875_0, n10868_0, n10861_0, n10854_0, n10840_0, n10810_1, n10784_1, n10781_0, n6738, n6726, n5758/**/, n5750, n5742}), .out(n13837), .config_in(config_chain[32453:32448]), .config_rst(config_rst)); 
buffer_wire buffer_13837 (.in(n13837), .out(n13837_0));
mux3 mux_8672 (.in({n9801_0, n9800_0, n5452}), .out(n13838), .config_in(config_chain[32455:32454]), .config_rst(config_rst)); 
buffer_wire buffer_13838 (.in(n13838), .out(n13838_0));
mux16 mux_8673 (.in({n13919_1, n10127_0/**/, n10098_0, n10095_0, n10089_0, n10072_0, n10066_0, n10063_0, n10036_1, n10011_0, n10002_1, n6440, n6432, n5464, n5456, n5448}), .out(n13839), .config_in(config_chain[32461:32456]), .config_rst(config_rst)); 
buffer_wire buffer_13839 (.in(n13839), .out(n13839_0));
mux3 mux_8674 (.in({n9823_0, n9822_0/**/, n5452}), .out(n13840), .config_in(config_chain[32463:32462]), .config_rst(config_rst)); 
buffer_wire buffer_13840 (.in(n13840), .out(n13840_0));
mux15 mux_8675 (.in({n13941_1, n10383_0, n10355_0, n10348_0, n10343_0/**/, n10336_0, n10324_0, n10309_0, n10294_1, n10265_0, n6542, n6534, n5562, n5554, n5546}), .out(n13841), .config_in(config_chain[32469:32464]), .config_rst(config_rst)); 
buffer_wire buffer_13841 (.in(n13841), .out(n13841_0));
mux3 mux_8676 (.in({n9843_0, n9842_0/**/, n5452}), .out(n13842), .config_in(config_chain[32471:32470]), .config_rst(config_rst)); 
buffer_wire buffer_13842 (.in(n13842), .out(n13842_0));
mux15 mux_8677 (.in({n13963_1, n10643_0, n10622_0, n10607_0, n10593_0, n10586_0, n10581_0, n10574_0, n10552_1, n10523_0, n6640/**/, n6632, n5660, n5652, n5644}), .out(n13843), .config_in(config_chain[32477:32472]), .config_rst(config_rst)); 
buffer_wire buffer_13843 (.in(n13843), .out(n13843_0));
mux3 mux_8678 (.in({n9863_0, n9782_1/**/, n5456}), .out(n13844), .config_in(config_chain[32479:32478]), .config_rst(config_rst)); 
buffer_wire buffer_13844 (.in(n13844), .out(n13844_0));
mux15 mux_8679 (.in({n13985_1/**/, n10905_0, n10883_0, n10876_0, n10862_0, n10847_0, n10833_0, n10826_0, n10812_1, n10783_0, n6738, n6730, n5758, n5750, n5742}), .out(n13845), .config_in(config_chain[32485:32480]), .config_rst(config_rst)); 
buffer_wire buffer_13845 (.in(n13845), .out(n13845_0));
mux3 mux_8680 (.in({n9803_0, n9802_0, n5456}), .out(n13846), .config_in(config_chain[32487:32486]), .config_rst(config_rst)); 
buffer_wire buffer_13846 (.in(n13846), .out(n13846_0));
mux15 mux_8681 (.in({n13921_1, n10125_0, n10109_0, n10092_0, n10086_0, n10083_0, n10060_0, n10057_0/**/, n10038_1, n10004_1, n6440, n6432, n5464, n5456, n5448}), .out(n13847), .config_in(config_chain[32493:32488]), .config_rst(config_rst)); 
buffer_wire buffer_13847 (.in(n13847), .out(n13847_0));
mux3 mux_8682 (.in({n9825_0, n9824_0/**/, n5456}), .out(n13848), .config_in(config_chain[32495:32494]), .config_rst(config_rst)); 
buffer_wire buffer_13848 (.in(n13848), .out(n13848_0));
mux15 mux_8683 (.in({n13943_1, n10381_0, n10363_0, n10356_0, n10344_0, n10329_0, n10317_0, n10310_0/**/, n10296_1, n10267_0, n6542, n6534, n6526, n5554, n5546}), .out(n13849), .config_in(config_chain[32501:32496]), .config_rst(config_rst)); 
buffer_wire buffer_13849 (.in(n13849), .out(n13849_0));
mux3 mux_8684 (.in({n9845_0, n9844_0/**/, n5456}), .out(n13850), .config_in(config_chain[32503:32502]), .config_rst(config_rst)); 
buffer_wire buffer_13850 (.in(n13850), .out(n13850_0));
mux15 mux_8685 (.in({n13965_1, n10641_0, n10615_0, n10608_0/**/, n10601_0, n10594_0, n10582_0, n10567_0, n10554_1, n10525_0, n6640, n6632, n6624, n5652, n5644}), .out(n13851), .config_in(config_chain[32509:32504]), .config_rst(config_rst)); 
buffer_wire buffer_13851 (.in(n13851), .out(n13851_0));
mux3 mux_8686 (.in({n9865_0/**/, n9784_1, n5456}), .out(n13852), .config_in(config_chain[32511:32510]), .config_rst(config_rst)); 
buffer_wire buffer_13852 (.in(n13852), .out(n13852_0));
mux15 mux_8687 (.in({n13987_1, n10903_0, n10884_0/**/, n10869_0, n10855_0, n10848_0, n10841_0, n10834_0, n10814_1, n10785_0, n6738, n6730, n6722, n5750, n5742}), .out(n13853), .config_in(config_chain[32517:32512]), .config_rst(config_rst)); 
buffer_wire buffer_13853 (.in(n13853), .out(n13853_0));
mux3 mux_8688 (.in({n9805_0, n9804_0, n5460}), .out(n13854), .config_in(config_chain[32519:32518]), .config_rst(config_rst)); 
buffer_wire buffer_13854 (.in(n13854), .out(n13854_0));
mux15 mux_8689 (.in({n13923_1, n10123_0, n10106_0, n10103_0, n10080_0/**/, n10077_0, n10071_0, n10054_0, n10040_1, n10006_1, n6440, n6432, n5464, n5456, n5448}), .out(n13855), .config_in(config_chain[32525:32520]), .config_rst(config_rst)); 
buffer_wire buffer_13855 (.in(n13855), .out(n13855_0));
mux3 mux_8690 (.in({n9827_0, n9826_0/**/, n5460}), .out(n13856), .config_in(config_chain[32527:32526]), .config_rst(config_rst)); 
buffer_wire buffer_13856 (.in(n13856), .out(n13856_0));
mux14 mux_8691 (.in({n13945_1, n10379_0, n10364_0, n10349_0, n10337_0, n10330_0, n10325_0, n10318_0, n10298_1, n6542/**/, n6534, n6526, n5558, n5546}), .out(n13857), .config_in(config_chain[32533:32528]), .config_rst(config_rst)); 
buffer_wire buffer_13857 (.in(n13857), .out(n13857_0));
mux3 mux_8692 (.in({n9847_0, n9846_0, n5460}), .out(n13858), .config_in(config_chain[32535:32534]), .config_rst(config_rst)); 
buffer_wire buffer_13858 (.in(n13858), .out(n13858_0));
mux14 mux_8693 (.in({n13967_1, n10639_0/**/, n10623_0, n10616_0, n10602_0, n10587_0, n10575_0, n10568_0, n10556_1, n6640, n6632, n6624, n5656, n5644}), .out(n13859), .config_in(config_chain[32541:32536]), .config_rst(config_rst)); 
buffer_wire buffer_13859 (.in(n13859), .out(n13859_0));
mux3 mux_8694 (.in({n9867_0, n9786_1, n5460}), .out(n13860), .config_in(config_chain[32543:32542]), .config_rst(config_rst)); 
buffer_wire buffer_13860 (.in(n13860), .out(n13860_0));
mux14 mux_8695 (.in({n13989_1, n10901_0, n10877_0, n10870_0, n10863_0, n10856_0, n10842_0, n10827_0, n10816_1, n6738, n6730, n6722/**/, n5754, n5742}), .out(n13861), .config_in(config_chain[32549:32544]), .config_rst(config_rst)); 
buffer_wire buffer_13861 (.in(n13861), .out(n13861_0));
mux3 mux_8696 (.in({n9807_0, n9806_0, n5460}), .out(n13862), .config_in(config_chain[32551:32550]), .config_rst(config_rst)); 
buffer_wire buffer_13862 (.in(n13862), .out(n13862_0));
mux15 mux_8697 (.in({n13925_1/**/, n10121_0, n10100_0, n10097_0, n10091_0, n10074_0, n10068_0, n10065_0, n10042_1, n10008_1, n6440, n6432, n5464, n5456, n5448}), .out(n13863), .config_in(config_chain[32557:32552]), .config_rst(config_rst)); 
buffer_wire buffer_13863 (.in(n13863), .out(n13863_0));
mux3 mux_8698 (.in({n9829_0, n9828_0/**/, n5464}), .out(n13864), .config_in(config_chain[32559:32558]), .config_rst(config_rst)); 
buffer_wire buffer_13864 (.in(n13864), .out(n13864_0));
mux14 mux_8699 (.in({n13947_1, n10377_0, n10357_0, n10350_0, n10345_0, n10338_0, n10326_0, n10311_0, n10300_1/**/, n6542, n6534, n6526, n5558, n5550}), .out(n13865), .config_in(config_chain[32565:32560]), .config_rst(config_rst)); 
buffer_wire buffer_13865 (.in(n13865), .out(n13865_0));
mux3 mux_8700 (.in({n9849_0, n9848_0, n5464}), .out(n13866), .config_in(config_chain[32567:32566]), .config_rst(config_rst)); 
buffer_wire buffer_13866 (.in(n13866), .out(n13866_0));
mux14 mux_8701 (.in({n13969_1, n10637_0, n10624_0, n10609_0, n10595_0/**/, n10588_0, n10583_0, n10576_0, n10558_1, n6640, n6632, n6624, n5656, n5648}), .out(n13867), .config_in(config_chain[32573:32568]), .config_rst(config_rst)); 
buffer_wire buffer_13867 (.in(n13867), .out(n13867_0));
mux3 mux_8702 (.in({n9869_0, n9788_1/**/, n5464}), .out(n13868), .config_in(config_chain[32575:32574]), .config_rst(config_rst)); 
buffer_wire buffer_13868 (.in(n13868), .out(n13868_0));
mux14 mux_8703 (.in({n13991_1, n10899_0, n10885_0, n10878_0, n10864_0, n10849_0, n10835_0, n10828_0, n10818_1, n6738/**/, n6730, n6722, n5754, n5746}), .out(n13869), .config_in(config_chain[32581:32576]), .config_rst(config_rst)); 
buffer_wire buffer_13869 (.in(n13869), .out(n13869_0));
mux3 mux_8704 (.in({n9809_0, n9808_0, n5464}), .out(n13870), .config_in(config_chain[32583:32582]), .config_rst(config_rst)); 
buffer_wire buffer_13870 (.in(n13870), .out(n13870_0));
mux15 mux_8705 (.in({n13927_1, n10119_0, n10111_0, n10094_0, n10088_0, n10085_0, n10062_0/**/, n10059_0, n10044_1, n10010_1, n6444, n6436, n6428, n5460, n5452}), .out(n13871), .config_in(config_chain[32589:32584]), .config_rst(config_rst)); 
buffer_wire buffer_13871 (.in(n13871), .out(n13871_0));
mux3 mux_8706 (.in({n9831_0, n9830_0/**/, n5464}), .out(n13872), .config_in(config_chain[32591:32590]), .config_rst(config_rst)); 
buffer_wire buffer_13872 (.in(n13872), .out(n13872_0));
mux13 mux_8707 (.in({n13949_1/**/, n10375_0, n10365_0, n10358_0, n10346_0, n10331_0, n10319_0, n10312_0, n10302_1, n6534, n6526, n5558, n5550}), .out(n13873), .config_in(config_chain[32597:32592]), .config_rst(config_rst)); 
buffer_wire buffer_13873 (.in(n13873), .out(n13873_0));
mux3 mux_8708 (.in({n9851_0, n9850_0, n6428}), .out(n13874), .config_in(config_chain[32599:32598]), .config_rst(config_rst)); 
buffer_wire buffer_13874 (.in(n13874), .out(n13874_0));
mux13 mux_8709 (.in({n13971_1, n10635_0, n10617_0, n10610_0, n10603_0, n10596_0/**/, n10584_0, n10569_0, n10560_1, n6632, n6624, n5656, n5648}), .out(n13875), .config_in(config_chain[32605:32600]), .config_rst(config_rst)); 
buffer_wire buffer_13875 (.in(n13875), .out(n13875_0));
mux3 mux_8710 (.in({n9871_0, n9790_1, n6428}), .out(n13876), .config_in(config_chain[32607:32606]), .config_rst(config_rst)); 
buffer_wire buffer_13876 (.in(n13876), .out(n13876_0));
mux13 mux_8711 (.in({n13993_1, n10897_0, n10886_0, n10871_0, n10857_0, n10850_0, n10843_0, n10836_0, n10820_1, n6730, n6722, n5754, n5746}), .out(n13877), .config_in(config_chain[32613:32608]), .config_rst(config_rst)); 
buffer_wire buffer_13877 (.in(n13877), .out(n13877_0));
mux3 mux_8712 (.in({n9811_0, n9810_0, n6428}), .out(n13878), .config_in(config_chain[32615:32614]), .config_rst(config_rst)); 
buffer_wire buffer_13878 (.in(n13878), .out(n13878_0));
mux15 mux_8713 (.in({n13929_1, n10117_0, n10108_0, n10105_0, n10082_0, n10079_0, n10056_0, n10053_0, n10046_1, n10001_0, n6444, n6436, n6428, n5460, n5452}), .out(n13879), .config_in(config_chain[32621:32616]), .config_rst(config_rst)); 
buffer_wire buffer_13879 (.in(n13879), .out(n13879_0));
mux3 mux_8714 (.in({n9833_0, n9832_0/**/, n6428}), .out(n13880), .config_in(config_chain[32623:32622]), .config_rst(config_rst)); 
buffer_wire buffer_13880 (.in(n13880), .out(n13880_0));
mux13 mux_8715 (.in({n13951_1, n10373_0, n10366_0, n10351_0, n10339_0, n10332_0, n10327_0, n10320_0, n10304_1, n6538/**/, n6526, n5558, n5550}), .out(n13881), .config_in(config_chain[32629:32624]), .config_rst(config_rst)); 
buffer_wire buffer_13881 (.in(n13881), .out(n13881_0));
mux3 mux_8716 (.in({n9853_0/**/, n9852_0, n6428}), .out(n13882), .config_in(config_chain[32631:32630]), .config_rst(config_rst)); 
buffer_wire buffer_13882 (.in(n13882), .out(n13882_0));
mux13 mux_8717 (.in({n13973_1, n10633_0, n10625_0, n10618_0, n10604_0, n10589_0/**/, n10577_0, n10570_0, n10562_1, n6636, n6624, n5656, n5648}), .out(n13883), .config_in(config_chain[32637:32632]), .config_rst(config_rst)); 
buffer_wire buffer_13883 (.in(n13883), .out(n13883_0));
mux3 mux_8718 (.in({n9873_0, n9792_1/**/, n6432}), .out(n13884), .config_in(config_chain[32639:32638]), .config_rst(config_rst)); 
buffer_wire buffer_13884 (.in(n13884), .out(n13884_0));
mux13 mux_8719 (.in({n13995_1, n10895_0, n10879_0, n10872_0, n10865_0, n10858_0, n10844_0/**/, n10829_0, n10822_1, n6734, n6722, n5754, n5746}), .out(n13885), .config_in(config_chain[32645:32640]), .config_rst(config_rst)); 
buffer_wire buffer_13885 (.in(n13885), .out(n13885_0));
mux3 mux_8720 (.in({n9813_0, n9812_0, n6432}), .out(n13886), .config_in(config_chain[32647:32646]), .config_rst(config_rst)); 
buffer_wire buffer_13886 (.in(n13886), .out(n13886_0));
mux15 mux_8721 (.in({n13931_1, n10115_0, n10102_0, n10099_0, n10076_0, n10073_0, n10070_0, n10067_0, n10048_1, n10003_0, n6444, n6436, n6428, n5460, n5452}), .out(n13887), .config_in(config_chain[32653:32648]), .config_rst(config_rst)); 
buffer_wire buffer_13887 (.in(n13887), .out(n13887_0));
mux3 mux_8722 (.in({n9835_0, n9834_0, n6432}), .out(n13888), .config_in(config_chain[32655:32654]), .config_rst(config_rst)); 
buffer_wire buffer_13888 (.in(n13888), .out(n13888_0));
mux13 mux_8723 (.in({n13953_1, n10371_0, n10359_0, n10352_0, n10347_0, n10340_0, n10313_0, n10306_1, n10258_1, n6538, n6530, n5558/**/, n5550}), .out(n13889), .config_in(config_chain[32661:32656]), .config_rst(config_rst)); 
buffer_wire buffer_13889 (.in(n13889), .out(n13889_0));
mux3 mux_8724 (.in({n9855_0, n9854_0/**/, n6432}), .out(n13890), .config_in(config_chain[32663:32662]), .config_rst(config_rst)); 
buffer_wire buffer_13890 (.in(n13890), .out(n13890_0));
mux13 mux_8725 (.in({n13975_1, n10631_0, n10626_0, n10611_0, n10597_0, n10590_0, n10585_0, n10578_0, n10564_1, n6636, n6628, n5656, n5648}), .out(n13891), .config_in(config_chain[32669:32664]), .config_rst(config_rst)); 
buffer_wire buffer_13891 (.in(n13891), .out(n13891_0));
mux3 mux_8726 (.in({n9875_0, n9794_1, n6432}), .out(n13892), .config_in(config_chain[32671:32670]), .config_rst(config_rst)); 
buffer_wire buffer_13892 (.in(n13892), .out(n13892_0));
mux13 mux_8727 (.in({n13997_1, n10893_0, n10887_0, n10880_0, n10866_0, n10851_0, n10837_0, n10830_0, n10824_1, n6734, n6726, n5754, n5746}), .out(n13893), .config_in(config_chain[32677:32672]), .config_rst(config_rst)); 
buffer_wire buffer_13893 (.in(n13893), .out(n13893_0));
mux3 mux_8728 (.in({n9815_0, n9814_0, n6436}), .out(n13894), .config_in(config_chain[32679:32678]), .config_rst(config_rst)); 
buffer_wire buffer_13894 (.in(n13894), .out(n13894_0));
mux15 mux_8729 (.in({n13933_1, n10113_0, n10096_0, n10093_0, n10090_0, n10087_0, n10064_0, n10061_0/**/, n10050_1, n10005_0, n6444, n6436, n6428, n5460, n5452}), .out(n13895), .config_in(config_chain[32685:32680]), .config_rst(config_rst)); 
buffer_wire buffer_13895 (.in(n13895), .out(n13895_0));
mux3 mux_8730 (.in({n9837_0, n9836_0/**/, n6436}), .out(n13896), .config_in(config_chain[32687:32686]), .config_rst(config_rst)); 
buffer_wire buffer_13896 (.in(n13896), .out(n13896_0));
mux13 mux_8731 (.in({n13955_1, n10369_0, n10367_0, n10360_0, n10333_0, n10321_0, n10314_0, n10260_1, n10256_1, n6538, n6530, n5562, n5550/**/}), .out(n13897), .config_in(config_chain[32693:32688]), .config_rst(config_rst)); 
buffer_wire buffer_13897 (.in(n13897), .out(n13897_0));
mux3 mux_8732 (.in({n9857_0, n9856_0/**/, n6436}), .out(n13898), .config_in(config_chain[32695:32694]), .config_rst(config_rst)); 
buffer_wire buffer_13898 (.in(n13898), .out(n13898_0));
mux13 mux_8733 (.in({n13977_1/**/, n10629_0, n10619_0, n10612_0, n10605_0, n10598_0, n10571_0, n10518_1, n10516_1, n6636, n6628, n5660, n5648}), .out(n13899), .config_in(config_chain[32701:32696]), .config_rst(config_rst)); 
buffer_wire buffer_13899 (.in(n13899), .out(n13899_0));
mux3 mux_8734 (.in({n9877_0, n9796_1, n6436}), .out(n13900), .config_in(config_chain[32703:32702]), .config_rst(config_rst)); 
buffer_wire buffer_13900 (.in(n13900), .out(n13900_0));
mux13 mux_8735 (.in({n13999_1, n10891_0/**/, n10888_0, n10873_0, n10859_0, n10852_0, n10845_0, n10838_0, n10778_1, n6734, n6726, n5758, n5746}), .out(n13901), .config_in(config_chain[32709:32704]), .config_rst(config_rst)); 
buffer_wire buffer_13901 (.in(n13901), .out(n13901_0));
mux3 mux_8736 (.in({n9817_0, n9816_0, n6436}), .out(n13902), .config_in(config_chain[32711:32710]), .config_rst(config_rst)); 
buffer_wire buffer_13902 (.in(n13902), .out(n13902_0));
mux15 mux_8737 (.in({n13935_1, n10131_0, n10110_0/**/, n10107_0, n10084_0, n10081_0, n10058_0, n10055_0, n10032_1, n10007_0, n6444, n6436, n6428, n5460, n5452}), .out(n13903), .config_in(config_chain[32717:32712]), .config_rst(config_rst)); 
buffer_wire buffer_13903 (.in(n13903), .out(n13903_0));
mux3 mux_8738 (.in({n9747_0, n9746_1, n6440}), .out(n13904), .config_in(config_chain[32719:32718]), .config_rst(config_rst)); 
buffer_wire buffer_13904 (.in(n13904), .out(n13904_0));
mux13 mux_8739 (.in({n13957_2, n10389_0, n10353_0, n10341_0, n10334_0, n10322_0, n10288_1, n10262_1, n10259_0, n6538, n6530, n5562, n5554}), .out(n13905), .config_in(config_chain[32725:32720]), .config_rst(config_rst)); 
buffer_wire buffer_13905 (.in(n13905), .out(n13905_0));
mux3 mux_8740 (.in({n9749_0, n9748_1, n6440}), .out(n13906), .config_in(config_chain[32727:32726]), .config_rst(config_rst)); 
buffer_wire buffer_13906 (.in(n13906), .out(n13906_0));
mux13 mux_8741 (.in({n13979_1, n10649_0, n10627_0, n10620_0, n10591_0, n10579_0, n10572_0/**/, n10546_1, n10520_1, n6636, n6628, n5660, n5652}), .out(n13907), .config_in(config_chain[32733:32728]), .config_rst(config_rst)); 
buffer_wire buffer_13907 (.in(n13907), .out(n13907_0));
mux3 mux_8742 (.in({n9751_0, n9750_1, n6440}), .out(n13908), .config_in(config_chain[32735:32734]), .config_rst(config_rst)); 
buffer_wire buffer_13908 (.in(n13908), .out(n13908_0));
mux13 mux_8743 (.in({n14001_1, n10911_0, n10881_0, n10874_0, n10867_0, n10860_0, n10831_0, n10806_1/**/, n10780_1, n6734, n6726, n5758, n5750}), .out(n13909), .config_in(config_chain[32741:32736]), .config_rst(config_rst)); 
buffer_wire buffer_13909 (.in(n13909), .out(n13909_0));
mux3 mux_8744 (.in({n9753_0/**/, n9752_1, n6440}), .out(n13910), .config_in(config_chain[32743:32742]), .config_rst(config_rst)); 
buffer_wire buffer_13910 (.in(n13910), .out(n13910_0));
mux13 mux_8745 (.in({n14023_1, n11175_0, n11152_0, n11137_0, n11123_0, n11116_0, n11109_0, n11102_0, n11068_1/**/, n6832, n6824, n5856, n5848}), .out(n13911), .config_in(config_chain[32749:32744]), .config_rst(config_rst)); 
buffer_wire buffer_13911 (.in(n13911), .out(n13911_0));
mux3 mux_8746 (.in({n9755_0, n9754_1, n6440}), .out(n13912), .config_in(config_chain[32751:32750]), .config_rst(config_rst)); 
buffer_wire buffer_13912 (.in(n13912), .out(n13912_0));
mux13 mux_8747 (.in({n14045_0, n11441_0, n11403_0, n11396_0, n11389_0, n11382_0, n11368_0, n11353_0, n11332_1, n6930, n6922/**/, n5954, n5946}), .out(n13913), .config_in(config_chain[32757:32752]), .config_rst(config_rst)); 
buffer_wire buffer_13913 (.in(n13913), .out(n13913_0));
mux3 mux_8748 (.in({n9757_0, n9756_1, n6444}), .out(n13914), .config_in(config_chain[32759:32758]), .config_rst(config_rst)); 
buffer_wire buffer_13914 (.in(n13914), .out(n13914_0));
mux13 mux_8749 (.in({n14067_0, n11707_0, n11678_0/**/, n11647_0, n11640_0, n11633_0, n11626_0, n11598_1, n11597_0, n7028, n7020, n6052, n6044}), .out(n13915), .config_in(config_chain[32765:32760]), .config_rst(config_rst)); 
buffer_wire buffer_13915 (.in(n13915), .out(n13915_0));
mux16 mux_8750 (.in({n13830_0/**/, n10115_0, n10105_0, n10100_0, n10079_0, n10074_0, n10068_0, n10053_0, n10032_1, n10008_1, n10001_0, n6538, n6530, n5562, n5554, n5546}), .out(n13916), .config_in(config_chain[32771:32766]), .config_rst(config_rst)); 
buffer_wire buffer_13916 (.in(n13916), .out(n13916_0));
mux15 mux_8751 (.in({n14003_1, n11173_0, n11145_0, n11138_0, n11131_0, n11124_0, n11095_0, n11088_0, n11070_1, n11044_1, n6832, n6824, n5856, n5848, n5840/**/}), .out(n13917), .config_in(config_chain[32777:32772]), .config_rst(config_rst)); 
buffer_wire buffer_13917 (.in(n13917), .out(n13917_0));
mux16 mux_8752 (.in({n13838_0, n10117_0, n10099_0, n10094_0, n10088_0, n10073_0, n10067_0, n10062_0, n10050_1/**/, n10010_1, n10003_0, n6538, n6530, n5562, n5554, n5546}), .out(n13918), .config_in(config_chain[32783:32778]), .config_rst(config_rst)); 
buffer_wire buffer_13918 (.in(n13918), .out(n13918_0));
mux15 mux_8753 (.in({n14005_1, n11171_0, n11153_0, n11146_0, n11117_0, n11110_0, n11103_0, n11096_0, n11072_1, n11046_1, n6836, n6824, n5856, n5848, n5840/**/}), .out(n13919), .config_in(config_chain[32789:32784]), .config_rst(config_rst)); 
buffer_wire buffer_13919 (.in(n13919), .out(n13919_0));
mux15 mux_8754 (.in({n13846_0, n10119_0, n10108_0/**/, n10093_0, n10087_0, n10082_0, n10061_0, n10056_0, n10048_1, n10005_0, n6538, n6530, n5562, n5554, n5546}), .out(n13920), .config_in(config_chain[32795:32790]), .config_rst(config_rst)); 
buffer_wire buffer_13920 (.in(n13920), .out(n13920_0));
mux15 mux_8755 (.in({n14007_1, n11169_0, n11139_0, n11132_0, n11125_0, n11118_0, n11104_0, n11089_0, n11074_1, n11045_0, n6836, n6828, n5856, n5848, n5840/**/}), .out(n13921), .config_in(config_chain[32801:32796]), .config_rst(config_rst)); 
buffer_wire buffer_13921 (.in(n13921), .out(n13921_0));
mux15 mux_8756 (.in({n13854_0, n10121_0, n10107_0, n10102_0, n10081_0/**/, n10076_0, n10070_0, n10055_0, n10046_1, n10007_0, n6538, n6530, n5562, n5554, n5546}), .out(n13922), .config_in(config_chain[32807:32802]), .config_rst(config_rst)); 
buffer_wire buffer_13922 (.in(n13922), .out(n13922_0));
mux15 mux_8757 (.in({n14009_1, n11167_0, n11147_0, n11140_0, n11126_0, n11111_0, n11097_0, n11090_0, n11076_1, n11047_0, n6836, n6828/**/, n6820, n5848, n5840}), .out(n13923), .config_in(config_chain[32813:32808]), .config_rst(config_rst)); 
buffer_wire buffer_13923 (.in(n13923), .out(n13923_0));
mux15 mux_8758 (.in({n13862_0, n10123_0, n10101_0, n10096_0, n10090_0, n10075_0, n10069_0, n10064_0, n10044_1, n10009_0, n6538/**/, n6530, n5562, n5554, n5546}), .out(n13924), .config_in(config_chain[32819:32814]), .config_rst(config_rst)); 
buffer_wire buffer_13924 (.in(n13924), .out(n13924_0));
mux14 mux_8759 (.in({n14011_1/**/, n11165_0, n11148_0, n11133_0, n11119_0, n11112_0, n11105_0, n11098_0, n11078_1, n6836, n6828, n6820, n5852, n5840}), .out(n13925), .config_in(config_chain[32825:32820]), .config_rst(config_rst)); 
buffer_wire buffer_13925 (.in(n13925), .out(n13925_0));
mux15 mux_8760 (.in({n13870_0, n10125_0, n10110_0, n10095_0, n10089_0, n10084_0, n10063_0, n10058_0, n10042_1, n10011_0, n6542, n6534, n6526, n5558, n5550/**/}), .out(n13926), .config_in(config_chain[32831:32826]), .config_rst(config_rst)); 
buffer_wire buffer_13926 (.in(n13926), .out(n13926_0));
mux14 mux_8761 (.in({n14013_1, n11163_0, n11141_0, n11134_0, n11127_0, n11120_0, n11106_0, n11091_0, n11080_1, n6836, n6828/**/, n6820, n5852, n5844}), .out(n13927), .config_in(config_chain[32837:32832]), .config_rst(config_rst)); 
buffer_wire buffer_13927 (.in(n13927), .out(n13927_0));
mux15 mux_8762 (.in({n13878_0, n10127_0, n10109_0, n10104_0, n10083_0, n10078_0, n10057_0, n10052_0, n10040_1/**/, n10000_1, n6542, n6534, n6526, n5558, n5550}), .out(n13928), .config_in(config_chain[32843:32838]), .config_rst(config_rst)); 
buffer_wire buffer_13928 (.in(n13928), .out(n13928_0));
mux13 mux_8763 (.in({n14015_1, n11161_0, n11149_0, n11142_0, n11128_0, n11113_0, n11099_0/**/, n11092_0, n11082_1, n6828, n6820, n5852, n5844}), .out(n13929), .config_in(config_chain[32849:32844]), .config_rst(config_rst)); 
buffer_wire buffer_13929 (.in(n13929), .out(n13929_0));
mux15 mux_8764 (.in({n13886_0, n10129_0, n10103_0, n10098_0, n10077_0, n10072_0, n10071_0, n10066_0, n10038_1, n10002_1, n6542, n6534, n6526, n5558, n5550/**/}), .out(n13930), .config_in(config_chain[32855:32850]), .config_rst(config_rst)); 
buffer_wire buffer_13930 (.in(n13930), .out(n13930_0));
mux13 mux_8765 (.in({n14017_1, n11159_0, n11150_0, n11135_0, n11121_0, n11114_0, n11107_0, n11100_0, n11084_1, n6832, n6820, n5852/**/, n5844}), .out(n13931), .config_in(config_chain[32861:32856]), .config_rst(config_rst)); 
buffer_wire buffer_13931 (.in(n13931), .out(n13931_0));
mux15 mux_8766 (.in({n13894_0, n10131_0, n10097_0, n10092_0, n10091_0, n10086_0, n10065_0, n10060_0, n10036_1, n10004_1, n6542, n6534, n6526, n5558/**/, n5550}), .out(n13932), .config_in(config_chain[32867:32862]), .config_rst(config_rst)); 
buffer_wire buffer_13932 (.in(n13932), .out(n13932_0));
mux13 mux_8767 (.in({n14019_1, n11157_0/**/, n11143_0, n11136_0, n11129_0, n11122_0, n11108_0, n11093_0, n11086_1, n6832, n6824, n5852, n5844}), .out(n13933), .config_in(config_chain[32873:32868]), .config_rst(config_rst)); 
buffer_wire buffer_13933 (.in(n13933), .out(n13933_0));
mux15 mux_8768 (.in({n13902_0, n10113_0, n10111_0, n10106_0, n10085_0, n10080_0/**/, n10059_0, n10054_0, n10034_1, n10006_1, n6542, n6534, n6526, n5558, n5550}), .out(n13934), .config_in(config_chain[32879:32874]), .config_rst(config_rst)); 
buffer_wire buffer_13934 (.in(n13934), .out(n13934_0));
mux13 mux_8769 (.in({n14021_1, n11155_0, n11151_0, n11144_0, n11130_0, n11115_0, n11101_0, n11094_0, n11042_1, n6832, n6824, n5856/**/, n5844}), .out(n13935), .config_in(config_chain[32885:32880]), .config_rst(config_rst)); 
buffer_wire buffer_13935 (.in(n13935), .out(n13935_0));
mux15 mux_8770 (.in({n13824_0, n10371_0, n10360_0, n10355_0, n10343_0, n10314_0/**/, n10309_0, n10288_1, n10265_0, n10260_1, n6636, n6628, n5660, n5652, n5644}), .out(n13936), .config_in(config_chain[32891:32886]), .config_rst(config_rst)); 
buffer_wire buffer_13936 (.in(n13936), .out(n13936_0));
mux15 mux_8771 (.in({n14025_0/**/, n11439_0, n11418_0, n11411_0, n11404_0, n11390_0, n11375_0, n11361_0, n11354_0, n11334_1, n6930, n6922, n5954, n5946, n5938}), .out(n13937), .config_in(config_chain[32897:32892]), .config_rst(config_rst)); 
buffer_wire buffer_13937 (.in(n13937), .out(n13937_0));
mux15 mux_8772 (.in({n13832_0/**/, n10373_0, n10363_0, n10334_0, n10329_0, n10322_0, n10317_0, n10267_0, n10262_1, n10256_1, n6640, n6628, n5660, n5652, n5644}), .out(n13938), .config_in(config_chain[32903:32898]), .config_rst(config_rst)); 
buffer_wire buffer_13938 (.in(n13938), .out(n13938_0));
mux15 mux_8773 (.in({n14027_0, n11437_0, n11412_0, n11397_0, n11383_0, n11376_0, n11369_0, n11362_0, n11336_1, n11310_1, n6934/**/, n6922, n5954, n5946, n5938}), .out(n13939), .config_in(config_chain[32909:32904]), .config_rst(config_rst)); 
buffer_wire buffer_13939 (.in(n13939), .out(n13939_0));
mux15 mux_8774 (.in({n13840_0, n10375_0, n10354_0, n10349_0, n10342_0, n10337_0, n10325_0, n10308_0, n10306_1, n10264_1, n6640, n6632, n5660/**/, n5652, n5644}), .out(n13940), .config_in(config_chain[32915:32910]), .config_rst(config_rst)); 
buffer_wire buffer_13940 (.in(n13940), .out(n13940_0));
mux15 mux_8775 (.in({n14029_0, n11435_0/**/, n11419_0, n11405_0, n11398_0, n11391_0, n11384_0, n11370_0, n11355_0, n11338_1, n6934, n6926, n5954, n5946, n5938}), .out(n13941), .config_in(config_chain[32921:32916]), .config_rst(config_rst)); 
buffer_wire buffer_13941 (.in(n13941), .out(n13941_0));
mux15 mux_8776 (.in({n13848_0, n10377_0, n10362_0, n10357_0, n10345_0, n10328_0, n10316_0, n10311_0, n10304_1/**/, n10266_1, n6640, n6632, n6624, n5652, n5644}), .out(n13942), .config_in(config_chain[32927:32922]), .config_rst(config_rst)); 
buffer_wire buffer_13942 (.in(n13942), .out(n13942_0));
mux15 mux_8777 (.in({n14031_0/**/, n11433_0, n11413_0, n11406_0, n11392_0, n11377_0, n11363_0, n11356_0, n11340_1, n11311_0, n6934, n6926, n6918, n5946, n5938}), .out(n13943), .config_in(config_chain[32933:32928]), .config_rst(config_rst)); 
buffer_wire buffer_13943 (.in(n13943), .out(n13943_0));
mux14 mux_8778 (.in({n13856_0/**/, n10379_0, n10365_0, n10348_0, n10336_0, n10331_0, n10324_0, n10319_0, n10302_1, n6640, n6632, n6624, n5656, n5644}), .out(n13944), .config_in(config_chain[32939:32934]), .config_rst(config_rst)); 
buffer_wire buffer_13944 (.in(n13944), .out(n13944_0));
mux14 mux_8779 (.in({n14033_0, n11431_0, n11414_0, n11399_0, n11385_0, n11378_0, n11371_0, n11364_0/**/, n11342_1, n6934, n6926, n6918, n5950, n5938}), .out(n13945), .config_in(config_chain[32945:32940]), .config_rst(config_rst)); 
buffer_wire buffer_13945 (.in(n13945), .out(n13945_0));
mux14 mux_8780 (.in({n13864_0/**/, n10381_0, n10356_0, n10351_0, n10344_0, n10339_0, n10327_0, n10310_0, n10300_1, n6640, n6632, n6624, n5656, n5648}), .out(n13946), .config_in(config_chain[32951:32946]), .config_rst(config_rst)); 
buffer_wire buffer_13946 (.in(n13946), .out(n13946_0));
mux14 mux_8781 (.in({n14035_0, n11429_0, n11407_0, n11400_0, n11393_0, n11386_0, n11372_0, n11357_0, n11344_1/**/, n6934, n6926, n6918, n5950, n5942}), .out(n13947), .config_in(config_chain[32957:32952]), .config_rst(config_rst)); 
buffer_wire buffer_13947 (.in(n13947), .out(n13947_0));
mux13 mux_8782 (.in({n13872_0/**/, n10383_0, n10364_0, n10359_0, n10347_0, n10330_0, n10318_0, n10313_0, n10298_1, n6632, n6624, n5656, n5648}), .out(n13948), .config_in(config_chain[32963:32958]), .config_rst(config_rst)); 
buffer_wire buffer_13948 (.in(n13948), .out(n13948_0));
mux13 mux_8783 (.in({n14037_0, n11427_0/**/, n11415_0, n11408_0, n11394_0, n11379_0, n11365_0, n11358_0, n11346_1, n6926, n6918, n5950, n5942}), .out(n13949), .config_in(config_chain[32969:32964]), .config_rst(config_rst)); 
buffer_wire buffer_13949 (.in(n13949), .out(n13949_0));
mux13 mux_8784 (.in({n13880_0/**/, n10385_0, n10367_0, n10350_0, n10338_0, n10333_0, n10326_0, n10321_0, n10296_1, n6636, n6624, n5656, n5648}), .out(n13950), .config_in(config_chain[32975:32970]), .config_rst(config_rst)); 
buffer_wire buffer_13950 (.in(n13950), .out(n13950_0));
mux13 mux_8785 (.in({n14039_0, n11425_0, n11416_0, n11401_0, n11387_0, n11380_0, n11373_0, n11366_0, n11348_1/**/, n6930, n6918, n5950, n5942}), .out(n13951), .config_in(config_chain[32981:32976]), .config_rst(config_rst)); 
buffer_wire buffer_13951 (.in(n13951), .out(n13951_0));
mux13 mux_8786 (.in({n13888_0, n10387_0, n10358_0, n10353_0, n10346_0, n10341_0, n10312_0, n10294_1, n10259_0, n6636, n6628, n5656, n5648}), .out(n13952), .config_in(config_chain[32987:32982]), .config_rst(config_rst)); 
buffer_wire buffer_13952 (.in(n13952), .out(n13952_0));
mux13 mux_8787 (.in({n14041_0, n11423_0, n11409_0, n11402_0, n11395_0, n11388_0, n11359_0, n11352_1, n11350_1, n6930, n6922/**/, n5950, n5942}), .out(n13953), .config_in(config_chain[32993:32988]), .config_rst(config_rst)); 
buffer_wire buffer_13953 (.in(n13953), .out(n13953_0));
mux13 mux_8788 (.in({n13896_0, n10389_0, n10366_0, n10361_0/**/, n10332_0, n10320_0, n10315_0, n10292_1, n10261_0, n6636, n6628, n5660, n5648}), .out(n13954), .config_in(config_chain[32999:32994]), .config_rst(config_rst)); 
buffer_wire buffer_13954 (.in(n13954), .out(n13954_0));
mux13 mux_8789 (.in({n14043_0, n11421_0, n11417_0/**/, n11410_0, n11381_0, n11374_0, n11367_0, n11360_0, n11308_1, n6930, n6922, n5954, n5942}), .out(n13955), .config_in(config_chain[33005:33000]), .config_rst(config_rst)); 
buffer_wire buffer_13955 (.in(n13955), .out(n13955_0));
mux13 mux_8790 (.in({n13904_0, n10369_0, n10352_0, n10340_0/**/, n10335_0, n10323_0, n10290_1, n10263_0, n10258_1, n6636, n6628, n5660, n5652}), .out(n13956), .config_in(config_chain[33011:33006]), .config_rst(config_rst)); 
buffer_wire buffer_13956 (.in(n13956), .out(n13956_0));
mux3 mux_8791 (.in({n12091_0, n12090_1, n7224}), .out(n13957), .config_in(config_chain[33013:33012]), .config_rst(config_rst)); 
buffer_wire buffer_13957 (.in(n13957), .out(n13957_0));
mux15 mux_8792 (.in({n13826_0, n10631_0, n10612_0, n10607_0, n10598_0, n10593_0, n10581_0, n10546_1/**/, n10523_0, n10518_1, n6734, n6726, n5758, n5750, n5742}), .out(n13958), .config_in(config_chain[33019:33014]), .config_rst(config_rst)); 
buffer_wire buffer_13958 (.in(n13958), .out(n13958_0));
mux15 mux_8793 (.in({n14047_0, n11705_0, n11671_0, n11664_0/**/, n11662_0, n11655_0, n11648_0, n11634_0, n11619_0, n11600_1, n7028, n7020, n6052, n6044, n6036}), .out(n13959), .config_in(config_chain[33025:33020]), .config_rst(config_rst)); 
buffer_wire buffer_13959 (.in(n13959), .out(n13959_0));
mux15 mux_8794 (.in({n13834_0, n10633_0, n10620_0, n10615_0, n10601_0, n10572_0, n10567_0/**/, n10525_0, n10520_1, n10516_1, n6738, n6726, n5758, n5750, n5742}), .out(n13960), .config_in(config_chain[33031:33026]), .config_rst(config_rst)); 
buffer_wire buffer_13960 (.in(n13960), .out(n13960_0));
mux15 mux_8795 (.in({n14049_0, n11703_0, n11684_0, n11679_0, n11672_0, n11656_0, n11641_0, n11627_0, n11620_0, n11602_1, n7032/**/, n7020, n6052, n6044, n6036}), .out(n13961), .config_in(config_chain[33037:33032]), .config_rst(config_rst)); 
buffer_wire buffer_13961 (.in(n13961), .out(n13961_0));
mux15 mux_8796 (.in({n13842_0, n10635_0, n10623_0, n10606_0, n10592_0/**/, n10587_0, n10580_0, n10575_0, n10564_1, n10522_1, n6738, n6730, n5758, n5750, n5742}), .out(n13962), .config_in(config_chain[33043:33038]), .config_rst(config_rst)); 
buffer_wire buffer_13962 (.in(n13962), .out(n13962_0));
mux15 mux_8797 (.in({n14051_0/**/, n11701_0, n11680_0, n11665_0, n11663_0, n11649_0, n11642_0, n11635_0, n11628_0, n11604_1, n7032, n7024, n6052, n6044, n6036}), .out(n13963), .config_in(config_chain[33049:33044]), .config_rst(config_rst)); 
buffer_wire buffer_13963 (.in(n13963), .out(n13963_0));
mux15 mux_8798 (.in({n13850_0, n10637_0, n10614_0, n10609_0, n10600_0/**/, n10595_0, n10583_0, n10566_0, n10562_1, n10524_1, n6738, n6730, n6722, n5750, n5742}), .out(n13964), .config_in(config_chain[33055:33050]), .config_rst(config_rst)); 
buffer_wire buffer_13964 (.in(n13964), .out(n13964_0));
mux15 mux_8799 (.in({n14053_0, n11699_0, n11685_0, n11673_0, n11666_0, n11657_0, n11650_0/**/, n11636_0, n11621_0, n11606_1, n7032, n7024, n7016, n6044, n6036}), .out(n13965), .config_in(config_chain[33061:33056]), .config_rst(config_rst)); 
buffer_wire buffer_13965 (.in(n13965), .out(n13965_0));
mux14 mux_8800 (.in({n13858_0, n10639_0, n10622_0, n10617_0, n10603_0, n10586_0, n10574_0, n10569_0, n10560_1, n6738, n6730, n6722/**/, n5754, n5742}), .out(n13966), .config_in(config_chain[33067:33062]), .config_rst(config_rst)); 
buffer_wire buffer_13966 (.in(n13966), .out(n13966_0));
mux14 mux_8801 (.in({n14055_0/**/, n11697_0, n11681_0, n11674_0, n11658_0, n11643_0, n11629_0, n11622_0, n11608_1, n7032, n7024, n7016, n6048, n6036}), .out(n13967), .config_in(config_chain[33073:33068]), .config_rst(config_rst)); 
buffer_wire buffer_13967 (.in(n13967), .out(n13967_0));
mux14 mux_8802 (.in({n13866_0, n10641_0, n10625_0, n10608_0, n10594_0/**/, n10589_0, n10582_0, n10577_0, n10558_1, n6738, n6730, n6722, n5754, n5746}), .out(n13968), .config_in(config_chain[33079:33074]), .config_rst(config_rst)); 
buffer_wire buffer_13968 (.in(n13968), .out(n13968_0));
mux14 mux_8803 (.in({n14057_0/**/, n11695_0, n11682_0, n11667_0, n11651_0, n11644_0, n11637_0, n11630_0, n11610_1, n7032, n7024, n7016, n6048, n6040}), .out(n13969), .config_in(config_chain[33085:33080]), .config_rst(config_rst)); 
buffer_wire buffer_13969 (.in(n13969), .out(n13969_0));
mux13 mux_8804 (.in({n13874_0, n10643_0, n10616_0, n10611_0, n10602_0, n10597_0, n10585_0, n10568_0, n10556_1/**/, n6730, n6722, n5754, n5746}), .out(n13970), .config_in(config_chain[33091:33086]), .config_rst(config_rst)); 
buffer_wire buffer_13970 (.in(n13970), .out(n13970_0));
mux13 mux_8805 (.in({n14059_0, n11693_0, n11675_0, n11668_0, n11659_0, n11652_0, n11638_0, n11623_0, n11612_1, n7024/**/, n7016, n6048, n6040}), .out(n13971), .config_in(config_chain[33097:33092]), .config_rst(config_rst)); 
buffer_wire buffer_13971 (.in(n13971), .out(n13971_0));
mux13 mux_8806 (.in({n13882_0, n10645_0, n10624_0, n10619_0, n10605_0, n10588_0, n10576_0/**/, n10571_0, n10554_1, n6734, n6722, n5754, n5746}), .out(n13972), .config_in(config_chain[33103:33098]), .config_rst(config_rst)); 
buffer_wire buffer_13972 (.in(n13972), .out(n13972_0));
mux13 mux_8807 (.in({n14061_0, n11691_0, n11683_0/**/, n11676_0, n11660_0, n11645_0, n11631_0, n11624_0, n11614_1, n7028, n7016, n6048, n6040}), .out(n13973), .config_in(config_chain[33109:33104]), .config_rst(config_rst)); 
buffer_wire buffer_13973 (.in(n13973), .out(n13973_0));
mux13 mux_8808 (.in({n13890_0, n10647_0, n10627_0, n10610_0, n10596_0, n10591_0, n10584_0, n10579_0/**/, n10552_1, n6734, n6726, n5754, n5746}), .out(n13974), .config_in(config_chain[33115:33110]), .config_rst(config_rst)); 
buffer_wire buffer_13974 (.in(n13974), .out(n13974_0));
mux13 mux_8809 (.in({n14063_0, n11689_0, n11669_0, n11653_0, n11646_0, n11639_0, n11632_0, n11616_1, n11596_1/**/, n7028, n7020, n6048, n6040}), .out(n13975), .config_in(config_chain[33121:33116]), .config_rst(config_rst)); 
buffer_wire buffer_13975 (.in(n13975), .out(n13975_0));
mux13 mux_8810 (.in({n13898_0, n10649_0, n10618_0, n10613_0, n10604_0, n10599_0, n10570_0, n10550_1/**/, n10519_0, n6734, n6726, n5758, n5746}), .out(n13976), .config_in(config_chain[33127:33122]), .config_rst(config_rst)); 
buffer_wire buffer_13976 (.in(n13976), .out(n13976_0));
mux13 mux_8811 (.in({n14065_0, n11687_0/**/, n11677_0, n11670_0, n11661_0, n11654_0, n11625_0, n11618_1, n11574_1, n7028, n7020, n6052, n6040}), .out(n13977), .config_in(config_chain[33133:33128]), .config_rst(config_rst)); 
buffer_wire buffer_13977 (.in(n13977), .out(n13977_0));
mux13 mux_8812 (.in({n13906_0, n10629_0, n10626_0, n10621_0, n10590_0, n10578_0, n10573_0, n10548_1, n10521_0/**/, n6734, n6726, n5758, n5750}), .out(n13978), .config_in(config_chain[33139:33134]), .config_rst(config_rst)); 
buffer_wire buffer_13978 (.in(n13978), .out(n13978_0));
mux3 mux_8813 (.in({n12093_0, n12092_1, n7224}), .out(n13979), .config_in(config_chain[33141:33140]), .config_rst(config_rst)); 
buffer_wire buffer_13979 (.in(n13979), .out(n13979_0));
mux15 mux_8814 (.in({n13828_1, n10893_0, n10888_0, n10883_0, n10852_0, n10847_0/**/, n10838_0, n10833_0, n10806_1, n10783_0, n6832, n6824, n5856, n5848, n5840}), .out(n13980), .config_in(config_chain[33147:33142]), .config_rst(config_rst)); 
buffer_wire buffer_13980 (.in(n13980), .out(n13980_0));
mux16 mux_8815 (.in({n14069_0, n11967_0, n11934_0, n11931_0, n11927_0, n11923_0, n11906_0, n11896_0, n11893_0, n11864_1/**/, n11828_1, n7126, n7118, n6150, n6142, n6134}), .out(n13981), .config_in(config_chain[33153:33148]), .config_rst(config_rst)); 
buffer_wire buffer_13981 (.in(n13981), .out(n13981_0));
mux15 mux_8816 (.in({n13836_1, n10895_0, n10874_0, n10869_0, n10860_0, n10855_0, n10841_0, n10785_0, n10780_1, n10778_1, n6836, n6824, n5856, n5848, n5840/**/}), .out(n13982), .config_in(config_chain[33159:33154]), .config_rst(config_rst)); 
buffer_wire buffer_13982 (.in(n13982), .out(n13982_0));
mux16 mux_8817 (.in({n14071_0, n11965_0, n11949_0, n11945_0/**/, n11928_0, n11920_0, n11917_0, n11890_0, n11887_0, n11866_1, n11860_1, n7126, n7118, n6150, n6142, n6134}), .out(n13983), .config_in(config_chain[33165:33160]), .config_rst(config_rst)); 
buffer_wire buffer_13983 (.in(n13983), .out(n13983_0));
mux15 mux_8818 (.in({n13844_1/**/, n10897_0, n10882_0, n10877_0, n10863_0, n10846_0, n10832_0, n10827_0, n10824_1, n10782_1, n6836, n6828, n5856, n5848, n5840}), .out(n13984), .config_in(config_chain[33171:33166]), .config_rst(config_rst)); 
buffer_wire buffer_13984 (.in(n13984), .out(n13984_0));
mux15 mux_8819 (.in({n14073_0, n11963_0, n11942_0, n11939_0, n11914_0, n11911_0, n11901_0, n11884_0/**/, n11882_1, n11868_1, n7126, n7118, n6150, n6142, n6134}), .out(n13985), .config_in(config_chain[33177:33172]), .config_rst(config_rst)); 
buffer_wire buffer_13985 (.in(n13985), .out(n13985_0));
mux15 mux_8820 (.in({n13852_1, n10899_0, n10885_0, n10868_0, n10854_0, n10849_0, n10840_0, n10835_0, n10822_1, n10784_1, n6836, n6828/**/, n6820, n5848, n5840}), .out(n13986), .config_in(config_chain[33183:33178]), .config_rst(config_rst)); 
buffer_wire buffer_13986 (.in(n13986), .out(n13986_0));
mux15 mux_8821 (.in({n14075_0, n11961_0, n11936_0, n11933_0, n11925_0, n11908_0, n11904_0, n11898_0, n11895_0, n11870_1/**/, n7126, n7118, n6150, n6142, n6134}), .out(n13987), .config_in(config_chain[33189:33184]), .config_rst(config_rst)); 
buffer_wire buffer_13987 (.in(n13987), .out(n13987_0));
mux14 mux_8822 (.in({n13860_1, n10901_0, n10876_0, n10871_0, n10862_0, n10857_0, n10843_0, n10826_0, n10820_1, n6836/**/, n6828, n6820, n5852, n5840}), .out(n13988), .config_in(config_chain[33195:33190]), .config_rst(config_rst)); 
buffer_wire buffer_13988 (.in(n13988), .out(n13988_0));
mux15 mux_8823 (.in({n14077_0, n11959_0, n11947_0, n11930_0, n11926_0/**/, n11922_0, n11919_0, n11892_0, n11889_0, n11872_1, n7126, n7118, n6150, n6142, n6134}), .out(n13989), .config_in(config_chain[33201:33196]), .config_rst(config_rst)); 
buffer_wire buffer_13989 (.in(n13989), .out(n13989_0));
mux14 mux_8824 (.in({n13868_1, n10903_0, n10884_0, n10879_0, n10865_0, n10848_0, n10834_0, n10829_0, n10818_1, n6836, n6828, n6820, n5852, n5844}), .out(n13990), .config_in(config_chain[33207:33202]), .config_rst(config_rst)); 
buffer_wire buffer_13990 (.in(n13990), .out(n13990_0));
mux15 mux_8825 (.in({n14079_0, n11957_0, n11948_0, n11944_0, n11941_0, n11916_0/**/, n11913_0, n11903_0, n11886_0, n11874_1, n7130, n7122, n7114, n6146, n6138}), .out(n13991), .config_in(config_chain[33213:33208]), .config_rst(config_rst)); 
buffer_wire buffer_13991 (.in(n13991), .out(n13991_0));
mux13 mux_8826 (.in({n13876_1, n10905_0/**/, n10887_0, n10870_0, n10856_0, n10851_0, n10842_0, n10837_0, n10816_1, n6828, n6820, n5852, n5844}), .out(n13992), .config_in(config_chain[33219:33214]), .config_rst(config_rst)); 
buffer_wire buffer_13992 (.in(n13992), .out(n13992_0));
mux15 mux_8827 (.in({n14081_0/**/, n11955_0, n11938_0, n11935_0, n11910_0, n11907_0, n11900_0, n11897_0, n11876_1, n11829_0, n7130, n7122, n7114, n6146, n6138}), .out(n13993), .config_in(config_chain[33225:33220]), .config_rst(config_rst)); 
buffer_wire buffer_13993 (.in(n13993), .out(n13993_0));
mux13 mux_8828 (.in({n13884_1, n10907_0, n10878_0, n10873_0, n10864_0, n10859_0/**/, n10845_0, n10828_0, n10814_1, n6832, n6820, n5852, n5844}), .out(n13994), .config_in(config_chain[33231:33226]), .config_rst(config_rst)); 
buffer_wire buffer_13994 (.in(n13994), .out(n13994_0));
mux15 mux_8829 (.in({n14083_0, n11953_0/**/, n11932_0, n11929_0, n11924_0, n11921_0, n11894_0, n11891_0, n11878_1, n11861_0, n7130, n7122, n7114, n6146, n6138}), .out(n13995), .config_in(config_chain[33237:33232]), .config_rst(config_rst)); 
buffer_wire buffer_13995 (.in(n13995), .out(n13995_0));
mux13 mux_8830 (.in({n13892_1, n10909_0, n10886_0, n10881_0, n10867_0, n10850_0, n10836_0, n10831_0, n10812_1, n6832/**/, n6824, n5852, n5844}), .out(n13996), .config_in(config_chain[33243:33238]), .config_rst(config_rst)); 
buffer_wire buffer_13996 (.in(n13996), .out(n13996_0));
mux15 mux_8831 (.in({n14085_0, n11951_0, n11946_0, n11943_0, n11918_0, n11915_0, n11888_0, n11885_0, n11883_0, n11880_1, n7130, n7122, n7114, n6146, n6138}), .out(n13997), .config_in(config_chain[33249:33244]), .config_rst(config_rst)); 
buffer_wire buffer_13997 (.in(n13997), .out(n13997_0));
mux13 mux_8832 (.in({n13900_1, n10911_0, n10889_0, n10872_0, n10858_0, n10853_0, n10844_0, n10839_0, n10810_1, n6832, n6824, n5856, n5844/**/}), .out(n13998), .config_in(config_chain[33255:33250]), .config_rst(config_rst)); 
buffer_wire buffer_13998 (.in(n13998), .out(n13998_0));
mux15 mux_8833 (.in({n14087_0, n11969_0, n11940_0, n11937_0, n11912_0, n11909_0, n11905_0, n11902_0, n11899_0, n11862_1, n7130, n7122, n7114, n6146, n6138/**/}), .out(n13999), .config_in(config_chain[33261:33256]), .config_rst(config_rst)); 
buffer_wire buffer_13999 (.in(n13999), .out(n13999_0));
mux13 mux_8834 (.in({n13908_1, n10891_0, n10880_0, n10875_0, n10866_0, n10861_0/**/, n10830_0, n10808_1, n10781_0, n6832, n6824, n5856, n5848}), .out(n14000), .config_in(config_chain[33267:33262]), .config_rst(config_rst)); 
buffer_wire buffer_14000 (.in(n14000), .out(n14000_0));
mux3 mux_8835 (.in({n12123_0, n12122_1, n7224}), .out(n14001), .config_in(config_chain[33269:33268]), .config_rst(config_rst)); 
buffer_wire buffer_14001 (.in(n14001), .out(n14001_0));
mux15 mux_8836 (.in({n13916_1, n11157_0, n11144_0, n11139_0, n11130_0, n11125_0, n11094_0, n11089_0, n11068_1, n11045_0, n6930, n6922/**/, n5954, n5946, n5938}), .out(n14002), .config_in(config_chain[33275:33270]), .config_rst(config_rst)); 
buffer_wire buffer_14002 (.in(n14002), .out(n14002_0));
mux4 mux_8837 (.in({n12211_0, n12124_1/**/, n7228, n6232}), .out(n14003), .config_in(config_chain[33277:33276]), .config_rst(config_rst)); 
buffer_wire buffer_14003 (.in(n14003), .out(n14003_0));
mux15 mux_8838 (.in({n13918_1, n11159_0, n11152_0, n11147_0, n11116_0, n11111_0, n11102_0, n11097_0/**/, n11047_0, n11042_1, n6934, n6922, n5954, n5946, n5938}), .out(n14004), .config_in(config_chain[33283:33278]), .config_rst(config_rst)); 
buffer_wire buffer_14004 (.in(n14004), .out(n14004_0));
mux3 mux_8839 (.in({n12213_0, n12126_1/**/, n6236}), .out(n14005), .config_in(config_chain[33285:33284]), .config_rst(config_rst)); 
buffer_wire buffer_14005 (.in(n14005), .out(n14005_0));
mux15 mux_8840 (.in({n13920_1, n11161_0, n11138_0, n11133_0, n11124_0, n11119_0, n11105_0, n11088_0, n11086_1, n11044_1, n6934, n6926, n5954/**/, n5946, n5938}), .out(n14006), .config_in(config_chain[33291:33286]), .config_rst(config_rst)); 
buffer_wire buffer_14006 (.in(n14006), .out(n14006_0));
mux3 mux_8841 (.in({n12215_0, n12128_1/**/, n6240}), .out(n14007), .config_in(config_chain[33293:33292]), .config_rst(config_rst)); 
buffer_wire buffer_14007 (.in(n14007), .out(n14007_0));
mux15 mux_8842 (.in({n13922_1, n11163_0, n11146_0, n11141_0, n11127_0, n11110_0, n11096_0, n11091_0, n11084_1/**/, n11046_1, n6934, n6926, n6918, n5946, n5938}), .out(n14008), .config_in(config_chain[33299:33294]), .config_rst(config_rst)); 
buffer_wire buffer_14008 (.in(n14008), .out(n14008_0));
mux3 mux_8843 (.in({n12217_0, n12130_1/**/, n6244}), .out(n14009), .config_in(config_chain[33301:33300]), .config_rst(config_rst)); 
buffer_wire buffer_14009 (.in(n14009), .out(n14009_0));
mux14 mux_8844 (.in({n13924_1, n11165_0, n11149_0/**/, n11132_0, n11118_0, n11113_0, n11104_0, n11099_0, n11082_1, n6934, n6926, n6918, n5950, n5938}), .out(n14010), .config_in(config_chain[33307:33302]), .config_rst(config_rst)); 
buffer_wire buffer_14010 (.in(n14010), .out(n14010_0));
mux3 mux_8845 (.in({n12219_0, n12132_1/**/, n6244}), .out(n14011), .config_in(config_chain[33309:33308]), .config_rst(config_rst)); 
buffer_wire buffer_14011 (.in(n14011), .out(n14011_0));
mux14 mux_8846 (.in({n13926_1, n11167_0, n11140_0, n11135_0, n11126_0, n11121_0, n11107_0/**/, n11090_0, n11080_1, n6934, n6926, n6918, n5950, n5942}), .out(n14012), .config_in(config_chain[33315:33310]), .config_rst(config_rst)); 
buffer_wire buffer_14012 (.in(n14012), .out(n14012_0));
mux3 mux_8847 (.in({n12221_0, n12134_1, n6248}), .out(n14013), .config_in(config_chain[33317:33316]), .config_rst(config_rst)); 
buffer_wire buffer_14013 (.in(n14013), .out(n14013_0));
mux13 mux_8848 (.in({n13928_1, n11169_0/**/, n11148_0, n11143_0, n11129_0, n11112_0, n11098_0, n11093_0, n11078_1, n6926, n6918, n5950, n5942}), .out(n14014), .config_in(config_chain[33323:33318]), .config_rst(config_rst)); 
buffer_wire buffer_14014 (.in(n14014), .out(n14014_0));
mux3 mux_8849 (.in({n12223_0, n12136_1, n7212}), .out(n14015), .config_in(config_chain[33325:33324]), .config_rst(config_rst)); 
buffer_wire buffer_14015 (.in(n14015), .out(n14015_0));
mux13 mux_8850 (.in({n13930_1, n11171_0, n11151_0, n11134_0, n11120_0, n11115_0, n11106_0, n11101_0, n11076_1, n6930/**/, n6918, n5950, n5942}), .out(n14016), .config_in(config_chain[33331:33326]), .config_rst(config_rst)); 
buffer_wire buffer_14016 (.in(n14016), .out(n14016_0));
mux3 mux_8851 (.in({n12225_0, n12138_1/**/, n7216}), .out(n14017), .config_in(config_chain[33333:33332]), .config_rst(config_rst)); 
buffer_wire buffer_14017 (.in(n14017), .out(n14017_0));
mux13 mux_8852 (.in({n13932_1, n11173_0, n11142_0, n11137_0, n11128_0, n11123_0, n11109_0, n11092_0, n11074_1/**/, n6930, n6922, n5950, n5942}), .out(n14018), .config_in(config_chain[33339:33334]), .config_rst(config_rst)); 
buffer_wire buffer_14018 (.in(n14018), .out(n14018_0));
mux3 mux_8853 (.in({n12227_0, n12140_1, n7220}), .out(n14019), .config_in(config_chain[33341:33340]), .config_rst(config_rst)); 
buffer_wire buffer_14019 (.in(n14019), .out(n14019_0));
mux13 mux_8854 (.in({n13934_1, n11175_0, n11150_0, n11145_0, n11131_0, n11114_0, n11100_0, n11095_0/**/, n11072_1, n6930, n6922, n5954, n5942}), .out(n14020), .config_in(config_chain[33347:33342]), .config_rst(config_rst)); 
buffer_wire buffer_14020 (.in(n14020), .out(n14020_0));
mux3 mux_8855 (.in({n12229_0, n12142_1, n7220}), .out(n14021), .config_in(config_chain[33349:33348]), .config_rst(config_rst)); 
buffer_wire buffer_14021 (.in(n14021), .out(n14021_0));
mux13 mux_8856 (.in({n13910_1, n11155_0, n11153_0, n11136_0, n11122_0, n11117_0, n11108_0, n11103_0, n11070_1, n6930, n6922/**/, n5954, n5946}), .out(n14022), .config_in(config_chain[33355:33350]), .config_rst(config_rst)); 
buffer_wire buffer_14022 (.in(n14022), .out(n14022_0));
mux3 mux_8857 (.in({n12145_0, n12144_1, n7224}), .out(n14023), .config_in(config_chain[33357:33356]), .config_rst(config_rst)); 
buffer_wire buffer_14023 (.in(n14023), .out(n14023_0));
mux15 mux_8858 (.in({n13936_1/**/, n11423_0, n11419_0, n11410_0, n11405_0, n11391_0, n11374_0, n11360_0, n11355_0, n11332_1, n7028, n7020, n6052, n6044, n6036}), .out(n14024), .config_in(config_chain[33363:33358]), .config_rst(config_rst)); 
buffer_wire buffer_14024 (.in(n14024), .out(n14024_0));
mux4 mux_8859 (.in({n12147_0, n12146_0, n7228/**/, n6232}), .out(n14025), .config_in(config_chain[33365:33364]), .config_rst(config_rst)); 
buffer_wire buffer_14025 (.in(n14025), .out(n14025_0));
mux15 mux_8860 (.in({n13938_1/**/, n11425_0, n11413_0, n11396_0, n11382_0, n11377_0, n11368_0, n11363_0, n11311_0, n11308_1, n7032, n7020, n6052, n6044, n6036}), .out(n14026), .config_in(config_chain[33371:33366]), .config_rst(config_rst)); 
buffer_wire buffer_14026 (.in(n14026), .out(n14026_0));
mux3 mux_8861 (.in({n12149_0, n12148_0, n6232}), .out(n14027), .config_in(config_chain[33373:33372]), .config_rst(config_rst)); 
buffer_wire buffer_14027 (.in(n14027), .out(n14027_0));
mux15 mux_8862 (.in({n13940_1, n11427_0, n11418_0, n11404_0, n11399_0, n11390_0, n11385_0, n11371_0, n11354_0, n11350_1, n7032, n7024, n6052, n6044, n6036/**/}), .out(n14028), .config_in(config_chain[33379:33374]), .config_rst(config_rst)); 
buffer_wire buffer_14028 (.in(n14028), .out(n14028_0));
mux3 mux_8863 (.in({n12151_0, n12150_0/**/, n6236}), .out(n14029), .config_in(config_chain[33381:33380]), .config_rst(config_rst)); 
buffer_wire buffer_14029 (.in(n14029), .out(n14029_0));
mux15 mux_8864 (.in({n13942_1, n11429_0, n11412_0, n11407_0, n11393_0, n11376_0, n11362_0, n11357_0, n11348_1/**/, n11310_1, n7032, n7024, n7016, n6044, n6036}), .out(n14030), .config_in(config_chain[33387:33382]), .config_rst(config_rst)); 
buffer_wire buffer_14030 (.in(n14030), .out(n14030_0));
mux3 mux_8865 (.in({n12153_0, n12152_0/**/, n6240}), .out(n14031), .config_in(config_chain[33389:33388]), .config_rst(config_rst)); 
buffer_wire buffer_14031 (.in(n14031), .out(n14031_0));
mux14 mux_8866 (.in({n13944_1/**/, n11431_0, n11415_0, n11398_0, n11384_0, n11379_0, n11370_0, n11365_0, n11346_1, n7032, n7024, n7016, n6048, n6036}), .out(n14032), .config_in(config_chain[33395:33390]), .config_rst(config_rst)); 
buffer_wire buffer_14032 (.in(n14032), .out(n14032_0));
mux3 mux_8867 (.in({n12155_0, n12154_0, n6244}), .out(n14033), .config_in(config_chain[33397:33396]), .config_rst(config_rst)); 
buffer_wire buffer_14033 (.in(n14033), .out(n14033_0));
mux14 mux_8868 (.in({n13946_1/**/, n11433_0, n11406_0, n11401_0, n11392_0, n11387_0, n11373_0, n11356_0, n11344_1, n7032, n7024, n7016, n6048, n6040}), .out(n14034), .config_in(config_chain[33403:33398]), .config_rst(config_rst)); 
buffer_wire buffer_14034 (.in(n14034), .out(n14034_0));
mux3 mux_8869 (.in({n12157_0, n12156_0, n6248}), .out(n14035), .config_in(config_chain[33405:33404]), .config_rst(config_rst)); 
buffer_wire buffer_14035 (.in(n14035), .out(n14035_0));
mux13 mux_8870 (.in({n13948_1/**/, n11435_0, n11414_0, n11409_0, n11395_0, n11378_0, n11364_0, n11359_0, n11342_1, n7024, n7016, n6048, n6040}), .out(n14036), .config_in(config_chain[33411:33406]), .config_rst(config_rst)); 
buffer_wire buffer_14036 (.in(n14036), .out(n14036_0));
mux3 mux_8871 (.in({n12159_0, n12158_0/**/, n6248}), .out(n14037), .config_in(config_chain[33413:33412]), .config_rst(config_rst)); 
buffer_wire buffer_14037 (.in(n14037), .out(n14037_0));
mux13 mux_8872 (.in({n13950_1/**/, n11437_0, n11417_0, n11400_0, n11386_0, n11381_0, n11372_0, n11367_0, n11340_1, n7028, n7016, n6048, n6040}), .out(n14038), .config_in(config_chain[33419:33414]), .config_rst(config_rst)); 
buffer_wire buffer_14038 (.in(n14038), .out(n14038_0));
mux3 mux_8873 (.in({n12161_0, n12160_0, n7212}), .out(n14039), .config_in(config_chain[33421:33420]), .config_rst(config_rst)); 
buffer_wire buffer_14039 (.in(n14039), .out(n14039_0));
mux13 mux_8874 (.in({n13952_1, n11439_0, n11408_0, n11403_0, n11394_0, n11389_0, n11358_0, n11353_0, n11338_1, n7028/**/, n7020, n6048, n6040}), .out(n14040), .config_in(config_chain[33427:33422]), .config_rst(config_rst)); 
buffer_wire buffer_14040 (.in(n14040), .out(n14040_0));
mux3 mux_8875 (.in({n12163_0/**/, n12162_0, n7216}), .out(n14041), .config_in(config_chain[33429:33428]), .config_rst(config_rst)); 
buffer_wire buffer_14041 (.in(n14041), .out(n14041_0));
mux13 mux_8876 (.in({n13954_1, n11441_0, n11416_0, n11411_0, n11380_0, n11375_0, n11366_0, n11361_0, n11336_1, n7028, n7020, n6052, n6040}), .out(n14042), .config_in(config_chain[33435:33430]), .config_rst(config_rst)); 
buffer_wire buffer_14042 (.in(n14042), .out(n14042_0));
mux3 mux_8877 (.in({n12165_0, n12164_0/**/, n7220}), .out(n14043), .config_in(config_chain[33437:33436]), .config_rst(config_rst)); 
buffer_wire buffer_14043 (.in(n14043), .out(n14043_0));
mux13 mux_8878 (.in({n13912_1, n11421_0, n11402_0/**/, n11397_0, n11388_0, n11383_0, n11369_0, n11352_1, n11334_1, n7028, n7020, n6052, n6044}), .out(n14044), .config_in(config_chain[33443:33438]), .config_rst(config_rst)); 
buffer_wire buffer_14044 (.in(n14044), .out(n14044_0));
mux3 mux_8879 (.in({n12167_0, n12166_0, n7224}), .out(n14045), .config_in(config_chain[33445:33444]), .config_rst(config_rst)); 
buffer_wire buffer_14045 (.in(n14045), .out(n14045_0));
mux15 mux_8880 (.in({n13958_1, n11689_0, n11670_0/**/, n11665_0, n11663_0, n11654_0, n11649_0, n11635_0, n11618_1, n11598_1, n7126, n7118, n6150, n6142, n6134}), .out(n14046), .config_in(config_chain[33451:33446]), .config_rst(config_rst)); 
buffer_wire buffer_14046 (.in(n14046), .out(n14046_0));
mux4 mux_8881 (.in({n12169_0, n12168_0/**/, n7228, n6232}), .out(n14047), .config_in(config_chain[33453:33452]), .config_rst(config_rst)); 
buffer_wire buffer_14047 (.in(n14047), .out(n14047_0));
mux15 mux_8882 (.in({n13960_1, n11691_0, n11685_0, n11678_0, n11673_0/**/, n11657_0, n11640_0, n11626_0, n11621_0, n11574_1, n7130, n7118, n6150, n6142, n6134}), .out(n14048), .config_in(config_chain[33459:33454]), .config_rst(config_rst)); 
buffer_wire buffer_14048 (.in(n14048), .out(n14048_0));
mux3 mux_8883 (.in({n12171_0, n12170_0/**/, n6236}), .out(n14049), .config_in(config_chain[33461:33460]), .config_rst(config_rst)); 
buffer_wire buffer_14049 (.in(n14049), .out(n14049_0));
mux15 mux_8884 (.in({n13962_1, n11693_0, n11681_0, n11664_0, n11662_0, n11648_0, n11643_0, n11634_0, n11629_0, n11616_1, n7130, n7122, n6150/**/, n6142, n6134}), .out(n14050), .config_in(config_chain[33467:33462]), .config_rst(config_rst)); 
buffer_wire buffer_14050 (.in(n14050), .out(n14050_0));
mux3 mux_8885 (.in({n12173_0, n12172_0/**/, n6236}), .out(n14051), .config_in(config_chain[33469:33468]), .config_rst(config_rst)); 
buffer_wire buffer_14051 (.in(n14051), .out(n14051_0));
mux15 mux_8886 (.in({n13964_1, n11695_0, n11684_0, n11672_0, n11667_0, n11656_0, n11651_0, n11637_0, n11620_0, n11614_1, n7130/**/, n7122, n7114, n6142, n6134}), .out(n14052), .config_in(config_chain[33475:33470]), .config_rst(config_rst)); 
buffer_wire buffer_14052 (.in(n14052), .out(n14052_0));
mux3 mux_8887 (.in({n12175_0/**/, n12174_0, n6240}), .out(n14053), .config_in(config_chain[33477:33476]), .config_rst(config_rst)); 
buffer_wire buffer_14053 (.in(n14053), .out(n14053_0));
mux14 mux_8888 (.in({n13966_1, n11697_0, n11680_0, n11675_0, n11659_0, n11642_0, n11628_0/**/, n11623_0, n11612_1, n7130, n7122, n7114, n6146, n6134}), .out(n14054), .config_in(config_chain[33483:33478]), .config_rst(config_rst)); 
buffer_wire buffer_14054 (.in(n14054), .out(n14054_0));
mux3 mux_8889 (.in({n12177_0, n12176_0/**/, n6244}), .out(n14055), .config_in(config_chain[33485:33484]), .config_rst(config_rst)); 
buffer_wire buffer_14055 (.in(n14055), .out(n14055_0));
mux14 mux_8890 (.in({n13968_1, n11699_0, n11683_0, n11666_0, n11650_0, n11645_0, n11636_0, n11631_0, n11610_1/**/, n7130, n7122, n7114, n6146, n6138}), .out(n14056), .config_in(config_chain[33491:33486]), .config_rst(config_rst)); 
buffer_wire buffer_14056 (.in(n14056), .out(n14056_0));
mux3 mux_8891 (.in({n12179_0, n12178_0/**/, n6248}), .out(n14057), .config_in(config_chain[33493:33492]), .config_rst(config_rst)); 
buffer_wire buffer_14057 (.in(n14057), .out(n14057_0));
mux13 mux_8892 (.in({n13970_1, n11701_0, n11674_0, n11669_0/**/, n11658_0, n11653_0, n11639_0, n11622_0, n11608_1, n7122, n7114, n6146, n6138}), .out(n14058), .config_in(config_chain[33499:33494]), .config_rst(config_rst)); 
buffer_wire buffer_14058 (.in(n14058), .out(n14058_0));
mux3 mux_8893 (.in({n12181_0, n12180_0, n7212}), .out(n14059), .config_in(config_chain[33501:33500]), .config_rst(config_rst)); 
buffer_wire buffer_14059 (.in(n14059), .out(n14059_0));
mux13 mux_8894 (.in({n13972_1, n11703_0, n11682_0/**/, n11677_0, n11661_0, n11644_0, n11630_0, n11625_0, n11606_1, n7126, n7114, n6146, n6138}), .out(n14060), .config_in(config_chain[33507:33502]), .config_rst(config_rst)); 
buffer_wire buffer_14060 (.in(n14060), .out(n14060_0));
mux3 mux_8895 (.in({n12183_0, n12182_0, n7212}), .out(n14061), .config_in(config_chain[33509:33508]), .config_rst(config_rst)); 
buffer_wire buffer_14061 (.in(n14061), .out(n14061_0));
mux13 mux_8896 (.in({n13974_1/**/, n11705_0, n11668_0, n11652_0, n11647_0, n11638_0, n11633_0, n11604_1, n11597_0, n7126, n7118, n6146, n6138}), .out(n14062), .config_in(config_chain[33515:33510]), .config_rst(config_rst)); 
buffer_wire buffer_14062 (.in(n14062), .out(n14062_0));
mux3 mux_8897 (.in({n12185_0, n12184_0/**/, n7216}), .out(n14063), .config_in(config_chain[33517:33516]), .config_rst(config_rst)); 
buffer_wire buffer_14063 (.in(n14063), .out(n14063_0));
mux13 mux_8898 (.in({n13976_1, n11707_0, n11676_0, n11671_0/**/, n11660_0, n11655_0, n11624_0, n11619_0, n11602_1, n7126, n7118, n6150, n6138}), .out(n14064), .config_in(config_chain[33523:33518]), .config_rst(config_rst)); 
buffer_wire buffer_14064 (.in(n14064), .out(n14064_0));
mux3 mux_8899 (.in({n12187_0, n12186_0, n7220/**/}), .out(n14065), .config_in(config_chain[33525:33524]), .config_rst(config_rst)); 
buffer_wire buffer_14065 (.in(n14065), .out(n14065_0));
mux13 mux_8900 (.in({n13914_2, n11687_0, n11679_0/**/, n11646_0, n11641_0, n11632_0, n11627_0, n11600_1, n11596_1, n7126, n7118, n6150, n6142}), .out(n14066), .config_in(config_chain[33531:33526]), .config_rst(config_rst)); 
buffer_wire buffer_14066 (.in(n14066), .out(n14066_0));
mux3 mux_8901 (.in({n12189_0, n12188_0, n7228}), .out(n14067), .config_in(config_chain[33533:33532]), .config_rst(config_rst)); 
buffer_wire buffer_14067 (.in(n14067), .out(n14067_0));
mux16 mux_8902 (.in({n13980_1, n11953_0, n11935_0, n11930_0, n11926_0, n11922_0, n11907_0, n11897_0, n11892_0, n11862_1, n11829_0, n7224, n7216, n6248, n6240, n6232}), .out(n14068), .config_in(config_chain[33539:33534]), .config_rst(config_rst)); 
buffer_wire buffer_14068 (.in(n14068), .out(n14068_0));
mux4 mux_8903 (.in({n12191_0, n12190_0, n7228, n6232}), .out(n14069), .config_in(config_chain[33541:33540]), .config_rst(config_rst)); 
buffer_wire buffer_14069 (.in(n14069), .out(n14069_0));
mux16 mux_8904 (.in({n13982_1, n11955_0, n11948_0/**/, n11944_0, n11929_0, n11921_0, n11916_0, n11891_0, n11886_0, n11880_1, n11861_0, n7224, n7216, n6248, n6240, n6232}), .out(n14070), .config_in(config_chain[33547:33542]), .config_rst(config_rst)); 
buffer_wire buffer_14070 (.in(n14070), .out(n14070_0));
mux3 mux_8905 (.in({n12193_0, n12192_0, n6236}), .out(n14071), .config_in(config_chain[33549:33548]), .config_rst(config_rst)); 
buffer_wire buffer_14071 (.in(n14071), .out(n14071_0));
mux15 mux_8906 (.in({n13984_1, n11957_0, n11943_0, n11938_0, n11915_0, n11910_0, n11900_0, n11885_0, n11883_0, n11878_1, n7224, n7216, n6248, n6240, n6232}), .out(n14072), .config_in(config_chain[33555:33550]), .config_rst(config_rst)); 
buffer_wire buffer_14072 (.in(n14072), .out(n14072_0));
mux3 mux_8907 (.in({n12195_0, n12194_0, n6240}), .out(n14073), .config_in(config_chain[33557:33556]), .config_rst(config_rst)); 
buffer_wire buffer_14073 (.in(n14073), .out(n14073_0));
mux15 mux_8908 (.in({n13986_1, n11959_0, n11937_0, n11932_0, n11924_0, n11909_0, n11905_0, n11899_0, n11894_0, n11876_1, n7224, n7216, n6248, n6240, n6232}), .out(n14074), .config_in(config_chain[33563:33558]), .config_rst(config_rst)); 
buffer_wire buffer_14074 (.in(n14074), .out(n14074_0));
mux3 mux_8909 (.in({n12197_0, n12196_0, n6240}), .out(n14075), .config_in(config_chain[33565:33564]), .config_rst(config_rst)); 
buffer_wire buffer_14075 (.in(n14075), .out(n14075_0));
mux15 mux_8910 (.in({n13988_1, n11961_0, n11946_0, n11931_0, n11927_0, n11923_0, n11918_0, n11893_0, n11888_0, n11874_1, n7224, n7216, n6248, n6240, n6232}), .out(n14076), .config_in(config_chain[33571:33566]), .config_rst(config_rst)); 
buffer_wire buffer_14076 (.in(n14076), .out(n14076_0));
mux3 mux_8911 (.in({n12199_0, n12198_0, n6244}), .out(n14077), .config_in(config_chain[33573:33572]), .config_rst(config_rst)); 
buffer_wire buffer_14077 (.in(n14077), .out(n14077_0));
mux15 mux_8912 (.in({n13990_1, n11963_0, n11949_0, n11945_0, n11940_0, n11917_0, n11912_0, n11902_0/**/, n11887_0, n11872_1, n7228, n7220, n7212, n6244, n6236}), .out(n14078), .config_in(config_chain[33579:33574]), .config_rst(config_rst)); 
buffer_wire buffer_14078 (.in(n14078), .out(n14078_0));
mux3 mux_8913 (.in({n12201_0, n12200_0, n6248}), .out(n14079), .config_in(config_chain[33581:33580]), .config_rst(config_rst)); 
buffer_wire buffer_14079 (.in(n14079), .out(n14079_0));
mux15 mux_8914 (.in({n13992_1, n11965_0, n11939_0, n11934_0, n11911_0, n11906_0, n11901_0/**/, n11896_0, n11870_1, n11828_1, n7228, n7220, n7212, n6244, n6236}), .out(n14080), .config_in(config_chain[33587:33582]), .config_rst(config_rst)); 
buffer_wire buffer_14080 (.in(n14080), .out(n14080_0));
mux3 mux_8915 (.in({n12203_0/**/, n12202_0, n7212}), .out(n14081), .config_in(config_chain[33589:33588]), .config_rst(config_rst)); 
buffer_wire buffer_14081 (.in(n14081), .out(n14081_0));
mux15 mux_8916 (.in({n13994_1, n11967_0, n11933_0, n11928_0, n11925_0, n11920_0, n11895_0, n11890_0, n11868_1, n11860_1, n7228, n7220, n7212, n6244, n6236}), .out(n14082), .config_in(config_chain[33595:33590]), .config_rst(config_rst)); 
buffer_wire buffer_14082 (.in(n14082), .out(n14082_0));
mux3 mux_8917 (.in({n12205_0/**/, n12204_0, n7216}), .out(n14083), .config_in(config_chain[33597:33596]), .config_rst(config_rst)); 
buffer_wire buffer_14083 (.in(n14083), .out(n14083_0));
mux15 mux_8918 (.in({n13996_1, n11969_0, n11947_0, n11942_0, n11919_0, n11914_0, n11889_0, n11884_0, n11882_1, n11866_1, n7228, n7220, n7212, n6244, n6236}), .out(n14084), .config_in(config_chain[33603:33598]), .config_rst(config_rst)); 
buffer_wire buffer_14084 (.in(n14084), .out(n14084_0));
mux3 mux_8919 (.in({n12207_0, n12206_0, n7216}), .out(n14085), .config_in(config_chain[33605:33604]), .config_rst(config_rst)); 
buffer_wire buffer_14085 (.in(n14085), .out(n14085_0));
mux15 mux_8920 (.in({n13998_1, n11951_0, n11941_0, n11936_0, n11913_0, n11908_0, n11904_0, n11903_0, n11898_0, n11864_1, n7228, n7220, n7212, n6244, n6236}), .out(n14086), .config_in(config_chain[33611:33606]), .config_rst(config_rst)); 
buffer_wire buffer_14086 (.in(n14086), .out(n14086_0));
mux3 mux_8921 (.in({n12209_0, n12208_0/**/, n7220}), .out(n14087), .config_in(config_chain[33613:33612]), .config_rst(config_rst)); 
buffer_wire buffer_14087 (.in(n14087), .out(n14087_0));
mux4 mux_8922 (.in({n9819_0, n9818_0, n7422, n6426}), .out(n14088), .config_in(config_chain[33615:33614]), .config_rst(config_rst)); 
buffer_wire buffer_14088 (.in(n14088), .out(n14088_0));
mux15 mux_8923 (.in({n14181_1, n10151_0, n10125_0, n10118_0/**/, n10106_0, n10079_0, n10072_0, n10054_1, n10008_2, n10005_0, n7418, n7410, n6442, n6434, n6426}), .out(n14089), .config_in(config_chain[33621:33616]), .config_rst(config_rst)); 
buffer_wire buffer_14089 (.in(n14089), .out(n14089_0));
mux4 mux_8924 (.in({n9839_0, n9838_0, n7422, n6426}), .out(n14090), .config_in(config_chain[33623:33622]), .config_rst(config_rst)); 
buffer_wire buffer_14090 (.in(n14090), .out(n14090_0));
mux15 mux_8925 (.in({n14203_1, n10409_0, n10375_0, n10368_0, n10361_0, n10354_0, n10342_0, n10310_1, n10264_2, n10261_0, n7516, n7508, n6540, n6532, n6524}), .out(n14091), .config_in(config_chain[33629:33624]), .config_rst(config_rst)); 
buffer_wire buffer_14091 (.in(n14091), .out(n14091_0));
mux4 mux_8926 (.in({n9859_0, n9858_0/**/, n7422, n6426}), .out(n14092), .config_in(config_chain[33631:33630]), .config_rst(config_rst)); 
buffer_wire buffer_14092 (.in(n14092), .out(n14092_0));
mux15 mux_8927 (.in({n14225_1, n10669_0, n10649_0, n10642_0, n10613_0, n10606_0, n10599_0, n10592_0, n10568_1, n10522_2, n7614, n7606, n6638, n6630, n6622}), .out(n14093), .config_in(config_chain[33637:33632]), .config_rst(config_rst)); 
buffer_wire buffer_14093 (.in(n14093), .out(n14093_0));
mux4 mux_8928 (.in({n9879_0, n9798_1, n7422, n6426}), .out(n14094), .config_in(config_chain[33639:33638]), .config_rst(config_rst)); 
buffer_wire buffer_14094 (.in(n14094), .out(n14094_0));
mux15 mux_8929 (.in({n14247_1, n10931_0, n10903_0, n10896_0, n10889_0, n10882_0, n10853_0, n10846_0/**/, n10828_1, n10782_2, n7712, n7704, n6736, n6728, n6720}), .out(n14095), .config_in(config_chain[33645:33640]), .config_rst(config_rst)); 
buffer_wire buffer_14095 (.in(n14095), .out(n14095_0));
mux3 mux_8930 (.in({n9821_0, n9820_0/**/, n6426}), .out(n14096), .config_in(config_chain[33647:33646]), .config_rst(config_rst)); 
buffer_wire buffer_14096 (.in(n14096), .out(n14096_0));
mux15 mux_8931 (.in({n14183_1, n10149_0, n10126_0, n10099_0, n10092_0/**/, n10087_0, n10080_0, n10056_1, n10010_2, n10007_0, n7422, n7410, n6442, n6434, n6426}), .out(n14097), .config_in(config_chain[33653:33648]), .config_rst(config_rst)); 
buffer_wire buffer_14097 (.in(n14097), .out(n14097_0));
mux3 mux_8932 (.in({n9841_0, n9840_0, n6430}), .out(n14098), .config_in(config_chain[33655:33654]), .config_rst(config_rst)); 
buffer_wire buffer_14098 (.in(n14098), .out(n14098_0));
mux15 mux_8933 (.in({n14205_1, n10407_0, n10383_0, n10376_0, n10362_0, n10335_0, n10328_0, n10312_1, n10266_2, n10263_0, n7520, n7508, n6540, n6532, n6524/**/}), .out(n14099), .config_in(config_chain[33661:33656]), .config_rst(config_rst)); 
buffer_wire buffer_14099 (.in(n14099), .out(n14099_0));
mux3 mux_8934 (.in({n9861_0, n9860_0/**/, n6430}), .out(n14100), .config_in(config_chain[33663:33662]), .config_rst(config_rst)); 
buffer_wire buffer_14100 (.in(n14100), .out(n14100_0));
mux15 mux_8935 (.in({n14227_1, n10667_0, n10635_0/**/, n10628_0, n10621_0, n10614_0, n10600_0, n10570_1, n10524_2, n10521_0, n7618, n7606, n6638, n6630, n6622}), .out(n14101), .config_in(config_chain[33669:33664]), .config_rst(config_rst)); 
buffer_wire buffer_14101 (.in(n14101), .out(n14101_0));
mux3 mux_8936 (.in({n9881_0, n9800_1/**/, n6430}), .out(n14102), .config_in(config_chain[33671:33670]), .config_rst(config_rst)); 
buffer_wire buffer_14102 (.in(n14102), .out(n14102_0));
mux15 mux_8937 (.in({n14249_1, n10929_0, n10911_0, n10904_0, n10875_0, n10868_0, n10861_0, n10854_0, n10830_1/**/, n10784_2, n7716, n7704, n6736, n6728, n6720}), .out(n14103), .config_in(config_chain[33677:33672]), .config_rst(config_rst)); 
buffer_wire buffer_14103 (.in(n14103), .out(n14103_0));
mux3 mux_8938 (.in({n9823_0, n9822_0, n6430}), .out(n14104), .config_in(config_chain[33679:33678]), .config_rst(config_rst)); 
buffer_wire buffer_14104 (.in(n14104), .out(n14104_0));
mux15 mux_8939 (.in({n14185_1, n10147_0/**/, n10119_0, n10112_0, n10107_0, n10100_0, n10088_0, n10073_0, n10058_1, n10009_0, n7422, n7414, n6442, n6434, n6426}), .out(n14105), .config_in(config_chain[33685:33680]), .config_rst(config_rst)); 
buffer_wire buffer_14105 (.in(n14105), .out(n14105_0));
mux3 mux_8940 (.in({n9843_0, n9842_0, n6430}), .out(n14106), .config_in(config_chain[33687:33686]), .config_rst(config_rst)); 
buffer_wire buffer_14106 (.in(n14106), .out(n14106_0));
mux15 mux_8941 (.in({n14207_1, n10405_0, n10384_0, n10369_0, n10355_0, n10348_0, n10343_0, n10336_0, n10314_1, n10265_0, n7520, n7512, n6540/**/, n6532, n6524}), .out(n14107), .config_in(config_chain[33693:33688]), .config_rst(config_rst)); 
buffer_wire buffer_14107 (.in(n14107), .out(n14107_0));
mux3 mux_8942 (.in({n9863_0, n9862_0, n6434}), .out(n14108), .config_in(config_chain[33695:33694]), .config_rst(config_rst)); 
buffer_wire buffer_14108 (.in(n14108), .out(n14108_0));
mux15 mux_8943 (.in({n14229_1, n10665_0, n10643_0, n10636_0, n10622_0, n10607_0, n10593_0, n10586_0, n10572_1/**/, n10523_0, n7618, n7610, n6638, n6630, n6622}), .out(n14109), .config_in(config_chain[33701:33696]), .config_rst(config_rst)); 
buffer_wire buffer_14109 (.in(n14109), .out(n14109_0));
mux3 mux_8944 (.in({n9883_0, n9802_1, n6434}), .out(n14110), .config_in(config_chain[33703:33702]), .config_rst(config_rst)); 
buffer_wire buffer_14110 (.in(n14110), .out(n14110_0));
mux15 mux_8945 (.in({n14251_1, n10927_0, n10897_0, n10890_0, n10883_0, n10876_0, n10862_0, n10847_0, n10832_1, n10783_0, n7716, n7708, n6736, n6728, n6720}), .out(n14111), .config_in(config_chain[33709:33704]), .config_rst(config_rst)); 
buffer_wire buffer_14111 (.in(n14111), .out(n14111_0));
mux3 mux_8946 (.in({n9825_0, n9824_0/**/, n6434}), .out(n14112), .config_in(config_chain[33711:33710]), .config_rst(config_rst)); 
buffer_wire buffer_14112 (.in(n14112), .out(n14112_0));
mux15 mux_8947 (.in({n14187_1, n10145_0, n10127_0, n10120_0/**/, n10108_0, n10093_0, n10081_0, n10074_0, n10060_1, n10011_0, n7422, n7414, n7406, n6434, n6426}), .out(n14113), .config_in(config_chain[33717:33712]), .config_rst(config_rst)); 
buffer_wire buffer_14113 (.in(n14113), .out(n14113_0));
mux3 mux_8948 (.in({n9845_0, n9844_0, n6434}), .out(n14114), .config_in(config_chain[33719:33718]), .config_rst(config_rst)); 
buffer_wire buffer_14114 (.in(n14114), .out(n14114_0));
mux15 mux_8949 (.in({n14209_1, n10403_0, n10377_0, n10370_0, n10363_0, n10356_0, n10344_0, n10329_0, n10316_1/**/, n10267_0, n7520, n7512, n7504, n6532, n6524}), .out(n14115), .config_in(config_chain[33725:33720]), .config_rst(config_rst)); 
buffer_wire buffer_14115 (.in(n14115), .out(n14115_0));
mux3 mux_8950 (.in({n9865_0, n9864_0, n6434}), .out(n14116), .config_in(config_chain[33727:33726]), .config_rst(config_rst)); 
buffer_wire buffer_14116 (.in(n14116), .out(n14116_0));
mux15 mux_8951 (.in({n14231_1, n10663_0, n10644_0, n10629_0, n10615_0, n10608_0, n10601_0, n10594_0, n10574_1, n10525_0, n7618, n7610, n7602/**/, n6630, n6622}), .out(n14117), .config_in(config_chain[33733:33728]), .config_rst(config_rst)); 
buffer_wire buffer_14117 (.in(n14117), .out(n14117_0));
mux3 mux_8952 (.in({n9885_0, n9804_1/**/, n6438}), .out(n14118), .config_in(config_chain[33735:33734]), .config_rst(config_rst)); 
buffer_wire buffer_14118 (.in(n14118), .out(n14118_0));
mux15 mux_8953 (.in({n14253_1, n10925_0, n10905_0, n10898_0, n10884_0, n10869_0, n10855_0/**/, n10848_0, n10834_1, n10785_0, n7716, n7708, n7700, n6728, n6720}), .out(n14119), .config_in(config_chain[33741:33736]), .config_rst(config_rst)); 
buffer_wire buffer_14119 (.in(n14119), .out(n14119_0));
mux3 mux_8954 (.in({n9827_0, n9826_0/**/, n6438}), .out(n14120), .config_in(config_chain[33743:33742]), .config_rst(config_rst)); 
buffer_wire buffer_14120 (.in(n14120), .out(n14120_0));
mux14 mux_8955 (.in({n14189_1, n10143_0, n10128_0, n10113_0, n10101_0, n10094_0, n10089_0, n10082_0, n10062_1, n7422, n7414, n7406, n6438, n6426}), .out(n14121), .config_in(config_chain[33749:33744]), .config_rst(config_rst)); 
buffer_wire buffer_14121 (.in(n14121), .out(n14121_0));
mux3 mux_8956 (.in({n9847_0, n9846_0, n6438}), .out(n14122), .config_in(config_chain[33751:33750]), .config_rst(config_rst)); 
buffer_wire buffer_14122 (.in(n14122), .out(n14122_0));
mux14 mux_8957 (.in({n14211_1/**/, n10401_0, n10385_0, n10378_0, n10364_0, n10349_0, n10337_0, n10330_0, n10318_1, n7520, n7512, n7504, n6536, n6524}), .out(n14123), .config_in(config_chain[33757:33752]), .config_rst(config_rst)); 
buffer_wire buffer_14123 (.in(n14123), .out(n14123_0));
mux3 mux_8958 (.in({n9867_0, n9866_0/**/, n6438}), .out(n14124), .config_in(config_chain[33759:33758]), .config_rst(config_rst)); 
buffer_wire buffer_14124 (.in(n14124), .out(n14124_0));
mux14 mux_8959 (.in({n14233_1, n10661_0, n10637_0, n10630_0, n10623_0, n10616_0, n10602_0, n10587_0, n10576_1, n7618, n7610, n7602, n6634, n6622}), .out(n14125), .config_in(config_chain[33765:33760]), .config_rst(config_rst)); 
buffer_wire buffer_14125 (.in(n14125), .out(n14125_0));
mux3 mux_8960 (.in({n9887_0, n9806_1, n6438}), .out(n14126), .config_in(config_chain[33767:33766]), .config_rst(config_rst)); 
buffer_wire buffer_14126 (.in(n14126), .out(n14126_0));
mux14 mux_8961 (.in({n14255_1, n10923_0, n10906_0, n10891_0, n10877_0, n10870_0/**/, n10863_0, n10856_0, n10836_1, n7716, n7708, n7700, n6732, n6720}), .out(n14127), .config_in(config_chain[33773:33768]), .config_rst(config_rst)); 
buffer_wire buffer_14127 (.in(n14127), .out(n14127_0));
mux3 mux_8962 (.in({n9829_0, n9828_0/**/, n6442}), .out(n14128), .config_in(config_chain[33775:33774]), .config_rst(config_rst)); 
buffer_wire buffer_14128 (.in(n14128), .out(n14128_0));
mux14 mux_8963 (.in({n14191_1, n10141_0, n10121_0, n10114_0, n10109_0, n10102_0, n10090_0, n10075_0, n10064_1, n7422, n7414, n7406, n6438, n6430/**/}), .out(n14129), .config_in(config_chain[33781:33776]), .config_rst(config_rst)); 
buffer_wire buffer_14129 (.in(n14129), .out(n14129_0));
mux3 mux_8964 (.in({n9849_0, n9848_0/**/, n6442}), .out(n14130), .config_in(config_chain[33783:33782]), .config_rst(config_rst)); 
buffer_wire buffer_14130 (.in(n14130), .out(n14130_0));
mux14 mux_8965 (.in({n14213_1, n10399_0, n10386_0, n10371_0, n10357_0, n10350_0, n10345_0, n10338_0, n10320_1, n7520, n7512, n7504, n6536/**/, n6528}), .out(n14131), .config_in(config_chain[33789:33784]), .config_rst(config_rst)); 
buffer_wire buffer_14131 (.in(n14131), .out(n14131_0));
mux3 mux_8966 (.in({n9869_0, n9868_0/**/, n6442}), .out(n14132), .config_in(config_chain[33791:33790]), .config_rst(config_rst)); 
buffer_wire buffer_14132 (.in(n14132), .out(n14132_0));
mux14 mux_8967 (.in({n14235_1, n10659_0, n10645_0, n10638_0, n10624_0, n10609_0, n10595_0, n10588_0, n10578_1, n7618/**/, n7610, n7602, n6634, n6626}), .out(n14133), .config_in(config_chain[33797:33792]), .config_rst(config_rst)); 
buffer_wire buffer_14133 (.in(n14133), .out(n14133_0));
mux3 mux_8968 (.in({n9889_0, n9808_1/**/, n6442}), .out(n14134), .config_in(config_chain[33799:33798]), .config_rst(config_rst)); 
buffer_wire buffer_14134 (.in(n14134), .out(n14134_0));
mux14 mux_8969 (.in({n14257_1, n10921_0, n10899_0, n10892_0, n10885_0, n10878_0, n10864_0, n10849_0, n10838_1, n7716, n7708/**/, n7700, n6732, n6724}), .out(n14135), .config_in(config_chain[33805:33800]), .config_rst(config_rst)); 
buffer_wire buffer_14135 (.in(n14135), .out(n14135_0));
mux3 mux_8970 (.in({n9831_0, n9830_0/**/, n6442}), .out(n14136), .config_in(config_chain[33807:33806]), .config_rst(config_rst)); 
buffer_wire buffer_14136 (.in(n14136), .out(n14136_0));
mux13 mux_8971 (.in({n14193_1, n10139_0/**/, n10129_0, n10122_0, n10110_0, n10095_0, n10083_0, n10076_0, n10066_1, n7414, n7406, n6438, n6430}), .out(n14137), .config_in(config_chain[33813:33808]), .config_rst(config_rst)); 
buffer_wire buffer_14137 (.in(n14137), .out(n14137_0));
mux3 mux_8972 (.in({n9851_0, n9850_0, n7406}), .out(n14138), .config_in(config_chain[33815:33814]), .config_rst(config_rst)); 
buffer_wire buffer_14138 (.in(n14138), .out(n14138_0));
mux13 mux_8973 (.in({n14215_1, n10397_0, n10379_0, n10372_0, n10365_0, n10358_0, n10346_0, n10331_0, n10322_1, n7512, n7504, n6536, n6528}), .out(n14139), .config_in(config_chain[33821:33816]), .config_rst(config_rst)); 
buffer_wire buffer_14139 (.in(n14139), .out(n14139_0));
mux3 mux_8974 (.in({n9871_0, n9870_0/**/, n7406}), .out(n14140), .config_in(config_chain[33823:33822]), .config_rst(config_rst)); 
buffer_wire buffer_14140 (.in(n14140), .out(n14140_0));
mux13 mux_8975 (.in({n14237_1, n10657_0/**/, n10646_0, n10631_0, n10617_0, n10610_0, n10603_0, n10596_0, n10580_1, n7610, n7602, n6634, n6626}), .out(n14141), .config_in(config_chain[33829:33824]), .config_rst(config_rst)); 
buffer_wire buffer_14141 (.in(n14141), .out(n14141_0));
mux3 mux_8976 (.in({n9891_0, n9810_1/**/, n7406}), .out(n14142), .config_in(config_chain[33831:33830]), .config_rst(config_rst)); 
buffer_wire buffer_14142 (.in(n14142), .out(n14142_0));
mux13 mux_8977 (.in({n14259_1, n10919_0, n10907_0, n10900_0, n10886_0, n10871_0, n10857_0, n10850_0/**/, n10840_1, n7708, n7700, n6732, n6724}), .out(n14143), .config_in(config_chain[33837:33832]), .config_rst(config_rst)); 
buffer_wire buffer_14143 (.in(n14143), .out(n14143_0));
mux3 mux_8978 (.in({n9833_0, n9832_0/**/, n7406}), .out(n14144), .config_in(config_chain[33839:33838]), .config_rst(config_rst)); 
buffer_wire buffer_14144 (.in(n14144), .out(n14144_0));
mux13 mux_8979 (.in({n14195_1, n10137_0, n10130_0, n10115_0, n10103_0, n10096_0, n10091_0, n10084_0, n10068_1, n7418, n7406, n6438, n6430}), .out(n14145), .config_in(config_chain[33845:33840]), .config_rst(config_rst)); 
buffer_wire buffer_14145 (.in(n14145), .out(n14145_0));
mux3 mux_8980 (.in({n9853_0, n9852_0, n7406}), .out(n14146), .config_in(config_chain[33847:33846]), .config_rst(config_rst)); 
buffer_wire buffer_14146 (.in(n14146), .out(n14146_0));
mux13 mux_8981 (.in({n14217_1, n10395_0, n10387_0, n10380_0, n10366_0, n10351_0, n10339_0, n10332_0, n10324_1/**/, n7516, n7504, n6536, n6528}), .out(n14147), .config_in(config_chain[33853:33848]), .config_rst(config_rst)); 
buffer_wire buffer_14147 (.in(n14147), .out(n14147_0));
mux3 mux_8982 (.in({n9873_0, n9872_0, n7410}), .out(n14148), .config_in(config_chain[33855:33854]), .config_rst(config_rst)); 
buffer_wire buffer_14148 (.in(n14148), .out(n14148_0));
mux13 mux_8983 (.in({n14239_1, n10655_0, n10639_0, n10632_0, n10625_0, n10618_0, n10604_0, n10589_0, n10582_1/**/, n7614, n7602, n6634, n6626}), .out(n14149), .config_in(config_chain[33861:33856]), .config_rst(config_rst)); 
buffer_wire buffer_14149 (.in(n14149), .out(n14149_0));
mux3 mux_8984 (.in({n9893_0/**/, n9812_1, n7410}), .out(n14150), .config_in(config_chain[33863:33862]), .config_rst(config_rst)); 
buffer_wire buffer_14150 (.in(n14150), .out(n14150_0));
mux13 mux_8985 (.in({n14261_1, n10917_0, n10908_0, n10893_0, n10879_0, n10872_0, n10865_0, n10858_0, n10842_1, n7712, n7700, n6732, n6724/**/}), .out(n14151), .config_in(config_chain[33869:33864]), .config_rst(config_rst)); 
buffer_wire buffer_14151 (.in(n14151), .out(n14151_0));
mux3 mux_8986 (.in({n9835_0, n9834_0, n7410}), .out(n14152), .config_in(config_chain[33871:33870]), .config_rst(config_rst)); 
buffer_wire buffer_14152 (.in(n14152), .out(n14152_0));
mux13 mux_8987 (.in({n14197_1, n10135_0, n10123_0, n10116_0, n10111_0, n10104_0, n10077_0, n10070_1, n10002_2, n7418, n7410, n6438, n6430}), .out(n14153), .config_in(config_chain[33877:33872]), .config_rst(config_rst)); 
buffer_wire buffer_14153 (.in(n14153), .out(n14153_0));
mux3 mux_8988 (.in({n9855_0, n9854_0, n7410}), .out(n14154), .config_in(config_chain[33879:33878]), .config_rst(config_rst)); 
buffer_wire buffer_14154 (.in(n14154), .out(n14154_0));
mux13 mux_8989 (.in({n14219_1, n10393_0, n10388_0, n10373_0, n10359_0, n10352_0, n10347_0, n10340_0, n10326_1, n7516, n7508, n6536, n6528}), .out(n14155), .config_in(config_chain[33885:33880]), .config_rst(config_rst)); 
buffer_wire buffer_14155 (.in(n14155), .out(n14155_0));
mux3 mux_8990 (.in({n9875_0, n9874_0, n7410}), .out(n14156), .config_in(config_chain[33887:33886]), .config_rst(config_rst)); 
buffer_wire buffer_14156 (.in(n14156), .out(n14156_0));
mux13 mux_8991 (.in({n14241_1, n10653_0, n10647_0, n10640_0, n10626_0, n10611_0, n10597_0, n10590_0, n10584_1, n7614, n7606, n6634, n6626}), .out(n14157), .config_in(config_chain[33893:33888]), .config_rst(config_rst)); 
buffer_wire buffer_14157 (.in(n14157), .out(n14157_0));
mux3 mux_8992 (.in({n9895_0, n9814_1/**/, n7414}), .out(n14158), .config_in(config_chain[33895:33894]), .config_rst(config_rst)); 
buffer_wire buffer_14158 (.in(n14158), .out(n14158_0));
mux13 mux_8993 (.in({n14263_1, n10915_0, n10901_0, n10894_0, n10887_0, n10880_0, n10866_0, n10851_0, n10844_1, n7712/**/, n7704, n6732, n6724}), .out(n14159), .config_in(config_chain[33901:33896]), .config_rst(config_rst)); 
buffer_wire buffer_14159 (.in(n14159), .out(n14159_0));
mux3 mux_8994 (.in({n9837_0, n9836_0, n7414}), .out(n14160), .config_in(config_chain[33903:33902]), .config_rst(config_rst)); 
buffer_wire buffer_14160 (.in(n14160), .out(n14160_0));
mux13 mux_8995 (.in({n14199_1, n10133_0, n10131_0, n10124_0, n10097_0, n10085_0, n10078_0/**/, n10004_2, n10000_2, n7418, n7410, n6442, n6430}), .out(n14161), .config_in(config_chain[33909:33904]), .config_rst(config_rst)); 
buffer_wire buffer_14161 (.in(n14161), .out(n14161_0));
mux3 mux_8996 (.in({n9857_0, n9856_0, n7414}), .out(n14162), .config_in(config_chain[33911:33910]), .config_rst(config_rst)); 
buffer_wire buffer_14162 (.in(n14162), .out(n14162_0));
mux13 mux_8997 (.in({n14221_1, n10391_0, n10381_0, n10374_0, n10367_0, n10360_0, n10333_0, n10260_2, n10258_2, n7516, n7508, n6540, n6528}), .out(n14163), .config_in(config_chain[33917:33912]), .config_rst(config_rst)); 
buffer_wire buffer_14163 (.in(n14163), .out(n14163_0));
mux3 mux_8998 (.in({n9877_0, n9876_0, n7414}), .out(n14164), .config_in(config_chain[33919:33918]), .config_rst(config_rst)); 
buffer_wire buffer_14164 (.in(n14164), .out(n14164_0));
mux13 mux_8999 (.in({n14243_1, n10651_0, n10648_0, n10633_0, n10619_0, n10612_0, n10605_0, n10598_0, n10518_2, n7614, n7606, n6638, n6626}), .out(n14165), .config_in(config_chain[33925:33920]), .config_rst(config_rst)); 
buffer_wire buffer_14165 (.in(n14165), .out(n14165_0));
mux3 mux_9000 (.in({n9897_0/**/, n9816_1, n7414}), .out(n14166), .config_in(config_chain[33927:33926]), .config_rst(config_rst)); 
buffer_wire buffer_14166 (.in(n14166), .out(n14166_0));
mux13 mux_9001 (.in({n14265_1, n10913_0, n10909_0, n10902_0, n10888_0, n10873_0, n10859_0, n10852_0, n10780_2, n7712, n7704, n6736, n6724}), .out(n14167), .config_in(config_chain[33933:33928]), .config_rst(config_rst)); 
buffer_wire buffer_14167 (.in(n14167), .out(n14167_0));
mux3 mux_9002 (.in({n9747_0, n9746_2, n7418}), .out(n14168), .config_in(config_chain[33935:33934]), .config_rst(config_rst)); 
buffer_wire buffer_14168 (.in(n14168), .out(n14168_0));
mux13 mux_9003 (.in({n14201_2, n10153_0, n10117_0, n10105_0, n10098_0, n10086_0, n10052_1, n10006_2, n10003_0/**/, n7418, n7410, n6442, n6434}), .out(n14169), .config_in(config_chain[33941:33936]), .config_rst(config_rst)); 
buffer_wire buffer_14169 (.in(n14169), .out(n14169_0));
mux3 mux_9004 (.in({n9749_0, n9748_2, n7418}), .out(n14170), .config_in(config_chain[33943:33942]), .config_rst(config_rst)); 
buffer_wire buffer_14170 (.in(n14170), .out(n14170_0));
mux13 mux_9005 (.in({n14223_2, n10411_0, n10389_0, n10382_0, n10353_0, n10341_0, n10334_0, n10308_1, n10262_2, n7516, n7508, n6540, n6532}), .out(n14171), .config_in(config_chain[33949:33944]), .config_rst(config_rst)); 
buffer_wire buffer_14171 (.in(n14171), .out(n14171_0));
mux3 mux_9006 (.in({n9751_0, n9750_2, n7418}), .out(n14172), .config_in(config_chain[33951:33950]), .config_rst(config_rst)); 
buffer_wire buffer_14172 (.in(n14172), .out(n14172_0));
mux13 mux_9007 (.in({n14245_1, n10671_0, n10641_0, n10634_0, n10627_0, n10620_0, n10591_0, n10566_1/**/, n10520_2, n7614, n7606, n6638, n6630}), .out(n14173), .config_in(config_chain[33957:33952]), .config_rst(config_rst)); 
buffer_wire buffer_14173 (.in(n14173), .out(n14173_0));
mux3 mux_9008 (.in({n9753_0/**/, n9752_2, n7418}), .out(n14174), .config_in(config_chain[33959:33958]), .config_rst(config_rst)); 
buffer_wire buffer_14174 (.in(n14174), .out(n14174_0));
mux13 mux_9009 (.in({n14267_1/**/, n10933_0, n10910_0, n10895_0, n10881_0, n10874_0, n10867_0, n10860_0, n10826_1, n7712, n7704, n6736, n6728}), .out(n14175), .config_in(config_chain[33965:33960]), .config_rst(config_rst)); 
buffer_wire buffer_14175 (.in(n14175), .out(n14175_0));
mux3 mux_9010 (.in({n9755_0, n9754_2, n7418}), .out(n14176), .config_in(config_chain[33967:33966]), .config_rst(config_rst)); 
buffer_wire buffer_14176 (.in(n14176), .out(n14176_0));
mux13 mux_9011 (.in({n14289_1, n11197_0, n11159_0, n11152_0, n11145_0, n11138_0, n11124_0, n11109_0, n11088_1/**/, n7810, n7802, n6834, n6826}), .out(n14177), .config_in(config_chain[33973:33968]), .config_rst(config_rst)); 
buffer_wire buffer_14177 (.in(n14177), .out(n14177_0));
mux3 mux_9012 (.in({n9757_0, n9756_2, n7422}), .out(n14178), .config_in(config_chain[33975:33974]), .config_rst(config_rst)); 
buffer_wire buffer_14178 (.in(n14178), .out(n14178_0));
mux13 mux_9013 (.in({n14311_0, n11463_0, n11434_0, n11403_0, n11396_0, n11389_0, n11382_0, n11354_1, n11353_0, n7908, n7900, n6932, n6924}), .out(n14179), .config_in(config_chain[33981:33976]), .config_rst(config_rst)); 
buffer_wire buffer_14179 (.in(n14179), .out(n14179_0));
mux15 mux_9014 (.in({n14088_0, n10135_0, n10124_0/**/, n10119_0, n10107_0, n10078_0, n10073_0, n10052_1, n10009_0, n10004_2, n7516, n7508, n6540, n6532, n6524}), .out(n14180), .config_in(config_chain[33987:33982]), .config_rst(config_rst)); 
buffer_wire buffer_14180 (.in(n14180), .out(n14180_0));
mux15 mux_9015 (.in({n14269_1/**/, n11195_0, n11174_0, n11167_0, n11160_0, n11146_0, n11131_0, n11117_0, n11110_0, n11090_1, n7810, n7802, n6834, n6826, n6818}), .out(n14181), .config_in(config_chain[33993:33988]), .config_rst(config_rst)); 
buffer_wire buffer_14181 (.in(n14181), .out(n14181_0));
mux15 mux_9016 (.in({n14096_0, n10137_0, n10127_0, n10098_0, n10093_0, n10086_0, n10081_0, n10011_0, n10006_2, n10000_2, n7520/**/, n7508, n6540, n6532, n6524}), .out(n14182), .config_in(config_chain[33999:33994]), .config_rst(config_rst)); 
buffer_wire buffer_14182 (.in(n14182), .out(n14182_0));
mux15 mux_9017 (.in({n14271_1, n11193_0, n11168_0, n11153_0, n11139_0, n11132_0, n11125_0, n11118_0, n11092_1, n11046_2, n7814/**/, n7802, n6834, n6826, n6818}), .out(n14183), .config_in(config_chain[34005:34000]), .config_rst(config_rst)); 
buffer_wire buffer_14183 (.in(n14183), .out(n14183_0));
mux15 mux_9018 (.in({n14104_0, n10139_0, n10118_0, n10113_0, n10106_0, n10101_0, n10089_0, n10072_0, n10070_1/**/, n10008_2, n7520, n7512, n6540, n6532, n6524}), .out(n14184), .config_in(config_chain[34011:34006]), .config_rst(config_rst)); 
buffer_wire buffer_14184 (.in(n14184), .out(n14184_0));
mux15 mux_9019 (.in({n14273_1, n11191_0, n11175_0, n11161_0, n11154_0/**/, n11147_0, n11140_0, n11126_0, n11111_0, n11094_1, n7814, n7806, n6834, n6826, n6818}), .out(n14185), .config_in(config_chain[34017:34012]), .config_rst(config_rst)); 
buffer_wire buffer_14185 (.in(n14185), .out(n14185_0));
mux15 mux_9020 (.in({n14112_0, n10141_0, n10126_0, n10121_0, n10109_0, n10092_0, n10080_0, n10075_0, n10068_1/**/, n10010_2, n7520, n7512, n7504, n6532, n6524}), .out(n14186), .config_in(config_chain[34023:34018]), .config_rst(config_rst)); 
buffer_wire buffer_14186 (.in(n14186), .out(n14186_0));
mux15 mux_9021 (.in({n14275_1, n11189_0, n11169_0/**/, n11162_0, n11148_0, n11133_0, n11119_0, n11112_0, n11096_1, n11047_0, n7814, n7806, n7798, n6826, n6818}), .out(n14187), .config_in(config_chain[34029:34024]), .config_rst(config_rst)); 
buffer_wire buffer_14187 (.in(n14187), .out(n14187_0));
mux14 mux_9022 (.in({n14120_0/**/, n10143_0, n10129_0, n10112_0, n10100_0, n10095_0, n10088_0, n10083_0, n10066_1, n7520, n7512, n7504, n6536, n6524}), .out(n14188), .config_in(config_chain[34035:34030]), .config_rst(config_rst)); 
buffer_wire buffer_14188 (.in(n14188), .out(n14188_0));
mux14 mux_9023 (.in({n14277_1, n11187_0, n11170_0, n11155_0, n11141_0, n11134_0, n11127_0, n11120_0, n11098_1, n7814, n7806, n7798, n6830, n6818}), .out(n14189), .config_in(config_chain[34041:34036]), .config_rst(config_rst)); 
buffer_wire buffer_14189 (.in(n14189), .out(n14189_0));
mux14 mux_9024 (.in({n14128_0, n10145_0, n10120_0, n10115_0, n10108_0, n10103_0, n10091_0, n10074_0, n10064_1, n7520, n7512, n7504/**/, n6536, n6528}), .out(n14190), .config_in(config_chain[34047:34042]), .config_rst(config_rst)); 
buffer_wire buffer_14190 (.in(n14190), .out(n14190_0));
mux14 mux_9025 (.in({n14279_1, n11185_0, n11163_0, n11156_0, n11149_0, n11142_0, n11128_0, n11113_0, n11100_1, n7814, n7806/**/, n7798, n6830, n6822}), .out(n14191), .config_in(config_chain[34053:34048]), .config_rst(config_rst)); 
buffer_wire buffer_14191 (.in(n14191), .out(n14191_0));
mux13 mux_9026 (.in({n14136_0, n10147_0, n10128_0/**/, n10123_0, n10111_0, n10094_0, n10082_0, n10077_0, n10062_1, n7512, n7504, n6536, n6528}), .out(n14192), .config_in(config_chain[34059:34054]), .config_rst(config_rst)); 
buffer_wire buffer_14192 (.in(n14192), .out(n14192_0));
mux13 mux_9027 (.in({n14281_1, n11183_0, n11171_0, n11164_0, n11150_0, n11135_0, n11121_0, n11114_0, n11102_1, n7806, n7798, n6830/**/, n6822}), .out(n14193), .config_in(config_chain[34065:34060]), .config_rst(config_rst)); 
buffer_wire buffer_14193 (.in(n14193), .out(n14193_0));
mux13 mux_9028 (.in({n14144_0/**/, n10149_0, n10131_0, n10114_0, n10102_0, n10097_0, n10090_0, n10085_0, n10060_1, n7516, n7504, n6536, n6528}), .out(n14194), .config_in(config_chain[34071:34066]), .config_rst(config_rst)); 
buffer_wire buffer_14194 (.in(n14194), .out(n14194_0));
mux13 mux_9029 (.in({n14283_1, n11181_0, n11172_0, n11157_0, n11143_0, n11136_0, n11129_0, n11122_0, n11104_1/**/, n7810, n7798, n6830, n6822}), .out(n14195), .config_in(config_chain[34077:34072]), .config_rst(config_rst)); 
buffer_wire buffer_14195 (.in(n14195), .out(n14195_0));
mux13 mux_9030 (.in({n14152_0, n10151_0, n10122_0, n10117_0, n10110_0, n10105_0, n10076_0, n10058_1/**/, n10003_0, n7516, n7508, n6536, n6528}), .out(n14196), .config_in(config_chain[34083:34078]), .config_rst(config_rst)); 
buffer_wire buffer_14196 (.in(n14196), .out(n14196_0));
mux13 mux_9031 (.in({n14285_1, n11179_0, n11165_0, n11158_0, n11151_0, n11144_0, n11115_0, n11108_1/**/, n11106_1, n7810, n7802, n6830, n6822}), .out(n14197), .config_in(config_chain[34089:34084]), .config_rst(config_rst)); 
buffer_wire buffer_14197 (.in(n14197), .out(n14197_0));
mux13 mux_9032 (.in({n14160_0, n10153_0, n10130_0, n10125_0, n10096_0, n10084_0, n10079_0, n10056_1/**/, n10005_0, n7516, n7508, n6540, n6528}), .out(n14198), .config_in(config_chain[34095:34090]), .config_rst(config_rst)); 
buffer_wire buffer_14198 (.in(n14198), .out(n14198_0));
mux13 mux_9033 (.in({n14287_1, n11177_0, n11173_0, n11166_0, n11137_0, n11130_0, n11123_0, n11116_0, n11044_2, n7810, n7802, n6834, n6822}), .out(n14199), .config_in(config_chain[34101:34096]), .config_rst(config_rst)); 
buffer_wire buffer_14199 (.in(n14199), .out(n14199_0));
mux13 mux_9034 (.in({n14168_0, n10133_0, n10116_0/**/, n10104_0, n10099_0, n10087_0, n10054_1, n10007_0, n10002_2, n7516, n7508, n6540, n6532}), .out(n14200), .config_in(config_chain[34107:34102]), .config_rst(config_rst)); 
buffer_wire buffer_14200 (.in(n14200), .out(n14200_0));
mux3 mux_9035 (.in({n12091_0/**/, n12090_2, n8202}), .out(n14201), .config_in(config_chain[34109:34108]), .config_rst(config_rst)); 
buffer_wire buffer_14201 (.in(n14201), .out(n14201_0));
mux15 mux_9036 (.in({n14090_0, n10393_0, n10374_0, n10369_0, n10360_0, n10355_0, n10343_0, n10308_1, n10265_0, n10260_2, n7614, n7606, n6638, n6630, n6622}), .out(n14202), .config_in(config_chain[34115:34110]), .config_rst(config_rst)); 
buffer_wire buffer_14202 (.in(n14202), .out(n14202_0));
mux15 mux_9037 (.in({n14291_0, n11461_0/**/, n11427_0, n11420_0, n11418_0, n11411_0, n11404_0, n11390_0, n11375_0, n11356_1, n7908, n7900, n6932, n6924, n6916}), .out(n14203), .config_in(config_chain[34121:34116]), .config_rst(config_rst)); 
buffer_wire buffer_14203 (.in(n14203), .out(n14203_0));
mux15 mux_9038 (.in({n14098_0, n10395_0, n10382_0, n10377_0, n10363_0/**/, n10334_0, n10329_0, n10267_0, n10262_2, n10258_2, n7618, n7606, n6638, n6630, n6622}), .out(n14204), .config_in(config_chain[34127:34122]), .config_rst(config_rst)); 
buffer_wire buffer_14204 (.in(n14204), .out(n14204_0));
mux15 mux_9039 (.in({n14293_0, n11459_0, n11440_0, n11435_0, n11428_0, n11412_0, n11397_0, n11383_0, n11376_0, n11358_1/**/, n7912, n7900, n6932, n6924, n6916}), .out(n14205), .config_in(config_chain[34133:34128]), .config_rst(config_rst)); 
buffer_wire buffer_14205 (.in(n14205), .out(n14205_0));
mux15 mux_9040 (.in({n14106_0, n10397_0, n10385_0, n10368_0/**/, n10354_0, n10349_0, n10342_0, n10337_0, n10326_1, n10264_2, n7618, n7610, n6638, n6630, n6622}), .out(n14206), .config_in(config_chain[34139:34134]), .config_rst(config_rst)); 
buffer_wire buffer_14206 (.in(n14206), .out(n14206_0));
mux15 mux_9041 (.in({n14295_0/**/, n11457_0, n11436_0, n11421_0, n11419_0, n11405_0, n11398_0, n11391_0, n11384_0, n11360_1, n7912, n7904, n6932, n6924, n6916}), .out(n14207), .config_in(config_chain[34145:34140]), .config_rst(config_rst)); 
buffer_wire buffer_14207 (.in(n14207), .out(n14207_0));
mux15 mux_9042 (.in({n14114_0, n10399_0, n10376_0, n10371_0, n10362_0, n10357_0, n10345_0, n10328_0, n10324_1, n10266_2, n7618, n7610, n7602, n6630, n6622}), .out(n14208), .config_in(config_chain[34151:34146]), .config_rst(config_rst)); 
buffer_wire buffer_14208 (.in(n14208), .out(n14208_0));
mux15 mux_9043 (.in({n14297_0, n11455_0, n11441_0, n11429_0, n11422_0, n11413_0, n11406_0, n11392_0, n11377_0, n11362_1/**/, n7912, n7904, n7896, n6924, n6916}), .out(n14209), .config_in(config_chain[34157:34152]), .config_rst(config_rst)); 
buffer_wire buffer_14209 (.in(n14209), .out(n14209_0));
mux14 mux_9044 (.in({n14122_0, n10401_0, n10384_0, n10379_0, n10365_0, n10348_0, n10336_0, n10331_0, n10322_1/**/, n7618, n7610, n7602, n6634, n6622}), .out(n14210), .config_in(config_chain[34163:34158]), .config_rst(config_rst)); 
buffer_wire buffer_14210 (.in(n14210), .out(n14210_0));
mux14 mux_9045 (.in({n14299_0, n11453_0, n11437_0, n11430_0, n11414_0/**/, n11399_0, n11385_0, n11378_0, n11364_1, n7912, n7904, n7896, n6928, n6916}), .out(n14211), .config_in(config_chain[34169:34164]), .config_rst(config_rst)); 
buffer_wire buffer_14211 (.in(n14211), .out(n14211_0));
mux14 mux_9046 (.in({n14130_0, n10403_0, n10387_0, n10370_0, n10356_0, n10351_0, n10344_0, n10339_0, n10320_1, n7618, n7610/**/, n7602, n6634, n6626}), .out(n14212), .config_in(config_chain[34175:34170]), .config_rst(config_rst)); 
buffer_wire buffer_14212 (.in(n14212), .out(n14212_0));
mux14 mux_9047 (.in({n14301_0, n11451_0, n11438_0, n11423_0, n11407_0, n11400_0, n11393_0, n11386_0, n11366_1, n7912/**/, n7904, n7896, n6928, n6920}), .out(n14213), .config_in(config_chain[34181:34176]), .config_rst(config_rst)); 
buffer_wire buffer_14213 (.in(n14213), .out(n14213_0));
mux13 mux_9048 (.in({n14138_0, n10405_0, n10378_0, n10373_0, n10364_0, n10359_0, n10347_0, n10330_0, n10318_1, n7610, n7602/**/, n6634, n6626}), .out(n14214), .config_in(config_chain[34187:34182]), .config_rst(config_rst)); 
buffer_wire buffer_14214 (.in(n14214), .out(n14214_0));
mux13 mux_9049 (.in({n14303_0, n11449_0, n11431_0, n11424_0, n11415_0, n11408_0, n11394_0, n11379_0, n11368_1, n7904, n7896, n6928, n6920/**/}), .out(n14215), .config_in(config_chain[34193:34188]), .config_rst(config_rst)); 
buffer_wire buffer_14215 (.in(n14215), .out(n14215_0));
mux13 mux_9050 (.in({n14146_0, n10407_0, n10386_0, n10381_0, n10367_0, n10350_0/**/, n10338_0, n10333_0, n10316_1, n7614, n7602, n6634, n6626}), .out(n14216), .config_in(config_chain[34199:34194]), .config_rst(config_rst)); 
buffer_wire buffer_14216 (.in(n14216), .out(n14216_0));
mux13 mux_9051 (.in({n14305_0, n11447_0, n11439_0, n11432_0/**/, n11416_0, n11401_0, n11387_0, n11380_0, n11370_1, n7908, n7896, n6928, n6920}), .out(n14217), .config_in(config_chain[34205:34200]), .config_rst(config_rst)); 
buffer_wire buffer_14217 (.in(n14217), .out(n14217_0));
mux13 mux_9052 (.in({n14154_0, n10409_0, n10389_0, n10372_0, n10358_0, n10353_0, n10346_0, n10341_0, n10314_1, n7614, n7606, n6634, n6626}), .out(n14218), .config_in(config_chain[34211:34206]), .config_rst(config_rst)); 
buffer_wire buffer_14218 (.in(n14218), .out(n14218_0));
mux13 mux_9053 (.in({n14307_0, n11445_0, n11425_0, n11409_0, n11402_0, n11395_0, n11388_0, n11372_1, n11352_1, n7908, n7900, n6928, n6920}), .out(n14219), .config_in(config_chain[34217:34212]), .config_rst(config_rst)); 
buffer_wire buffer_14219 (.in(n14219), .out(n14219_0));
mux13 mux_9054 (.in({n14162_0, n10411_0, n10380_0, n10375_0/**/, n10366_0, n10361_0, n10332_0, n10312_1, n10261_0, n7614, n7606, n6638, n6626}), .out(n14220), .config_in(config_chain[34223:34218]), .config_rst(config_rst)); 
buffer_wire buffer_14220 (.in(n14220), .out(n14220_0));
mux13 mux_9055 (.in({n14309_0/**/, n11443_0, n11433_0, n11426_0, n11417_0, n11410_0, n11381_0, n11374_1, n11310_2, n7908, n7900, n6932, n6920}), .out(n14221), .config_in(config_chain[34229:34224]), .config_rst(config_rst)); 
buffer_wire buffer_14221 (.in(n14221), .out(n14221_0));
mux13 mux_9056 (.in({n14170_0, n10391_0, n10388_0, n10383_0, n10352_0, n10340_0, n10335_0, n10310_1, n10263_0, n7614, n7606, n6638, n6630}), .out(n14222), .config_in(config_chain[34235:34230]), .config_rst(config_rst)); 
buffer_wire buffer_14222 (.in(n14222), .out(n14222_0));
mux3 mux_9057 (.in({n12093_0, n12092_2, n8202}), .out(n14223), .config_in(config_chain[34237:34236]), .config_rst(config_rst)); 
buffer_wire buffer_14223 (.in(n14223), .out(n14223_0));
mux15 mux_9058 (.in({n14092_0/**/, n10653_0, n10648_0, n10643_0, n10612_0, n10607_0, n10598_0, n10593_0, n10566_1, n10523_0, n7712, n7704, n6736, n6728, n6720}), .out(n14224), .config_in(config_chain[34243:34238]), .config_rst(config_rst)); 
buffer_wire buffer_14224 (.in(n14224), .out(n14224_0));
mux16 mux_9059 (.in({n14313_0/**/, n11725_0, n11692_0, n11689_0, n11685_0, n11681_0, n11664_0, n11654_0, n11651_0, n11622_1, n11596_1, n8006, n7998, n7030, n7022, n7014}), .out(n14225), .config_in(config_chain[34249:34244]), .config_rst(config_rst)); 
buffer_wire buffer_14225 (.in(n14225), .out(n14225_0));
mux15 mux_9060 (.in({n14100_0/**/, n10655_0, n10634_0, n10629_0, n10620_0, n10615_0, n10601_0, n10525_0, n10520_2, n10518_2, n7716, n7704, n6736, n6728, n6720}), .out(n14226), .config_in(config_chain[34255:34250]), .config_rst(config_rst)); 
buffer_wire buffer_14226 (.in(n14226), .out(n14226_0));
mux16 mux_9061 (.in({n14315_0, n11723_0, n11707_0, n11703_0, n11686_0/**/, n11678_0, n11675_0, n11648_0, n11645_0, n11624_1, n11618_1, n8006, n7998, n7030, n7022, n7014}), .out(n14227), .config_in(config_chain[34261:34256]), .config_rst(config_rst)); 
buffer_wire buffer_14227 (.in(n14227), .out(n14227_0));
mux15 mux_9062 (.in({n14108_0, n10657_0, n10642_0, n10637_0, n10623_0, n10606_0, n10592_0, n10587_0/**/, n10584_1, n10522_2, n7716, n7708, n6736, n6728, n6720}), .out(n14228), .config_in(config_chain[34267:34262]), .config_rst(config_rst)); 
buffer_wire buffer_14228 (.in(n14228), .out(n14228_0));
mux15 mux_9063 (.in({n14317_0, n11721_0, n11700_0, n11697_0, n11672_0, n11669_0, n11659_0, n11642_0, n11640_1, n11626_1, n8006, n7998, n7030, n7022, n7014}), .out(n14229), .config_in(config_chain[34273:34268]), .config_rst(config_rst)); 
buffer_wire buffer_14229 (.in(n14229), .out(n14229_0));
mux15 mux_9064 (.in({n14116_0, n10659_0, n10645_0, n10628_0, n10614_0, n10609_0, n10600_0, n10595_0, n10582_1, n10524_2, n7716/**/, n7708, n7700, n6728, n6720}), .out(n14230), .config_in(config_chain[34279:34274]), .config_rst(config_rst)); 
buffer_wire buffer_14230 (.in(n14230), .out(n14230_0));
mux15 mux_9065 (.in({n14319_0, n11719_0/**/, n11694_0, n11691_0, n11683_0, n11666_0, n11662_0, n11656_0, n11653_0, n11628_1, n8006, n7998, n7030, n7022, n7014}), .out(n14231), .config_in(config_chain[34285:34280]), .config_rst(config_rst)); 
buffer_wire buffer_14231 (.in(n14231), .out(n14231_0));
mux14 mux_9066 (.in({n14124_0, n10661_0, n10636_0/**/, n10631_0, n10622_0, n10617_0, n10603_0, n10586_0, n10580_1, n7716, n7708, n7700, n6732, n6720}), .out(n14232), .config_in(config_chain[34291:34286]), .config_rst(config_rst)); 
buffer_wire buffer_14232 (.in(n14232), .out(n14232_0));
mux15 mux_9067 (.in({n14321_0, n11717_0, n11705_0/**/, n11688_0, n11684_0, n11680_0, n11677_0, n11650_0, n11647_0, n11630_1, n8006, n7998, n7030, n7022, n7014}), .out(n14233), .config_in(config_chain[34297:34292]), .config_rst(config_rst)); 
buffer_wire buffer_14233 (.in(n14233), .out(n14233_0));
mux14 mux_9068 (.in({n14132_0/**/, n10663_0, n10644_0, n10639_0, n10625_0, n10608_0, n10594_0, n10589_0, n10578_1, n7716, n7708, n7700, n6732, n6724}), .out(n14234), .config_in(config_chain[34303:34298]), .config_rst(config_rst)); 
buffer_wire buffer_14234 (.in(n14234), .out(n14234_0));
mux15 mux_9069 (.in({n14323_0, n11715_0, n11706_0, n11702_0, n11699_0, n11674_0, n11671_0, n11661_0/**/, n11644_0, n11632_1, n8010, n8002, n7994, n7026, n7018}), .out(n14235), .config_in(config_chain[34309:34304]), .config_rst(config_rst)); 
buffer_wire buffer_14235 (.in(n14235), .out(n14235_0));
mux13 mux_9070 (.in({n14140_0, n10665_0, n10647_0, n10630_0/**/, n10616_0, n10611_0, n10602_0, n10597_0, n10576_1, n7708, n7700, n6732, n6724}), .out(n14236), .config_in(config_chain[34315:34310]), .config_rst(config_rst)); 
buffer_wire buffer_14236 (.in(n14236), .out(n14236_0));
mux15 mux_9071 (.in({n14325_0, n11713_0, n11696_0, n11693_0, n11668_0, n11665_0/**/, n11658_0, n11655_0, n11634_1, n11597_0, n8010, n8002, n7994, n7026, n7018}), .out(n14237), .config_in(config_chain[34321:34316]), .config_rst(config_rst)); 
buffer_wire buffer_14237 (.in(n14237), .out(n14237_0));
mux13 mux_9072 (.in({n14148_0, n10667_0, n10638_0, n10633_0, n10624_0, n10619_0, n10605_0, n10588_0, n10574_1, n7712, n7700, n6732, n6724}), .out(n14238), .config_in(config_chain[34327:34322]), .config_rst(config_rst)); 
buffer_wire buffer_14238 (.in(n14238), .out(n14238_0));
mux15 mux_9073 (.in({n14327_0, n11711_0, n11690_0, n11687_0, n11682_0/**/, n11679_0, n11652_0, n11649_0, n11636_1, n11619_0, n8010, n8002, n7994, n7026, n7018}), .out(n14239), .config_in(config_chain[34333:34328]), .config_rst(config_rst)); 
buffer_wire buffer_14239 (.in(n14239), .out(n14239_0));
mux13 mux_9074 (.in({n14156_0, n10669_0, n10646_0, n10641_0/**/, n10627_0, n10610_0, n10596_0, n10591_0, n10572_1, n7712, n7704, n6732, n6724}), .out(n14240), .config_in(config_chain[34339:34334]), .config_rst(config_rst)); 
buffer_wire buffer_14240 (.in(n14240), .out(n14240_0));
mux15 mux_9075 (.in({n14329_0, n11709_0, n11704_0, n11701_0, n11676_0, n11673_0, n11646_0, n11643_0, n11641_0, n11638_1, n8010, n8002, n7994, n7026, n7018}), .out(n14241), .config_in(config_chain[34345:34340]), .config_rst(config_rst)); 
buffer_wire buffer_14241 (.in(n14241), .out(n14241_0));
mux13 mux_9076 (.in({n14164_0, n10671_0, n10649_0, n10632_0, n10618_0, n10613_0, n10604_0, n10599_0, n10570_1, n7712, n7704, n6736/**/, n6724}), .out(n14242), .config_in(config_chain[34351:34346]), .config_rst(config_rst)); 
buffer_wire buffer_14242 (.in(n14242), .out(n14242_0));
mux15 mux_9077 (.in({n14331_0, n11727_0, n11698_0, n11695_0, n11670_0, n11667_0, n11663_0, n11660_0, n11657_0, n11620_1, n8010/**/, n8002, n7994, n7026, n7018}), .out(n14243), .config_in(config_chain[34357:34352]), .config_rst(config_rst)); 
buffer_wire buffer_14243 (.in(n14243), .out(n14243_0));
mux13 mux_9078 (.in({n14172_0, n10651_0, n10640_0, n10635_0, n10626_0, n10621_0, n10590_0/**/, n10568_1, n10521_0, n7712, n7704, n6736, n6728}), .out(n14244), .config_in(config_chain[34363:34358]), .config_rst(config_rst)); 
buffer_wire buffer_14244 (.in(n14244), .out(n14244_0));
mux3 mux_9079 (.in({n12123_0, n12122_1, n8202}), .out(n14245), .config_in(config_chain[34365:34364]), .config_rst(config_rst)); 
buffer_wire buffer_14245 (.in(n14245), .out(n14245_0));
mux15 mux_9080 (.in({n14094_1, n10915_0, n10902_0, n10897_0, n10888_0, n10883_0, n10852_0, n10847_0, n10826_1, n10783_0, n7810, n7802, n6834/**/, n6826, n6818}), .out(n14246), .config_in(config_chain[34371:34366]), .config_rst(config_rst)); 
buffer_wire buffer_14246 (.in(n14246), .out(n14246_0));
mux16 mux_9081 (.in({n14333_0, n11987_0, n11962_0, n11959_0, n11934_0, n11931_0, n11927_0, n11923_0, n11906_0/**/, n11886_1, n11828_2, n8104, n8096, n7128, n7120, n7112}), .out(n14247), .config_in(config_chain[34377:34372]), .config_rst(config_rst)); 
buffer_wire buffer_14247 (.in(n14247), .out(n14247_0));
mux15 mux_9082 (.in({n14102_1, n10917_0, n10910_0, n10905_0, n10874_0, n10869_0, n10860_0, n10855_0, n10785_0, n10780_2, n7814, n7802, n6834, n6826, n6818/**/}), .out(n14248), .config_in(config_chain[34383:34378]), .config_rst(config_rst)); 
buffer_wire buffer_14248 (.in(n14248), .out(n14248_0));
mux16 mux_9083 (.in({n14335_0, n11985_0, n11956_0, n11953_0, n11949_0, n11945_0, n11928_0, n11920_0/**/, n11917_0, n11888_1, n11860_1, n8104, n8096, n7128, n7120, n7112}), .out(n14249), .config_in(config_chain[34389:34384]), .config_rst(config_rst)); 
buffer_wire buffer_14249 (.in(n14249), .out(n14249_0));
mux15 mux_9084 (.in({n14110_1, n10919_0, n10896_0, n10891_0, n10882_0, n10877_0, n10863_0, n10846_0, n10844_1, n10782_2, n7814, n7806, n6834, n6826, n6818/**/}), .out(n14250), .config_in(config_chain[34395:34390]), .config_rst(config_rst)); 
buffer_wire buffer_14250 (.in(n14250), .out(n14250_0));
mux15 mux_9085 (.in({n14337_0, n11983_0, n11967_0, n11950_0, n11942_0, n11939_0, n11914_0, n11911_0, n11890_1/**/, n11882_1, n8104, n8096, n7128, n7120, n7112}), .out(n14251), .config_in(config_chain[34401:34396]), .config_rst(config_rst)); 
buffer_wire buffer_14251 (.in(n14251), .out(n14251_0));
mux15 mux_9086 (.in({n14118_1, n10921_0, n10904_0, n10899_0, n10885_0, n10868_0, n10854_0, n10849_0, n10842_1/**/, n10784_2, n7814, n7806, n7798, n6826, n6818}), .out(n14252), .config_in(config_chain[34407:34402]), .config_rst(config_rst)); 
buffer_wire buffer_14252 (.in(n14252), .out(n14252_0));
mux15 mux_9087 (.in({n14339_0, n11981_0/**/, n11964_0, n11961_0, n11936_0, n11933_0, n11925_0, n11908_0, n11904_1, n11892_1, n8104, n8096, n7128, n7120, n7112}), .out(n14253), .config_in(config_chain[34413:34408]), .config_rst(config_rst)); 
buffer_wire buffer_14253 (.in(n14253), .out(n14253_0));
mux14 mux_9088 (.in({n14126_1, n10923_0, n10907_0, n10890_0, n10876_0/**/, n10871_0, n10862_0, n10857_0, n10840_1, n7814, n7806, n7798, n6830, n6818}), .out(n14254), .config_in(config_chain[34419:34414]), .config_rst(config_rst)); 
buffer_wire buffer_14254 (.in(n14254), .out(n14254_0));
mux15 mux_9089 (.in({n14341_0/**/, n11979_0, n11958_0, n11955_0, n11947_0, n11930_0, n11926_0, n11922_0, n11919_0, n11894_1, n8104, n8096, n7128, n7120, n7112}), .out(n14255), .config_in(config_chain[34425:34420]), .config_rst(config_rst)); 
buffer_wire buffer_14255 (.in(n14255), .out(n14255_0));
mux14 mux_9090 (.in({n14134_1, n10925_0, n10898_0, n10893_0, n10884_0, n10879_0, n10865_0, n10848_0, n10838_1, n7814, n7806, n7798/**/, n6830, n6822}), .out(n14256), .config_in(config_chain[34431:34426]), .config_rst(config_rst)); 
buffer_wire buffer_14256 (.in(n14256), .out(n14256_0));
mux15 mux_9091 (.in({n14343_0, n11977_0, n11969_0/**/, n11952_0, n11948_0, n11944_0, n11941_0, n11916_0, n11913_0, n11896_1, n8108, n8100, n8092, n7124, n7116}), .out(n14257), .config_in(config_chain[34437:34432]), .config_rst(config_rst)); 
buffer_wire buffer_14257 (.in(n14257), .out(n14257_0));
mux13 mux_9092 (.in({n14142_1, n10927_0, n10906_0, n10901_0, n10887_0, n10870_0, n10856_0, n10851_0, n10836_1, n7806, n7798/**/, n6830, n6822}), .out(n14258), .config_in(config_chain[34443:34438]), .config_rst(config_rst)); 
buffer_wire buffer_14258 (.in(n14258), .out(n14258_0));
mux15 mux_9093 (.in({n14345_0, n11975_0, n11966_0, n11963_0, n11938_0, n11935_0, n11910_0, n11907_0/**/, n11898_1, n11829_0, n8108, n8100, n8092, n7124, n7116}), .out(n14259), .config_in(config_chain[34449:34444]), .config_rst(config_rst)); 
buffer_wire buffer_14259 (.in(n14259), .out(n14259_0));
mux13 mux_9094 (.in({n14150_1, n10929_0/**/, n10909_0, n10892_0, n10878_0, n10873_0, n10864_0, n10859_0, n10834_1, n7810, n7798, n6830, n6822}), .out(n14260), .config_in(config_chain[34455:34450]), .config_rst(config_rst)); 
buffer_wire buffer_14260 (.in(n14260), .out(n14260_0));
mux15 mux_9095 (.in({n14347_0, n11973_0, n11960_0, n11957_0, n11932_0, n11929_0, n11924_0, n11921_0, n11900_1, n11861_0, n8108/**/, n8100, n8092, n7124, n7116}), .out(n14261), .config_in(config_chain[34461:34456]), .config_rst(config_rst)); 
buffer_wire buffer_14261 (.in(n14261), .out(n14261_0));
mux13 mux_9096 (.in({n14158_1/**/, n10931_0, n10900_0, n10895_0, n10886_0, n10881_0, n10867_0, n10850_0, n10832_1, n7810, n7802, n6830, n6822}), .out(n14262), .config_in(config_chain[34467:34462]), .config_rst(config_rst)); 
buffer_wire buffer_14262 (.in(n14262), .out(n14262_0));
mux15 mux_9097 (.in({n14349_0, n11971_0, n11954_0, n11951_0, n11946_0, n11943_0, n11918_0/**/, n11915_0, n11902_1, n11883_0, n8108, n8100, n8092, n7124, n7116}), .out(n14263), .config_in(config_chain[34473:34468]), .config_rst(config_rst)); 
buffer_wire buffer_14263 (.in(n14263), .out(n14263_0));
mux13 mux_9098 (.in({n14166_1, n10933_0, n10908_0, n10903_0, n10889_0, n10872_0, n10858_0, n10853_0, n10830_1, n7810, n7802, n6834/**/, n6822}), .out(n14264), .config_in(config_chain[34479:34474]), .config_rst(config_rst)); 
buffer_wire buffer_14264 (.in(n14264), .out(n14264_0));
mux15 mux_9099 (.in({n14351_0, n11989_0, n11968_0, n11965_0, n11940_0, n11937_0, n11912_0/**/, n11909_0, n11905_0, n11884_1, n8108, n8100, n8092, n7124, n7116}), .out(n14265), .config_in(config_chain[34485:34480]), .config_rst(config_rst)); 
buffer_wire buffer_14265 (.in(n14265), .out(n14265_0));
mux13 mux_9100 (.in({n14174_1, n10913_0, n10911_0, n10894_0, n10880_0, n10875_0, n10866_0, n10861_0, n10828_1/**/, n7810, n7802, n6834, n6826}), .out(n14266), .config_in(config_chain[34491:34486]), .config_rst(config_rst)); 
buffer_wire buffer_14266 (.in(n14266), .out(n14266_0));
mux3 mux_9101 (.in({n12145_0, n12144_1/**/, n8202}), .out(n14267), .config_in(config_chain[34493:34492]), .config_rst(config_rst)); 
buffer_wire buffer_14267 (.in(n14267), .out(n14267_0));
mux15 mux_9102 (.in({n14180_1, n11179_0, n11175_0, n11166_0, n11161_0, n11147_0, n11130_0, n11116_0, n11111_0/**/, n11088_1, n7908, n7900, n6932, n6924, n6916}), .out(n14268), .config_in(config_chain[34499:34494]), .config_rst(config_rst)); 
buffer_wire buffer_14268 (.in(n14268), .out(n14268_0));
mux4 mux_9103 (.in({n12231_0, n12146_1, n8206/**/, n7210}), .out(n14269), .config_in(config_chain[34501:34500]), .config_rst(config_rst)); 
buffer_wire buffer_14269 (.in(n14269), .out(n14269_0));
mux15 mux_9104 (.in({n14182_1, n11181_0, n11169_0, n11152_0/**/, n11138_0, n11133_0, n11124_0, n11119_0, n11047_0, n11044_2, n7912, n7900, n6932, n6924, n6916}), .out(n14270), .config_in(config_chain[34507:34502]), .config_rst(config_rst)); 
buffer_wire buffer_14270 (.in(n14270), .out(n14270_0));
mux3 mux_9105 (.in({n12233_0, n12148_1/**/, n7210}), .out(n14271), .config_in(config_chain[34509:34508]), .config_rst(config_rst)); 
buffer_wire buffer_14271 (.in(n14271), .out(n14271_0));
mux15 mux_9106 (.in({n14184_1, n11183_0, n11174_0, n11160_0, n11155_0, n11146_0, n11141_0, n11127_0, n11110_0, n11106_1, n7912, n7904, n6932/**/, n6924, n6916}), .out(n14272), .config_in(config_chain[34515:34510]), .config_rst(config_rst)); 
buffer_wire buffer_14272 (.in(n14272), .out(n14272_0));
mux3 mux_9107 (.in({n12235_0/**/, n12150_1, n7214}), .out(n14273), .config_in(config_chain[34517:34516]), .config_rst(config_rst)); 
buffer_wire buffer_14273 (.in(n14273), .out(n14273_0));
mux15 mux_9108 (.in({n14186_1, n11185_0, n11168_0, n11163_0, n11149_0, n11132_0, n11118_0, n11113_0, n11104_1/**/, n11046_2, n7912, n7904, n7896, n6924, n6916}), .out(n14274), .config_in(config_chain[34523:34518]), .config_rst(config_rst)); 
buffer_wire buffer_14274 (.in(n14274), .out(n14274_0));
mux3 mux_9109 (.in({n12237_0/**/, n12152_1, n7218}), .out(n14275), .config_in(config_chain[34525:34524]), .config_rst(config_rst)); 
buffer_wire buffer_14275 (.in(n14275), .out(n14275_0));
mux14 mux_9110 (.in({n14188_1/**/, n11187_0, n11171_0, n11154_0, n11140_0, n11135_0, n11126_0, n11121_0, n11102_1, n7912, n7904, n7896, n6928, n6916}), .out(n14276), .config_in(config_chain[34531:34526]), .config_rst(config_rst)); 
buffer_wire buffer_14276 (.in(n14276), .out(n14276_0));
mux3 mux_9111 (.in({n12239_0, n12154_1, n7222}), .out(n14277), .config_in(config_chain[34533:34532]), .config_rst(config_rst)); 
buffer_wire buffer_14277 (.in(n14277), .out(n14277_0));
mux14 mux_9112 (.in({n14190_1, n11189_0, n11162_0, n11157_0, n11148_0/**/, n11143_0, n11129_0, n11112_0, n11100_1, n7912, n7904, n7896, n6928, n6920}), .out(n14278), .config_in(config_chain[34539:34534]), .config_rst(config_rst)); 
buffer_wire buffer_14278 (.in(n14278), .out(n14278_0));
mux3 mux_9113 (.in({n12241_0, n12156_1/**/, n7226}), .out(n14279), .config_in(config_chain[34541:34540]), .config_rst(config_rst)); 
buffer_wire buffer_14279 (.in(n14279), .out(n14279_0));
mux13 mux_9114 (.in({n14192_1, n11191_0, n11170_0, n11165_0, n11151_0, n11134_0, n11120_0, n11115_0, n11098_1, n7904/**/, n7896, n6928, n6920}), .out(n14280), .config_in(config_chain[34547:34542]), .config_rst(config_rst)); 
buffer_wire buffer_14280 (.in(n14280), .out(n14280_0));
mux3 mux_9115 (.in({n12243_0, n12158_1, n7226/**/}), .out(n14281), .config_in(config_chain[34549:34548]), .config_rst(config_rst)); 
buffer_wire buffer_14281 (.in(n14281), .out(n14281_0));
mux13 mux_9116 (.in({n14194_1/**/, n11193_0, n11173_0, n11156_0, n11142_0, n11137_0, n11128_0, n11123_0, n11096_1, n7908, n7896, n6928, n6920}), .out(n14282), .config_in(config_chain[34555:34550]), .config_rst(config_rst)); 
buffer_wire buffer_14282 (.in(n14282), .out(n14282_0));
mux3 mux_9117 (.in({n12245_0, n12160_1/**/, n8190}), .out(n14283), .config_in(config_chain[34557:34556]), .config_rst(config_rst)); 
buffer_wire buffer_14283 (.in(n14283), .out(n14283_0));
mux13 mux_9118 (.in({n14196_1, n11195_0, n11164_0, n11159_0, n11150_0, n11145_0, n11114_0, n11109_0, n11094_1, n7908, n7900, n6928, n6920/**/}), .out(n14284), .config_in(config_chain[34563:34558]), .config_rst(config_rst)); 
buffer_wire buffer_14284 (.in(n14284), .out(n14284_0));
mux3 mux_9119 (.in({n12247_0/**/, n12162_1, n8194}), .out(n14285), .config_in(config_chain[34565:34564]), .config_rst(config_rst)); 
buffer_wire buffer_14285 (.in(n14285), .out(n14285_0));
mux13 mux_9120 (.in({n14198_1, n11197_0, n11172_0, n11167_0, n11136_0/**/, n11131_0, n11122_0, n11117_0, n11092_1, n7908, n7900, n6932, n6920}), .out(n14286), .config_in(config_chain[34571:34566]), .config_rst(config_rst)); 
buffer_wire buffer_14286 (.in(n14286), .out(n14286_0));
mux3 mux_9121 (.in({n12249_0, n12164_1, n8198/**/}), .out(n14287), .config_in(config_chain[34573:34572]), .config_rst(config_rst)); 
buffer_wire buffer_14287 (.in(n14287), .out(n14287_0));
mux13 mux_9122 (.in({n14176_1, n11177_0, n11158_0, n11153_0, n11144_0, n11139_0, n11125_0, n11108_1, n11090_1, n7908, n7900, n6932, n6924}), .out(n14288), .config_in(config_chain[34579:34574]), .config_rst(config_rst)); 
buffer_wire buffer_14288 (.in(n14288), .out(n14288_0));
mux3 mux_9123 (.in({n12167_0, n12166_1, n8202}), .out(n14289), .config_in(config_chain[34581:34580]), .config_rst(config_rst)); 
buffer_wire buffer_14289 (.in(n14289), .out(n14289_0));
mux15 mux_9124 (.in({n14202_1, n11445_0, n11426_0, n11421_0, n11419_0, n11410_0, n11405_0/**/, n11391_0, n11374_1, n11354_1, n8006, n7998, n7030, n7022, n7014}), .out(n14290), .config_in(config_chain[34587:34582]), .config_rst(config_rst)); 
buffer_wire buffer_14290 (.in(n14290), .out(n14290_0));
mux4 mux_9125 (.in({n12169_0, n12168_0, n8206, n7210}), .out(n14291), .config_in(config_chain[34589:34588]), .config_rst(config_rst)); 
buffer_wire buffer_14291 (.in(n14291), .out(n14291_0));
mux15 mux_9126 (.in({n14204_1, n11447_0, n11441_0, n11434_0, n11429_0, n11413_0, n11396_0, n11382_0, n11377_0/**/, n11310_2, n8010, n7998, n7030, n7022, n7014}), .out(n14292), .config_in(config_chain[34595:34590]), .config_rst(config_rst)); 
buffer_wire buffer_14292 (.in(n14292), .out(n14292_0));
mux3 mux_9127 (.in({n12171_0, n12170_0, n7214}), .out(n14293), .config_in(config_chain[34597:34596]), .config_rst(config_rst)); 
buffer_wire buffer_14293 (.in(n14293), .out(n14293_0));
mux15 mux_9128 (.in({n14206_1, n11449_0, n11437_0, n11420_0/**/, n11418_0, n11404_0, n11399_0, n11390_0, n11385_0, n11372_1, n8010, n8002, n7030, n7022, n7014}), .out(n14294), .config_in(config_chain[34603:34598]), .config_rst(config_rst)); 
buffer_wire buffer_14294 (.in(n14294), .out(n14294_0));
mux3 mux_9129 (.in({n12173_0, n12172_0/**/, n7214}), .out(n14295), .config_in(config_chain[34605:34604]), .config_rst(config_rst)); 
buffer_wire buffer_14295 (.in(n14295), .out(n14295_0));
mux15 mux_9130 (.in({n14208_1, n11451_0, n11440_0, n11428_0, n11423_0, n11412_0, n11407_0, n11393_0, n11376_0, n11370_1/**/, n8010, n8002, n7994, n7022, n7014}), .out(n14296), .config_in(config_chain[34611:34606]), .config_rst(config_rst)); 
buffer_wire buffer_14296 (.in(n14296), .out(n14296_0));
mux3 mux_9131 (.in({n12175_0, n12174_0, n7218}), .out(n14297), .config_in(config_chain[34613:34612]), .config_rst(config_rst)); 
buffer_wire buffer_14297 (.in(n14297), .out(n14297_0));
mux14 mux_9132 (.in({n14210_1, n11453_0, n11436_0, n11431_0, n11415_0, n11398_0, n11384_0, n11379_0, n11368_1, n8010, n8002, n7994, n7026, n7014}), .out(n14298), .config_in(config_chain[34619:34614]), .config_rst(config_rst)); 
buffer_wire buffer_14298 (.in(n14298), .out(n14298_0));
mux3 mux_9133 (.in({n12177_0, n12176_0/**/, n7222}), .out(n14299), .config_in(config_chain[34621:34620]), .config_rst(config_rst)); 
buffer_wire buffer_14299 (.in(n14299), .out(n14299_0));
mux14 mux_9134 (.in({n14212_1, n11455_0, n11439_0, n11422_0, n11406_0/**/, n11401_0, n11392_0, n11387_0, n11366_1, n8010, n8002, n7994, n7026, n7018}), .out(n14300), .config_in(config_chain[34627:34622]), .config_rst(config_rst)); 
buffer_wire buffer_14300 (.in(n14300), .out(n14300_0));
mux3 mux_9135 (.in({n12179_0/**/, n12178_0, n7226}), .out(n14301), .config_in(config_chain[34629:34628]), .config_rst(config_rst)); 
buffer_wire buffer_14301 (.in(n14301), .out(n14301_0));
mux13 mux_9136 (.in({n14214_1, n11457_0, n11430_0, n11425_0, n11414_0, n11409_0, n11395_0, n11378_0, n11364_1, n8002, n7994, n7026/**/, n7018}), .out(n14302), .config_in(config_chain[34635:34630]), .config_rst(config_rst)); 
buffer_wire buffer_14302 (.in(n14302), .out(n14302_0));
mux3 mux_9137 (.in({n12181_0, n12180_0, n8190}), .out(n14303), .config_in(config_chain[34637:34636]), .config_rst(config_rst)); 
buffer_wire buffer_14303 (.in(n14303), .out(n14303_0));
mux13 mux_9138 (.in({n14216_1, n11459_0, n11438_0, n11433_0, n11417_0, n11400_0, n11386_0, n11381_0, n11362_1, n8006/**/, n7994, n7026, n7018}), .out(n14304), .config_in(config_chain[34643:34638]), .config_rst(config_rst)); 
buffer_wire buffer_14304 (.in(n14304), .out(n14304_0));
mux3 mux_9139 (.in({n12183_0, n12182_0, n8190}), .out(n14305), .config_in(config_chain[34645:34644]), .config_rst(config_rst)); 
buffer_wire buffer_14305 (.in(n14305), .out(n14305_0));
mux13 mux_9140 (.in({n14218_1, n11461_0, n11424_0/**/, n11408_0, n11403_0, n11394_0, n11389_0, n11360_1, n11353_0, n8006, n7998, n7026, n7018}), .out(n14306), .config_in(config_chain[34651:34646]), .config_rst(config_rst)); 
buffer_wire buffer_14306 (.in(n14306), .out(n14306_0));
mux3 mux_9141 (.in({n12185_0, n12184_0, n8194}), .out(n14307), .config_in(config_chain[34653:34652]), .config_rst(config_rst)); 
buffer_wire buffer_14307 (.in(n14307), .out(n14307_0));
mux13 mux_9142 (.in({n14220_1, n11463_0, n11432_0, n11427_0/**/, n11416_0, n11411_0, n11380_0, n11375_0, n11358_1, n8006, n7998, n7030, n7018}), .out(n14308), .config_in(config_chain[34659:34654]), .config_rst(config_rst)); 
buffer_wire buffer_14308 (.in(n14308), .out(n14308_0));
mux3 mux_9143 (.in({n12187_0/**/, n12186_0, n8198}), .out(n14309), .config_in(config_chain[34661:34660]), .config_rst(config_rst)); 
buffer_wire buffer_14309 (.in(n14309), .out(n14309_0));
mux13 mux_9144 (.in({n14178_1, n11443_0, n11435_0/**/, n11402_0, n11397_0, n11388_0, n11383_0, n11356_1, n11352_1, n8006, n7998, n7030, n7022}), .out(n14310), .config_in(config_chain[34667:34662]), .config_rst(config_rst)); 
buffer_wire buffer_14310 (.in(n14310), .out(n14310_0));
mux3 mux_9145 (.in({n12189_0, n12188_0/**/, n8206}), .out(n14311), .config_in(config_chain[34669:34668]), .config_rst(config_rst)); 
buffer_wire buffer_14311 (.in(n14311), .out(n14311_0));
mux16 mux_9146 (.in({n14224_1/**/, n11711_0, n11693_0, n11688_0, n11684_0, n11680_0, n11665_0, n11655_0, n11650_0, n11620_1, n11597_0, n8104, n8096, n7128, n7120, n7112}), .out(n14312), .config_in(config_chain[34675:34670]), .config_rst(config_rst)); 
buffer_wire buffer_14312 (.in(n14312), .out(n14312_0));
mux4 mux_9147 (.in({n12191_0, n12190_0/**/, n8206, n7210}), .out(n14313), .config_in(config_chain[34677:34676]), .config_rst(config_rst)); 
buffer_wire buffer_14313 (.in(n14313), .out(n14313_0));
mux16 mux_9148 (.in({n14226_1, n11713_0/**/, n11706_0, n11702_0, n11687_0, n11679_0, n11674_0, n11649_0, n11644_0, n11638_1, n11619_0, n8104, n8096, n7128, n7120, n7112}), .out(n14314), .config_in(config_chain[34683:34678]), .config_rst(config_rst)); 
buffer_wire buffer_14314 (.in(n14314), .out(n14314_0));
mux3 mux_9149 (.in({n12193_0, n12192_0/**/, n7214}), .out(n14315), .config_in(config_chain[34685:34684]), .config_rst(config_rst)); 
buffer_wire buffer_14315 (.in(n14315), .out(n14315_0));
mux15 mux_9150 (.in({n14228_1, n11715_0, n11701_0, n11696_0, n11673_0, n11668_0, n11658_0, n11643_0, n11641_0, n11636_1, n8104, n8096, n7128, n7120, n7112}), .out(n14316), .config_in(config_chain[34691:34686]), .config_rst(config_rst)); 
buffer_wire buffer_14316 (.in(n14316), .out(n14316_0));
mux3 mux_9151 (.in({n12195_0, n12194_0/**/, n7218}), .out(n14317), .config_in(config_chain[34693:34692]), .config_rst(config_rst)); 
buffer_wire buffer_14317 (.in(n14317), .out(n14317_0));
mux15 mux_9152 (.in({n14230_1, n11717_0, n11695_0, n11690_0/**/, n11682_0, n11667_0, n11663_0, n11657_0, n11652_0, n11634_1, n8104, n8096, n7128, n7120, n7112}), .out(n14318), .config_in(config_chain[34699:34694]), .config_rst(config_rst)); 
buffer_wire buffer_14318 (.in(n14318), .out(n14318_0));
mux3 mux_9153 (.in({n12197_0, n12196_0, n7218}), .out(n14319), .config_in(config_chain[34701:34700]), .config_rst(config_rst)); 
buffer_wire buffer_14319 (.in(n14319), .out(n14319_0));
mux15 mux_9154 (.in({n14232_1/**/, n11719_0, n11704_0, n11689_0, n11685_0, n11681_0, n11676_0, n11651_0, n11646_0, n11632_1, n8104, n8096, n7128, n7120, n7112}), .out(n14320), .config_in(config_chain[34707:34702]), .config_rst(config_rst)); 
buffer_wire buffer_14320 (.in(n14320), .out(n14320_0));
mux3 mux_9155 (.in({n12199_0, n12198_0, n7222}), .out(n14321), .config_in(config_chain[34709:34708]), .config_rst(config_rst)); 
buffer_wire buffer_14321 (.in(n14321), .out(n14321_0));
mux15 mux_9156 (.in({n14234_1, n11721_0, n11707_0, n11703_0, n11698_0, n11675_0, n11670_0, n11660_0, n11645_0, n11630_1/**/, n8108, n8100, n8092, n7124, n7116}), .out(n14322), .config_in(config_chain[34715:34710]), .config_rst(config_rst)); 
buffer_wire buffer_14322 (.in(n14322), .out(n14322_0));
mux3 mux_9157 (.in({n12201_0, n12200_0, n7226}), .out(n14323), .config_in(config_chain[34717:34716]), .config_rst(config_rst)); 
buffer_wire buffer_14323 (.in(n14323), .out(n14323_0));
mux15 mux_9158 (.in({n14236_1, n11723_0/**/, n11697_0, n11692_0, n11669_0, n11664_0, n11659_0, n11654_0, n11628_1, n11596_1, n8108, n8100, n8092, n7124, n7116}), .out(n14324), .config_in(config_chain[34723:34718]), .config_rst(config_rst)); 
buffer_wire buffer_14324 (.in(n14324), .out(n14324_0));
mux3 mux_9159 (.in({n12203_0, n12202_0, n8190}), .out(n14325), .config_in(config_chain[34725:34724]), .config_rst(config_rst)); 
buffer_wire buffer_14325 (.in(n14325), .out(n14325_0));
mux15 mux_9160 (.in({n14238_1, n11725_0, n11691_0/**/, n11686_0, n11683_0, n11678_0, n11653_0, n11648_0, n11626_1, n11618_1, n8108, n8100, n8092, n7124, n7116}), .out(n14326), .config_in(config_chain[34731:34726]), .config_rst(config_rst)); 
buffer_wire buffer_14326 (.in(n14326), .out(n14326_0));
mux3 mux_9161 (.in({n12205_0, n12204_0, n8194}), .out(n14327), .config_in(config_chain[34733:34732]), .config_rst(config_rst)); 
buffer_wire buffer_14327 (.in(n14327), .out(n14327_0));
mux15 mux_9162 (.in({n14240_1, n11727_0, n11705_0, n11700_0, n11677_0, n11672_0, n11647_0, n11642_0, n11640_1/**/, n11624_1, n8108, n8100, n8092, n7124, n7116}), .out(n14328), .config_in(config_chain[34739:34734]), .config_rst(config_rst)); 
buffer_wire buffer_14328 (.in(n14328), .out(n14328_0));
mux3 mux_9163 (.in({n12207_0, n12206_0, n8194}), .out(n14329), .config_in(config_chain[34741:34740]), .config_rst(config_rst)); 
buffer_wire buffer_14329 (.in(n14329), .out(n14329_0));
mux15 mux_9164 (.in({n14242_1, n11709_0, n11699_0, n11694_0, n11671_0, n11666_0, n11662_0/**/, n11661_0, n11656_0, n11622_1, n8108, n8100, n8092, n7124, n7116}), .out(n14330), .config_in(config_chain[34747:34742]), .config_rst(config_rst)); 
buffer_wire buffer_14330 (.in(n14330), .out(n14330_0));
mux3 mux_9165 (.in({n12209_0/**/, n12208_0, n8198}), .out(n14331), .config_in(config_chain[34749:34748]), .config_rst(config_rst)); 
buffer_wire buffer_14331 (.in(n14331), .out(n14331_0));
mux16 mux_9166 (.in({n14246_1, n11973_0, n11963_0, n11958_0, n11935_0, n11930_0, n11926_0, n11922_0/**/, n11907_0, n11884_1, n11829_0, n8202, n8194, n7226, n7218, n7210}), .out(n14332), .config_in(config_chain[34755:34750]), .config_rst(config_rst)); 
buffer_wire buffer_14332 (.in(n14332), .out(n14332_0));
mux4 mux_9167 (.in({n12211_0, n12210_0, n8206, n7210}), .out(n14333), .config_in(config_chain[34757:34756]), .config_rst(config_rst)); 
buffer_wire buffer_14333 (.in(n14333), .out(n14333_0));
mux16 mux_9168 (.in({n14248_1, n11975_0, n11957_0, n11952_0, n11948_0, n11944_0, n11929_0, n11921_0/**/, n11916_0, n11902_1, n11861_0, n8202, n8194, n7226, n7218, n7210}), .out(n14334), .config_in(config_chain[34763:34758]), .config_rst(config_rst)); 
buffer_wire buffer_14334 (.in(n14334), .out(n14334_0));
mux3 mux_9169 (.in({n12213_0, n12212_0, n7214}), .out(n14335), .config_in(config_chain[34765:34764]), .config_rst(config_rst)); 
buffer_wire buffer_14335 (.in(n14335), .out(n14335_0));
mux15 mux_9170 (.in({n14250_1, n11977_0, n11966_0, n11951_0, n11943_0, n11938_0/**/, n11915_0, n11910_0, n11900_1, n11883_0, n8202, n8194, n7226, n7218, n7210}), .out(n14336), .config_in(config_chain[34771:34766]), .config_rst(config_rst)); 
buffer_wire buffer_14336 (.in(n14336), .out(n14336_0));
mux3 mux_9171 (.in({n12215_0/**/, n12214_0, n7218}), .out(n14337), .config_in(config_chain[34773:34772]), .config_rst(config_rst)); 
buffer_wire buffer_14337 (.in(n14337), .out(n14337_0));
mux15 mux_9172 (.in({n14252_1, n11979_0, n11965_0, n11960_0, n11937_0, n11932_0, n11924_0, n11909_0, n11905_0, n11898_1, n8202, n8194, n7226, n7218, n7210}), .out(n14338), .config_in(config_chain[34779:34774]), .config_rst(config_rst)); 
buffer_wire buffer_14338 (.in(n14338), .out(n14338_0));
mux3 mux_9173 (.in({n12217_0, n12216_0/**/, n7222}), .out(n14339), .config_in(config_chain[34781:34780]), .config_rst(config_rst)); 
buffer_wire buffer_14339 (.in(n14339), .out(n14339_0));
mux15 mux_9174 (.in({n14254_1, n11981_0, n11959_0, n11954_0, n11946_0, n11931_0, n11927_0, n11923_0, n11918_0, n11896_1, n8202, n8194, n7226, n7218, n7210}), .out(n14340), .config_in(config_chain[34787:34782]), .config_rst(config_rst)); 
buffer_wire buffer_14340 (.in(n14340), .out(n14340_0));
mux3 mux_9175 (.in({n12219_0, n12218_0/**/, n7222}), .out(n14341), .config_in(config_chain[34789:34788]), .config_rst(config_rst)); 
buffer_wire buffer_14341 (.in(n14341), .out(n14341_0));
mux15 mux_9176 (.in({n14256_1, n11983_0, n11968_0, n11953_0, n11949_0, n11945_0/**/, n11940_0, n11917_0, n11912_0, n11894_1, n8206, n8198, n8190, n7222, n7214}), .out(n14342), .config_in(config_chain[34795:34790]), .config_rst(config_rst)); 
buffer_wire buffer_14342 (.in(n14342), .out(n14342_0));
mux3 mux_9177 (.in({n12221_0, n12220_0, n7226}), .out(n14343), .config_in(config_chain[34797:34796]), .config_rst(config_rst)); 
buffer_wire buffer_14343 (.in(n14343), .out(n14343_0));
mux15 mux_9178 (.in({n14258_1, n11985_0, n11967_0, n11962_0, n11939_0, n11934_0, n11911_0, n11906_0/**/, n11892_1, n11828_2, n8206, n8198, n8190, n7222, n7214}), .out(n14344), .config_in(config_chain[34803:34798]), .config_rst(config_rst)); 
buffer_wire buffer_14344 (.in(n14344), .out(n14344_0));
mux3 mux_9179 (.in({n12223_0, n12222_0, n8190}), .out(n14345), .config_in(config_chain[34805:34804]), .config_rst(config_rst)); 
buffer_wire buffer_14345 (.in(n14345), .out(n14345_0));
mux15 mux_9180 (.in({n14260_1, n11987_0, n11961_0, n11956_0, n11933_0, n11928_0, n11925_0/**/, n11920_0, n11890_1, n11860_1, n8206, n8198, n8190, n7222, n7214}), .out(n14346), .config_in(config_chain[34811:34806]), .config_rst(config_rst)); 
buffer_wire buffer_14346 (.in(n14346), .out(n14346_0));
mux3 mux_9181 (.in({n12225_0, n12224_0, n8194}), .out(n14347), .config_in(config_chain[34813:34812]), .config_rst(config_rst)); 
buffer_wire buffer_14347 (.in(n14347), .out(n14347_0));
mux15 mux_9182 (.in({n14262_1, n11989_0, n11955_0/**/, n11950_0, n11947_0, n11942_0, n11919_0, n11914_0, n11888_1, n11882_1, n8206, n8198, n8190, n7222, n7214}), .out(n14348), .config_in(config_chain[34819:34814]), .config_rst(config_rst)); 
buffer_wire buffer_14348 (.in(n14348), .out(n14348_0));
mux3 mux_9183 (.in({n12227_0, n12226_0, n8198}), .out(n14349), .config_in(config_chain[34821:34820]), .config_rst(config_rst)); 
buffer_wire buffer_14349 (.in(n14349), .out(n14349_0));
mux15 mux_9184 (.in({n14264_1, n11971_0, n11969_0, n11964_0, n11941_0, n11936_0, n11913_0, n11908_0, n11904_1, n11886_1, n8206, n8198, n8190/**/, n7222, n7214}), .out(n14350), .config_in(config_chain[34827:34822]), .config_rst(config_rst)); 
buffer_wire buffer_14350 (.in(n14350), .out(n14350_0));
mux3 mux_9185 (.in({n12229_0, n12228_0, n8198}), .out(n14351), .config_in(config_chain[34829:34828]), .config_rst(config_rst)); 
buffer_wire buffer_14351 (.in(n14351), .out(n14351_0));
mux4 mux_9186 (.in({n9899_0, n9818_1, n8400, n7404}), .out(n14352), .config_in(config_chain[34831:34830]), .config_rst(config_rst)); 
buffer_wire buffer_14352 (.in(n14352), .out(n14352_0));
mux15 mux_9187 (.in({n14511_1, n10953_0, n10932_0, n10925_0, n10918_0, n10904_0, n10889_0, n10875_0, n10868_0, n10848_1, n8690, n8682, n7714, n7706, n7698}), .out(n14353), .config_in(config_chain[34837:34832]), .config_rst(config_rst)); 
buffer_wire buffer_14353 (.in(n14353), .out(n14353_0));
mux4 mux_9188 (.in({n9839_0, n9838_0, n8400, n7404}), .out(n14354), .config_in(config_chain[34839:34838]), .config_rst(config_rst)); 
buffer_wire buffer_14354 (.in(n14354), .out(n14354_0));
mux15 mux_9189 (.in({n14445_1, n10173_0, n10139_0, n10132_0, n10125_0, n10118_0, n10106_0, n10074_1, n10008_2, n10005_0, n8396, n8388, n7420, n7412, n7404}), .out(n14355), .config_in(config_chain[34845:34840]), .config_rst(config_rst)); 
buffer_wire buffer_14355 (.in(n14355), .out(n14355_0));
mux4 mux_9190 (.in({n9859_0, n9858_0, n8400, n7404}), .out(n14356), .config_in(config_chain[34847:34846]), .config_rst(config_rst)); 
buffer_wire buffer_14356 (.in(n14356), .out(n14356_0));
mux15 mux_9191 (.in({n14467_1, n10431_0, n10411_0, n10404_0, n10375_0, n10368_0, n10361_0, n10354_0, n10330_1, n10264_2, n8494, n8486, n7518, n7510, n7502}), .out(n14357), .config_in(config_chain[34853:34848]), .config_rst(config_rst)); 
buffer_wire buffer_14357 (.in(n14357), .out(n14357_0));
mux4 mux_9192 (.in({n9879_0, n9878_0/**/, n8400, n7404}), .out(n14358), .config_in(config_chain[34855:34854]), .config_rst(config_rst)); 
buffer_wire buffer_14358 (.in(n14358), .out(n14358_0));
mux15 mux_9193 (.in({n14489_1, n10691_0, n10663_0, n10656_0, n10649_0, n10642_0, n10613_0, n10606_0, n10588_1, n10522_2, n8592, n8584, n7616, n7608, n7600}), .out(n14359), .config_in(config_chain[34861:34856]), .config_rst(config_rst)); 
buffer_wire buffer_14359 (.in(n14359), .out(n14359_0));
mux3 mux_9194 (.in({n9901_0, n9820_1/**/, n7404}), .out(n14360), .config_in(config_chain[34863:34862]), .config_rst(config_rst)); 
buffer_wire buffer_14360 (.in(n14360), .out(n14360_0));
mux15 mux_9195 (.in({n14513_1, n10951_0, n10926_0/**/, n10911_0, n10897_0, n10890_0, n10883_0, n10876_0, n10850_1, n10784_2, n8694, n8682, n7714, n7706, n7698}), .out(n14361), .config_in(config_chain[34869:34864]), .config_rst(config_rst)); 
buffer_wire buffer_14361 (.in(n14361), .out(n14361_0));
mux3 mux_9196 (.in({n9841_0, n9840_0, n7408}), .out(n14362), .config_in(config_chain[34871:34870]), .config_rst(config_rst)); 
buffer_wire buffer_14362 (.in(n14362), .out(n14362_0));
mux15 mux_9197 (.in({n14447_1, n10171_0, n10147_0, n10140_0, n10126_0, n10099_0, n10092_0, n10076_1, n10010_2, n10007_0, n8400, n8388, n7420, n7412, n7404}), .out(n14363), .config_in(config_chain[34877:34872]), .config_rst(config_rst)); 
buffer_wire buffer_14363 (.in(n14363), .out(n14363_0));
mux3 mux_9198 (.in({n9861_0, n9860_0, n7408}), .out(n14364), .config_in(config_chain[34879:34878]), .config_rst(config_rst)); 
buffer_wire buffer_14364 (.in(n14364), .out(n14364_0));
mux15 mux_9199 (.in({n14469_1, n10429_0, n10397_0, n10390_0/**/, n10383_0, n10376_0, n10362_0, n10332_1, n10266_2, n10263_0, n8498, n8486, n7518, n7510, n7502}), .out(n14365), .config_in(config_chain[34885:34880]), .config_rst(config_rst)); 
buffer_wire buffer_14365 (.in(n14365), .out(n14365_0));
mux3 mux_9200 (.in({n9881_0, n9880_0/**/, n7408}), .out(n14366), .config_in(config_chain[34887:34886]), .config_rst(config_rst)); 
buffer_wire buffer_14366 (.in(n14366), .out(n14366_0));
mux15 mux_9201 (.in({n14491_1, n10689_0, n10671_0, n10664_0, n10635_0, n10628_0, n10621_0, n10614_0, n10590_1, n10524_2, n8596, n8584, n7616, n7608, n7600}), .out(n14367), .config_in(config_chain[34893:34888]), .config_rst(config_rst)); 
buffer_wire buffer_14367 (.in(n14367), .out(n14367_0));
mux3 mux_9202 (.in({n9903_0, n9822_1, n7408}), .out(n14368), .config_in(config_chain[34895:34894]), .config_rst(config_rst)); 
buffer_wire buffer_14368 (.in(n14368), .out(n14368_0));
mux15 mux_9203 (.in({n14515_1, n10949_0, n10933_0, n10919_0, n10912_0, n10905_0, n10898_0, n10884_0, n10869_0, n10852_1, n8694, n8686, n7714, n7706, n7698}), .out(n14369), .config_in(config_chain[34901:34896]), .config_rst(config_rst)); 
buffer_wire buffer_14369 (.in(n14369), .out(n14369_0));
mux3 mux_9204 (.in({n9843_0, n9842_0, n7408}), .out(n14370), .config_in(config_chain[34903:34902]), .config_rst(config_rst)); 
buffer_wire buffer_14370 (.in(n14370), .out(n14370_0));
mux15 mux_9205 (.in({n14449_1, n10169_0, n10148_0, n10133_0, n10119_0, n10112_0, n10107_0, n10100_0, n10078_1, n10009_0, n8400, n8392, n7420, n7412, n7404}), .out(n14371), .config_in(config_chain[34909:34904]), .config_rst(config_rst)); 
buffer_wire buffer_14371 (.in(n14371), .out(n14371_0));
mux3 mux_9206 (.in({n9863_0, n9862_0, n7412}), .out(n14372), .config_in(config_chain[34911:34910]), .config_rst(config_rst)); 
buffer_wire buffer_14372 (.in(n14372), .out(n14372_0));
mux15 mux_9207 (.in({n14471_1, n10427_0, n10405_0, n10398_0, n10384_0, n10369_0, n10355_0, n10348_0, n10334_1, n10265_0, n8498, n8490, n7518, n7510, n7502}), .out(n14373), .config_in(config_chain[34917:34912]), .config_rst(config_rst)); 
buffer_wire buffer_14373 (.in(n14373), .out(n14373_0));
mux3 mux_9208 (.in({n9883_0, n9882_0/**/, n7412}), .out(n14374), .config_in(config_chain[34919:34918]), .config_rst(config_rst)); 
buffer_wire buffer_14374 (.in(n14374), .out(n14374_0));
mux15 mux_9209 (.in({n14493_1/**/, n10687_0, n10657_0, n10650_0, n10643_0, n10636_0, n10622_0, n10607_0, n10592_1, n10523_0, n8596, n8588, n7616, n7608, n7600}), .out(n14375), .config_in(config_chain[34925:34920]), .config_rst(config_rst)); 
buffer_wire buffer_14375 (.in(n14375), .out(n14375_0));
mux3 mux_9210 (.in({n9905_0, n9824_1/**/, n7412}), .out(n14376), .config_in(config_chain[34927:34926]), .config_rst(config_rst)); 
buffer_wire buffer_14376 (.in(n14376), .out(n14376_0));
mux15 mux_9211 (.in({n14517_1, n10947_0, n10927_0, n10920_0, n10906_0, n10891_0, n10877_0, n10870_0, n10854_1/**/, n10785_0, n8694, n8686, n8678, n7706, n7698}), .out(n14377), .config_in(config_chain[34933:34928]), .config_rst(config_rst)); 
buffer_wire buffer_14377 (.in(n14377), .out(n14377_0));
mux3 mux_9212 (.in({n9845_0, n9844_0, n7412}), .out(n14378), .config_in(config_chain[34935:34934]), .config_rst(config_rst)); 
buffer_wire buffer_14378 (.in(n14378), .out(n14378_0));
mux15 mux_9213 (.in({n14451_1, n10167_0, n10141_0, n10134_0, n10127_0, n10120_0, n10108_0, n10093_0, n10080_1/**/, n10011_0, n8400, n8392, n8384, n7412, n7404}), .out(n14379), .config_in(config_chain[34941:34936]), .config_rst(config_rst)); 
buffer_wire buffer_14379 (.in(n14379), .out(n14379_0));
mux3 mux_9214 (.in({n9865_0, n9864_0, n7412}), .out(n14380), .config_in(config_chain[34943:34942]), .config_rst(config_rst)); 
buffer_wire buffer_14380 (.in(n14380), .out(n14380_0));
mux15 mux_9215 (.in({n14473_1, n10425_0, n10406_0, n10391_0, n10377_0, n10370_0, n10363_0, n10356_0/**/, n10336_1, n10267_0, n8498, n8490, n8482, n7510, n7502}), .out(n14381), .config_in(config_chain[34949:34944]), .config_rst(config_rst)); 
buffer_wire buffer_14381 (.in(n14381), .out(n14381_0));
mux3 mux_9216 (.in({n9885_0, n9884_0, n7416}), .out(n14382), .config_in(config_chain[34951:34950]), .config_rst(config_rst)); 
buffer_wire buffer_14382 (.in(n14382), .out(n14382_0));
mux15 mux_9217 (.in({n14495_1, n10685_0, n10665_0, n10658_0, n10644_0/**/, n10629_0, n10615_0, n10608_0, n10594_1, n10525_0, n8596, n8588, n8580, n7608, n7600}), .out(n14383), .config_in(config_chain[34957:34952]), .config_rst(config_rst)); 
buffer_wire buffer_14383 (.in(n14383), .out(n14383_0));
mux3 mux_9218 (.in({n9907_0, n9826_1/**/, n7416}), .out(n14384), .config_in(config_chain[34959:34958]), .config_rst(config_rst)); 
buffer_wire buffer_14384 (.in(n14384), .out(n14384_0));
mux14 mux_9219 (.in({n14519_1, n10945_0, n10928_0, n10913_0, n10899_0, n10892_0, n10885_0, n10878_0, n10856_1, n8694, n8686, n8678, n7710/**/, n7698}), .out(n14385), .config_in(config_chain[34965:34960]), .config_rst(config_rst)); 
buffer_wire buffer_14385 (.in(n14385), .out(n14385_0));
mux3 mux_9220 (.in({n9847_0, n9846_0, n7416}), .out(n14386), .config_in(config_chain[34967:34966]), .config_rst(config_rst)); 
buffer_wire buffer_14386 (.in(n14386), .out(n14386_0));
mux14 mux_9221 (.in({n14453_1, n10165_0, n10149_0, n10142_0, n10128_0, n10113_0, n10101_0, n10094_0, n10082_1, n8400, n8392, n8384, n7416, n7404}), .out(n14387), .config_in(config_chain[34973:34968]), .config_rst(config_rst)); 
buffer_wire buffer_14387 (.in(n14387), .out(n14387_0));
mux3 mux_9222 (.in({n9867_0, n9866_0, n7416}), .out(n14388), .config_in(config_chain[34975:34974]), .config_rst(config_rst)); 
buffer_wire buffer_14388 (.in(n14388), .out(n14388_0));
mux14 mux_9223 (.in({n14475_1, n10423_0, n10399_0, n10392_0, n10385_0, n10378_0, n10364_0, n10349_0, n10338_1, n8498, n8490, n8482, n7514, n7502}), .out(n14389), .config_in(config_chain[34981:34976]), .config_rst(config_rst)); 
buffer_wire buffer_14389 (.in(n14389), .out(n14389_0));
mux3 mux_9224 (.in({n9887_0, n9886_0, n7416}), .out(n14390), .config_in(config_chain[34983:34982]), .config_rst(config_rst)); 
buffer_wire buffer_14390 (.in(n14390), .out(n14390_0));
mux14 mux_9225 (.in({n14497_1, n10683_0, n10666_0, n10651_0, n10637_0, n10630_0, n10623_0, n10616_0, n10596_1, n8596, n8588, n8580, n7612, n7600}), .out(n14391), .config_in(config_chain[34989:34984]), .config_rst(config_rst)); 
buffer_wire buffer_14391 (.in(n14391), .out(n14391_0));
mux3 mux_9226 (.in({n9909_0, n9828_1/**/, n7420}), .out(n14392), .config_in(config_chain[34991:34990]), .config_rst(config_rst)); 
buffer_wire buffer_14392 (.in(n14392), .out(n14392_0));
mux14 mux_9227 (.in({n14521_1, n10943_0, n10921_0, n10914_0/**/, n10907_0, n10900_0, n10886_0, n10871_0, n10858_1, n8694, n8686, n8678, n7710, n7702}), .out(n14393), .config_in(config_chain[34997:34992]), .config_rst(config_rst)); 
buffer_wire buffer_14393 (.in(n14393), .out(n14393_0));
mux3 mux_9228 (.in({n9849_0, n9848_0, n7420}), .out(n14394), .config_in(config_chain[34999:34998]), .config_rst(config_rst)); 
buffer_wire buffer_14394 (.in(n14394), .out(n14394_0));
mux14 mux_9229 (.in({n14455_1, n10163_0, n10150_0, n10135_0, n10121_0, n10114_0, n10109_0, n10102_0, n10084_1, n8400, n8392, n8384, n7416, n7408}), .out(n14395), .config_in(config_chain[35005:35000]), .config_rst(config_rst)); 
buffer_wire buffer_14395 (.in(n14395), .out(n14395_0));
mux3 mux_9230 (.in({n9869_0, n9868_0, n7420}), .out(n14396), .config_in(config_chain[35007:35006]), .config_rst(config_rst)); 
buffer_wire buffer_14396 (.in(n14396), .out(n14396_0));
mux14 mux_9231 (.in({n14477_1, n10421_0, n10407_0, n10400_0, n10386_0, n10371_0/**/, n10357_0, n10350_0, n10340_1, n8498, n8490, n8482, n7514, n7506}), .out(n14397), .config_in(config_chain[35013:35008]), .config_rst(config_rst)); 
buffer_wire buffer_14397 (.in(n14397), .out(n14397_0));
mux3 mux_9232 (.in({n9889_0, n9888_0, n7420}), .out(n14398), .config_in(config_chain[35015:35014]), .config_rst(config_rst)); 
buffer_wire buffer_14398 (.in(n14398), .out(n14398_0));
mux14 mux_9233 (.in({n14499_1, n10681_0, n10659_0/**/, n10652_0, n10645_0, n10638_0, n10624_0, n10609_0, n10598_1, n8596, n8588, n8580, n7612, n7604}), .out(n14399), .config_in(config_chain[35021:35016]), .config_rst(config_rst)); 
buffer_wire buffer_14399 (.in(n14399), .out(n14399_0));
mux3 mux_9234 (.in({n9911_0, n9830_1/**/, n7420}), .out(n14400), .config_in(config_chain[35023:35022]), .config_rst(config_rst)); 
buffer_wire buffer_14400 (.in(n14400), .out(n14400_0));
mux13 mux_9235 (.in({n14523_1, n10941_0, n10929_0, n10922_0, n10908_0, n10893_0, n10879_0, n10872_0, n10860_1, n8686, n8678, n7710, n7702}), .out(n14401), .config_in(config_chain[35029:35024]), .config_rst(config_rst)); 
buffer_wire buffer_14401 (.in(n14401), .out(n14401_0));
mux3 mux_9236 (.in({n9851_0, n9850_0, n8384}), .out(n14402), .config_in(config_chain[35031:35030]), .config_rst(config_rst)); 
buffer_wire buffer_14402 (.in(n14402), .out(n14402_0));
mux13 mux_9237 (.in({n14457_1, n10161_0, n10143_0, n10136_0, n10129_0, n10122_0, n10110_0, n10095_0, n10086_1, n8392, n8384, n7416, n7408}), .out(n14403), .config_in(config_chain[35037:35032]), .config_rst(config_rst)); 
buffer_wire buffer_14403 (.in(n14403), .out(n14403_0));
mux3 mux_9238 (.in({n9871_0, n9870_0, n8384}), .out(n14404), .config_in(config_chain[35039:35038]), .config_rst(config_rst)); 
buffer_wire buffer_14404 (.in(n14404), .out(n14404_0));
mux13 mux_9239 (.in({n14479_1, n10419_0, n10408_0, n10393_0, n10379_0, n10372_0, n10365_0, n10358_0, n10342_1, n8490, n8482, n7514, n7506}), .out(n14405), .config_in(config_chain[35045:35040]), .config_rst(config_rst)); 
buffer_wire buffer_14405 (.in(n14405), .out(n14405_0));
mux3 mux_9240 (.in({n9891_0, n9890_0, n8384}), .out(n14406), .config_in(config_chain[35047:35046]), .config_rst(config_rst)); 
buffer_wire buffer_14406 (.in(n14406), .out(n14406_0));
mux13 mux_9241 (.in({n14501_1, n10679_0, n10667_0, n10660_0/**/, n10646_0, n10631_0, n10617_0, n10610_0, n10600_1, n8588, n8580, n7612, n7604}), .out(n14407), .config_in(config_chain[35053:35048]), .config_rst(config_rst)); 
buffer_wire buffer_14407 (.in(n14407), .out(n14407_0));
mux3 mux_9242 (.in({n9913_0, n9832_1/**/, n8384}), .out(n14408), .config_in(config_chain[35055:35054]), .config_rst(config_rst)); 
buffer_wire buffer_14408 (.in(n14408), .out(n14408_0));
mux13 mux_9243 (.in({n14525_1, n10939_0, n10930_0, n10915_0, n10901_0, n10894_0, n10887_0, n10880_0, n10862_1/**/, n8690, n8678, n7710, n7702}), .out(n14409), .config_in(config_chain[35061:35056]), .config_rst(config_rst)); 
buffer_wire buffer_14409 (.in(n14409), .out(n14409_0));
mux3 mux_9244 (.in({n9853_0, n9852_0, n8384}), .out(n14410), .config_in(config_chain[35063:35062]), .config_rst(config_rst)); 
buffer_wire buffer_14410 (.in(n14410), .out(n14410_0));
mux13 mux_9245 (.in({n14459_1, n10159_0, n10151_0, n10144_0, n10130_0, n10115_0, n10103_0, n10096_0, n10088_1, n8396, n8384, n7416, n7408}), .out(n14411), .config_in(config_chain[35069:35064]), .config_rst(config_rst)); 
buffer_wire buffer_14411 (.in(n14411), .out(n14411_0));
mux3 mux_9246 (.in({n9873_0, n9872_0, n8388}), .out(n14412), .config_in(config_chain[35071:35070]), .config_rst(config_rst)); 
buffer_wire buffer_14412 (.in(n14412), .out(n14412_0));
mux13 mux_9247 (.in({n14481_1/**/, n10417_0, n10401_0, n10394_0, n10387_0, n10380_0, n10366_0, n10351_0, n10344_1, n8494, n8482, n7514, n7506}), .out(n14413), .config_in(config_chain[35077:35072]), .config_rst(config_rst)); 
buffer_wire buffer_14413 (.in(n14413), .out(n14413_0));
mux3 mux_9248 (.in({n9893_0, n9892_0, n8388}), .out(n14414), .config_in(config_chain[35079:35078]), .config_rst(config_rst)); 
buffer_wire buffer_14414 (.in(n14414), .out(n14414_0));
mux13 mux_9249 (.in({n14503_1, n10677_0, n10668_0, n10653_0, n10639_0, n10632_0, n10625_0, n10618_0, n10602_1, n8592, n8580, n7612/**/, n7604}), .out(n14415), .config_in(config_chain[35085:35080]), .config_rst(config_rst)); 
buffer_wire buffer_14415 (.in(n14415), .out(n14415_0));
mux3 mux_9250 (.in({n9915_0, n9834_1, n8388}), .out(n14416), .config_in(config_chain[35087:35086]), .config_rst(config_rst)); 
buffer_wire buffer_14416 (.in(n14416), .out(n14416_0));
mux13 mux_9251 (.in({n14527_1/**/, n10937_0, n10923_0, n10916_0, n10909_0, n10902_0, n10873_0, n10866_1, n10864_1, n8690, n8682, n7710, n7702}), .out(n14417), .config_in(config_chain[35093:35088]), .config_rst(config_rst)); 
buffer_wire buffer_14417 (.in(n14417), .out(n14417_0));
mux3 mux_9252 (.in({n9855_0, n9854_0, n8388}), .out(n14418), .config_in(config_chain[35095:35094]), .config_rst(config_rst)); 
buffer_wire buffer_14418 (.in(n14418), .out(n14418_0));
mux13 mux_9253 (.in({n14461_1, n10157_0, n10152_0, n10137_0, n10123_0, n10116_0, n10111_0, n10104_0, n10090_1/**/, n8396, n8388, n7416, n7408}), .out(n14419), .config_in(config_chain[35101:35096]), .config_rst(config_rst)); 
buffer_wire buffer_14419 (.in(n14419), .out(n14419_0));
mux3 mux_9254 (.in({n9875_0, n9874_0, n8388}), .out(n14420), .config_in(config_chain[35103:35102]), .config_rst(config_rst)); 
buffer_wire buffer_14420 (.in(n14420), .out(n14420_0));
mux13 mux_9255 (.in({n14483_1, n10415_0/**/, n10409_0, n10402_0, n10388_0, n10373_0, n10359_0, n10352_0, n10346_1, n8494, n8486, n7514, n7506}), .out(n14421), .config_in(config_chain[35109:35104]), .config_rst(config_rst)); 
buffer_wire buffer_14421 (.in(n14421), .out(n14421_0));
mux3 mux_9256 (.in({n9895_0, n9894_0, n8392}), .out(n14422), .config_in(config_chain[35111:35110]), .config_rst(config_rst)); 
buffer_wire buffer_14422 (.in(n14422), .out(n14422_0));
mux13 mux_9257 (.in({n14505_1, n10675_0, n10661_0, n10654_0, n10647_0, n10640_0, n10626_0, n10611_0, n10604_1, n8592, n8584, n7612, n7604}), .out(n14423), .config_in(config_chain[35117:35112]), .config_rst(config_rst)); 
buffer_wire buffer_14423 (.in(n14423), .out(n14423_0));
mux3 mux_9258 (.in({n9917_0, n9836_1/**/, n8392}), .out(n14424), .config_in(config_chain[35119:35118]), .config_rst(config_rst)); 
buffer_wire buffer_14424 (.in(n14424), .out(n14424_0));
mux13 mux_9259 (.in({n14529_1, n10935_0, n10931_0, n10924_0, n10895_0, n10888_0, n10881_0, n10874_0, n10782_2, n8690, n8682, n7714/**/, n7702}), .out(n14425), .config_in(config_chain[35125:35120]), .config_rst(config_rst)); 
buffer_wire buffer_14425 (.in(n14425), .out(n14425_0));
mux3 mux_9260 (.in({n9857_0, n9856_0, n8392}), .out(n14426), .config_in(config_chain[35127:35126]), .config_rst(config_rst)); 
buffer_wire buffer_14426 (.in(n14426), .out(n14426_0));
mux13 mux_9261 (.in({n14463_1, n10155_0, n10145_0, n10138_0, n10131_0, n10124_0, n10097_0, n10004_2, n10002_2, n8396, n8388, n7420, n7408}), .out(n14427), .config_in(config_chain[35133:35128]), .config_rst(config_rst)); 
buffer_wire buffer_14427 (.in(n14427), .out(n14427_0));
mux3 mux_9262 (.in({n9877_0, n9876_0, n8392}), .out(n14428), .config_in(config_chain[35135:35134]), .config_rst(config_rst)); 
buffer_wire buffer_14428 (.in(n14428), .out(n14428_0));
mux13 mux_9263 (.in({n14485_1, n10413_0, n10410_0, n10395_0, n10381_0, n10374_0, n10367_0, n10360_0, n10260_2, n8494, n8486, n7518, n7506/**/}), .out(n14429), .config_in(config_chain[35141:35136]), .config_rst(config_rst)); 
buffer_wire buffer_14429 (.in(n14429), .out(n14429_0));
mux3 mux_9264 (.in({n9897_0, n9896_0, n8392}), .out(n14430), .config_in(config_chain[35143:35142]), .config_rst(config_rst)); 
buffer_wire buffer_14430 (.in(n14430), .out(n14430_0));
mux13 mux_9265 (.in({n14507_1, n10673_0, n10669_0, n10662_0, n10648_0, n10633_0, n10619_0, n10612_0, n10520_2, n8592, n8584, n7616, n7604}), .out(n14431), .config_in(config_chain[35149:35144]), .config_rst(config_rst)); 
buffer_wire buffer_14431 (.in(n14431), .out(n14431_0));
mux3 mux_9266 (.in({n9919_0/**/, n9746_2, n8396}), .out(n14432), .config_in(config_chain[35151:35150]), .config_rst(config_rst)); 
buffer_wire buffer_14432 (.in(n14432), .out(n14432_0));
mux3 mux_9267 (.in({n12091_0, n12090_2, n9180}), .out(n14433), .config_in(config_chain[35153:35152]), .config_rst(config_rst)); 
buffer_wire buffer_14433 (.in(n14433), .out(n14433_0));
mux3 mux_9268 (.in({n9749_0, n9748_2, n8396}), .out(n14434), .config_in(config_chain[35155:35154]), .config_rst(config_rst)); 
buffer_wire buffer_14434 (.in(n14434), .out(n14434_0));
mux13 mux_9269 (.in({n14465_2, n10175_0, n10153_0, n10146_0, n10117_0, n10105_0, n10098_0, n10072_1, n10006_2, n8396, n8388, n7420, n7412}), .out(n14435), .config_in(config_chain[35161:35156]), .config_rst(config_rst)); 
buffer_wire buffer_14435 (.in(n14435), .out(n14435_0));
mux3 mux_9270 (.in({n9751_0, n9750_2, n8396}), .out(n14436), .config_in(config_chain[35163:35162]), .config_rst(config_rst)); 
buffer_wire buffer_14436 (.in(n14436), .out(n14436_0));
mux13 mux_9271 (.in({n14487_2, n10433_0, n10403_0, n10396_0, n10389_0, n10382_0, n10353_0, n10328_1, n10262_2, n8494, n8486, n7518, n7510}), .out(n14437), .config_in(config_chain[35169:35164]), .config_rst(config_rst)); 
buffer_wire buffer_14437 (.in(n14437), .out(n14437_0));
mux3 mux_9272 (.in({n9753_0, n9752_2, n8396}), .out(n14438), .config_in(config_chain[35171:35170]), .config_rst(config_rst)); 
buffer_wire buffer_14438 (.in(n14438), .out(n14438_0));
mux13 mux_9273 (.in({n14509_1, n10693_0, n10670_0, n10655_0, n10641_0, n10634_0, n10627_0, n10620_0, n10586_1, n8592, n8584, n7616, n7608}), .out(n14439), .config_in(config_chain[35177:35172]), .config_rst(config_rst)); 
buffer_wire buffer_14439 (.in(n14439), .out(n14439_0));
mux3 mux_9274 (.in({n9755_0, n9754_2, n8396}), .out(n14440), .config_in(config_chain[35179:35178]), .config_rst(config_rst)); 
buffer_wire buffer_14440 (.in(n14440), .out(n14440_0));
mux13 mux_9275 (.in({n14531_1/**/, n10955_0, n10917_0, n10910_0, n10903_0, n10896_0, n10882_0, n10867_0, n10846_1, n8690, n8682, n7714, n7706}), .out(n14441), .config_in(config_chain[35185:35180]), .config_rst(config_rst)); 
buffer_wire buffer_14441 (.in(n14441), .out(n14441_0));
mux3 mux_9276 (.in({n9757_0, n9756_2, n8400}), .out(n14442), .config_in(config_chain[35187:35186]), .config_rst(config_rst)); 
buffer_wire buffer_14442 (.in(n14442), .out(n14442_0));
mux13 mux_9277 (.in({n14553_1, n11219_0, n11190_0, n11159_0, n11152_0, n11145_0, n11138_0, n11110_1/**/, n11109_0, n8788, n8780, n7812, n7804}), .out(n14443), .config_in(config_chain[35193:35188]), .config_rst(config_rst)); 
buffer_wire buffer_14443 (.in(n14443), .out(n14443_0));
mux15 mux_9278 (.in({n14354_0, n10157_0, n10138_0, n10133_0, n10124_0, n10119_0, n10107_0, n10072_1/**/, n10009_0, n10004_2, n8494, n8486, n7518, n7510, n7502}), .out(n14444), .config_in(config_chain[35199:35194]), .config_rst(config_rst)); 
buffer_wire buffer_14444 (.in(n14444), .out(n14444_0));
mux15 mux_9279 (.in({n14533_1, n11217_0, n11183_0, n11176_0, n11174_0, n11167_0, n11160_0, n11146_0, n11131_0, n11112_1/**/, n8788, n8780, n7812, n7804, n7796}), .out(n14445), .config_in(config_chain[35205:35200]), .config_rst(config_rst)); 
buffer_wire buffer_14445 (.in(n14445), .out(n14445_0));
mux15 mux_9280 (.in({n14362_0, n10159_0, n10146_0, n10141_0, n10127_0, n10098_0/**/, n10093_0, n10011_0, n10006_2, n10002_2, n8498, n8486, n7518, n7510, n7502}), .out(n14446), .config_in(config_chain[35211:35206]), .config_rst(config_rst)); 
buffer_wire buffer_14446 (.in(n14446), .out(n14446_0));
mux15 mux_9281 (.in({n14535_1, n11215_0, n11196_0, n11191_0, n11184_0, n11168_0/**/, n11153_0, n11139_0, n11132_0, n11114_1, n8792, n8780, n7812, n7804, n7796}), .out(n14447), .config_in(config_chain[35217:35212]), .config_rst(config_rst)); 
buffer_wire buffer_14447 (.in(n14447), .out(n14447_0));
mux15 mux_9282 (.in({n14370_0, n10161_0, n10149_0, n10132_0, n10118_0, n10113_0, n10106_0/**/, n10101_0, n10090_1, n10008_2, n8498, n8490, n7518, n7510, n7502}), .out(n14448), .config_in(config_chain[35223:35218]), .config_rst(config_rst)); 
buffer_wire buffer_14448 (.in(n14448), .out(n14448_0));
mux15 mux_9283 (.in({n14537_1/**/, n11213_0, n11192_0, n11177_0, n11175_0, n11161_0, n11154_0, n11147_0, n11140_0, n11116_1, n8792, n8784, n7812, n7804, n7796}), .out(n14449), .config_in(config_chain[35229:35224]), .config_rst(config_rst)); 
buffer_wire buffer_14449 (.in(n14449), .out(n14449_0));
mux15 mux_9284 (.in({n14378_0, n10163_0, n10140_0/**/, n10135_0, n10126_0, n10121_0, n10109_0, n10092_0, n10088_1, n10010_2, n8498, n8490, n8482, n7510, n7502}), .out(n14450), .config_in(config_chain[35235:35230]), .config_rst(config_rst)); 
buffer_wire buffer_14450 (.in(n14450), .out(n14450_0));
mux15 mux_9285 (.in({n14539_1, n11211_0, n11197_0, n11185_0, n11178_0, n11169_0, n11162_0, n11148_0, n11133_0, n11118_1, n8792/**/, n8784, n8776, n7804, n7796}), .out(n14451), .config_in(config_chain[35241:35236]), .config_rst(config_rst)); 
buffer_wire buffer_14451 (.in(n14451), .out(n14451_0));
mux14 mux_9286 (.in({n14386_0, n10165_0, n10148_0, n10143_0, n10129_0, n10112_0, n10100_0, n10095_0, n10086_1, n8498, n8490, n8482, n7514, n7502}), .out(n14452), .config_in(config_chain[35247:35242]), .config_rst(config_rst)); 
buffer_wire buffer_14452 (.in(n14452), .out(n14452_0));
mux14 mux_9287 (.in({n14541_1/**/, n11209_0, n11193_0, n11186_0, n11170_0, n11155_0, n11141_0, n11134_0, n11120_1, n8792, n8784, n8776, n7808, n7796}), .out(n14453), .config_in(config_chain[35253:35248]), .config_rst(config_rst)); 
buffer_wire buffer_14453 (.in(n14453), .out(n14453_0));
mux14 mux_9288 (.in({n14394_0, n10167_0, n10151_0, n10134_0, n10120_0, n10115_0, n10108_0, n10103_0/**/, n10084_1, n8498, n8490, n8482, n7514, n7506}), .out(n14454), .config_in(config_chain[35259:35254]), .config_rst(config_rst)); 
buffer_wire buffer_14454 (.in(n14454), .out(n14454_0));
mux14 mux_9289 (.in({n14543_1, n11207_0/**/, n11194_0, n11179_0, n11163_0, n11156_0, n11149_0, n11142_0, n11122_1, n8792, n8784, n8776, n7808, n7800}), .out(n14455), .config_in(config_chain[35265:35260]), .config_rst(config_rst)); 
buffer_wire buffer_14455 (.in(n14455), .out(n14455_0));
mux13 mux_9290 (.in({n14402_0, n10169_0, n10142_0, n10137_0, n10128_0, n10123_0, n10111_0, n10094_0, n10082_1/**/, n8490, n8482, n7514, n7506}), .out(n14456), .config_in(config_chain[35271:35266]), .config_rst(config_rst)); 
buffer_wire buffer_14456 (.in(n14456), .out(n14456_0));
mux13 mux_9291 (.in({n14545_1, n11205_0, n11187_0, n11180_0, n11171_0, n11164_0, n11150_0, n11135_0/**/, n11124_1, n8784, n8776, n7808, n7800}), .out(n14457), .config_in(config_chain[35277:35272]), .config_rst(config_rst)); 
buffer_wire buffer_14457 (.in(n14457), .out(n14457_0));
mux13 mux_9292 (.in({n14410_0, n10171_0, n10150_0/**/, n10145_0, n10131_0, n10114_0, n10102_0, n10097_0, n10080_1, n8494, n8482, n7514, n7506}), .out(n14458), .config_in(config_chain[35283:35278]), .config_rst(config_rst)); 
buffer_wire buffer_14458 (.in(n14458), .out(n14458_0));
mux13 mux_9293 (.in({n14547_1, n11203_0, n11195_0, n11188_0, n11172_0/**/, n11157_0, n11143_0, n11136_0, n11126_1, n8788, n8776, n7808, n7800}), .out(n14459), .config_in(config_chain[35289:35284]), .config_rst(config_rst)); 
buffer_wire buffer_14459 (.in(n14459), .out(n14459_0));
mux13 mux_9294 (.in({n14418_0, n10173_0, n10153_0, n10136_0/**/, n10122_0, n10117_0, n10110_0, n10105_0, n10078_1, n8494, n8486, n7514, n7506}), .out(n14460), .config_in(config_chain[35295:35290]), .config_rst(config_rst)); 
buffer_wire buffer_14460 (.in(n14460), .out(n14460_0));
mux13 mux_9295 (.in({n14549_1, n11201_0, n11181_0, n11165_0, n11158_0/**/, n11151_0, n11144_0, n11128_1, n11108_1, n8788, n8780, n7808, n7800}), .out(n14461), .config_in(config_chain[35301:35296]), .config_rst(config_rst)); 
buffer_wire buffer_14461 (.in(n14461), .out(n14461_0));
mux13 mux_9296 (.in({n14426_0, n10175_0, n10144_0, n10139_0, n10130_0, n10125_0, n10096_0/**/, n10076_1, n10005_0, n8494, n8486, n7518, n7506}), .out(n14462), .config_in(config_chain[35307:35302]), .config_rst(config_rst)); 
buffer_wire buffer_14462 (.in(n14462), .out(n14462_0));
mux13 mux_9297 (.in({n14551_1, n11199_0, n11189_0/**/, n11182_0, n11173_0, n11166_0, n11137_0, n11130_1, n11046_2, n8788, n8780, n7812, n7800}), .out(n14463), .config_in(config_chain[35313:35308]), .config_rst(config_rst)); 
buffer_wire buffer_14463 (.in(n14463), .out(n14463_0));
mux13 mux_9298 (.in({n14434_0, n10155_0, n10152_0, n10147_0, n10116_0/**/, n10104_0, n10099_0, n10074_1, n10007_0, n8494, n8486, n7518, n7510}), .out(n14464), .config_in(config_chain[35319:35314]), .config_rst(config_rst)); 
buffer_wire buffer_14464 (.in(n14464), .out(n14464_0));
mux3 mux_9299 (.in({n12093_0, n12092_2, n9180}), .out(n14465), .config_in(config_chain[35321:35320]), .config_rst(config_rst)); 
buffer_wire buffer_14465 (.in(n14465), .out(n14465_0));
mux15 mux_9300 (.in({n14356_0, n10415_0, n10410_0, n10405_0, n10374_0, n10369_0, n10360_0, n10355_0, n10328_1, n10265_0, n8592, n8584, n7616, n7608, n7600}), .out(n14466), .config_in(config_chain[35327:35322]), .config_rst(config_rst)); 
buffer_wire buffer_14466 (.in(n14466), .out(n14466_0));
mux16 mux_9301 (.in({n14555_0, n11481_0, n11448_0/**/, n11445_0, n11441_0, n11437_0, n11420_0, n11410_0, n11407_0, n11378_1, n11352_1, n8886, n8878, n7910, n7902, n7894}), .out(n14467), .config_in(config_chain[35333:35328]), .config_rst(config_rst)); 
buffer_wire buffer_14467 (.in(n14467), .out(n14467_0));
mux15 mux_9302 (.in({n14364_0, n10417_0, n10396_0, n10391_0/**/, n10382_0, n10377_0, n10363_0, n10267_0, n10262_2, n10260_2, n8596, n8584, n7616, n7608, n7600}), .out(n14468), .config_in(config_chain[35339:35334]), .config_rst(config_rst)); 
buffer_wire buffer_14468 (.in(n14468), .out(n14468_0));
mux16 mux_9303 (.in({n14557_0, n11479_0, n11463_0, n11459_0, n11442_0, n11434_0, n11431_0, n11404_0, n11401_0, n11380_1, n11374_1/**/, n8886, n8878, n7910, n7902, n7894}), .out(n14469), .config_in(config_chain[35345:35340]), .config_rst(config_rst)); 
buffer_wire buffer_14469 (.in(n14469), .out(n14469_0));
mux15 mux_9304 (.in({n14372_0, n10419_0, n10404_0, n10399_0, n10385_0, n10368_0, n10354_0, n10349_0, n10346_1/**/, n10264_2, n8596, n8588, n7616, n7608, n7600}), .out(n14470), .config_in(config_chain[35351:35346]), .config_rst(config_rst)); 
buffer_wire buffer_14470 (.in(n14470), .out(n14470_0));
mux15 mux_9305 (.in({n14559_0, n11477_0, n11456_0, n11453_0, n11428_0, n11425_0, n11415_0, n11398_0, n11396_1, n11382_1, n8886, n8878, n7910, n7902, n7894}), .out(n14471), .config_in(config_chain[35357:35352]), .config_rst(config_rst)); 
buffer_wire buffer_14471 (.in(n14471), .out(n14471_0));
mux15 mux_9306 (.in({n14380_0, n10421_0, n10407_0, n10390_0, n10376_0, n10371_0, n10362_0, n10357_0, n10344_1, n10266_2, n8596/**/, n8588, n8580, n7608, n7600}), .out(n14472), .config_in(config_chain[35363:35358]), .config_rst(config_rst)); 
buffer_wire buffer_14472 (.in(n14472), .out(n14472_0));
mux15 mux_9307 (.in({n14561_0, n11475_0, n11450_0, n11447_0, n11439_0, n11422_0, n11418_0, n11412_0, n11409_0, n11384_1, n8886/**/, n8878, n7910, n7902, n7894}), .out(n14473), .config_in(config_chain[35369:35364]), .config_rst(config_rst)); 
buffer_wire buffer_14473 (.in(n14473), .out(n14473_0));
mux14 mux_9308 (.in({n14388_0, n10423_0, n10398_0/**/, n10393_0, n10384_0, n10379_0, n10365_0, n10348_0, n10342_1, n8596, n8588, n8580, n7612, n7600}), .out(n14474), .config_in(config_chain[35375:35370]), .config_rst(config_rst)); 
buffer_wire buffer_14474 (.in(n14474), .out(n14474_0));
mux15 mux_9309 (.in({n14563_0, n11473_0, n11461_0, n11444_0, n11440_0, n11436_0/**/, n11433_0, n11406_0, n11403_0, n11386_1, n8886, n8878, n7910, n7902, n7894}), .out(n14475), .config_in(config_chain[35381:35376]), .config_rst(config_rst)); 
buffer_wire buffer_14475 (.in(n14475), .out(n14475_0));
mux14 mux_9310 (.in({n14396_0, n10425_0/**/, n10406_0, n10401_0, n10387_0, n10370_0, n10356_0, n10351_0, n10340_1, n8596, n8588, n8580, n7612, n7604}), .out(n14476), .config_in(config_chain[35387:35382]), .config_rst(config_rst)); 
buffer_wire buffer_14476 (.in(n14476), .out(n14476_0));
mux15 mux_9311 (.in({n14565_0, n11471_0, n11462_0, n11458_0, n11455_0, n11430_0, n11427_0, n11417_0, n11400_0, n11388_1, n8890, n8882, n8874, n7906, n7898}), .out(n14477), .config_in(config_chain[35393:35388]), .config_rst(config_rst)); 
buffer_wire buffer_14477 (.in(n14477), .out(n14477_0));
mux13 mux_9312 (.in({n14404_0, n10427_0, n10409_0, n10392_0/**/, n10378_0, n10373_0, n10364_0, n10359_0, n10338_1, n8588, n8580, n7612, n7604}), .out(n14478), .config_in(config_chain[35399:35394]), .config_rst(config_rst)); 
buffer_wire buffer_14478 (.in(n14478), .out(n14478_0));
mux15 mux_9313 (.in({n14567_0/**/, n11469_0, n11452_0, n11449_0, n11424_0, n11421_0, n11414_0, n11411_0, n11390_1, n11353_0, n8890, n8882, n8874, n7906, n7898}), .out(n14479), .config_in(config_chain[35405:35400]), .config_rst(config_rst)); 
buffer_wire buffer_14479 (.in(n14479), .out(n14479_0));
mux13 mux_9314 (.in({n14412_0, n10429_0, n10400_0, n10395_0, n10386_0, n10381_0, n10367_0, n10350_0, n10336_1/**/, n8592, n8580, n7612, n7604}), .out(n14480), .config_in(config_chain[35411:35406]), .config_rst(config_rst)); 
buffer_wire buffer_14480 (.in(n14480), .out(n14480_0));
mux15 mux_9315 (.in({n14569_0, n11467_0, n11446_0, n11443_0, n11438_0, n11435_0, n11408_0, n11405_0, n11392_1/**/, n11375_0, n8890, n8882, n8874, n7906, n7898}), .out(n14481), .config_in(config_chain[35417:35412]), .config_rst(config_rst)); 
buffer_wire buffer_14481 (.in(n14481), .out(n14481_0));
mux13 mux_9316 (.in({n14420_0, n10431_0, n10408_0, n10403_0, n10389_0, n10372_0, n10358_0, n10353_0, n10334_1, n8592, n8584, n7612/**/, n7604}), .out(n14482), .config_in(config_chain[35423:35418]), .config_rst(config_rst)); 
buffer_wire buffer_14482 (.in(n14482), .out(n14482_0));
mux15 mux_9317 (.in({n14571_0, n11465_0, n11460_0, n11457_0, n11432_0/**/, n11429_0, n11402_0, n11399_0, n11397_0, n11394_1, n8890, n8882, n8874, n7906, n7898}), .out(n14483), .config_in(config_chain[35429:35424]), .config_rst(config_rst)); 
buffer_wire buffer_14483 (.in(n14483), .out(n14483_0));
mux13 mux_9318 (.in({n14428_0, n10433_0, n10411_0, n10394_0, n10380_0/**/, n10375_0, n10366_0, n10361_0, n10332_1, n8592, n8584, n7616, n7604}), .out(n14484), .config_in(config_chain[35435:35430]), .config_rst(config_rst)); 
buffer_wire buffer_14484 (.in(n14484), .out(n14484_0));
mux15 mux_9319 (.in({n14573_0, n11483_0, n11454_0, n11451_0, n11426_0, n11423_0, n11419_0, n11416_0/**/, n11413_0, n11376_1, n8890, n8882, n8874, n7906, n7898}), .out(n14485), .config_in(config_chain[35441:35436]), .config_rst(config_rst)); 
buffer_wire buffer_14485 (.in(n14485), .out(n14485_0));
mux13 mux_9320 (.in({n14436_0, n10413_0/**/, n10402_0, n10397_0, n10388_0, n10383_0, n10352_0, n10330_1, n10263_0, n8592, n8584, n7616, n7608}), .out(n14486), .config_in(config_chain[35447:35442]), .config_rst(config_rst)); 
buffer_wire buffer_14486 (.in(n14486), .out(n14486_0));
mux3 mux_9321 (.in({n12123_0, n12122_2, n9180}), .out(n14487), .config_in(config_chain[35449:35448]), .config_rst(config_rst)); 
buffer_wire buffer_14487 (.in(n14487), .out(n14487_0));
mux15 mux_9322 (.in({n14358_0, n10675_0, n10662_0, n10657_0, n10648_0/**/, n10643_0, n10612_0, n10607_0, n10586_1, n10523_0, n8690, n8682, n7714, n7706, n7698}), .out(n14488), .config_in(config_chain[35455:35450]), .config_rst(config_rst)); 
buffer_wire buffer_14488 (.in(n14488), .out(n14488_0));
mux16 mux_9323 (.in({n14575_0, n11745_0, n11720_0, n11717_0, n11692_0, n11689_0, n11685_0, n11681_0, n11664_0, n11644_1, n11596_2, n8984, n8976, n8008, n8000, n7992}), .out(n14489), .config_in(config_chain[35461:35456]), .config_rst(config_rst)); 
buffer_wire buffer_14489 (.in(n14489), .out(n14489_0));
mux15 mux_9324 (.in({n14366_0, n10677_0, n10670_0/**/, n10665_0, n10634_0, n10629_0, n10620_0, n10615_0, n10525_0, n10520_2, n8694, n8682, n7714, n7706, n7698}), .out(n14490), .config_in(config_chain[35467:35462]), .config_rst(config_rst)); 
buffer_wire buffer_14490 (.in(n14490), .out(n14490_0));
mux16 mux_9325 (.in({n14577_0, n11743_0, n11714_0/**/, n11711_0, n11707_0, n11703_0, n11686_0, n11678_0, n11675_0, n11646_1, n11618_1, n8984, n8976, n8008, n8000, n7992}), .out(n14491), .config_in(config_chain[35473:35468]), .config_rst(config_rst)); 
buffer_wire buffer_14491 (.in(n14491), .out(n14491_0));
mux15 mux_9326 (.in({n14374_0, n10679_0, n10656_0, n10651_0, n10642_0, n10637_0, n10623_0, n10606_0, n10604_1, n10522_2, n8694/**/, n8686, n7714, n7706, n7698}), .out(n14492), .config_in(config_chain[35479:35474]), .config_rst(config_rst)); 
buffer_wire buffer_14492 (.in(n14492), .out(n14492_0));
mux15 mux_9327 (.in({n14579_0/**/, n11741_0, n11725_0, n11708_0, n11700_0, n11697_0, n11672_0, n11669_0, n11648_1, n11640_1, n8984, n8976, n8008, n8000, n7992}), .out(n14493), .config_in(config_chain[35485:35480]), .config_rst(config_rst)); 
buffer_wire buffer_14493 (.in(n14493), .out(n14493_0));
mux15 mux_9328 (.in({n14382_0, n10681_0, n10664_0, n10659_0, n10645_0, n10628_0, n10614_0, n10609_0, n10602_1, n10524_2, n8694, n8686, n8678/**/, n7706, n7698}), .out(n14494), .config_in(config_chain[35491:35486]), .config_rst(config_rst)); 
buffer_wire buffer_14494 (.in(n14494), .out(n14494_0));
mux15 mux_9329 (.in({n14581_0, n11739_0, n11722_0, n11719_0, n11694_0/**/, n11691_0, n11683_0, n11666_0, n11662_1, n11650_1, n8984, n8976, n8008, n8000, n7992}), .out(n14495), .config_in(config_chain[35497:35492]), .config_rst(config_rst)); 
buffer_wire buffer_14495 (.in(n14495), .out(n14495_0));
mux14 mux_9330 (.in({n14390_0, n10683_0, n10667_0, n10650_0/**/, n10636_0, n10631_0, n10622_0, n10617_0, n10600_1, n8694, n8686, n8678, n7710, n7698}), .out(n14496), .config_in(config_chain[35503:35498]), .config_rst(config_rst)); 
buffer_wire buffer_14496 (.in(n14496), .out(n14496_0));
mux15 mux_9331 (.in({n14583_0, n11737_0, n11716_0, n11713_0, n11705_0, n11688_0, n11684_0, n11680_0, n11677_0, n11652_1/**/, n8984, n8976, n8008, n8000, n7992}), .out(n14497), .config_in(config_chain[35509:35504]), .config_rst(config_rst)); 
buffer_wire buffer_14497 (.in(n14497), .out(n14497_0));
mux14 mux_9332 (.in({n14398_0, n10685_0, n10658_0, n10653_0, n10644_0, n10639_0, n10625_0, n10608_0, n10598_1, n8694, n8686, n8678, n7710, n7702}), .out(n14498), .config_in(config_chain[35515:35510]), .config_rst(config_rst)); 
buffer_wire buffer_14498 (.in(n14498), .out(n14498_0));
mux15 mux_9333 (.in({n14585_0, n11735_0, n11727_0, n11710_0, n11706_0, n11702_0, n11699_0/**/, n11674_0, n11671_0, n11654_1, n8988, n8980, n8972, n8004, n7996}), .out(n14499), .config_in(config_chain[35521:35516]), .config_rst(config_rst)); 
buffer_wire buffer_14499 (.in(n14499), .out(n14499_0));
mux13 mux_9334 (.in({n14406_0, n10687_0, n10666_0, n10661_0, n10647_0, n10630_0, n10616_0, n10611_0, n10596_1, n8686/**/, n8678, n7710, n7702}), .out(n14500), .config_in(config_chain[35527:35522]), .config_rst(config_rst)); 
buffer_wire buffer_14500 (.in(n14500), .out(n14500_0));
mux15 mux_9335 (.in({n14587_0, n11733_0, n11724_0, n11721_0, n11696_0, n11693_0, n11668_0, n11665_0, n11656_1, n11597_0, n8988, n8980/**/, n8972, n8004, n7996}), .out(n14501), .config_in(config_chain[35533:35528]), .config_rst(config_rst)); 
buffer_wire buffer_14501 (.in(n14501), .out(n14501_0));
mux13 mux_9336 (.in({n14414_0, n10689_0, n10669_0, n10652_0, n10638_0, n10633_0, n10624_0, n10619_0, n10594_1, n8690, n8678, n7710, n7702}), .out(n14502), .config_in(config_chain[35539:35534]), .config_rst(config_rst)); 
buffer_wire buffer_14502 (.in(n14502), .out(n14502_0));
mux15 mux_9337 (.in({n14589_0, n11731_0, n11718_0, n11715_0, n11690_0, n11687_0, n11682_0, n11679_0, n11658_1/**/, n11619_0, n8988, n8980, n8972, n8004, n7996}), .out(n14503), .config_in(config_chain[35545:35540]), .config_rst(config_rst)); 
buffer_wire buffer_14503 (.in(n14503), .out(n14503_0));
mux13 mux_9338 (.in({n14422_0, n10691_0/**/, n10660_0, n10655_0, n10646_0, n10641_0, n10627_0, n10610_0, n10592_1, n8690, n8682, n7710, n7702}), .out(n14504), .config_in(config_chain[35551:35546]), .config_rst(config_rst)); 
buffer_wire buffer_14504 (.in(n14504), .out(n14504_0));
mux15 mux_9339 (.in({n14591_0, n11729_0, n11712_0, n11709_0, n11704_0, n11701_0, n11676_0, n11673_0, n11660_1, n11641_0, n8988/**/, n8980, n8972, n8004, n7996}), .out(n14505), .config_in(config_chain[35557:35552]), .config_rst(config_rst)); 
buffer_wire buffer_14505 (.in(n14505), .out(n14505_0));
mux13 mux_9340 (.in({n14430_0, n10693_0, n10668_0/**/, n10663_0, n10649_0, n10632_0, n10618_0, n10613_0, n10590_1, n8690, n8682, n7714, n7702}), .out(n14506), .config_in(config_chain[35563:35558]), .config_rst(config_rst)); 
buffer_wire buffer_14506 (.in(n14506), .out(n14506_0));
mux15 mux_9341 (.in({n14593_0, n11747_0, n11726_0, n11723_0, n11698_0/**/, n11695_0, n11670_0, n11667_0, n11663_0, n11642_1, n8988, n8980, n8972, n8004, n7996}), .out(n14507), .config_in(config_chain[35569:35564]), .config_rst(config_rst)); 
buffer_wire buffer_14507 (.in(n14507), .out(n14507_0));
mux13 mux_9342 (.in({n14438_0, n10673_0, n10671_0, n10654_0, n10640_0, n10635_0, n10626_0, n10621_0, n10588_1/**/, n8690, n8682, n7714, n7706}), .out(n14508), .config_in(config_chain[35575:35570]), .config_rst(config_rst)); 
buffer_wire buffer_14508 (.in(n14508), .out(n14508_0));
mux3 mux_9343 (.in({n12145_0, n12144_1/**/, n9180}), .out(n14509), .config_in(config_chain[35577:35576]), .config_rst(config_rst)); 
buffer_wire buffer_14509 (.in(n14509), .out(n14509_0));
mux15 mux_9344 (.in({n14352_1, n10937_0, n10933_0, n10924_0, n10919_0, n10905_0, n10888_0, n10874_0, n10869_0, n10846_1, n8788, n8780, n7812, n7804, n7796}), .out(n14510), .config_in(config_chain[35583:35578]), .config_rst(config_rst)); 
buffer_wire buffer_14510 (.in(n14510), .out(n14510_0));
mux16 mux_9345 (.in({n14595_0, n12007_0, n11982_0, n11979_0, n11956_0, n11953_0, n11945_0, n11928_0, n11927_0, n11908_1, n11828_2, n9082, n9074, n8106, n8098, n8090}), .out(n14511), .config_in(config_chain[35589:35584]), .config_rst(config_rst)); 
buffer_wire buffer_14511 (.in(n14511), .out(n14511_0));
mux15 mux_9346 (.in({n14360_1/**/, n10939_0, n10927_0, n10910_0, n10896_0, n10891_0, n10882_0, n10877_0, n10785_0, n10782_2, n8792, n8780, n7812, n7804, n7796}), .out(n14512), .config_in(config_chain[35595:35590]), .config_rst(config_rst)); 
buffer_wire buffer_14512 (.in(n14512), .out(n14512_0));
mux16 mux_9347 (.in({n14597_0, n12005_0, n11976_0, n11973_0, n11967_0, n11950_0, n11949_0, n11942_0, n11939_0, n11910_1, n11860_2, n9082, n9074, n8106, n8098, n8090/**/}), .out(n14513), .config_in(config_chain[35601:35596]), .config_rst(config_rst)); 
buffer_wire buffer_14513 (.in(n14513), .out(n14513_0));
mux15 mux_9348 (.in({n14368_1, n10941_0, n10932_0, n10918_0, n10913_0, n10904_0, n10899_0, n10885_0, n10868_0/**/, n10864_1, n8792, n8784, n7812, n7804, n7796}), .out(n14514), .config_in(config_chain[35607:35602]), .config_rst(config_rst)); 
buffer_wire buffer_14514 (.in(n14514), .out(n14514_0));
mux15 mux_9349 (.in({n14599_0, n12003_0, n11987_0, n11970_0, n11964_0, n11961_0, n11936_0, n11933_0, n11912_1, n11882_1, n9082/**/, n9074, n8106, n8098, n8090}), .out(n14515), .config_in(config_chain[35613:35608]), .config_rst(config_rst)); 
buffer_wire buffer_14515 (.in(n14515), .out(n14515_0));
mux15 mux_9350 (.in({n14376_1, n10943_0, n10926_0, n10921_0, n10907_0/**/, n10890_0, n10876_0, n10871_0, n10862_1, n10784_2, n8792, n8784, n8776, n7804, n7796}), .out(n14516), .config_in(config_chain[35619:35614]), .config_rst(config_rst)); 
buffer_wire buffer_14516 (.in(n14516), .out(n14516_0));
mux15 mux_9351 (.in({n14601_0, n12001_0, n11984_0, n11981_0, n11958_0, n11955_0, n11947_0, n11930_0, n11914_1, n11904_1, n9082/**/, n9074, n8106, n8098, n8090}), .out(n14517), .config_in(config_chain[35625:35620]), .config_rst(config_rst)); 
buffer_wire buffer_14517 (.in(n14517), .out(n14517_0));
mux14 mux_9352 (.in({n14384_1, n10945_0, n10929_0, n10912_0/**/, n10898_0, n10893_0, n10884_0, n10879_0, n10860_1, n8792, n8784, n8776, n7808, n7796}), .out(n14518), .config_in(config_chain[35631:35626]), .config_rst(config_rst)); 
buffer_wire buffer_14518 (.in(n14518), .out(n14518_0));
mux15 mux_9353 (.in({n14603_0, n11999_0/**/, n11978_0, n11975_0, n11969_0, n11952_0, n11944_0, n11941_0, n11926_1, n11916_1, n9082, n9074, n8106, n8098, n8090}), .out(n14519), .config_in(config_chain[35637:35632]), .config_rst(config_rst)); 
buffer_wire buffer_14519 (.in(n14519), .out(n14519_0));
mux14 mux_9354 (.in({n14392_1, n10947_0, n10920_0, n10915_0, n10906_0, n10901_0, n10887_0, n10870_0, n10858_1, n8792, n8784/**/, n8776, n7808, n7800}), .out(n14520), .config_in(config_chain[35643:35638]), .config_rst(config_rst)); 
buffer_wire buffer_14520 (.in(n14520), .out(n14520_0));
mux15 mux_9355 (.in({n14605_0, n11997_0, n11989_0, n11972_0, n11966_0, n11963_0, n11948_0, n11938_0, n11935_0, n11918_1, n9086/**/, n9078, n9070, n8102, n8094}), .out(n14521), .config_in(config_chain[35649:35644]), .config_rst(config_rst)); 
buffer_wire buffer_14521 (.in(n14521), .out(n14521_0));
mux13 mux_9356 (.in({n14400_1/**/, n10949_0, n10928_0, n10923_0, n10909_0, n10892_0, n10878_0, n10873_0, n10856_1, n8784, n8776, n7808, n7800}), .out(n14522), .config_in(config_chain[35655:35650]), .config_rst(config_rst)); 
buffer_wire buffer_14522 (.in(n14522), .out(n14522_0));
mux15 mux_9357 (.in({n14607_0, n11995_0/**/, n11986_0, n11983_0, n11960_0, n11957_0, n11932_0, n11929_0, n11920_1, n11829_0, n9086, n9078, n9070, n8102, n8094}), .out(n14523), .config_in(config_chain[35661:35656]), .config_rst(config_rst)); 
buffer_wire buffer_14523 (.in(n14523), .out(n14523_0));
mux13 mux_9358 (.in({n14408_1/**/, n10951_0, n10931_0, n10914_0, n10900_0, n10895_0, n10886_0, n10881_0, n10854_1, n8788, n8776, n7808, n7800}), .out(n14524), .config_in(config_chain[35667:35662]), .config_rst(config_rst)); 
buffer_wire buffer_14524 (.in(n14524), .out(n14524_0));
mux15 mux_9359 (.in({n14609_0, n11993_0, n11980_0, n11977_0, n11954_0, n11951_0, n11946_0, n11943_0, n11922_1/**/, n11861_0, n9086, n9078, n9070, n8102, n8094}), .out(n14525), .config_in(config_chain[35673:35668]), .config_rst(config_rst)); 
buffer_wire buffer_14525 (.in(n14525), .out(n14525_0));
mux13 mux_9360 (.in({n14416_1, n10953_0, n10922_0, n10917_0, n10908_0, n10903_0, n10872_0, n10867_0, n10852_1/**/, n8788, n8780, n7808, n7800}), .out(n14526), .config_in(config_chain[35679:35674]), .config_rst(config_rst)); 
buffer_wire buffer_14526 (.in(n14526), .out(n14526_0));
mux15 mux_9361 (.in({n14611_0, n11991_0, n11974_0, n11971_0, n11968_0, n11965_0, n11940_0, n11937_0, n11924_1/**/, n11883_0, n9086, n9078, n9070, n8102, n8094}), .out(n14527), .config_in(config_chain[35685:35680]), .config_rst(config_rst)); 
buffer_wire buffer_14527 (.in(n14527), .out(n14527_0));
mux13 mux_9362 (.in({n14424_1, n10955_0, n10930_0, n10925_0, n10894_0, n10889_0, n10880_0, n10875_0, n10850_1, n8788, n8780, n7812/**/, n7800}), .out(n14528), .config_in(config_chain[35691:35686]), .config_rst(config_rst)); 
buffer_wire buffer_14528 (.in(n14528), .out(n14528_0));
mux15 mux_9363 (.in({n14613_0, n12009_0, n11988_0, n11985_0, n11962_0, n11959_0, n11934_0, n11931_0, n11906_1/**/, n11905_0, n9086, n9078, n9070, n8102, n8094}), .out(n14529), .config_in(config_chain[35697:35692]), .config_rst(config_rst)); 
buffer_wire buffer_14529 (.in(n14529), .out(n14529_0));
mux13 mux_9364 (.in({n14440_1, n10935_0/**/, n10916_0, n10911_0, n10902_0, n10897_0, n10883_0, n10866_1, n10848_1, n8788, n8780, n7812, n7804}), .out(n14530), .config_in(config_chain[35703:35698]), .config_rst(config_rst)); 
buffer_wire buffer_14530 (.in(n14530), .out(n14530_0));
mux3 mux_9365 (.in({n12167_0, n12166_1/**/, n9180}), .out(n14531), .config_in(config_chain[35705:35704]), .config_rst(config_rst)); 
buffer_wire buffer_14531 (.in(n14531), .out(n14531_0));
mux15 mux_9366 (.in({n14444_1, n11201_0, n11182_0, n11177_0, n11175_0, n11166_0, n11161_0, n11147_0, n11130_1, n11110_1, n8886, n8878/**/, n7910, n7902, n7894}), .out(n14532), .config_in(config_chain[35711:35706]), .config_rst(config_rst)); 
buffer_wire buffer_14532 (.in(n14532), .out(n14532_0));
mux4 mux_9367 (.in({n12251_0, n12168_1, n9184, n8188}), .out(n14533), .config_in(config_chain[35713:35712]), .config_rst(config_rst)); 
buffer_wire buffer_14533 (.in(n14533), .out(n14533_0));
mux15 mux_9368 (.in({n14446_1, n11203_0, n11197_0, n11190_0/**/, n11185_0, n11169_0, n11152_0, n11138_0, n11133_0, n11046_2, n8890, n8878, n7910, n7902, n7894}), .out(n14534), .config_in(config_chain[35719:35714]), .config_rst(config_rst)); 
buffer_wire buffer_14534 (.in(n14534), .out(n14534_0));
mux3 mux_9369 (.in({n12253_0, n12170_1, n8192}), .out(n14535), .config_in(config_chain[35721:35720]), .config_rst(config_rst)); 
buffer_wire buffer_14535 (.in(n14535), .out(n14535_0));
mux15 mux_9370 (.in({n14448_1, n11205_0, n11193_0, n11176_0, n11174_0, n11160_0, n11155_0, n11146_0, n11141_0, n11128_1, n8890/**/, n8882, n7910, n7902, n7894}), .out(n14536), .config_in(config_chain[35727:35722]), .config_rst(config_rst)); 
buffer_wire buffer_14536 (.in(n14536), .out(n14536_0));
mux3 mux_9371 (.in({n12255_0, n12172_1/**/, n8192}), .out(n14537), .config_in(config_chain[35729:35728]), .config_rst(config_rst)); 
buffer_wire buffer_14537 (.in(n14537), .out(n14537_0));
mux15 mux_9372 (.in({n14450_1/**/, n11207_0, n11196_0, n11184_0, n11179_0, n11168_0, n11163_0, n11149_0, n11132_0, n11126_1, n8890, n8882, n8874, n7902, n7894}), .out(n14538), .config_in(config_chain[35735:35730]), .config_rst(config_rst)); 
buffer_wire buffer_14538 (.in(n14538), .out(n14538_0));
mux3 mux_9373 (.in({n12257_0, n12174_1, n8196}), .out(n14539), .config_in(config_chain[35737:35736]), .config_rst(config_rst)); 
buffer_wire buffer_14539 (.in(n14539), .out(n14539_0));
mux14 mux_9374 (.in({n14452_1, n11209_0, n11192_0/**/, n11187_0, n11171_0, n11154_0, n11140_0, n11135_0, n11124_1, n8890, n8882, n8874, n7906, n7894}), .out(n14540), .config_in(config_chain[35743:35738]), .config_rst(config_rst)); 
buffer_wire buffer_14540 (.in(n14540), .out(n14540_0));
mux3 mux_9375 (.in({n12259_0, n12176_1/**/, n8200}), .out(n14541), .config_in(config_chain[35745:35744]), .config_rst(config_rst)); 
buffer_wire buffer_14541 (.in(n14541), .out(n14541_0));
mux14 mux_9376 (.in({n14454_1, n11211_0, n11195_0, n11178_0, n11162_0, n11157_0, n11148_0, n11143_0, n11122_1/**/, n8890, n8882, n8874, n7906, n7898}), .out(n14542), .config_in(config_chain[35751:35746]), .config_rst(config_rst)); 
buffer_wire buffer_14542 (.in(n14542), .out(n14542_0));
mux3 mux_9377 (.in({n12261_0, n12178_1/**/, n8204}), .out(n14543), .config_in(config_chain[35753:35752]), .config_rst(config_rst)); 
buffer_wire buffer_14543 (.in(n14543), .out(n14543_0));
mux13 mux_9378 (.in({n14456_1, n11213_0, n11186_0, n11181_0, n11170_0/**/, n11165_0, n11151_0, n11134_0, n11120_1, n8882, n8874, n7906, n7898}), .out(n14544), .config_in(config_chain[35759:35754]), .config_rst(config_rst)); 
buffer_wire buffer_14544 (.in(n14544), .out(n14544_0));
mux3 mux_9379 (.in({n12263_0/**/, n12180_1, n9168}), .out(n14545), .config_in(config_chain[35761:35760]), .config_rst(config_rst)); 
buffer_wire buffer_14545 (.in(n14545), .out(n14545_0));
mux13 mux_9380 (.in({n14458_1, n11215_0, n11194_0, n11189_0, n11173_0, n11156_0, n11142_0, n11137_0, n11118_1/**/, n8886, n8874, n7906, n7898}), .out(n14546), .config_in(config_chain[35767:35762]), .config_rst(config_rst)); 
buffer_wire buffer_14546 (.in(n14546), .out(n14546_0));
mux3 mux_9381 (.in({n12265_0, n12182_1, n9168}), .out(n14547), .config_in(config_chain[35769:35768]), .config_rst(config_rst)); 
buffer_wire buffer_14547 (.in(n14547), .out(n14547_0));
mux13 mux_9382 (.in({n14460_1, n11217_0, n11180_0, n11164_0, n11159_0, n11150_0, n11145_0, n11116_1, n11109_0, n8886, n8878, n7906, n7898/**/}), .out(n14548), .config_in(config_chain[35775:35770]), .config_rst(config_rst)); 
buffer_wire buffer_14548 (.in(n14548), .out(n14548_0));
mux3 mux_9383 (.in({n12267_0/**/, n12184_1, n9172}), .out(n14549), .config_in(config_chain[35777:35776]), .config_rst(config_rst)); 
buffer_wire buffer_14549 (.in(n14549), .out(n14549_0));
mux13 mux_9384 (.in({n14462_1, n11219_0, n11188_0, n11183_0, n11172_0, n11167_0, n11136_0, n11131_0, n11114_1, n8886, n8878/**/, n7910, n7898}), .out(n14550), .config_in(config_chain[35783:35778]), .config_rst(config_rst)); 
buffer_wire buffer_14550 (.in(n14550), .out(n14550_0));
mux3 mux_9385 (.in({n12269_0, n12186_1/**/, n9176}), .out(n14551), .config_in(config_chain[35785:35784]), .config_rst(config_rst)); 
buffer_wire buffer_14551 (.in(n14551), .out(n14551_0));
mux13 mux_9386 (.in({n14442_1, n11199_0, n11191_0, n11158_0, n11153_0, n11144_0, n11139_0, n11112_1/**/, n11108_1, n8886, n8878, n7910, n7902}), .out(n14552), .config_in(config_chain[35791:35786]), .config_rst(config_rst)); 
buffer_wire buffer_14552 (.in(n14552), .out(n14552_0));
mux3 mux_9387 (.in({n12189_0, n12188_1, n9184}), .out(n14553), .config_in(config_chain[35793:35792]), .config_rst(config_rst)); 
buffer_wire buffer_14553 (.in(n14553), .out(n14553_0));
mux16 mux_9388 (.in({n14466_1, n11467_0, n11449_0, n11444_0, n11440_0, n11436_0/**/, n11421_0, n11411_0, n11406_0, n11376_1, n11353_0, n8984, n8976, n8008, n8000, n7992}), .out(n14554), .config_in(config_chain[35799:35794]), .config_rst(config_rst)); 
buffer_wire buffer_14554 (.in(n14554), .out(n14554_0));
mux4 mux_9389 (.in({n12191_0, n12190_0, n9184, n8188}), .out(n14555), .config_in(config_chain[35801:35800]), .config_rst(config_rst)); 
buffer_wire buffer_14555 (.in(n14555), .out(n14555_0));
mux16 mux_9390 (.in({n14468_1, n11469_0, n11462_0/**/, n11458_0, n11443_0, n11435_0, n11430_0, n11405_0, n11400_0, n11394_1, n11375_0, n8984, n8976, n8008, n8000, n7992}), .out(n14556), .config_in(config_chain[35807:35802]), .config_rst(config_rst)); 
buffer_wire buffer_14556 (.in(n14556), .out(n14556_0));
mux3 mux_9391 (.in({n12193_0, n12192_0, n8192}), .out(n14557), .config_in(config_chain[35809:35808]), .config_rst(config_rst)); 
buffer_wire buffer_14557 (.in(n14557), .out(n14557_0));
mux15 mux_9392 (.in({n14470_1, n11471_0, n11457_0, n11452_0, n11429_0, n11424_0/**/, n11414_0, n11399_0, n11397_0, n11392_1, n8984, n8976, n8008, n8000, n7992}), .out(n14558), .config_in(config_chain[35815:35810]), .config_rst(config_rst)); 
buffer_wire buffer_14558 (.in(n14558), .out(n14558_0));
mux3 mux_9393 (.in({n12195_0/**/, n12194_0, n8196}), .out(n14559), .config_in(config_chain[35817:35816]), .config_rst(config_rst)); 
buffer_wire buffer_14559 (.in(n14559), .out(n14559_0));
mux15 mux_9394 (.in({n14472_1, n11473_0, n11451_0, n11446_0, n11438_0, n11423_0, n11419_0, n11413_0, n11408_0, n11390_1, n8984, n8976, n8008/**/, n8000, n7992}), .out(n14560), .config_in(config_chain[35823:35818]), .config_rst(config_rst)); 
buffer_wire buffer_14560 (.in(n14560), .out(n14560_0));
mux3 mux_9395 (.in({n12197_0, n12196_0, n8196}), .out(n14561), .config_in(config_chain[35825:35824]), .config_rst(config_rst)); 
buffer_wire buffer_14561 (.in(n14561), .out(n14561_0));
mux15 mux_9396 (.in({n14474_1, n11475_0, n11460_0, n11445_0, n11441_0, n11437_0, n11432_0, n11407_0, n11402_0, n11388_1, n8984, n8976, n8008, n8000, n7992}), .out(n14562), .config_in(config_chain[35831:35826]), .config_rst(config_rst)); 
buffer_wire buffer_14562 (.in(n14562), .out(n14562_0));
mux3 mux_9397 (.in({n12199_0, n12198_0, n8200/**/}), .out(n14563), .config_in(config_chain[35833:35832]), .config_rst(config_rst)); 
buffer_wire buffer_14563 (.in(n14563), .out(n14563_0));
mux15 mux_9398 (.in({n14476_1, n11477_0, n11463_0, n11459_0, n11454_0, n11431_0, n11426_0, n11416_0, n11401_0, n11386_1/**/, n8988, n8980, n8972, n8004, n7996}), .out(n14564), .config_in(config_chain[35839:35834]), .config_rst(config_rst)); 
buffer_wire buffer_14564 (.in(n14564), .out(n14564_0));
mux3 mux_9399 (.in({n12201_0, n12200_0/**/, n8204}), .out(n14565), .config_in(config_chain[35841:35840]), .config_rst(config_rst)); 
buffer_wire buffer_14565 (.in(n14565), .out(n14565_0));
mux15 mux_9400 (.in({n14478_1, n11479_0, n11453_0, n11448_0, n11425_0, n11420_0, n11415_0, n11410_0, n11384_1/**/, n11352_1, n8988, n8980, n8972, n8004, n7996}), .out(n14566), .config_in(config_chain[35847:35842]), .config_rst(config_rst)); 
buffer_wire buffer_14566 (.in(n14566), .out(n14566_0));
mux3 mux_9401 (.in({n12203_0, n12202_0/**/, n9168}), .out(n14567), .config_in(config_chain[35849:35848]), .config_rst(config_rst)); 
buffer_wire buffer_14567 (.in(n14567), .out(n14567_0));
mux15 mux_9402 (.in({n14480_1, n11481_0, n11447_0, n11442_0/**/, n11439_0, n11434_0, n11409_0, n11404_0, n11382_1, n11374_1, n8988, n8980, n8972, n8004, n7996}), .out(n14568), .config_in(config_chain[35855:35850]), .config_rst(config_rst)); 
buffer_wire buffer_14568 (.in(n14568), .out(n14568_0));
mux3 mux_9403 (.in({n12205_0/**/, n12204_0, n9172}), .out(n14569), .config_in(config_chain[35857:35856]), .config_rst(config_rst)); 
buffer_wire buffer_14569 (.in(n14569), .out(n14569_0));
mux15 mux_9404 (.in({n14482_1, n11483_0, n11461_0, n11456_0, n11433_0/**/, n11428_0, n11403_0, n11398_0, n11396_1, n11380_1, n8988, n8980, n8972, n8004, n7996}), .out(n14570), .config_in(config_chain[35863:35858]), .config_rst(config_rst)); 
buffer_wire buffer_14570 (.in(n14570), .out(n14570_0));
mux3 mux_9405 (.in({n12207_0, n12206_0, n9172}), .out(n14571), .config_in(config_chain[35865:35864]), .config_rst(config_rst)); 
buffer_wire buffer_14571 (.in(n14571), .out(n14571_0));
mux15 mux_9406 (.in({n14484_1, n11465_0, n11455_0/**/, n11450_0, n11427_0, n11422_0, n11418_0, n11417_0, n11412_0, n11378_1, n8988, n8980, n8972, n8004, n7996}), .out(n14572), .config_in(config_chain[35871:35866]), .config_rst(config_rst)); 
buffer_wire buffer_14572 (.in(n14572), .out(n14572_0));
mux3 mux_9407 (.in({n12209_0, n12208_0/**/, n9176}), .out(n14573), .config_in(config_chain[35873:35872]), .config_rst(config_rst)); 
buffer_wire buffer_14573 (.in(n14573), .out(n14573_0));
mux16 mux_9408 (.in({n14488_1/**/, n11731_0, n11721_0, n11716_0, n11693_0, n11688_0, n11684_0, n11680_0, n11665_0, n11642_1, n11597_0, n9082, n9074, n8106, n8098, n8090}), .out(n14574), .config_in(config_chain[35879:35874]), .config_rst(config_rst)); 
buffer_wire buffer_14574 (.in(n14574), .out(n14574_0));
mux4 mux_9409 (.in({n12211_0, n12210_0, n9184, n8188}), .out(n14575), .config_in(config_chain[35881:35880]), .config_rst(config_rst)); 
buffer_wire buffer_14575 (.in(n14575), .out(n14575_0));
mux16 mux_9410 (.in({n14490_1/**/, n11733_0, n11715_0, n11710_0, n11706_0, n11702_0, n11687_0, n11679_0, n11674_0, n11660_1, n11619_0, n9082, n9074, n8106, n8098, n8090}), .out(n14576), .config_in(config_chain[35887:35882]), .config_rst(config_rst)); 
buffer_wire buffer_14576 (.in(n14576), .out(n14576_0));
mux3 mux_9411 (.in({n12213_0, n12212_0, n8192}), .out(n14577), .config_in(config_chain[35889:35888]), .config_rst(config_rst)); 
buffer_wire buffer_14577 (.in(n14577), .out(n14577_0));
mux15 mux_9412 (.in({n14492_1, n11735_0, n11724_0, n11709_0, n11701_0, n11696_0, n11673_0, n11668_0, n11658_1/**/, n11641_0, n9082, n9074, n8106, n8098, n8090}), .out(n14578), .config_in(config_chain[35895:35890]), .config_rst(config_rst)); 
buffer_wire buffer_14578 (.in(n14578), .out(n14578_0));
mux3 mux_9413 (.in({n12215_0, n12214_0/**/, n8196}), .out(n14579), .config_in(config_chain[35897:35896]), .config_rst(config_rst)); 
buffer_wire buffer_14579 (.in(n14579), .out(n14579_0));
mux15 mux_9414 (.in({n14494_1, n11737_0, n11723_0, n11718_0, n11695_0, n11690_0, n11682_0, n11667_0, n11663_0, n11656_1, n9082/**/, n9074, n8106, n8098, n8090}), .out(n14580), .config_in(config_chain[35903:35898]), .config_rst(config_rst)); 
buffer_wire buffer_14580 (.in(n14580), .out(n14580_0));
mux3 mux_9415 (.in({n12217_0, n12216_0, n8200}), .out(n14581), .config_in(config_chain[35905:35904]), .config_rst(config_rst)); 
buffer_wire buffer_14581 (.in(n14581), .out(n14581_0));
mux15 mux_9416 (.in({n14496_1, n11739_0, n11717_0, n11712_0, n11704_0, n11689_0, n11685_0, n11681_0, n11676_0, n11654_1, n9082, n9074, n8106, n8098, n8090/**/}), .out(n14582), .config_in(config_chain[35911:35906]), .config_rst(config_rst)); 
buffer_wire buffer_14582 (.in(n14582), .out(n14582_0));
mux3 mux_9417 (.in({n12219_0, n12218_0, n8200}), .out(n14583), .config_in(config_chain[35913:35912]), .config_rst(config_rst)); 
buffer_wire buffer_14583 (.in(n14583), .out(n14583_0));
mux15 mux_9418 (.in({n14498_1, n11741_0, n11726_0, n11711_0, n11707_0, n11703_0/**/, n11698_0, n11675_0, n11670_0, n11652_1, n9086, n9078, n9070, n8102, n8094}), .out(n14584), .config_in(config_chain[35919:35914]), .config_rst(config_rst)); 
buffer_wire buffer_14584 (.in(n14584), .out(n14584_0));
mux3 mux_9419 (.in({n12221_0/**/, n12220_0, n8204}), .out(n14585), .config_in(config_chain[35921:35920]), .config_rst(config_rst)); 
buffer_wire buffer_14585 (.in(n14585), .out(n14585_0));
mux15 mux_9420 (.in({n14500_1, n11743_0, n11725_0, n11720_0, n11697_0, n11692_0/**/, n11669_0, n11664_0, n11650_1, n11596_2, n9086, n9078, n9070, n8102, n8094}), .out(n14586), .config_in(config_chain[35927:35922]), .config_rst(config_rst)); 
buffer_wire buffer_14586 (.in(n14586), .out(n14586_0));
mux3 mux_9421 (.in({n12223_0, n12222_0, n9168}), .out(n14587), .config_in(config_chain[35929:35928]), .config_rst(config_rst)); 
buffer_wire buffer_14587 (.in(n14587), .out(n14587_0));
mux15 mux_9422 (.in({n14502_1, n11745_0, n11719_0, n11714_0, n11691_0, n11686_0, n11683_0, n11678_0, n11648_1, n11618_1, n9086, n9078, n9070, n8102, n8094}), .out(n14588), .config_in(config_chain[35935:35930]), .config_rst(config_rst)); 
buffer_wire buffer_14588 (.in(n14588), .out(n14588_0));
mux3 mux_9423 (.in({n12225_0, n12224_0/**/, n9172}), .out(n14589), .config_in(config_chain[35937:35936]), .config_rst(config_rst)); 
buffer_wire buffer_14589 (.in(n14589), .out(n14589_0));
mux15 mux_9424 (.in({n14504_1, n11747_0, n11713_0, n11708_0, n11705_0, n11700_0, n11677_0, n11672_0/**/, n11646_1, n11640_1, n9086, n9078, n9070, n8102, n8094}), .out(n14590), .config_in(config_chain[35943:35938]), .config_rst(config_rst)); 
buffer_wire buffer_14590 (.in(n14590), .out(n14590_0));
mux3 mux_9425 (.in({n12227_0, n12226_0/**/, n9176}), .out(n14591), .config_in(config_chain[35945:35944]), .config_rst(config_rst)); 
buffer_wire buffer_14591 (.in(n14591), .out(n14591_0));
mux15 mux_9426 (.in({n14506_1, n11729_0/**/, n11727_0, n11722_0, n11699_0, n11694_0, n11671_0, n11666_0, n11662_1, n11644_1, n9086, n9078, n9070, n8102, n8094}), .out(n14592), .config_in(config_chain[35951:35946]), .config_rst(config_rst)); 
buffer_wire buffer_14592 (.in(n14592), .out(n14592_0));
mux3 mux_9427 (.in({n12229_0, n12228_0, n9176}), .out(n14593), .config_in(config_chain[35953:35952]), .config_rst(config_rst)); 
buffer_wire buffer_14593 (.in(n14593), .out(n14593_0));
mux16 mux_9428 (.in({n14510_1, n11993_0, n11983_0, n11978_0/**/, n11957_0, n11952_0, n11944_0, n11929_0, n11926_1, n11906_1, n11829_0, n9180, n9172, n8204, n8196, n8188}), .out(n14594), .config_in(config_chain[35959:35954]), .config_rst(config_rst)); 
buffer_wire buffer_14594 (.in(n14594), .out(n14594_0));
mux4 mux_9429 (.in({n12231_0, n12230_0, n9184, n8188}), .out(n14595), .config_in(config_chain[35961:35960]), .config_rst(config_rst)); 
buffer_wire buffer_14595 (.in(n14595), .out(n14595_0));
mux16 mux_9430 (.in({n14512_1, n11995_0, n11977_0, n11972_0, n11966_0, n11951_0, n11948_0/**/, n11943_0, n11938_0, n11924_1, n11861_0, n9180, n9172, n8204, n8196, n8188}), .out(n14596), .config_in(config_chain[35967:35962]), .config_rst(config_rst)); 
buffer_wire buffer_14596 (.in(n14596), .out(n14596_0));
mux3 mux_9431 (.in({n12233_0, n12232_0, n8188}), .out(n14597), .config_in(config_chain[35969:35968]), .config_rst(config_rst)); 
buffer_wire buffer_14597 (.in(n14597), .out(n14597_0));
mux15 mux_9432 (.in({n14514_1, n11997_0, n11986_0, n11971_0, n11965_0, n11960_0, n11937_0/**/, n11932_0, n11922_1, n11883_0, n9180, n9172, n8204, n8196, n8188}), .out(n14598), .config_in(config_chain[35975:35970]), .config_rst(config_rst)); 
buffer_wire buffer_14598 (.in(n14598), .out(n14598_0));
mux3 mux_9433 (.in({n12235_0, n12234_0, n8192}), .out(n14599), .config_in(config_chain[35977:35976]), .config_rst(config_rst)); 
buffer_wire buffer_14599 (.in(n14599), .out(n14599_0));
mux15 mux_9434 (.in({n14516_1, n11999_0, n11985_0, n11980_0, n11959_0, n11954_0, n11946_0, n11931_0/**/, n11920_1, n11905_0, n9180, n9172, n8204, n8196, n8188}), .out(n14600), .config_in(config_chain[35983:35978]), .config_rst(config_rst)); 
buffer_wire buffer_14600 (.in(n14600), .out(n14600_0));
mux3 mux_9435 (.in({n12237_0, n12236_0, n8196}), .out(n14601), .config_in(config_chain[35985:35984]), .config_rst(config_rst)); 
buffer_wire buffer_14601 (.in(n14601), .out(n14601_0));
mux15 mux_9436 (.in({n14518_1, n12001_0, n11979_0, n11974_0, n11968_0, n11953_0, n11945_0, n11940_0, n11927_0, n11918_1, n9180, n9172, n8204, n8196, n8188}), .out(n14602), .config_in(config_chain[35991:35986]), .config_rst(config_rst)); 
buffer_wire buffer_14602 (.in(n14602), .out(n14602_0));
mux3 mux_9437 (.in({n12239_0/**/, n12238_0, n8200}), .out(n14603), .config_in(config_chain[35993:35992]), .config_rst(config_rst)); 
buffer_wire buffer_14603 (.in(n14603), .out(n14603_0));
mux15 mux_9438 (.in({n14520_1, n12003_0, n11988_0, n11973_0, n11967_0, n11962_0, n11949_0/**/, n11939_0, n11934_0, n11916_1, n9184, n9176, n9168, n8200, n8192}), .out(n14604), .config_in(config_chain[35999:35994]), .config_rst(config_rst)); 
buffer_wire buffer_14604 (.in(n14604), .out(n14604_0));
mux3 mux_9439 (.in({n12241_0, n12240_0, n8204}), .out(n14605), .config_in(config_chain[36001:36000]), .config_rst(config_rst)); 
buffer_wire buffer_14605 (.in(n14605), .out(n14605_0));
mux15 mux_9440 (.in({n14522_1, n12005_0, n11987_0, n11982_0, n11961_0, n11956_0, n11933_0, n11928_0, n11914_1, n11828_2, n9184, n9176, n9168, n8200, n8192}), .out(n14606), .config_in(config_chain[36007:36002]), .config_rst(config_rst)); 
buffer_wire buffer_14606 (.in(n14606), .out(n14606_0));
mux3 mux_9441 (.in({n12243_0, n12242_0, n8204}), .out(n14607), .config_in(config_chain[36009:36008]), .config_rst(config_rst)); 
buffer_wire buffer_14607 (.in(n14607), .out(n14607_0));
mux15 mux_9442 (.in({n14524_1, n12007_0, n11981_0, n11976_0, n11955_0, n11950_0, n11947_0, n11942_0, n11912_1, n11860_2, n9184, n9176, n9168, n8200, n8192}), .out(n14608), .config_in(config_chain[36015:36010]), .config_rst(config_rst)); 
buffer_wire buffer_14608 (.in(n14608), .out(n14608_0));
mux3 mux_9443 (.in({n12245_0, n12244_0, n9168}), .out(n14609), .config_in(config_chain[36017:36016]), .config_rst(config_rst)); 
buffer_wire buffer_14609 (.in(n14609), .out(n14609_0));
mux15 mux_9444 (.in({n14526_1, n12009_0, n11975_0, n11970_0, n11969_0, n11964_0, n11941_0, n11936_0, n11910_1, n11882_1, n9184, n9176, n9168, n8200, n8192}), .out(n14610), .config_in(config_chain[36023:36018]), .config_rst(config_rst)); 
buffer_wire buffer_14610 (.in(n14610), .out(n14610_0));
mux3 mux_9445 (.in({n12247_0, n12246_0, n9172}), .out(n14611), .config_in(config_chain[36025:36024]), .config_rst(config_rst)); 
buffer_wire buffer_14611 (.in(n14611), .out(n14611_0));
mux15 mux_9446 (.in({n14528_1, n11991_0, n11989_0, n11984_0, n11963_0, n11958_0/**/, n11935_0, n11930_0, n11908_1, n11904_1, n9184, n9176, n9168, n8200, n8192}), .out(n14612), .config_in(config_chain[36031:36026]), .config_rst(config_rst)); 
buffer_wire buffer_14612 (.in(n14612), .out(n14612_0));
mux3 mux_9447 (.in({n12249_0, n12248_0, n9176}), .out(n14613), .config_in(config_chain[36033:36032]), .config_rst(config_rst)); 
buffer_wire buffer_14613 (.in(n14613), .out(n14613_0));
mux3 mux_9448 (.in({n9898_0/**/, n9271, n8382}), .out(n14614), .config_in(config_chain[36035:36034]), .config_rst(config_rst)); 
buffer_wire buffer_14614 (.in(n14614), .out(n14614_0));
mux12 mux_9449 (.in({n14751_1, n10676_0, n10660_0, n10644_0, n10606_1, n10522_2, n9373, n9364, n9358, n8594, n8586, n8578}), .out(n14615), .config_in(config_chain[36041:36036]), .config_rst(config_rst)); 
buffer_wire buffer_14615 (.in(n14615), .out(n14615_0));
mux3 mux_9450 (.in({n9756_2, n9271, n8382}), .out(n14616), .config_in(config_chain[36043:36042]), .config_rst(config_rst)); 
buffer_wire buffer_14616 (.in(n14616), .out(n14616_0));
mux12 mux_9451 (.in({n14773_1, n10954_0, n10934_0/**/, n10916_0, n10900_0, n10884_1, n9421, n9412, n9406, n8692, n8684, n8676}), .out(n14617), .config_in(config_chain[36049:36044]), .config_rst(config_rst)); 
buffer_wire buffer_14617 (.in(n14617), .out(n14617_0));
mux3 mux_9452 (.in({n9754_2, n9271, n8382}), .out(n14618), .config_in(config_chain[36051:36050]), .config_rst(config_rst)); 
buffer_wire buffer_14618 (.in(n14618), .out(n14618_0));
mux12 mux_9453 (.in({n14707_1, n10170_0, n10132_0, n10116_0, n10102_1/**/, n10008_2, n9277, n9268, n9262, n8398, n8390, n8382}), .out(n14619), .config_in(config_chain[36057:36052]), .config_rst(config_rst)); 
buffer_wire buffer_14619 (.in(n14619), .out(n14619_0));
mux3 mux_9454 (.in({n9752_2, n9271, n8382}), .out(n14620), .config_in(config_chain[36059:36058]), .config_rst(config_rst)); 
buffer_wire buffer_14620 (.in(n14620), .out(n14620_0));
mux12 mux_9455 (.in({n14729_1, n10422_0/**/, n10406_0, n10368_0, n10352_1, n10264_2, n9325, n9316, n9310, n8496, n8488, n8480}), .out(n14621), .config_in(config_chain[36065:36060]), .config_rst(config_rst)); 
buffer_wire buffer_14621 (.in(n14621), .out(n14621_0));
mux3 mux_9456 (.in({n9750_2, n9274, n8382}), .out(n14622), .config_in(config_chain[36067:36066]), .config_rst(config_rst)); 
buffer_wire buffer_14622 (.in(n14622), .out(n14622_0));
mux12 mux_9457 (.in({n14753_1, n10682_0, n10666_0/**/, n10628_0, n10612_1, n10524_2, n9373, n9367, n9358, n8594, n8586, n8578}), .out(n14623), .config_in(config_chain[36073:36068]), .config_rst(config_rst)); 
buffer_wire buffer_14623 (.in(n14623), .out(n14623_0));
mux3 mux_9458 (.in({n9748_2, n9274, n8386}), .out(n14624), .config_in(config_chain[36075:36074]), .config_rst(config_rst)); 
buffer_wire buffer_14624 (.in(n14624), .out(n14624_0));
mux12 mux_9459 (.in({n14775_1, n10940_0, n10922_0, n10906_0, n10868_1, n10784_2, n9421, n9415, n9406, n8692, n8684, n8676/**/}), .out(n14625), .config_in(config_chain[36081:36076]), .config_rst(config_rst)); 
buffer_wire buffer_14625 (.in(n14625), .out(n14625_0));
mux3 mux_9460 (.in({n9918_0, n9274, n8386}), .out(n14626), .config_in(config_chain[36083:36082]), .config_rst(config_rst)); 
buffer_wire buffer_14626 (.in(n14626), .out(n14626_0));
mux12 mux_9461 (.in({n14709_1, n10154_0, n10138_0/**/, n10122_0, n10108_1, n10010_2, n9277, n9271, n9262, n8398, n8390, n8382}), .out(n14627), .config_in(config_chain[36089:36084]), .config_rst(config_rst)); 
buffer_wire buffer_14627 (.in(n14627), .out(n14627_0));
mux3 mux_9462 (.in({n9896_0/**/, n9274, n8386}), .out(n14628), .config_in(config_chain[36091:36090]), .config_rst(config_rst)); 
buffer_wire buffer_14628 (.in(n14628), .out(n14628_0));
mux12 mux_9463 (.in({n14731_1, n10428_0/**/, n10390_0, n10374_0, n10358_1, n10266_2, n9325, n9319, n9310, n8496, n8488, n8480}), .out(n14629), .config_in(config_chain[36097:36092]), .config_rst(config_rst)); 
buffer_wire buffer_14629 (.in(n14629), .out(n14629_0));
mux3 mux_9464 (.in({n9876_0/**/, n9274, n8386}), .out(n14630), .config_in(config_chain[36099:36098]), .config_rst(config_rst)); 
buffer_wire buffer_14630 (.in(n14630), .out(n14630_0));
mux11 mux_9465 (.in({n14755_1, n10688_0, n10650_0, n10634_0, n10618_1, n9373, n9367, n9361, n8594, n8586, n8578}), .out(n14631), .config_in(config_chain[36105:36100]), .config_rst(config_rst)); 
buffer_wire buffer_14631 (.in(n14631), .out(n14631_0));
mux3 mux_9466 (.in({n9856_1, n9277, n8386}), .out(n14632), .config_in(config_chain[36107:36106]), .config_rst(config_rst)); 
buffer_wire buffer_14632 (.in(n14632), .out(n14632_0));
mux11 mux_9467 (.in({n14777_1, n10946_0, n10928_0/**/, n10890_0, n10874_1, n9421, n9415, n9409, n8692, n8684, n8676}), .out(n14633), .config_in(config_chain[36113:36108]), .config_rst(config_rst)); 
buffer_wire buffer_14633 (.in(n14633), .out(n14633_0));
mux3 mux_9468 (.in({n9916_0, n9277, n8390}), .out(n14634), .config_in(config_chain[36115:36114]), .config_rst(config_rst)); 
buffer_wire buffer_14634 (.in(n14634), .out(n14634_0));
mux11 mux_9469 (.in({n14711_1, n10160_0, n10144_0, n10128_0, n10092_1, n9277, n9271, n9265, n8398, n8390, n8382}), .out(n14635), .config_in(config_chain[36121:36116]), .config_rst(config_rst)); 
buffer_wire buffer_14635 (.in(n14635), .out(n14635_0));
mux3 mux_9470 (.in({n9894_0/**/, n9277, n8390}), .out(n14636), .config_in(config_chain[36123:36122]), .config_rst(config_rst)); 
buffer_wire buffer_14636 (.in(n14636), .out(n14636_0));
mux11 mux_9471 (.in({n14733_1, n10412_0, n10396_0, n10380_0, n10364_1, n9325, n9319, n9313, n8496, n8488, n8480}), .out(n14637), .config_in(config_chain[36129:36124]), .config_rst(config_rst)); 
buffer_wire buffer_14637 (.in(n14637), .out(n14637_0));
mux3 mux_9472 (.in({n9874_0/**/, n9277, n8390}), .out(n14638), .config_in(config_chain[36131:36130]), .config_rst(config_rst)); 
buffer_wire buffer_14638 (.in(n14638), .out(n14638_0));
mux11 mux_9473 (.in({n14757_1, n10672_0, n10656_0/**/, n10640_0, n10624_1, n9373, n9367, n9361, n9355, n8586, n8578}), .out(n14639), .config_in(config_chain[36137:36132]), .config_rst(config_rst)); 
buffer_wire buffer_14639 (.in(n14639), .out(n14639_0));
mux3 mux_9474 (.in({n9854_1, n9277, n8390}), .out(n14640), .config_in(config_chain[36139:36138]), .config_rst(config_rst)); 
buffer_wire buffer_14640 (.in(n14640), .out(n14640_0));
mux11 mux_9475 (.in({n14779_1, n10952_0, n10912_0, n10896_0, n10880_1/**/, n9421, n9415, n9409, n9403, n8684, n8676}), .out(n14641), .config_in(config_chain[36145:36140]), .config_rst(config_rst)); 
buffer_wire buffer_14641 (.in(n14641), .out(n14641_0));
mux3 mux_9476 (.in({n9914_0/**/, n9280, n8390}), .out(n14642), .config_in(config_chain[36147:36146]), .config_rst(config_rst)); 
buffer_wire buffer_14642 (.in(n14642), .out(n14642_0));
mux11 mux_9477 (.in({n14713_1, n10166_0, n10150_0, n10112_0, n10098_1, n9277, n9271, n9265, n9259, n8390, n8382}), .out(n14643), .config_in(config_chain[36153:36148]), .config_rst(config_rst)); 
buffer_wire buffer_14643 (.in(n14643), .out(n14643_0));
mux3 mux_9478 (.in({n9892_0/**/, n9280, n8394}), .out(n14644), .config_in(config_chain[36155:36154]), .config_rst(config_rst)); 
buffer_wire buffer_14644 (.in(n14644), .out(n14644_0));
mux11 mux_9479 (.in({n14735_1, n10418_0, n10402_0, n10386_0, n10348_1/**/, n9325, n9319, n9313, n9307, n8488, n8480}), .out(n14645), .config_in(config_chain[36161:36156]), .config_rst(config_rst)); 
buffer_wire buffer_14645 (.in(n14645), .out(n14645_0));
mux3 mux_9480 (.in({n9872_0, n9280, n8394}), .out(n14646), .config_in(config_chain[36163:36162]), .config_rst(config_rst)); 
buffer_wire buffer_14646 (.in(n14646), .out(n14646_0));
mux11 mux_9481 (.in({n14759_1, n10678_0/**/, n10662_0, n10646_0, n10608_1, n9373, n9367, n9361, n9355, n8590, n8578}), .out(n14647), .config_in(config_chain[36169:36164]), .config_rst(config_rst)); 
buffer_wire buffer_14647 (.in(n14647), .out(n14647_0));
mux3 mux_9482 (.in({n9852_1/**/, n9280, n8394}), .out(n14648), .config_in(config_chain[36171:36170]), .config_rst(config_rst)); 
buffer_wire buffer_14648 (.in(n14648), .out(n14648_0));
mux11 mux_9483 (.in({n14781_1, n10936_0, n10918_0, n10902_0, n10886_1, n9421, n9415, n9409, n9403, n8688, n8676/**/}), .out(n14649), .config_in(config_chain[36177:36172]), .config_rst(config_rst)); 
buffer_wire buffer_14649 (.in(n14649), .out(n14649_0));
mux3 mux_9484 (.in({n9912_0/**/, n9280, n8394}), .out(n14650), .config_in(config_chain[36179:36178]), .config_rst(config_rst)); 
buffer_wire buffer_14650 (.in(n14650), .out(n14650_0));
mux11 mux_9485 (.in({n14715_1, n10172_0, n10134_0, n10118_0, n10104_1, n9277, n9271, n9265, n9259, n8394, n8382}), .out(n14651), .config_in(config_chain[36185:36180]), .config_rst(config_rst)); 
buffer_wire buffer_14651 (.in(n14651), .out(n14651_0));
mux2 mux_9486 (.in({n9890_0, n8394}), .out(n14652), .config_in(config_chain[36186:36186]), .config_rst(config_rst)); 
buffer_wire buffer_14652 (.in(n14652), .out(n14652_0));
mux11 mux_9487 (.in({n14737_1, n10424_0, n10408_0, n10370_0, n10354_1, n9325, n9319, n9313, n9307, n8492, n8480}), .out(n14653), .config_in(config_chain[36192:36187]), .config_rst(config_rst)); 
buffer_wire buffer_14653 (.in(n14653), .out(n14653_0));
mux2 mux_9488 (.in({n9870_0, n8398}), .out(n14654), .config_in(config_chain[36193:36193]), .config_rst(config_rst)); 
buffer_wire buffer_14654 (.in(n14654), .out(n14654_0));
mux11 mux_9489 (.in({n14761_1, n10684_0, n10668_0, n10630_0, n10614_1, n9376, n9367, n9361, n9355, n8590, n8582}), .out(n14655), .config_in(config_chain[36199:36194]), .config_rst(config_rst)); 
buffer_wire buffer_14655 (.in(n14655), .out(n14655_0));
mux2 mux_9490 (.in({n9850_1/**/, n8398}), .out(n14656), .config_in(config_chain[36200:36200]), .config_rst(config_rst)); 
buffer_wire buffer_14656 (.in(n14656), .out(n14656_0));
mux11 mux_9491 (.in({n14783_1, n10942_0, n10924_0, n10908_0, n10870_1/**/, n9424, n9415, n9409, n9403, n8688, n8680}), .out(n14657), .config_in(config_chain[36206:36201]), .config_rst(config_rst)); 
buffer_wire buffer_14657 (.in(n14657), .out(n14657_0));
mux2 mux_9492 (.in({n9910_0/**/, n8398}), .out(n14658), .config_in(config_chain[36207:36207]), .config_rst(config_rst)); 
buffer_wire buffer_14658 (.in(n14658), .out(n14658_0));
mux11 mux_9493 (.in({n14717_1, n10156_0, n10140_0, n10124_0, n10110_1, n9280, n9271, n9265, n9259, n8394, n8386}), .out(n14659), .config_in(config_chain[36213:36208]), .config_rst(config_rst)); 
buffer_wire buffer_14659 (.in(n14659), .out(n14659_0));
mux2 mux_9494 (.in({n9888_0/**/, n8398}), .out(n14660), .config_in(config_chain[36214:36214]), .config_rst(config_rst)); 
buffer_wire buffer_14660 (.in(n14660), .out(n14660_0));
mux11 mux_9495 (.in({n14739_1, n10430_0, n10392_0, n10376_0/**/, n10360_1, n9328, n9319, n9313, n9307, n8492, n8484}), .out(n14661), .config_in(config_chain[36220:36215]), .config_rst(config_rst)); 
buffer_wire buffer_14661 (.in(n14661), .out(n14661_0));
mux2 mux_9496 (.in({n9868_0, n8398}), .out(n14662), .config_in(config_chain[36221:36221]), .config_rst(config_rst)); 
buffer_wire buffer_14662 (.in(n14662), .out(n14662_0));
mux11 mux_9497 (.in({n14763_1, n10690_0/**/, n10652_0, n10636_0, n10620_1, n9376, n9370, n9361, n9355, n8590, n8582}), .out(n14663), .config_in(config_chain[36227:36222]), .config_rst(config_rst)); 
buffer_wire buffer_14663 (.in(n14663), .out(n14663_0));
mux2 mux_9498 (.in({n9848_1, n9259}), .out(n14664), .config_in(config_chain[36228:36228]), .config_rst(config_rst)); 
buffer_wire buffer_14664 (.in(n14664), .out(n14664_0));
mux11 mux_9499 (.in({n14785_1, n10948_0, n10930_0, n10892_0, n10876_1, n9424, n9418, n9409, n9403, n8688, n8680/**/}), .out(n14665), .config_in(config_chain[36234:36229]), .config_rst(config_rst)); 
buffer_wire buffer_14665 (.in(n14665), .out(n14665_0));
mux2 mux_9500 (.in({n9908_0/**/, n9259}), .out(n14666), .config_in(config_chain[36235:36235]), .config_rst(config_rst)); 
buffer_wire buffer_14666 (.in(n14666), .out(n14666_0));
mux11 mux_9501 (.in({n14719_1, n10162_0, n10146_0, n10130_0, n10094_1, n9280, n9274, n9265, n9259, n8394, n8386}), .out(n14667), .config_in(config_chain[36241:36236]), .config_rst(config_rst)); 
buffer_wire buffer_14667 (.in(n14667), .out(n14667_0));
mux2 mux_9502 (.in({n9886_0/**/, n9259}), .out(n14668), .config_in(config_chain[36242:36242]), .config_rst(config_rst)); 
buffer_wire buffer_14668 (.in(n14668), .out(n14668_0));
mux11 mux_9503 (.in({n14741_1, n10414_0, n10398_0, n10382_0, n10366_1, n9328, n9322, n9313, n9307, n8492, n8484}), .out(n14669), .config_in(config_chain[36248:36243]), .config_rst(config_rst)); 
buffer_wire buffer_14669 (.in(n14669), .out(n14669_0));
mux2 mux_9504 (.in({n9866_0, n9259}), .out(n14670), .config_in(config_chain[36249:36249]), .config_rst(config_rst)); 
buffer_wire buffer_14670 (.in(n14670), .out(n14670_0));
mux11 mux_9505 (.in({n14765_1, n10674_0/**/, n10658_0, n10642_0, n10626_1, n9376, n9370, n9364, n9355, n8590, n8582}), .out(n14671), .config_in(config_chain[36255:36250]), .config_rst(config_rst)); 
buffer_wire buffer_14671 (.in(n14671), .out(n14671_0));
mux2 mux_9506 (.in({n9846_1/**/, n9259}), .out(n14672), .config_in(config_chain[36256:36256]), .config_rst(config_rst)); 
buffer_wire buffer_14672 (.in(n14672), .out(n14672_0));
mux11 mux_9507 (.in({n14787_1/**/, n10914_0, n10898_0, n10882_1, n10866_1, n9424, n9418, n9412, n9403, n8688, n8680}), .out(n14673), .config_in(config_chain[36262:36257]), .config_rst(config_rst)); 
buffer_wire buffer_14673 (.in(n14673), .out(n14673_0));
mux2 mux_9508 (.in({n9906_0, n9262}), .out(n14674), .config_in(config_chain[36263:36263]), .config_rst(config_rst)); 
buffer_wire buffer_14674 (.in(n14674), .out(n14674_0));
mux11 mux_9509 (.in({n14721_1, n10168_0, n10152_0, n10114_0, n10100_1, n9280, n9274, n9268, n9259, n8394, n8386}), .out(n14675), .config_in(config_chain[36269:36264]), .config_rst(config_rst)); 
buffer_wire buffer_14675 (.in(n14675), .out(n14675_0));
mux2 mux_9510 (.in({n9884_0/**/, n9262}), .out(n14676), .config_in(config_chain[36270:36270]), .config_rst(config_rst)); 
buffer_wire buffer_14676 (.in(n14676), .out(n14676_0));
mux11 mux_9511 (.in({n14743_1, n10420_0, n10404_0, n10388_0/**/, n10350_1, n9328, n9322, n9316, n9307, n8492, n8484}), .out(n14677), .config_in(config_chain[36276:36271]), .config_rst(config_rst)); 
buffer_wire buffer_14677 (.in(n14677), .out(n14677_0));
mux2 mux_9512 (.in({n9864_0, n9262}), .out(n14678), .config_in(config_chain[36277:36277]), .config_rst(config_rst)); 
buffer_wire buffer_14678 (.in(n14678), .out(n14678_0));
mux11 mux_9513 (.in({n14767_1, n10680_0, n10664_0/**/, n10648_0, n10610_1, n9376, n9370, n9364, n9358, n8590, n8582}), .out(n14679), .config_in(config_chain[36283:36278]), .config_rst(config_rst)); 
buffer_wire buffer_14679 (.in(n14679), .out(n14679_0));
mux2 mux_9514 (.in({n9844_1, n9262}), .out(n14680), .config_in(config_chain[36284:36284]), .config_rst(config_rst)); 
buffer_wire buffer_14680 (.in(n14680), .out(n14680_0));
mux11 mux_9515 (.in({n14789_1, n10938_0/**/, n10920_0, n10904_0, n10888_1, n9424, n9418, n9412, n9406, n8688, n8680}), .out(n14681), .config_in(config_chain[36290:36285]), .config_rst(config_rst)); 
buffer_wire buffer_14681 (.in(n14681), .out(n14681_0));
mux2 mux_9516 (.in({n9904_0/**/, n9262}), .out(n14682), .config_in(config_chain[36291:36291]), .config_rst(config_rst)); 
buffer_wire buffer_14682 (.in(n14682), .out(n14682_0));
mux11 mux_9517 (.in({n14723_1, n10174_0, n10136_0, n10120_0, n10106_1, n9280, n9274, n9268, n9262, n8394, n8386}), .out(n14683), .config_in(config_chain[36297:36292]), .config_rst(config_rst)); 
buffer_wire buffer_14683 (.in(n14683), .out(n14683_0));
mux2 mux_9518 (.in({n9882_0, n9265}), .out(n14684), .config_in(config_chain[36298:36298]), .config_rst(config_rst)); 
buffer_wire buffer_14684 (.in(n14684), .out(n14684_0));
mux11 mux_9519 (.in({n14745_1, n10426_0, n10410_0, n10372_0, n10356_1, n9328, n9322, n9316, n9310, n8492, n8484}), .out(n14685), .config_in(config_chain[36304:36299]), .config_rst(config_rst)); 
buffer_wire buffer_14685 (.in(n14685), .out(n14685_0));
mux2 mux_9520 (.in({n9862_0/**/, n9265}), .out(n14686), .config_in(config_chain[36305:36305]), .config_rst(config_rst)); 
buffer_wire buffer_14686 (.in(n14686), .out(n14686_0));
mux11 mux_9521 (.in({n14769_1, n10686_0, n10670_0, n10632_0, n10616_1, n9376, n9370, n9364, n9358, n8594, n8582}), .out(n14687), .config_in(config_chain[36311:36306]), .config_rst(config_rst)); 
buffer_wire buffer_14687 (.in(n14687), .out(n14687_0));
mux2 mux_9522 (.in({n9842_1, n9265}), .out(n14688), .config_in(config_chain[36312:36312]), .config_rst(config_rst)); 
buffer_wire buffer_14688 (.in(n14688), .out(n14688_0));
mux11 mux_9523 (.in({n14791_1, n10944_0, n10926_0, n10910_0, n10872_1, n9424, n9418, n9412, n9406, n8692, n8680}), .out(n14689), .config_in(config_chain[36318:36313]), .config_rst(config_rst)); 
buffer_wire buffer_14689 (.in(n14689), .out(n14689_0));
mux2 mux_9524 (.in({n9902_0, n9265}), .out(n14690), .config_in(config_chain[36319:36319]), .config_rst(config_rst)); 
buffer_wire buffer_14690 (.in(n14690), .out(n14690_0));
mux11 mux_9525 (.in({n14725_1, n10158_0, n10142_0, n10126_0, n10004_2, n9280, n9274, n9268, n9262, n8398, n8386}), .out(n14691), .config_in(config_chain[36325:36320]), .config_rst(config_rst)); 
buffer_wire buffer_14691 (.in(n14691), .out(n14691_0));
mux2 mux_9526 (.in({n9880_0, n9265}), .out(n14692), .config_in(config_chain[36326:36326]), .config_rst(config_rst)); 
buffer_wire buffer_14692 (.in(n14692), .out(n14692_0));
mux11 mux_9527 (.in({n14747_1, n10432_0, n10394_0, n10378_0, n10362_1, n9328, n9322, n9316, n9310, n8496, n8484}), .out(n14693), .config_in(config_chain[36332:36327]), .config_rst(config_rst)); 
buffer_wire buffer_14693 (.in(n14693), .out(n14693_0));
mux2 mux_9528 (.in({n9860_0, n9268}), .out(n14694), .config_in(config_chain[36333:36333]), .config_rst(config_rst)); 
buffer_wire buffer_14694 (.in(n14694), .out(n14694_0));
mux2 mux_9529 (.in({n12092_2/**/, n9652}), .out(n14695), .config_in(config_chain[36334:36334]), .config_rst(config_rst)); 
buffer_wire buffer_14695 (.in(n14695), .out(n14695_0));
mux2 mux_9530 (.in({n9840_1, n9268}), .out(n14696), .config_in(config_chain[36335:36335]), .config_rst(config_rst)); 
buffer_wire buffer_14696 (.in(n14696), .out(n14696_0));
mux2 mux_9531 (.in({n12122_2, n9652}), .out(n14697), .config_in(config_chain[36336:36336]), .config_rst(config_rst)); 
buffer_wire buffer_14697 (.in(n14697), .out(n14697_0));
mux2 mux_9532 (.in({n9900_0, n9268}), .out(n14698), .config_in(config_chain[36337:36337]), .config_rst(config_rst)); 
buffer_wire buffer_14698 (.in(n14698), .out(n14698_0));
mux10 mux_9533 (.in({n14727_2, n10164_0/**/, n10148_0, n10096_1, n10006_2, n9274, n9268, n9262, n8398, n8390}), .out(n14699), .config_in(config_chain[36343:36338]), .config_rst(config_rst)); 
buffer_wire buffer_14699 (.in(n14699), .out(n14699_0));
mux2 mux_9534 (.in({n9878_0, n9268}), .out(n14700), .config_in(config_chain[36344:36344]), .config_rst(config_rst)); 
buffer_wire buffer_14700 (.in(n14700), .out(n14700_0));
mux10 mux_9535 (.in({n14749_2, n10416_0, n10400_0, n10384_0, n10262_2, n9322, n9316, n9310, n8496, n8488}), .out(n14701), .config_in(config_chain[36350:36345]), .config_rst(config_rst)); 
buffer_wire buffer_14701 (.in(n14701), .out(n14701_0));
mux2 mux_9536 (.in({n9858_0, n9268}), .out(n14702), .config_in(config_chain[36351:36351]), .config_rst(config_rst)); 
buffer_wire buffer_14702 (.in(n14702), .out(n14702_0));
mux10 mux_9537 (.in({n14771_1, n10692_0, n10654_0, n10638_0, n10622_1, n9370, n9364, n9358, n8594, n8586}), .out(n14703), .config_in(config_chain[36357:36352]), .config_rst(config_rst)); 
buffer_wire buffer_14703 (.in(n14703), .out(n14703_0));
mux2 mux_9538 (.in({n9838_1/**/, n9271}), .out(n14704), .config_in(config_chain[36358:36358]), .config_rst(config_rst)); 
buffer_wire buffer_14704 (.in(n14704), .out(n14704_0));
mux10 mux_9539 (.in({n14793_1, n10950_0/**/, n10932_0, n10894_0, n10878_1, n9418, n9412, n9406, n8692, n8684}), .out(n14705), .config_in(config_chain[36364:36359]), .config_rst(config_rst)); 
buffer_wire buffer_14705 (.in(n14705), .out(n14705_0));
mux12 mux_9540 (.in({n14618_0, n10170_0, n10132_0/**/, n10116_0, n10102_1, n10008_2, n9325, n9316, n9310, n8496, n8488, n8480}), .out(n14706), .config_in(config_chain[36370:36365]), .config_rst(config_rst)); 
buffer_wire buffer_14706 (.in(n14706), .out(n14706_0));
mux13 mux_9541 (.in({n14795_1, n11186_0, n11176_0, n11146_1, n11136_1, n11108_1, n9472, n9466/**/, n9460, n9454, n8790, n8782, n8774}), .out(n14707), .config_in(config_chain[36376:36371]), .config_rst(config_rst)); 
buffer_wire buffer_14707 (.in(n14707), .out(n14707_0));
mux12 mux_9542 (.in({n14626_0, n10154_0, n10138_0/**/, n10122_0, n10108_1, n10010_2, n9325, n9319, n9310, n8496, n8488, n8480}), .out(n14708), .config_in(config_chain[36382:36377]), .config_rst(config_rst)); 
buffer_wire buffer_14708 (.in(n14708), .out(n14708_0));
mux13 mux_9543 (.in({n14797_1, n11208_0, n11198_0, n11168_0, n11158_0, n11130_1, n9472, n9466/**/, n9460, n9454, n8790, n8782, n8774}), .out(n14709), .config_in(config_chain[36388:36383]), .config_rst(config_rst)); 
buffer_wire buffer_14709 (.in(n14709), .out(n14709_0));
mux11 mux_9544 (.in({n14634_0, n10160_0, n10144_0/**/, n10128_0, n10092_1, n9325, n9319, n9313, n8496, n8488, n8480}), .out(n14710), .config_in(config_chain[36394:36389]), .config_rst(config_rst)); 
buffer_wire buffer_14710 (.in(n14710), .out(n14710_0));
mux13 mux_9545 (.in({n14799_1, n11192_0, n11182_0, n11152_1, n11142_1, n11132_1, n9472, n9466/**/, n9460, n9454, n8790, n8782, n8774}), .out(n14711), .config_in(config_chain[36400:36395]), .config_rst(config_rst)); 
buffer_wire buffer_14711 (.in(n14711), .out(n14711_0));
mux11 mux_9546 (.in({n14642_0, n10166_0, n10150_0, n10112_0/**/, n10098_1, n9325, n9319, n9313, n9307, n8488, n8480}), .out(n14712), .config_in(config_chain[36406:36401]), .config_rst(config_rst)); 
buffer_wire buffer_14712 (.in(n14712), .out(n14712_0));
mux13 mux_9547 (.in({n14801_1, n11214_0, n11204_0, n11174_0, n11164_0, n11154_0, n9472, n9466/**/, n9460, n9454, n8790, n8782, n8774}), .out(n14713), .config_in(config_chain[36412:36407]), .config_rst(config_rst)); 
buffer_wire buffer_14713 (.in(n14713), .out(n14713_0));
mux11 mux_9548 (.in({n14650_0/**/, n10172_0, n10134_0, n10118_0, n10104_1, n9325, n9319, n9313, n9307, n8492, n8480}), .out(n14714), .config_in(config_chain[36418:36413]), .config_rst(config_rst)); 
buffer_wire buffer_14714 (.in(n14714), .out(n14714_0));
mux13 mux_9549 (.in({n14803_1, n11196_0, n11188_0, n11178_0, n11148_1, n11138_1, n9472, n9466/**/, n9460, n9454, n8790, n8782, n8774}), .out(n14715), .config_in(config_chain[36424:36419]), .config_rst(config_rst)); 
buffer_wire buffer_14715 (.in(n14715), .out(n14715_0));
mux11 mux_9550 (.in({n14658_0, n10156_0, n10140_0/**/, n10124_0, n10110_1, n9328, n9319, n9313, n9307, n8492, n8484}), .out(n14716), .config_in(config_chain[36430:36425]), .config_rst(config_rst)); 
buffer_wire buffer_14716 (.in(n14716), .out(n14716_0));
mux12 mux_9551 (.in({n14805_1, n11218_0, n11210_0, n11200_0/**/, n11170_0, n11160_0, n9469, n9463, n9457, n9451, n8786, n8778}), .out(n14717), .config_in(config_chain[36436:36431]), .config_rst(config_rst)); 
buffer_wire buffer_14717 (.in(n14717), .out(n14717_0));
mux11 mux_9552 (.in({n14666_0, n10162_0, n10146_0, n10130_0, n10094_1/**/, n9328, n9322, n9313, n9307, n8492, n8484}), .out(n14718), .config_in(config_chain[36442:36437]), .config_rst(config_rst)); 
buffer_wire buffer_14718 (.in(n14718), .out(n14718_0));
mux11 mux_9553 (.in({n14807_1, n11194_0/**/, n11184_0, n11144_1, n11134_1, n9469, n9463, n9457, n9451, n8786, n8778}), .out(n14719), .config_in(config_chain[36448:36443]), .config_rst(config_rst)); 
buffer_wire buffer_14719 (.in(n14719), .out(n14719_0));
mux11 mux_9554 (.in({n14674_0, n10168_0/**/, n10152_0, n10114_0, n10100_1, n9328, n9322, n9316, n9307, n8492, n8484}), .out(n14720), .config_in(config_chain[36454:36449]), .config_rst(config_rst)); 
buffer_wire buffer_14720 (.in(n14720), .out(n14720_0));
mux11 mux_9555 (.in({n14809_1, n11216_0, n11206_0, n11166_0/**/, n11156_0, n9469, n9463, n9457, n9451, n8786, n8778}), .out(n14721), .config_in(config_chain[36460:36455]), .config_rst(config_rst)); 
buffer_wire buffer_14721 (.in(n14721), .out(n14721_0));
mux11 mux_9556 (.in({n14682_0/**/, n10174_0, n10136_0, n10120_0, n10106_1, n9328, n9322, n9316, n9310, n8492, n8484}), .out(n14722), .config_in(config_chain[36466:36461]), .config_rst(config_rst)); 
buffer_wire buffer_14722 (.in(n14722), .out(n14722_0));
mux11 mux_9557 (.in({n14811_1, n11190_0, n11180_0, n11150_1, n11140_1, n9469, n9463, n9457, n9451, n8786/**/, n8778}), .out(n14723), .config_in(config_chain[36472:36467]), .config_rst(config_rst)); 
buffer_wire buffer_14723 (.in(n14723), .out(n14723_0));
mux11 mux_9558 (.in({n14690_0, n10158_0, n10142_0/**/, n10126_0, n10004_2, n9328, n9322, n9316, n9310, n8496, n8484}), .out(n14724), .config_in(config_chain[36478:36473]), .config_rst(config_rst)); 
buffer_wire buffer_14724 (.in(n14724), .out(n14724_0));
mux11 mux_9559 (.in({n14813_1, n11212_0, n11202_0, n11172_0, n11162_0/**/, n9469, n9463, n9457, n9451, n8786, n8778}), .out(n14725), .config_in(config_chain[36484:36479]), .config_rst(config_rst)); 
buffer_wire buffer_14725 (.in(n14725), .out(n14725_0));
mux10 mux_9560 (.in({n14698_0, n10164_0, n10148_0/**/, n10096_1, n10006_2, n9322, n9316, n9310, n8496, n8488}), .out(n14726), .config_in(config_chain[36490:36485]), .config_rst(config_rst)); 
buffer_wire buffer_14726 (.in(n14726), .out(n14726_0));
mux2 mux_9561 (.in({n12144_2, n9652}), .out(n14727), .config_in(config_chain[36491:36491]), .config_rst(config_rst)); 
buffer_wire buffer_14727 (.in(n14727), .out(n14727_0));
mux12 mux_9562 (.in({n14620_0, n10422_0/**/, n10406_0, n10368_0, n10352_1, n10264_2, n9373, n9364, n9358, n8594, n8586, n8578}), .out(n14728), .config_in(config_chain[36497:36492]), .config_rst(config_rst)); 
buffer_wire buffer_14728 (.in(n14728), .out(n14728_0));
mux13 mux_9563 (.in({n14815_0, n11478_0/**/, n11468_0, n11430_0, n11420_0, n11352_2, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14729), .config_in(config_chain[36503:36498]), .config_rst(config_rst)); 
buffer_wire buffer_14729 (.in(n14729), .out(n14729_0));
mux12 mux_9564 (.in({n14628_0/**/, n10428_0, n10390_0, n10374_0, n10358_1, n10266_2, n9373, n9367, n9358, n8594, n8586, n8578}), .out(n14730), .config_in(config_chain[36509:36504]), .config_rst(config_rst)); 
buffer_wire buffer_14730 (.in(n14730), .out(n14730_0));
mux13 mux_9565 (.in({n14817_0, n11452_0/**/, n11442_0, n11412_1, n11402_1, n11374_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14731), .config_in(config_chain[36515:36510]), .config_rst(config_rst)); 
buffer_wire buffer_14731 (.in(n14731), .out(n14731_0));
mux11 mux_9566 (.in({n14636_0, n10412_0/**/, n10396_0, n10380_0, n10364_1, n9373, n9367, n9361, n8594, n8586, n8578}), .out(n14732), .config_in(config_chain[36521:36516]), .config_rst(config_rst)); 
buffer_wire buffer_14732 (.in(n14732), .out(n14732_0));
mux13 mux_9567 (.in({n14819_0, n11474_0, n11464_0, n11436_0/**/, n11426_0, n11396_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14733), .config_in(config_chain[36527:36522]), .config_rst(config_rst)); 
buffer_wire buffer_14733 (.in(n14733), .out(n14733_0));
mux11 mux_9568 (.in({n14644_0, n10418_0, n10402_0/**/, n10386_0, n10348_1, n9373, n9367, n9361, n9355, n8586, n8578}), .out(n14734), .config_in(config_chain[36533:36528]), .config_rst(config_rst)); 
buffer_wire buffer_14734 (.in(n14734), .out(n14734_0));
mux13 mux_9569 (.in({n14821_0, n11458_0, n11448_0, n11418_1, n11408_1, n11398_1/**/, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14735), .config_in(config_chain[36539:36534]), .config_rst(config_rst)); 
buffer_wire buffer_14735 (.in(n14735), .out(n14735_0));
mux11 mux_9570 (.in({n14652_0, n10424_0, n10408_0, n10370_0, n10354_1/**/, n9373, n9367, n9361, n9355, n8590, n8578}), .out(n14736), .config_in(config_chain[36545:36540]), .config_rst(config_rst)); 
buffer_wire buffer_14736 (.in(n14736), .out(n14736_0));
mux13 mux_9571 (.in({n14823_0, n11480_0, n11470_0, n11440_0, n11432_0/**/, n11422_0, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14737), .config_in(config_chain[36551:36546]), .config_rst(config_rst)); 
buffer_wire buffer_14737 (.in(n14737), .out(n14737_0));
mux11 mux_9572 (.in({n14660_0, n10430_0, n10392_0, n10376_0/**/, n10360_1, n9376, n9367, n9361, n9355, n8590, n8582}), .out(n14738), .config_in(config_chain[36557:36552]), .config_rst(config_rst)); 
buffer_wire buffer_14738 (.in(n14738), .out(n14738_0));
mux12 mux_9573 (.in({n14825_0, n11462_0, n11454_0, n11444_0, n11414_1, n11404_1, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14739), .config_in(config_chain[36563:36558]), .config_rst(config_rst)); 
buffer_wire buffer_14739 (.in(n14739), .out(n14739_0));
mux11 mux_9574 (.in({n14668_0, n10414_0/**/, n10398_0, n10382_0, n10366_1, n9376, n9370, n9361, n9355, n8590, n8582}), .out(n14740), .config_in(config_chain[36569:36564]), .config_rst(config_rst)); 
buffer_wire buffer_14740 (.in(n14740), .out(n14740_0));
mux11 mux_9575 (.in({n14827_0, n11476_0, n11466_0/**/, n11438_0, n11428_0, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14741), .config_in(config_chain[36575:36570]), .config_rst(config_rst)); 
buffer_wire buffer_14741 (.in(n14741), .out(n14741_0));
mux11 mux_9576 (.in({n14676_0, n10420_0/**/, n10404_0, n10388_0, n10350_1, n9376, n9370, n9364, n9355, n8590, n8582}), .out(n14742), .config_in(config_chain[36581:36576]), .config_rst(config_rst)); 
buffer_wire buffer_14742 (.in(n14742), .out(n14742_0));
mux11 mux_9577 (.in({n14829_0, n11460_0, n11450_0/**/, n11410_1, n11400_1, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14743), .config_in(config_chain[36587:36582]), .config_rst(config_rst)); 
buffer_wire buffer_14743 (.in(n14743), .out(n14743_0));
mux11 mux_9578 (.in({n14684_0, n10426_0/**/, n10410_0, n10372_0, n10356_1, n9376, n9370, n9364, n9358, n8590, n8582}), .out(n14744), .config_in(config_chain[36593:36588]), .config_rst(config_rst)); 
buffer_wire buffer_14744 (.in(n14744), .out(n14744_0));
mux11 mux_9579 (.in({n14831_0, n11482_0/**/, n11472_0, n11434_0, n11424_0, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14745), .config_in(config_chain[36599:36594]), .config_rst(config_rst)); 
buffer_wire buffer_14745 (.in(n14745), .out(n14745_0));
mux11 mux_9580 (.in({n14692_0, n10432_0, n10394_0, n10378_0, n10362_1/**/, n9376, n9370, n9364, n9358, n8594, n8582}), .out(n14746), .config_in(config_chain[36605:36600]), .config_rst(config_rst)); 
buffer_wire buffer_14746 (.in(n14746), .out(n14746_0));
mux11 mux_9581 (.in({n14833_0, n11456_0, n11446_0/**/, n11416_1, n11406_1, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14747), .config_in(config_chain[36611:36606]), .config_rst(config_rst)); 
buffer_wire buffer_14747 (.in(n14747), .out(n14747_0));
mux10 mux_9582 (.in({n14700_0, n10416_0, n10400_0/**/, n10384_0, n10262_2, n9370, n9364, n9358, n8594, n8586}), .out(n14748), .config_in(config_chain[36617:36612]), .config_rst(config_rst)); 
buffer_wire buffer_14748 (.in(n14748), .out(n14748_0));
mux2 mux_9583 (.in({n12166_1/**/, n9652}), .out(n14749), .config_in(config_chain[36618:36618]), .config_rst(config_rst)); 
buffer_wire buffer_14749 (.in(n14749), .out(n14749_0));
mux12 mux_9584 (.in({n14614_0/**/, n10676_0, n10660_0, n10644_0, n10606_1, n10522_2, n9421, n9412, n9406, n8692, n8684, n8676}), .out(n14750), .config_in(config_chain[36624:36619]), .config_rst(config_rst)); 
buffer_wire buffer_14750 (.in(n14750), .out(n14750_0));
mux13 mux_9585 (.in({n14835_0, n11722_0/**/, n11712_0, n11674_1, n11664_1, n11596_2, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14751), .config_in(config_chain[36630:36625]), .config_rst(config_rst)); 
buffer_wire buffer_14751 (.in(n14751), .out(n14751_0));
mux12 mux_9586 (.in({n14622_0, n10682_0, n10666_0, n10628_0, n10612_1, n10524_2, n9421, n9415, n9406, n8692, n8684, n8676/**/}), .out(n14752), .config_in(config_chain[36636:36631]), .config_rst(config_rst)); 
buffer_wire buffer_14752 (.in(n14752), .out(n14752_0));
mux13 mux_9587 (.in({n14837_0, n11742_0/**/, n11732_0, n11696_0, n11686_0, n11618_2, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14753), .config_in(config_chain[36642:36637]), .config_rst(config_rst)); 
buffer_wire buffer_14753 (.in(n14753), .out(n14753_0));
mux11 mux_9588 (.in({n14630_0, n10688_0/**/, n10650_0, n10634_0, n10618_1, n9421, n9415, n9409, n8692, n8684, n8676}), .out(n14754), .config_in(config_chain[36648:36643]), .config_rst(config_rst)); 
buffer_wire buffer_14754 (.in(n14754), .out(n14754_0));
mux13 mux_9589 (.in({n14839_0, n11718_0, n11708_0/**/, n11680_1, n11670_1, n11640_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14755), .config_in(config_chain[36654:36649]), .config_rst(config_rst)); 
buffer_wire buffer_14755 (.in(n14755), .out(n14755_0));
mux11 mux_9590 (.in({n14638_0, n10672_0, n10656_0, n10640_0, n10624_1, n9421, n9415, n9409, n9403, n8684, n8676/**/}), .out(n14756), .config_in(config_chain[36660:36655]), .config_rst(config_rst)); 
buffer_wire buffer_14756 (.in(n14756), .out(n14756_0));
mux13 mux_9591 (.in({n14841_0, n11738_0, n11728_0, n11702_0/**/, n11692_0, n11662_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14757), .config_in(config_chain[36666:36661]), .config_rst(config_rst)); 
buffer_wire buffer_14757 (.in(n14757), .out(n14757_0));
mux11 mux_9592 (.in({n14646_0, n10678_0, n10662_0, n10646_0, n10608_1, n9421, n9415, n9409, n9403, n8688, n8676}), .out(n14758), .config_in(config_chain[36672:36667]), .config_rst(config_rst)); 
buffer_wire buffer_14758 (.in(n14758), .out(n14758_0));
mux13 mux_9593 (.in({n14843_0, n11724_0, n11714_0, n11684_1, n11676_1, n11666_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14759), .config_in(config_chain[36678:36673]), .config_rst(config_rst)); 
buffer_wire buffer_14759 (.in(n14759), .out(n14759_0));
mux11 mux_9594 (.in({n14654_0, n10684_0/**/, n10668_0, n10630_0, n10614_1, n9424, n9415, n9409, n9403, n8688, n8680}), .out(n14760), .config_in(config_chain[36684:36679]), .config_rst(config_rst)); 
buffer_wire buffer_14760 (.in(n14760), .out(n14760_0));
mux12 mux_9595 (.in({n14845_0, n11744_0/**/, n11734_0, n11706_0, n11698_0, n11688_0, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14761), .config_in(config_chain[36690:36685]), .config_rst(config_rst)); 
buffer_wire buffer_14761 (.in(n14761), .out(n14761_0));
mux11 mux_9596 (.in({n14662_0, n10690_0/**/, n10652_0, n10636_0, n10620_1, n9424, n9418, n9409, n9403, n8688, n8680}), .out(n14762), .config_in(config_chain[36696:36691]), .config_rst(config_rst)); 
buffer_wire buffer_14762 (.in(n14762), .out(n14762_0));
mux11 mux_9597 (.in({n14847_0, n11720_0, n11710_0, n11682_1/**/, n11672_1, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14763), .config_in(config_chain[36702:36697]), .config_rst(config_rst)); 
buffer_wire buffer_14763 (.in(n14763), .out(n14763_0));
mux11 mux_9598 (.in({n14670_0, n10674_0, n10658_0, n10642_0, n10626_1, n9424, n9418, n9412, n9403, n8688, n8680/**/}), .out(n14764), .config_in(config_chain[36708:36703]), .config_rst(config_rst)); 
buffer_wire buffer_14764 (.in(n14764), .out(n14764_0));
mux11 mux_9599 (.in({n14849_0, n11740_0, n11730_0, n11704_0, n11694_0, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14765), .config_in(config_chain[36714:36709]), .config_rst(config_rst)); 
buffer_wire buffer_14765 (.in(n14765), .out(n14765_0));
mux11 mux_9600 (.in({n14678_0, n10680_0/**/, n10664_0, n10648_0, n10610_1, n9424, n9418, n9412, n9406, n8688, n8680}), .out(n14766), .config_in(config_chain[36720:36715]), .config_rst(config_rst)); 
buffer_wire buffer_14766 (.in(n14766), .out(n14766_0));
mux11 mux_9601 (.in({n14851_0, n11726_0, n11716_0, n11678_1, n11668_1, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14767), .config_in(config_chain[36726:36721]), .config_rst(config_rst)); 
buffer_wire buffer_14767 (.in(n14767), .out(n14767_0));
mux11 mux_9602 (.in({n14686_0, n10686_0, n10670_0, n10632_0, n10616_1, n9424, n9418, n9412, n9406, n8692, n8680/**/}), .out(n14768), .config_in(config_chain[36732:36727]), .config_rst(config_rst)); 
buffer_wire buffer_14768 (.in(n14768), .out(n14768_0));
mux11 mux_9603 (.in({n14853_0, n11746_0, n11736_0/**/, n11700_0, n11690_0, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14769), .config_in(config_chain[36738:36733]), .config_rst(config_rst)); 
buffer_wire buffer_14769 (.in(n14769), .out(n14769_0));
mux10 mux_9604 (.in({n14702_0, n10692_0/**/, n10654_0, n10638_0, n10622_1, n9418, n9412, n9406, n8692, n8684}), .out(n14770), .config_in(config_chain[36744:36739]), .config_rst(config_rst)); 
buffer_wire buffer_14770 (.in(n14770), .out(n14770_0));
mux2 mux_9605 (.in({n12188_1, n9652}), .out(n14771), .config_in(config_chain[36745:36745]), .config_rst(config_rst)); 
buffer_wire buffer_14771 (.in(n14771), .out(n14771_0));
mux12 mux_9606 (.in({n14616_1, n10954_0, n10934_0, n10916_0, n10900_0, n10884_1, n9469, n9460, n9454, n8790, n8782, n8774/**/}), .out(n14772), .config_in(config_chain[36751:36746]), .config_rst(config_rst)); 
buffer_wire buffer_14772 (.in(n14772), .out(n14772_0));
mux13 mux_9607 (.in({n14855_0, n12000_0, n11990_0, n11964_0, n11954_0, n11828_2, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14773), .config_in(config_chain[36757:36752]), .config_rst(config_rst)); 
buffer_wire buffer_14773 (.in(n14773), .out(n14773_0));
mux12 mux_9608 (.in({n14624_1, n10940_0/**/, n10922_0, n10906_0, n10868_1, n10784_2, n9469, n9463, n9454, n8790, n8782, n8774}), .out(n14774), .config_in(config_chain[36763:36758]), .config_rst(config_rst)); 
buffer_wire buffer_14774 (.in(n14774), .out(n14774_0));
mux13 mux_9609 (.in({n14857_0, n11984_0, n11974_0/**/, n11938_1, n11928_1, n11860_2, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14775), .config_in(config_chain[36769:36764]), .config_rst(config_rst)); 
buffer_wire buffer_14775 (.in(n14775), .out(n14775_0));
mux11 mux_9610 (.in({n14632_1, n10946_0, n10928_0, n10890_0, n10874_1, n9469, n9463, n9457, n8790, n8782, n8774/**/}), .out(n14776), .config_in(config_chain[36775:36770]), .config_rst(config_rst)); 
buffer_wire buffer_14776 (.in(n14776), .out(n14776_0));
mux13 mux_9611 (.in({n14859_0, n12006_0, n11996_0, n11960_0, n11950_0/**/, n11882_2, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14777), .config_in(config_chain[36781:36776]), .config_rst(config_rst)); 
buffer_wire buffer_14777 (.in(n14777), .out(n14777_0));
mux11 mux_9612 (.in({n14640_1, n10952_0, n10912_0, n10896_0/**/, n10880_1, n9469, n9463, n9457, n9451, n8782, n8774}), .out(n14778), .config_in(config_chain[36787:36782]), .config_rst(config_rst)); 
buffer_wire buffer_14778 (.in(n14778), .out(n14778_0));
mux13 mux_9613 (.in({n14861_0, n11980_0/**/, n11970_0, n11944_1, n11934_1, n11904_1, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14779), .config_in(config_chain[36793:36788]), .config_rst(config_rst)); 
buffer_wire buffer_14779 (.in(n14779), .out(n14779_0));
mux11 mux_9614 (.in({n14648_1, n10936_0, n10918_0, n10902_0, n10886_1/**/, n9469, n9463, n9457, n9451, n8786, n8774}), .out(n14780), .config_in(config_chain[36799:36794]), .config_rst(config_rst)); 
buffer_wire buffer_14780 (.in(n14780), .out(n14780_0));
mux13 mux_9615 (.in({n14863_0, n12002_0/**/, n11992_0, n11966_0, n11956_0, n11926_1, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14781), .config_in(config_chain[36805:36800]), .config_rst(config_rst)); 
buffer_wire buffer_14781 (.in(n14781), .out(n14781_0));
mux11 mux_9616 (.in({n14656_1, n10942_0, n10924_0/**/, n10908_0, n10870_1, n9472, n9463, n9457, n9451, n8786, n8778}), .out(n14782), .config_in(config_chain[36811:36806]), .config_rst(config_rst)); 
buffer_wire buffer_14782 (.in(n14782), .out(n14782_0));
mux12 mux_9617 (.in({n14865_0, n11986_0, n11976_0, n11948_1, n11940_1, n11930_1, n9613, n9607, n9601, n9595, n9080/**/, n9072}), .out(n14783), .config_in(config_chain[36817:36812]), .config_rst(config_rst)); 
buffer_wire buffer_14783 (.in(n14783), .out(n14783_0));
mux11 mux_9618 (.in({n14664_1, n10948_0/**/, n10930_0, n10892_0, n10876_1, n9472, n9466, n9457, n9451, n8786, n8778}), .out(n14784), .config_in(config_chain[36823:36818]), .config_rst(config_rst)); 
buffer_wire buffer_14784 (.in(n14784), .out(n14784_0));
mux11 mux_9619 (.in({n14867_0, n12008_0, n11998_0/**/, n11962_0, n11952_0, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14785), .config_in(config_chain[36829:36824]), .config_rst(config_rst)); 
buffer_wire buffer_14785 (.in(n14785), .out(n14785_0));
mux11 mux_9620 (.in({n14672_1, n10914_0, n10898_0, n10882_1, n10866_1, n9472, n9466/**/, n9460, n9451, n8786, n8778}), .out(n14786), .config_in(config_chain[36835:36830]), .config_rst(config_rst)); 
buffer_wire buffer_14786 (.in(n14786), .out(n14786_0));
mux11 mux_9621 (.in({n14869_0, n11982_0, n11972_0, n11946_1, n11936_1, n9613, n9607, n9601, n9595, n9080, n9072/**/}), .out(n14787), .config_in(config_chain[36841:36836]), .config_rst(config_rst)); 
buffer_wire buffer_14787 (.in(n14787), .out(n14787_0));
mux11 mux_9622 (.in({n14680_1, n10938_0, n10920_0, n10904_0, n10888_1, n9472, n9466/**/, n9460, n9454, n8786, n8778}), .out(n14788), .config_in(config_chain[36847:36842]), .config_rst(config_rst)); 
buffer_wire buffer_14788 (.in(n14788), .out(n14788_0));
mux11 mux_9623 (.in({n14871_0, n12004_0, n11994_0, n11968_0, n11958_0/**/, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14789), .config_in(config_chain[36853:36848]), .config_rst(config_rst)); 
buffer_wire buffer_14789 (.in(n14789), .out(n14789_0));
mux11 mux_9624 (.in({n14688_1, n10944_0, n10926_0, n10910_0, n10872_1, n9472, n9466/**/, n9460, n9454, n8790, n8778}), .out(n14790), .config_in(config_chain[36859:36854]), .config_rst(config_rst)); 
buffer_wire buffer_14790 (.in(n14790), .out(n14790_0));
mux11 mux_9625 (.in({n14873_0, n11988_0, n11978_0, n11942_1, n11932_1, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14791), .config_in(config_chain[36865:36860]), .config_rst(config_rst)); 
buffer_wire buffer_14791 (.in(n14791), .out(n14791_0));
mux10 mux_9626 (.in({n14704_1, n10950_0, n10932_0, n10894_0, n10878_1, n9466/**/, n9460, n9454, n8790, n8782}), .out(n14792), .config_in(config_chain[36871:36866]), .config_rst(config_rst)); 
buffer_wire buffer_14792 (.in(n14792), .out(n14792_0));
mux2 mux_9627 (.in({n12230_0/**/, n9655}), .out(n14793), .config_in(config_chain[36872:36872]), .config_rst(config_rst)); 
buffer_wire buffer_14793 (.in(n14793), .out(n14793_0));
mux13 mux_9628 (.in({n14706_1/**/, n11186_0, n11176_0, n11146_1, n11136_1, n11108_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14794), .config_in(config_chain[36878:36873]), .config_rst(config_rst)); 
buffer_wire buffer_14794 (.in(n14794), .out(n14794_0));
mux3 mux_9629 (.in({n12210_0, n9655, n9166}), .out(n14795), .config_in(config_chain[36880:36879]), .config_rst(config_rst)); 
buffer_wire buffer_14795 (.in(n14795), .out(n14795_0));
mux13 mux_9630 (.in({n14708_1, n11208_0, n11198_0, n11168_0/**/, n11158_0, n11130_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14796), .config_in(config_chain[36886:36881]), .config_rst(config_rst)); 
buffer_wire buffer_14796 (.in(n14796), .out(n14796_0));
mux3 mux_9631 (.in({n12212_0/**/, n9658, n9170}), .out(n14797), .config_in(config_chain[36888:36887]), .config_rst(config_rst)); 
buffer_wire buffer_14797 (.in(n14797), .out(n14797_0));
mux13 mux_9632 (.in({n14710_1/**/, n11192_0, n11182_0, n11152_1, n11142_1, n11132_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14798), .config_in(config_chain[36894:36889]), .config_rst(config_rst)); 
buffer_wire buffer_14798 (.in(n14798), .out(n14798_0));
mux3 mux_9633 (.in({n12214_0/**/, n9661, n9174}), .out(n14799), .config_in(config_chain[36896:36895]), .config_rst(config_rst)); 
buffer_wire buffer_14799 (.in(n14799), .out(n14799_0));
mux13 mux_9634 (.in({n14712_1, n11214_0, n11204_0, n11174_0, n11164_0, n11154_0, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14800), .config_in(config_chain[36902:36897]), .config_rst(config_rst)); 
buffer_wire buffer_14800 (.in(n14800), .out(n14800_0));
mux3 mux_9635 (.in({n12216_0, n9664, n9174}), .out(n14801), .config_in(config_chain[36904:36903]), .config_rst(config_rst)); 
buffer_wire buffer_14801 (.in(n14801), .out(n14801_0));
mux13 mux_9636 (.in({n14714_1, n11196_0, n11188_0, n11178_0, n11148_1, n11138_1, n9520, n9514, n9508, n9502, n8888, n8880, n8872}), .out(n14802), .config_in(config_chain[36910:36905]), .config_rst(config_rst)); 
buffer_wire buffer_14802 (.in(n14802), .out(n14802_0));
mux3 mux_9637 (.in({n12218_0, n9664, n9178}), .out(n14803), .config_in(config_chain[36912:36911]), .config_rst(config_rst)); 
buffer_wire buffer_14803 (.in(n14803), .out(n14803_0));
mux12 mux_9638 (.in({n14716_1/**/, n11218_0, n11210_0, n11200_0, n11170_0, n11160_0, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14804), .config_in(config_chain[36918:36913]), .config_rst(config_rst)); 
buffer_wire buffer_14804 (.in(n14804), .out(n14804_0));
mux2 mux_9639 (.in({n12220_0, n9182}), .out(n14805), .config_in(config_chain[36919:36919]), .config_rst(config_rst)); 
buffer_wire buffer_14805 (.in(n14805), .out(n14805_0));
mux11 mux_9640 (.in({n14718_1, n11194_0, n11184_0, n11144_1, n11134_1/**/, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14806), .config_in(config_chain[36925:36920]), .config_rst(config_rst)); 
buffer_wire buffer_14806 (.in(n14806), .out(n14806_0));
mux2 mux_9641 (.in({n12222_0/**/, n9643}), .out(n14807), .config_in(config_chain[36926:36926]), .config_rst(config_rst)); 
buffer_wire buffer_14807 (.in(n14807), .out(n14807_0));
mux11 mux_9642 (.in({n14720_1/**/, n11216_0, n11206_0, n11166_0, n11156_0, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14808), .config_in(config_chain[36932:36927]), .config_rst(config_rst)); 
buffer_wire buffer_14808 (.in(n14808), .out(n14808_0));
mux2 mux_9643 (.in({n12224_0, n9646}), .out(n14809), .config_in(config_chain[36933:36933]), .config_rst(config_rst)); 
buffer_wire buffer_14809 (.in(n14809), .out(n14809_0));
mux11 mux_9644 (.in({n14722_1/**/, n11190_0, n11180_0, n11150_1, n11140_1, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14810), .config_in(config_chain[36939:36934]), .config_rst(config_rst)); 
buffer_wire buffer_14810 (.in(n14810), .out(n14810_0));
mux2 mux_9645 (.in({n12226_0, n9646}), .out(n14811), .config_in(config_chain[36940:36940]), .config_rst(config_rst)); 
buffer_wire buffer_14811 (.in(n14811), .out(n14811_0));
mux11 mux_9646 (.in({n14724_1, n11212_0/**/, n11202_0, n11172_0, n11162_0, n9517, n9511, n9505, n9499, n8884, n8876}), .out(n14812), .config_in(config_chain[36946:36941]), .config_rst(config_rst)); 
buffer_wire buffer_14812 (.in(n14812), .out(n14812_0));
mux2 mux_9647 (.in({n12228_0/**/, n9649}), .out(n14813), .config_in(config_chain[36947:36947]), .config_rst(config_rst)); 
buffer_wire buffer_14813 (.in(n14813), .out(n14813_0));
mux13 mux_9648 (.in({n14728_1/**/, n11478_0, n11468_0, n11430_0, n11420_0, n11352_2, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14814), .config_in(config_chain[36953:36948]), .config_rst(config_rst)); 
buffer_wire buffer_14814 (.in(n14814), .out(n14814_0));
mux3 mux_9649 (.in({n12232_0, n9655, n9166}), .out(n14815), .config_in(config_chain[36955:36954]), .config_rst(config_rst)); 
buffer_wire buffer_14815 (.in(n14815), .out(n14815_0));
mux13 mux_9650 (.in({n14730_1, n11452_0, n11442_0, n11412_1/**/, n11402_1, n11374_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14816), .config_in(config_chain[36961:36956]), .config_rst(config_rst)); 
buffer_wire buffer_14816 (.in(n14816), .out(n14816_0));
mux3 mux_9651 (.in({n12234_0, n9658, n9170}), .out(n14817), .config_in(config_chain[36963:36962]), .config_rst(config_rst)); 
buffer_wire buffer_14817 (.in(n14817), .out(n14817_0));
mux13 mux_9652 (.in({n14732_1, n11474_0/**/, n11464_0, n11436_0, n11426_0, n11396_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14818), .config_in(config_chain[36969:36964]), .config_rst(config_rst)); 
buffer_wire buffer_14818 (.in(n14818), .out(n14818_0));
mux3 mux_9653 (.in({n12236_0, n9661, n9174}), .out(n14819), .config_in(config_chain[36971:36970]), .config_rst(config_rst)); 
buffer_wire buffer_14819 (.in(n14819), .out(n14819_0));
mux13 mux_9654 (.in({n14734_1, n11458_0, n11448_0/**/, n11418_1, n11408_1, n11398_1, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14820), .config_in(config_chain[36977:36972]), .config_rst(config_rst)); 
buffer_wire buffer_14820 (.in(n14820), .out(n14820_0));
mux3 mux_9655 (.in({n12238_0, n9664, n9178}), .out(n14821), .config_in(config_chain[36979:36978]), .config_rst(config_rst)); 
buffer_wire buffer_14821 (.in(n14821), .out(n14821_0));
mux13 mux_9656 (.in({n14736_1, n11480_0, n11470_0, n11440_0, n11432_0, n11422_0, n9568, n9562, n9556, n9550, n8986, n8978, n8970}), .out(n14822), .config_in(config_chain[36985:36980]), .config_rst(config_rst)); 
buffer_wire buffer_14822 (.in(n14822), .out(n14822_0));
mux2 mux_9657 (.in({n12240_0/**/, n9178}), .out(n14823), .config_in(config_chain[36986:36986]), .config_rst(config_rst)); 
buffer_wire buffer_14823 (.in(n14823), .out(n14823_0));
mux12 mux_9658 (.in({n14738_1, n11462_0, n11454_0, n11444_0, n11414_1, n11404_1, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14824), .config_in(config_chain[36992:36987]), .config_rst(config_rst)); 
buffer_wire buffer_14824 (.in(n14824), .out(n14824_0));
mux2 mux_9659 (.in({n12242_0, n9182}), .out(n14825), .config_in(config_chain[36993:36993]), .config_rst(config_rst)); 
buffer_wire buffer_14825 (.in(n14825), .out(n14825_0));
mux11 mux_9660 (.in({n14740_1, n11476_0, n11466_0, n11438_0, n11428_0/**/, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14826), .config_in(config_chain[36999:36994]), .config_rst(config_rst)); 
buffer_wire buffer_14826 (.in(n14826), .out(n14826_0));
mux2 mux_9661 (.in({n12244_0/**/, n9643}), .out(n14827), .config_in(config_chain[37000:37000]), .config_rst(config_rst)); 
buffer_wire buffer_14827 (.in(n14827), .out(n14827_0));
mux11 mux_9662 (.in({n14742_1, n11460_0/**/, n11450_0, n11410_1, n11400_1, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14828), .config_in(config_chain[37006:37001]), .config_rst(config_rst)); 
buffer_wire buffer_14828 (.in(n14828), .out(n14828_0));
mux2 mux_9663 (.in({n12246_0, n9646}), .out(n14829), .config_in(config_chain[37007:37007]), .config_rst(config_rst)); 
buffer_wire buffer_14829 (.in(n14829), .out(n14829_0));
mux11 mux_9664 (.in({n14744_1, n11482_0, n11472_0/**/, n11434_0, n11424_0, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14830), .config_in(config_chain[37013:37008]), .config_rst(config_rst)); 
buffer_wire buffer_14830 (.in(n14830), .out(n14830_0));
mux2 mux_9665 (.in({n12248_0, n9649}), .out(n14831), .config_in(config_chain[37014:37014]), .config_rst(config_rst)); 
buffer_wire buffer_14831 (.in(n14831), .out(n14831_0));
mux11 mux_9666 (.in({n14746_1, n11456_0, n11446_0, n11416_1, n11406_1/**/, n9565, n9559, n9553, n9547, n8982, n8974}), .out(n14832), .config_in(config_chain[37020:37015]), .config_rst(config_rst)); 
buffer_wire buffer_14832 (.in(n14832), .out(n14832_0));
mux2 mux_9667 (.in({n12090_2, n9649}), .out(n14833), .config_in(config_chain[37021:37021]), .config_rst(config_rst)); 
buffer_wire buffer_14833 (.in(n14833), .out(n14833_0));
mux13 mux_9668 (.in({n14750_1, n11722_0, n11712_0, n11674_1/**/, n11664_1, n11596_2, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14834), .config_in(config_chain[37027:37022]), .config_rst(config_rst)); 
buffer_wire buffer_14834 (.in(n14834), .out(n14834_0));
mux3 mux_9669 (.in({n12250_0, n9655, n9166}), .out(n14835), .config_in(config_chain[37029:37028]), .config_rst(config_rst)); 
buffer_wire buffer_14835 (.in(n14835), .out(n14835_0));
mux13 mux_9670 (.in({n14752_1, n11742_0, n11732_0, n11696_0, n11686_0, n11618_2, n9616, n9610, n9604, n9598, n9084, n9076, n9068/**/}), .out(n14836), .config_in(config_chain[37035:37030]), .config_rst(config_rst)); 
buffer_wire buffer_14836 (.in(n14836), .out(n14836_0));
mux3 mux_9671 (.in({n12252_0, n9658, n9166}), .out(n14837), .config_in(config_chain[37037:37036]), .config_rst(config_rst)); 
buffer_wire buffer_14837 (.in(n14837), .out(n14837_0));
mux13 mux_9672 (.in({n14754_1, n11718_0, n11708_0, n11680_1/**/, n11670_1, n11640_1, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14838), .config_in(config_chain[37043:37038]), .config_rst(config_rst)); 
buffer_wire buffer_14838 (.in(n14838), .out(n14838_0));
mux3 mux_9673 (.in({n12254_0, n9658, n9170}), .out(n14839), .config_in(config_chain[37045:37044]), .config_rst(config_rst)); 
buffer_wire buffer_14839 (.in(n14839), .out(n14839_0));
mux13 mux_9674 (.in({n14756_1, n11738_0, n11728_0, n11702_0, n11692_0, n11662_1, n9616, n9610, n9604, n9598, n9084, n9076, n9068}), .out(n14840), .config_in(config_chain[37051:37046]), .config_rst(config_rst)); 
buffer_wire buffer_14840 (.in(n14840), .out(n14840_0));
mux3 mux_9675 (.in({n12256_0/**/, n9661, n9174}), .out(n14841), .config_in(config_chain[37053:37052]), .config_rst(config_rst)); 
buffer_wire buffer_14841 (.in(n14841), .out(n14841_0));
mux13 mux_9676 (.in({n14758_1, n11724_0, n11714_0, n11684_1, n11676_1, n11666_1, n9616, n9610, n9604, n9598, n9084/**/, n9076, n9068}), .out(n14842), .config_in(config_chain[37059:37054]), .config_rst(config_rst)); 
buffer_wire buffer_14842 (.in(n14842), .out(n14842_0));
mux3 mux_9677 (.in({n12258_0, n9664, n9178}), .out(n14843), .config_in(config_chain[37061:37060]), .config_rst(config_rst)); 
buffer_wire buffer_14843 (.in(n14843), .out(n14843_0));
mux12 mux_9678 (.in({n14760_1, n11744_0, n11734_0, n11706_0, n11698_0, n11688_0, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14844), .config_in(config_chain[37067:37062]), .config_rst(config_rst)); 
buffer_wire buffer_14844 (.in(n14844), .out(n14844_0));
mux2 mux_9679 (.in({n12260_0/**/, n9182}), .out(n14845), .config_in(config_chain[37068:37068]), .config_rst(config_rst)); 
buffer_wire buffer_14845 (.in(n14845), .out(n14845_0));
mux11 mux_9680 (.in({n14762_1/**/, n11720_0, n11710_0, n11682_1, n11672_1, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14846), .config_in(config_chain[37074:37069]), .config_rst(config_rst)); 
buffer_wire buffer_14846 (.in(n14846), .out(n14846_0));
mux2 mux_9681 (.in({n12262_0, n9182}), .out(n14847), .config_in(config_chain[37075:37075]), .config_rst(config_rst)); 
buffer_wire buffer_14847 (.in(n14847), .out(n14847_0));
mux11 mux_9682 (.in({n14764_1, n11740_0, n11730_0, n11704_0, n11694_0, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14848), .config_in(config_chain[37081:37076]), .config_rst(config_rst)); 
buffer_wire buffer_14848 (.in(n14848), .out(n14848_0));
mux2 mux_9683 (.in({n12264_0/**/, n9643}), .out(n14849), .config_in(config_chain[37082:37082]), .config_rst(config_rst)); 
buffer_wire buffer_14849 (.in(n14849), .out(n14849_0));
mux11 mux_9684 (.in({n14766_1, n11726_0, n11716_0, n11678_1, n11668_1, n9613, n9607, n9601, n9595, n9080, n9072/**/}), .out(n14850), .config_in(config_chain[37088:37083]), .config_rst(config_rst)); 
buffer_wire buffer_14850 (.in(n14850), .out(n14850_0));
mux2 mux_9685 (.in({n12266_0, n9646}), .out(n14851), .config_in(config_chain[37089:37089]), .config_rst(config_rst)); 
buffer_wire buffer_14851 (.in(n14851), .out(n14851_0));
mux11 mux_9686 (.in({n14768_1, n11746_0, n11736_0, n11700_0, n11690_0, n9613, n9607, n9601, n9595, n9080, n9072}), .out(n14852), .config_in(config_chain[37095:37090]), .config_rst(config_rst)); 
buffer_wire buffer_14852 (.in(n14852), .out(n14852_0));
mux2 mux_9687 (.in({n12268_0/**/, n9649}), .out(n14853), .config_in(config_chain[37096:37096]), .config_rst(config_rst)); 
buffer_wire buffer_14853 (.in(n14853), .out(n14853_0));
mux13 mux_9688 (.in({n14772_1, n12000_0/**/, n11990_0, n11964_0, n11954_0, n11828_2, n9664, n9658, n9652, n9646, n9182, n9174, n9166}), .out(n14854), .config_in(config_chain[37102:37097]), .config_rst(config_rst)); 
buffer_wire buffer_14854 (.in(n14854), .out(n14854_0));
mux3 mux_9689 (.in({n12190_1, n9655, n9166}), .out(n14855), .config_in(config_chain[37104:37103]), .config_rst(config_rst)); 
buffer_wire buffer_14855 (.in(n14855), .out(n14855_0));
mux13 mux_9690 (.in({n14774_1, n11984_0/**/, n11974_0, n11938_1, n11928_1, n11860_2, n9664, n9658, n9652, n9646, n9182, n9174, n9166}), .out(n14856), .config_in(config_chain[37110:37105]), .config_rst(config_rst)); 
buffer_wire buffer_14856 (.in(n14856), .out(n14856_0));
mux3 mux_9691 (.in({n12192_1, n9658, n9170}), .out(n14857), .config_in(config_chain[37112:37111]), .config_rst(config_rst)); 
buffer_wire buffer_14857 (.in(n14857), .out(n14857_0));
mux13 mux_9692 (.in({n14776_1, n12006_0/**/, n11996_0, n11960_0, n11950_0, n11882_2, n9664, n9658, n9652, n9646, n9182, n9174, n9166}), .out(n14858), .config_in(config_chain[37118:37113]), .config_rst(config_rst)); 
buffer_wire buffer_14858 (.in(n14858), .out(n14858_0));
mux3 mux_9693 (.in({n12194_1, n9661, n9170}), .out(n14859), .config_in(config_chain[37120:37119]), .config_rst(config_rst)); 
buffer_wire buffer_14859 (.in(n14859), .out(n14859_0));
mux13 mux_9694 (.in({n14778_1, n11980_0, n11970_0/**/, n11944_1, n11934_1, n11904_1, n9664, n9658, n9652, n9646, n9182, n9174, n9166}), .out(n14860), .config_in(config_chain[37126:37121]), .config_rst(config_rst)); 
buffer_wire buffer_14860 (.in(n14860), .out(n14860_0));
mux3 mux_9695 (.in({n12196_1, n9661, n9174}), .out(n14861), .config_in(config_chain[37128:37127]), .config_rst(config_rst)); 
buffer_wire buffer_14861 (.in(n14861), .out(n14861_0));
mux13 mux_9696 (.in({n14780_1, n12002_0, n11992_0, n11966_0, n11956_0, n11926_1, n9664, n9658, n9652, n9646, n9182, n9174, n9166}), .out(n14862), .config_in(config_chain[37134:37129]), .config_rst(config_rst)); 
buffer_wire buffer_14862 (.in(n14862), .out(n14862_0));
mux3 mux_9697 (.in({n12198_1/**/, n9664, n9178}), .out(n14863), .config_in(config_chain[37136:37135]), .config_rst(config_rst)); 
buffer_wire buffer_14863 (.in(n14863), .out(n14863_0));
mux12 mux_9698 (.in({n14782_1, n11986_0, n11976_0, n11948_1, n11940_1, n11930_1/**/, n9661, n9655, n9649, n9643, n9178, n9170}), .out(n14864), .config_in(config_chain[37142:37137]), .config_rst(config_rst)); 
buffer_wire buffer_14864 (.in(n14864), .out(n14864_0));
mux2 mux_9699 (.in({n12200_1, n9182}), .out(n14865), .config_in(config_chain[37143:37143]), .config_rst(config_rst)); 
buffer_wire buffer_14865 (.in(n14865), .out(n14865_0));
mux11 mux_9700 (.in({n14784_1, n12008_0/**/, n11998_0, n11962_0, n11952_0, n9661, n9655, n9649, n9643, n9178, n9170}), .out(n14866), .config_in(config_chain[37149:37144]), .config_rst(config_rst)); 
buffer_wire buffer_14866 (.in(n14866), .out(n14866_0));
mux2 mux_9701 (.in({n12202_1, n9643}), .out(n14867), .config_in(config_chain[37150:37150]), .config_rst(config_rst)); 
buffer_wire buffer_14867 (.in(n14867), .out(n14867_0));
mux11 mux_9702 (.in({n14786_1/**/, n11982_0, n11972_0, n11946_1, n11936_1, n9661, n9655, n9649, n9643, n9178, n9170}), .out(n14868), .config_in(config_chain[37156:37151]), .config_rst(config_rst)); 
buffer_wire buffer_14868 (.in(n14868), .out(n14868_0));
mux2 mux_9703 (.in({n12204_1, n9643}), .out(n14869), .config_in(config_chain[37157:37157]), .config_rst(config_rst)); 
buffer_wire buffer_14869 (.in(n14869), .out(n14869_0));
mux11 mux_9704 (.in({n14788_1, n12004_0, n11994_0/**/, n11968_0, n11958_0, n9661, n9655, n9649, n9643, n9178, n9170}), .out(n14870), .config_in(config_chain[37163:37158]), .config_rst(config_rst)); 
buffer_wire buffer_14870 (.in(n14870), .out(n14870_0));
mux2 mux_9705 (.in({n12206_1, n9646}), .out(n14871), .config_in(config_chain[37164:37164]), .config_rst(config_rst)); 
buffer_wire buffer_14871 (.in(n14871), .out(n14871_0));
mux11 mux_9706 (.in({n14790_1/**/, n11988_0, n11978_0, n11942_1, n11932_1, n9661, n9655, n9649, n9643, n9178, n9170}), .out(n14872), .config_in(config_chain[37170:37165]), .config_rst(config_rst)); 
buffer_wire buffer_14872 (.in(n14872), .out(n14872_0));
mux2 mux_9707 (.in({n12208_1, n9649}), .out(n14873), .config_in(config_chain[37171:37171]), .config_rst(config_rst)); 
buffer_wire buffer_14873 (.in(n14873), .out(n14873_0));

wire [7:0]outpad_0_1;
assign outpad_0_1 = {n45, n42, n39, n36, n33, n30, n27, n24};
wire [7:0]inpad_0_1;
assign {n46, n43, n40, n37, n34, n31, n28, n25} = inpad_0_1;

io io_0_1 ( .outpad(outpad_0_1), .inpad(inpad_0_1), .io_ext(io_0_1_wire), .config_in(config_chain[37179:37172]), .config_rst(config_rst) );

wire [7:0]outpad_0_2;
assign outpad_0_2 = {n93, n90, n87, n84, n81, n78, n75, n72};
wire [7:0]inpad_0_2;
assign {n94, n91, n88, n85, n82, n79, n76, n73} = inpad_0_2;

io io_0_2 ( .outpad(outpad_0_2), .inpad(inpad_0_2), .io_ext(io_0_2_wire), .config_in(config_chain[37187:37180]), .config_rst(config_rst) );

wire [7:0]outpad_0_3;
assign outpad_0_3 = {n141, n138, n135, n132, n129, n126, n123, n120};
wire [7:0]inpad_0_3;
assign {n142, n139, n136, n133, n130, n127, n124, n121} = inpad_0_3;

io io_0_3 ( .outpad(outpad_0_3), .inpad(inpad_0_3), .io_ext(io_0_3_wire), .config_in(config_chain[37195:37188]), .config_rst(config_rst) );

wire [7:0]outpad_0_4;
assign outpad_0_4 = {n189, n186, n183, n180, n177, n174, n171, n168};
wire [7:0]inpad_0_4;
assign {n190, n187, n184, n181, n178, n175, n172, n169} = inpad_0_4;

io io_0_4 ( .outpad(outpad_0_4), .inpad(inpad_0_4), .io_ext(io_0_4_wire), .config_in(config_chain[37203:37196]), .config_rst(config_rst) );

wire [7:0]outpad_0_5;
assign outpad_0_5 = {n237, n234, n231, n228, n225, n222, n219, n216};
wire [7:0]inpad_0_5;
assign {n238, n235, n232, n229, n226, n223, n220, n217} = inpad_0_5;

io io_0_5 ( .outpad(outpad_0_5), .inpad(inpad_0_5), .io_ext(io_0_5_wire), .config_in(config_chain[37211:37204]), .config_rst(config_rst) );

wire [7:0]outpad_0_6;
assign outpad_0_6 = {n285, n282, n279, n276, n273, n270, n267, n264};
wire [7:0]inpad_0_6;
assign {n286, n283, n280, n277, n274, n271, n268, n265} = inpad_0_6;

io io_0_6 ( .outpad(outpad_0_6), .inpad(inpad_0_6), .io_ext(io_0_6_wire), .config_in(config_chain[37219:37212]), .config_rst(config_rst) );

wire [7:0]outpad_0_7;
assign outpad_0_7 = {n333, n330, n327, n324, n321, n318, n315, n312};
wire [7:0]inpad_0_7;
assign {n334, n331, n328, n325, n322, n319, n316, n313} = inpad_0_7;

io io_0_7 ( .outpad(outpad_0_7), .inpad(inpad_0_7), .io_ext(io_0_7_wire), .config_in(config_chain[37227:37220]), .config_rst(config_rst) );

wire [7:0]outpad_0_8;
assign outpad_0_8 = {n381, n378, n375, n372, n369, n366, n363, n360};
wire [7:0]inpad_0_8;
assign {n382, n379, n376, n373, n370, n367, n364, n361} = inpad_0_8;

io io_0_8 ( .outpad(outpad_0_8), .inpad(inpad_0_8), .io_ext(io_0_8_wire), .config_in(config_chain[37235:37228]), .config_rst(config_rst) );

wire [7:0]outpad_0_9;
assign outpad_0_9 = {n429, n426, n423, n420, n417, n414, n411, n408};
wire [7:0]inpad_0_9;
assign {n430, n427, n424, n421, n418, n415, n412, n409} = inpad_0_9;

io io_0_9 ( .outpad(outpad_0_9), .inpad(inpad_0_9), .io_ext(io_0_9_wire), .config_in(config_chain[37243:37236]), .config_rst(config_rst) );

wire [7:0]outpad_1_0;
assign outpad_1_0 = {n477, n474, n471, n468, n465, n462, n459, n456};
wire [7:0]inpad_1_0;
assign {n478, n475, n472, n469, n466, n463, n460, n457} = inpad_1_0;

io io_1_0 ( .outpad(outpad_1_0), .inpad(inpad_1_0), .io_ext(io_1_0_wire), .config_in(config_chain[37251:37244]), .config_rst(config_rst) );

wire [0:0]clk_1_1;
assign clk_1_1 = {fpga_clk};
wire [12:0]I1_1_1;
assign I1_1_1 = {n517, n516, n515, n514, n513, n512, n511, n510, n509, n508, n507, n506, n505};
wire [12:0]I2_1_1;
assign I2_1_1 = {n530, n529, n528, n527, n526, n525, n524, n523, n522, n521, n520, n519, n518};
wire [12:0]I3_1_1;
assign I3_1_1 = {n543, n542, n541, n540, n539, n538, n537, n536, n535, n534, n533, n532, n531};
wire [12:0]I4_1_1;
assign I4_1_1 = {n556, n555, n554, n553, n552, n551, n550, n549, n548, n547, n546, n545, n544};
wire [19:0]O_1_1;
assign {n576, n575, n574, n573, n572, n571, n570, n569, n568, n567, n566, n565, n564, n563, n562, n561, n560, n559, n558, n557} = O_1_1;

clb clb_1_1 ( .clk(clk_1_1), .reset(fpga_rst), .I4(I4_1_1), .I3(I3_1_1), .I2(I2_1_1), .I1(I1_1_1), .O(O_1_1), .config_in(config_chain[39211:37252]), .config_rst(config_rst) );

wire [0:0]clk_1_2;
assign clk_1_2 = {fpga_clk};
wire [12:0]I1_1_2;
assign I1_1_2 = {n615, n614, n613, n612, n611, n610, n609, n608, n607, n606, n605, n604, n603};
wire [12:0]I2_1_2;
assign I2_1_2 = {n628, n627, n626, n625, n624, n623, n622, n621, n620, n619, n618, n617, n616};
wire [12:0]I3_1_2;
assign I3_1_2 = {n641, n640, n639, n638, n637, n636, n635, n634, n633, n632, n631, n630, n629};
wire [12:0]I4_1_2;
assign I4_1_2 = {n654, n653, n652, n651, n650, n649, n648, n647, n646, n645, n644, n643, n642};
wire [19:0]O_1_2;
assign {n674, n673, n672, n671, n670, n669, n668, n667, n666, n665, n664, n663, n662, n661, n660, n659, n658, n657, n656, n655} = O_1_2;

clb clb_1_2 ( .clk(clk_1_2), .reset(fpga_rst), .I4(I4_1_2), .I3(I3_1_2), .I2(I2_1_2), .I1(I1_1_2), .O(O_1_2), .config_in(config_chain[41171:39212]), .config_rst(config_rst) );

wire [0:0]clk_1_3;
assign clk_1_3 = {fpga_clk};
wire [12:0]I1_1_3;
assign I1_1_3 = {n713, n712, n711, n710, n709, n708, n707, n706, n705, n704, n703, n702, n701};
wire [12:0]I2_1_3;
assign I2_1_3 = {n726, n725, n724, n723, n722, n721, n720, n719, n718, n717, n716, n715, n714};
wire [12:0]I3_1_3;
assign I3_1_3 = {n739, n738, n737, n736, n735, n734, n733, n732, n731, n730, n729, n728, n727};
wire [12:0]I4_1_3;
assign I4_1_3 = {n752, n751, n750, n749, n748, n747, n746, n745, n744, n743, n742, n741, n740};
wire [19:0]O_1_3;
assign {n772, n771, n770, n769, n768, n767, n766, n765, n764, n763, n762, n761, n760, n759, n758, n757, n756, n755, n754, n753} = O_1_3;

clb clb_1_3 ( .clk(clk_1_3), .reset(fpga_rst), .I4(I4_1_3), .I3(I3_1_3), .I2(I2_1_3), .I1(I1_1_3), .O(O_1_3), .config_in(config_chain[43131:41172]), .config_rst(config_rst) );

wire [0:0]clk_1_4;
assign clk_1_4 = {fpga_clk};
wire [12:0]I1_1_4;
assign I1_1_4 = {n811, n810, n809, n808, n807, n806, n805, n804, n803, n802, n801, n800, n799};
wire [12:0]I2_1_4;
assign I2_1_4 = {n824, n823, n822, n821, n820, n819, n818, n817, n816, n815, n814, n813, n812};
wire [12:0]I3_1_4;
assign I3_1_4 = {n837, n836, n835, n834, n833, n832, n831, n830, n829, n828, n827, n826, n825};
wire [12:0]I4_1_4;
assign I4_1_4 = {n850, n849, n848, n847, n846, n845, n844, n843, n842, n841, n840, n839, n838};
wire [19:0]O_1_4;
assign {n870, n869, n868, n867, n866, n865, n864, n863, n862, n861, n860, n859, n858, n857, n856, n855, n854, n853, n852, n851} = O_1_4;

clb clb_1_4 ( .clk(clk_1_4), .reset(fpga_rst), .I4(I4_1_4), .I3(I3_1_4), .I2(I2_1_4), .I1(I1_1_4), .O(O_1_4), .config_in(config_chain[45091:43132]), .config_rst(config_rst) );

wire [0:0]clk_1_5;
assign clk_1_5 = {fpga_clk};
wire [12:0]I1_1_5;
assign I1_1_5 = {n909, n908, n907, n906, n905, n904, n903, n902, n901, n900, n899, n898, n897};
wire [12:0]I2_1_5;
assign I2_1_5 = {n922, n921, n920, n919, n918, n917, n916, n915, n914, n913, n912, n911, n910};
wire [12:0]I3_1_5;
assign I3_1_5 = {n935, n934, n933, n932, n931, n930, n929, n928, n927, n926, n925, n924, n923};
wire [12:0]I4_1_5;
assign I4_1_5 = {n948, n947, n946, n945, n944, n943, n942, n941, n940, n939, n938, n937, n936};
wire [19:0]O_1_5;
assign {n968, n967, n966, n965, n964, n963, n962, n961, n960, n959, n958, n957, n956, n955, n954, n953, n952, n951, n950, n949} = O_1_5;

clb clb_1_5 ( .clk(clk_1_5), .reset(fpga_rst), .I4(I4_1_5), .I3(I3_1_5), .I2(I2_1_5), .I1(I1_1_5), .O(O_1_5), .config_in(config_chain[47051:45092]), .config_rst(config_rst) );

wire [0:0]clk_1_6;
assign clk_1_6 = {fpga_clk};
wire [12:0]I1_1_6;
assign I1_1_6 = {n1007, n1006, n1005, n1004, n1003, n1002, n1001, n1000, n999, n998, n997, n996, n995};
wire [12:0]I2_1_6;
assign I2_1_6 = {n1020, n1019, n1018, n1017, n1016, n1015, n1014, n1013, n1012, n1011, n1010, n1009, n1008};
wire [12:0]I3_1_6;
assign I3_1_6 = {n1033, n1032, n1031, n1030, n1029, n1028, n1027, n1026, n1025, n1024, n1023, n1022, n1021};
wire [12:0]I4_1_6;
assign I4_1_6 = {n1046, n1045, n1044, n1043, n1042, n1041, n1040, n1039, n1038, n1037, n1036, n1035, n1034};
wire [19:0]O_1_6;
assign {n1066, n1065, n1064, n1063, n1062, n1061, n1060, n1059, n1058, n1057, n1056, n1055, n1054, n1053, n1052, n1051, n1050, n1049, n1048, n1047} = O_1_6;

clb clb_1_6 ( .clk(clk_1_6), .reset(fpga_rst), .I4(I4_1_6), .I3(I3_1_6), .I2(I2_1_6), .I1(I1_1_6), .O(O_1_6), .config_in(config_chain[49011:47052]), .config_rst(config_rst) );

wire [0:0]clk_1_7;
assign clk_1_7 = {fpga_clk};
wire [12:0]I1_1_7;
assign I1_1_7 = {n1105, n1104, n1103, n1102, n1101, n1100, n1099, n1098, n1097, n1096, n1095, n1094, n1093};
wire [12:0]I2_1_7;
assign I2_1_7 = {n1118, n1117, n1116, n1115, n1114, n1113, n1112, n1111, n1110, n1109, n1108, n1107, n1106};
wire [12:0]I3_1_7;
assign I3_1_7 = {n1131, n1130, n1129, n1128, n1127, n1126, n1125, n1124, n1123, n1122, n1121, n1120, n1119};
wire [12:0]I4_1_7;
assign I4_1_7 = {n1144, n1143, n1142, n1141, n1140, n1139, n1138, n1137, n1136, n1135, n1134, n1133, n1132};
wire [19:0]O_1_7;
assign {n1164, n1163, n1162, n1161, n1160, n1159, n1158, n1157, n1156, n1155, n1154, n1153, n1152, n1151, n1150, n1149, n1148, n1147, n1146, n1145} = O_1_7;

clb clb_1_7 ( .clk(clk_1_7), .reset(fpga_rst), .I4(I4_1_7), .I3(I3_1_7), .I2(I2_1_7), .I1(I1_1_7), .O(O_1_7), .config_in(config_chain[50971:49012]), .config_rst(config_rst) );

wire [0:0]clk_1_8;
assign clk_1_8 = {fpga_clk};
wire [12:0]I1_1_8;
assign I1_1_8 = {n1203, n1202, n1201, n1200, n1199, n1198, n1197, n1196, n1195, n1194, n1193, n1192, n1191};
wire [12:0]I2_1_8;
assign I2_1_8 = {n1216, n1215, n1214, n1213, n1212, n1211, n1210, n1209, n1208, n1207, n1206, n1205, n1204};
wire [12:0]I3_1_8;
assign I3_1_8 = {n1229, n1228, n1227, n1226, n1225, n1224, n1223, n1222, n1221, n1220, n1219, n1218, n1217};
wire [12:0]I4_1_8;
assign I4_1_8 = {n1242, n1241, n1240, n1239, n1238, n1237, n1236, n1235, n1234, n1233, n1232, n1231, n1230};
wire [19:0]O_1_8;
assign {n1262, n1261, n1260, n1259, n1258, n1257, n1256, n1255, n1254, n1253, n1252, n1251, n1250, n1249, n1248, n1247, n1246, n1245, n1244, n1243} = O_1_8;

clb clb_1_8 ( .clk(clk_1_8), .reset(fpga_rst), .I4(I4_1_8), .I3(I3_1_8), .I2(I2_1_8), .I1(I1_1_8), .O(O_1_8), .config_in(config_chain[52931:50972]), .config_rst(config_rst) );

wire [0:0]clk_1_9;
assign clk_1_9 = {fpga_clk};
wire [12:0]I1_1_9;
assign I1_1_9 = {n1301, n1300, n1299, n1298, n1297, n1296, n1295, n1294, n1293, n1292, n1291, n1290, n1289};
wire [12:0]I2_1_9;
assign I2_1_9 = {n1314, n1313, n1312, n1311, n1310, n1309, n1308, n1307, n1306, n1305, n1304, n1303, n1302};
wire [12:0]I3_1_9;
assign I3_1_9 = {n1327, n1326, n1325, n1324, n1323, n1322, n1321, n1320, n1319, n1318, n1317, n1316, n1315};
wire [12:0]I4_1_9;
assign I4_1_9 = {n1340, n1339, n1338, n1337, n1336, n1335, n1334, n1333, n1332, n1331, n1330, n1329, n1328};
wire [19:0]O_1_9;
assign {n1360, n1359, n1358, n1357, n1356, n1355, n1354, n1353, n1352, n1351, n1350, n1349, n1348, n1347, n1346, n1345, n1344, n1343, n1342, n1341} = O_1_9;

clb clb_1_9 ( .clk(clk_1_9), .reset(fpga_rst), .I4(I4_1_9), .I3(I3_1_9), .I2(I2_1_9), .I1(I1_1_9), .O(O_1_9), .config_in(config_chain[54891:52932]), .config_rst(config_rst) );

wire [7:0]outpad_1_10;
assign outpad_1_10 = {n1407, n1404, n1401, n1398, n1395, n1392, n1389, n1386};
wire [7:0]inpad_1_10;
assign {n1408, n1405, n1402, n1399, n1396, n1393, n1390, n1387} = inpad_1_10;

io io_1_10 ( .outpad(outpad_1_10), .inpad(inpad_1_10), .io_ext(io_1_10_wire), .config_in(config_chain[54899:54892]), .config_rst(config_rst) );

wire [7:0]outpad_2_0;
assign outpad_2_0 = {n1455, n1452, n1449, n1446, n1443, n1440, n1437, n1434};
wire [7:0]inpad_2_0;
assign {n1456, n1453, n1450, n1447, n1444, n1441, n1438, n1435} = inpad_2_0;

io io_2_0 ( .outpad(outpad_2_0), .inpad(inpad_2_0), .io_ext(io_2_0_wire), .config_in(config_chain[54907:54900]), .config_rst(config_rst) );

wire [0:0]clk_2_1;
assign clk_2_1 = {fpga_clk};
wire [12:0]I1_2_1;
assign I1_2_1 = {n1495, n1494, n1493, n1492, n1491, n1490, n1489, n1488, n1487, n1486, n1485, n1484, n1483};
wire [12:0]I2_2_1;
assign I2_2_1 = {n1508, n1507, n1506, n1505, n1504, n1503, n1502, n1501, n1500, n1499, n1498, n1497, n1496};
wire [12:0]I3_2_1;
assign I3_2_1 = {n1521, n1520, n1519, n1518, n1517, n1516, n1515, n1514, n1513, n1512, n1511, n1510, n1509};
wire [12:0]I4_2_1;
assign I4_2_1 = {n1534, n1533, n1532, n1531, n1530, n1529, n1528, n1527, n1526, n1525, n1524, n1523, n1522};
wire [19:0]O_2_1;
assign {n1554, n1553, n1552, n1551, n1550, n1549, n1548, n1547, n1546, n1545, n1544, n1543, n1542, n1541, n1540, n1539, n1538, n1537, n1536, n1535} = O_2_1;

clb clb_2_1 ( .clk(clk_2_1), .reset(fpga_rst), .I4(I4_2_1), .I3(I3_2_1), .I2(I2_2_1), .I1(I1_2_1), .O(O_2_1), .config_in(config_chain[56867:54908]), .config_rst(config_rst) );

wire [0:0]clk_2_2;
assign clk_2_2 = {fpga_clk};
wire [12:0]I1_2_2;
assign I1_2_2 = {n1593, n1592, n1591, n1590, n1589, n1588, n1587, n1586, n1585, n1584, n1583, n1582, n1581};
wire [12:0]I2_2_2;
assign I2_2_2 = {n1606, n1605, n1604, n1603, n1602, n1601, n1600, n1599, n1598, n1597, n1596, n1595, n1594};
wire [12:0]I3_2_2;
assign I3_2_2 = {n1619, n1618, n1617, n1616, n1615, n1614, n1613, n1612, n1611, n1610, n1609, n1608, n1607};
wire [12:0]I4_2_2;
assign I4_2_2 = {n1632, n1631, n1630, n1629, n1628, n1627, n1626, n1625, n1624, n1623, n1622, n1621, n1620};
wire [19:0]O_2_2;
assign {n1652, n1651, n1650, n1649, n1648, n1647, n1646, n1645, n1644, n1643, n1642, n1641, n1640, n1639, n1638, n1637, n1636, n1635, n1634, n1633} = O_2_2;

clb clb_2_2 ( .clk(clk_2_2), .reset(fpga_rst), .I4(I4_2_2), .I3(I3_2_2), .I2(I2_2_2), .I1(I1_2_2), .O(O_2_2), .config_in(config_chain[58827:56868]), .config_rst(config_rst) );

wire [0:0]clk_2_3;
assign clk_2_3 = {fpga_clk};
wire [12:0]I1_2_3;
assign I1_2_3 = {n1691, n1690, n1689, n1688, n1687, n1686, n1685, n1684, n1683, n1682, n1681, n1680, n1679};
wire [12:0]I2_2_3;
assign I2_2_3 = {n1704, n1703, n1702, n1701, n1700, n1699, n1698, n1697, n1696, n1695, n1694, n1693, n1692};
wire [12:0]I3_2_3;
assign I3_2_3 = {n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, n1707, n1706, n1705};
wire [12:0]I4_2_3;
assign I4_2_3 = {n1730, n1729, n1728, n1727, n1726, n1725, n1724, n1723, n1722, n1721, n1720, n1719, n1718};
wire [19:0]O_2_3;
assign {n1750, n1749, n1748, n1747, n1746, n1745, n1744, n1743, n1742, n1741, n1740, n1739, n1738, n1737, n1736, n1735, n1734, n1733, n1732, n1731} = O_2_3;

clb clb_2_3 ( .clk(clk_2_3), .reset(fpga_rst), .I4(I4_2_3), .I3(I3_2_3), .I2(I2_2_3), .I1(I1_2_3), .O(O_2_3), .config_in(config_chain[60787:58828]), .config_rst(config_rst) );

wire [0:0]clk_2_4;
assign clk_2_4 = {fpga_clk};
wire [12:0]I1_2_4;
assign I1_2_4 = {n1789, n1788, n1787, n1786, n1785, n1784, n1783, n1782, n1781, n1780, n1779, n1778, n1777};
wire [12:0]I2_2_4;
assign I2_2_4 = {n1802, n1801, n1800, n1799, n1798, n1797, n1796, n1795, n1794, n1793, n1792, n1791, n1790};
wire [12:0]I3_2_4;
assign I3_2_4 = {n1815, n1814, n1813, n1812, n1811, n1810, n1809, n1808, n1807, n1806, n1805, n1804, n1803};
wire [12:0]I4_2_4;
assign I4_2_4 = {n1828, n1827, n1826, n1825, n1824, n1823, n1822, n1821, n1820, n1819, n1818, n1817, n1816};
wire [19:0]O_2_4;
assign {n1848, n1847, n1846, n1845, n1844, n1843, n1842, n1841, n1840, n1839, n1838, n1837, n1836, n1835, n1834, n1833, n1832, n1831, n1830, n1829} = O_2_4;

clb clb_2_4 ( .clk(clk_2_4), .reset(fpga_rst), .I4(I4_2_4), .I3(I3_2_4), .I2(I2_2_4), .I1(I1_2_4), .O(O_2_4), .config_in(config_chain[62747:60788]), .config_rst(config_rst) );

wire [0:0]clk_2_5;
assign clk_2_5 = {fpga_clk};
wire [12:0]I1_2_5;
assign I1_2_5 = {n1887, n1886, n1885, n1884, n1883, n1882, n1881, n1880, n1879, n1878, n1877, n1876, n1875};
wire [12:0]I2_2_5;
assign I2_2_5 = {n1900, n1899, n1898, n1897, n1896, n1895, n1894, n1893, n1892, n1891, n1890, n1889, n1888};
wire [12:0]I3_2_5;
assign I3_2_5 = {n1913, n1912, n1911, n1910, n1909, n1908, n1907, n1906, n1905, n1904, n1903, n1902, n1901};
wire [12:0]I4_2_5;
assign I4_2_5 = {n1926, n1925, n1924, n1923, n1922, n1921, n1920, n1919, n1918, n1917, n1916, n1915, n1914};
wire [19:0]O_2_5;
assign {n1946, n1945, n1944, n1943, n1942, n1941, n1940, n1939, n1938, n1937, n1936, n1935, n1934, n1933, n1932, n1931, n1930, n1929, n1928, n1927} = O_2_5;

clb clb_2_5 ( .clk(clk_2_5), .reset(fpga_rst), .I4(I4_2_5), .I3(I3_2_5), .I2(I2_2_5), .I1(I1_2_5), .O(O_2_5), .config_in(config_chain[64707:62748]), .config_rst(config_rst) );

wire [0:0]clk_2_6;
assign clk_2_6 = {fpga_clk};
wire [12:0]I1_2_6;
assign I1_2_6 = {n1985, n1984, n1983, n1982, n1981, n1980, n1979, n1978, n1977, n1976, n1975, n1974, n1973};
wire [12:0]I2_2_6;
assign I2_2_6 = {n1998, n1997, n1996, n1995, n1994, n1993, n1992, n1991, n1990, n1989, n1988, n1987, n1986};
wire [12:0]I3_2_6;
assign I3_2_6 = {n2011, n2010, n2009, n2008, n2007, n2006, n2005, n2004, n2003, n2002, n2001, n2000, n1999};
wire [12:0]I4_2_6;
assign I4_2_6 = {n2024, n2023, n2022, n2021, n2020, n2019, n2018, n2017, n2016, n2015, n2014, n2013, n2012};
wire [19:0]O_2_6;
assign {n2044, n2043, n2042, n2041, n2040, n2039, n2038, n2037, n2036, n2035, n2034, n2033, n2032, n2031, n2030, n2029, n2028, n2027, n2026, n2025} = O_2_6;

clb clb_2_6 ( .clk(clk_2_6), .reset(fpga_rst), .I4(I4_2_6), .I3(I3_2_6), .I2(I2_2_6), .I1(I1_2_6), .O(O_2_6), .config_in(config_chain[66667:64708]), .config_rst(config_rst) );

wire [0:0]clk_2_7;
assign clk_2_7 = {fpga_clk};
wire [12:0]I1_2_7;
assign I1_2_7 = {n2083, n2082, n2081, n2080, n2079, n2078, n2077, n2076, n2075, n2074, n2073, n2072, n2071};
wire [12:0]I2_2_7;
assign I2_2_7 = {n2096, n2095, n2094, n2093, n2092, n2091, n2090, n2089, n2088, n2087, n2086, n2085, n2084};
wire [12:0]I3_2_7;
assign I3_2_7 = {n2109, n2108, n2107, n2106, n2105, n2104, n2103, n2102, n2101, n2100, n2099, n2098, n2097};
wire [12:0]I4_2_7;
assign I4_2_7 = {n2122, n2121, n2120, n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, n2111, n2110};
wire [19:0]O_2_7;
assign {n2142, n2141, n2140, n2139, n2138, n2137, n2136, n2135, n2134, n2133, n2132, n2131, n2130, n2129, n2128, n2127, n2126, n2125, n2124, n2123} = O_2_7;

clb clb_2_7 ( .clk(clk_2_7), .reset(fpga_rst), .I4(I4_2_7), .I3(I3_2_7), .I2(I2_2_7), .I1(I1_2_7), .O(O_2_7), .config_in(config_chain[68627:66668]), .config_rst(config_rst) );

wire [0:0]clk_2_8;
assign clk_2_8 = {fpga_clk};
wire [12:0]I1_2_8;
assign I1_2_8 = {n2181, n2180, n2179, n2178, n2177, n2176, n2175, n2174, n2173, n2172, n2171, n2170, n2169};
wire [12:0]I2_2_8;
assign I2_2_8 = {n2194, n2193, n2192, n2191, n2190, n2189, n2188, n2187, n2186, n2185, n2184, n2183, n2182};
wire [12:0]I3_2_8;
assign I3_2_8 = {n2207, n2206, n2205, n2204, n2203, n2202, n2201, n2200, n2199, n2198, n2197, n2196, n2195};
wire [12:0]I4_2_8;
assign I4_2_8 = {n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, n2212, n2211, n2210, n2209, n2208};
wire [19:0]O_2_8;
assign {n2240, n2239, n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231, n2230, n2229, n2228, n2227, n2226, n2225, n2224, n2223, n2222, n2221} = O_2_8;

clb clb_2_8 ( .clk(clk_2_8), .reset(fpga_rst), .I4(I4_2_8), .I3(I3_2_8), .I2(I2_2_8), .I1(I1_2_8), .O(O_2_8), .config_in(config_chain[70587:68628]), .config_rst(config_rst) );

wire [0:0]clk_2_9;
assign clk_2_9 = {fpga_clk};
wire [12:0]I1_2_9;
assign I1_2_9 = {n2279, n2278, n2277, n2276, n2275, n2274, n2273, n2272, n2271, n2270, n2269, n2268, n2267};
wire [12:0]I2_2_9;
assign I2_2_9 = {n2292, n2291, n2290, n2289, n2288, n2287, n2286, n2285, n2284, n2283, n2282, n2281, n2280};
wire [12:0]I3_2_9;
assign I3_2_9 = {n2305, n2304, n2303, n2302, n2301, n2300, n2299, n2298, n2297, n2296, n2295, n2294, n2293};
wire [12:0]I4_2_9;
assign I4_2_9 = {n2318, n2317, n2316, n2315, n2314, n2313, n2312, n2311, n2310, n2309, n2308, n2307, n2306};
wire [19:0]O_2_9;
assign {n2338, n2337, n2336, n2335, n2334, n2333, n2332, n2331, n2330, n2329, n2328, n2327, n2326, n2325, n2324, n2323, n2322, n2321, n2320, n2319} = O_2_9;

clb clb_2_9 ( .clk(clk_2_9), .reset(fpga_rst), .I4(I4_2_9), .I3(I3_2_9), .I2(I2_2_9), .I1(I1_2_9), .O(O_2_9), .config_in(config_chain[72547:70588]), .config_rst(config_rst) );

wire [7:0]outpad_2_10;
assign outpad_2_10 = {n2385, n2382, n2379, n2376, n2373, n2370, n2367, n2364};
wire [7:0]inpad_2_10;
assign {n2386, n2383, n2380, n2377, n2374, n2371, n2368, n2365} = inpad_2_10;

io io_2_10 ( .outpad(outpad_2_10), .inpad(inpad_2_10), .io_ext(io_2_10_wire), .config_in(config_chain[72555:72548]), .config_rst(config_rst) );

wire [7:0]outpad_3_0;
assign outpad_3_0 = {n2433, n2430, n2427, n2424, n2421, n2418, n2415, n2412};
wire [7:0]inpad_3_0;
assign {n2434, n2431, n2428, n2425, n2422, n2419, n2416, n2413} = inpad_3_0;

io io_3_0 ( .outpad(outpad_3_0), .inpad(inpad_3_0), .io_ext(io_3_0_wire), .config_in(config_chain[72563:72556]), .config_rst(config_rst) );

wire [0:0]clk_3_1;
assign clk_3_1 = {fpga_clk};
wire [12:0]I1_3_1;
assign I1_3_1 = {n2473, n2472, n2471, n2470, n2469, n2468, n2467, n2466, n2465, n2464, n2463, n2462, n2461};
wire [12:0]I2_3_1;
assign I2_3_1 = {n2486, n2485, n2484, n2483, n2482, n2481, n2480, n2479, n2478, n2477, n2476, n2475, n2474};
wire [12:0]I3_3_1;
assign I3_3_1 = {n2499, n2498, n2497, n2496, n2495, n2494, n2493, n2492, n2491, n2490, n2489, n2488, n2487};
wire [12:0]I4_3_1;
assign I4_3_1 = {n2512, n2511, n2510, n2509, n2508, n2507, n2506, n2505, n2504, n2503, n2502, n2501, n2500};
wire [19:0]O_3_1;
assign {n2532, n2531, n2530, n2529, n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2520, n2519, n2518, n2517, n2516, n2515, n2514, n2513} = O_3_1;

clb clb_3_1 ( .clk(clk_3_1), .reset(fpga_rst), .I4(I4_3_1), .I3(I3_3_1), .I2(I2_3_1), .I1(I1_3_1), .O(O_3_1), .config_in(config_chain[74523:72564]), .config_rst(config_rst) );

wire [0:0]clk_3_2;
assign clk_3_2 = {fpga_clk};
wire [12:0]I1_3_2;
assign I1_3_2 = {n2571, n2570, n2569, n2568, n2567, n2566, n2565, n2564, n2563, n2562, n2561, n2560, n2559};
wire [12:0]I2_3_2;
assign I2_3_2 = {n2584, n2583, n2582, n2581, n2580, n2579, n2578, n2577, n2576, n2575, n2574, n2573, n2572};
wire [12:0]I3_3_2;
assign I3_3_2 = {n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588, n2587, n2586, n2585};
wire [12:0]I4_3_2;
assign I4_3_2 = {n2610, n2609, n2608, n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598};
wire [19:0]O_3_2;
assign {n2630, n2629, n2628, n2627, n2626, n2625, n2624, n2623, n2622, n2621, n2620, n2619, n2618, n2617, n2616, n2615, n2614, n2613, n2612, n2611} = O_3_2;

clb clb_3_2 ( .clk(clk_3_2), .reset(fpga_rst), .I4(I4_3_2), .I3(I3_3_2), .I2(I2_3_2), .I1(I1_3_2), .O(O_3_2), .config_in(config_chain[76483:74524]), .config_rst(config_rst) );

wire [0:0]clk_3_3;
assign clk_3_3 = {fpga_clk};
wire [12:0]I1_3_3;
assign I1_3_3 = {n2669, n2668, n2667, n2666, n2665, n2664, n2663, n2662, n2661, n2660, n2659, n2658, n2657};
wire [12:0]I2_3_3;
assign I2_3_3 = {n2682, n2681, n2680, n2679, n2678, n2677, n2676, n2675, n2674, n2673, n2672, n2671, n2670};
wire [12:0]I3_3_3;
assign I3_3_3 = {n2695, n2694, n2693, n2692, n2691, n2690, n2689, n2688, n2687, n2686, n2685, n2684, n2683};
wire [12:0]I4_3_3;
assign I4_3_3 = {n2708, n2707, n2706, n2705, n2704, n2703, n2702, n2701, n2700, n2699, n2698, n2697, n2696};
wire [19:0]O_3_3;
assign {n2728, n2727, n2726, n2725, n2724, n2723, n2722, n2721, n2720, n2719, n2718, n2717, n2716, n2715, n2714, n2713, n2712, n2711, n2710, n2709} = O_3_3;

clb clb_3_3 ( .clk(clk_3_3), .reset(fpga_rst), .I4(I4_3_3), .I3(I3_3_3), .I2(I2_3_3), .I1(I1_3_3), .O(O_3_3), .config_in(config_chain[78443:76484]), .config_rst(config_rst) );

wire [0:0]clk_3_4;
assign clk_3_4 = {fpga_clk};
wire [12:0]I1_3_4;
assign I1_3_4 = {n2767, n2766, n2765, n2764, n2763, n2762, n2761, n2760, n2759, n2758, n2757, n2756, n2755};
wire [12:0]I2_3_4;
assign I2_3_4 = {n2780, n2779, n2778, n2777, n2776, n2775, n2774, n2773, n2772, n2771, n2770, n2769, n2768};
wire [12:0]I3_3_4;
assign I3_3_4 = {n2793, n2792, n2791, n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2783, n2782, n2781};
wire [12:0]I4_3_4;
assign I4_3_4 = {n2806, n2805, n2804, n2803, n2802, n2801, n2800, n2799, n2798, n2797, n2796, n2795, n2794};
wire [19:0]O_3_4;
assign {n2826, n2825, n2824, n2823, n2822, n2821, n2820, n2819, n2818, n2817, n2816, n2815, n2814, n2813, n2812, n2811, n2810, n2809, n2808, n2807} = O_3_4;

clb clb_3_4 ( .clk(clk_3_4), .reset(fpga_rst), .I4(I4_3_4), .I3(I3_3_4), .I2(I2_3_4), .I1(I1_3_4), .O(O_3_4), .config_in(config_chain[80403:78444]), .config_rst(config_rst) );

wire [0:0]clk_3_5;
assign clk_3_5 = {fpga_clk};
wire [12:0]I1_3_5;
assign I1_3_5 = {n2865, n2864, n2863, n2862, n2861, n2860, n2859, n2858, n2857, n2856, n2855, n2854, n2853};
wire [12:0]I2_3_5;
assign I2_3_5 = {n2878, n2877, n2876, n2875, n2874, n2873, n2872, n2871, n2870, n2869, n2868, n2867, n2866};
wire [12:0]I3_3_5;
assign I3_3_5 = {n2891, n2890, n2889, n2888, n2887, n2886, n2885, n2884, n2883, n2882, n2881, n2880, n2879};
wire [12:0]I4_3_5;
assign I4_3_5 = {n2904, n2903, n2902, n2901, n2900, n2899, n2898, n2897, n2896, n2895, n2894, n2893, n2892};
wire [19:0]O_3_5;
assign {n2924, n2923, n2922, n2921, n2920, n2919, n2918, n2917, n2916, n2915, n2914, n2913, n2912, n2911, n2910, n2909, n2908, n2907, n2906, n2905} = O_3_5;

clb clb_3_5 ( .clk(clk_3_5), .reset(fpga_rst), .I4(I4_3_5), .I3(I3_3_5), .I2(I2_3_5), .I1(I1_3_5), .O(O_3_5), .config_in(config_chain[82363:80404]), .config_rst(config_rst) );

wire [0:0]clk_3_6;
assign clk_3_6 = {fpga_clk};
wire [12:0]I1_3_6;
assign I1_3_6 = {n2963, n2962, n2961, n2960, n2959, n2958, n2957, n2956, n2955, n2954, n2953, n2952, n2951};
wire [12:0]I2_3_6;
assign I2_3_6 = {n2976, n2975, n2974, n2973, n2972, n2971, n2970, n2969, n2968, n2967, n2966, n2965, n2964};
wire [12:0]I3_3_6;
assign I3_3_6 = {n2989, n2988, n2987, n2986, n2985, n2984, n2983, n2982, n2981, n2980, n2979, n2978, n2977};
wire [12:0]I4_3_6;
assign I4_3_6 = {n3002, n3001, n3000, n2999, n2998, n2997, n2996, n2995, n2994, n2993, n2992, n2991, n2990};
wire [19:0]O_3_6;
assign {n3022, n3021, n3020, n3019, n3018, n3017, n3016, n3015, n3014, n3013, n3012, n3011, n3010, n3009, n3008, n3007, n3006, n3005, n3004, n3003} = O_3_6;

clb clb_3_6 ( .clk(clk_3_6), .reset(fpga_rst), .I4(I4_3_6), .I3(I3_3_6), .I2(I2_3_6), .I1(I1_3_6), .O(O_3_6), .config_in(config_chain[84323:82364]), .config_rst(config_rst) );

wire [0:0]clk_3_7;
assign clk_3_7 = {fpga_clk};
wire [12:0]I1_3_7;
assign I1_3_7 = {n3061, n3060, n3059, n3058, n3057, n3056, n3055, n3054, n3053, n3052, n3051, n3050, n3049};
wire [12:0]I2_3_7;
assign I2_3_7 = {n3074, n3073, n3072, n3071, n3070, n3069, n3068, n3067, n3066, n3065, n3064, n3063, n3062};
wire [12:0]I3_3_7;
assign I3_3_7 = {n3087, n3086, n3085, n3084, n3083, n3082, n3081, n3080, n3079, n3078, n3077, n3076, n3075};
wire [12:0]I4_3_7;
assign I4_3_7 = {n3100, n3099, n3098, n3097, n3096, n3095, n3094, n3093, n3092, n3091, n3090, n3089, n3088};
wire [19:0]O_3_7;
assign {n3120, n3119, n3118, n3117, n3116, n3115, n3114, n3113, n3112, n3111, n3110, n3109, n3108, n3107, n3106, n3105, n3104, n3103, n3102, n3101} = O_3_7;

clb clb_3_7 ( .clk(clk_3_7), .reset(fpga_rst), .I4(I4_3_7), .I3(I3_3_7), .I2(I2_3_7), .I1(I1_3_7), .O(O_3_7), .config_in(config_chain[86283:84324]), .config_rst(config_rst) );

wire [0:0]clk_3_8;
assign clk_3_8 = {fpga_clk};
wire [12:0]I1_3_8;
assign I1_3_8 = {n3159, n3158, n3157, n3156, n3155, n3154, n3153, n3152, n3151, n3150, n3149, n3148, n3147};
wire [12:0]I2_3_8;
assign I2_3_8 = {n3172, n3171, n3170, n3169, n3168, n3167, n3166, n3165, n3164, n3163, n3162, n3161, n3160};
wire [12:0]I3_3_8;
assign I3_3_8 = {n3185, n3184, n3183, n3182, n3181, n3180, n3179, n3178, n3177, n3176, n3175, n3174, n3173};
wire [12:0]I4_3_8;
assign I4_3_8 = {n3198, n3197, n3196, n3195, n3194, n3193, n3192, n3191, n3190, n3189, n3188, n3187, n3186};
wire [19:0]O_3_8;
assign {n3218, n3217, n3216, n3215, n3214, n3213, n3212, n3211, n3210, n3209, n3208, n3207, n3206, n3205, n3204, n3203, n3202, n3201, n3200, n3199} = O_3_8;

clb clb_3_8 ( .clk(clk_3_8), .reset(fpga_rst), .I4(I4_3_8), .I3(I3_3_8), .I2(I2_3_8), .I1(I1_3_8), .O(O_3_8), .config_in(config_chain[88243:86284]), .config_rst(config_rst) );

wire [0:0]clk_3_9;
assign clk_3_9 = {fpga_clk};
wire [12:0]I1_3_9;
assign I1_3_9 = {n3257, n3256, n3255, n3254, n3253, n3252, n3251, n3250, n3249, n3248, n3247, n3246, n3245};
wire [12:0]I2_3_9;
assign I2_3_9 = {n3270, n3269, n3268, n3267, n3266, n3265, n3264, n3263, n3262, n3261, n3260, n3259, n3258};
wire [12:0]I3_3_9;
assign I3_3_9 = {n3283, n3282, n3281, n3280, n3279, n3278, n3277, n3276, n3275, n3274, n3273, n3272, n3271};
wire [12:0]I4_3_9;
assign I4_3_9 = {n3296, n3295, n3294, n3293, n3292, n3291, n3290, n3289, n3288, n3287, n3286, n3285, n3284};
wire [19:0]O_3_9;
assign {n3316, n3315, n3314, n3313, n3312, n3311, n3310, n3309, n3308, n3307, n3306, n3305, n3304, n3303, n3302, n3301, n3300, n3299, n3298, n3297} = O_3_9;

clb clb_3_9 ( .clk(clk_3_9), .reset(fpga_rst), .I4(I4_3_9), .I3(I3_3_9), .I2(I2_3_9), .I1(I1_3_9), .O(O_3_9), .config_in(config_chain[90203:88244]), .config_rst(config_rst) );

wire [7:0]outpad_3_10;
assign outpad_3_10 = {n3363, n3360, n3357, n3354, n3351, n3348, n3345, n3342};
wire [7:0]inpad_3_10;
assign {n3364, n3361, n3358, n3355, n3352, n3349, n3346, n3343} = inpad_3_10;

io io_3_10 ( .outpad(outpad_3_10), .inpad(inpad_3_10), .io_ext(io_3_10_wire), .config_in(config_chain[90211:90204]), .config_rst(config_rst) );

wire [7:0]outpad_4_0;
assign outpad_4_0 = {n3411, n3408, n3405, n3402, n3399, n3396, n3393, n3390};
wire [7:0]inpad_4_0;
assign {n3412, n3409, n3406, n3403, n3400, n3397, n3394, n3391} = inpad_4_0;

io io_4_0 ( .outpad(outpad_4_0), .inpad(inpad_4_0), .io_ext(io_4_0_wire), .config_in(config_chain[90219:90212]), .config_rst(config_rst) );

wire [0:0]clk_4_1;
assign clk_4_1 = {fpga_clk};
wire [12:0]I1_4_1;
assign I1_4_1 = {n3451, n3450, n3449, n3448, n3447, n3446, n3445, n3444, n3443, n3442, n3441, n3440, n3439};
wire [12:0]I2_4_1;
assign I2_4_1 = {n3464, n3463, n3462, n3461, n3460, n3459, n3458, n3457, n3456, n3455, n3454, n3453, n3452};
wire [12:0]I3_4_1;
assign I3_4_1 = {n3477, n3476, n3475, n3474, n3473, n3472, n3471, n3470, n3469, n3468, n3467, n3466, n3465};
wire [12:0]I4_4_1;
assign I4_4_1 = {n3490, n3489, n3488, n3487, n3486, n3485, n3484, n3483, n3482, n3481, n3480, n3479, n3478};
wire [19:0]O_4_1;
assign {n3510, n3509, n3508, n3507, n3506, n3505, n3504, n3503, n3502, n3501, n3500, n3499, n3498, n3497, n3496, n3495, n3494, n3493, n3492, n3491} = O_4_1;

clb clb_4_1 ( .clk(clk_4_1), .reset(fpga_rst), .I4(I4_4_1), .I3(I3_4_1), .I2(I2_4_1), .I1(I1_4_1), .O(O_4_1), .config_in(config_chain[92179:90220]), .config_rst(config_rst) );

wire [0:0]clk_4_2;
assign clk_4_2 = {fpga_clk};
wire [12:0]I1_4_2;
assign I1_4_2 = {n3549, n3548, n3547, n3546, n3545, n3544, n3543, n3542, n3541, n3540, n3539, n3538, n3537};
wire [12:0]I2_4_2;
assign I2_4_2 = {n3562, n3561, n3560, n3559, n3558, n3557, n3556, n3555, n3554, n3553, n3552, n3551, n3550};
wire [12:0]I3_4_2;
assign I3_4_2 = {n3575, n3574, n3573, n3572, n3571, n3570, n3569, n3568, n3567, n3566, n3565, n3564, n3563};
wire [12:0]I4_4_2;
assign I4_4_2 = {n3588, n3587, n3586, n3585, n3584, n3583, n3582, n3581, n3580, n3579, n3578, n3577, n3576};
wire [19:0]O_4_2;
assign {n3608, n3607, n3606, n3605, n3604, n3603, n3602, n3601, n3600, n3599, n3598, n3597, n3596, n3595, n3594, n3593, n3592, n3591, n3590, n3589} = O_4_2;

clb clb_4_2 ( .clk(clk_4_2), .reset(fpga_rst), .I4(I4_4_2), .I3(I3_4_2), .I2(I2_4_2), .I1(I1_4_2), .O(O_4_2), .config_in(config_chain[94139:92180]), .config_rst(config_rst) );

wire [0:0]clk_4_3;
assign clk_4_3 = {fpga_clk};
wire [12:0]I1_4_3;
assign I1_4_3 = {n3647, n3646, n3645, n3644, n3643, n3642, n3641, n3640, n3639, n3638, n3637, n3636, n3635};
wire [12:0]I2_4_3;
assign I2_4_3 = {n3660, n3659, n3658, n3657, n3656, n3655, n3654, n3653, n3652, n3651, n3650, n3649, n3648};
wire [12:0]I3_4_3;
assign I3_4_3 = {n3673, n3672, n3671, n3670, n3669, n3668, n3667, n3666, n3665, n3664, n3663, n3662, n3661};
wire [12:0]I4_4_3;
assign I4_4_3 = {n3686, n3685, n3684, n3683, n3682, n3681, n3680, n3679, n3678, n3677, n3676, n3675, n3674};
wire [19:0]O_4_3;
assign {n3706, n3705, n3704, n3703, n3702, n3701, n3700, n3699, n3698, n3697, n3696, n3695, n3694, n3693, n3692, n3691, n3690, n3689, n3688, n3687} = O_4_3;

clb clb_4_3 ( .clk(clk_4_3), .reset(fpga_rst), .I4(I4_4_3), .I3(I3_4_3), .I2(I2_4_3), .I1(I1_4_3), .O(O_4_3), .config_in(config_chain[96099:94140]), .config_rst(config_rst) );

wire [0:0]clk_4_4;
assign clk_4_4 = {fpga_clk};
wire [12:0]I1_4_4;
assign I1_4_4 = {n3745, n3744, n3743, n3742, n3741, n3740, n3739, n3738, n3737, n3736, n3735, n3734, n3733};
wire [12:0]I2_4_4;
assign I2_4_4 = {n3758, n3757, n3756, n3755, n3754, n3753, n3752, n3751, n3750, n3749, n3748, n3747, n3746};
wire [12:0]I3_4_4;
assign I3_4_4 = {n3771, n3770, n3769, n3768, n3767, n3766, n3765, n3764, n3763, n3762, n3761, n3760, n3759};
wire [12:0]I4_4_4;
assign I4_4_4 = {n3784, n3783, n3782, n3781, n3780, n3779, n3778, n3777, n3776, n3775, n3774, n3773, n3772};
wire [19:0]O_4_4;
assign {n3804, n3803, n3802, n3801, n3800, n3799, n3798, n3797, n3796, n3795, n3794, n3793, n3792, n3791, n3790, n3789, n3788, n3787, n3786, n3785} = O_4_4;

clb clb_4_4 ( .clk(clk_4_4), .reset(fpga_rst), .I4(I4_4_4), .I3(I3_4_4), .I2(I2_4_4), .I1(I1_4_4), .O(O_4_4), .config_in(config_chain[98059:96100]), .config_rst(config_rst) );

wire [0:0]clk_4_5;
assign clk_4_5 = {fpga_clk};
wire [12:0]I1_4_5;
assign I1_4_5 = {n3843, n3842, n3841, n3840, n3839, n3838, n3837, n3836, n3835, n3834, n3833, n3832, n3831};
wire [12:0]I2_4_5;
assign I2_4_5 = {n3856, n3855, n3854, n3853, n3852, n3851, n3850, n3849, n3848, n3847, n3846, n3845, n3844};
wire [12:0]I3_4_5;
assign I3_4_5 = {n3869, n3868, n3867, n3866, n3865, n3864, n3863, n3862, n3861, n3860, n3859, n3858, n3857};
wire [12:0]I4_4_5;
assign I4_4_5 = {n3882, n3881, n3880, n3879, n3878, n3877, n3876, n3875, n3874, n3873, n3872, n3871, n3870};
wire [19:0]O_4_5;
assign {n3902, n3901, n3900, n3899, n3898, n3897, n3896, n3895, n3894, n3893, n3892, n3891, n3890, n3889, n3888, n3887, n3886, n3885, n3884, n3883} = O_4_5;

clb clb_4_5 ( .clk(clk_4_5), .reset(fpga_rst), .I4(I4_4_5), .I3(I3_4_5), .I2(I2_4_5), .I1(I1_4_5), .O(O_4_5), .config_in(config_chain[100019:98060]), .config_rst(config_rst) );

wire [0:0]clk_4_6;
assign clk_4_6 = {fpga_clk};
wire [12:0]I1_4_6;
assign I1_4_6 = {n3941, n3940, n3939, n3938, n3937, n3936, n3935, n3934, n3933, n3932, n3931, n3930, n3929};
wire [12:0]I2_4_6;
assign I2_4_6 = {n3954, n3953, n3952, n3951, n3950, n3949, n3948, n3947, n3946, n3945, n3944, n3943, n3942};
wire [12:0]I3_4_6;
assign I3_4_6 = {n3967, n3966, n3965, n3964, n3963, n3962, n3961, n3960, n3959, n3958, n3957, n3956, n3955};
wire [12:0]I4_4_6;
assign I4_4_6 = {n3980, n3979, n3978, n3977, n3976, n3975, n3974, n3973, n3972, n3971, n3970, n3969, n3968};
wire [19:0]O_4_6;
assign {n4000, n3999, n3998, n3997, n3996, n3995, n3994, n3993, n3992, n3991, n3990, n3989, n3988, n3987, n3986, n3985, n3984, n3983, n3982, n3981} = O_4_6;

clb clb_4_6 ( .clk(clk_4_6), .reset(fpga_rst), .I4(I4_4_6), .I3(I3_4_6), .I2(I2_4_6), .I1(I1_4_6), .O(O_4_6), .config_in(config_chain[101979:100020]), .config_rst(config_rst) );

wire [0:0]clk_4_7;
assign clk_4_7 = {fpga_clk};
wire [12:0]I1_4_7;
assign I1_4_7 = {n4039, n4038, n4037, n4036, n4035, n4034, n4033, n4032, n4031, n4030, n4029, n4028, n4027};
wire [12:0]I2_4_7;
assign I2_4_7 = {n4052, n4051, n4050, n4049, n4048, n4047, n4046, n4045, n4044, n4043, n4042, n4041, n4040};
wire [12:0]I3_4_7;
assign I3_4_7 = {n4065, n4064, n4063, n4062, n4061, n4060, n4059, n4058, n4057, n4056, n4055, n4054, n4053};
wire [12:0]I4_4_7;
assign I4_4_7 = {n4078, n4077, n4076, n4075, n4074, n4073, n4072, n4071, n4070, n4069, n4068, n4067, n4066};
wire [19:0]O_4_7;
assign {n4098, n4097, n4096, n4095, n4094, n4093, n4092, n4091, n4090, n4089, n4088, n4087, n4086, n4085, n4084, n4083, n4082, n4081, n4080, n4079} = O_4_7;

clb clb_4_7 ( .clk(clk_4_7), .reset(fpga_rst), .I4(I4_4_7), .I3(I3_4_7), .I2(I2_4_7), .I1(I1_4_7), .O(O_4_7), .config_in(config_chain[103939:101980]), .config_rst(config_rst) );

wire [0:0]clk_4_8;
assign clk_4_8 = {fpga_clk};
wire [12:0]I1_4_8;
assign I1_4_8 = {n4137, n4136, n4135, n4134, n4133, n4132, n4131, n4130, n4129, n4128, n4127, n4126, n4125};
wire [12:0]I2_4_8;
assign I2_4_8 = {n4150, n4149, n4148, n4147, n4146, n4145, n4144, n4143, n4142, n4141, n4140, n4139, n4138};
wire [12:0]I3_4_8;
assign I3_4_8 = {n4163, n4162, n4161, n4160, n4159, n4158, n4157, n4156, n4155, n4154, n4153, n4152, n4151};
wire [12:0]I4_4_8;
assign I4_4_8 = {n4176, n4175, n4174, n4173, n4172, n4171, n4170, n4169, n4168, n4167, n4166, n4165, n4164};
wire [19:0]O_4_8;
assign {n4196, n4195, n4194, n4193, n4192, n4191, n4190, n4189, n4188, n4187, n4186, n4185, n4184, n4183, n4182, n4181, n4180, n4179, n4178, n4177} = O_4_8;

clb clb_4_8 ( .clk(clk_4_8), .reset(fpga_rst), .I4(I4_4_8), .I3(I3_4_8), .I2(I2_4_8), .I1(I1_4_8), .O(O_4_8), .config_in(config_chain[105899:103940]), .config_rst(config_rst) );

wire [0:0]clk_4_9;
assign clk_4_9 = {fpga_clk};
wire [12:0]I1_4_9;
assign I1_4_9 = {n4235, n4234, n4233, n4232, n4231, n4230, n4229, n4228, n4227, n4226, n4225, n4224, n4223};
wire [12:0]I2_4_9;
assign I2_4_9 = {n4248, n4247, n4246, n4245, n4244, n4243, n4242, n4241, n4240, n4239, n4238, n4237, n4236};
wire [12:0]I3_4_9;
assign I3_4_9 = {n4261, n4260, n4259, n4258, n4257, n4256, n4255, n4254, n4253, n4252, n4251, n4250, n4249};
wire [12:0]I4_4_9;
assign I4_4_9 = {n4274, n4273, n4272, n4271, n4270, n4269, n4268, n4267, n4266, n4265, n4264, n4263, n4262};
wire [19:0]O_4_9;
assign {n4294, n4293, n4292, n4291, n4290, n4289, n4288, n4287, n4286, n4285, n4284, n4283, n4282, n4281, n4280, n4279, n4278, n4277, n4276, n4275} = O_4_9;

clb clb_4_9 ( .clk(clk_4_9), .reset(fpga_rst), .I4(I4_4_9), .I3(I3_4_9), .I2(I2_4_9), .I1(I1_4_9), .O(O_4_9), .config_in(config_chain[107859:105900]), .config_rst(config_rst) );

wire [7:0]outpad_4_10;
assign outpad_4_10 = {n4341, n4338, n4335, n4332, n4329, n4326, n4323, n4320};
wire [7:0]inpad_4_10;
assign {n4342, n4339, n4336, n4333, n4330, n4327, n4324, n4321} = inpad_4_10;

io io_4_10 ( .outpad(outpad_4_10), .inpad(inpad_4_10), .io_ext(io_4_10_wire), .config_in(config_chain[107867:107860]), .config_rst(config_rst) );

wire [7:0]outpad_5_0;
assign outpad_5_0 = {n4389, n4386, n4383, n4380, n4377, n4374, n4371, n4368};
wire [7:0]inpad_5_0;
assign {n4390, n4387, n4384, n4381, n4378, n4375, n4372, n4369} = inpad_5_0;

io io_5_0 ( .outpad(outpad_5_0), .inpad(inpad_5_0), .io_ext(io_5_0_wire), .config_in(config_chain[107875:107868]), .config_rst(config_rst) );

wire [0:0]clk_5_1;
assign clk_5_1 = {fpga_clk};
wire [12:0]I1_5_1;
assign I1_5_1 = {n4429, n4428, n4427, n4426, n4425, n4424, n4423, n4422, n4421, n4420, n4419, n4418, n4417};
wire [12:0]I2_5_1;
assign I2_5_1 = {n4442, n4441, n4440, n4439, n4438, n4437, n4436, n4435, n4434, n4433, n4432, n4431, n4430};
wire [12:0]I3_5_1;
assign I3_5_1 = {n4455, n4454, n4453, n4452, n4451, n4450, n4449, n4448, n4447, n4446, n4445, n4444, n4443};
wire [12:0]I4_5_1;
assign I4_5_1 = {n4468, n4467, n4466, n4465, n4464, n4463, n4462, n4461, n4460, n4459, n4458, n4457, n4456};
wire [19:0]O_5_1;
assign {n4488, n4487, n4486, n4485, n4484, n4483, n4482, n4481, n4480, n4479, n4478, n4477, n4476, n4475, n4474, n4473, n4472, n4471, n4470, n4469} = O_5_1;

clb clb_5_1 ( .clk(clk_5_1), .reset(fpga_rst), .I4(I4_5_1), .I3(I3_5_1), .I2(I2_5_1), .I1(I1_5_1), .O(O_5_1), .config_in(config_chain[109835:107876]), .config_rst(config_rst) );

wire [0:0]clk_5_2;
assign clk_5_2 = {fpga_clk};
wire [12:0]I1_5_2;
assign I1_5_2 = {n4527, n4526, n4525, n4524, n4523, n4522, n4521, n4520, n4519, n4518, n4517, n4516, n4515};
wire [12:0]I2_5_2;
assign I2_5_2 = {n4540, n4539, n4538, n4537, n4536, n4535, n4534, n4533, n4532, n4531, n4530, n4529, n4528};
wire [12:0]I3_5_2;
assign I3_5_2 = {n4553, n4552, n4551, n4550, n4549, n4548, n4547, n4546, n4545, n4544, n4543, n4542, n4541};
wire [12:0]I4_5_2;
assign I4_5_2 = {n4566, n4565, n4564, n4563, n4562, n4561, n4560, n4559, n4558, n4557, n4556, n4555, n4554};
wire [19:0]O_5_2;
assign {n4586, n4585, n4584, n4583, n4582, n4581, n4580, n4579, n4578, n4577, n4576, n4575, n4574, n4573, n4572, n4571, n4570, n4569, n4568, n4567} = O_5_2;

clb clb_5_2 ( .clk(clk_5_2), .reset(fpga_rst), .I4(I4_5_2), .I3(I3_5_2), .I2(I2_5_2), .I1(I1_5_2), .O(O_5_2), .config_in(config_chain[111795:109836]), .config_rst(config_rst) );

wire [0:0]clk_5_3;
assign clk_5_3 = {fpga_clk};
wire [12:0]I1_5_3;
assign I1_5_3 = {n4625, n4624, n4623, n4622, n4621, n4620, n4619, n4618, n4617, n4616, n4615, n4614, n4613};
wire [12:0]I2_5_3;
assign I2_5_3 = {n4638, n4637, n4636, n4635, n4634, n4633, n4632, n4631, n4630, n4629, n4628, n4627, n4626};
wire [12:0]I3_5_3;
assign I3_5_3 = {n4651, n4650, n4649, n4648, n4647, n4646, n4645, n4644, n4643, n4642, n4641, n4640, n4639};
wire [12:0]I4_5_3;
assign I4_5_3 = {n4664, n4663, n4662, n4661, n4660, n4659, n4658, n4657, n4656, n4655, n4654, n4653, n4652};
wire [19:0]O_5_3;
assign {n4684, n4683, n4682, n4681, n4680, n4679, n4678, n4677, n4676, n4675, n4674, n4673, n4672, n4671, n4670, n4669, n4668, n4667, n4666, n4665} = O_5_3;

clb clb_5_3 ( .clk(clk_5_3), .reset(fpga_rst), .I4(I4_5_3), .I3(I3_5_3), .I2(I2_5_3), .I1(I1_5_3), .O(O_5_3), .config_in(config_chain[113755:111796]), .config_rst(config_rst) );

wire [0:0]clk_5_4;
assign clk_5_4 = {fpga_clk};
wire [12:0]I1_5_4;
assign I1_5_4 = {n4723, n4722, n4721, n4720, n4719, n4718, n4717, n4716, n4715, n4714, n4713, n4712, n4711};
wire [12:0]I2_5_4;
assign I2_5_4 = {n4736, n4735, n4734, n4733, n4732, n4731, n4730, n4729, n4728, n4727, n4726, n4725, n4724};
wire [12:0]I3_5_4;
assign I3_5_4 = {n4749, n4748, n4747, n4746, n4745, n4744, n4743, n4742, n4741, n4740, n4739, n4738, n4737};
wire [12:0]I4_5_4;
assign I4_5_4 = {n4762, n4761, n4760, n4759, n4758, n4757, n4756, n4755, n4754, n4753, n4752, n4751, n4750};
wire [19:0]O_5_4;
assign {n4782, n4781, n4780, n4779, n4778, n4777, n4776, n4775, n4774, n4773, n4772, n4771, n4770, n4769, n4768, n4767, n4766, n4765, n4764, n4763} = O_5_4;

clb clb_5_4 ( .clk(clk_5_4), .reset(fpga_rst), .I4(I4_5_4), .I3(I3_5_4), .I2(I2_5_4), .I1(I1_5_4), .O(O_5_4), .config_in(config_chain[115715:113756]), .config_rst(config_rst) );

wire [0:0]clk_5_5;
assign clk_5_5 = {fpga_clk};
wire [12:0]I1_5_5;
assign I1_5_5 = {n4821, n4820, n4819, n4818, n4817, n4816, n4815, n4814, n4813, n4812, n4811, n4810, n4809};
wire [12:0]I2_5_5;
assign I2_5_5 = {n4834, n4833, n4832, n4831, n4830, n4829, n4828, n4827, n4826, n4825, n4824, n4823, n4822};
wire [12:0]I3_5_5;
assign I3_5_5 = {n4847, n4846, n4845, n4844, n4843, n4842, n4841, n4840, n4839, n4838, n4837, n4836, n4835};
wire [12:0]I4_5_5;
assign I4_5_5 = {n4860, n4859, n4858, n4857, n4856, n4855, n4854, n4853, n4852, n4851, n4850, n4849, n4848};
wire [19:0]O_5_5;
assign {n4880, n4879, n4878, n4877, n4876, n4875, n4874, n4873, n4872, n4871, n4870, n4869, n4868, n4867, n4866, n4865, n4864, n4863, n4862, n4861} = O_5_5;

clb clb_5_5 ( .clk(clk_5_5), .reset(fpga_rst), .I4(I4_5_5), .I3(I3_5_5), .I2(I2_5_5), .I1(I1_5_5), .O(O_5_5), .config_in(config_chain[117675:115716]), .config_rst(config_rst) );

wire [0:0]clk_5_6;
assign clk_5_6 = {fpga_clk};
wire [12:0]I1_5_6;
assign I1_5_6 = {n4919, n4918, n4917, n4916, n4915, n4914, n4913, n4912, n4911, n4910, n4909, n4908, n4907};
wire [12:0]I2_5_6;
assign I2_5_6 = {n4932, n4931, n4930, n4929, n4928, n4927, n4926, n4925, n4924, n4923, n4922, n4921, n4920};
wire [12:0]I3_5_6;
assign I3_5_6 = {n4945, n4944, n4943, n4942, n4941, n4940, n4939, n4938, n4937, n4936, n4935, n4934, n4933};
wire [12:0]I4_5_6;
assign I4_5_6 = {n4958, n4957, n4956, n4955, n4954, n4953, n4952, n4951, n4950, n4949, n4948, n4947, n4946};
wire [19:0]O_5_6;
assign {n4978, n4977, n4976, n4975, n4974, n4973, n4972, n4971, n4970, n4969, n4968, n4967, n4966, n4965, n4964, n4963, n4962, n4961, n4960, n4959} = O_5_6;

clb clb_5_6 ( .clk(clk_5_6), .reset(fpga_rst), .I4(I4_5_6), .I3(I3_5_6), .I2(I2_5_6), .I1(I1_5_6), .O(O_5_6), .config_in(config_chain[119635:117676]), .config_rst(config_rst) );

wire [0:0]clk_5_7;
assign clk_5_7 = {fpga_clk};
wire [12:0]I1_5_7;
assign I1_5_7 = {n5017, n5016, n5015, n5014, n5013, n5012, n5011, n5010, n5009, n5008, n5007, n5006, n5005};
wire [12:0]I2_5_7;
assign I2_5_7 = {n5030, n5029, n5028, n5027, n5026, n5025, n5024, n5023, n5022, n5021, n5020, n5019, n5018};
wire [12:0]I3_5_7;
assign I3_5_7 = {n5043, n5042, n5041, n5040, n5039, n5038, n5037, n5036, n5035, n5034, n5033, n5032, n5031};
wire [12:0]I4_5_7;
assign I4_5_7 = {n5056, n5055, n5054, n5053, n5052, n5051, n5050, n5049, n5048, n5047, n5046, n5045, n5044};
wire [19:0]O_5_7;
assign {n5076, n5075, n5074, n5073, n5072, n5071, n5070, n5069, n5068, n5067, n5066, n5065, n5064, n5063, n5062, n5061, n5060, n5059, n5058, n5057} = O_5_7;

clb clb_5_7 ( .clk(clk_5_7), .reset(fpga_rst), .I4(I4_5_7), .I3(I3_5_7), .I2(I2_5_7), .I1(I1_5_7), .O(O_5_7), .config_in(config_chain[121595:119636]), .config_rst(config_rst) );

wire [0:0]clk_5_8;
assign clk_5_8 = {fpga_clk};
wire [12:0]I1_5_8;
assign I1_5_8 = {n5115, n5114, n5113, n5112, n5111, n5110, n5109, n5108, n5107, n5106, n5105, n5104, n5103};
wire [12:0]I2_5_8;
assign I2_5_8 = {n5128, n5127, n5126, n5125, n5124, n5123, n5122, n5121, n5120, n5119, n5118, n5117, n5116};
wire [12:0]I3_5_8;
assign I3_5_8 = {n5141, n5140, n5139, n5138, n5137, n5136, n5135, n5134, n5133, n5132, n5131, n5130, n5129};
wire [12:0]I4_5_8;
assign I4_5_8 = {n5154, n5153, n5152, n5151, n5150, n5149, n5148, n5147, n5146, n5145, n5144, n5143, n5142};
wire [19:0]O_5_8;
assign {n5174, n5173, n5172, n5171, n5170, n5169, n5168, n5167, n5166, n5165, n5164, n5163, n5162, n5161, n5160, n5159, n5158, n5157, n5156, n5155} = O_5_8;

clb clb_5_8 ( .clk(clk_5_8), .reset(fpga_rst), .I4(I4_5_8), .I3(I3_5_8), .I2(I2_5_8), .I1(I1_5_8), .O(O_5_8), .config_in(config_chain[123555:121596]), .config_rst(config_rst) );

wire [0:0]clk_5_9;
assign clk_5_9 = {fpga_clk};
wire [12:0]I1_5_9;
assign I1_5_9 = {n5213, n5212, n5211, n5210, n5209, n5208, n5207, n5206, n5205, n5204, n5203, n5202, n5201};
wire [12:0]I2_5_9;
assign I2_5_9 = {n5226, n5225, n5224, n5223, n5222, n5221, n5220, n5219, n5218, n5217, n5216, n5215, n5214};
wire [12:0]I3_5_9;
assign I3_5_9 = {n5239, n5238, n5237, n5236, n5235, n5234, n5233, n5232, n5231, n5230, n5229, n5228, n5227};
wire [12:0]I4_5_9;
assign I4_5_9 = {n5252, n5251, n5250, n5249, n5248, n5247, n5246, n5245, n5244, n5243, n5242, n5241, n5240};
wire [19:0]O_5_9;
assign {n5272, n5271, n5270, n5269, n5268, n5267, n5266, n5265, n5264, n5263, n5262, n5261, n5260, n5259, n5258, n5257, n5256, n5255, n5254, n5253} = O_5_9;

clb clb_5_9 ( .clk(clk_5_9), .reset(fpga_rst), .I4(I4_5_9), .I3(I3_5_9), .I2(I2_5_9), .I1(I1_5_9), .O(O_5_9), .config_in(config_chain[125515:123556]), .config_rst(config_rst) );

wire [7:0]outpad_5_10;
assign outpad_5_10 = {n5319, n5316, n5313, n5310, n5307, n5304, n5301, n5298};
wire [7:0]inpad_5_10;
assign {n5320, n5317, n5314, n5311, n5308, n5305, n5302, n5299} = inpad_5_10;

io io_5_10 ( .outpad(outpad_5_10), .inpad(inpad_5_10), .io_ext(io_5_10_wire), .config_in(config_chain[125523:125516]), .config_rst(config_rst) );

wire [7:0]outpad_6_0;
assign outpad_6_0 = {n5367, n5364, n5361, n5358, n5355, n5352, n5349, n5346};
wire [7:0]inpad_6_0;
assign {n5368, n5365, n5362, n5359, n5356, n5353, n5350, n5347} = inpad_6_0;

io io_6_0 ( .outpad(outpad_6_0), .inpad(inpad_6_0), .io_ext(io_6_0_wire), .config_in(config_chain[125531:125524]), .config_rst(config_rst) );

wire [0:0]clk_6_1;
assign clk_6_1 = {fpga_clk};
wire [12:0]I1_6_1;
assign I1_6_1 = {n5407, n5406, n5405, n5404, n5403, n5402, n5401, n5400, n5399, n5398, n5397, n5396, n5395};
wire [12:0]I2_6_1;
assign I2_6_1 = {n5420, n5419, n5418, n5417, n5416, n5415, n5414, n5413, n5412, n5411, n5410, n5409, n5408};
wire [12:0]I3_6_1;
assign I3_6_1 = {n5433, n5432, n5431, n5430, n5429, n5428, n5427, n5426, n5425, n5424, n5423, n5422, n5421};
wire [12:0]I4_6_1;
assign I4_6_1 = {n5446, n5445, n5444, n5443, n5442, n5441, n5440, n5439, n5438, n5437, n5436, n5435, n5434};
wire [19:0]O_6_1;
assign {n5466, n5465, n5464, n5463, n5462, n5461, n5460, n5459, n5458, n5457, n5456, n5455, n5454, n5453, n5452, n5451, n5450, n5449, n5448, n5447} = O_6_1;

clb clb_6_1 ( .clk(clk_6_1), .reset(fpga_rst), .I4(I4_6_1), .I3(I3_6_1), .I2(I2_6_1), .I1(I1_6_1), .O(O_6_1), .config_in(config_chain[127491:125532]), .config_rst(config_rst) );

wire [0:0]clk_6_2;
assign clk_6_2 = {fpga_clk};
wire [12:0]I1_6_2;
assign I1_6_2 = {n5505, n5504, n5503, n5502, n5501, n5500, n5499, n5498, n5497, n5496, n5495, n5494, n5493};
wire [12:0]I2_6_2;
assign I2_6_2 = {n5518, n5517, n5516, n5515, n5514, n5513, n5512, n5511, n5510, n5509, n5508, n5507, n5506};
wire [12:0]I3_6_2;
assign I3_6_2 = {n5531, n5530, n5529, n5528, n5527, n5526, n5525, n5524, n5523, n5522, n5521, n5520, n5519};
wire [12:0]I4_6_2;
assign I4_6_2 = {n5544, n5543, n5542, n5541, n5540, n5539, n5538, n5537, n5536, n5535, n5534, n5533, n5532};
wire [19:0]O_6_2;
assign {n5564, n5563, n5562, n5561, n5560, n5559, n5558, n5557, n5556, n5555, n5554, n5553, n5552, n5551, n5550, n5549, n5548, n5547, n5546, n5545} = O_6_2;

clb clb_6_2 ( .clk(clk_6_2), .reset(fpga_rst), .I4(I4_6_2), .I3(I3_6_2), .I2(I2_6_2), .I1(I1_6_2), .O(O_6_2), .config_in(config_chain[129451:127492]), .config_rst(config_rst) );

wire [0:0]clk_6_3;
assign clk_6_3 = {fpga_clk};
wire [12:0]I1_6_3;
assign I1_6_3 = {n5603, n5602, n5601, n5600, n5599, n5598, n5597, n5596, n5595, n5594, n5593, n5592, n5591};
wire [12:0]I2_6_3;
assign I2_6_3 = {n5616, n5615, n5614, n5613, n5612, n5611, n5610, n5609, n5608, n5607, n5606, n5605, n5604};
wire [12:0]I3_6_3;
assign I3_6_3 = {n5629, n5628, n5627, n5626, n5625, n5624, n5623, n5622, n5621, n5620, n5619, n5618, n5617};
wire [12:0]I4_6_3;
assign I4_6_3 = {n5642, n5641, n5640, n5639, n5638, n5637, n5636, n5635, n5634, n5633, n5632, n5631, n5630};
wire [19:0]O_6_3;
assign {n5662, n5661, n5660, n5659, n5658, n5657, n5656, n5655, n5654, n5653, n5652, n5651, n5650, n5649, n5648, n5647, n5646, n5645, n5644, n5643} = O_6_3;

clb clb_6_3 ( .clk(clk_6_3), .reset(fpga_rst), .I4(I4_6_3), .I3(I3_6_3), .I2(I2_6_3), .I1(I1_6_3), .O(O_6_3), .config_in(config_chain[131411:129452]), .config_rst(config_rst) );

wire [0:0]clk_6_4;
assign clk_6_4 = {fpga_clk};
wire [12:0]I1_6_4;
assign I1_6_4 = {n5701, n5700, n5699, n5698, n5697, n5696, n5695, n5694, n5693, n5692, n5691, n5690, n5689};
wire [12:0]I2_6_4;
assign I2_6_4 = {n5714, n5713, n5712, n5711, n5710, n5709, n5708, n5707, n5706, n5705, n5704, n5703, n5702};
wire [12:0]I3_6_4;
assign I3_6_4 = {n5727, n5726, n5725, n5724, n5723, n5722, n5721, n5720, n5719, n5718, n5717, n5716, n5715};
wire [12:0]I4_6_4;
assign I4_6_4 = {n5740, n5739, n5738, n5737, n5736, n5735, n5734, n5733, n5732, n5731, n5730, n5729, n5728};
wire [19:0]O_6_4;
assign {n5760, n5759, n5758, n5757, n5756, n5755, n5754, n5753, n5752, n5751, n5750, n5749, n5748, n5747, n5746, n5745, n5744, n5743, n5742, n5741} = O_6_4;

clb clb_6_4 ( .clk(clk_6_4), .reset(fpga_rst), .I4(I4_6_4), .I3(I3_6_4), .I2(I2_6_4), .I1(I1_6_4), .O(O_6_4), .config_in(config_chain[133371:131412]), .config_rst(config_rst) );

wire [0:0]clk_6_5;
assign clk_6_5 = {fpga_clk};
wire [12:0]I1_6_5;
assign I1_6_5 = {n5799, n5798, n5797, n5796, n5795, n5794, n5793, n5792, n5791, n5790, n5789, n5788, n5787};
wire [12:0]I2_6_5;
assign I2_6_5 = {n5812, n5811, n5810, n5809, n5808, n5807, n5806, n5805, n5804, n5803, n5802, n5801, n5800};
wire [12:0]I3_6_5;
assign I3_6_5 = {n5825, n5824, n5823, n5822, n5821, n5820, n5819, n5818, n5817, n5816, n5815, n5814, n5813};
wire [12:0]I4_6_5;
assign I4_6_5 = {n5838, n5837, n5836, n5835, n5834, n5833, n5832, n5831, n5830, n5829, n5828, n5827, n5826};
wire [19:0]O_6_5;
assign {n5858, n5857, n5856, n5855, n5854, n5853, n5852, n5851, n5850, n5849, n5848, n5847, n5846, n5845, n5844, n5843, n5842, n5841, n5840, n5839} = O_6_5;

clb clb_6_5 ( .clk(clk_6_5), .reset(fpga_rst), .I4(I4_6_5), .I3(I3_6_5), .I2(I2_6_5), .I1(I1_6_5), .O(O_6_5), .config_in(config_chain[135331:133372]), .config_rst(config_rst) );

wire [0:0]clk_6_6;
assign clk_6_6 = {fpga_clk};
wire [12:0]I1_6_6;
assign I1_6_6 = {n5897, n5896, n5895, n5894, n5893, n5892, n5891, n5890, n5889, n5888, n5887, n5886, n5885};
wire [12:0]I2_6_6;
assign I2_6_6 = {n5910, n5909, n5908, n5907, n5906, n5905, n5904, n5903, n5902, n5901, n5900, n5899, n5898};
wire [12:0]I3_6_6;
assign I3_6_6 = {n5923, n5922, n5921, n5920, n5919, n5918, n5917, n5916, n5915, n5914, n5913, n5912, n5911};
wire [12:0]I4_6_6;
assign I4_6_6 = {n5936, n5935, n5934, n5933, n5932, n5931, n5930, n5929, n5928, n5927, n5926, n5925, n5924};
wire [19:0]O_6_6;
assign {n5956, n5955, n5954, n5953, n5952, n5951, n5950, n5949, n5948, n5947, n5946, n5945, n5944, n5943, n5942, n5941, n5940, n5939, n5938, n5937} = O_6_6;

clb clb_6_6 ( .clk(clk_6_6), .reset(fpga_rst), .I4(I4_6_6), .I3(I3_6_6), .I2(I2_6_6), .I1(I1_6_6), .O(O_6_6), .config_in(config_chain[137291:135332]), .config_rst(config_rst) );

wire [0:0]clk_6_7;
assign clk_6_7 = {fpga_clk};
wire [12:0]I1_6_7;
assign I1_6_7 = {n5995, n5994, n5993, n5992, n5991, n5990, n5989, n5988, n5987, n5986, n5985, n5984, n5983};
wire [12:0]I2_6_7;
assign I2_6_7 = {n6008, n6007, n6006, n6005, n6004, n6003, n6002, n6001, n6000, n5999, n5998, n5997, n5996};
wire [12:0]I3_6_7;
assign I3_6_7 = {n6021, n6020, n6019, n6018, n6017, n6016, n6015, n6014, n6013, n6012, n6011, n6010, n6009};
wire [12:0]I4_6_7;
assign I4_6_7 = {n6034, n6033, n6032, n6031, n6030, n6029, n6028, n6027, n6026, n6025, n6024, n6023, n6022};
wire [19:0]O_6_7;
assign {n6054, n6053, n6052, n6051, n6050, n6049, n6048, n6047, n6046, n6045, n6044, n6043, n6042, n6041, n6040, n6039, n6038, n6037, n6036, n6035} = O_6_7;

clb clb_6_7 ( .clk(clk_6_7), .reset(fpga_rst), .I4(I4_6_7), .I3(I3_6_7), .I2(I2_6_7), .I1(I1_6_7), .O(O_6_7), .config_in(config_chain[139251:137292]), .config_rst(config_rst) );

wire [0:0]clk_6_8;
assign clk_6_8 = {fpga_clk};
wire [12:0]I1_6_8;
assign I1_6_8 = {n6093, n6092, n6091, n6090, n6089, n6088, n6087, n6086, n6085, n6084, n6083, n6082, n6081};
wire [12:0]I2_6_8;
assign I2_6_8 = {n6106, n6105, n6104, n6103, n6102, n6101, n6100, n6099, n6098, n6097, n6096, n6095, n6094};
wire [12:0]I3_6_8;
assign I3_6_8 = {n6119, n6118, n6117, n6116, n6115, n6114, n6113, n6112, n6111, n6110, n6109, n6108, n6107};
wire [12:0]I4_6_8;
assign I4_6_8 = {n6132, n6131, n6130, n6129, n6128, n6127, n6126, n6125, n6124, n6123, n6122, n6121, n6120};
wire [19:0]O_6_8;
assign {n6152, n6151, n6150, n6149, n6148, n6147, n6146, n6145, n6144, n6143, n6142, n6141, n6140, n6139, n6138, n6137, n6136, n6135, n6134, n6133} = O_6_8;

clb clb_6_8 ( .clk(clk_6_8), .reset(fpga_rst), .I4(I4_6_8), .I3(I3_6_8), .I2(I2_6_8), .I1(I1_6_8), .O(O_6_8), .config_in(config_chain[141211:139252]), .config_rst(config_rst) );

wire [0:0]clk_6_9;
assign clk_6_9 = {fpga_clk};
wire [12:0]I1_6_9;
assign I1_6_9 = {n6191, n6190, n6189, n6188, n6187, n6186, n6185, n6184, n6183, n6182, n6181, n6180, n6179};
wire [12:0]I2_6_9;
assign I2_6_9 = {n6204, n6203, n6202, n6201, n6200, n6199, n6198, n6197, n6196, n6195, n6194, n6193, n6192};
wire [12:0]I3_6_9;
assign I3_6_9 = {n6217, n6216, n6215, n6214, n6213, n6212, n6211, n6210, n6209, n6208, n6207, n6206, n6205};
wire [12:0]I4_6_9;
assign I4_6_9 = {n6230, n6229, n6228, n6227, n6226, n6225, n6224, n6223, n6222, n6221, n6220, n6219, n6218};
wire [19:0]O_6_9;
assign {n6250, n6249, n6248, n6247, n6246, n6245, n6244, n6243, n6242, n6241, n6240, n6239, n6238, n6237, n6236, n6235, n6234, n6233, n6232, n6231} = O_6_9;

clb clb_6_9 ( .clk(clk_6_9), .reset(fpga_rst), .I4(I4_6_9), .I3(I3_6_9), .I2(I2_6_9), .I1(I1_6_9), .O(O_6_9), .config_in(config_chain[143171:141212]), .config_rst(config_rst) );

wire [7:0]outpad_6_10;
assign outpad_6_10 = {n6297, n6294, n6291, n6288, n6285, n6282, n6279, n6276};
wire [7:0]inpad_6_10;
assign {n6298, n6295, n6292, n6289, n6286, n6283, n6280, n6277} = inpad_6_10;

io io_6_10 ( .outpad(outpad_6_10), .inpad(inpad_6_10), .io_ext(io_6_10_wire), .config_in(config_chain[143179:143172]), .config_rst(config_rst) );

wire [7:0]outpad_7_0;
assign outpad_7_0 = {n6345, n6342, n6339, n6336, n6333, n6330, n6327, n6324};
wire [7:0]inpad_7_0;
assign {n6346, n6343, n6340, n6337, n6334, n6331, n6328, n6325} = inpad_7_0;

io io_7_0 ( .outpad(outpad_7_0), .inpad(inpad_7_0), .io_ext(io_7_0_wire), .config_in(config_chain[143187:143180]), .config_rst(config_rst) );

wire [0:0]clk_7_1;
assign clk_7_1 = {fpga_clk};
wire [12:0]I1_7_1;
assign I1_7_1 = {n6385, n6384, n6383, n6382, n6381, n6380, n6379, n6378, n6377, n6376, n6375, n6374, n6373};
wire [12:0]I2_7_1;
assign I2_7_1 = {n6398, n6397, n6396, n6395, n6394, n6393, n6392, n6391, n6390, n6389, n6388, n6387, n6386};
wire [12:0]I3_7_1;
assign I3_7_1 = {n6411, n6410, n6409, n6408, n6407, n6406, n6405, n6404, n6403, n6402, n6401, n6400, n6399};
wire [12:0]I4_7_1;
assign I4_7_1 = {n6424, n6423, n6422, n6421, n6420, n6419, n6418, n6417, n6416, n6415, n6414, n6413, n6412};
wire [19:0]O_7_1;
assign {n6444, n6443, n6442, n6441, n6440, n6439, n6438, n6437, n6436, n6435, n6434, n6433, n6432, n6431, n6430, n6429, n6428, n6427, n6426, n6425} = O_7_1;

clb clb_7_1 ( .clk(clk_7_1), .reset(fpga_rst), .I4(I4_7_1), .I3(I3_7_1), .I2(I2_7_1), .I1(I1_7_1), .O(O_7_1), .config_in(config_chain[145147:143188]), .config_rst(config_rst) );

wire [0:0]clk_7_2;
assign clk_7_2 = {fpga_clk};
wire [12:0]I1_7_2;
assign I1_7_2 = {n6483, n6482, n6481, n6480, n6479, n6478, n6477, n6476, n6475, n6474, n6473, n6472, n6471};
wire [12:0]I2_7_2;
assign I2_7_2 = {n6496, n6495, n6494, n6493, n6492, n6491, n6490, n6489, n6488, n6487, n6486, n6485, n6484};
wire [12:0]I3_7_2;
assign I3_7_2 = {n6509, n6508, n6507, n6506, n6505, n6504, n6503, n6502, n6501, n6500, n6499, n6498, n6497};
wire [12:0]I4_7_2;
assign I4_7_2 = {n6522, n6521, n6520, n6519, n6518, n6517, n6516, n6515, n6514, n6513, n6512, n6511, n6510};
wire [19:0]O_7_2;
assign {n6542, n6541, n6540, n6539, n6538, n6537, n6536, n6535, n6534, n6533, n6532, n6531, n6530, n6529, n6528, n6527, n6526, n6525, n6524, n6523} = O_7_2;

clb clb_7_2 ( .clk(clk_7_2), .reset(fpga_rst), .I4(I4_7_2), .I3(I3_7_2), .I2(I2_7_2), .I1(I1_7_2), .O(O_7_2), .config_in(config_chain[147107:145148]), .config_rst(config_rst) );

wire [0:0]clk_7_3;
assign clk_7_3 = {fpga_clk};
wire [12:0]I1_7_3;
assign I1_7_3 = {n6581, n6580, n6579, n6578, n6577, n6576, n6575, n6574, n6573, n6572, n6571, n6570, n6569};
wire [12:0]I2_7_3;
assign I2_7_3 = {n6594, n6593, n6592, n6591, n6590, n6589, n6588, n6587, n6586, n6585, n6584, n6583, n6582};
wire [12:0]I3_7_3;
assign I3_7_3 = {n6607, n6606, n6605, n6604, n6603, n6602, n6601, n6600, n6599, n6598, n6597, n6596, n6595};
wire [12:0]I4_7_3;
assign I4_7_3 = {n6620, n6619, n6618, n6617, n6616, n6615, n6614, n6613, n6612, n6611, n6610, n6609, n6608};
wire [19:0]O_7_3;
assign {n6640, n6639, n6638, n6637, n6636, n6635, n6634, n6633, n6632, n6631, n6630, n6629, n6628, n6627, n6626, n6625, n6624, n6623, n6622, n6621} = O_7_3;

clb clb_7_3 ( .clk(clk_7_3), .reset(fpga_rst), .I4(I4_7_3), .I3(I3_7_3), .I2(I2_7_3), .I1(I1_7_3), .O(O_7_3), .config_in(config_chain[149067:147108]), .config_rst(config_rst) );

wire [0:0]clk_7_4;
assign clk_7_4 = {fpga_clk};
wire [12:0]I1_7_4;
assign I1_7_4 = {n6679, n6678, n6677, n6676, n6675, n6674, n6673, n6672, n6671, n6670, n6669, n6668, n6667};
wire [12:0]I2_7_4;
assign I2_7_4 = {n6692, n6691, n6690, n6689, n6688, n6687, n6686, n6685, n6684, n6683, n6682, n6681, n6680};
wire [12:0]I3_7_4;
assign I3_7_4 = {n6705, n6704, n6703, n6702, n6701, n6700, n6699, n6698, n6697, n6696, n6695, n6694, n6693};
wire [12:0]I4_7_4;
assign I4_7_4 = {n6718, n6717, n6716, n6715, n6714, n6713, n6712, n6711, n6710, n6709, n6708, n6707, n6706};
wire [19:0]O_7_4;
assign {n6738, n6737, n6736, n6735, n6734, n6733, n6732, n6731, n6730, n6729, n6728, n6727, n6726, n6725, n6724, n6723, n6722, n6721, n6720, n6719} = O_7_4;

clb clb_7_4 ( .clk(clk_7_4), .reset(fpga_rst), .I4(I4_7_4), .I3(I3_7_4), .I2(I2_7_4), .I1(I1_7_4), .O(O_7_4), .config_in(config_chain[151027:149068]), .config_rst(config_rst) );

wire [0:0]clk_7_5;
assign clk_7_5 = {fpga_clk};
wire [12:0]I1_7_5;
assign I1_7_5 = {n6777, n6776, n6775, n6774, n6773, n6772, n6771, n6770, n6769, n6768, n6767, n6766, n6765};
wire [12:0]I2_7_5;
assign I2_7_5 = {n6790, n6789, n6788, n6787, n6786, n6785, n6784, n6783, n6782, n6781, n6780, n6779, n6778};
wire [12:0]I3_7_5;
assign I3_7_5 = {n6803, n6802, n6801, n6800, n6799, n6798, n6797, n6796, n6795, n6794, n6793, n6792, n6791};
wire [12:0]I4_7_5;
assign I4_7_5 = {n6816, n6815, n6814, n6813, n6812, n6811, n6810, n6809, n6808, n6807, n6806, n6805, n6804};
wire [19:0]O_7_5;
assign {n6836, n6835, n6834, n6833, n6832, n6831, n6830, n6829, n6828, n6827, n6826, n6825, n6824, n6823, n6822, n6821, n6820, n6819, n6818, n6817} = O_7_5;

clb clb_7_5 ( .clk(clk_7_5), .reset(fpga_rst), .I4(I4_7_5), .I3(I3_7_5), .I2(I2_7_5), .I1(I1_7_5), .O(O_7_5), .config_in(config_chain[152987:151028]), .config_rst(config_rst) );

wire [0:0]clk_7_6;
assign clk_7_6 = {fpga_clk};
wire [12:0]I1_7_6;
assign I1_7_6 = {n6875, n6874, n6873, n6872, n6871, n6870, n6869, n6868, n6867, n6866, n6865, n6864, n6863};
wire [12:0]I2_7_6;
assign I2_7_6 = {n6888, n6887, n6886, n6885, n6884, n6883, n6882, n6881, n6880, n6879, n6878, n6877, n6876};
wire [12:0]I3_7_6;
assign I3_7_6 = {n6901, n6900, n6899, n6898, n6897, n6896, n6895, n6894, n6893, n6892, n6891, n6890, n6889};
wire [12:0]I4_7_6;
assign I4_7_6 = {n6914, n6913, n6912, n6911, n6910, n6909, n6908, n6907, n6906, n6905, n6904, n6903, n6902};
wire [19:0]O_7_6;
assign {n6934, n6933, n6932, n6931, n6930, n6929, n6928, n6927, n6926, n6925, n6924, n6923, n6922, n6921, n6920, n6919, n6918, n6917, n6916, n6915} = O_7_6;

clb clb_7_6 ( .clk(clk_7_6), .reset(fpga_rst), .I4(I4_7_6), .I3(I3_7_6), .I2(I2_7_6), .I1(I1_7_6), .O(O_7_6), .config_in(config_chain[154947:152988]), .config_rst(config_rst) );

wire [0:0]clk_7_7;
assign clk_7_7 = {fpga_clk};
wire [12:0]I1_7_7;
assign I1_7_7 = {n6973, n6972, n6971, n6970, n6969, n6968, n6967, n6966, n6965, n6964, n6963, n6962, n6961};
wire [12:0]I2_7_7;
assign I2_7_7 = {n6986, n6985, n6984, n6983, n6982, n6981, n6980, n6979, n6978, n6977, n6976, n6975, n6974};
wire [12:0]I3_7_7;
assign I3_7_7 = {n6999, n6998, n6997, n6996, n6995, n6994, n6993, n6992, n6991, n6990, n6989, n6988, n6987};
wire [12:0]I4_7_7;
assign I4_7_7 = {n7012, n7011, n7010, n7009, n7008, n7007, n7006, n7005, n7004, n7003, n7002, n7001, n7000};
wire [19:0]O_7_7;
assign {n7032, n7031, n7030, n7029, n7028, n7027, n7026, n7025, n7024, n7023, n7022, n7021, n7020, n7019, n7018, n7017, n7016, n7015, n7014, n7013} = O_7_7;

clb clb_7_7 ( .clk(clk_7_7), .reset(fpga_rst), .I4(I4_7_7), .I3(I3_7_7), .I2(I2_7_7), .I1(I1_7_7), .O(O_7_7), .config_in(config_chain[156907:154948]), .config_rst(config_rst) );

wire [0:0]clk_7_8;
assign clk_7_8 = {fpga_clk};
wire [12:0]I1_7_8;
assign I1_7_8 = {n7071, n7070, n7069, n7068, n7067, n7066, n7065, n7064, n7063, n7062, n7061, n7060, n7059};
wire [12:0]I2_7_8;
assign I2_7_8 = {n7084, n7083, n7082, n7081, n7080, n7079, n7078, n7077, n7076, n7075, n7074, n7073, n7072};
wire [12:0]I3_7_8;
assign I3_7_8 = {n7097, n7096, n7095, n7094, n7093, n7092, n7091, n7090, n7089, n7088, n7087, n7086, n7085};
wire [12:0]I4_7_8;
assign I4_7_8 = {n7110, n7109, n7108, n7107, n7106, n7105, n7104, n7103, n7102, n7101, n7100, n7099, n7098};
wire [19:0]O_7_8;
assign {n7130, n7129, n7128, n7127, n7126, n7125, n7124, n7123, n7122, n7121, n7120, n7119, n7118, n7117, n7116, n7115, n7114, n7113, n7112, n7111} = O_7_8;

clb clb_7_8 ( .clk(clk_7_8), .reset(fpga_rst), .I4(I4_7_8), .I3(I3_7_8), .I2(I2_7_8), .I1(I1_7_8), .O(O_7_8), .config_in(config_chain[158867:156908]), .config_rst(config_rst) );

wire [0:0]clk_7_9;
assign clk_7_9 = {fpga_clk};
wire [12:0]I1_7_9;
assign I1_7_9 = {n7169, n7168, n7167, n7166, n7165, n7164, n7163, n7162, n7161, n7160, n7159, n7158, n7157};
wire [12:0]I2_7_9;
assign I2_7_9 = {n7182, n7181, n7180, n7179, n7178, n7177, n7176, n7175, n7174, n7173, n7172, n7171, n7170};
wire [12:0]I3_7_9;
assign I3_7_9 = {n7195, n7194, n7193, n7192, n7191, n7190, n7189, n7188, n7187, n7186, n7185, n7184, n7183};
wire [12:0]I4_7_9;
assign I4_7_9 = {n7208, n7207, n7206, n7205, n7204, n7203, n7202, n7201, n7200, n7199, n7198, n7197, n7196};
wire [19:0]O_7_9;
assign {n7228, n7227, n7226, n7225, n7224, n7223, n7222, n7221, n7220, n7219, n7218, n7217, n7216, n7215, n7214, n7213, n7212, n7211, n7210, n7209} = O_7_9;

clb clb_7_9 ( .clk(clk_7_9), .reset(fpga_rst), .I4(I4_7_9), .I3(I3_7_9), .I2(I2_7_9), .I1(I1_7_9), .O(O_7_9), .config_in(config_chain[160827:158868]), .config_rst(config_rst) );

wire [7:0]outpad_7_10;
assign outpad_7_10 = {n7275, n7272, n7269, n7266, n7263, n7260, n7257, n7254};
wire [7:0]inpad_7_10;
assign {n7276, n7273, n7270, n7267, n7264, n7261, n7258, n7255} = inpad_7_10;

io io_7_10 ( .outpad(outpad_7_10), .inpad(inpad_7_10), .io_ext(io_7_10_wire), .config_in(config_chain[160835:160828]), .config_rst(config_rst) );

wire [7:0]outpad_8_0;
assign outpad_8_0 = {n7323, n7320, n7317, n7314, n7311, n7308, n7305, n7302};
wire [7:0]inpad_8_0;
assign {n7324, n7321, n7318, n7315, n7312, n7309, n7306, n7303} = inpad_8_0;

io io_8_0 ( .outpad(outpad_8_0), .inpad(inpad_8_0), .io_ext(io_8_0_wire), .config_in(config_chain[160843:160836]), .config_rst(config_rst) );

wire [0:0]clk_8_1;
assign clk_8_1 = {fpga_clk};
wire [12:0]I1_8_1;
assign I1_8_1 = {n7363, n7362, n7361, n7360, n7359, n7358, n7357, n7356, n7355, n7354, n7353, n7352, n7351};
wire [12:0]I2_8_1;
assign I2_8_1 = {n7376, n7375, n7374, n7373, n7372, n7371, n7370, n7369, n7368, n7367, n7366, n7365, n7364};
wire [12:0]I3_8_1;
assign I3_8_1 = {n7389, n7388, n7387, n7386, n7385, n7384, n7383, n7382, n7381, n7380, n7379, n7378, n7377};
wire [12:0]I4_8_1;
assign I4_8_1 = {n7402, n7401, n7400, n7399, n7398, n7397, n7396, n7395, n7394, n7393, n7392, n7391, n7390};
wire [19:0]O_8_1;
assign {n7422, n7421, n7420, n7419, n7418, n7417, n7416, n7415, n7414, n7413, n7412, n7411, n7410, n7409, n7408, n7407, n7406, n7405, n7404, n7403} = O_8_1;

clb clb_8_1 ( .clk(clk_8_1), .reset(fpga_rst), .I4(I4_8_1), .I3(I3_8_1), .I2(I2_8_1), .I1(I1_8_1), .O(O_8_1), .config_in(config_chain[162803:160844]), .config_rst(config_rst) );

wire [0:0]clk_8_2;
assign clk_8_2 = {fpga_clk};
wire [12:0]I1_8_2;
assign I1_8_2 = {n7461, n7460, n7459, n7458, n7457, n7456, n7455, n7454, n7453, n7452, n7451, n7450, n7449};
wire [12:0]I2_8_2;
assign I2_8_2 = {n7474, n7473, n7472, n7471, n7470, n7469, n7468, n7467, n7466, n7465, n7464, n7463, n7462};
wire [12:0]I3_8_2;
assign I3_8_2 = {n7487, n7486, n7485, n7484, n7483, n7482, n7481, n7480, n7479, n7478, n7477, n7476, n7475};
wire [12:0]I4_8_2;
assign I4_8_2 = {n7500, n7499, n7498, n7497, n7496, n7495, n7494, n7493, n7492, n7491, n7490, n7489, n7488};
wire [19:0]O_8_2;
assign {n7520, n7519, n7518, n7517, n7516, n7515, n7514, n7513, n7512, n7511, n7510, n7509, n7508, n7507, n7506, n7505, n7504, n7503, n7502, n7501} = O_8_2;

clb clb_8_2 ( .clk(clk_8_2), .reset(fpga_rst), .I4(I4_8_2), .I3(I3_8_2), .I2(I2_8_2), .I1(I1_8_2), .O(O_8_2), .config_in(config_chain[164763:162804]), .config_rst(config_rst) );

wire [0:0]clk_8_3;
assign clk_8_3 = {fpga_clk};
wire [12:0]I1_8_3;
assign I1_8_3 = {n7559, n7558, n7557, n7556, n7555, n7554, n7553, n7552, n7551, n7550, n7549, n7548, n7547};
wire [12:0]I2_8_3;
assign I2_8_3 = {n7572, n7571, n7570, n7569, n7568, n7567, n7566, n7565, n7564, n7563, n7562, n7561, n7560};
wire [12:0]I3_8_3;
assign I3_8_3 = {n7585, n7584, n7583, n7582, n7581, n7580, n7579, n7578, n7577, n7576, n7575, n7574, n7573};
wire [12:0]I4_8_3;
assign I4_8_3 = {n7598, n7597, n7596, n7595, n7594, n7593, n7592, n7591, n7590, n7589, n7588, n7587, n7586};
wire [19:0]O_8_3;
assign {n7618, n7617, n7616, n7615, n7614, n7613, n7612, n7611, n7610, n7609, n7608, n7607, n7606, n7605, n7604, n7603, n7602, n7601, n7600, n7599} = O_8_3;

clb clb_8_3 ( .clk(clk_8_3), .reset(fpga_rst), .I4(I4_8_3), .I3(I3_8_3), .I2(I2_8_3), .I1(I1_8_3), .O(O_8_3), .config_in(config_chain[166723:164764]), .config_rst(config_rst) );

wire [0:0]clk_8_4;
assign clk_8_4 = {fpga_clk};
wire [12:0]I1_8_4;
assign I1_8_4 = {n7657, n7656, n7655, n7654, n7653, n7652, n7651, n7650, n7649, n7648, n7647, n7646, n7645};
wire [12:0]I2_8_4;
assign I2_8_4 = {n7670, n7669, n7668, n7667, n7666, n7665, n7664, n7663, n7662, n7661, n7660, n7659, n7658};
wire [12:0]I3_8_4;
assign I3_8_4 = {n7683, n7682, n7681, n7680, n7679, n7678, n7677, n7676, n7675, n7674, n7673, n7672, n7671};
wire [12:0]I4_8_4;
assign I4_8_4 = {n7696, n7695, n7694, n7693, n7692, n7691, n7690, n7689, n7688, n7687, n7686, n7685, n7684};
wire [19:0]O_8_4;
assign {n7716, n7715, n7714, n7713, n7712, n7711, n7710, n7709, n7708, n7707, n7706, n7705, n7704, n7703, n7702, n7701, n7700, n7699, n7698, n7697} = O_8_4;

clb clb_8_4 ( .clk(clk_8_4), .reset(fpga_rst), .I4(I4_8_4), .I3(I3_8_4), .I2(I2_8_4), .I1(I1_8_4), .O(O_8_4), .config_in(config_chain[168683:166724]), .config_rst(config_rst) );

wire [0:0]clk_8_5;
assign clk_8_5 = {fpga_clk};
wire [12:0]I1_8_5;
assign I1_8_5 = {n7755, n7754, n7753, n7752, n7751, n7750, n7749, n7748, n7747, n7746, n7745, n7744, n7743};
wire [12:0]I2_8_5;
assign I2_8_5 = {n7768, n7767, n7766, n7765, n7764, n7763, n7762, n7761, n7760, n7759, n7758, n7757, n7756};
wire [12:0]I3_8_5;
assign I3_8_5 = {n7781, n7780, n7779, n7778, n7777, n7776, n7775, n7774, n7773, n7772, n7771, n7770, n7769};
wire [12:0]I4_8_5;
assign I4_8_5 = {n7794, n7793, n7792, n7791, n7790, n7789, n7788, n7787, n7786, n7785, n7784, n7783, n7782};
wire [19:0]O_8_5;
assign {n7814, n7813, n7812, n7811, n7810, n7809, n7808, n7807, n7806, n7805, n7804, n7803, n7802, n7801, n7800, n7799, n7798, n7797, n7796, n7795} = O_8_5;

clb clb_8_5 ( .clk(clk_8_5), .reset(fpga_rst), .I4(I4_8_5), .I3(I3_8_5), .I2(I2_8_5), .I1(I1_8_5), .O(O_8_5), .config_in(config_chain[170643:168684]), .config_rst(config_rst) );

wire [0:0]clk_8_6;
assign clk_8_6 = {fpga_clk};
wire [12:0]I1_8_6;
assign I1_8_6 = {n7853, n7852, n7851, n7850, n7849, n7848, n7847, n7846, n7845, n7844, n7843, n7842, n7841};
wire [12:0]I2_8_6;
assign I2_8_6 = {n7866, n7865, n7864, n7863, n7862, n7861, n7860, n7859, n7858, n7857, n7856, n7855, n7854};
wire [12:0]I3_8_6;
assign I3_8_6 = {n7879, n7878, n7877, n7876, n7875, n7874, n7873, n7872, n7871, n7870, n7869, n7868, n7867};
wire [12:0]I4_8_6;
assign I4_8_6 = {n7892, n7891, n7890, n7889, n7888, n7887, n7886, n7885, n7884, n7883, n7882, n7881, n7880};
wire [19:0]O_8_6;
assign {n7912, n7911, n7910, n7909, n7908, n7907, n7906, n7905, n7904, n7903, n7902, n7901, n7900, n7899, n7898, n7897, n7896, n7895, n7894, n7893} = O_8_6;

clb clb_8_6 ( .clk(clk_8_6), .reset(fpga_rst), .I4(I4_8_6), .I3(I3_8_6), .I2(I2_8_6), .I1(I1_8_6), .O(O_8_6), .config_in(config_chain[172603:170644]), .config_rst(config_rst) );

wire [0:0]clk_8_7;
assign clk_8_7 = {fpga_clk};
wire [12:0]I1_8_7;
assign I1_8_7 = {n7951, n7950, n7949, n7948, n7947, n7946, n7945, n7944, n7943, n7942, n7941, n7940, n7939};
wire [12:0]I2_8_7;
assign I2_8_7 = {n7964, n7963, n7962, n7961, n7960, n7959, n7958, n7957, n7956, n7955, n7954, n7953, n7952};
wire [12:0]I3_8_7;
assign I3_8_7 = {n7977, n7976, n7975, n7974, n7973, n7972, n7971, n7970, n7969, n7968, n7967, n7966, n7965};
wire [12:0]I4_8_7;
assign I4_8_7 = {n7990, n7989, n7988, n7987, n7986, n7985, n7984, n7983, n7982, n7981, n7980, n7979, n7978};
wire [19:0]O_8_7;
assign {n8010, n8009, n8008, n8007, n8006, n8005, n8004, n8003, n8002, n8001, n8000, n7999, n7998, n7997, n7996, n7995, n7994, n7993, n7992, n7991} = O_8_7;

clb clb_8_7 ( .clk(clk_8_7), .reset(fpga_rst), .I4(I4_8_7), .I3(I3_8_7), .I2(I2_8_7), .I1(I1_8_7), .O(O_8_7), .config_in(config_chain[174563:172604]), .config_rst(config_rst) );

wire [0:0]clk_8_8;
assign clk_8_8 = {fpga_clk};
wire [12:0]I1_8_8;
assign I1_8_8 = {n8049, n8048, n8047, n8046, n8045, n8044, n8043, n8042, n8041, n8040, n8039, n8038, n8037};
wire [12:0]I2_8_8;
assign I2_8_8 = {n8062, n8061, n8060, n8059, n8058, n8057, n8056, n8055, n8054, n8053, n8052, n8051, n8050};
wire [12:0]I3_8_8;
assign I3_8_8 = {n8075, n8074, n8073, n8072, n8071, n8070, n8069, n8068, n8067, n8066, n8065, n8064, n8063};
wire [12:0]I4_8_8;
assign I4_8_8 = {n8088, n8087, n8086, n8085, n8084, n8083, n8082, n8081, n8080, n8079, n8078, n8077, n8076};
wire [19:0]O_8_8;
assign {n8108, n8107, n8106, n8105, n8104, n8103, n8102, n8101, n8100, n8099, n8098, n8097, n8096, n8095, n8094, n8093, n8092, n8091, n8090, n8089} = O_8_8;

clb clb_8_8 ( .clk(clk_8_8), .reset(fpga_rst), .I4(I4_8_8), .I3(I3_8_8), .I2(I2_8_8), .I1(I1_8_8), .O(O_8_8), .config_in(config_chain[176523:174564]), .config_rst(config_rst) );

wire [0:0]clk_8_9;
assign clk_8_9 = {fpga_clk};
wire [12:0]I1_8_9;
assign I1_8_9 = {n8147, n8146, n8145, n8144, n8143, n8142, n8141, n8140, n8139, n8138, n8137, n8136, n8135};
wire [12:0]I2_8_9;
assign I2_8_9 = {n8160, n8159, n8158, n8157, n8156, n8155, n8154, n8153, n8152, n8151, n8150, n8149, n8148};
wire [12:0]I3_8_9;
assign I3_8_9 = {n8173, n8172, n8171, n8170, n8169, n8168, n8167, n8166, n8165, n8164, n8163, n8162, n8161};
wire [12:0]I4_8_9;
assign I4_8_9 = {n8186, n8185, n8184, n8183, n8182, n8181, n8180, n8179, n8178, n8177, n8176, n8175, n8174};
wire [19:0]O_8_9;
assign {n8206, n8205, n8204, n8203, n8202, n8201, n8200, n8199, n8198, n8197, n8196, n8195, n8194, n8193, n8192, n8191, n8190, n8189, n8188, n8187} = O_8_9;

clb clb_8_9 ( .clk(clk_8_9), .reset(fpga_rst), .I4(I4_8_9), .I3(I3_8_9), .I2(I2_8_9), .I1(I1_8_9), .O(O_8_9), .config_in(config_chain[178483:176524]), .config_rst(config_rst) );

wire [7:0]outpad_8_10;
assign outpad_8_10 = {n8253, n8250, n8247, n8244, n8241, n8238, n8235, n8232};
wire [7:0]inpad_8_10;
assign {n8254, n8251, n8248, n8245, n8242, n8239, n8236, n8233} = inpad_8_10;

io io_8_10 ( .outpad(outpad_8_10), .inpad(inpad_8_10), .io_ext(io_8_10_wire), .config_in(config_chain[178491:178484]), .config_rst(config_rst) );

wire [7:0]outpad_9_0;
assign outpad_9_0 = {n8301, n8298, n8295, n8292, n8289, n8286, n8283, n8280};
wire [7:0]inpad_9_0;
assign {n8302, n8299, n8296, n8293, n8290, n8287, n8284, n8281} = inpad_9_0;

io io_9_0 ( .outpad(outpad_9_0), .inpad(inpad_9_0), .io_ext(io_9_0_wire), .config_in(config_chain[178499:178492]), .config_rst(config_rst) );

wire [0:0]clk_9_1;
assign clk_9_1 = {fpga_clk};
wire [12:0]I1_9_1;
assign I1_9_1 = {n8341, n8340, n8339, n8338, n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329};
wire [12:0]I2_9_1;
assign I2_9_1 = {n8354, n8353, n8352, n8351, n8350, n8349, n8348, n8347, n8346, n8345, n8344, n8343, n8342};
wire [12:0]I3_9_1;
assign I3_9_1 = {n8367, n8366, n8365, n8364, n8363, n8362, n8361, n8360, n8359, n8358, n8357, n8356, n8355};
wire [12:0]I4_9_1;
assign I4_9_1 = {n8380, n8379, n8378, n8377, n8376, n8375, n8374, n8373, n8372, n8371, n8370, n8369, n8368};
wire [19:0]O_9_1;
assign {n8400, n8399, n8398, n8397, n8396, n8395, n8394, n8393, n8392, n8391, n8390, n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381} = O_9_1;

clb clb_9_1 ( .clk(clk_9_1), .reset(fpga_rst), .I4(I4_9_1), .I3(I3_9_1), .I2(I2_9_1), .I1(I1_9_1), .O(O_9_1), .config_in(config_chain[180459:178500]), .config_rst(config_rst) );

wire [0:0]clk_9_2;
assign clk_9_2 = {fpga_clk};
wire [12:0]I1_9_2;
assign I1_9_2 = {n8439, n8438, n8437, n8436, n8435, n8434, n8433, n8432, n8431, n8430, n8429, n8428, n8427};
wire [12:0]I2_9_2;
assign I2_9_2 = {n8452, n8451, n8450, n8449, n8448, n8447, n8446, n8445, n8444, n8443, n8442, n8441, n8440};
wire [12:0]I3_9_2;
assign I3_9_2 = {n8465, n8464, n8463, n8462, n8461, n8460, n8459, n8458, n8457, n8456, n8455, n8454, n8453};
wire [12:0]I4_9_2;
assign I4_9_2 = {n8478, n8477, n8476, n8475, n8474, n8473, n8472, n8471, n8470, n8469, n8468, n8467, n8466};
wire [19:0]O_9_2;
assign {n8498, n8497, n8496, n8495, n8494, n8493, n8492, n8491, n8490, n8489, n8488, n8487, n8486, n8485, n8484, n8483, n8482, n8481, n8480, n8479} = O_9_2;

clb clb_9_2 ( .clk(clk_9_2), .reset(fpga_rst), .I4(I4_9_2), .I3(I3_9_2), .I2(I2_9_2), .I1(I1_9_2), .O(O_9_2), .config_in(config_chain[182419:180460]), .config_rst(config_rst) );

wire [0:0]clk_9_3;
assign clk_9_3 = {fpga_clk};
wire [12:0]I1_9_3;
assign I1_9_3 = {n8537, n8536, n8535, n8534, n8533, n8532, n8531, n8530, n8529, n8528, n8527, n8526, n8525};
wire [12:0]I2_9_3;
assign I2_9_3 = {n8550, n8549, n8548, n8547, n8546, n8545, n8544, n8543, n8542, n8541, n8540, n8539, n8538};
wire [12:0]I3_9_3;
assign I3_9_3 = {n8563, n8562, n8561, n8560, n8559, n8558, n8557, n8556, n8555, n8554, n8553, n8552, n8551};
wire [12:0]I4_9_3;
assign I4_9_3 = {n8576, n8575, n8574, n8573, n8572, n8571, n8570, n8569, n8568, n8567, n8566, n8565, n8564};
wire [19:0]O_9_3;
assign {n8596, n8595, n8594, n8593, n8592, n8591, n8590, n8589, n8588, n8587, n8586, n8585, n8584, n8583, n8582, n8581, n8580, n8579, n8578, n8577} = O_9_3;

clb clb_9_3 ( .clk(clk_9_3), .reset(fpga_rst), .I4(I4_9_3), .I3(I3_9_3), .I2(I2_9_3), .I1(I1_9_3), .O(O_9_3), .config_in(config_chain[184379:182420]), .config_rst(config_rst) );

wire [0:0]clk_9_4;
assign clk_9_4 = {fpga_clk};
wire [12:0]I1_9_4;
assign I1_9_4 = {n8635, n8634, n8633, n8632, n8631, n8630, n8629, n8628, n8627, n8626, n8625, n8624, n8623};
wire [12:0]I2_9_4;
assign I2_9_4 = {n8648, n8647, n8646, n8645, n8644, n8643, n8642, n8641, n8640, n8639, n8638, n8637, n8636};
wire [12:0]I3_9_4;
assign I3_9_4 = {n8661, n8660, n8659, n8658, n8657, n8656, n8655, n8654, n8653, n8652, n8651, n8650, n8649};
wire [12:0]I4_9_4;
assign I4_9_4 = {n8674, n8673, n8672, n8671, n8670, n8669, n8668, n8667, n8666, n8665, n8664, n8663, n8662};
wire [19:0]O_9_4;
assign {n8694, n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684, n8683, n8682, n8681, n8680, n8679, n8678, n8677, n8676, n8675} = O_9_4;

clb clb_9_4 ( .clk(clk_9_4), .reset(fpga_rst), .I4(I4_9_4), .I3(I3_9_4), .I2(I2_9_4), .I1(I1_9_4), .O(O_9_4), .config_in(config_chain[186339:184380]), .config_rst(config_rst) );

wire [0:0]clk_9_5;
assign clk_9_5 = {fpga_clk};
wire [12:0]I1_9_5;
assign I1_9_5 = {n8733, n8732, n8731, n8730, n8729, n8728, n8727, n8726, n8725, n8724, n8723, n8722, n8721};
wire [12:0]I2_9_5;
assign I2_9_5 = {n8746, n8745, n8744, n8743, n8742, n8741, n8740, n8739, n8738, n8737, n8736, n8735, n8734};
wire [12:0]I3_9_5;
assign I3_9_5 = {n8759, n8758, n8757, n8756, n8755, n8754, n8753, n8752, n8751, n8750, n8749, n8748, n8747};
wire [12:0]I4_9_5;
assign I4_9_5 = {n8772, n8771, n8770, n8769, n8768, n8767, n8766, n8765, n8764, n8763, n8762, n8761, n8760};
wire [19:0]O_9_5;
assign {n8792, n8791, n8790, n8789, n8788, n8787, n8786, n8785, n8784, n8783, n8782, n8781, n8780, n8779, n8778, n8777, n8776, n8775, n8774, n8773} = O_9_5;

clb clb_9_5 ( .clk(clk_9_5), .reset(fpga_rst), .I4(I4_9_5), .I3(I3_9_5), .I2(I2_9_5), .I1(I1_9_5), .O(O_9_5), .config_in(config_chain[188299:186340]), .config_rst(config_rst) );

wire [0:0]clk_9_6;
assign clk_9_6 = {fpga_clk};
wire [12:0]I1_9_6;
assign I1_9_6 = {n8831, n8830, n8829, n8828, n8827, n8826, n8825, n8824, n8823, n8822, n8821, n8820, n8819};
wire [12:0]I2_9_6;
assign I2_9_6 = {n8844, n8843, n8842, n8841, n8840, n8839, n8838, n8837, n8836, n8835, n8834, n8833, n8832};
wire [12:0]I3_9_6;
assign I3_9_6 = {n8857, n8856, n8855, n8854, n8853, n8852, n8851, n8850, n8849, n8848, n8847, n8846, n8845};
wire [12:0]I4_9_6;
assign I4_9_6 = {n8870, n8869, n8868, n8867, n8866, n8865, n8864, n8863, n8862, n8861, n8860, n8859, n8858};
wire [19:0]O_9_6;
assign {n8890, n8889, n8888, n8887, n8886, n8885, n8884, n8883, n8882, n8881, n8880, n8879, n8878, n8877, n8876, n8875, n8874, n8873, n8872, n8871} = O_9_6;

clb clb_9_6 ( .clk(clk_9_6), .reset(fpga_rst), .I4(I4_9_6), .I3(I3_9_6), .I2(I2_9_6), .I1(I1_9_6), .O(O_9_6), .config_in(config_chain[190259:188300]), .config_rst(config_rst) );

wire [0:0]clk_9_7;
assign clk_9_7 = {fpga_clk};
wire [12:0]I1_9_7;
assign I1_9_7 = {n8929, n8928, n8927, n8926, n8925, n8924, n8923, n8922, n8921, n8920, n8919, n8918, n8917};
wire [12:0]I2_9_7;
assign I2_9_7 = {n8942, n8941, n8940, n8939, n8938, n8937, n8936, n8935, n8934, n8933, n8932, n8931, n8930};
wire [12:0]I3_9_7;
assign I3_9_7 = {n8955, n8954, n8953, n8952, n8951, n8950, n8949, n8948, n8947, n8946, n8945, n8944, n8943};
wire [12:0]I4_9_7;
assign I4_9_7 = {n8968, n8967, n8966, n8965, n8964, n8963, n8962, n8961, n8960, n8959, n8958, n8957, n8956};
wire [19:0]O_9_7;
assign {n8988, n8987, n8986, n8985, n8984, n8983, n8982, n8981, n8980, n8979, n8978, n8977, n8976, n8975, n8974, n8973, n8972, n8971, n8970, n8969} = O_9_7;

clb clb_9_7 ( .clk(clk_9_7), .reset(fpga_rst), .I4(I4_9_7), .I3(I3_9_7), .I2(I2_9_7), .I1(I1_9_7), .O(O_9_7), .config_in(config_chain[192219:190260]), .config_rst(config_rst) );

wire [0:0]clk_9_8;
assign clk_9_8 = {fpga_clk};
wire [12:0]I1_9_8;
assign I1_9_8 = {n9027, n9026, n9025, n9024, n9023, n9022, n9021, n9020, n9019, n9018, n9017, n9016, n9015};
wire [12:0]I2_9_8;
assign I2_9_8 = {n9040, n9039, n9038, n9037, n9036, n9035, n9034, n9033, n9032, n9031, n9030, n9029, n9028};
wire [12:0]I3_9_8;
assign I3_9_8 = {n9053, n9052, n9051, n9050, n9049, n9048, n9047, n9046, n9045, n9044, n9043, n9042, n9041};
wire [12:0]I4_9_8;
assign I4_9_8 = {n9066, n9065, n9064, n9063, n9062, n9061, n9060, n9059, n9058, n9057, n9056, n9055, n9054};
wire [19:0]O_9_8;
assign {n9086, n9085, n9084, n9083, n9082, n9081, n9080, n9079, n9078, n9077, n9076, n9075, n9074, n9073, n9072, n9071, n9070, n9069, n9068, n9067} = O_9_8;

clb clb_9_8 ( .clk(clk_9_8), .reset(fpga_rst), .I4(I4_9_8), .I3(I3_9_8), .I2(I2_9_8), .I1(I1_9_8), .O(O_9_8), .config_in(config_chain[194179:192220]), .config_rst(config_rst) );

wire [0:0]clk_9_9;
assign clk_9_9 = {fpga_clk};
wire [12:0]I1_9_9;
assign I1_9_9 = {n9125, n9124, n9123, n9122, n9121, n9120, n9119, n9118, n9117, n9116, n9115, n9114, n9113};
wire [12:0]I2_9_9;
assign I2_9_9 = {n9138, n9137, n9136, n9135, n9134, n9133, n9132, n9131, n9130, n9129, n9128, n9127, n9126};
wire [12:0]I3_9_9;
assign I3_9_9 = {n9151, n9150, n9149, n9148, n9147, n9146, n9145, n9144, n9143, n9142, n9141, n9140, n9139};
wire [12:0]I4_9_9;
assign I4_9_9 = {n9164, n9163, n9162, n9161, n9160, n9159, n9158, n9157, n9156, n9155, n9154, n9153, n9152};
wire [19:0]O_9_9;
assign {n9184, n9183, n9182, n9181, n9180, n9179, n9178, n9177, n9176, n9175, n9174, n9173, n9172, n9171, n9170, n9169, n9168, n9167, n9166, n9165} = O_9_9;

clb clb_9_9 ( .clk(clk_9_9), .reset(fpga_rst), .I4(I4_9_9), .I3(I3_9_9), .I2(I2_9_9), .I1(I1_9_9), .O(O_9_9), .config_in(config_chain[196139:194180]), .config_rst(config_rst) );

wire [7:0]outpad_9_10;
assign outpad_9_10 = {n9231, n9228, n9225, n9222, n9219, n9216, n9213, n9210};
wire [7:0]inpad_9_10;
assign {n9232, n9229, n9226, n9223, n9220, n9217, n9214, n9211} = inpad_9_10;

io io_9_10 ( .outpad(outpad_9_10), .inpad(inpad_9_10), .io_ext(io_9_10_wire), .config_in(config_chain[196147:196140]), .config_rst(config_rst) );

wire [7:0]outpad_10_1;
assign outpad_10_1 = {n9279, n9276, n9273, n9270, n9267, n9264, n9261, n9258};
wire [7:0]inpad_10_1;
assign {n9280, n9277, n9274, n9271, n9268, n9265, n9262, n9259} = inpad_10_1;

io io_10_1 ( .outpad(outpad_10_1), .inpad(inpad_10_1), .io_ext(io_10_1_wire), .config_in(config_chain[196155:196148]), .config_rst(config_rst) );

wire [7:0]outpad_10_2;
assign outpad_10_2 = {n9327, n9324, n9321, n9318, n9315, n9312, n9309, n9306};
wire [7:0]inpad_10_2;
assign {n9328, n9325, n9322, n9319, n9316, n9313, n9310, n9307} = inpad_10_2;

io io_10_2 ( .outpad(outpad_10_2), .inpad(inpad_10_2), .io_ext(io_10_2_wire), .config_in(config_chain[196163:196156]), .config_rst(config_rst) );

wire [7:0]outpad_10_3;
assign outpad_10_3 = {n9375, n9372, n9369, n9366, n9363, n9360, n9357, n9354};
wire [7:0]inpad_10_3;
assign {n9376, n9373, n9370, n9367, n9364, n9361, n9358, n9355} = inpad_10_3;

io io_10_3 ( .outpad(outpad_10_3), .inpad(inpad_10_3), .io_ext(io_10_3_wire), .config_in(config_chain[196171:196164]), .config_rst(config_rst) );

wire [7:0]outpad_10_4;
assign outpad_10_4 = {n9423, n9420, n9417, n9414, n9411, n9408, n9405, n9402};
wire [7:0]inpad_10_4;
assign {n9424, n9421, n9418, n9415, n9412, n9409, n9406, n9403} = inpad_10_4;

io io_10_4 ( .outpad(outpad_10_4), .inpad(inpad_10_4), .io_ext(io_10_4_wire), .config_in(config_chain[196179:196172]), .config_rst(config_rst) );

wire [7:0]outpad_10_5;
assign outpad_10_5 = {n9471, n9468, n9465, n9462, n9459, n9456, n9453, n9450};
wire [7:0]inpad_10_5;
assign {n9472, n9469, n9466, n9463, n9460, n9457, n9454, n9451} = inpad_10_5;

io io_10_5 ( .outpad(outpad_10_5), .inpad(inpad_10_5), .io_ext(io_10_5_wire), .config_in(config_chain[196187:196180]), .config_rst(config_rst) );

wire [7:0]outpad_10_6;
assign outpad_10_6 = {n9519, n9516, n9513, n9510, n9507, n9504, n9501, n9498};
wire [7:0]inpad_10_6;
assign {n9520, n9517, n9514, n9511, n9508, n9505, n9502, n9499} = inpad_10_6;

io io_10_6 ( .outpad(outpad_10_6), .inpad(inpad_10_6), .io_ext(io_10_6_wire), .config_in(config_chain[196195:196188]), .config_rst(config_rst) );

wire [7:0]outpad_10_7;
assign outpad_10_7 = {n9567, n9564, n9561, n9558, n9555, n9552, n9549, n9546};
wire [7:0]inpad_10_7;
assign {n9568, n9565, n9562, n9559, n9556, n9553, n9550, n9547} = inpad_10_7;

io io_10_7 ( .outpad(outpad_10_7), .inpad(inpad_10_7), .io_ext(io_10_7_wire), .config_in(config_chain[196203:196196]), .config_rst(config_rst) );

wire [7:0]outpad_10_8;
assign outpad_10_8 = {n9615, n9612, n9609, n9606, n9603, n9600, n9597, n9594};
wire [7:0]inpad_10_8;
assign {n9616, n9613, n9610, n9607, n9604, n9601, n9598, n9595} = inpad_10_8;

io io_10_8 ( .outpad(outpad_10_8), .inpad(inpad_10_8), .io_ext(io_10_8_wire), .config_in(config_chain[196211:196204]), .config_rst(config_rst) );

wire [7:0]outpad_10_9;
assign outpad_10_9 = {n9663, n9660, n9657, n9654, n9651, n9648, n9645, n9642};
wire [7:0]inpad_10_9;
assign {n9664, n9661, n9658, n9655, n9652, n9649, n9646, n9643} = inpad_10_9;

io io_10_9 ( .outpad(outpad_10_9), .inpad(inpad_10_9), .io_ext(io_10_9_wire), .config_in(config_chain[196219:196212]), .config_rst(config_rst) );

config_helper config_helper( .config_in(config_in), .config_out(config_chain[`CONFIG_SIZE-1:0]), .clk(config_clk) );

endmodule

