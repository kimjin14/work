module dsip (
	pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_, pkey_243_, pcount_2_, 
	pkey_4_, pkey_132_, pkey_158_, pkey_169_, pkey_242_, pcount_1_, pkey_146_, pkey_168_, pkey_245_, pcount_0_, 
	pkey_6_, pkey_130_, pkey_145_, pkey_244_, pkey_9_, pkey_16_, pkey_27_, pkey_38_, pkey_49_, pkey_122_, 
	pkey_148_, pkey_153_, pkey_166_, pkey_221_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_48_, pkey_110_, 
	pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_, pkey_246_, pkey_253_, pkey_18_, pkey_29_, pkey_36_, 
	pkey_120_, pkey_155_, pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_, pkey_37_, pkey_46_, 
	pkey_112_, pkey_149_, pkey_156_, pkey_163_, pkey_211_, pkey_248_, pkey_56_, pkey_67_, pkey_78_, pkey_89_, 
	pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_, pkey_238_, pkey_57_, pkey_66_, pkey_88_, 
	pkey_114_, pkey_125_, pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_58_, pkey_69_, pkey_76_, pkey_115_, 
	pkey_124_, pkey_137_, pkey_160_, pkey_214_, pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_, 
	pkey_123_, pkey_138_, pkey_152_, pkey_222_, pkey_237_, pkey_251_, pkey_1_, pkey_96_, pkey_117_, pkey_140_, 
	pkey_216_, pkey_229_, pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_, pkey_217_, pkey_228_, 
	pkey_235_, pkey_3_, pkey_98_, pkey_128_, pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_, 
	pkey_2_, pkey_99_, pkey_134_, pkey_141_, pkey_219_, pkey_226_, pkey_233_, pkey_240_, pkey_70_, pkey_81_, 
	pkey_92_, pkey_180_, pkey_193_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, pclk, pkey_50_, 
	pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_, pstart_0_, pkey_51_, pkey_60_, pkey_109_, pkey_181_, 
	pkey_196_, pkey_208_, pkey_52_, pkey_74_, pkey_85_, pkey_104_, pkey_171_, pkey_197_, pkey_203_, pencrypt_0_, 
	pkey_53_, pkey_62_, pkey_75_, pkey_84_, pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_, pkey_72_, 
	pkey_83_, pkey_90_, pkey_106_, pkey_205_, pkey_64_, pkey_73_, pkey_82_, pkey_91_, pkey_105_, pkey_170_, 
	pkey_204_, pkey_12_, pkey_34_, pkey_45_, pkey_100_, pkey_188_, pkey_13_, pkey_22_, pkey_35_, pkey_44_, 
	pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_, pkey_102_, pkey_173_, pkey_201_, pkey_24_, 
	pkey_33_, pkey_42_, pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_, pkey_179_, pkey_184_, 
	pkey_40_, pkey_190_, pkey_10_, pkey_21_, pkey_177_, pkey_186_, pkey_11_, pkey_20_, pkey_178_, pkey_185_, 
	pkey_192_, pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_, pksi_115_, pksi_128_, pdata_ready_0_, 
	pksi_51_, pksi_60_, pksi_73_, pksi_82_, pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_, pksi_63_, 
	pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_, pksi_62_, pksi_71_, pksi_80_, pksi_97_, 
	pksi_114_, pksi_129_, pksi_54_, pksi_65_, pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_, pksi_191_, 
	pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_, pksi_56_, pksi_67_, pksi_74_, pksi_85_, 
	pksi_92_, pksi_117_, pksi_126_, pksi_57_, pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_, 
	pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_, pksi_24_, pksi_37_, pksi_46_, 
	pksi_109_, pnew_count_3_, pksi_16_, pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_, 
	pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_, pksi_43_, pksi_106_, pksi_111_, 
	pnew_count_0_, pksi_11_, pksi_20_, pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_, 
	pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_, pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, 
	pksi_3_, pksi_151_, pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_, pksi_189_, pksi_1_, 
	pksi_166_, pksi_179_, pksi_188_, pksi_0_, pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_, 
	pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_, pksi_141_, pksi_167_, pksi_174_, pksi_185_, 
	pksi_38_, pksi_49_, pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_, pksi_132_, pksi_169_, 
	pksi_176_, pksi_183_, pksi_58_, pksi_69_, pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_, 
	pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_, pksi_89_, pksi_135_, pksi_144_, pksi_157_, 
	pksi_171_, pksi_180_, pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_, pksi_172_, pksi_7_, 
	pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_, pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, 
	pksi_139_, pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_, pksi_161_);

input pcount_3_;
input pkey_5_;
input pkey_131_;
input pkey_144_;
input pkey_157_;
input pkey_230_;
input pkey_243_;
input pcount_2_;
input pkey_4_;
input pkey_132_;
input pkey_158_;
input pkey_169_;
input pkey_242_;
input pcount_1_;
input pkey_146_;
input pkey_168_;
input pkey_245_;
input pcount_0_;
input pkey_6_;
input pkey_130_;
input pkey_145_;
input pkey_244_;
input pkey_9_;
input pkey_16_;
input pkey_27_;
input pkey_38_;
input pkey_49_;
input pkey_122_;
input pkey_148_;
input pkey_153_;
input pkey_166_;
input pkey_221_;
input pkey_252_;
input pkey_8_;
input pkey_17_;
input pkey_26_;
input pkey_48_;
input pkey_110_;
input pkey_121_;
input pkey_147_;
input pkey_154_;
input pkey_165_;
input pkey_220_;
input pkey_246_;
input pkey_253_;
input pkey_18_;
input pkey_29_;
input pkey_36_;
input pkey_120_;
input pkey_155_;
input pkey_164_;
input pkey_210_;
input pkey_249_;
input pkey_254_;
input pkey_19_;
input pkey_28_;
input pkey_37_;
input pkey_46_;
input pkey_112_;
input pkey_149_;
input pkey_156_;
input pkey_163_;
input pkey_211_;
input pkey_248_;
input pkey_56_;
input pkey_67_;
input pkey_78_;
input pkey_89_;
input pkey_113_;
input pkey_126_;
input pkey_139_;
input pkey_162_;
input pkey_212_;
input pkey_225_;
input pkey_238_;
input pkey_57_;
input pkey_66_;
input pkey_88_;
input pkey_114_;
input pkey_125_;
input pkey_150_;
input pkey_161_;
input pkey_213_;
input pkey_224_;
input pkey_58_;
input pkey_69_;
input pkey_76_;
input pkey_115_;
input pkey_124_;
input pkey_137_;
input pkey_160_;
input pkey_214_;
input pkey_250_;
input pkey_59_;
input pkey_68_;
input pkey_77_;
input pkey_86_;
input pkey_116_;
input pkey_123_;
input pkey_138_;
input pkey_152_;
input pkey_222_;
input pkey_237_;
input pkey_251_;
input pkey_1_;
input pkey_96_;
input pkey_117_;
input pkey_140_;
input pkey_216_;
input pkey_229_;
input pkey_234_;
input pkey_0_;
input pkey_97_;
input pkey_118_;
input pkey_129_;
input pkey_136_;
input pkey_217_;
input pkey_228_;
input pkey_235_;
input pkey_3_;
input pkey_98_;
input pkey_128_;
input pkey_133_;
input pkey_142_;
input pkey_218_;
input pkey_227_;
input pkey_232_;
input pkey_241_;
input pkey_2_;
input pkey_99_;
input pkey_134_;
input pkey_141_;
input pkey_219_;
input pkey_226_;
input pkey_233_;
input pkey_240_;
input pkey_70_;
input pkey_81_;
input pkey_92_;
input pkey_180_;
input pkey_193_;
input pkey_80_;
input pkey_93_;
input pkey_107_;
input pkey_194_;
input pkey_206_;
input pclk;
input pkey_50_;
input pkey_61_;
input pkey_94_;
input pkey_182_;
input pkey_195_;
input pkey_209_;
input pstart_0_;
input pkey_51_;
input pkey_60_;
input pkey_109_;
input pkey_181_;
input pkey_196_;
input pkey_208_;
input pkey_52_;
input pkey_74_;
input pkey_85_;
input pkey_104_;
input pkey_171_;
input pkey_197_;
input pkey_203_;
input pencrypt_0_;
input pkey_53_;
input pkey_62_;
input pkey_75_;
input pkey_84_;
input pkey_172_;
input pkey_198_;
input pkey_202_;
input pkey_54_;
input pkey_65_;
input pkey_72_;
input pkey_83_;
input pkey_90_;
input pkey_106_;
input pkey_205_;
input pkey_64_;
input pkey_73_;
input pkey_82_;
input pkey_91_;
input pkey_105_;
input pkey_170_;
input pkey_204_;
input pkey_12_;
input pkey_34_;
input pkey_45_;
input pkey_100_;
input pkey_188_;
input pkey_13_;
input pkey_22_;
input pkey_35_;
input pkey_44_;
input pkey_176_;
input pkey_187_;
input pkey_14_;
input pkey_25_;
input pkey_32_;
input pkey_43_;
input pkey_102_;
input pkey_173_;
input pkey_201_;
input pkey_24_;
input pkey_33_;
input pkey_42_;
input pkey_101_;
input pkey_174_;
input pkey_189_;
input pkey_200_;
input pkey_30_;
input pkey_41_;
input pkey_179_;
input pkey_184_;
input pkey_40_;
input pkey_190_;
input pkey_10_;
input pkey_21_;
input pkey_177_;
input pkey_186_;
input pkey_11_;
input pkey_20_;
input pkey_178_;
input pkey_185_;
input pkey_192_;
output pksi_50_;
output pksi_61_;
output pksi_72_;
output pksi_83_;
output pksi_94_;
output pksi_102_;
output pksi_115_;
output pksi_128_;
output pdata_ready_0_;
output pksi_51_;
output pksi_60_;
output pksi_73_;
output pksi_82_;
output pksi_95_;
output pksi_101_;
output pksi_116_;
output pksi_127_;
output pksi_52_;
output pksi_63_;
output pksi_70_;
output pksi_81_;
output pksi_96_;
output pksi_100_;
output pksi_113_;
output pksi_53_;
output pksi_62_;
output pksi_71_;
output pksi_80_;
output pksi_97_;
output pksi_114_;
output pksi_129_;
output pksi_54_;
output pksi_65_;
output pksi_76_;
output pksi_87_;
output pksi_90_;
output pksi_119_;
output pksi_124_;
output pksi_191_;
output pksi_55_;
output pksi_64_;
output pksi_77_;
output pksi_86_;
output pksi_91_;
output pksi_123_;
output pksi_56_;
output pksi_67_;
output pksi_74_;
output pksi_85_;
output pksi_92_;
output pksi_117_;
output pksi_126_;
output pksi_57_;
output pksi_66_;
output pksi_75_;
output pksi_84_;
output pksi_93_;
output pksi_118_;
output pksi_125_;
output pksi_190_;
output pksi_14_;
output pksi_25_;
output pksi_36_;
output pksi_47_;
output pksi_120_;
output pksi_15_;
output pksi_24_;
output pksi_37_;
output pksi_46_;
output pksi_109_;
output pnew_count_3_;
output pksi_16_;
output pksi_27_;
output pksi_34_;
output pksi_45_;
output pksi_108_;
output pksi_122_;
output pksi_17_;
output pksi_26_;
output pksi_35_;
output pksi_44_;
output pksi_107_;
output pksi_121_;
output pksi_10_;
output pksi_21_;
output pksi_32_;
output pksi_43_;
output pksi_106_;
output pksi_111_;
output pnew_count_0_;
output pksi_11_;
output pksi_20_;
output pksi_33_;
output pksi_42_;
output pksi_105_;
output pksi_112_;
output pksi_12_;
output pksi_23_;
output pksi_30_;
output pksi_41_;
output pksi_104_;
output pnew_count_2_;
output pksi_13_;
output pksi_22_;
output pksi_31_;
output pksi_40_;
output pksi_103_;
output pksi_110_;
output pnew_count_1_;
output pksi_3_;
output pksi_151_;
output pksi_164_;
output pksi_177_;
output pksi_2_;
output pksi_152_;
output pksi_163_;
output pksi_178_;
output pksi_189_;
output pksi_1_;
output pksi_166_;
output pksi_179_;
output pksi_188_;
output pksi_0_;
output pksi_150_;
output pksi_165_;
output pksi_187_;
output pksi_18_;
output pksi_29_;
output pksi_142_;
output pksi_168_;
output pksi_173_;
output pksi_186_;
output pksi_19_;
output pksi_28_;
output pksi_130_;
output pksi_141_;
output pksi_167_;
output pksi_174_;
output pksi_185_;
output pksi_38_;
output pksi_49_;
output pksi_131_;
output pksi_140_;
output pksi_175_;
output pksi_184_;
output pksi_39_;
output pksi_48_;
output pksi_132_;
output pksi_169_;
output pksi_176_;
output pksi_183_;
output pksi_58_;
output pksi_69_;
output pksi_133_;
output pksi_146_;
output pksi_159_;
output pksi_182_;
output pksi_59_;
output pksi_68_;
output pksi_134_;
output pksi_145_;
output pksi_170_;
output pksi_181_;
output pksi_9_;
output pksi_78_;
output pksi_89_;
output pksi_135_;
output pksi_144_;
output pksi_157_;
output pksi_171_;
output pksi_180_;
output pksi_8_;
output pksi_79_;
output pksi_88_;
output pksi_136_;
output pksi_143_;
output pksi_158_;
output pksi_172_;
output pksi_7_;
output pksi_98_;
output pksi_137_;
output pksi_155_;
output pksi_160_;
output pksi_6_;
output pksi_99_;
output pksi_138_;
output pksi_149_;
output pksi_156_;
output pksi_5_;
output pksi_139_;
output pksi_148_;
output pksi_153_;
output pksi_162_;
output pksi_4_;
output pksi_147_;
output pksi_154_;
output pksi_161_;
wire n_n2385;
wire n_n2397;
wire n_n2409;
wire n_n2424;
wire n_n2436;
wire n_n2449;
wire n_n2500;
wire n_n2512;
wire n_n2386;
wire n_n2395;
wire n_n2411;
wire n_n2423;
wire n_n2437;
wire n_n2447;
wire n_n2501;
wire n_n2511;
wire n_n2387;
wire n_n2399;
wire n_n2406;
wire n_n2422;
wire n_n2459;
wire n_n2471;
wire n_n2502;
wire n_n2515;
wire n_n2523;
wire n_n2388;
wire n_n2398;
wire n_n2407;
wire n_n2421;
wire n_n2460;
wire n_n2470;
wire n_n2503;
wire n_n2514;
wire n_n2275;
wire n_n2380;
wire n_n2392;
wire n_n2404;
wire n_n2419;
wire n_n2483;
wire n_n2496;
wire n_n2508;
wire n_n2521;
wire n_n2381;
wire n_n2391;
wire n_n2405;
wire n_n2418;
wire n_n2484;
wire n_n2494;
wire n_n2497;
wire n_n2522;
wire n_n2382;
wire n_n2394;
wire n_n2402;
wire n_n2417;
wire n_n2498;
wire n_n2510;
wire n_n2383;
wire n_n2393;
wire n_n2403;
wire n_n2415;
wire n_n2499;
wire n_n2509;
wire n_n2520;
wire n_n2270;
wire n_n2427;
wire n_n2439;
wire n_n2453;
wire n_n2465;
wire n_n2478;
wire n_n2491;
wire n_n2271;
wire n_n2428;
wire n_n2438;
wire n_n2454;
wire n_n2464;
wire n_n2479;
wire n_n2490;
wire n_n2273;
wire n_n2429;
wire n_n2442;
wire n_n2450;
wire n_n2463;
wire n_n2480;
wire n_n2493;
wire n_n2274;
wire n_n2431;
wire n_n2441;
wire n_n2451;
wire n_n2461;
wire n_n2482;
wire n_n2492;
wire n_n2265;
wire n_n2389;
wire n_n2401;
wire n_n2432;
wire n_n2444;
wire n_n2457;
wire n_n2469;
wire n_n2472;
wire n_n2487;
wire n_n2504;
wire n_n2518;
wire n_n2266;
wire n_n2390;
wire n_n2400;
wire n_n2433;
wire n_n2443;
wire n_n2458;
wire n_n2468;
wire n_n2473;
wire n_n2486;
wire n_n2505;
wire n_n2516;
wire n_n2267;
wire n_n2413;
wire n_n2426;
wire n_n2434;
wire n_n2446;
wire n_n2455;
wire n_n2467;
wire n_n2475;
wire n_n2489;
wire n_n2506;
wire n_n2269;
wire n_n2414;
wire n_n2425;
wire n_n2435;
wire n_n2445;
wire n_n2456;
wire n_n2466;
wire n_n2477;
wire n_n2488;
wire n_n2519;
wire n_n2323;
wire n_n2335;
wire n_n2348;
wire n_n2360;
wire n_n2373;
wire n_n2324;
wire n_n2334;
wire n_n2349;
wire n_n2359;
wire n_n2375;
wire n_n2325;
wire n_n2338;
wire n_n2346;
wire n_n2358;
wire n_n2376;
wire n_n2264;
wire n_n2326;
wire n_n2336;
wire n_n2347;
wire n_n2357;
wire n_n2377;
wire n_n2276;
wire n_n2290;
wire n_n2302;
wire n_n2315;
wire n_n2378;
wire n_n2278;
wire n_n2289;
wire n_n2303;
wire n_n2314;
wire n_n2379;
wire n_n2279;
wire n_n2292;
wire n_n2299;
wire n_n2313;
wire n_n2281;
wire n_n2291;
wire n_n2300;
wire n_n2312;
wire n_n2282;
wire n_n2294;
wire n_n2307;
wire n_n2319;
wire n_n2331;
wire n_n2345;
wire n_n2283;
wire n_n2293;
wire n_n2308;
wire n_n2318;
wire n_n2332;
wire n_n2344;
wire n_n2284;
wire n_n2296;
wire n_n2304;
wire n_n2317;
wire n_n2355;
wire n_n2367;
wire n_n2285;
wire n_n2295;
wire n_n2306;
wire n_n2316;
wire n_n2356;
wire n_n2366;
wire n_n2286;
wire n_n2298;
wire n_n2327;
wire n_n2340;
wire n_n2353;
wire n_n2364;
wire n_n2368;
wire n_n2287;
wire n_n2297;
wire n_n2328;
wire n_n2339;
wire n_n2354;
wire n_n2363;
wire n_n2370;
wire n_n2309;
wire n_n2322;
wire n_n2329;
wire n_n2343;
wire n_n2350;
wire n_n2362;
wire n_n2371;
wire n_n2311;
wire n_n2321;
wire n_n2330;
wire n_n2341;
wire n_n2351;
wire n_n2361;
wire n_n2372;
wire n_n200;
wire n_n204;
wire wire653;
wire n_n2530;
wire wire647;
wire wire655;
wire wire664;
wire wire669;
wire wire670;
wire wire673;
wire wire682;
wire wire684;
wire wire687;
wire wire689;
wire wire692;
wire wire693;
wire wire695;
wire wire698;
wire wire699;
wire wire701;
wire wire704;
wire wire705;
wire wire706;
wire wire710;
wire wire711;
wire wire714;
wire wire716;
wire wire717;
wire wire719;
wire wire722;
wire wire723;
wire wire725;
wire wire728;
wire wire729;
wire wire730;
wire wire734;
wire wire735;
wire wire736;
wire wire738;
wire wire741;
wire wire744;
wire wire746;
wire wire747;
wire wire749;
wire wire752;
wire wire753;
wire wire756;
wire wire758;
wire wire759;
wire wire761;
wire wire764;
wire wire765;
wire wire768;
wire wire770;
wire wire771;
wire wire772;
wire wire774;
wire wire777;
wire wire780;
wire wire782;
wire wire783;
wire wire784;
wire wire788;
wire wire789;
wire wire791;
wire wire794;
wire wire795;
wire wire797;
wire wire800;
wire wire801;
wire wire803;
wire wire806;
wire wire807;
wire wire809;
wire wire812;
wire wire813;
wire wire815;
wire wire818;
wire wire819;
wire wire822;
wire wire824;
wire wire825;
wire wire826;
wire wire828;
wire wire831;
wire wire833;
wire wire836;
wire wire837;
wire wire839;
wire wire842;
wire wire843;
wire wire845;
wire wire848;
wire wire849;
wire wire850;
wire wire854;
wire wire855;
wire wire857;
wire wire860;
wire wire861;
wire wire863;
wire wire866;
wire wire867;
wire wire869;
wire wire872;
wire wire873;
wire wire875;
wire wire878;
wire wire879;
wire wire881;
wire wire884;
wire wire885;
wire wire886;
wire wire889;
wire wire891;
wire wire893;
wire wire896;
wire wire897;
wire wire898;
wire wire902;
wire wire903;
wire wire905;
wire wire908;
wire wire909;
wire wire911;
wire wire914;
wire wire915;
wire wire917;
wire wire920;
wire wire921;
wire wire924;
wire wire926;
wire wire927;
wire wire929;
wire wire932;
wire wire933;
wire wire934;
wire wire936;
wire wire939;
wire wire941;
wire wire944;
wire wire945;
wire wire947;
wire wire950;
wire wire951;
wire wire953;
wire wire956;
wire wire957;
wire wire959;
wire wire962;
wire wire963;
wire wire964;
wire wire966;
wire wire969;
wire wire971;
wire wire974;
wire wire975;
wire wire977;
wire wire980;
wire wire981;
wire wire983;
wire wire986;
wire wire987;
wire wire989;
wire wire992;
wire wire993;
wire wire995;
wire wire998;
wire wire999;
wire wire1001;
wire wire1004;
wire wire1005;
wire wire1007;
wire wire1010;
wire wire1011;
wire wire1013;
wire wire1016;
wire wire1017;
wire wire1019;
wire wire1022;
wire wire1023;
wire wire1025;
wire wire1028;
wire wire1029;
wire wire1031;
wire wire1034;
wire wire1035;
wire wire1038;
wire wire1040;
wire wire1041;
wire wire1043;
wire wire1046;
wire wire1047;
wire wire1049;
wire wire1052;
wire wire1053;
wire wire1055;
wire wire1058;
wire wire1059;
wire wire1061;
wire wire1064;
wire wire1065;
wire wire1068;
wire wire1070;
wire wire1071;
wire wire1073;
wire wire1076;
wire wire1077;
wire wire1079;
wire wire1082;
wire wire1083;
wire wire1085;
wire wire1088;
wire wire1089;
wire wire1091;
wire wire1094;
wire wire1095;
wire wire1097;
wire wire1100;
wire wire1101;
wire wire1103;
wire wire1106;
wire wire1107;
wire wire1109;
wire wire1112;
wire wire1113;
wire wire1115;
wire wire1118;
wire wire1119;
wire wire1121;
wire wire1124;
wire wire1125;
wire wire1127;
wire wire1130;
wire wire1131;
wire wire1133;
wire wire1136;
wire wire1137;
wire wire1140;
wire wire1142;
wire wire1143;
wire wire1145;
wire wire1148;
wire wire1149;
wire wire1151;
wire wire1154;
wire wire1155;
wire wire1158;
wire wire1160;
wire wire1161;
wire wire1163;
wire wire1166;
wire wire1167;
wire wire1170;
wire wire1172;
wire wire1173;
wire wire1175;
wire wire1178;
wire wire1179;
wire wire1180;
wire wire1184;
wire wire1185;
wire wire1187;
wire wire1190;
wire wire1191;
wire wire1193;
wire wire1196;
wire wire1197;
wire wire1199;
wire wire1202;
wire wire1203;
wire wire1205;
wire wire1208;
wire wire1209;
wire wire1211;
wire wire1214;
wire wire1215;
wire wire1217;
wire wire1219;
wire wire1221;
wire wire1223;
wire wire1226;
wire wire1227;
wire wire1229;
wire wire1232;
wire wire1233;
wire wire1235;
wire wire1238;
wire wire1239;
wire wire1242;
wire wire1243;
wire wire1245;
wire wire1247;
wire wire1250;
wire wire1251;
wire wire1253;
wire wire1256;
wire wire1257;
wire wire1259;
wire wire1262;
wire wire1263;
wire wire1265;
wire wire1268;
wire wire1269;
wire wire1271;
wire wire1274;
wire wire1275;
wire wire1277;
wire wire1280;
wire wire1281;
wire wire1284;
wire wire1286;
wire wire1287;
wire wire1289;
wire wire1292;
wire wire1293;
wire wire1295;
wire wire1298;
wire wire1299;
wire wire1302;
wire wire1304;
wire wire1305;
wire wire1307;
wire wire1310;
wire wire1311;
wire wire1313;
wire wire1316;
wire wire1317;
wire wire1319;
wire wire1322;
wire wire1323;
wire wire1325;
wire wire1328;
wire wire1329;
wire wire1331;
wire wire1334;
wire wire1335;
wire wire1337;
wire wire1340;
wire wire1341;
wire wire1343;
wire wire1346;
wire wire1347;
wire wire1349;
wire wire1352;
wire wire1353;
wire wire1355;
wire wire1357;
wire wire1359;
wire wire1361;
wire wire1364;
wire wire1365;
wire wire1367;
wire wire1368;
wire wire1371;
wire wire1373;
wire wire1376;
wire wire1377;
wire wire1379;
wire wire1382;
wire wire1383;
wire wire1385;
wire wire1388;
wire wire1389;
wire wire1391;
wire wire1394;
wire wire1395;
wire wire1397;
wire wire1400;
wire wire1401;
wire wire1403;
wire wire1406;
wire wire1407;
wire wire1408;
wire wire1410;
wire wire1413;
wire wire1415;
wire wire1418;
wire wire1419;
wire wire1421;
wire wire1424;
wire wire1425;
wire wire1427;
wire wire1430;
wire wire1431;
wire wire1432;
wire wire1434;
wire wire1437;
wire wire1439;
wire wire1442;
wire wire1443;
wire wire1445;
wire wire1448;
wire wire1449;
wire wire1451;
wire wire1454;
wire wire1455;
wire wire1457;
wire wire1460;
wire wire1461;
wire wire1463;
wire wire1466;
wire wire1467;
wire wire1469;
wire wire1472;
wire wire1473;
wire wire1474;
wire wire1478;
wire wire1479;
wire wire1481;
wire wire1484;
wire wire1485;
wire wire1487;
wire wire1490;
wire wire1491;
wire wire1493;
wire wire1496;
wire wire1497;
wire wire1499;
wire wire1502;
wire wire1503;
wire wire1505;
wire wire1508;
wire wire1509;
wire wire1511;
wire wire1514;
wire wire1515;
wire wire1516;
wire wire1520;
wire wire1521;
wire wire1523;
wire wire1526;
wire wire1527;
wire wire1529;
wire wire1532;
wire wire1533;
wire wire1536;
wire wire1538;
wire wire1539;
wire wire1541;
wire wire1542;
wire wire1545;
wire wire1547;
wire wire1550;
wire wire1551;
wire wire1553;
wire wire1556;
wire wire1557;
wire wire1559;
wire wire1562;
wire wire1563;
wire wire1565;
wire wire1568;
wire wire1569;
wire wire1571;
wire wire1572;
wire wire1575;
wire wire1578;
wire wire1580;
wire wire1581;
wire wire1584;
wire wire1586;
wire wire1587;
wire wire1589;
wire wire1592;
wire wire1593;
wire wire1595;
wire wire1596;
wire wire1599;
wire wire1601;
wire wire1604;
wire wire1605;
wire wire1607;
wire wire1610;
wire wire1611;
wire wire1613;
wire wire1616;
wire wire1617;
wire wire1619;
wire wire1622;
wire wire1623;
wire wire1626;
wire wire1628;
wire wire1629;
wire wire1631;
wire wire1634;
wire wire1635;
wire wire1637;
wire wire1640;
wire wire1641;
wire wire1644;
wire wire1646;
wire wire1647;
wire wire1649;
wire wire1652;
wire wire1653;
wire wire1655;
wire wire1658;
wire wire1659;
wire wire1661;
wire wire1664;
wire wire1665;
wire wire1667;
wire wire1670;
wire wire1671;
wire wire1673;
wire wire1676;
wire wire1677;
wire wire1679;
wire wire1682;
wire wire1683;
wire wire1685;
wire wire1688;
wire wire1689;
wire wire1691;
wire wire1694;
wire wire1695;
wire wire1697;
wire wire1700;
wire wire1701;
wire wire1703;
wire wire1706;
wire wire1707;
wire wire1709;
wire wire1712;
wire wire1713;
wire wire1715;
wire wire1718;
wire wire1719;
wire wire1721;
wire wire1724;
wire wire1725;
wire wire1727;
wire wire1730;
wire wire1731;
wire wire1733;
wire wire1736;
wire wire1737;
wire wire1739;
wire wire1742;
wire wire1743;
wire wire1745;
wire wire1748;
wire wire1749;
wire wire1751;
wire wire1754;
wire wire1755;
wire wire1757;
wire wire1760;
wire wire1761;
wire wire1763;
wire wire1766;
wire wire1767;
wire wire1769;
wire wire1772;
wire wire1773;
wire wire1775;
wire wire1778;
wire wire1779;
wire wire1781;
wire wire1784;
wire wire1785;
wire wire1787;
wire wire1790;
wire wire1791;
wire wire1793;
wire wire1796;
wire wire1797;
wire wire1799;
wire wire1802;
wire wire1803;
wire wire1805;
wire wire1808;
wire wire1809;
wire wire1811;
wire wire1814;
wire wire1815;
wire wire1817;
wire wire1820;
wire wire1821;
wire wire1822;
wire wire1824;
wire wire1827;
wire wire1829;
wire wire1832;
wire wire1833;
wire wire1835;
wire wire1838;
wire wire1839;
wire wire1841;
wire wire1844;
wire wire1845;
wire wire1847;
wire wire1848;
wire wire1851;
wire wire1853;
wire wire1856;
wire wire1857;
wire wire1859;
wire wire1862;
wire wire1863;
wire wire1865;
wire wire1868;
wire wire1869;
wire wire1871;
wire wire1874;
wire wire1875;
wire wire1877;
wire wire1880;
wire wire1881;
wire wire1883;
wire wire1885;
wire wire1887;
wire wire1889;
wire wire1892;
wire wire1893;
wire wire1894;
wire wire1898;
wire wire1899;
wire wire1901;
wire wire1904;
wire wire1905;
wire wire1907;
wire wire1910;
wire wire1911;
wire wire1913;
wire wire1916;
wire wire1917;
wire wire1919;
wire wire1922;
wire wire1923;
wire wire1925;
wire wire1928;
wire wire1929;
wire wire1931;
wire wire1934;
wire wire1935;
wire wire1937;
wire wire1940;
wire wire1941;
wire wire1943;
wire wire1946;
wire wire1947;
wire wire1949;
wire wire1952;
wire wire1953;
wire wire1955;
wire wire1958;
wire wire1959;
wire wire1961;
wire wire1964;
wire wire1965;
wire wire1967;
wire wire1970;
wire wire1971;
wire wire1973;
wire wire1976;
wire wire1977;
wire wire1979;
wire wire1982;
wire wire1983;
wire wire1985;
wire wire1988;
wire wire1989;
wire wire1991;
wire wire1994;
wire wire1995;
wire wire1997;
wire wire2000;
wire wire2001;
wire wire2003;
wire wire2006;
wire wire2007;
wire wire2009;
wire wire2012;
wire wire2013;
wire wire2015;
wire wire2018;
wire wire2019;
wire wire2021;
wire wire2024;
wire wire2025;
wire wire6182;
wire wire6183;
wire wire6186;
wire wire6187;
wire wire6190;
wire wire6191;
wire wire6194;
wire wire6195;
wire wire6198;
wire wire6199;
wire wire6202;
wire wire6203;
wire wire6206;
wire wire6207;
wire wire6210;
wire wire6211;
wire wire6214;
wire wire6215;
wire wire6218;
wire wire6219;
wire wire6222;
wire wire6223;
wire wire6226;
wire wire6227;
wire wire6230;
wire wire6231;
wire wire6234;
wire wire6235;
wire wire6238;
wire wire6239;
wire wire6242;
wire wire6243;
wire wire6246;
wire wire6247;
wire wire6250;
wire wire6251;
wire wire6254;
wire wire6255;
wire wire6258;
wire wire6259;
wire wire6262;
wire wire6263;
wire wire6266;
wire wire6267;
wire wire6270;
wire wire6271;
wire wire6274;
wire wire6275;
wire wire6278;
wire wire6279;
wire wire6282;
wire wire6283;
wire wire6286;
wire wire6287;
wire wire6290;
wire wire6291;
wire wire6294;
wire wire6295;
wire wire6298;
wire wire6299;
wire wire6302;
wire wire6303;
wire wire6306;
wire wire6307;
wire wire6310;
wire wire6311;
wire wire6314;
wire wire6315;
wire wire6318;
wire wire6319;
wire wire6322;
wire wire6323;
wire wire6326;
wire wire6327;
wire wire6330;
wire wire6331;
wire wire6334;
wire wire6335;
wire wire6338;
wire wire6339;
wire wire6342;
wire wire6343;
wire wire6346;
wire wire6347;
wire wire6350;
wire wire6351;
wire wire6354;
wire wire6355;
wire wire6358;
wire wire6359;
wire wire6362;
wire wire6363;
wire wire6366;
wire wire6367;
wire wire6370;
wire wire6371;
wire wire6374;
wire wire6375;
wire wire6378;
wire wire6379;
wire wire6382;
wire wire6383;
wire wire6386;
wire wire6387;
wire wire6390;
wire wire6391;
wire wire6394;
wire wire6395;
wire wire6398;
wire wire6399;
wire wire6402;
wire wire6403;
wire wire6406;
wire wire6407;
wire wire6410;
wire wire6411;
wire wire6414;
wire wire6415;
wire wire6418;
wire wire6419;
wire wire6422;
wire wire6423;
wire wire6426;
wire wire6427;
wire wire6430;
wire wire6431;
wire wire6434;
wire wire6435;
wire wire6438;
wire wire6439;
wire wire6442;
wire wire6443;
wire wire6446;
wire wire6447;
wire wire6450;
wire wire6451;
wire wire6454;
wire wire6455;
wire wire6458;
wire wire6459;
wire wire6462;
wire wire6463;
wire wire6466;
wire wire6467;
wire wire6470;
wire wire6471;
wire wire6474;
wire wire6475;
wire wire6478;
wire wire6479;
wire wire6482;
wire wire6483;
wire wire6486;
wire wire6487;
wire wire6490;
wire wire6491;
wire wire6494;
wire wire6495;
wire wire6498;
wire wire6499;
wire wire6502;
wire wire6503;
wire wire6506;
wire wire6507;
wire wire6510;
wire wire6511;
wire wire6514;
wire wire6515;
wire wire6518;
wire wire6519;
wire wire6522;
wire wire6523;
wire wire6526;
wire wire6527;
wire wire6530;
wire wire6531;
wire wire6534;
wire wire6535;
wire wire6538;
wire wire6539;
wire wire6542;
wire wire6543;
wire wire6546;
wire wire6547;
wire wire6550;
wire wire6551;
wire wire6554;
wire wire6555;
wire wire6558;
wire wire6559;
wire wire6562;
wire wire6563;
wire wire6566;
wire wire6567;
wire wire6570;
wire wire6571;
wire wire6574;
wire wire6575;
wire wire6578;
wire wire6579;
wire wire6582;
wire wire6583;
wire wire6586;
wire wire6587;
wire wire6590;
wire wire6591;
wire wire6594;
wire wire6595;
wire wire6598;
wire wire6599;
wire wire6602;
wire wire6603;
wire wire6606;
wire wire6607;
wire wire6610;
wire wire6611;
wire wire6614;
wire wire6615;
wire wire6618;
wire wire6619;
wire wire6622;
wire wire6623;
wire wire6626;
wire wire6627;
wire wire6630;
wire wire6631;
wire wire6634;
wire wire6635;
wire wire6638;
wire wire6639;
wire wire6642;
wire wire6643;
wire wire6646;
wire wire6647;
wire wire6650;
wire wire6651;
wire wire6654;
wire wire6655;
wire wire6658;
wire wire6659;
wire wire6662;
wire wire6663;
wire wire6666;
wire wire6667;
wire wire6670;
wire wire6671;
wire wire6674;
wire wire6675;
wire wire6678;
wire wire6679;
wire wire6682;
wire wire6683;
wire wire6686;
wire wire6687;
wire wire6690;
wire wire6691;
wire wire6694;
wire wire6695;
wire wire6698;
wire wire6699;
wire wire6702;
wire wire6703;
wire wire6706;
wire wire6707;
wire wire6710;
wire wire6711;
wire wire6714;
wire wire6715;
wire wire6718;
wire wire6719;
wire wire6722;
wire wire6723;
wire wire6726;
wire wire6727;
wire wire6730;
wire wire6731;
wire wire6734;
wire wire6735;
wire wire6738;
wire wire6739;
wire wire6742;
wire wire6743;
wire wire6746;
wire wire6747;
wire wire6750;
wire wire6751;
wire wire6754;
wire wire6755;
wire wire6758;
wire wire6759;
wire wire6762;
wire wire6763;
wire wire6766;
wire wire6767;
wire wire6770;
wire wire6771;
wire wire6774;
wire wire6775;
wire wire6778;
wire wire6779;
wire wire6782;
wire wire6783;
wire wire6786;
wire wire6787;
wire wire6790;
wire wire6791;
wire wire6794;
wire wire6795;
wire wire6798;
wire wire6799;
wire wire6802;
wire wire6803;
wire wire6806;
wire wire6807;
wire wire6810;
wire wire6811;
wire wire6814;
wire wire6815;
wire wire6818;
wire wire6819;
wire wire6822;
wire wire6823;
wire wire6826;
wire wire6827;
wire wire6830;
wire wire6831;
wire wire6834;
wire wire6835;
wire wire6838;
wire wire6839;
wire wire6842;
wire wire6843;
wire wire6846;
wire wire6847;
wire wire6850;
wire wire6851;
wire wire6854;
wire wire6855;
wire wire6858;
wire wire6859;
wire wire6862;
wire wire6863;
wire wire6866;
wire wire6867;
wire wire6870;
wire wire6871;
wire wire6874;
wire wire6875;
wire wire6878;
wire wire6879;
wire wire6882;
wire wire6883;
wire wire6886;
wire wire6887;
wire wire6890;
wire wire6891;
wire wire6894;
wire wire6895;
wire wire6898;
wire wire6899;
wire wire6902;
wire wire6903;
wire wire6906;
wire wire6907;
wire wire6910;
wire wire6911;
wire wire6914;
wire wire6915;
wire wire6918;
wire wire6919;
wire wire6922;
wire wire6923;
wire wire6926;
wire wire6927;
wire wire6930;
wire wire6931;
wire wire6934;
wire wire6935;
wire wire6938;
wire wire6939;
wire wire6942;
wire wire6943;
wire wire6946;
wire wire6947;
wire wire6950;
wire wire6951;
wire wire6954;
wire wire6955;
wire wire6958;
wire wire6959;
wire wire6962;
wire wire6963;
wire wire6966;
wire wire6967;
wire wire6970;
wire wire6971;
wire wire6974;
wire wire6975;
wire wire6978;
wire wire6979;
wire wire6982;
wire wire6983;
wire wire6986;
wire wire6987;
wire wire6990;
wire wire6991;
wire wire6994;
wire wire6995;
wire wire6998;
wire wire6999;
wire wire7002;
wire wire7003;
wire wire7006;
wire wire7007;
wire wire7010;
wire wire7011;
wire wire7014;
wire wire7015;
wire wire7018;
wire wire7019;
wire wire7022;
wire wire7023;
wire wire7026;
wire wire7027;
wire wire7030;
wire wire7031;
wire wire7034;
wire wire7035;
wire wire7038;
wire wire7039;
wire wire7042;
wire wire7043;
wire wire7046;
wire wire7047;
wire wire7050;
wire wire7051;
wire wire7054;
wire wire7055;
wire wire7058;
wire wire7059;
wire wire7062;
wire wire7063;
wire wire7066;
wire wire7067;
wire wire7070;
wire wire7071;
wire wire7074;
wire wire7075;
wire wire7079;
wire wire7081;
wire wire7084;
reg pksi_17_;

reg pksi_185_;

reg n_n2410;

reg pksi_170_;

reg pksi_155_;

reg pksi_147_;

reg pksi_109_;

reg n_n2513;

reg pksi_19_;

reg n_n2396;

reg n_n2412;

reg n_n121;

reg pksi_148_;

reg n_n2448;

reg pksi_107_;

reg pksi_110_;

reg pksi_9_;

reg pksi_176_;

reg pksi_180_;

reg pksi_178_;

reg pksi_135_;

reg pksi_129_;

reg pksi_100_;

reg pksi_117_;

reg pksi_118_;

reg pksi_5_;

reg pksi_169_;

reg n_n2408;

reg pksi_184_;

reg pksi_125_;

reg pksi_138_;

reg pksi_114_;

reg pksi_99_;

reg pksi_85_;

reg pksi_14_;

reg pksi_4_;

reg pksi_186_;

reg n_n2420;

reg pksi_141_;

reg pksi_113_;

reg pksi_115_;

reg pksi_98_;

reg pksi_2_;

reg pksi_23_;

reg pksi_177_;

reg pksi_189_;

reg n_n2485;

reg n_n2495;

reg pksi_97_;

reg pksi_102_;

reg pksi_11_;

reg pksi_173_;

reg pksi_179_;

reg pksi_171_;

reg pksi_104_;

reg pksi_103_;

reg n_n2384;

reg pksi_183_;

reg pksi_172_;

reg n_n2416;

reg pksi_116_;

reg pksi_96_;

reg pksi_119_;

reg pksi_84_;

reg pksi_159_;

reg n_n2440;

reg pksi_160_;

reg pksi_128_;

reg pksi_127_;

reg pksi_142_;

reg n_n2272;

reg pksi_149_;

reg pksi_162_;

reg pksi_154_;

reg pksi_121_;

reg pksi_134_;

reg pksi_126_;

reg pksi_82_;

reg n_n2430;

reg pksi_153_;

reg pksi_165_;

reg pksi_137_;

reg n_n2481;

reg pksi_101_;

reg pksi_93_;

reg pksi_161_;

reg pksi_156_;

reg n_n2452;

reg n_n2462;

reg pksi_123_;

reg pksi_111_;

reg pksi_92_;

reg pksi_15_;

reg n_n109;

reg pksi_145_;

reg pksi_144_;

reg pksi_150_;

reg pksi_124_;

reg pksi_132_;

reg pksi_130_;

reg pksi_105_;

reg pksi_112_;

reg n_n10;

reg pksi_6_;

reg pksi_188_;

reg pksi_152_;

reg pksi_163_;

reg pksi_166_;

reg pksi_131_;

reg n_n2474;

reg pksi_136_;

reg pksi_108_;

reg n_n2517;

reg n_n2268;

reg pksi_175_;

reg pksi_190_;

reg pksi_164_;

reg pksi_158_;

reg pksi_167_;

reg pksi_133_;

reg n_n2476;

reg pksi_122_;

reg n_n2507;

reg pksi_75_;

reg pksi_182_;

reg pksi_174_;

reg pksi_157_;

reg pksi_151_;

reg pksi_146_;

reg pksi_140_;

reg pksi_120_;

reg n_n168;

reg pksi_106_;

reg pksi_57_;

reg pksi_36_;

reg pksi_38_;

reg pksi_28_;

reg n_n2374;

reg pksi_53_;

reg pksi_27_;

reg pksi_26_;

reg pksi_47_;

reg pksi_1_;

reg pksi_63_;

reg pksi_34_;

reg pksi_24_;

reg pksi_30_;

reg pksi_18_;

reg pksi_79_;

reg pksi_54_;

reg n_n2337;

reg pksi_46_;

reg pksi_39_;

reg pksi_8_;

reg n_n2277;

reg pksi_91_;

reg pksi_51_;

reg pksi_70_;

reg pksi_0_;

reg pksi_73_;

reg pksi_89_;

reg pksi_60_;

reg pksi_48_;

reg pksi_22_;

reg n_n2280;

reg pksi_77_;

reg pksi_64_;

reg pksi_56_;

reg pksi_80_;

reg pksi_81_;

reg n_n2301;

reg pksi_66_;

reg pksi_72_;

reg pksi_78_;

reg pksi_69_;

reg n_n2320;

reg pksi_40_;

reg pksi_32_;

reg pksi_94_;

reg pksi_87_;

reg pksi_61_;

reg pksi_59_;

reg n_n2333;

reg pksi_42_;

reg pksi_86_;

reg pksi_76_;

reg n_n2305;

reg pksi_50_;

reg pksi_33_;

reg pksi_12_;

reg pksi_74_;

reg pksi_95_;

reg pksi_58_;

reg pksi_62_;

reg pksi_29_;

reg pksi_3_;

reg pksi_83_;

reg pksi_68_;

reg pksi_71_;

reg pksi_37_;

reg pksi_41_;

reg n_n2365;

reg n_n2369;

reg n_n2288;

reg pksi_55_;

reg pksi_52_;

reg pksi_45_;

reg pksi_43_;

reg pksi_16_;

reg pksi_10_;

reg n_n2310;

reg pksi_67_;

reg pksi_31_;

reg pksi_25_;

reg pksi_35_;

reg pksi_20_;

reg pksi_21_;

reg pksi_49_;

reg pksi_65_;

reg pksi_44_;

reg n_n2342;

reg n_n2352;

reg pksi_7_;

reg pksi_13_;

always  @(posedge pclk)
	pksi_17_<=n_n2385;

 always  @(posedge pclk)
	pksi_185_<=n_n2397;

 always  @(posedge pclk)
	n_n2410<=n_n2409;

 always  @(posedge pclk)
	pksi_170_<=n_n2424;

 always  @(posedge pclk)
	pksi_155_<=n_n2436;

 always  @(posedge pclk)
	pksi_147_<=n_n2449;

 always  @(posedge pclk)
	pksi_109_<=n_n2500;

 always  @(posedge pclk)
	n_n2513<=n_n2512;

 always  @(posedge pclk)
	pksi_19_<=n_n2386;

 always  @(posedge pclk)
	n_n2396<=n_n2395;

 always  @(posedge pclk)
	n_n2412<=n_n2411;

 always  @(posedge pclk)
	n_n121<=n_n2423;

 always  @(posedge pclk)
	pksi_148_<=n_n2437;

 always  @(posedge pclk)
	n_n2448<=n_n2447;

 always  @(posedge pclk)
	pksi_107_<=n_n2501;

 always  @(posedge pclk)
	pksi_110_<=n_n2511;

 always  @(posedge pclk)
	pksi_9_<=n_n2387;

 always  @(posedge pclk)
	pksi_176_<=n_n2399;

 always  @(posedge pclk)
	pksi_180_<=n_n2406;

 always  @(posedge pclk)
	pksi_178_<=n_n2422;

 always  @(posedge pclk)
	pksi_135_<=n_n2459;

 always  @(posedge pclk)
	pksi_129_<=n_n2471;

 always  @(posedge pclk)
	pksi_100_<=n_n2502;

 always  @(posedge pclk)
	pksi_117_<=n_n2515;

 always  @(posedge pclk)
	pksi_118_<=n_n2523;

 always  @(posedge pclk)
	pksi_5_<=n_n2388;

 always  @(posedge pclk)
	pksi_169_<=n_n2398;

 always  @(posedge pclk)
	n_n2408<=n_n2407;

 always  @(posedge pclk)
	pksi_184_<=n_n2421;

 always  @(posedge pclk)
	pksi_125_<=n_n2460;

 always  @(posedge pclk)
	pksi_138_<=n_n2470;

 always  @(posedge pclk)
	pksi_114_<=n_n2503;

 always  @(posedge pclk)
	pksi_99_<=n_n2514;

 always  @(posedge pclk)
	pksi_85_<=n_n2275;

 always  @(posedge pclk)
	pksi_14_<=n_n2380;

 always  @(posedge pclk)
	pksi_4_<=n_n2392;

 always  @(posedge pclk)
	pksi_186_<=n_n2404;

 always  @(posedge pclk)
	n_n2420<=n_n2419;

 always  @(posedge pclk)
	pksi_141_<=n_n2483;

 always  @(posedge pclk)
	pksi_113_<=n_n2496;

 always  @(posedge pclk)
	pksi_115_<=n_n2508;

 always  @(posedge pclk)
	pksi_98_<=n_n2521;

 always  @(posedge pclk)
	pksi_2_<=n_n2381;

 always  @(posedge pclk)
	pksi_23_<=n_n2391;

 always  @(posedge pclk)
	pksi_177_<=n_n2405;

 always  @(posedge pclk)
	pksi_189_<=n_n2418;

 always  @(posedge pclk)
	n_n2485<=n_n2484;

 always  @(posedge pclk)
	n_n2495<=n_n2494;

 always  @(posedge pclk)
	pksi_97_<=n_n2497;

 always  @(posedge pclk)
	pksi_102_<=n_n2522;

 always  @(posedge pclk)
	pksi_11_<=n_n2382;

 always  @(posedge pclk)
	pksi_173_<=n_n2394;

 always  @(posedge pclk)
	pksi_179_<=n_n2402;

 always  @(posedge pclk)
	pksi_171_<=n_n2417;

 always  @(posedge pclk)
	pksi_104_<=n_n2498;

 always  @(posedge pclk)
	pksi_103_<=n_n2510;

 always  @(posedge pclk)
	n_n2384<=n_n2383;

 always  @(posedge pclk)
	pksi_183_<=n_n2393;

 always  @(posedge pclk)
	pksi_172_<=n_n2403;

 always  @(posedge pclk)
	n_n2416<=n_n2415;

 always  @(posedge pclk)
	pksi_116_<=n_n2499;

 always  @(posedge pclk)
	pksi_96_<=n_n2509;

 always  @(posedge pclk)
	pksi_119_<=n_n2520;

 always  @(posedge pclk)
	pksi_84_<=n_n2270;

 always  @(posedge pclk)
	pksi_159_<=n_n2427;

 always  @(posedge pclk)
	n_n2440<=n_n2439;

 always  @(posedge pclk)
	pksi_160_<=n_n2453;

 always  @(posedge pclk)
	pksi_128_<=n_n2465;

 always  @(posedge pclk)
	pksi_127_<=n_n2478;

 always  @(posedge pclk)
	pksi_142_<=n_n2491;

 always  @(posedge pclk)
	n_n2272<=n_n2271;

 always  @(posedge pclk)
	pksi_149_<=n_n2428;

 always  @(posedge pclk)
	pksi_162_<=n_n2438;

 always  @(posedge pclk)
	pksi_154_<=n_n2454;

 always  @(posedge pclk)
	pksi_121_<=n_n2464;

 always  @(posedge pclk)
	pksi_134_<=n_n2479;

 always  @(posedge pclk)
	pksi_126_<=n_n2490;

 always  @(posedge pclk)
	pksi_82_<=n_n2273;

 always  @(posedge pclk)
	n_n2430<=n_n2429;

 always  @(posedge pclk)
	pksi_153_<=n_n2442;

 always  @(posedge pclk)
	pksi_165_<=n_n2450;

 always  @(posedge pclk)
	pksi_137_<=n_n2463;

 always  @(posedge pclk)
	n_n2481<=n_n2480;

 always  @(posedge pclk)
	pksi_101_<=n_n2493;

 always  @(posedge pclk)
	pksi_93_<=n_n2274;

 always  @(posedge pclk)
	pksi_161_<=n_n2431;

 always  @(posedge pclk)
	pksi_156_<=n_n2441;

 always  @(posedge pclk)
	n_n2452<=n_n2451;

 always  @(posedge pclk)
	n_n2462<=n_n2461;

 always  @(posedge pclk)
	pksi_123_<=n_n2482;

 always  @(posedge pclk)
	pksi_111_<=n_n2492;

 always  @(posedge pclk)
	pksi_92_<=n_n2265;

 always  @(posedge pclk)
	pksi_15_<=n_n2389;

 always  @(posedge pclk)
	n_n109<=n_n2401;

 always  @(posedge pclk)
	pksi_145_<=n_n2432;

 always  @(posedge pclk)
	pksi_144_<=n_n2444;

 always  @(posedge pclk)
	pksi_150_<=n_n2457;

 always  @(posedge pclk)
	pksi_124_<=n_n2469;

 always  @(posedge pclk)
	pksi_132_<=n_n2472;

 always  @(posedge pclk)
	pksi_130_<=n_n2487;

 always  @(posedge pclk)
	pksi_105_<=n_n2504;

 always  @(posedge pclk)
	pksi_112_<=n_n2518;

 always  @(posedge pclk)
	n_n10<=n_n2266;

 always  @(posedge pclk)
	pksi_6_<=n_n2390;

 always  @(posedge pclk)
	pksi_188_<=n_n2400;

 always  @(posedge pclk)
	pksi_152_<=n_n2433;

 always  @(posedge pclk)
	pksi_163_<=n_n2443;

 always  @(posedge pclk)
	pksi_166_<=n_n2458;

 always  @(posedge pclk)
	pksi_131_<=n_n2468;

 always  @(posedge pclk)
	n_n2474<=n_n2473;

 always  @(posedge pclk)
	pksi_136_<=n_n2486;

 always  @(posedge pclk)
	pksi_108_<=n_n2505;

 always  @(posedge pclk)
	n_n2517<=n_n2516;

 always  @(posedge pclk)
	n_n2268<=n_n2267;

 always  @(posedge pclk)
	pksi_175_<=n_n2413;

 always  @(posedge pclk)
	pksi_190_<=n_n2426;

 always  @(posedge pclk)
	pksi_164_<=n_n2434;

 always  @(posedge pclk)
	pksi_158_<=n_n2446;

 always  @(posedge pclk)
	pksi_167_<=n_n2455;

 always  @(posedge pclk)
	pksi_133_<=n_n2467;

 always  @(posedge pclk)
	n_n2476<=n_n2475;

 always  @(posedge pclk)
	pksi_122_<=n_n2489;

 always  @(posedge pclk)
	n_n2507<=n_n2506;

 always  @(posedge pclk)
	pksi_75_<=n_n2269;

 always  @(posedge pclk)
	pksi_182_<=n_n2414;

 always  @(posedge pclk)
	pksi_174_<=n_n2425;

 always  @(posedge pclk)
	pksi_157_<=n_n2435;

 always  @(posedge pclk)
	pksi_151_<=n_n2445;

 always  @(posedge pclk)
	pksi_146_<=n_n2456;

 always  @(posedge pclk)
	pksi_140_<=n_n2466;

 always  @(posedge pclk)
	pksi_120_<=n_n2477;

 always  @(posedge pclk)
	n_n168<=n_n2488;

 always  @(posedge pclk)
	pksi_106_<=n_n2519;

 always  @(posedge pclk)
	pksi_57_<=n_n2323;

 always  @(posedge pclk)
	pksi_36_<=n_n2335;

 always  @(posedge pclk)
	pksi_38_<=n_n2348;

 always  @(posedge pclk)
	pksi_28_<=n_n2360;

 always  @(posedge pclk)
	n_n2374<=n_n2373;

 always  @(posedge pclk)
	pksi_53_<=n_n2324;

 always  @(posedge pclk)
	pksi_27_<=n_n2334;

 always  @(posedge pclk)
	pksi_26_<=n_n2349;

 always  @(posedge pclk)
	pksi_47_<=n_n2359;

 always  @(posedge pclk)
	pksi_1_<=n_n2375;

 always  @(posedge pclk)
	pksi_63_<=n_n2325;

 always  @(posedge pclk)
	pksi_34_<=n_n2338;

 always  @(posedge pclk)
	pksi_24_<=n_n2346;

 always  @(posedge pclk)
	pksi_30_<=n_n2358;

 always  @(posedge pclk)
	pksi_18_<=n_n2376;

 always  @(posedge pclk)
	pksi_79_<=n_n2264;

 always  @(posedge pclk)
	pksi_54_<=n_n2326;

 always  @(posedge pclk)
	n_n2337<=n_n2336;

 always  @(posedge pclk)
	pksi_46_<=n_n2347;

 always  @(posedge pclk)
	pksi_39_<=n_n2357;

 always  @(posedge pclk)
	pksi_8_<=n_n2377;

 always  @(posedge pclk)
	n_n2277<=n_n2276;

 always  @(posedge pclk)
	pksi_91_<=n_n2290;

 always  @(posedge pclk)
	pksi_51_<=n_n2302;

 always  @(posedge pclk)
	pksi_70_<=n_n2315;

 always  @(posedge pclk)
	pksi_0_<=n_n2378;

 always  @(posedge pclk)
	pksi_73_<=n_n2278;

 always  @(posedge pclk)
	pksi_89_<=n_n2289;

 always  @(posedge pclk)
	pksi_60_<=n_n2303;

 always  @(posedge pclk)
	pksi_48_<=n_n2314;

 always  @(posedge pclk)
	pksi_22_<=n_n2379;

 always  @(posedge pclk)
	n_n2280<=n_n2279;

 always  @(posedge pclk)
	pksi_77_<=n_n2292;

 always  @(posedge pclk)
	pksi_64_<=n_n2299;

 always  @(posedge pclk)
	pksi_56_<=n_n2313;

 always  @(posedge pclk)
	pksi_80_<=n_n2281;

 always  @(posedge pclk)
	pksi_81_<=n_n2291;

 always  @(posedge pclk)
	n_n2301<=n_n2300;

 always  @(posedge pclk)
	pksi_66_<=n_n2312;

 always  @(posedge pclk)
	pksi_72_<=n_n2282;

 always  @(posedge pclk)
	pksi_78_<=n_n2294;

 always  @(posedge pclk)
	pksi_69_<=n_n2307;

 always  @(posedge pclk)
	n_n2320<=n_n2319;

 always  @(posedge pclk)
	pksi_40_<=n_n2331;

 always  @(posedge pclk)
	pksi_32_<=n_n2345;

 always  @(posedge pclk)
	pksi_94_<=n_n2283;

 always  @(posedge pclk)
	pksi_87_<=n_n2293;

 always  @(posedge pclk)
	pksi_61_<=n_n2308;

 always  @(posedge pclk)
	pksi_59_<=n_n2318;

 always  @(posedge pclk)
	n_n2333<=n_n2332;

 always  @(posedge pclk)
	pksi_42_<=n_n2344;

 always  @(posedge pclk)
	pksi_86_<=n_n2284;

 always  @(posedge pclk)
	pksi_76_<=n_n2296;

 always  @(posedge pclk)
	n_n2305<=n_n2304;

 always  @(posedge pclk)
	pksi_50_<=n_n2317;

 always  @(posedge pclk)
	pksi_33_<=n_n2355;

 always  @(posedge pclk)
	pksi_12_<=n_n2367;

 always  @(posedge pclk)
	pksi_74_<=n_n2285;

 always  @(posedge pclk)
	pksi_95_<=n_n2295;

 always  @(posedge pclk)
	pksi_58_<=n_n2306;

 always  @(posedge pclk)
	pksi_62_<=n_n2316;

 always  @(posedge pclk)
	pksi_29_<=n_n2356;

 always  @(posedge pclk)
	pksi_3_<=n_n2366;

 always  @(posedge pclk)
	pksi_83_<=n_n2286;

 always  @(posedge pclk)
	pksi_68_<=n_n2298;

 always  @(posedge pclk)
	pksi_71_<=n_n2327;

 always  @(posedge pclk)
	pksi_37_<=n_n2340;

 always  @(posedge pclk)
	pksi_41_<=n_n2353;

 always  @(posedge pclk)
	n_n2365<=n_n2364;

 always  @(posedge pclk)
	n_n2369<=n_n2368;

 always  @(posedge pclk)
	n_n2288<=n_n2287;

 always  @(posedge pclk)
	pksi_55_<=n_n2297;

 always  @(posedge pclk)
	pksi_52_<=n_n2328;

 always  @(posedge pclk)
	pksi_45_<=n_n2339;

 always  @(posedge pclk)
	pksi_43_<=n_n2354;

 always  @(posedge pclk)
	pksi_16_<=n_n2363;

 always  @(posedge pclk)
	pksi_10_<=n_n2370;

 always  @(posedge pclk)
	n_n2310<=n_n2309;

 always  @(posedge pclk)
	pksi_67_<=n_n2322;

 always  @(posedge pclk)
	pksi_31_<=n_n2329;

 always  @(posedge pclk)
	pksi_25_<=n_n2343;

 always  @(posedge pclk)
	pksi_35_<=n_n2350;

 always  @(posedge pclk)
	pksi_20_<=n_n2362;

 always  @(posedge pclk)
	pksi_21_<=n_n2371;

 always  @(posedge pclk)
	pksi_49_<=n_n2311;

 always  @(posedge pclk)
	pksi_65_<=n_n2321;

 always  @(posedge pclk)
	pksi_44_<=n_n2330;

 always  @(posedge pclk)
	n_n2342<=n_n2341;

 always  @(posedge pclk)
	n_n2352<=n_n2351;

 always  @(posedge pclk)
	pksi_7_<=n_n2361;

 always  @(posedge pclk)
	pksi_13_<=n_n2372;

 assign pdata_ready_0_ = ( n_n204  &  wire653 ) | ( n_n200  &  wire7079 ) ;
 assign pnew_count_3_ = ( wire669 ) | ( wire670 ) | ( pstart_0_  &  (~ pencrypt_0_) ) ;
 assign pnew_count_0_ = ( (~ pcount_0_)  &  (~ pstart_0_) ) | ( pstart_0_  &  (~ pencrypt_0_) ) ;
 assign pnew_count_2_ = ( wire7084 ) | ( pcount_2_  &  (~ wire647) ) ;
 assign pnew_count_1_ = ( pstart_0_  &  (~ pencrypt_0_) ) | ( pcount_1_  &  pcount_0_  &  (~ pencrypt_0_) ) | ( (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) | ( (~ pcount_1_)  &  pcount_0_  &  (~ pstart_0_)  &  pencrypt_0_ ) | ( pcount_1_  &  (~ pcount_0_)  &  (~ pstart_0_)  &  pencrypt_0_ ) ;
 assign n_n2385 = ( wire2021 ) | ( wire2024 ) | ( wire2025 ) | ( wire6183 ) ;
 assign n_n2397 = ( wire2015 ) | ( wire2018 ) | ( wire2019 ) | ( wire6187 ) ;
 assign n_n2409 = ( wire2009 ) | ( wire2012 ) | ( wire2013 ) | ( wire6191 ) ;
 assign n_n2424 = ( wire2003 ) | ( wire2006 ) | ( wire2007 ) | ( wire6195 ) ;
 assign n_n2436 = ( wire1997 ) | ( wire2000 ) | ( wire2001 ) | ( wire6199 ) ;
 assign n_n2449 = ( wire1991 ) | ( wire1994 ) | ( wire1995 ) | ( wire6203 ) ;
 assign n_n2500 = ( wire1985 ) | ( wire1988 ) | ( wire1989 ) | ( wire6207 ) ;
 assign n_n2512 = ( wire1979 ) | ( wire1982 ) | ( wire1983 ) | ( wire6211 ) ;
 assign n_n2386 = ( wire1973 ) | ( wire1976 ) | ( wire1977 ) | ( wire6215 ) ;
 assign n_n2395 = ( wire1967 ) | ( wire1970 ) | ( wire1971 ) | ( wire6219 ) ;
 assign n_n2411 = ( wire1961 ) | ( wire1964 ) | ( wire1965 ) | ( wire6223 ) ;
 assign n_n2423 = ( wire1955 ) | ( wire1958 ) | ( wire1959 ) | ( wire6227 ) ;
 assign n_n2437 = ( wire1949 ) | ( wire1952 ) | ( wire1953 ) | ( wire6231 ) ;
 assign n_n2447 = ( wire1943 ) | ( wire1946 ) | ( wire1947 ) | ( wire6235 ) ;
 assign n_n2501 = ( wire1937 ) | ( wire1940 ) | ( wire1941 ) | ( wire6239 ) ;
 assign n_n2511 = ( wire1931 ) | ( wire1934 ) | ( wire1935 ) | ( wire6243 ) ;
 assign n_n2387 = ( wire1925 ) | ( wire1928 ) | ( wire1929 ) | ( wire6247 ) ;
 assign n_n2399 = ( wire1919 ) | ( wire1922 ) | ( wire1923 ) | ( wire6251 ) ;
 assign n_n2406 = ( wire1913 ) | ( wire1916 ) | ( wire1917 ) | ( wire6255 ) ;
 assign n_n2422 = ( wire1907 ) | ( wire1910 ) | ( wire1911 ) | ( wire6259 ) ;
 assign n_n2459 = ( wire1901 ) | ( wire1904 ) | ( wire1905 ) | ( wire6263 ) ;
 assign n_n2471 = ( wire1894 ) | ( wire1898 ) | ( wire1899 ) | ( wire6267 ) ;
 assign n_n2502 = ( wire1889 ) | ( wire1892 ) | ( wire1893 ) | ( wire6271 ) ;
 assign n_n2515 = ( wire1883 ) | ( wire1885 ) | ( wire1887 ) | ( wire6275 ) ;
 assign n_n2523 = ( wire1877 ) | ( wire1880 ) | ( wire1881 ) | ( wire6279 ) ;
 assign n_n2388 = ( wire1871 ) | ( wire1874 ) | ( wire1875 ) | ( wire6283 ) ;
 assign n_n2398 = ( wire1865 ) | ( wire1868 ) | ( wire1869 ) | ( wire6287 ) ;
 assign n_n2407 = ( wire1859 ) | ( wire1862 ) | ( wire1863 ) | ( wire6291 ) ;
 assign n_n2421 = ( wire1853 ) | ( wire1856 ) | ( wire1857 ) | ( wire6295 ) ;
 assign n_n2460 = ( wire1847 ) | ( wire1848 ) | ( wire1851 ) | ( wire6299 ) ;
 assign n_n2470 = ( wire1841 ) | ( wire1844 ) | ( wire1845 ) | ( wire6303 ) ;
 assign n_n2503 = ( wire1835 ) | ( wire1838 ) | ( wire1839 ) | ( wire6307 ) ;
 assign n_n2514 = ( wire1829 ) | ( wire1832 ) | ( wire1833 ) | ( wire6311 ) ;
 assign n_n2275 = ( wire1822 ) | ( wire1824 ) | ( wire1827 ) | ( wire6315 ) ;
 assign n_n2380 = ( wire1817 ) | ( wire1820 ) | ( wire1821 ) | ( wire6319 ) ;
 assign n_n2392 = ( wire1811 ) | ( wire1814 ) | ( wire1815 ) | ( wire6323 ) ;
 assign n_n2404 = ( wire1805 ) | ( wire1808 ) | ( wire1809 ) | ( wire6327 ) ;
 assign n_n2419 = ( wire1799 ) | ( wire1802 ) | ( wire1803 ) | ( wire6331 ) ;
 assign n_n2483 = ( wire1793 ) | ( wire1796 ) | ( wire1797 ) | ( wire6335 ) ;
 assign n_n2496 = ( wire1787 ) | ( wire1790 ) | ( wire1791 ) | ( wire6339 ) ;
 assign n_n2508 = ( wire1781 ) | ( wire1784 ) | ( wire1785 ) | ( wire6343 ) ;
 assign n_n2521 = ( wire1775 ) | ( wire1778 ) | ( wire1779 ) | ( wire6347 ) ;
 assign n_n2381 = ( wire1769 ) | ( wire1772 ) | ( wire1773 ) | ( wire6351 ) ;
 assign n_n2391 = ( wire1763 ) | ( wire1766 ) | ( wire1767 ) | ( wire6355 ) ;
 assign n_n2405 = ( wire1757 ) | ( wire1760 ) | ( wire1761 ) | ( wire6359 ) ;
 assign n_n2418 = ( wire1751 ) | ( wire1754 ) | ( wire1755 ) | ( wire6363 ) ;
 assign n_n2484 = ( wire1745 ) | ( wire1748 ) | ( wire1749 ) | ( wire6367 ) ;
 assign n_n2494 = ( wire1739 ) | ( wire1742 ) | ( wire1743 ) | ( wire6371 ) ;
 assign n_n2497 = ( wire1733 ) | ( wire1736 ) | ( wire1737 ) | ( wire6375 ) ;
 assign n_n2522 = ( wire1727 ) | ( wire1730 ) | ( wire1731 ) | ( wire6379 ) ;
 assign n_n2382 = ( wire1721 ) | ( wire1724 ) | ( wire1725 ) | ( wire6383 ) ;
 assign n_n2394 = ( wire1715 ) | ( wire1718 ) | ( wire1719 ) | ( wire6387 ) ;
 assign n_n2402 = ( wire1709 ) | ( wire1712 ) | ( wire1713 ) | ( wire6391 ) ;
 assign n_n2417 = ( wire1703 ) | ( wire1706 ) | ( wire1707 ) | ( wire6395 ) ;
 assign n_n2498 = ( wire1697 ) | ( wire1700 ) | ( wire1701 ) | ( wire6399 ) ;
 assign n_n2510 = ( wire1691 ) | ( wire1694 ) | ( wire1695 ) | ( wire6403 ) ;
 assign n_n2383 = ( wire1685 ) | ( wire1688 ) | ( wire1689 ) | ( wire6407 ) ;
 assign n_n2393 = ( wire1679 ) | ( wire1682 ) | ( wire1683 ) | ( wire6411 ) ;
 assign n_n2403 = ( wire1673 ) | ( wire1676 ) | ( wire1677 ) | ( wire6415 ) ;
 assign n_n2415 = ( wire1667 ) | ( wire1670 ) | ( wire1671 ) | ( wire6419 ) ;
 assign n_n2499 = ( wire1661 ) | ( wire1664 ) | ( wire1665 ) | ( wire6423 ) ;
 assign n_n2509 = ( wire1655 ) | ( wire1658 ) | ( wire1659 ) | ( wire6427 ) ;
 assign n_n2520 = ( wire1649 ) | ( wire1652 ) | ( wire1653 ) | ( wire6431 ) ;
 assign n_n2270 = ( wire1644 ) | ( wire1646 ) | ( wire1647 ) | ( wire6435 ) ;
 assign n_n2427 = ( wire1637 ) | ( wire1640 ) | ( wire1641 ) | ( wire6439 ) ;
 assign n_n2439 = ( wire1631 ) | ( wire1634 ) | ( wire1635 ) | ( wire6443 ) ;
 assign n_n2453 = ( wire1626 ) | ( wire1628 ) | ( wire1629 ) | ( wire6447 ) ;
 assign n_n2465 = ( wire1619 ) | ( wire1622 ) | ( wire1623 ) | ( wire6451 ) ;
 assign n_n2478 = ( wire1613 ) | ( wire1616 ) | ( wire1617 ) | ( wire6455 ) ;
 assign n_n2491 = ( wire1607 ) | ( wire1610 ) | ( wire1611 ) | ( wire6459 ) ;
 assign n_n2271 = ( wire1601 ) | ( wire1604 ) | ( wire1605 ) | ( wire6463 ) ;
 assign n_n2428 = ( wire1595 ) | ( wire1596 ) | ( wire1599 ) | ( wire6467 ) ;
 assign n_n2438 = ( wire1589 ) | ( wire1592 ) | ( wire1593 ) | ( wire6471 ) ;
 assign n_n2454 = ( wire1584 ) | ( wire1586 ) | ( wire1587 ) | ( wire6475 ) ;
 assign n_n2464 = ( wire1578 ) | ( wire1580 ) | ( wire1581 ) | ( wire6479 ) ;
 assign n_n2479 = ( wire1571 ) | ( wire1572 ) | ( wire1575 ) | ( wire6483 ) ;
 assign n_n2490 = ( wire1565 ) | ( wire1568 ) | ( wire1569 ) | ( wire6487 ) ;
 assign n_n2273 = ( wire1559 ) | ( wire1562 ) | ( wire1563 ) | ( wire6491 ) ;
 assign n_n2429 = ( wire1553 ) | ( wire1556 ) | ( wire1557 ) | ( wire6495 ) ;
 assign n_n2442 = ( wire1547 ) | ( wire1550 ) | ( wire1551 ) | ( wire6499 ) ;
 assign n_n2450 = ( wire1541 ) | ( wire1542 ) | ( wire1545 ) | ( wire6503 ) ;
 assign n_n2463 = ( wire1536 ) | ( wire1538 ) | ( wire1539 ) | ( wire6507 ) ;
 assign n_n2480 = ( wire1529 ) | ( wire1532 ) | ( wire1533 ) | ( wire6511 ) ;
 assign n_n2493 = ( wire1523 ) | ( wire1526 ) | ( wire1527 ) | ( wire6515 ) ;
 assign n_n2274 = ( wire1516 ) | ( wire1520 ) | ( wire1521 ) | ( wire6519 ) ;
 assign n_n2431 = ( wire1511 ) | ( wire1514 ) | ( wire1515 ) | ( wire6523 ) ;
 assign n_n2441 = ( wire1505 ) | ( wire1508 ) | ( wire1509 ) | ( wire6527 ) ;
 assign n_n2451 = ( wire1499 ) | ( wire1502 ) | ( wire1503 ) | ( wire6531 ) ;
 assign n_n2461 = ( wire1493 ) | ( wire1496 ) | ( wire1497 ) | ( wire6535 ) ;
 assign n_n2482 = ( wire1487 ) | ( wire1490 ) | ( wire1491 ) | ( wire6539 ) ;
 assign n_n2492 = ( wire1481 ) | ( wire1484 ) | ( wire1485 ) | ( wire6543 ) ;
 assign n_n2265 = ( wire1474 ) | ( wire1478 ) | ( wire1479 ) | ( wire6547 ) ;
 assign n_n2389 = ( wire1469 ) | ( wire1472 ) | ( wire1473 ) | ( wire6551 ) ;
 assign n_n2401 = ( wire1463 ) | ( wire1466 ) | ( wire1467 ) | ( wire6555 ) ;
 assign n_n2432 = ( wire1457 ) | ( wire1460 ) | ( wire1461 ) | ( wire6559 ) ;
 assign n_n2444 = ( wire1451 ) | ( wire1454 ) | ( wire1455 ) | ( wire6563 ) ;
 assign n_n2457 = ( wire1445 ) | ( wire1448 ) | ( wire1449 ) | ( wire6567 ) ;
 assign n_n2469 = ( wire1439 ) | ( wire1442 ) | ( wire1443 ) | ( wire6571 ) ;
 assign n_n2472 = ( wire1432 ) | ( wire1434 ) | ( wire1437 ) | ( wire6575 ) ;
 assign n_n2487 = ( wire1427 ) | ( wire1430 ) | ( wire1431 ) | ( wire6579 ) ;
 assign n_n2504 = ( wire1421 ) | ( wire1424 ) | ( wire1425 ) | ( wire6583 ) ;
 assign n_n2518 = ( wire1415 ) | ( wire1418 ) | ( wire1419 ) | ( wire6587 ) ;
 assign n_n2266 = ( wire1408 ) | ( wire1410 ) | ( wire1413 ) | ( wire6591 ) ;
 assign n_n2390 = ( wire1403 ) | ( wire1406 ) | ( wire1407 ) | ( wire6595 ) ;
 assign n_n2400 = ( wire1397 ) | ( wire1400 ) | ( wire1401 ) | ( wire6599 ) ;
 assign n_n2433 = ( wire1391 ) | ( wire1394 ) | ( wire1395 ) | ( wire6603 ) ;
 assign n_n2443 = ( wire1385 ) | ( wire1388 ) | ( wire1389 ) | ( wire6607 ) ;
 assign n_n2458 = ( wire1379 ) | ( wire1382 ) | ( wire1383 ) | ( wire6611 ) ;
 assign n_n2468 = ( wire1373 ) | ( wire1376 ) | ( wire1377 ) | ( wire6615 ) ;
 assign n_n2473 = ( wire1367 ) | ( wire1368 ) | ( wire1371 ) | ( wire6619 ) ;
 assign n_n2486 = ( wire1361 ) | ( wire1364 ) | ( wire1365 ) | ( wire6623 ) ;
 assign n_n2505 = ( wire1355 ) | ( wire1357 ) | ( wire1359 ) | ( wire6627 ) ;
 assign n_n2516 = ( wire1349 ) | ( wire1352 ) | ( wire1353 ) | ( wire6631 ) ;
 assign n_n2267 = ( wire1343 ) | ( wire1346 ) | ( wire1347 ) | ( wire6635 ) ;
 assign n_n2413 = ( wire1337 ) | ( wire1340 ) | ( wire1341 ) | ( wire6639 ) ;
 assign n_n2426 = ( wire1331 ) | ( wire1334 ) | ( wire1335 ) | ( wire6643 ) ;
 assign n_n2434 = ( wire1325 ) | ( wire1328 ) | ( wire1329 ) | ( wire6647 ) ;
 assign n_n2446 = ( wire1319 ) | ( wire1322 ) | ( wire1323 ) | ( wire6651 ) ;
 assign n_n2455 = ( wire1313 ) | ( wire1316 ) | ( wire1317 ) | ( wire6655 ) ;
 assign n_n2467 = ( wire1307 ) | ( wire1310 ) | ( wire1311 ) | ( wire6659 ) ;
 assign n_n2475 = ( wire1302 ) | ( wire1304 ) | ( wire1305 ) | ( wire6663 ) ;
 assign n_n2489 = ( wire1295 ) | ( wire1298 ) | ( wire1299 ) | ( wire6667 ) ;
 assign n_n2506 = ( wire1289 ) | ( wire1292 ) | ( wire1293 ) | ( wire6671 ) ;
 assign n_n2269 = ( wire1284 ) | ( wire1286 ) | ( wire1287 ) | ( wire6675 ) ;
 assign n_n2414 = ( wire1277 ) | ( wire1280 ) | ( wire1281 ) | ( wire6679 ) ;
 assign n_n2425 = ( wire1271 ) | ( wire1274 ) | ( wire1275 ) | ( wire6683 ) ;
 assign n_n2435 = ( wire1265 ) | ( wire1268 ) | ( wire1269 ) | ( wire6687 ) ;
 assign n_n2445 = ( wire1259 ) | ( wire1262 ) | ( wire1263 ) | ( wire6691 ) ;
 assign n_n2456 = ( wire1253 ) | ( wire1256 ) | ( wire1257 ) | ( wire6695 ) ;
 assign n_n2466 = ( wire1247 ) | ( wire1250 ) | ( wire1251 ) | ( wire6699 ) ;
 assign n_n2477 = ( wire1242 ) | ( wire1243 ) | ( wire1245 ) | ( wire6703 ) ;
 assign n_n2488 = ( wire1235 ) | ( wire1238 ) | ( wire1239 ) | ( wire6707 ) ;
 assign n_n2519 = ( wire1229 ) | ( wire1232 ) | ( wire1233 ) | ( wire6711 ) ;
 assign n_n2323 = ( wire1223 ) | ( wire1226 ) | ( wire1227 ) | ( wire6715 ) ;
 assign n_n2335 = ( wire1217 ) | ( wire1219 ) | ( wire1221 ) | ( wire6719 ) ;
 assign n_n2348 = ( wire1211 ) | ( wire1214 ) | ( wire1215 ) | ( wire6723 ) ;
 assign n_n2360 = ( wire1205 ) | ( wire1208 ) | ( wire1209 ) | ( wire6727 ) ;
 assign n_n2373 = ( wire1199 ) | ( wire1202 ) | ( wire1203 ) | ( wire6731 ) ;
 assign n_n2324 = ( wire1193 ) | ( wire1196 ) | ( wire1197 ) | ( wire6735 ) ;
 assign n_n2334 = ( wire1187 ) | ( wire1190 ) | ( wire1191 ) | ( wire6739 ) ;
 assign n_n2349 = ( wire1180 ) | ( wire1184 ) | ( wire1185 ) | ( wire6743 ) ;
 assign n_n2359 = ( wire1175 ) | ( wire1178 ) | ( wire1179 ) | ( wire6747 ) ;
 assign n_n2375 = ( wire1170 ) | ( wire1172 ) | ( wire1173 ) | ( wire6751 ) ;
 assign n_n2325 = ( wire1163 ) | ( wire1166 ) | ( wire1167 ) | ( wire6755 ) ;
 assign n_n2338 = ( wire1158 ) | ( wire1160 ) | ( wire1161 ) | ( wire6759 ) ;
 assign n_n2346 = ( wire1151 ) | ( wire1154 ) | ( wire1155 ) | ( wire6763 ) ;
 assign n_n2358 = ( wire1145 ) | ( wire1148 ) | ( wire1149 ) | ( wire6767 ) ;
 assign n_n2376 = ( wire1140 ) | ( wire1142 ) | ( wire1143 ) | ( wire6771 ) ;
 assign n_n2264 = ( wire1133 ) | ( wire1136 ) | ( wire1137 ) | ( wire6775 ) ;
 assign n_n2326 = ( wire1127 ) | ( wire1130 ) | ( wire1131 ) | ( wire6779 ) ;
 assign n_n2336 = ( wire1121 ) | ( wire1124 ) | ( wire1125 ) | ( wire6783 ) ;
 assign n_n2347 = ( wire1115 ) | ( wire1118 ) | ( wire1119 ) | ( wire6787 ) ;
 assign n_n2357 = ( wire1109 ) | ( wire1112 ) | ( wire1113 ) | ( wire6791 ) ;
 assign n_n2377 = ( wire1103 ) | ( wire1106 ) | ( wire1107 ) | ( wire6795 ) ;
 assign n_n2276 = ( wire1097 ) | ( wire1100 ) | ( wire1101 ) | ( wire6799 ) ;
 assign n_n2290 = ( wire1091 ) | ( wire1094 ) | ( wire1095 ) | ( wire6803 ) ;
 assign n_n2302 = ( wire1085 ) | ( wire1088 ) | ( wire1089 ) | ( wire6807 ) ;
 assign n_n2315 = ( wire1079 ) | ( wire1082 ) | ( wire1083 ) | ( wire6811 ) ;
 assign n_n2378 = ( wire1073 ) | ( wire1076 ) | ( wire1077 ) | ( wire6815 ) ;
 assign n_n2278 = ( wire1068 ) | ( wire1070 ) | ( wire1071 ) | ( wire6819 ) ;
 assign n_n2289 = ( wire1061 ) | ( wire1064 ) | ( wire1065 ) | ( wire6823 ) ;
 assign n_n2303 = ( wire1055 ) | ( wire1058 ) | ( wire1059 ) | ( wire6827 ) ;
 assign n_n2314 = ( wire1049 ) | ( wire1052 ) | ( wire1053 ) | ( wire6831 ) ;
 assign n_n2379 = ( wire1043 ) | ( wire1046 ) | ( wire1047 ) | ( wire6835 ) ;
 assign n_n2279 = ( wire1038 ) | ( wire1040 ) | ( wire1041 ) | ( wire6839 ) ;
 assign n_n2292 = ( wire1031 ) | ( wire1034 ) | ( wire1035 ) | ( wire6843 ) ;
 assign n_n2299 = ( wire1025 ) | ( wire1028 ) | ( wire1029 ) | ( wire6847 ) ;
 assign n_n2313 = ( wire1019 ) | ( wire1022 ) | ( wire1023 ) | ( wire6851 ) ;
 assign n_n2281 = ( wire1013 ) | ( wire1016 ) | ( wire1017 ) | ( wire6855 ) ;
 assign n_n2291 = ( wire1007 ) | ( wire1010 ) | ( wire1011 ) | ( wire6859 ) ;
 assign n_n2300 = ( wire1001 ) | ( wire1004 ) | ( wire1005 ) | ( wire6863 ) ;
 assign n_n2312 = ( wire995 ) | ( wire998 ) | ( wire999 ) | ( wire6867 ) ;
 assign n_n2282 = ( wire989 ) | ( wire992 ) | ( wire993 ) | ( wire6871 ) ;
 assign n_n2294 = ( wire983 ) | ( wire986 ) | ( wire987 ) | ( wire6875 ) ;
 assign n_n2307 = ( wire977 ) | ( wire980 ) | ( wire981 ) | ( wire6879 ) ;
 assign n_n2319 = ( wire971 ) | ( wire974 ) | ( wire975 ) | ( wire6883 ) ;
 assign n_n2331 = ( wire964 ) | ( wire966 ) | ( wire969 ) | ( wire6887 ) ;
 assign n_n2345 = ( wire959 ) | ( wire962 ) | ( wire963 ) | ( wire6891 ) ;
 assign n_n2283 = ( wire953 ) | ( wire956 ) | ( wire957 ) | ( wire6895 ) ;
 assign n_n2293 = ( wire947 ) | ( wire950 ) | ( wire951 ) | ( wire6899 ) ;
 assign n_n2308 = ( wire941 ) | ( wire944 ) | ( wire945 ) | ( wire6903 ) ;
 assign n_n2318 = ( wire934 ) | ( wire936 ) | ( wire939 ) | ( wire6907 ) ;
 assign n_n2332 = ( wire929 ) | ( wire932 ) | ( wire933 ) | ( wire6911 ) ;
 assign n_n2344 = ( wire924 ) | ( wire926 ) | ( wire927 ) | ( wire6915 ) ;
 assign n_n2284 = ( wire917 ) | ( wire920 ) | ( wire921 ) | ( wire6919 ) ;
 assign n_n2296 = ( wire911 ) | ( wire914 ) | ( wire915 ) | ( wire6923 ) ;
 assign n_n2304 = ( wire905 ) | ( wire908 ) | ( wire909 ) | ( wire6927 ) ;
 assign n_n2317 = ( wire898 ) | ( wire902 ) | ( wire903 ) | ( wire6931 ) ;
 assign n_n2355 = ( wire893 ) | ( wire896 ) | ( wire897 ) | ( wire6935 ) ;
 assign n_n2367 = ( wire886 ) | ( wire889 ) | ( wire891 ) | ( wire6939 ) ;
 assign n_n2285 = ( wire881 ) | ( wire884 ) | ( wire885 ) | ( wire6943 ) ;
 assign n_n2295 = ( wire875 ) | ( wire878 ) | ( wire879 ) | ( wire6947 ) ;
 assign n_n2306 = ( wire869 ) | ( wire872 ) | ( wire873 ) | ( wire6951 ) ;
 assign n_n2316 = ( wire863 ) | ( wire866 ) | ( wire867 ) | ( wire6955 ) ;
 assign n_n2356 = ( wire857 ) | ( wire860 ) | ( wire861 ) | ( wire6959 ) ;
 assign n_n2366 = ( wire850 ) | ( wire854 ) | ( wire855 ) | ( wire6963 ) ;
 assign n_n2286 = ( wire845 ) | ( wire848 ) | ( wire849 ) | ( wire6967 ) ;
 assign n_n2298 = ( wire839 ) | ( wire842 ) | ( wire843 ) | ( wire6971 ) ;
 assign n_n2327 = ( wire833 ) | ( wire836 ) | ( wire837 ) | ( wire6975 ) ;
 assign n_n2340 = ( wire826 ) | ( wire828 ) | ( wire831 ) | ( wire6979 ) ;
 assign n_n2353 = ( wire822 ) | ( wire824 ) | ( wire825 ) | ( wire6983 ) ;
 assign n_n2364 = ( wire815 ) | ( wire818 ) | ( wire819 ) | ( wire6987 ) ;
 assign n_n2368 = ( wire809 ) | ( wire812 ) | ( wire813 ) | ( wire6991 ) ;
 assign n_n2287 = ( wire803 ) | ( wire806 ) | ( wire807 ) | ( wire6995 ) ;
 assign n_n2297 = ( wire797 ) | ( wire800 ) | ( wire801 ) | ( wire6999 ) ;
 assign n_n2328 = ( wire791 ) | ( wire794 ) | ( wire795 ) | ( wire7003 ) ;
 assign n_n2339 = ( wire784 ) | ( wire788 ) | ( wire789 ) | ( wire7007 ) ;
 assign n_n2354 = ( wire780 ) | ( wire782 ) | ( wire783 ) | ( wire7011 ) ;
 assign n_n2363 = ( wire772 ) | ( wire774 ) | ( wire777 ) | ( wire7015 ) ;
 assign n_n2370 = ( wire768 ) | ( wire770 ) | ( wire771 ) | ( wire7019 ) ;
 assign n_n2309 = ( wire761 ) | ( wire764 ) | ( wire765 ) | ( wire7023 ) ;
 assign n_n2322 = ( wire756 ) | ( wire758 ) | ( wire759 ) | ( wire7027 ) ;
 assign n_n2329 = ( wire749 ) | ( wire752 ) | ( wire753 ) | ( wire7031 ) ;
 assign n_n2343 = ( wire744 ) | ( wire746 ) | ( wire747 ) | ( wire7035 ) ;
 assign n_n2350 = ( wire736 ) | ( wire738 ) | ( wire741 ) | ( wire7039 ) ;
 assign n_n2362 = ( wire730 ) | ( wire734 ) | ( wire735 ) | ( wire7043 ) ;
 assign n_n2371 = ( wire725 ) | ( wire728 ) | ( wire729 ) | ( wire7047 ) ;
 assign n_n2311 = ( wire719 ) | ( wire722 ) | ( wire723 ) | ( wire7051 ) ;
 assign n_n2321 = ( wire714 ) | ( wire716 ) | ( wire717 ) | ( wire7055 ) ;
 assign n_n2330 = ( wire706 ) | ( wire710 ) | ( wire711 ) | ( wire7059 ) ;
 assign n_n2341 = ( wire701 ) | ( wire704 ) | ( wire705 ) | ( wire7063 ) ;
 assign n_n2351 = ( wire695 ) | ( wire698 ) | ( wire699 ) | ( wire7067 ) ;
 assign n_n2361 = ( wire689 ) | ( wire692 ) | ( wire693 ) | ( wire7071 ) ;
 assign n_n2372 = ( wire682 ) | ( wire684 ) | ( wire687 ) | ( wire7075 ) ;
 assign n_n200 = ( (~ pcount_3_)  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) | ( pcount_3_  &  pcount_2_  &  pcount_1_  &  (~ pcount_0_) ) | ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_) ) ;
 assign n_n204 = ( (~ pcount_3_)  &  (~ pcount_2_)  &  (~ pcount_1_) ) | ( (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_) ) | ( pcount_3_  &  pcount_2_  &  pcount_1_  &  pcount_0_ ) ;
 assign wire653 = ( pcount_1_  &  pcount_0_  &  (~ pstart_0_)  &  pencrypt_0_ ) ;
 assign n_n2530 = ( (~ pstart_0_) ) | ( pencrypt_0_ ) ;
 assign wire647 = ( pstart_0_  &  pencrypt_0_ ) | ( pcount_1_  &  pcount_0_  &  pencrypt_0_ ) | ( (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) ;
 assign wire655 = ( (~ pstart_0_)  &  pencrypt_0_ ) ;
 assign pksi_90_ = ( n_n10 ) ;
 assign pksi_191_ = ( n_n121 ) ;
 assign pksi_187_ = ( n_n121 ) ;
 assign pksi_168_ = ( n_n109 ) ;
 assign pksi_181_ = ( n_n109 ) ;
 assign pksi_88_ = ( n_n10 ) ;
 assign pksi_143_ = ( n_n168 ) ;
 assign pksi_139_ = ( n_n168 ) ;
 assign wire664 = ( (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) ;
 assign wire669 = ( (~ pcount_3_)  &  wire673 ) | ( (~ pcount_3_)  &  pcount_2_  &  wire653 ) ;
 assign wire670 = ( pcount_3_  &  (~ wire647) ) | ( pcount_3_  &  wire7081 ) ;
 assign wire673 = ( (~ pcount_2_)  &  (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pencrypt_0_) ) ;
 assign wire682 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2374  &  n_n204 ) ;
 assign wire684 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_1_  &  (~ n_n204) ) ;
 assign wire687 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_10_  &  (~ n_n200) ) ;
 assign wire689 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_16_  &  (~ n_n204) ) ;
 assign wire692 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_20_  &  n_n204 ) ;
 assign wire693 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_47_  &  (~ n_n200) ) ;
 assign wire695 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_43_  &  (~ n_n204) ) ;
 assign wire698 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_41_  &  n_n204 ) ;
 assign wire699 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_26_  &  (~ n_n200) ) ;
 assign wire701 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_42_  &  (~ n_n204) ) ;
 assign wire704 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_25_  &  n_n204 ) ;
 assign wire705 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_45_  &  (~ n_n200) ) ;
 assign wire706 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2333  &  (~ n_n204) ) ;
 assign wire710 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_40_  &  n_n204 ) ;
 assign wire711 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_52_  &  (~ n_n200) ) ;
 assign wire714 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_57_  &  (~ n_n204) ) ;
 assign wire716 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_67_  &  n_n204 ) ;
 assign wire717 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_59_  &  (~ n_n200) ) ;
 assign wire719 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_56_  &  (~ n_n204) ) ;
 assign wire722 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_66_  &  n_n204 ) ;
 assign wire723 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_61_  &  (~ n_n200) ) ;
 assign wire725 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2374  &  (~ n_n204) ) ;
 assign wire728 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_10_  &  n_n200 ) ;
 assign wire729 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_13_  &  n_n204 ) ;
 assign wire730 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2365  &  (~ n_n204) ) ;
 assign wire734 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_16_  &  n_n204 ) ;
 assign wire735 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_28_  &  (~ n_n200) ) ;
 assign wire736 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2352  &  n_n204 ) ;
 assign wire738 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_41_  &  (~ n_n204) ) ;
 assign wire741 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_38_  &  (~ n_n200) ) ;
 assign wire744 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_32_  &  (~ n_n204) ) ;
 assign wire746 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_42_  &  n_n204 ) ;
 assign wire747 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_37_  &  (~ n_n200) ) ;
 assign wire749 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_40_  &  (~ n_n204) ) ;
 assign wire752 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_44_  &  n_n204 ) ;
 assign wire753 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_71_  &  (~ n_n200) ) ;
 assign wire756 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_53_  &  (~ n_n204) ) ;
 assign wire758 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_65_  &  n_n200 ) ;
 assign wire759 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_57_  &  n_n204 ) ;
 assign wire761 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_66_  &  (~ n_n204) ) ;
 assign wire764 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_49_  &  n_n204 ) ;
 assign wire765 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_69_  &  (~ n_n200) ) ;
 assign wire768 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_13_  &  (~ n_n204) ) ;
 assign wire770 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_21_  &  n_n204 ) ;
 assign wire771 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_12_  &  (~ n_n200) ) ;
 assign wire772 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2365  &  n_n204 ) ;
 assign wire774 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_3_  &  (~ n_n204) ) ;
 assign wire777 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_7_  &  (~ n_n200) ) ;
 assign wire780 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_29_  &  (~ n_n204) ) ;
 assign wire782 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_41_  &  n_n200 ) ;
 assign wire783 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_33_  &  n_n204 ) ;
 assign wire784 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2342  &  (~ n_n204) ) ;
 assign wire788 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_34_  &  n_n200 ) ;
 assign wire789 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_37_  &  n_n204 ) ;
 assign wire791 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_44_  &  (~ n_n204) ) ;
 assign wire794 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_31_  &  n_n204 ) ;
 assign wire795 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_54_  &  (~ n_n200) ) ;
 assign wire797 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_64_  &  (~ n_n204) ) ;
 assign wire800 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_68_  &  n_n204 ) ;
 assign wire801 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_95_  &  (~ n_n200) ) ;
 assign wire803 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_91_  &  (~ n_n204) ) ;
 assign wire806 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_89_  &  n_n204 ) ;
 assign wire807 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_74_  &  (~ n_n200) ) ;
 assign wire809 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_21_  &  (~ n_n204) ) ;
 assign wire812 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_10_  &  n_n204 ) ;
 assign wire813 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_3_  &  (~ n_n200) ) ;
 assign wire815 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_12_  &  (~ n_n204) ) ;
 assign wire818 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_3_  &  n_n204 ) ;
 assign wire819 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_20_  &  (~ n_n200) ) ;
 assign wire822 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_33_  &  (~ n_n204) ) ;
 assign wire824 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_43_  &  n_n204 ) ;
 assign wire825 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_35_  &  (~ n_n200) ) ;
 assign wire826 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2342  &  n_n204 ) ;
 assign wire828 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_25_  &  (~ n_n204) ) ;
 assign wire831 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_34_  &  (~ n_n200) ) ;
 assign wire833 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_31_  &  (~ n_n204) ) ;
 assign wire836 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_52_  &  n_n204 ) ;
 assign wire837 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_63_  &  (~ n_n200) ) ;
 assign wire839 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2301  &  (~ n_n204) ) ;
 assign wire842 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_64_  &  n_n204 ) ;
 assign wire843 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_76_  &  (~ n_n200) ) ;
 assign wire845 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_89_  &  (~ n_n204) ) ;
 assign wire848 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2288  &  n_n204 ) ;
 assign wire849 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_86_  &  (~ n_n200) ) ;
 assign wire850 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2369  &  (~ n_n204) ) ;
 assign wire854 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_12_  &  n_n204 ) ;
 assign wire855 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_16_  &  (~ n_n200) ) ;
 assign wire857 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_30_  &  (~ n_n204) ) ;
 assign wire860 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_39_  &  n_n204 ) ;
 assign wire861 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_43_  &  (~ n_n200) ) ;
 assign wire863 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_59_  &  (~ n_n204) ) ;
 assign wire866 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_50_  &  n_n204 ) ;
 assign wire867 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_48_  &  (~ n_n200) ) ;
 assign wire869 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_61_  &  (~ n_n204) ) ;
 assign wire872 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_69_  &  n_n204 ) ;
 assign wire873 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_60_  &  (~ n_n200) ) ;
 assign wire875 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_55_  &  (~ n_n204) ) ;
 assign wire878 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_76_  &  n_n204 ) ;
 assign wire879 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_87_  &  (~ n_n200) ) ;
 assign wire881 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2288  &  (~ n_n204) ) ;
 assign wire884 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_83_  &  n_n204 ) ;
 assign wire885 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_94_  &  (~ n_n200) ) ;
 assign wire886 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2369  &  n_n204 ) ;
 assign wire889 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_10_  &  (~ n_n204) ) ;
 assign wire891 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_3_  &  n_n200 ) ;
 assign wire893 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_39_  &  (~ n_n204) ) ;
 assign wire896 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_29_  &  n_n204 ) ;
 assign wire897 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_41_  &  (~ n_n200) ) ;
 assign wire898 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2320  &  (~ n_n204) ) ;
 assign wire902 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_59_  &  n_n204 ) ;
 assign wire903 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_70_  &  (~ n_n200) ) ;
 assign wire905 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_69_  &  (~ n_n204) ) ;
 assign wire908 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_58_  &  n_n204 ) ;
 assign wire909 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_51_  &  (~ n_n200) ) ;
 assign wire911 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_68_  &  (~ n_n204) ) ;
 assign wire914 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_55_  &  n_n204 ) ;
 assign wire915 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_78_  &  (~ n_n200) ) ;
 assign wire917 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_83_  &  (~ n_n204) ) ;
 assign wire920 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_74_  &  n_n204 ) ;
 assign wire921 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_72_  &  (~ n_n200) ) ;
 assign wire924 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_24_  &  (~ n_n204) ) ;
 assign wire926 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_25_  &  n_n200 ) ;
 assign wire927 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_32_  &  n_n204 ) ;
 assign wire929 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_36_  &  (~ n_n204) ) ;
 assign wire932 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_27_  &  n_n204 ) ;
 assign wire933 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_44_  &  (~ n_n200) ) ;
 assign wire934 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2320  &  n_n204 ) ;
 assign wire936 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_65_  &  (~ n_n204) ) ;
 assign wire939 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_62_  &  (~ n_n200) ) ;
 assign wire941 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_49_  &  (~ n_n204) ) ;
 assign wire944 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2310  &  n_n204 ) ;
 assign wire945 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_58_  &  (~ n_n200) ) ;
 assign wire947 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_95_  &  (~ n_n204) ) ;
 assign wire950 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_78_  &  n_n204 ) ;
 assign wire951 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_81_  &  (~ n_n200) ) ;
 assign wire953 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_74_  &  (~ n_n204) ) ;
 assign wire956 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_86_  &  n_n204 ) ;
 assign wire957 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_80_  &  (~ n_n200) ) ;
 assign wire959 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_46_  &  (~ n_n204) ) ;
 assign wire962 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_24_  &  n_n204 ) ;
 assign wire963 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_25_  &  (~ n_n200) ) ;
 assign wire964 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2333  &  n_n204 ) ;
 assign wire966 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_27_  &  (~ n_n204) ) ;
 assign wire969 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_31_  &  (~ n_n200) ) ;
 assign wire971 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_67_  &  (~ n_n204) ) ;
 assign wire974 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_65_  &  n_n204 ) ;
 assign wire975 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_50_  &  (~ n_n200) ) ;
 assign wire977 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2310  &  (~ n_n204) ) ;
 assign wire980 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2305  &  (~ n_n200) ) ;
 assign wire981 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_61_  &  n_n204 ) ;
 assign wire983 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_76_  &  (~ n_n204) ) ;
 assign wire986 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_95_  &  n_n204 ) ;
 assign wire987 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_77_  &  (~ n_n200) ) ;
 assign wire989 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_86_  &  (~ n_n204) ) ;
 assign wire992 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2280  &  (~ n_n200) ) ;
 assign wire993 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_94_  &  n_n204 ) ;
 assign wire995 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_48_  &  (~ n_n204) ) ;
 assign wire998 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_56_  &  n_n204 ) ;
 assign wire999 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2310  &  (~ n_n200) ) ;
 assign wire1001 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_60_  &  (~ n_n204) ) ;
 assign wire1004 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_51_  &  n_n204 ) ;
 assign wire1005 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_68_  &  (~ n_n200) ) ;
 assign wire1007 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_87_  &  (~ n_n204) ) ;
 assign wire1010 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_77_  &  n_n204 ) ;
 assign wire1011 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_89_  &  (~ n_n200) ) ;
 assign wire1013 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_94_  &  (~ n_n204) ) ;
 assign wire1016 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_72_  &  n_n204 ) ;
 assign wire1017 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_73_  &  (~ n_n200) ) ;
 assign wire1019 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_70_  &  (~ n_n204) ) ;
 assign wire1022 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_48_  &  n_n204 ) ;
 assign wire1023 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_49_  &  (~ n_n200) ) ;
 assign wire1025 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_51_  &  (~ n_n204) ) ;
 assign wire1028 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2301  &  n_n204 ) ;
 assign wire1029 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_55_  &  (~ n_n200) ) ;
 assign wire1031 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_78_  &  (~ n_n204) ) ;
 assign wire1034 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_87_  &  n_n204 ) ;
 assign wire1035 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_91_  &  (~ n_n200) ) ;
 assign wire1038 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_72_  &  (~ n_n204) ) ;
 assign wire1040 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_73_  &  n_n200 ) ;
 assign wire1041 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_80_  &  n_n204 ) ;
 assign wire1043 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_2_  &  (~ n_n204) ) ;
 assign wire1046 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_14_  &  n_n204 ) ;
 assign wire1047 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_8_  &  (~ n_n200) ) ;
 assign wire1049 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_62_  &  (~ n_n204) ) ;
 assign wire1052 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_70_  &  n_n204 ) ;
 assign wire1053 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_66_  &  (~ n_n200) ) ;
 assign wire1055 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_58_  &  (~ n_n204) ) ;
 assign wire1058 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2305  &  n_n204 ) ;
 assign wire1059 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2301  &  (~ n_n200) ) ;
 assign wire1061 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_81_  &  (~ n_n204) ) ;
 assign wire1064 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_91_  &  n_n204 ) ;
 assign wire1065 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_83_  &  (~ n_n200) ) ;
 assign wire1068 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_80_  &  (~ n_n204) ) ;
 assign wire1070 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2280  &  n_n204 ) ;
 assign wire1071 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_85_  &  (~ n_n200) ) ;
 assign wire1073 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_14_  &  (~ n_n204) ) ;
 assign wire1076 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_22_  &  n_n204 ) ;
 assign wire1077 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_18_  &  (~ n_n200) ) ;
 assign wire1079 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_50_  &  (~ n_n204) ) ;
 assign wire1082 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_62_  &  n_n204 ) ;
 assign wire1083 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_56_  &  (~ n_n200) ) ;
 assign wire1085 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2305  &  (~ n_n204) ) ;
 assign wire1088 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_60_  &  n_n204 ) ;
 assign wire1089 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_64_  &  (~ n_n200) ) ;
 assign wire1091 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_77_  &  (~ n_n204) ) ;
 assign wire1094 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_81_  &  n_n204 ) ;
 assign wire1095 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2288  &  (~ n_n200) ) ;
 assign wire1097 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2280  &  (~ n_n204) ) ;
 assign wire1100 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_73_  &  n_n204 ) ;
 assign wire1101 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_93_  &  (~ n_n200) ) ;
 assign wire1103 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_22_  &  (~ n_n204) ) ;
 assign wire1106 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_0_  &  n_n204 ) ;
 assign wire1107 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_1_  &  (~ n_n200) ) ;
 assign wire1109 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_47_  &  (~ n_n204) ) ;
 assign wire1112 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_30_  &  n_n204 ) ;
 assign wire1113 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_33_  &  (~ n_n200) ) ;
 assign wire1115 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_26_  &  (~ n_n204) ) ;
 assign wire1118 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_38_  &  n_n204 ) ;
 assign wire1119 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_32_  &  (~ n_n200) ) ;
 assign wire1121 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_45_  &  (~ n_n204) ) ;
 assign wire1124 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_34_  &  n_n204 ) ;
 assign wire1125 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_27_  &  (~ n_n200) ) ;
 assign wire1127 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_52_  &  (~ n_n204) ) ;
 assign wire1130 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_71_  &  n_n204 ) ;
 assign wire1131 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_53_  &  (~ n_n200) ) ;
 assign wire1133 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n10  &  (~ n_n204) ) ;
 assign wire1136 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_92_  &  n_n204 ) ;
 assign wire1137 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_23_  &  (~ n_n200) ) ;
 assign wire1140 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_0_  &  (~ n_n204) ) ;
 assign wire1142 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_1_  &  n_n200 ) ;
 assign wire1143 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_8_  &  n_n204 ) ;
 assign wire1145 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_28_  &  (~ n_n204) ) ;
 assign wire1148 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_47_  &  n_n204 ) ;
 assign wire1149 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_29_  &  (~ n_n200) ) ;
 assign wire1151 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_38_  &  (~ n_n204) ) ;
 assign wire1154 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_46_  &  n_n204 ) ;
 assign wire1155 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_42_  &  (~ n_n200) ) ;
 assign wire1158 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_37_  &  (~ n_n204) ) ;
 assign wire1160 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_45_  &  n_n204 ) ;
 assign wire1161 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_36_  &  (~ n_n200) ) ;
 assign wire1163 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_71_  &  (~ n_n204) ) ;
 assign wire1166 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_54_  &  n_n204 ) ;
 assign wire1167 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_57_  &  (~ n_n200) ) ;
 assign wire1170 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_8_  &  (~ n_n204) ) ;
 assign wire1172 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_18_  &  n_n204 ) ;
 assign wire1173 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_13_  &  (~ n_n200) ) ;
 assign wire1175 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_7_  &  (~ n_n204) ) ;
 assign wire1178 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_28_  &  n_n204 ) ;
 assign wire1179 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_39_  &  (~ n_n200) ) ;
 assign wire1180 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2352  &  (~ n_n204) ) ;
 assign wire1184 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_35_  &  n_n204 ) ;
 assign wire1185 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_46_  &  (~ n_n200) ) ;
 assign wire1187 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2337  &  (~ n_n204) ) ;
 assign wire1190 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_36_  &  n_n204 ) ;
 assign wire1191 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_40_  &  (~ n_n200) ) ;
 assign wire1193 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_54_  &  (~ n_n204) ) ;
 assign wire1196 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_63_  &  n_n204 ) ;
 assign wire1197 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_67_  &  (~ n_n200) ) ;
 assign wire1199 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_18_  &  (~ n_n204) ) ;
 assign wire1202 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_1_  &  n_n204 ) ;
 assign wire1203 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_21_  &  (~ n_n200) ) ;
 assign wire1205 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_20_  &  (~ n_n204) ) ;
 assign wire1208 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_7_  &  n_n204 ) ;
 assign wire1209 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_30_  &  (~ n_n200) ) ;
 assign wire1211 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_35_  &  (~ n_n204) ) ;
 assign wire1214 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_26_  &  n_n204 ) ;
 assign wire1215 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_24_  &  (~ n_n200) ) ;
 assign wire1217 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2337  &  n_n204 ) ;
 assign wire1219 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_34_  &  (~ n_n204) ) ;
 assign wire1221 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_27_  &  n_n200 ) ;
 assign wire1223 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_63_  &  (~ n_n204) ) ;
 assign wire1226 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_53_  &  n_n204 ) ;
 assign wire1227 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_65_  &  (~ n_n200) ) ;
 assign wire1229 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_98_  &  (~ n_n204) ) ;
 assign wire1232 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_112_  &  n_n200 ) ;
 assign wire1233 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_119_  &  n_n204 ) ;
 assign wire1235 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_126_  &  (~ n_n204) ) ;
 assign wire1238 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_122_  &  n_n204 ) ;
 assign wire1239 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_136_  &  (~ n_n200) ) ;
 assign wire1242 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_134_  &  (~ n_n204) ) ;
 assign wire1243 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2476  &  n_n200 ) ;
 assign wire1245 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_127_  &  n_n204 ) ;
 assign wire1247 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_131_  &  (~ n_n204) ) ;
 assign wire1250 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_133_  &  n_n204 ) ;
 assign wire1251 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_121_  &  (~ n_n200) ) ;
 assign wire1253 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_166_  &  (~ n_n204) ) ;
 assign wire1256 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_150_  &  n_n204 ) ;
 assign wire1257 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_154_  &  (~ n_n200) ) ;
 assign wire1259 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2448  &  (~ n_n204) ) ;
 assign wire1262 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_158_  &  n_n204 ) ;
 assign wire1263 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_163_  &  (~ n_n200) ) ;
 assign wire1265 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_148_  &  (~ n_n204) ) ;
 assign wire1268 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_155_  &  n_n204 ) ;
 assign wire1269 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_152_  &  (~ n_n200) ) ;
 assign wire1271 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_159_  &  (~ n_n204) ) ;
 assign wire1274 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_190_  &  n_n204 ) ;
 assign wire1275 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n121  &  (~ n_n200) ) ;
 assign wire1277 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_171_  &  (~ n_n204) ) ;
 assign wire1280 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2416  &  n_n204 ) ;
 assign wire1281 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2412  &  (~ n_n200) ) ;
 assign wire1284 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2272  &  (~ n_n204) ) ;
 assign wire1286 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_84_  &  n_n204 ) ;
 assign wire1287 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n10  &  (~ n_n200) ) ;
 assign wire1289 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_96_  &  (~ n_n204) ) ;
 assign wire1292 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_115_  &  n_n204 ) ;
 assign wire1293 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_105_  &  (~ n_n200) ) ;
 assign wire1295 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_142_  &  (~ n_n204) ) ;
 assign wire1298 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_126_  &  n_n204 ) ;
 assign wire1299 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_130_  &  (~ n_n200) ) ;
 assign wire1302 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_127_  &  (~ n_n204) ) ;
 assign wire1304 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_120_  &  n_n204 ) ;
 assign wire1305 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_132_  &  (~ n_n200) ) ;
 assign wire1307 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_124_  &  (~ n_n204) ) ;
 assign wire1310 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_131_  &  n_n204 ) ;
 assign wire1311 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_128_  &  (~ n_n200) ) ;
 assign wire1313 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_150_  &  (~ n_n204) ) ;
 assign wire1316 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_146_  &  n_n204 ) ;
 assign wire1317 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_160_  &  (~ n_n200) ) ;
 assign wire1319 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_147_  &  (~ n_n204) ) ;
 assign wire1322 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2448  &  n_n204 ) ;
 assign wire1323 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_144_  &  (~ n_n200) ) ;
 assign wire1325 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_155_  &  (~ n_n204) ) ;
 assign wire1328 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_157_  &  n_n204 ) ;
 assign wire1329 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_145_  &  (~ n_n200) ) ;
 assign wire1331 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_149_  &  (~ n_n204) ) ;
 assign wire1334 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_159_  &  n_n204 ) ;
 assign wire1335 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_170_  &  (~ n_n200) ) ;
 assign wire1337 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2416  &  (~ n_n204) ) ;
 assign wire1340 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_182_  &  n_n204 ) ;
 assign wire1341 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2410  &  (~ n_n200) ) ;
 assign wire1343 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_84_  &  (~ n_n204) ) ;
 assign wire1346 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_75_  &  n_n204 ) ;
 assign wire1347 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_92_  &  (~ n_n200) ) ;
 assign wire1349 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_106_  &  (~ n_n204) ) ;
 assign wire1352 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_112_  &  n_n204 ) ;
 assign wire1353 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_99_  &  (~ n_n200) ) ;
 assign wire1355 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_115_  &  (~ n_n204) ) ;
 assign wire1357 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2507  &  n_n204 ) ;
 assign wire1359 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_114_  &  (~ n_n200) ) ;
 assign wire1361 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n168  &  (~ n_n204) ) ;
 assign wire1364 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_130_  &  n_n204 ) ;
 assign wire1365 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_141_  &  (~ n_n200) ) ;
 assign wire1367 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_120_  &  (~ n_n204) ) ;
 assign wire1368 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2476  &  n_n204 ) ;
 assign wire1371 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_129_  &  (~ n_n200) ) ;
 assign wire1373 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_138_  &  (~ n_n204) ) ;
 assign wire1376 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_124_  &  n_n204 ) ;
 assign wire1377 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_140_  &  (~ n_n200) ) ;
 assign wire1379 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_125_  &  (~ n_n204) ) ;
 assign wire1382 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_135_  &  n_n204 ) ;
 assign wire1383 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_146_  &  (~ n_n200) ) ;
 assign wire1385 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_151_  &  (~ n_n204) ) ;
 assign wire1388 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_144_  &  n_n204 ) ;
 assign wire1389 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_156_  &  (~ n_n200) ) ;
 assign wire1391 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_157_  &  (~ n_n204) ) ;
 assign wire1394 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_164_  &  n_n204 ) ;
 assign wire1395 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_161_  &  (~ n_n200) ) ;
 assign wire1397 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_179_  &  (~ n_n204) ) ;
 assign wire1400 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n109  &  n_n204 ) ;
 assign wire1401 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_169_  &  (~ n_n200) ) ;
 assign wire1403 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_4_  &  (~ n_n204) ) ;
 assign wire1406 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_23_  &  n_n204 ) ;
 assign wire1407 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_5_  &  (~ n_n200) ) ;
 assign wire1408 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2268  &  n_n204 ) ;
 assign wire1410 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_75_  &  (~ n_n204) ) ;
 assign wire1413 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_79_  &  (~ n_n200) ) ;
 assign wire1415 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_119_  &  (~ n_n204) ) ;
 assign wire1418 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_106_  &  n_n204 ) ;
 assign wire1419 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_117_  &  (~ n_n200) ) ;
 assign wire1421 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2507  &  (~ n_n204) ) ;
 assign wire1424 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_108_  &  n_n204 ) ;
 assign wire1425 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_100_  &  (~ n_n200) ) ;
 assign wire1427 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_122_  &  (~ n_n204) ) ;
 assign wire1430 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2485  &  (~ n_n200) ) ;
 assign wire1431 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n168  &  n_n204 ) ;
 assign wire1432 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2474  &  n_n204 ) ;
 assign wire1434 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2476  &  (~ n_n204) ) ;
 assign wire1437 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_138_  &  (~ n_n200) ) ;
 assign wire1439 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_129_  &  (~ n_n204) ) ;
 assign wire1442 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_138_  &  n_n204 ) ;
 assign wire1443 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_133_  &  (~ n_n200) ) ;
 assign wire1445 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_135_  &  (~ n_n204) ) ;
 assign wire1448 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_166_  &  n_n204 ) ;
 assign wire1449 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_167_  &  (~ n_n200) ) ;
 assign wire1451 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_158_  &  (~ n_n204) ) ;
 assign wire1454 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_151_  &  n_n204 ) ;
 assign wire1455 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_153_  &  (~ n_n200) ) ;
 assign wire1457 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_164_  &  (~ n_n204) ) ;
 assign wire1460 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_161_  &  n_n200 ) ;
 assign wire1461 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_152_  &  n_n204 ) ;
 assign wire1463 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_172_  &  (~ n_n204) ) ;
 assign wire1466 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_179_  &  n_n204 ) ;
 assign wire1467 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_176_  &  (~ n_n200) ) ;
 assign wire1469 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_23_  &  (~ n_n204) ) ;
 assign wire1472 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_6_  &  n_n204 ) ;
 assign wire1473 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_9_  &  (~ n_n200) ) ;
 assign wire1474 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2268  &  (~ n_n204) ) ;
 assign wire1478 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n10  &  n_n204 ) ;
 assign wire1479 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_4_  &  (~ n_n200) ) ;
 assign wire1481 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2495  &  (~ n_n204) ) ;
 assign wire1484 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_101_  &  n_n204 ) ;
 assign wire1485 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_126_  &  (~ n_n200) ) ;
 assign wire1487 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2485  &  (~ n_n204) ) ;
 assign wire1490 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_141_  &  n_n204 ) ;
 assign wire1491 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_134_  &  (~ n_n200) ) ;
 assign wire1493 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_121_  &  (~ n_n204) ) ;
 assign wire1496 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_137_  &  n_n204 ) ;
 assign wire1497 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_135_  &  (~ n_n200) ) ;
 assign wire1499 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_154_  &  (~ n_n204) ) ;
 assign wire1502 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_160_  &  n_n204 ) ;
 assign wire1503 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_147_  &  (~ n_n200) ) ;
 assign wire1505 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_163_  &  (~ n_n204) ) ;
 assign wire1508 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_153_  &  n_n204 ) ;
 assign wire1509 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_162_  &  (~ n_n200) ) ;
 assign wire1511 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_152_  &  (~ n_n204) ) ;
 assign wire1514 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_145_  &  n_n204 ) ;
 assign wire1515 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_149_  &  (~ n_n200) ) ;
 assign wire1516 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2277  &  (~ n_n204) ) ;
 assign wire1520 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2272  &  (~ n_n200) ) ;
 assign wire1521 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_85_  &  n_n204 ) ;
 assign wire1523 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_113_  &  (~ n_n204) ) ;
 assign wire1526 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2495  &  n_n204 ) ;
 assign wire1527 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_142_  &  (~ n_n200) ) ;
 assign wire1529 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_141_  &  (~ n_n204) ) ;
 assign wire1532 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_123_  &  n_n204 ) ;
 assign wire1533 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_127_  &  (~ n_n200) ) ;
 assign wire1536 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_128_  &  (~ n_n204) ) ;
 assign wire1538 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_121_  &  n_n204 ) ;
 assign wire1539 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_125_  &  (~ n_n200) ) ;
 assign wire1541 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2452  &  n_n204 ) ;
 assign wire1542 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_160_  &  (~ n_n204) ) ;
 assign wire1545 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2448  &  (~ n_n200) ) ;
 assign wire1547 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_144_  &  (~ n_n204) ) ;
 assign wire1550 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2440  &  (~ n_n200) ) ;
 assign wire1551 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_163_  &  n_n204 ) ;
 assign wire1553 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_145_  &  (~ n_n204) ) ;
 assign wire1556 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_161_  &  n_n204 ) ;
 assign wire1557 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_159_  &  (~ n_n200) ) ;
 assign wire1559 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_85_  &  (~ n_n204) ) ;
 assign wire1562 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_93_  &  n_n204 ) ;
 assign wire1563 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_84_  &  (~ n_n200) ) ;
 assign wire1565 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_111_  &  (~ n_n204) ) ;
 assign wire1568 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_142_  &  n_n204 ) ;
 assign wire1569 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n168  &  (~ n_n200) ) ;
 assign wire1571 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_123_  &  (~ n_n204) ) ;
 assign wire1572 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2481  &  n_n204 ) ;
 assign wire1575 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_120_  &  (~ n_n200) ) ;
 assign wire1578 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_140_  &  (~ n_n204) ) ;
 assign wire1580 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_137_  &  n_n200 ) ;
 assign wire1581 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_128_  &  n_n204 ) ;
 assign wire1584 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_146_  &  (~ n_n204) ) ;
 assign wire1586 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_160_  &  n_n200 ) ;
 assign wire1587 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_167_  &  n_n204 ) ;
 assign wire1589 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_156_  &  (~ n_n204) ) ;
 assign wire1592 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2440  &  n_n204 ) ;
 assign wire1593 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_155_  &  (~ n_n200) ) ;
 assign wire1595 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_161_  &  (~ n_n204) ) ;
 assign wire1596 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2430  &  n_n204 ) ;
 assign wire1599 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_190_  &  (~ n_n200) ) ;
 assign wire1601 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_93_  &  (~ n_n204) ) ;
 assign wire1604 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_82_  &  n_n204 ) ;
 assign wire1605 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_75_  &  (~ n_n200) ) ;
 assign wire1607 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_101_  &  (~ n_n204) ) ;
 assign wire1610 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_111_  &  n_n204 ) ;
 assign wire1611 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_122_  &  (~ n_n200) ) ;
 assign wire1613 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2481  &  (~ n_n204) ) ;
 assign wire1616 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_120_  &  n_n200 ) ;
 assign wire1617 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_134_  &  n_n204 ) ;
 assign wire1619 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_133_  &  (~ n_n204) ) ;
 assign wire1622 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_140_  &  n_n204 ) ;
 assign wire1623 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_137_  &  (~ n_n200) ) ;
 assign wire1626 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_167_  &  (~ n_n204) ) ;
 assign wire1628 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_154_  &  n_n204 ) ;
 assign wire1629 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_165_  &  (~ n_n200) ) ;
 assign wire1631 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_153_  &  (~ n_n204) ) ;
 assign wire1634 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_156_  &  n_n204 ) ;
 assign wire1635 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_148_  &  (~ n_n200) ) ;
 assign wire1637 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2430  &  (~ n_n204) ) ;
 assign wire1640 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_149_  &  n_n204 ) ;
 assign wire1641 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_174_  &  (~ n_n200) ) ;
 assign wire1644 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_82_  &  (~ n_n204) ) ;
 assign wire1646 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_75_  &  n_n200 ) ;
 assign wire1647 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2272  &  n_n204 ) ;
 assign wire1649 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_102_  &  (~ n_n204) ) ;
 assign wire1652 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_98_  &  n_n204 ) ;
 assign wire1653 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_112_  &  (~ n_n200) ) ;
 assign wire1655 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_110_  &  (~ n_n204) ) ;
 assign wire1658 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_115_  &  n_n200 ) ;
 assign wire1659 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_103_  &  n_n204 ) ;
 assign wire1661 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_107_  &  (~ n_n204) ) ;
 assign wire1664 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_109_  &  n_n204 ) ;
 assign wire1665 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_97_  &  (~ n_n200) ) ;
 assign wire1667 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_189_  &  (~ n_n204) ) ;
 assign wire1670 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_171_  &  n_n204 ) ;
 assign wire1671 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_175_  &  (~ n_n200) ) ;
 assign wire1673 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_177_  &  (~ n_n204) ) ;
 assign wire1676 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_186_  &  n_n204 ) ;
 assign wire1677 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n109  &  (~ n_n200) ) ;
 assign wire1679 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2396  &  (~ n_n204) ) ;
 assign wire1682 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_173_  &  n_n204 ) ;
 assign wire1683 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_102_  &  (~ n_n200) ) ;
 assign wire1685 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_19_  &  (~ n_n204) ) ;
 assign wire1688 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_17_  &  n_n204 ) ;
 assign wire1689 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_2_  &  (~ n_n200) ) ;
 assign wire1691 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2513  &  (~ n_n204) ) ;
 assign wire1694 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_110_  &  n_n204 ) ;
 assign wire1695 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_115_  &  (~ n_n200) ) ;
 assign wire1697 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_109_  &  (~ n_n204) ) ;
 assign wire1700 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_116_  &  n_n204 ) ;
 assign wire1701 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_113_  &  (~ n_n200) ) ;
 assign wire1703 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2420  &  (~ n_n204) ) ;
 assign wire1706 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_189_  &  n_n204 ) ;
 assign wire1707 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_182_  &  (~ n_n200) ) ;
 assign wire1709 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_186_  &  (~ n_n204) ) ;
 assign wire1712 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_172_  &  n_n204 ) ;
 assign wire1713 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_188_  &  (~ n_n200) ) ;
 assign wire1715 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_185_  &  (~ n_n204) ) ;
 assign wire1718 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2396  &  n_n204 ) ;
 assign wire1719 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_118_  &  (~ n_n200) ) ;
 assign wire1721 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_17_  &  (~ n_n204) ) ;
 assign wire1724 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2384  &  n_n204 ) ;
 assign wire1725 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_14_  &  (~ n_n200) ) ;
 assign wire1727 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_183_  &  (~ n_n204) ) ;
 assign wire1730 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_118_  &  n_n204 ) ;
 assign wire1731 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_119_  &  (~ n_n200) ) ;
 assign wire1733 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_116_  &  (~ n_n204) ) ;
 assign wire1736 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2495  &  (~ n_n200) ) ;
 assign wire1737 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_104_  &  n_n204 ) ;
 assign wire1739 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_97_  &  (~ n_n204) ) ;
 assign wire1742 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_113_  &  n_n204 ) ;
 assign wire1743 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_111_  &  (~ n_n200) ) ;
 assign wire1745 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_130_  &  (~ n_n204) ) ;
 assign wire1748 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_136_  &  n_n204 ) ;
 assign wire1749 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_123_  &  (~ n_n200) ) ;
 assign wire1751 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_184_  &  (~ n_n204) ) ;
 assign wire1754 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2416  &  (~ n_n200) ) ;
 assign wire1755 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2420  &  n_n204 ) ;
 assign wire1757 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2408  &  (~ n_n204) ) ;
 assign wire1760 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_180_  &  n_n204 ) ;
 assign wire1761 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_172_  &  (~ n_n200) ) ;
 assign wire1763 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_79_  &  (~ n_n204) ) ;
 assign wire1766 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_4_  &  n_n204 ) ;
 assign wire1767 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_15_  &  (~ n_n200) ) ;
 assign wire1769 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2384  &  (~ n_n204) ) ;
 assign wire1772 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_11_  &  n_n204 ) ;
 assign wire1773 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_22_  &  (~ n_n200) ) ;
 assign wire1775 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_118_  &  (~ n_n204) ) ;
 assign wire1778 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_102_  &  n_n204 ) ;
 assign wire1779 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_106_  &  (~ n_n200) ) ;
 assign wire1781 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_103_  &  (~ n_n204) ) ;
 assign wire1784 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_96_  &  n_n204 ) ;
 assign wire1785 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_108_  &  (~ n_n200) ) ;
 assign wire1787 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_104_  &  (~ n_n204) ) ;
 assign wire1790 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_97_  &  n_n204 ) ;
 assign wire1791 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_101_  &  (~ n_n200) ) ;
 assign wire1793 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_136_  &  (~ n_n204) ) ;
 assign wire1796 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_123_  &  n_n200 ) ;
 assign wire1797 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2485  &  n_n204 ) ;
 assign wire1799 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_178_  &  (~ n_n204) ) ;
 assign wire1802 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_184_  &  n_n204 ) ;
 assign wire1803 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_171_  &  (~ n_n200) ) ;
 assign wire1805 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_180_  &  (~ n_n204) ) ;
 assign wire1808 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_177_  &  n_n204 ) ;
 assign wire1809 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_179_  &  (~ n_n200) ) ;
 assign wire1811 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_92_  &  (~ n_n204) ) ;
 assign wire1814 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_79_  &  n_n204 ) ;
 assign wire1815 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_6_  &  (~ n_n200) ) ;
 assign wire1817 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_11_  &  (~ n_n204) ) ;
 assign wire1820 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_2_  &  n_n204 ) ;
 assign wire1821 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_0_  &  (~ n_n200) ) ;
 assign wire1822 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2277  &  n_n204 ) ;
 assign wire1824 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_73_  &  (~ n_n204) ) ;
 assign wire1827 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_82_  &  (~ n_n200) ) ;
 assign wire1829 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2517  &  (~ n_n204) ) ;
 assign wire1832 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_117_  &  n_n204 ) ;
 assign wire1833 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_110_  &  (~ n_n200) ) ;
 assign wire1835 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_108_  &  (~ n_n204) ) ;
 assign wire1838 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_105_  &  n_n204 ) ;
 assign wire1839 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_107_  &  (~ n_n200) ) ;
 assign wire1841 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_132_  &  (~ n_n204) ) ;
 assign wire1844 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_129_  &  n_n204 ) ;
 assign wire1845 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_131_  &  (~ n_n200) ) ;
 assign wire1847 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2462  &  n_n204 ) ;
 assign wire1848 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_137_  &  (~ n_n204) ) ;
 assign wire1851 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_166_  &  (~ n_n200) ) ;
 assign wire1853 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n121  &  (~ n_n204) ) ;
 assign wire1856 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_178_  &  n_n204 ) ;
 assign wire1857 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_189_  &  (~ n_n200) ) ;
 assign wire1859 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2412  &  (~ n_n204) ) ;
 assign wire1862 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2410  &  n_n204 ) ;
 assign wire1863 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_177_  &  (~ n_n200) ) ;
 assign wire1865 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_188_  &  (~ n_n204) ) ;
 assign wire1868 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_176_  &  n_n204 ) ;
 assign wire1869 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2396  &  (~ n_n200) ) ;
 assign wire1871 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_6_  &  (~ n_n204) ) ;
 assign wire1874 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_15_  &  n_n204 ) ;
 assign wire1875 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_19_  &  (~ n_n200) ) ;
 assign wire1877 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_173_  &  (~ n_n204) ) ;
 assign wire1880 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_183_  &  n_n204 ) ;
 assign wire1881 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_98_  &  (~ n_n200) ) ;
 assign wire1883 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_112_  &  (~ n_n204) ) ;
 assign wire1885 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2517  &  n_n204 ) ;
 assign wire1887 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2513  &  (~ n_n200) ) ;
 assign wire1889 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_105_  &  (~ n_n204) ) ;
 assign wire1892 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_114_  &  n_n204 ) ;
 assign wire1893 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_109_  &  (~ n_n200) ) ;
 assign wire1894 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2474  &  (~ n_n204) ) ;
 assign wire1898 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_132_  &  n_n204 ) ;
 assign wire1899 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_124_  &  (~ n_n200) ) ;
 assign wire1901 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2462  &  (~ n_n204) ) ;
 assign wire1904 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_125_  &  n_n204 ) ;
 assign wire1905 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_150_  &  (~ n_n200) ) ;
 assign wire1907 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_170_  &  (~ n_n204) ) ;
 assign wire1910 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2420  &  (~ n_n200) ) ;
 assign wire1911 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n121  &  n_n204 ) ;
 assign wire1913 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2410  &  (~ n_n204) ) ;
 assign wire1916 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2408  &  n_n204 ) ;
 assign wire1917 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_186_  &  (~ n_n200) ) ;
 assign wire1919 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n109  &  (~ n_n204) ) ;
 assign wire1922 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_188_  &  n_n204 ) ;
 assign wire1923 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_185_  &  (~ n_n200) ) ;
 assign wire1925 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_15_  &  (~ n_n204) ) ;
 assign wire1928 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_5_  &  n_n204 ) ;
 assign wire1929 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_17_  &  (~ n_n200) ) ;
 assign wire1931 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_99_  &  (~ n_n204) ) ;
 assign wire1934 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2513  &  n_n204 ) ;
 assign wire1935 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_96_  &  (~ n_n200) ) ;
 assign wire1937 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_114_  &  (~ n_n204) ) ;
 assign wire1940 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_100_  &  n_n204 ) ;
 assign wire1941 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_116_  &  (~ n_n200) ) ;
 assign wire1943 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_165_  &  (~ n_n204) ) ;
 assign wire1946 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_147_  &  n_n204 ) ;
 assign wire1947 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_151_  &  (~ n_n200) ) ;
 assign wire1949 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2440  &  (~ n_n204) ) ;
 assign wire1952 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_162_  &  n_n204 ) ;
 assign wire1953 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_157_  &  (~ n_n200) ) ;
 assign wire1955 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_174_  &  (~ n_n204) ) ;
 assign wire1958 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_170_  &  n_n204 ) ;
 assign wire1959 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_184_  &  (~ n_n200) ) ;
 assign wire1961 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_182_  &  (~ n_n204) ) ;
 assign wire1964 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2408  &  (~ n_n200) ) ;
 assign wire1965 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_175_  &  n_n204 ) ;
 assign wire1967 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_169_  &  (~ n_n204) ) ;
 assign wire1970 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_185_  &  n_n204 ) ;
 assign wire1971 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_183_  &  (~ n_n200) ) ;
 assign wire1973 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_5_  &  (~ n_n204) ) ;
 assign wire1976 = ( (~ pstart_0_)  &  pencrypt_0_  &  n_n2384  &  (~ n_n200) ) ;
 assign wire1977 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_9_  &  n_n204 ) ;
 assign wire1979 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_117_  &  (~ n_n204) ) ;
 assign wire1982 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_99_  &  n_n204 ) ;
 assign wire1983 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_103_  &  (~ n_n200) ) ;
 assign wire1985 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_100_  &  (~ n_n204) ) ;
 assign wire1988 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_107_  &  n_n204 ) ;
 assign wire1989 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_104_  &  (~ n_n200) ) ;
 assign wire1991 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2452  &  (~ n_n204) ) ;
 assign wire1994 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_165_  &  n_n204 ) ;
 assign wire1995 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_158_  &  (~ n_n200) ) ;
 assign wire1997 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_162_  &  (~ n_n204) ) ;
 assign wire2000 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_148_  &  n_n204 ) ;
 assign wire2001 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_164_  &  (~ n_n200) ) ;
 assign wire2003 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_190_  &  (~ n_n204) ) ;
 assign wire2006 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_174_  &  n_n204 ) ;
 assign wire2007 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_178_  &  (~ n_n200) ) ;
 assign wire2009 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_175_  &  (~ n_n204) ) ;
 assign wire2012 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  n_n2412  &  n_n204 ) ;
 assign wire2013 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_180_  &  (~ n_n200) ) ;
 assign wire2015 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_176_  &  (~ n_n204) ) ;
 assign wire2018 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_169_  &  n_n204 ) ;
 assign wire2019 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_173_  &  (~ n_n200) ) ;
 assign wire2021 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_9_  &  (~ n_n204) ) ;
 assign wire2024 = ( (~ pstart_0_)  &  (~ pencrypt_0_)  &  pksi_19_  &  n_n204 ) ;
 assign wire2025 = ( (~ pstart_0_)  &  pencrypt_0_  &  pksi_11_  &  (~ n_n200) ) ;
 assign wire6182 = ( pkey_57_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_0_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6183 = ( wire6182 ) | ( n_n2384  &  n_n200  &  wire655 ) ;
 assign wire6186 = ( pkey_211_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_219_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6187 = ( wire6186 ) | ( n_n2396  &  n_n200  &  wire655 ) ;
 assign wire6190 = ( pkey_213_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_205_ ) ;
 assign wire6191 = ( wire6190 ) | ( n_n2408  &  n_n200  &  wire655 ) ;
 assign wire6194 = ( pkey_230_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_238_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6195 = ( wire6194 ) | ( n_n121  &  n_n200  &  wire655 ) ;
 assign wire6198 = ( pkey_156_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_164_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6199 = ( wire6198 ) | ( pksi_157_  &  n_n200  &  wire655 ) ;
 assign wire6202 = ( pstart_0_  &  pkey_181_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_189_ ) ;
 assign wire6203 = ( wire6202 ) | ( n_n2448  &  n_n200  &  wire655 ) ;
 assign wire6206 = ( pkey_28_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_20_ ) ;
 assign wire6207 = ( wire6206 ) | ( pksi_116_  &  n_n200  &  wire655 ) ;
 assign wire6210 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_53_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_45_ ) ;
 assign wire6211 = ( wire6210 ) | ( pksi_110_  &  n_n200  &  wire655 ) ;
 assign wire6214 = ( pkey_0_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_8_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6215 = ( wire6214 ) | ( pksi_17_  &  n_n200  &  wire655 ) ;
 assign wire6218 = ( pstart_0_  &  pkey_203_  &  pencrypt_0_ ) | ( pkey_211_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6219 = ( wire6218 ) | ( pksi_173_  &  n_n200  &  wire655 ) ;
 assign wire6222 = ( pkey_213_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_221_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6223 = ( wire6222 ) | ( n_n2410  &  n_n200  &  wire655 ) ;
 assign wire6226 = ( pkey_222_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_230_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6227 = ( wire6226 ) | ( pksi_178_  &  n_n200  &  wire655 ) ;
 assign wire6230 = ( pkey_164_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_172_ ) ;
 assign wire6231 = ( wire6230 ) | ( pksi_155_  &  n_n200  &  wire655 ) ;
 assign wire6234 = ( pstart_0_  &  pkey_181_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_173_ ) ;
 assign wire6235 = ( wire6234 ) | ( pksi_158_  &  n_n200  &  wire655 ) ;
 assign wire6238 = ( pkey_28_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_36_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6239 = ( wire6238 ) | ( pksi_109_  &  n_n200  &  wire655 ) ;
 assign wire6242 = ( pkey_37_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_45_ ) ;
 assign wire6243 = ( wire6242 ) | ( pksi_103_  &  n_n200  &  wire655 ) ;
 assign wire6246 = ( pkey_8_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_16_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6247 = ( wire6246 ) | ( pksi_19_  &  n_n200  &  wire655 ) ;
 assign wire6250 = ( pstart_0_  &  pkey_196_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_204_ ) ;
 assign wire6251 = ( wire6250 ) | ( pksi_169_  &  n_n200  &  wire655 ) ;
 assign wire6254 = ( pkey_252_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_197_  &  (~ pencrypt_0_) ) ;
 assign wire6255 = ( wire6254 ) | ( pksi_177_  &  n_n200  &  wire655 ) ;
 assign wire6258 = ( pkey_214_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_222_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6259 = ( wire6258 ) | ( pksi_184_  &  n_n200  &  wire655 ) ;
 assign wire6262 = ( pkey_67_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_190_ ) ;
 assign wire6263 = ( wire6262 ) | ( pksi_166_  &  n_n200  &  wire655 ) ;
 assign wire6266 = ( pkey_116_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_124_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6267 = ( wire6266 ) | ( pksi_138_  &  n_n200  &  wire655 ) ;
 assign wire6270 = ( pkey_36_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_44_ ) ;
 assign wire6271 = ( wire6270 ) | ( pksi_107_  &  n_n200  &  wire655 ) ;
 assign wire6274 = ( pkey_61_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_6_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6275 = ( wire6274 ) | ( pksi_99_  &  n_n200  &  wire655 ) ;
 assign wire6278 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_62_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_54_ ) ;
 assign wire6279 = ( wire6278 ) | ( pksi_102_  &  n_n200  &  wire655 ) ;
 assign wire6282 = ( pkey_16_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_24_ ) ;
 assign wire6283 = ( wire6282 ) | ( pksi_9_  &  n_n200  &  wire655 ) ;
 assign wire6286 = ( pkey_219_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_196_  &  (~ pencrypt_0_) ) ;
 assign wire6287 = ( wire6286 ) | ( pksi_185_  &  n_n200  &  wire655 ) ;
 assign wire6290 = ( pstart_0_  &  pkey_197_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_205_ ) ;
 assign wire6291 = ( wire6290 ) | ( pksi_180_  &  n_n200  &  wire655 ) ;
 assign wire6294 = ( pkey_206_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_214_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6295 = ( wire6294 ) | ( n_n2420  &  n_n200  &  wire655 ) ;
 assign wire6298 = ( pkey_67_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_75_ ) ;
 assign wire6299 = ( wire6298 ) | ( pksi_135_  &  n_n200  &  wire655 ) ;
 assign wire6302 = ( pkey_116_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_44_ ) ;
 assign wire6303 = ( wire6302 ) | ( pksi_124_  &  n_n200  &  wire655 ) ;
 assign wire6306 = ( pstart_0_  &  pkey_52_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_44_ ) ;
 assign wire6307 = ( wire6306 ) | ( pksi_100_  &  n_n200  &  wire655 ) ;
 assign wire6310 = ( pkey_61_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_53_ ) ;
 assign wire6311 = ( wire6310 ) | ( n_n2513  &  n_n200  &  wire655 ) ;
 assign wire6314 = ( pkey_226_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_234_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6315 = ( wire6314 ) | ( pksi_93_  &  n_n200  &  wire655 ) ;
 assign wire6318 = ( pstart_0_  &  pencrypt_0_  &  pkey_25_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_33_ ) ;
 assign wire6319 = ( wire6318 ) | ( pksi_22_  &  n_n200  &  wire655 ) ;
 assign wire6322 = ( pkey_48_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_56_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6323 = ( wire6322 ) | ( pksi_23_  &  n_n200  &  wire655 ) ;
 assign wire6326 = ( pkey_244_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_172_ ) ;
 assign wire6327 = ( wire6326 ) | ( pksi_172_  &  n_n200  &  wire655 ) ;
 assign wire6330 = ( pkey_206_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_198_ ) ;
 assign wire6331 = ( wire6330 ) | ( pksi_189_  &  n_n200  &  wire655 ) ;
 assign wire6334 = ( pkey_125_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_70_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6335 = ( wire6334 ) | ( n_n2481  &  (~ n_n200)  &  wire655 ) ;
 assign wire6338 = ( pkey_19_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_27_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6339 = ( wire6338 ) | ( n_n2495  &  n_n200  &  wire655 ) ;
 assign wire6342 = ( pstart_0_  &  pencrypt_0_  &  pkey_13_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_21_ ) ;
 assign wire6343 = ( wire6342 ) | ( n_n2507  &  n_n200  &  wire655 ) ;
 assign wire6346 = ( pkey_38_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_46_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6347 = ( wire6346 ) | ( pksi_119_  &  n_n200  &  wire655 ) ;
 assign wire6350 = ( pstart_0_  &  pencrypt_0_  &  pkey_33_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_41_ ) ;
 assign wire6351 = ( wire6350 ) | ( pksi_14_  &  n_n200  &  wire655 ) ;
 assign wire6354 = ( pkey_48_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_40_ ) ;
 assign wire6355 = ( wire6354 ) | ( pksi_6_  &  n_n200  &  wire655 ) ;
 assign wire6358 = ( pkey_244_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_252_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6359 = ( wire6358 ) | ( pksi_186_  &  n_n200  &  wire655 ) ;
 assign wire6362 = ( pkey_253_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_198_ ) ;
 assign wire6363 = ( wire6362 ) | ( pksi_171_  &  n_n200  &  wire655 ) ;
 assign wire6366 = ( pkey_70_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_78_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6367 = ( wire6366 ) | ( pksi_141_  &  n_n200  &  wire655 ) ;
 assign wire6370 = ( pkey_19_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_11_ ) ;
 assign wire6371 = ( wire6370 ) | ( pksi_101_  &  n_n200  &  wire655 ) ;
 assign wire6374 = ( pkey_27_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_4_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6375 = ( wire6374 ) | ( pksi_113_  &  n_n200  &  wire655 ) ;
 assign wire6378 = ( pkey_46_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_54_ ) ;
 assign wire6379 = ( wire6378 ) | ( pksi_98_  &  n_n200  &  wire655 ) ;
 assign wire6382 = ( pkey_49_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_41_ ) ;
 assign wire6383 = ( wire6382 ) | ( pksi_2_  &  n_n200  &  wire655 ) ;
 assign wire6386 = ( pkey_195_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_203_  &  (~ pencrypt_0_) ) ;
 assign wire6387 = ( wire6386 ) | ( pksi_183_  &  n_n200  &  wire655 ) ;
 assign wire6390 = ( pkey_220_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_228_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6391 = ( wire6390 ) | ( n_n109  &  n_n200  &  wire655 ) ;
 assign wire6394 = ( pkey_245_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_253_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6395 = ( wire6394 ) | ( n_n2416  &  n_n200  &  wire655 ) ;
 assign wire6398 = ( pkey_4_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_12_ ) ;
 assign wire6399 = ( wire6398 ) | ( pksi_97_  &  n_n200  &  wire655 ) ;
 assign wire6402 = ( pkey_29_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_37_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6403 = ( wire6402 ) | ( pksi_96_  &  n_n200  &  wire655 ) ;
 assign wire6406 = ( pkey_49_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_57_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6407 = ( wire6406 ) | ( pksi_11_  &  n_n200  &  wire655 ) ;
 assign wire6410 = ( pkey_195_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_62_ ) ;
 assign wire6411 = ( wire6410 ) | ( pksi_118_  &  n_n200  &  wire655 ) ;
 assign wire6414 = ( pkey_228_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_172_ ) ;
 assign wire6415 = ( wire6414 ) | ( pksi_179_  &  n_n200  &  wire655 ) ;
 assign wire6418 = ( pkey_237_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_245_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6419 = ( wire6418 ) | ( pksi_182_  &  n_n200  &  wire655 ) ;
 assign wire6422 = ( pstart_0_  &  pencrypt_0_  &  pkey_12_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_20_ ) ;
 assign wire6423 = ( wire6422 ) | ( pksi_104_  &  n_n200  &  wire655 ) ;
 assign wire6426 = ( pkey_29_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_21_ ) ;
 assign wire6427 = ( wire6426 ) | ( n_n2507  &  (~ n_n200)  &  wire655 ) ;
 assign wire6430 = ( pkey_38_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_30_ ) ;
 assign wire6431 = ( wire6430 ) | ( pksi_106_  &  n_n200  &  wire655 ) ;
 assign wire6434 = ( pkey_194_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_202_ ) ;
 assign wire6435 = ( wire6434 ) | ( n_n2268  &  (~ n_n200)  &  wire655 ) ;
 assign wire6438 = ( pkey_254_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_131_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6439 = ( wire6438 ) | ( pksi_190_  &  n_n200  &  wire655 ) ;
 assign wire6442 = ( pkey_180_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_188_ ) ;
 assign wire6443 = ( wire6442 ) | ( pksi_162_  &  n_n200  &  wire655 ) ;
 assign wire6446 = ( pkey_142_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_150_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6447 = ( wire6446 ) | ( n_n2452  &  n_n200  &  wire655 ) ;
 assign wire6450 = ( pkey_68_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_76_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6451 = ( wire6450 ) | ( pksi_121_  &  n_n200  &  wire655 ) ;
 assign wire6454 = ( pkey_93_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_101_ ) ;
 assign wire6455 = ( wire6454 ) | ( n_n2476  &  (~ n_n200)  &  wire655 ) ;
 assign wire6458 = ( pkey_118_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_126_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6459 = ( wire6458 ) | ( pksi_126_  &  n_n200  &  wire655 ) ;
 assign wire6462 = ( pkey_210_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_202_ ) ;
 assign wire6463 = ( wire6462 ) | ( pksi_84_  &  n_n200  &  wire655 ) ;
 assign wire6466 = ( pkey_131_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_139_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6467 = ( wire6466 ) | ( pksi_159_  &  n_n200  &  wire655 ) ;
 assign wire6470 = ( pkey_180_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_172_ ) ;
 assign wire6471 = ( wire6470 ) | ( pksi_148_  &  n_n200  &  wire655 ) ;
 assign wire6474 = ( pkey_150_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_158_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6475 = ( wire6474 ) | ( n_n2452  &  (~ n_n200)  &  wire655 ) ;
 assign wire6478 = ( pkey_68_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_91_ ) ;
 assign wire6479 = ( wire6478 ) | ( n_n2462  &  (~ n_n200)  &  wire655 ) ;
 assign wire6482 = ( pstart_0_  &  pkey_109_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_101_ ) ;
 assign wire6483 = ( wire6482 ) | ( pksi_127_  &  n_n200  &  wire655 ) ;
 assign wire6486 = ( pkey_110_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_118_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6487 = ( wire6486 ) | ( pksi_122_  &  n_n200  &  wire655 ) ;
 assign wire6490 = ( pkey_210_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_218_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6491 = ( wire6490 ) | ( n_n2272  &  n_n200  &  wire655 ) ;
 assign wire6494 = ( pkey_139_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_147_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6495 = ( wire6494 ) | ( pksi_149_  &  n_n200  &  wire655 ) ;
 assign wire6498 = ( pkey_133_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_141_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6499 = ( wire6498 ) | ( pksi_156_  &  n_n200  &  wire655 ) ;
 assign wire6502 = ( pkey_134_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_189_ ) ;
 assign wire6503 = ( wire6502 ) | ( pksi_147_  &  n_n200  &  wire655 ) ;
 assign wire6506 = ( pstart_0_  &  pencrypt_0_  &  pkey_83_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_91_ ) ;
 assign wire6507 = ( wire6506 ) | ( n_n2462  &  n_n200  &  wire655 ) ;
 assign wire6510 = ( pstart_0_  &  pkey_109_  &  pencrypt_0_ ) | ( pkey_117_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6511 = ( wire6510 ) | ( pksi_134_  &  n_n200  &  wire655 ) ;
 assign wire6514 = ( pkey_3_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_11_ ) ;
 assign wire6515 = ( wire6514 ) | ( pksi_111_  &  n_n200  &  wire655 ) ;
 assign wire6518 = ( pkey_218_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_226_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6519 = ( wire6518 ) | ( pksi_82_  &  n_n200  &  wire655 ) ;
 assign wire6522 = ( pkey_147_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_155_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6523 = ( wire6522 ) | ( n_n2430  &  n_n200  &  wire655 ) ;
 assign wire6526 = ( pkey_133_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_188_ ) ;
 assign wire6527 = ( wire6526 ) | ( n_n2440  &  n_n200  &  wire655 ) ;
 assign wire6530 = ( pkey_134_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_142_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6531 = ( wire6530 ) | ( pksi_165_  &  n_n200  &  wire655 ) ;
 assign wire6534 = ( pstart_0_  &  pencrypt_0_  &  pkey_75_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_83_ ) ;
 assign wire6535 = ( wire6534 ) | ( pksi_125_  &  n_n200  &  wire655 ) ;
 assign wire6538 = ( pkey_117_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_125_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6539 = ( wire6538 ) | ( n_n2481  &  n_n200  &  wire655 ) ;
 assign wire6542 = ( pkey_126_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_3_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6543 = ( wire6542 ) | ( pksi_142_  &  n_n200  &  wire655 ) ;
 assign wire6546 = ( pkey_227_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_235_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6547 = ( wire6546 ) | ( pksi_79_  &  n_n200  &  wire655 ) ;
 assign wire6550 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_32_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_24_ ) ;
 assign wire6551 = ( wire6550 ) | ( pksi_5_  &  n_n200  &  wire655 ) ;
 assign wire6554 = ( pkey_212_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_220_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6555 = ( wire6554 ) | ( pksi_188_  &  n_n200  &  wire655 ) ;
 assign wire6558 = ( pkey_155_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_132_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6559 = ( wire6558 ) | ( n_n2430  &  (~ n_n200)  &  wire655 ) ;
 assign wire6562 = ( pkey_149_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_157_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6563 = ( wire6562 ) | ( pksi_163_  &  n_n200  &  wire655 ) ;
 assign wire6566 = ( pkey_182_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_174_ ) ;
 assign wire6567 = ( wire6566 ) | ( pksi_146_  &  n_n200  &  wire655 ) ;
 assign wire6570 = ( pstart_0_  &  pencrypt_0_  &  pkey_100_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_44_ ) ;
 assign wire6571 = ( wire6570 ) | ( pksi_131_  &  n_n200  &  wire655 ) ;
 assign wire6574 = ( pkey_124_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_69_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6575 = ( wire6574 ) | ( pksi_129_  &  n_n200  &  wire655 ) ;
 assign wire6578 = ( pkey_86_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_94_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6579 = ( wire6578 ) | ( pksi_136_  &  n_n200  &  wire655 ) ;
 assign wire6582 = ( pstart_0_  &  pkey_52_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_60_  &  (~ pencrypt_0_) ) ;
 assign wire6583 = ( wire6582 ) | ( pksi_114_  &  n_n200  &  wire655 ) ;
 assign wire6586 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_22_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_14_ ) ;
 assign wire6587 = ( wire6586 ) | ( n_n2517  &  n_n200  &  wire655 ) ;
 assign wire6590 = ( pkey_235_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_243_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6591 = ( wire6590 ) | ( pksi_92_  &  n_n200  &  wire655 ) ;
 assign wire6594 = ( pstart_0_  &  pencrypt_0_  &  pkey_32_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_40_ ) ;
 assign wire6595 = ( wire6594 ) | ( pksi_15_  &  n_n200  &  wire655 ) ;
 assign wire6598 = ( pkey_212_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_204_ ) ;
 assign wire6599 = ( wire6598 ) | ( pksi_176_  &  n_n200  &  wire655 ) ;
 assign wire6602 = ( pkey_132_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_140_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6603 = ( wire6602 ) | ( pksi_145_  &  n_n200  &  wire655 ) ;
 assign wire6606 = ( pkey_141_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_149_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6607 = ( wire6606 ) | ( pksi_153_  &  n_n200  &  wire655 ) ;
 assign wire6610 = ( pkey_182_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_190_ ) ;
 assign wire6611 = ( wire6610 ) | ( pksi_150_  &  n_n200  &  wire655 ) ;
 assign wire6614 = ( pkey_92_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_100_ ) ;
 assign wire6615 = ( wire6614 ) | ( pksi_133_  &  n_n200  &  wire655 ) ;
 assign wire6618 = ( pkey_69_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_77_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6619 = ( wire6618 ) | ( pksi_132_  &  n_n200  &  wire655 ) ;
 assign wire6622 = ( pkey_78_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_86_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6623 = ( wire6622 ) | ( n_n2485  &  n_n200  &  wire655 ) ;
 assign wire6626 = ( pstart_0_  &  pkey_60_  &  pencrypt_0_ ) | ( pkey_5_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6627 = ( wire6626 ) | ( pksi_105_  &  n_n200  &  wire655 ) ;
 assign wire6630 = ( pkey_6_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_14_ ) ;
 assign wire6631 = ( wire6630 ) | ( pksi_117_  &  n_n200  &  wire655 ) ;
 assign wire6634 = ( pkey_243_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_251_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6635 = ( wire6634 ) | ( n_n10  &  n_n200  &  wire655 ) ;
 assign wire6638 = ( pkey_221_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_229_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6639 = ( wire6638 ) | ( n_n2412  &  n_n200  &  wire655 ) ;
 assign wire6642 = ( pkey_246_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_254_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6643 = ( wire6642 ) | ( pksi_174_  &  n_n200  &  wire655 ) ;
 assign wire6646 = ( pkey_140_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_148_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6647 = ( wire6646 ) | ( pksi_152_  &  n_n200  &  wire655 ) ;
 assign wire6650 = ( pkey_165_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_173_ ) ;
 assign wire6651 = ( wire6650 ) | ( pksi_151_  &  n_n200  &  wire655 ) ;
 assign wire6654 = ( pkey_158_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_166_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6655 = ( wire6654 ) | ( pksi_154_  &  n_n200  &  wire655 ) ;
 assign wire6658 = ( pkey_92_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_84_ ) ;
 assign wire6659 = ( wire6658 ) | ( pksi_140_  &  n_n200  &  wire655 ) ;
 assign wire6662 = ( pkey_77_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_85_  &  (~ pencrypt_0_) ) ;
 assign wire6663 = ( wire6662 ) | ( n_n2474  &  n_n200  &  wire655 ) ;
 assign wire6666 = ( pkey_110_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_102_ ) ;
 assign wire6667 = ( wire6666 ) | ( n_n168  &  n_n200  &  wire655 ) ;
 assign wire6670 = ( pkey_5_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_13_ ) ;
 assign wire6671 = ( wire6670 ) | ( pksi_108_  &  n_n200  &  wire655 ) ;
 assign wire6674 = ( pkey_251_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_194_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6675 = ( wire6674 ) | ( n_n2268  &  n_n200  &  wire655 ) ;
 assign wire6678 = ( pkey_229_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_237_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6679 = ( wire6678 ) | ( pksi_175_  &  n_n200  &  wire655 ) ;
 assign wire6682 = ( pkey_238_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_246_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6683 = ( wire6682 ) | ( pksi_170_  &  n_n200  &  wire655 ) ;
 assign wire6686 = ( pkey_148_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_156_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6687 = ( wire6686 ) | ( pksi_164_  &  n_n200  &  wire655 ) ;
 assign wire6690 = ( pkey_157_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_165_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6691 = ( wire6690 ) | ( pksi_144_  &  n_n200  &  wire655 ) ;
 assign wire6694 = ( pkey_166_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_174_ ) ;
 assign wire6695 = ( wire6694 ) | ( pksi_167_  &  n_n200  &  wire655 ) ;
 assign wire6698 = ( pkey_76_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_84_ ) ;
 assign wire6699 = ( wire6698 ) | ( pksi_128_  &  n_n200  &  wire655 ) ;
 assign wire6702 = ( pstart_0_  &  pkey_85_  &  pencrypt_0_ ) | ( pkey_93_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6703 = ( wire6702 ) | ( n_n2474  &  (~ n_n200)  &  wire655 ) ;
 assign wire6706 = ( pkey_94_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_102_ ) ;
 assign wire6707 = ( wire6706 ) | ( pksi_130_  &  n_n200  &  wire655 ) ;
 assign wire6710 = ( pstart_0_  &  pencrypt_0_  &  pkey_22_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_30_ ) ;
 assign wire6711 = ( wire6710 ) | ( n_n2517  &  (~ n_n200)  &  wire655 ) ;
 assign wire6714 = ( pkey_136_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_144_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6715 = ( wire6714 ) | ( pksi_67_  &  n_n200  &  wire655 ) ;
 assign wire6718 = ( pkey_66_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_74_  &  (~ pencrypt_0_) ) ;
 assign wire6719 = ( wire6718 ) | ( n_n2333  &  (~ n_n200)  &  wire655 ) ;
 assign wire6722 = ( pkey_89_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_97_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6723 = ( wire6722 ) | ( pksi_46_  &  n_n200  &  wire655 ) ;
 assign wire6726 = ( pkey_112_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_120_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6727 = ( wire6726 ) | ( pksi_47_  &  n_n200  &  wire655 ) ;
 assign wire6730 = ( pkey_50_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_42_ ) ;
 assign wire6731 = ( wire6730 ) | ( pksi_13_  &  n_n200  &  wire655 ) ;
 assign wire6734 = ( pkey_144_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_152_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6735 = ( wire6734 ) | ( pksi_57_  &  n_n200  &  wire655 ) ;
 assign wire6738 = ( pkey_123_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_66_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6739 = ( wire6738 ) | ( n_n2333  &  n_n200  &  wire655 ) ;
 assign wire6742 = ( pkey_97_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_105_ ) ;
 assign wire6743 = ( wire6742 ) | ( pksi_38_  &  n_n200  &  wire655 ) ;
 assign wire6746 = ( pstart_0_  &  pkey_104_  &  pencrypt_0_ ) | ( pkey_112_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6747 = ( wire6746 ) | ( pksi_30_  &  n_n200  &  wire655 ) ;
 assign wire6750 = ( pkey_50_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_58_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6751 = ( wire6750 ) | ( n_n2374  &  n_n200  &  wire655 ) ;
 assign wire6754 = ( pkey_152_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_160_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6755 = ( wire6754 ) | ( pksi_53_  &  n_n200  &  wire655 ) ;
 assign wire6758 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_90_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_82_ ) ;
 assign wire6759 = ( wire6758 ) | ( n_n2337  &  n_n200  &  wire655 ) ;
 assign wire6762 = ( pkey_81_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_73_ ) ;
 assign wire6763 = ( wire6762 ) | ( pksi_32_  &  n_n200  &  wire655 ) ;
 assign wire6766 = ( pkey_96_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_104_  &  (~ pencrypt_0_) ) ;
 assign wire6767 = ( wire6766 ) | ( pksi_39_  &  n_n200  &  wire655 ) ;
 assign wire6770 = ( pkey_58_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_1_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6771 = ( wire6770 ) | ( n_n2374  &  (~ n_n200)  &  wire655 ) ;
 assign wire6774 = ( pkey_56_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_227_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6775 = ( wire6774 ) | ( pksi_4_  &  n_n200  &  wire655 ) ;
 assign wire6778 = ( pkey_160_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_168_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6779 = ( wire6778 ) | ( pksi_63_  &  n_n200  &  wire655 ) ;
 assign wire6782 = ( pstart_0_  &  pkey_74_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_82_ ) ;
 assign wire6783 = ( wire6782 ) | ( pksi_36_  &  n_n200  &  wire655 ) ;
 assign wire6786 = ( pkey_81_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_89_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6787 = ( wire6786 ) | ( pksi_24_  &  n_n200  &  wire655 ) ;
 assign wire6790 = ( pkey_88_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_96_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6791 = ( wire6790 ) | ( pksi_29_  &  n_n200  &  wire655 ) ;
 assign wire6794 = ( pkey_1_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_9_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6795 = ( wire6794 ) | ( pksi_18_  &  n_n200  &  wire655 ) ;
 assign wire6798 = ( pkey_234_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_242_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6799 = ( wire6798 ) | ( pksi_85_  &  n_n200  &  wire655 ) ;
 assign wire6802 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_200_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_192_ ) ;
 assign wire6803 = ( wire6802 ) | ( pksi_89_  &  n_n200  &  wire655 ) ;
 assign wire6806 = ( pkey_130_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_187_ ) ;
 assign wire6807 = ( wire6806 ) | ( n_n2301  &  n_n200  &  wire655 ) ;
 assign wire6810 = ( pkey_145_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_153_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6811 = ( wire6810 ) | ( pksi_48_  &  n_n200  &  wire655 ) ;
 assign wire6814 = ( pkey_9_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_17_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6815 = ( wire6814 ) | ( pksi_8_  &  n_n200  &  wire655 ) ;
 assign wire6818 = ( pkey_242_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_250_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6819 = ( wire6818 ) | ( n_n2277  &  n_n200  &  wire655 ) ;
 assign wire6822 = ( pkey_249_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_192_ ) ;
 assign wire6823 = ( wire6822 ) | ( n_n2288  &  n_n200  &  wire655 ) ;
 assign wire6826 = ( pkey_130_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_138_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6827 = ( wire6826 ) | ( pksi_51_  &  n_n200  &  wire655 ) ;
 assign wire6830 = ( pkey_137_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_145_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6831 = ( wire6830 ) | ( pksi_56_  &  n_n200  &  wire655 ) ;
 assign wire6834 = ( pkey_17_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_25_ ) ;
 assign wire6835 = ( wire6834 ) | ( pksi_0_  &  n_n200  &  wire655 ) ;
 assign wire6838 = ( pkey_250_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_193_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6839 = ( wire6838 ) | ( n_n2277  &  (~ n_n200)  &  wire655 ) ;
 assign wire6842 = ( pstart_0_  &  pkey_208_  &  pencrypt_0_ ) | ( pkey_216_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6843 = ( wire6842 ) | ( pksi_81_  &  n_n200  &  wire655 ) ;
 assign wire6846 = ( pstart_0_  &  pkey_171_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_179_ ) ;
 assign wire6847 = ( wire6846 ) | ( pksi_68_  &  n_n200  &  wire655 ) ;
 assign wire6850 = ( pkey_129_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_137_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6851 = ( wire6850 ) | ( pksi_66_  &  n_n200  &  wire655 ) ;
 assign wire6854 = ( pkey_193_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_201_ ) ;
 assign wire6855 = ( wire6854 ) | ( n_n2280  &  n_n200  &  wire655 ) ;
 assign wire6858 = ( pstart_0_  &  pkey_208_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_200_ ) ;
 assign wire6859 = ( wire6858 ) | ( pksi_91_  &  n_n200  &  wire655 ) ;
 assign wire6862 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_187_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_179_ ) ;
 assign wire6863 = ( wire6862 ) | ( pksi_64_  &  n_n200  &  wire655 ) ;
 assign wire6866 = ( pkey_129_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_186_ ) ;
 assign wire6867 = ( wire6866 ) | ( pksi_49_  &  n_n200  &  wire655 ) ;
 assign wire6870 = ( pkey_209_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_201_ ) ;
 assign wire6871 = ( wire6870 ) | ( pksi_80_  &  n_n200  &  wire655 ) ;
 assign wire6874 = ( pkey_224_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_232_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6875 = ( wire6874 ) | ( pksi_87_  &  n_n200  &  wire655 ) ;
 assign wire6878 = ( pkey_154_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_162_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6879 = ( wire6878 ) | ( pksi_58_  &  n_n200  &  wire655 ) ;
 assign wire6882 = ( pstart_0_  &  pencrypt_0_  &  pkey_177_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_185_ ) ;
 assign wire6883 = ( wire6882 ) | ( pksi_59_  &  n_n200  &  wire655 ) ;
 assign wire6886 = ( pkey_107_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_115_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6887 = ( wire6886 ) | ( pksi_44_  &  n_n200  &  wire655 ) ;
 assign wire6890 = ( pstart_0_  &  pencrypt_0_  &  pkey_65_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_73_ ) ;
 assign wire6891 = ( wire6890 ) | ( pksi_42_  &  n_n200  &  wire655 ) ;
 assign wire6894 = ( pkey_209_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_217_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6895 = ( wire6894 ) | ( pksi_72_  &  n_n200  &  wire655 ) ;
 assign wire6898 = ( pkey_216_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_224_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6899 = ( wire6898 ) | ( pksi_77_  &  n_n200  &  wire655 ) ;
 assign wire6902 = ( pkey_162_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_170_ ) ;
 assign wire6903 = ( wire6902 ) | ( pksi_69_  &  n_n200  &  wire655 ) ;
 assign wire6906 = ( pkey_169_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_177_ ) ;
 assign wire6907 = ( wire6906 ) | ( pksi_50_  &  n_n200  &  wire655 ) ;
 assign wire6910 = ( pkey_115_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_123_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6911 = ( wire6910 ) | ( pksi_40_  &  n_n200  &  wire655 ) ;
 assign wire6914 = ( pkey_122_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_65_ ) ;
 assign wire6915 = ( wire6914 ) | ( n_n2342  &  (~ n_n200)  &  wire655 ) ;
 assign wire6918 = ( pkey_217_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_225_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6919 = ( wire6918 ) | ( pksi_94_  &  n_n200  &  wire655 ) ;
 assign wire6922 = ( pkey_240_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_248_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6923 = ( wire6922 ) | ( pksi_95_  &  n_n200  &  wire655 ) ;
 assign wire6926 = ( pkey_138_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_146_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6927 = ( wire6926 ) | ( pksi_60_  &  n_n200  &  wire655 ) ;
 assign wire6930 = ( pkey_161_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_169_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6931 = ( wire6930 ) | ( pksi_62_  &  n_n200  &  wire655 ) ;
 assign wire6934 = ( pkey_80_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_72_ ) ;
 assign wire6935 = ( wire6934 ) | ( pksi_43_  &  n_n200  &  wire655 ) ;
 assign wire6938 = ( pkey_2_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_10_ ) ;
 assign wire6939 = ( wire6938 ) | ( n_n2365  &  (~ n_n200)  &  wire655 ) ;
 assign wire6942 = ( pkey_225_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_233_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6943 = ( wire6942 ) | ( pksi_86_  &  n_n200  &  wire655 ) ;
 assign wire6946 = ( pkey_232_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_240_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6947 = ( wire6946 ) | ( pksi_78_  &  n_n200  &  wire655 ) ;
 assign wire6950 = ( pkey_146_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_154_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6951 = ( wire6950 ) | ( n_n2305  &  n_n200  &  wire655 ) ;
 assign wire6954 = ( pkey_153_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_161_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6955 = ( wire6954 ) | ( pksi_70_  &  n_n200  &  wire655 ) ;
 assign wire6958 = ( pkey_80_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_88_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6959 = ( wire6958 ) | ( pksi_33_  &  n_n200  &  wire655 ) ;
 assign wire6962 = ( pkey_59_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_2_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6963 = ( wire6962 ) | ( n_n2365  &  n_n200  &  wire655 ) ;
 assign wire6966 = ( pkey_233_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_241_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6967 = ( wire6966 ) | ( pksi_74_  &  n_n200  &  wire655 ) ;
 assign wire6970 = ( pkey_163_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  pkey_171_  &  (~ pencrypt_0_) ) ;
 assign wire6971 = ( wire6970 ) | ( pksi_55_  &  n_n200  &  wire655 ) ;
 assign wire6974 = ( pkey_168_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_176_ ) ;
 assign wire6975 = ( wire6974 ) | ( pksi_54_  &  n_n200  &  wire655 ) ;
 assign wire6978 = ( pkey_98_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_106_ ) ;
 assign wire6979 = ( wire6978 ) | ( pksi_45_  &  n_n200  &  wire655 ) ;
 assign wire6982 = ( pkey_121_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_64_ ) ;
 assign wire6983 = ( wire6982 ) | ( n_n2352  &  n_n200  &  wire655 ) ;
 assign wire6986 = ( pstart_0_  &  pkey_51_  &  pencrypt_0_ ) | ( pkey_59_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6987 = ( wire6986 ) | ( pksi_16_  &  n_n200  &  wire655 ) ;
 assign wire6990 = ( pkey_18_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_10_ ) ;
 assign wire6991 = ( wire6990 ) | ( pksi_12_  &  n_n200  &  wire655 ) ;
 assign wire6994 = ( pkey_241_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_249_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6995 = ( wire6994 ) | ( pksi_83_  &  n_n200  &  wire655 ) ;
 assign wire6998 = ( pkey_248_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_163_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire6999 = ( wire6998 ) | ( pksi_76_  &  n_n200  &  wire655 ) ;
 assign wire7002 = ( pstart_0_  &  pencrypt_0_  &  pkey_176_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_184_ ) ;
 assign wire7003 = ( wire7002 ) | ( pksi_71_  &  n_n200  &  wire655 ) ;
 assign wire7006 = ( pkey_98_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_90_ ) ;
 assign wire7007 = ( wire7006 ) | ( n_n2337  &  (~ n_n200)  &  wire655 ) ;
 assign wire7010 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_72_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_64_ ) ;
 assign wire7011 = ( wire7010 ) | ( n_n2352  &  (~ n_n200)  &  wire655 ) ;
 assign wire7014 = ( pstart_0_  &  pkey_51_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_43_ ) ;
 assign wire7015 = ( wire7014 ) | ( pksi_20_  &  n_n200  &  wire655 ) ;
 assign wire7018 = ( pkey_18_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_26_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7019 = ( wire7018 ) | ( n_n2369  &  n_n200  &  wire655 ) ;
 assign wire7022 = ( pstart_0_  &  pencrypt_0_  &  pkey_170_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_178_ ) ;
 assign wire7023 = ( wire7022 ) | ( pksi_61_  &  n_n200  &  wire655 ) ;
 assign wire7026 = ( pkey_128_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_136_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7027 = ( wire7026 ) | ( n_n2320  &  (~ n_n200)  &  wire655 ) ;
 assign wire7030 = ( pkey_99_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_184_ ) ;
 assign wire7031 = ( wire7030 ) | ( pksi_52_  &  n_n200  &  wire655 ) ;
 assign wire7034 = ( pkey_114_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_122_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7035 = ( wire7034 ) | ( n_n2342  &  n_n200  &  wire655 ) ;
 assign wire7038 = ( pkey_113_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_105_ ) ;
 assign wire7039 = ( wire7038 ) | ( pksi_26_  &  n_n200  &  wire655 ) ;
 assign wire7042 = ( pstart_0_  &  pencrypt_0_  &  pkey_35_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_43_ ) ;
 assign wire7043 = ( wire7042 ) | ( pksi_7_  &  n_n200  &  wire655 ) ;
 assign wire7046 = ( pkey_26_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_34_ ) ;
 assign wire7047 = ( wire7046 ) | ( n_n2369  &  (~ n_n200)  &  wire655 ) ;
 assign wire7050 = ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_186_ ) | ( pstart_0_  &  pencrypt_0_  &  pkey_178_ ) ;
 assign wire7051 = ( wire7050 ) | ( n_n2310  &  n_n200  &  wire655 ) ;
 assign wire7054 = ( pkey_128_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_185_ ) ;
 assign wire7055 = ( wire7054 ) | ( n_n2320  &  n_n200  &  wire655 ) ;
 assign wire7058 = ( pkey_99_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_107_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7059 = ( wire7058 ) | ( pksi_31_  &  n_n200  &  wire655 ) ;
 assign wire7062 = ( pkey_114_  &  pstart_0_  &  (~ pencrypt_0_) ) | ( pstart_0_  &  pencrypt_0_  &  pkey_106_ ) ;
 assign wire7063 = ( wire7062 ) | ( pksi_37_  &  n_n200  &  wire655 ) ;
 assign wire7066 = ( pkey_113_  &  pstart_0_  &  pencrypt_0_ ) | ( pkey_121_  &  pstart_0_  &  (~ pencrypt_0_) ) ;
 assign wire7067 = ( wire7066 ) | ( pksi_35_  &  n_n200  &  wire655 ) ;
 assign wire7070 = ( pkey_120_  &  pstart_0_  &  pencrypt_0_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_35_ ) ;
 assign wire7071 = ( wire7070 ) | ( pksi_28_  &  n_n200  &  wire655 ) ;
 assign wire7074 = ( pstart_0_  &  pencrypt_0_  &  pkey_34_ ) | ( pstart_0_  &  (~ pencrypt_0_)  &  pkey_42_ ) ;
 assign wire7075 = ( wire7074 ) | ( pksi_21_  &  n_n200  &  wire655 ) ;
 assign wire7079 = ( (~ pcount_1_)  &  (~ pcount_0_)  &  (~ pstart_0_)  &  (~ pencrypt_0_) ) ;
 assign wire7081 = ( pcount_2_  &  (~ pencrypt_0_) ) | ( (~ pcount_2_)  &  (~ pstart_0_)  &  pencrypt_0_ ) ;
 assign wire7084 = ( (~ n_n2530) ) | ( wire664 ) | ( (~ pcount_2_)  &  wire653 ) ;


endmodule

