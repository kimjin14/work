module s38584 (
	pg115, pg126, pg116, pg125, pg5, pg135, pg127, pg100, 
	pg6751, pg99, pg6750, pg120, pg134, pg113, pg124, pg114, pg92, pg6748, 
	pg91, pg6749, pclk, pg6746, pg84, pg6747, pg6744, pg6745, pg6753, pg6752, 
	pg56, pg57, pg64, pg73, pg36, pg54, pg72, pg90, pg35, pg44, 
	pg53, pg8342, pg8353, pg8870, pg9048, pg9741, pg13272, pg13906, pg28030, pg28041, 
	pg33533, pg34437, pg8132, pg8783, pg9555, pg12184, pg13068, pg13099, pg31521, pg33435, 
	pg34425, pg7260, pg8344, pg8784, pg14167, pg17320, pg18101, pg30327, pg31793, pg34435, 
	pg8398, pg8785, pg18100, pg20899, pg34436, pg8786, pg14828, pg20557, pg20654, pg21727, 
	pg24171, pg24182, pg26876, pg30329, pg33894, pg34239, pg7243, pg7540, pg8235, pg8787, 
	pg12470, pg17819, pg19334, pg24172, pg24181, pg26877, pg32454, pg34597, pg8403, pg8788, 
	pg9497, pg13926, pg14189, pg14451, pg23190, pg24151, pg24162, pg24180, pg26801, pg33874, 
	pg34237, pg7245, pg8215, pg8789, pg10122, pg12919, pg16924, pg17291, pg20763, pg24161, 
	pg24170, pg28042, pg34238, pg12833, pg14705, pg14738, pg14749, pg16693, pg16718, pg17423, 
	pg18097, pg24164, pg24175, pg29211, pg34235, pg18098, pg20901, pg23652, pg24163, pg24176, 
	pg24185, pg29210, pg34201, pg34236, pg11388, pg17577, pg17674, pg17760, pg18099, pg20652, 
	pg24166, pg24173, pg24184, pg29213, pg29220, pg34233, pg34972, pg14597, pg14694, pg17813, 
	pg21292, pg24165, pg24174, pg24183, pg29212, pg29221, pg32975, pg34234, pg34788, pg11678, 
	pg12923, pg14518, pg14662, pg14673, pg17607, pg17715, pg19357, pg24168, pg24179, pg25219, 
	pg29215, pg30332, pg34956, pg16627, pg23612, pg24167, pg29214, pg34232, pg14635, pg17519, 
	pg17580, pg24177, pg25167, pg29217, pg30330, pg34240, pg12832, pg16722, pg24169, pg24178, 
	pg29216, pg30331, pg34221, pg7916, pg8919, pg11447, pg13881, pg16624, pg17711, pg17722, 
	pg20049, pg25259, pg25583, pg29219, pg33948, pg33959, pg34927, pg8918, pg11770, pg16874, 
	pg17604, pg21245, pg25584, pg29218, pg33949, pg34917, pg25585, pg32185, pg33946, pg34839, 
	pg8839, pg16603, pg16656, pg16744, pg17646, pg17743, pg17778, pg17787, pg18092, pg25586, 
	pg33947, pg34919, pg11418, pg16686, pg17845, pg21176, pg25114, pg25590, pg34383, pg34923, 
	pg12368, pg13895, pg14779, pg17639, pg17688, pg18094, pg18881, pg23683, pg33079, pg33945, 
	pg34913, pg10527, pg13865, pg16659, pg17649, pg17678, pg17685, pg17739, pg17764, pg18095, 
	pg33935, pg34925, pg11349, pg13259, pg16748, pg16775, pg17316, pg17404, pg17871, pg18096, 
	pg21270, pg25582, pg34915, pg8416, pg9617, pg31863, pg33659, pg33950, pg7257, pg8920, 
	pg9251, pg9817, pg13966, pg14217, pg27831, pg31861, pg34921, pg8291, pg12238, pg12300, 
	pg14096, pg14201, pg14421, pg16955, pg17400, pg26875, pg31862, pg32429, pg8283, pg8915, 
	pg9019, pg9682, pg12350, pg12422, pg13049, pg13085, pg14125, pg14147, pg25587, pg31665, 
	pg8279, pg21698, pg25588, pg31860, pg8719, pg8917, pg9615, pg9680, pg9743, pg23002, 
	pg25589, pg28753, pg31656, pg33636, pg7946, pg8178, pg8277, pg8358, pg8475, pg8916, 
	pg9553, pg10306, pg10500, pg13039, pg23759);

input pg115;
input pg126;
input pg116;
input pg125;
input pg5;
input pg135;
input pg127;
input pg100;
input pg6751;
input pg99;
input pg6750;
input pg120;
input pg134;
input pg113;
input pg124;
input pg114;
input pg92;
input pg6748;
input pg91;
input pg6749;
input pclk;
input pg6746;
input pg84;
input pg6747;
input pg6744;
input pg6745;
input pg6753;
input pg6752;
input pg56;
input pg57;
input pg64;
input pg73;
input pg36;
input pg54;
input pg72;
input pg90;
input pg35;
input pg44;
input pg53;
output pg8342;
output pg8353;
output pg8870;
output pg9048;
output pg9741;
output pg13272;
output pg13906;
output pg28030;
output pg28041;
output pg33533;
output pg34437;
output pg8132;
output pg8783;
output pg9555;
output pg12184;
output pg13068;
output pg13099;
output pg31521;
output pg33435;
output pg34425;
output pg7260;
output pg8344;
output pg8784;
output pg14167;
output pg17320;
output pg18101;
output pg30327;
output pg31793;
output pg34435;
output pg8398;
output pg8785;
output pg18100;
output pg20899;
output pg34436;
output pg8786;
output pg14828;
output pg20557;
output pg20654;
output pg21727;
output pg24171;
output pg24182;
output pg26876;
output pg30329;
output pg33894;
output pg34239;
output pg7243;
output pg7540;
output pg8235;
output pg8787;
output pg12470;
output pg17819;
output pg19334;
output pg24172;
output pg24181;
output pg26877;
output pg32454;
output pg34597;
output pg8403;
output pg8788;
output pg9497;
output pg13926;
output pg14189;
output pg14451;
output pg23190;
output pg24151;
output pg24162;
output pg24180;
output pg26801;
output pg33874;
output pg34237;
output pg7245;
output pg8215;
output pg8789;
output pg10122;
output pg12919;
output pg16924;
output pg17291;
output pg20763;
output pg24161;
output pg24170;
output pg28042;
output pg34238;
output pg12833;
output pg14705;
output pg14738;
output pg14749;
output pg16693;
output pg16718;
output pg17423;
output pg18097;
output pg24164;
output pg24175;
output pg29211;
output pg34235;
output pg18098;
output pg20901;
output pg23652;
output pg24163;
output pg24176;
output pg24185;
output pg29210;
output pg34201;
output pg34236;
output pg11388;
output pg17577;
output pg17674;
output pg17760;
output pg18099;
output pg20652;
output pg24166;
output pg24173;
output pg24184;
output pg29213;
output pg29220;
output pg34233;
output pg34972;
output pg14597;
output pg14694;
output pg17813;
output pg21292;
output pg24165;
output pg24174;
output pg24183;
output pg29212;
output pg29221;
output pg32975;
output pg34234;
output pg34788;
output pg11678;
output pg12923;
output pg14518;
output pg14662;
output pg14673;
output pg17607;
output pg17715;
output pg19357;
output pg24168;
output pg24179;
output pg25219;
output pg29215;
output pg30332;
output pg34956;
output pg16627;
output pg23612;
output pg24167;
output pg29214;
output pg34232;
output pg14635;
output pg17519;
output pg17580;
output pg24177;
output pg25167;
output pg29217;
output pg30330;
output pg34240;
output pg12832;
output pg16722;
output pg24169;
output pg24178;
output pg29216;
output pg30331;
output pg34221;
output pg7916;
output pg8919;
output pg11447;
output pg13881;
output pg16624;
output pg17711;
output pg17722;
output pg20049;
output pg25259;
output pg25583;
output pg29219;
output pg33948;
output pg33959;
output pg34927;
output pg8918;
output pg11770;
output pg16874;
output pg17604;
output pg21245;
output pg25584;
output pg29218;
output pg33949;
output pg34917;
output pg25585;
output pg32185;
output pg33946;
output pg34839;
output pg8839;
output pg16603;
output pg16656;
output pg16744;
output pg17646;
output pg17743;
output pg17778;
output pg17787;
output pg18092;
output pg25586;
output pg33947;
output pg34919;
output pg11418;
output pg16686;
output pg17845;
output pg21176;
output pg25114;
output pg25590;
output pg34383;
output pg34923;
output pg12368;
output pg13895;
output pg14779;
output pg17639;
output pg17688;
output pg18094;
output pg18881;
output pg23683;
output pg33079;
output pg33945;
output pg34913;
output pg10527;
output pg13865;
output pg16659;
output pg17649;
output pg17678;
output pg17685;
output pg17739;
output pg17764;
output pg18095;
output pg33935;
output pg34925;
output pg11349;
output pg13259;
output pg16748;
output pg16775;
output pg17316;
output pg17404;
output pg17871;
output pg18096;
output pg21270;
output pg25582;
output pg34915;
output pg8416;
output pg9617;
output pg31863;
output pg33659;
output pg33950;
output pg7257;
output pg8920;
output pg9251;
output pg9817;
output pg13966;
output pg14217;
output pg27831;
output pg31861;
output pg34921;
output pg8291;
output pg12238;
output pg12300;
output pg14096;
output pg14201;
output pg14421;
output pg16955;
output pg17400;
output pg26875;
output pg31862;
output pg32429;
output pg8283;
output pg8915;
output pg9019;
output pg9682;
output pg12350;
output pg12422;
output pg13049;
output pg13085;
output pg14125;
output pg14147;
output pg25587;
output pg31665;
output pg8279;
output pg21698;
output pg25588;
output pg31860;
output pg8719;
output pg8917;
output pg9615;
output pg9680;
output pg9743;
output pg23002;
output pg25589;
output pg28753;
output pg31656;
output pg33636;
output pg7946;
output pg8178;
output pg8277;
output pg8358;
output pg8475;
output pg8916;
output pg9553;
output pg10306;
output pg10500;
output pg13039;
output pg23759;
wire ng33063;
wire ng34455;
wire ng24264;
wire ng26917;
wire ng33013;
wire ng26951;
wire ng24281;
wire ng30338;
wire ng30403;
wire ng34610;
wire ng33537;
wire ng25595;
wire ng34446;
wire ng34266;
wire ng24205;
wire ng26907;
wire ng33962;
wire ng32983;
wire ng34030;
wire ng24277;
wire ng34605;
wire ng29283;
wire ng33033;
wire ng25678;
wire ng34598;
wire ng33553;
wire ng33023;
wire ng25600;
wire ng24207;
wire ng34249;
wire ng30343;
wire ng30551;
wire ng24341;
wire ng30546;
wire ng29294;
wire ng26893;
wire ng29238;
wire ng24347;
wire ng29270;
wire ng26883;
wire ng25609;
wire ng25662;
wire ng33581;
wire ng34803;
wire ng30334;
wire ng33964;
wire ng34600;
wire ng33608;
wire ng24263;
wire ng33980;
wire ng30353;
wire ng29302;
wire ng33996;
wire ng32992;
wire ng26889;
wire ng34445;
wire ng30537;
wire ng25670;
wire ng28044;
wire ng29242;
wire ng34799;
wire ng30346;
wire ng33994;
wire ng34601;
wire ng34722;
wire ng30454;
wire ng24258;
wire ng30492;
wire ng30437;
wire ng25687;
wire ng29257;
wire ng25682;
wire ng33987;
wire ng30424;
wire ng34727;
wire ng29303;
wire ng32981;
wire ng30526;
wire ng33997;
wire ng29296;
wire ng33042;
wire ng25697;
wire ng30444;
wire ng29230;
wire ng30438;
wire ng24278;
wire ng25654;
wire ng30558;
wire ng33601;
wire ng29275;
wire ng29237;
wire ng29306;
wire ng30350;
wire ng33985;
wire ng30377;
wire ng24208;
wire ng26884;
wire ng25701;
wire ng24348;
wire ng33559;
wire ng30392;
wire ng25667;
wire ng33050;
wire ng25610;
wire ng29309;
wire ng33062;
wire ng24240;
wire ng29264;
wire ng28063;
wire ng34639;
wire ng30549;
wire ng26924;
wire ng34020;
wire ng33970;
wire ng33594;
wire ng30488;
wire ng34604;
wire ng30469;
wire ng26912;
wire ng24204;
wire ng34467;
wire ng34613;
wire ng24349;
wire ng21898;
wire ng26927;
wire ng30507;
wire ng28092;
wire ng26914;
wire ng26948;
wire ng30430;
wire ng34037;
wire ng26952;
wire ng26939;
wire ng30355;
wire ng33620;
wire ng34024;
wire ng29233;
wire ng33040;
wire ng34630;
wire ng33617;
wire ng24260;
wire ng21897;
wire ng25598;
wire ng32977;
wire ng25656;
wire ng28051;
wire ng30528;
wire ng33588;
wire ng34795;
wire ng26946;
wire ng28099;
wire ng30502;
wire ng26899;
wire ng33573;
wire ng30481;
wire ng26955;
wire ng34250;
wire ng25703;
wire ng26922;
wire ng30451;
wire ng30337;
wire ng31902;
wire ng25611;
wire ng33989;
wire ng30486;
wire ng31903;
wire ng30362;
wire ng34801;
wire ng29269;
wire ng33967;
wire ng33055;
wire ng24201;
wire ng25591;
wire ng25714;
wire ng30411;
wire ng28050;
wire ng34458;
wire ng28072;
wire ng33961;
wire ng24238;
wire ng33038;
wire ng25761;
wire ng30468;
wire ng28057;
wire ng26910;
wire ng24266;
wire ng30509;
wire ng25756;
wire ng24215;
wire ng34009;
wire ng34725;
wire ng34017;
wire ng30442;
wire ng34264;
wire ng25630;
wire ng30562;
wire ng34616;
wire ng33070;
wire ng29289;
wire ng25628;
wire ng33555;
wire ng29281;
wire ng24352;
wire ng34791;
wire ng29284;
wire ng30426;
wire ng30515;
wire ng33068;
wire ng34443;
wire ng26944;
wire ng31898;
wire ng25705;
wire ng34026;
wire ng30457;
wire ng30390;
wire ng30404;
wire ng29236;
wire ng21895;
wire ng24269;
wire ng34448;
wire ng25650;
wire ng33036;
wire ng30341;
wire ng30540;
wire ng34730;
wire ng25763;
wire ng24282;
wire ng34451;
wire ng25729;
wire ng34980;
wire ng24254;
wire ng29235;
wire ng34003;
wire ng25715;
wire ng33149;
wire ng33197;
wire ng28089;
wire ng30463;
wire ng33562;
wire ng33546;
wire ng24272;
wire ng34628;
wire ng34027;
wire ng28055;
wire ng31865;
wire ng32985;
wire ng26931;
wire ng29244;
wire ng34439;
wire ng34849;
wire ng34459;
wire ng30363;
wire ng24247;
wire ng30365;
wire ng29300;
wire ng33591;
wire ng33626;
wire ng29305;
wire ng33570;
wire ng30484;
wire ng34256;
wire ng34011;
wire ng33590;
wire ng29240;
wire ng25699;
wire ng26934;
wire ng25636;
wire ng30344;
wire ng34633;
wire ng30399;
wire ng30561;
wire ng30520;
wire ng30409;
wire ng34805;
wire ng33599;
wire ng30410;
wire ng31895;
wire ng34619;
wire ng25664;
wire ng25653;
wire ng30412;
wire ng25681;
wire ng30395;
wire ng30380;
wire ng30405;
wire ng30476;
wire ng33560;
wire ng24236;
wire ng33029;
wire ng24280;
wire ng30370;
wire ng25749;
wire ng30538;
wire ng34025;
wire ng31899;
wire ng30531;
wire ng33619;
wire ng26903;
wire ng29268;
wire ng33067;
wire ng26923;
wire ng28085;
wire ng33583;
wire ng26909;
wire ng24355;
wire ng29304;
wire ng26926;
wire ng34796;
wire ng33598;
wire ng30559;
wire ng28087;
wire ng33012;
wire ng28060;
wire ng33540;
wire ng33627;
wire ng34615;
wire ng34040;
wire ng29267;
wire ng34251;
wire ng29243;
wire ng26950;
wire ng25634;
wire ng29227;
wire ng26896;
wire ng25764;
wire ng29286;
wire ng28091;
wire ng33545;
wire ng29297;
wire ng33577;
wire ng30357;
wire ng30544;
wire ng30358;
wire ng30367;
wire ng31866;
wire ng25683;
wire ng29246;
wire ng25734;
wire ng21892;
wire ng25706;
wire ng28093;
wire ng33016;
wire ng24353;
wire ng25655;
wire ng34642;
wire ng25704;
wire ng33008;
wire ng30421;
wire ng33007;
wire ng25730;
wire ng25624;
wire ng34255;
wire ng30371;
wire ng26900;
wire ng33607;
wire ng26904;
wire ng34626;
wire ng29293;
wire ng34268;
wire ng29271;
wire ng28083;
wire ng26886;
wire ng33576;
wire ng29266;
wire ng34260;
wire ng33618;
wire ng34640;
wire ng30445;
wire ng30514;
wire ng30356;
wire ng25685;
wire ng30525;
wire ng30342;
wire ng30560;
wire ng33567;
wire ng29290;
wire ng25602;
wire ng33544;
wire ng34606;
wire ng34013;
wire ng30441;
wire ng33977;
wire ng34621;
wire ng26908;
wire ng34257;
wire ng29299;
wire ng30470;
wire ng26954;
wire ng21901;
wire ng33574;
wire ng34607;
wire ng33011;
wire ng26965;
wire ng30429;
wire ng25619;
wire ng30414;
wire ng33541;
wire ng33615;
wire ng33548;
wire ng33053;
wire ng25750;
wire ng34622;
wire ng25720;
wire ng34804;
wire ng30543;
wire ng34005;
wire ng30383;
wire ng34647;
wire ng29255;
wire ng30523;
wire ng24211;
wire ng33556;
wire ng24214;
wire ng25700;
wire ng25691;
wire ng29261;
wire ng27511;
wire ng33561;
wire ng34641;
wire ng29245;
wire ng30435;
wire ng34006;
wire ng34038;
wire ng21899;
wire ng30391;
wire ng29228;
wire ng25696;
wire ng34029;
wire ng26929;
wire ng30548;
wire ng30364;
wire ng30431;
wire ng33003;
wire ng33014;
wire ng25631;
wire ng26916;
wire ng24246;
wire ng32987;
wire ng33558;
wire ng34468;
wire ng34732;
wire ng25626;
wire ng33592;
wire ng25762;
wire ng25597;
wire ng33986;
wire ng25690;
wire ng29288;
wire ng33212;
wire ng33586;
wire ng30373;
wire ng29229;
wire ng34614;
wire ng33611;
wire ng33041;
wire ng32997;
wire ng29226;
wire ng26966;
wire ng34034;
wire ng24253;
wire ng26920;
wire ng30369;
wire ng25721;
wire ng21891;
wire ng30506;
wire ng25747;
wire ng30440;
wire ng33597;
wire ng30475;
wire ng33034;
wire ng30472;
wire ng34634;
wire ng26890;
wire ng34797;
wire ng32982;
wire ng34629;
wire ng33031;
wire ng32989;
wire ng28069;
wire ng25615;
wire ng25719;
wire ng30493;
wire ng25639;
wire ng30448;
wire ng25593;
wire ng34254;
wire ng34631;
wire ng30467;
wire ng34465;
wire ng33578;
wire ng25702;
wire ng34650;
wire ng24202;
wire ng26919;
wire ng28049;
wire ng33998;
wire ng26913;
wire ng28059;
wire ng24342;
wire ng34010;
wire ng28096;
wire ng24273;
wire ng26928;
wire ng25596;
wire ng28056;
wire ng28053;
wire ng29260;
wire ng34261;
wire ng24345;
wire ng30458;
wire ng24276;
wire ng30483;
wire ng32978;
wire ng33976;
wire ng34729;
wire ng26947;
wire ng25625;
wire ng33552;
wire ng25622;
wire ng26892;
wire ng25757;
wire ng26901;
wire ng33058;
wire ng33534;
wire ng26932;
wire ng33035;
wire ng33060;
wire ng24233;
wire ng25612;
wire ng24335;
wire ng31900;
wire ng34624;
wire ng30345;
wire ng26895;
wire ng21900;
wire ng33045;
wire ng25744;
wire ng30532;
wire ng25708;
wire ng24257;
wire ng34450;
wire ng30471;
wire ng33542;
wire ng31904;
wire ng28088;
wire ng25698;
wire ng34728;
wire ng30461;
wire ng34618;
wire ng33609;
wire ng29259;
wire ng30361;
wire ng24338;
wire ng26958;
wire ng33981;
wire ng30381;
wire ng24337;
wire ng30499;
wire ng24239;
wire ng26897;
wire ng26891;
wire ng33024;
wire ng34447;
wire ng33971;
wire ng29295;
wire ng30402;
wire ng26961;
wire ng30487;
wire ng30552;
wire ng25677;
wire ng26949;
wire ng26967;
wire ng33018;
wire ng30452;
wire ng34611;
wire ng30556;
wire ng30415;
wire ng29307;
wire ng30413;
wire ng30433;
wire ng30511;
wire ng28086;
wire ng34039;
wire ng30340;
wire ng30512;
wire ng24234;
wire ng34793;
wire ng24241;
wire ng30359;
wire ng33176;
wire ng33047;
wire ng25638;
wire ng34466;
wire ng30563;
wire ng34612;
wire ng34449;
wire ng30400;
wire ng30407;
wire ng30500;
wire ng34911;
wire ng32994;
wire ng34035;
wire ng34259;
wire ng34800;
wire ng30504;
wire ng24210;
wire ng34462;
wire ng26915;
wire ng30436;
wire ng31894;
wire ng33039;
wire ng24261;
wire ng33623;
wire ng30530;
wire ng30524;
wire ng25716;
wire ng32976;
wire ng34719;
wire ng34262;
wire ng30485;
wire ng30460;
wire ng33009;
wire ng26956;
wire ng33536;
wire ng32980;
wire ng29253;
wire ng34456;
wire ng30379;
wire ng30382;
wire ng34018;
wire ng30443;
wire ng33988;
wire ng34265;
wire ng33572;
wire ng34016;
wire ng29247;
wire ng25637;
wire ng30397;
wire ng30351;
wire ng26918;
wire ng30408;
wire ng30503;
wire ng24298;
wire ng25742;
wire ng25635;
wire ng33044;
wire ng30394;
wire ng33568;
wire ng24271;
wire ng33963;
wire ng34636;
wire ng29298;
wire ng30474;
wire ng34625;
wire ng34798;
wire ng24350;
wire ng33613;
wire ng29265;
wire ng29276;
wire ng33059;
wire ng29278;
wire ng34253;
wire ng30542;
wire ng28102;
wire ng24268;
wire ng30349;
wire ng33219;
wire ng30422;
wire ng33587;
wire ng33603;
wire ng26888;
wire ng34453;
wire ng34021;
wire ng34440;
wire ng34794;
wire ng33164;
wire ng26968;
wire ng29285;
wire ng33582;
wire ng24231;
wire ng33065;
wire ng30522;
wire ng24334;
wire ng34000;
wire ng28071;
wire ng33566;
wire ng34635;
wire ng30398;
wire ng31871;
wire ng33000;
wire ng29241;
wire ng29234;
wire ng25733;
wire ng29222;
wire ng25686;
wire ng30385;
wire ng34623;
wire ng34457;
wire ng34441;
wire ng30420;
wire ng34790;
wire ng34627;
wire ng34806;
wire ng34637;
wire ng34263;
wire ng34041;
wire ng28090;
wire ng25669;
wire ng28084;
wire ng33593;
wire ng34638;
wire ng33975;
wire ng25648;
wire ng32979;
wire ng24242;
wire ng32990;
wire ng26894;
wire ng34792;
wire ng24262;
wire ng25627;
wire ng29272;
wire ng34033;
wire ng29292;
wire ng33984;
wire ng24213;
wire ng30518;
wire ng30456;
wire ng33017;
wire ng28052;
wire ng30347;
wire ng34004;
wire ng34850;
wire ng33604;
wire ng33600;
wire ng26969;
wire ng33969;
wire ng26880;
wire ng26902;
wire ng34599;
wire ng25617;
wire ng25614;
wire ng26962;
wire ng34269;
wire ng33606;
wire ng33596;
wire ng34620;
wire ng30536;
wire ng26882;
wire ng25632;
wire ng28054;
wire ng33992;
wire ng28048;
wire ng24343;
wire ng26964;
wire ng33982;
wire ng33625;
wire ng29282;
wire ng28070;
wire ng24250;
wire ng34643;
wire ng24237;
wire ng24206;
wire ng30480;
wire ng30455;
wire ng25748;
wire ng30336;
wire ng30497;
wire ng32986;
wire ng34880;
wire ng24245;
wire ng33037;
wire ng33999;
wire ng29250;
wire ng33019;
wire ng33595;
wire ng34022;
wire ng30557;
wire ng33032;
wire ng33602;
wire ng33612;
wire ng26906;
wire ng30450;
wire ng30339;
wire ng34464;
wire ng30428;
wire ng34028;
wire ng30401;
wire ng33569;
wire ng30501;
wire ng33204;
wire ng34720;
wire ng28043;
wire ng26930;
wire ng25592;
wire ng33622;
wire ng26938;
wire ng28058;
wire ng33054;
wire ng30464;
wire ng34731;
wire ng33551;
wire ng33048;
wire ng26925;
wire ng30465;
wire ng29274;
wire ng34002;
wire ng25649;
wire ng26887;
wire ng29308;
wire ng33621;
wire ng30449;
wire ng31864;
wire ng32988;
wire ng30535;
wire ng32993;
wire ng34019;
wire ng25663;
wire ng25594;
wire ng33624;
wire ng33539;
wire ng30348;
wire ng30335;
wire ng24251;
wire ng29239;
wire ng33584;
wire ng30419;
wire ng28047;
wire ng33027;
wire ng29273;
wire ng25601;
wire ng34442;
wire ng30539;
wire ng33187;
wire ng26905;
wire ng30459;
wire ng30378;
wire ng26970;
wire ng33610;
wire ng31870;
wire ng34463;
wire ng33575;
wire ng26957;
wire ng28045;
wire ng33614;
wire ng26898;
wire ng28066;
wire ng24203;
wire ng29224;
wire ng30375;
wire ng33015;
wire ng30529;
wire ng33990;
wire ng25605;
wire ng30406;
wire ng34721;
wire ng25695;
wire ng34808;
wire ng26921;
wire ng34724;
wire ng33021;
wire ng33557;
wire ng33563;
wire ng29225;
wire ng32984;
wire ng30508;
wire ng34444;
wire ng30547;
wire ng28073;
wire ng25735;
wire ng30417;
wire ng33547;
wire ng33549;
wire ng25707;
wire ng33001;
wire ng31901;
wire ng33616;
wire ng30434;
wire ng30479;
wire ng34258;
wire ng18597;
wire ng30473;
wire ng34735;
wire ng34007;
wire ng26963;
wire ng25676;
wire ng30453;
wire ng24336;
wire ng32996;
wire ng30521;
wire ng30510;
wire ng30495;
wire ng34023;
wire ng24209;
wire ng33972;
wire ng33993;
wire ng30366;
wire ng34014;
wire ng26940;
wire ng30555;
wire ng30418;
wire ng33960;
wire ng30517;
wire ng30553;
wire ng25629;
wire ng30462;
wire ng33978;
wire ng33589;
wire ng34726;
wire ng33006;
wire ng30516;
wire ng34603;
wire ng25618;
wire ng26933;
wire ng24346;
wire ng32991;
wire ng30368;
wire ng24243;
wire ng31896;
wire ng30423;
wire ng25722;
wire ng34454;
wire ng32995;
wire ng28105;
wire ng33057;
wire ng25758;
wire ng30478;
wire ng29251;
wire ng28082;
wire ng24249;
wire ng21896;
wire ng24270;
wire ng33580;
wire ng33564;
wire ng29232;
wire ng34008;
wire ng33565;
wire ng24351;
wire ng30396;
wire ng33979;
wire ng30386;
wire ng30376;
wire ng24339;
wire ng30550;
wire ng34608;
wire ng29249;
wire ng33010;
wire ng29280;
wire ng30491;
wire ng29256;
wire ng34461;
wire ng29231;
wire ng34723;
wire ng24252;
wire ng34252;
wire ng34015;
wire ng30427;
wire ng33535;
wire ng25621;
wire ng33028;
wire ng33543;
wire ng30489;
wire ng24256;
wire ng21894;
wire ng30534;
wire ng34807;
wire ng29258;
wire ng30352;
wire ng29301;
wire ng34452;
wire ng31869;
wire ng25599;
wire ng33046;
wire ng34031;
wire ng30490;
wire ng34644;
wire ng25604;
wire ng34881;
wire ng33966;
wire ng34460;
wire ng24235;
wire ng33991;
wire ng24279;
wire ng30388;
wire ng33005;
wire ng33064;
wire ng33550;
wire ng30360;
wire ng34036;
wire ng24267;
wire ng29291;
wire ng33538;
wire ng30416;
wire ng24216;
wire ng24344;
wire ng33973;
wire ng30374;
wire ng29254;
wire ng33002;
wire ng21893;
wire ng30466;
wire ng29262;
wire ng30482;
wire ng28074;
wire ng24248;
wire ng33968;
wire ng25736;
wire ng34733;
wire ng29223;
wire ng29263;
wire ng34609;
wire ng34032;
wire ng34602;
wire ng34012;
wire ng30477;
wire ng30354;
wire ng26945;
wire ng34617;
wire ng24232;
wire ng29248;
wire ng24340;
wire ng30533;
wire ng33049;
wire ng31868;
wire ng30513;
wire ng33052;
wire ng34632;
wire ng33579;
wire ng32998;
wire ng24255;
wire ng30446;
wire ng33974;
wire ng33026;
wire ng30384;
wire ng34267;
wire ng34438;
wire ng33983;
wire ng25623;
wire ng28046;
wire ng24200;
wire ng30333;
wire ng33605;
wire ng33069;
wire ng30505;
wire ng34882;
wire ng30393;
wire ng30494;
wire ng26971;
wire ng25613;
wire ng30425;
wire ng32999;
wire ng30387;
wire ng33554;
wire ng25668;
wire ng33022;
wire ng34001;
wire ng25684;
wire ng24244;
wire ng33004;
wire ng25616;
wire ng34734;
wire ng30527;
wire ng31897;
wire ng30389;
wire ng24354;
wire ng30432;
wire ng31867;
wire ng30496;
wire ng34646;
wire ng33571;
wire ng25743;
wire ng30439;
wire ng34802;
wire ng29252;
wire ng24275;
wire ng33585;
wire ng30545;
wire ng30554;
wire ng33043;
wire ng24259;
wire ng33965;
wire ng25728;
wire ng30541;
wire ng30447;
wire ng31872;
wire ng30372;
wire ng24274;
wire ng26881;
wire ng25633;
wire ng34645;
wire ng30498;
wire ng30519;
wire ng29287;
wire ng33995;
wire ng20841;
wire ng21193;
wire ng20982;
wire ni24685;
wire ng19968;
wire ng20014;
wire ng19919;
wire ng21127;
wire ng21256;
wire ng19422;
wire ng19402;
wire ng19984;
wire ng26365;
wire ng17657;
wire ng17700;
wire ni31106;
wire ng30937;
wire ng31021;
wire ng31376;
wire ng30673;
wire ng30614;
wire ni31271;
wire ng30735;
wire ng28180;
wire ni31191;
wire ni31121;
wire ni31141;
wire ni30330;
wire ni31221;
wire ng31327;
wire ng17694;
wire ng17727;
wire ng31566;
wire ng31710;
wire ng34237;
wire ng33496;
wire ni31171;
wire ng31070;
wire ni31843;
wire ng34235;
wire ng25590;
wire ng26977;
wire ng18935;
wire ng27903;
wire ng22472;
wire ng26390;
wire ng24591;
wire ng13977;
wire ng29503;
wire ng29676;
wire ng30590;
wire ng8806;
wire ng10632;
wire ng23590;
wire ng27635;
wire ng28761;
wire ng27602;
wire ng11676;
wire ng31134;
wire ng23042;
wire ng25917;
wire ng14868;
wire ng10160;
wire ng23666;
wire ng10939;
wire ng13378;
wire ng13385;
wire ng11607;
wire ng30304;
wire ng25385;
wire ng23699;
wire ng30300;
wire ng22369;
wire ng27775;
wire ng15036;
wire ng12692;
wire ng20000;
wire ng25300;
wire ng12371;
wire ng24609;
wire ng14058;
wire ng14885;
wire ng20887;
wire ng12735;
wire ng30311;
wire ng17625;
wire ng12377;
wire ng31003;
wire ng28336;
wire ng16173;
wire ng28010;
wire ng13307;
wire ng15039;
wire ng14683;
wire ng25371;
wire ng14858;
wire ng11626;
wire ng11537;
wire ng7142;
wire ng14905;
wire ng10925;
wire ng24468;
wire ng26759;
wire ng34162;
wire ng10312;
wire ng12609;
wire ng12515;
wire ng8958;
wire ng11534;
wire ng10715;
wire ng13315;
wire ng12824;
wire ng14697;
wire ng28140;
wire ng27972;
wire ng22432;
wire ng12437;
wire ng25473;
wire ng10491;
wire ng14947;
wire ng17766;
wire ng17613;
wire ng17747;
wire ng17724;
wire ng17690;
wire ng24374;
wire ng20875;
wire ng23932;
wire ng31509;
wire ng12571;
wire ng14735;
wire ng9694;
wire ng26314;
wire ng27494;
wire ni18740;
wire ng10967;
wire ng12512;
wire ng12632;
wire ng14950;
wire ng26770;
wire ng17424;
wire ng11012;
wire ng11797;
wire ng11261;
wire ng10831;
wire ng29737;
wire ng11194;
wire ng11350;
wire ng13700;
wire ng13765;
wire ng24457;
wire ng26725;
wire ng12026;
wire ng14367;
wire ng11960;
wire ng11804;
wire ng11173;
wire ng21024;
wire ng11389;
wire ng13806;
wire ng29672;
wire ng14708;
wire ng17653;
wire ng24688;
wire ng30583;
wire ng11780;
wire ng22342;
wire ng25275;
wire ng10511;
wire ng10902;
wire ng16244;
wire ng16194;
wire ng17725;
wire ng16283;
wire ng16205;
wire ng12333;
wire ng25776;
wire ng31009;
wire ng22457;
wire ng25470;
wire ng13273;
wire ng10961;
wire ng16539;
wire ng16486;
wire ng25317;
wire ng11473;
wire ng13892;
wire ng10671;
wire ng13861;
wire ng12581;
wire ng11185;
wire ng14822;
wire ng25382;
wire ng14291;
wire ng17297;
wire ng8864;
wire ng11514;
wire ng11155;
wire ng11755;
wire ng20739;
wire ng10808;
wire ng13217;
wire ng24875;
wire ng12716;
wire ng8906;
wire ng11480;
wire ng15737;
wire ng25911;
wire ng34703;
wire ng8967;
wire ng14996;
wire ng29186;
wire ng22417;
wire ng10421;
wire ng14741;
wire ng12911;
wire ng13242;
wire ng27440;
wire ng17401;
wire ng10341;
wire ng14861;
wire ni18785;
wire ng12289;
wire ng21277;
wire ng10929;
wire ng14015;
wire ng14271;
wire ng22992;
wire ng28903;
wire ng14021;
wire ng12641;
wire ng12915;
wire ng28880;
wire ng23733;
wire ng29488;
wire ng25349;
wire ng10207;
wire ng11915;
wire ng27999;
wire ng14306;
wire ng8417;
wire ng16246;
wire ng23112;
wire ng14782;
wire ng23280;
wire ng29501;
wire ng30293;
wire ng28846;
wire ng14727;
wire ng14755;
wire ng19063;
wire ng15674;
wire ng25290;
wire ng13923;
wire ng16187;
wire ng28349;
wire ng29008;
wire ng12228;
wire ng10909;
wire ng13336;
wire ng27833;
wire ng12432;
wire ng14678;
wire ng32212;
wire ng22862;
wire ng14142;
wire ng8359;
wire ng8751;
wire ng11893;
wire ng15695;
wire ng19140;
wire ng25429;
wire ng25389;
wire ng7661;
wire ng10695;
wire ng14908;
wire ng24478;
wire ng26793;
wire ng29313;
wire ng12405;
wire ng14656;
wire ng25233;
wire ng27020;
wire ng28144;
wire ng13156;
wire ng25357;
wire ng12812;
wire ng14855;
wire ng11729;
wire ng13951;
wire ng10999;
wire ng24471;
wire ng31971;
wire ng13983;
wire ng11747;
wire ng14101;
wire ng25779;
wire ng10281;
wire ng14927;
wire ng12772;
wire ng14723;
wire ng23309;
wire ng14768;
wire ng29657;
wire ng28973;
wire ng23204;
wire ng7675;
wire ng7352;
wire ng14506;
wire ng11160;
wire ng21012;
wire ng11405;
wire ng14133;
wire ng23978;
wire ng27395;
wire ng28739;
wire ng22498;
wire ng12629;
wire ng25341;
wire ng27629;
wire ng14438;
wire ng11432;
wire ng30576;
wire ng12301;
wire ng27474;
wire ng27445;
wire ng17405;
wire ng10721;
wire ng23067;
wire ng12798;
wire ng14764;
wire ng24460;
wire ng26737;
wire ni17529;
wire ng12483;
wire ng9649;
wire ng11320;
wire ng26218;
wire ng11773;
wire ng11834;
wire ng11283;
wire ng11527;
wire ng13955;
wire ng14902;
wire ng24447;
wire ng26703;
wire ng13134;
wire ng26195;
wire ng11130;
wire ng34550;
wire ng13948;
wire ng25498;
wire ng25439;
wire ng13986;
wire ng12453;
wire ng14807;
wire ng28652;
wire ng13960;
wire ng11435;
wire ng14008;
wire ng27421;
wire ng17321;
wire ng12680;
wire ng15014;
wire ng25467;
wire ng25495;
wire ng25144;
wire ng23560;
wire ng27670;
wire ng30286;
wire ng25435;
wire ng10266;
wire ng12402;
wire ng13284;
wire ng14981;
wire ng20248;
wire ng17264;
wire ng14279;
wire ng13963;
wire ng12933;
wire ng14665;
wire ng26625;
wire ng31950;
wire ng11148;
wire ng10887;
wire ng14720;
wire ng7567;
wire ng30314;
wire ng29719;
wire ng26994;
wire ng23630;
wire ng13570;
wire ng10224;
wire ng14075;
wire ng14999;
wire ng8347;
wire ng10823;
wire ng12374;
wire ng22384;
wire ng25309;
wire ng25396;
wire ng14713;
wire ng20682;
wire ng28982;
wire ng14915;
wire ng11939;
wire ng28833;
wire ng7601;
wire ng15748;
wire ng11869;
wire ng14048;
wire ng12505;
wire ng10838;
wire ng14758;
wire ng13889;
wire ng12622;
wire ng10874;
wire ng24411;
wire ng26166;
wire ng13846;
wire ng14899;
wire ng12471;
wire ng14170;
wire ng8691;
wire ng23618;
wire ng14988;
wire ng10733;
wire ng10756;
wire ng15018;
wire ng28768;
wire ng11483;
wire ng10666;
wire ng10893;
wire ng14848;
wire ng11292;
wire ni27429;
wire ng25851;
wire ng29073;
wire ng28353;
wire ng25888;
wire ng23890;
wire ng13346;
wire ng9762;
wire ng28927;
wire ng15033;
wire ng12667;
wire ng20375;
wire ng26256;
wire ng26212;
wire ng24627;
wire ng14864;
wire ng31997;
wire ng11171;
wire ng30307;
wire ng28789;
wire ng8728;
wire ng20905;
wire ng20751;
wire ng29110;
wire ng33394;
wire ng25337;
wire ng13291;
wire ng13873;
wire ng13980;
wire ng25400;
wire ng23553;
wire ng23657;
wire ng29036;
wire ng25895;
wire ng25426;
wire ng13756;
wire ng27796;
wire ng29496;
wire ng11003;
wire ng10862;
wire ng11245;
wire ng25448;
wire ng14069;
wire ng14959;
wire ng12925;
wire ng25432;
wire ng11123;
wire ng12443;
wire ng14659;
wire ng27469;
wire ng28444;
wire ng29001;
wire ng29486;
wire ng11178;
wire ng11584;
wire ng13920;
wire ng14688;
wire ng12578;
wire ng11571;
wire ng25531;
wire ng10588;
wire ng31783;
wire ng11006;
wire ng13330;
wire ng14627;
wire ng14974;
wire ng14041;
wire ng27617;
wire ng28626;
wire ng14776;
wire ng13517;
wire ng11916;
wire ng14825;
wire ng23972;
wire ng14640;
wire ng23324;
wire ng16846;
wire ng14247;
wire ng12479;
wire ng10869;
wire ng14761;
wire ng28220;
wire ng23286;
wire ng14098;
wire ng27738;
wire ng7598;
wire ng13211;
wire ng22654;
wire ng26171;
wire ng15591;
wire ng14085;
wire ng28853;
wire ng11419;
wire ng11255;
wire ng14018;
wire ng11139;
wire ng14051;
wire ng24433;
wire ng26673;
wire ng14813;
wire ng11111;
wire ng12239;
wire ng12423;
wire ng9586;
wire ng15042;
wire ng12492;
wire ng14127;
wire ng7620;
wire ng14879;
wire ng28962;
wire ng14953;
wire ng27933;
wire ng27854;
wire ng11978;
wire ng29722;
wire ng14055;
wire ng14968;
wire ng11937;
wire ng13929;
wire ng30298;
wire ng14797;
wire ng28020;
wire ng29489;
wire ng14679;
wire ng9724;
wire ng27882;
wire ng10185;
wire ng13260;
wire ng8933;
wire ng23554;
wire ng10878;
wire ng15585;
wire ng27416;
wire ng26148;
wire ng26213;
wire ng11763;
wire ng23909;
wire ng7304;
wire ng14956;
wire ng29702;
wire ng13121;
wire ng12540;
wire ng25514;
wire ng14984;
wire ng14130;
wire ng14151;
wire ng14752;
wire ng25492;
wire ng8721;
wire ng28799;
wire ng28471;
wire ng28892;
wire ng23586;
wire ng14211;
wire ng29730;
wire ng24380;
wire ng10699;
wire ng10918;
wire ng14892;
wire ng11956;
wire ng25537;
wire ng12450;
wire ng8984;
wire ng14943;
wire ng17317;
wire ng12558;
wire ng13486;
wire ng28484;
wire ng10890;
wire ni30751;
wire ng14157;
wire ng14918;
wire ng14154;
wire ng13500;
wire ng14732;
wire ng10649;
wire ng17292;
wire ng16696;
wire ng14800;
wire ng11737;
wire ng9755;
wire ng14841;
wire ng14024;
wire ng22585;
wire ng12351;
wire ng11846;
wire ng16272;
wire ng28458;
wire ng11144;
wire ng14773;
wire ng14227;
wire ng23532;
wire ng10948;
wire ng14082;
wire ng14895;
wire ng14933;
wire ng23342;
wire ng24444;
wire ng26694;
wire ng11326;
wire ng10124;
wire ng11149;
wire ng13597;
wire ng13898;
wire ng14691;
wire ng29482;
wire ng14011;
wire ng23949;
wire ng14851;
wire ng13990;
wire ng26236;
wire ng23975;
wire ng13657;
wire ng14804;
wire ng12729;
wire ng14817;
wire ng14712;
wire ng13539;
wire ng13464;
wire ng28504;
wire ng29694;
wire ng28942;
wire ng28440;
wire ng14611;
wire ng9640;
wire ng8476;
wire ng15021;
wire ng30605;
wire ng15024;
wire ng29495;
wire ng14116;
wire ng14110;
wire ng9700;
wire ng16757;
wire ng17217;
wire ng14317;
wire ng14993;
wire ng13915;
wire ng15008;
wire ng14940;
wire ng16663;
wire ng25476;
wire ng33851;
wire ng21284;
wire ng14810;
wire ng29485;
wire ng14642;
wire ng34056;
wire ng34051;
wire ng34424;
wire ng16728;
wire ng9835;
wire ni30745;
wire ng12332;
wire wire3134;
wire wire3137;
wire wire3138;
wire wire3139;
wire wire3140;
wire wire3141;
wire wire3148;
wire wire3149;
wire wire3150;
wire wire3151;
wire wire3152;
wire wire3155;
wire wire3156;
wire wire3157;
wire wire3158;
wire wire3159;
wire wire3160;
wire wire3161;
wire wire3162;
wire wire3163;
wire wire3164;
wire wire3165;
wire wire3166;
wire wire3167;
wire wire3170;
wire wire3171;
wire wire3172;
wire wire3173;
wire wire3174;
wire wire3175;
wire wire3176;
wire wire3177;
wire wire3183;
wire wire3184;
wire wire3185;
wire wire3186;
wire wire3187;
wire wire3189;
wire wire3190;
wire wire3191;
wire wire3192;
wire wire3203;
wire wire3205;
wire wire3209;
wire wire3212;
wire wire3215;
wire wire3228;
wire wire3229;
wire wire3230;
wire wire3234;
wire wire3237;
wire wire3240;
wire wire3253;
wire wire3256;
wire wire3257;
wire wire3258;
wire wire3267;
wire wire3268;
wire wire3269;
wire wire3271;
wire wire3272;
wire wire3274;
wire wire3276;
wire wire3278;
wire wire3281;
wire wire3284;
wire wire3285;
wire wire3289;
wire wire3292;
wire wire3295;
wire wire3298;
wire wire3304;
wire wire3307;
wire wire3326;
wire wire3327;
wire wire3336;
wire wire3337;
wire wire3343;
wire wire3344;
wire wire3349;
wire wire3350;
wire wire3351;
wire wire3356;
wire wire3367;
wire wire3368;
wire wire3369;
wire wire3370;
wire wire3376;
wire wire3382;
wire wire3383;
wire wire3384;
wire wire3385;
wire wire3389;
wire wire3393;
wire wire3394;
wire wire3395;
wire wire3396;
wire wire3399;
wire wire3402;
wire wire3407;
wire wire3408;
wire wire3409;
wire wire3411;
wire wire3412;
wire wire3418;
wire wire3422;
wire wire3426;
wire wire3431;
wire wire3432;
wire wire3435;
wire wire3442;
wire wire3443;
wire wire3444;
wire wire3453;
wire wire3456;
wire wire3462;
wire wire3464;
wire wire3465;
wire wire3466;
wire wire3467;
wire wire3468;
wire wire3470;
wire wire3471;
wire wire3485;
wire wire3492;
wire wire3495;
wire wire3497;
wire wire3498;
wire wire3501;
wire wire3504;
wire wire3505;
wire wire3506;
wire wire3507;
wire wire3521;
wire wire3522;
wire wire3526;
wire wire3530;
wire wire3533;
wire wire3541;
wire wire3545;
wire wire3546;
wire wire3547;
wire wire3548;
wire wire3549;
wire wire3551;
wire wire3553;
wire wire3560;
wire wire3562;
wire wire3563;
wire wire3565;
wire wire3571;
wire wire3574;
wire wire3578;
wire wire3584;
wire wire3585;
wire wire3594;
wire wire3595;
wire wire3600;
wire wire3601;
wire wire3607;
wire wire3608;
wire wire3616;
wire wire3617;
wire wire3618;
wire wire3619;
wire wire3629;
wire wire3632;
wire wire3635;
wire wire3642;
wire wire3643;
wire wire3644;
wire wire3649;
wire wire3653;
wire wire3657;
wire wire3658;
wire wire3659;
wire wire3667;
wire wire3676;
wire wire3677;
wire wire3678;
wire wire3688;
wire wire3691;
wire wire3693;
wire wire3694;
wire wire3695;
wire wire3696;
wire wire3704;
wire wire3705;
wire wire3712;
wire wire3719;
wire wire3720;
wire wire3721;
wire wire3722;
wire wire3723;
wire wire3727;
wire wire3729;
wire wire3730;
wire wire3736;
wire wire3746;
wire wire3747;
wire wire3752;
wire wire3755;
wire wire3756;
wire wire3757;
wire wire3758;
wire wire3760;
wire wire3761;
wire wire3762;
wire wire3763;
wire wire3768;
wire wire3769;
wire wire3771;
wire wire3772;
wire wire3780;
wire wire3782;
wire wire3786;
wire wire3787;
wire wire3791;
wire wire3801;
wire wire3802;
wire wire3804;
wire wire3805;
wire wire3810;
wire wire3816;
wire wire3821;
wire wire3827;
wire wire3828;
wire wire3829;
wire wire3837;
wire wire3838;
wire wire3845;
wire wire3849;
wire wire3853;
wire wire3854;
wire wire3855;
wire wire3856;
wire wire3860;
wire wire3868;
wire wire3874;
wire wire3880;
wire wire3883;
wire wire3886;
wire wire3889;
wire wire3892;
wire wire3894;
wire wire3895;
wire wire3897;
wire wire3902;
wire wire3903;
wire wire3905;
wire wire3906;
wire wire3910;
wire wire3912;
wire wire3915;
wire wire3918;
wire wire3921;
wire wire3922;
wire wire3924;
wire wire3926;
wire wire3927;
wire wire3928;
wire wire3929;
wire wire3932;
wire wire3939;
wire wire3940;
wire wire3946;
wire wire3952;
wire wire3955;
wire wire3958;
wire wire3961;
wire wire3962;
wire wire3967;
wire wire3969;
wire wire3974;
wire wire3975;
wire wire3976;
wire wire3977;
wire wire3978;
wire wire3979;
wire wire3980;
wire wire3984;
wire wire3988;
wire wire3991;
wire wire3994;
wire wire3998;
wire wire4001;
wire wire4003;
wire wire4007;
wire wire4011;
wire wire4012;
wire wire4016;
wire wire4017;
wire wire4018;
wire wire4019;
wire wire4025;
wire wire4034;
wire wire4041;
wire wire4044;
wire wire4045;
wire wire4047;
wire wire4050;
wire wire4051;
wire wire4053;
wire wire4064;
wire wire4068;
wire wire4069;
wire wire4094;
wire wire4095;
wire wire4099;
wire wire4100;
wire wire4101;
wire wire4106;
wire wire4107;
wire wire4108;
wire wire4109;
wire wire4112;
wire wire4115;
wire wire4118;
wire wire4124;
wire wire4127;
wire wire4133;
wire wire4137;
wire wire4144;
wire wire4145;
wire wire4154;
wire wire4156;
wire wire4157;
wire wire4158;
wire wire4168;
wire wire4172;
wire wire4175;
wire wire4176;
wire wire4177;
wire wire4189;
wire wire4190;
wire wire4191;
wire wire4193;
wire wire4197;
wire wire4199;
wire wire4200;
wire wire4204;
wire wire4207;
wire wire4210;
wire wire4220;
wire wire4221;
wire wire4226;
wire wire4227;
wire wire4228;
wire wire4233;
wire wire4234;
wire wire4235;
wire wire4236;
wire wire4242;
wire wire4248;
wire wire4253;
wire wire4254;
wire wire4278;
wire wire4279;
wire wire4283;
wire wire4288;
wire wire4291;
wire wire4300;
wire wire4303;
wire wire4306;
wire wire4308;
wire wire4309;
wire wire4314;
wire wire4315;
wire wire4316;
wire wire4319;
wire wire4320;
wire wire4332;
wire wire4333;
wire wire4334;
wire wire4335;
wire wire4336;
wire wire4339;
wire wire4343;
wire wire4355;
wire wire4359;
wire wire4361;
wire wire4362;
wire wire4366;
wire wire4367;
wire wire4368;
wire wire4378;
wire wire4403;
wire wire4404;
wire wire4406;
wire wire4414;
wire wire4415;
wire wire4417;
wire wire4421;
wire wire4429;
wire wire4430;
wire wire4431;
wire wire4439;
wire wire4445;
wire wire4446;
wire wire4456;
wire wire4457;
wire wire4462;
wire wire4466;
wire wire4467;
wire wire4470;
wire wire4477;
wire wire4478;
wire wire4486;
wire wire4488;
wire wire4489;
wire wire4493;
wire wire4494;
wire wire4495;
wire wire4499;
wire wire4505;
wire wire4506;
wire wire4509;
wire wire4514;
wire wire4515;
wire wire4517;
wire wire4518;
wire wire4525;
wire wire4528;
wire wire4530;
wire wire4531;
wire wire4532;
wire wire4533;
wire wire4534;
wire wire4537;
wire wire4538;
wire wire4539;
wire wire4540;
wire wire4541;
wire wire4550;
wire wire4570;
wire wire4574;
wire wire4577;
wire wire4578;
wire wire4581;
wire wire4582;
wire wire4583;
wire wire4584;
wire wire4590;
wire wire4595;
wire wire4596;
wire wire4598;
wire wire4600;
wire wire4604;
wire wire4608;
wire wire4623;
wire wire4626;
wire wire4630;
wire wire4633;
wire wire4652;
wire wire4653;
wire wire4659;
wire wire4660;
wire wire4663;
wire wire4664;
wire wire4669;
wire wire4673;
wire wire4676;
wire wire4677;
wire wire4681;
wire wire4683;
wire wire4684;
wire wire4685;
wire wire4689;
wire wire4692;
wire wire4693;
wire wire4708;
wire wire4711;
wire wire4712;
wire wire4715;
wire wire4721;
wire wire4722;
wire wire4724;
wire wire4725;
wire wire4729;
wire wire4736;
wire wire4740;
wire wire4741;
wire wire4745;
wire wire4749;
wire wire4757;
wire wire4759;
wire wire4760;
wire wire4761;
wire wire4764;
wire wire4765;
wire wire4766;
wire wire4767;
wire wire4768;
wire wire4769;
wire wire4783;
wire wire4794;
wire wire4795;
wire wire4796;
wire wire4797;
wire wire4798;
wire wire4826;
wire wire4827;
wire wire4828;
wire wire4834;
wire wire4836;
wire wire4839;
wire wire4842;
wire wire4843;
wire wire4857;
wire wire4860;
wire wire4861;
wire wire4863;
wire wire4870;
wire wire4873;
wire wire4878;
wire wire4879;
wire wire4882;
wire wire4883;
wire wire4884;
wire wire4885;
wire wire4888;
wire wire4889;
wire wire4892;
wire wire4893;
wire wire4895;
wire wire4899;
wire wire4903;
wire wire4906;
wire wire4908;
wire wire4909;
wire wire4912;
wire wire4913;
wire wire4914;
wire wire4915;
wire wire4916;
wire wire4929;
wire wire4930;
wire wire4934;
wire wire4937;
wire wire4941;
wire wire4944;
wire wire4945;
wire wire4952;
wire wire4955;
wire wire4958;
wire wire4972;
wire wire4982;
wire wire4988;
wire wire4993;
wire wire4999;
wire wire5002;
wire wire5005;
wire wire5008;
wire wire5011;
wire wire5018;
wire wire5021;
wire wire5024;
wire wire5036;
wire wire5064;
wire wire5067;
wire wire5070;
wire wire5076;
wire wire5079;
wire wire5082;
wire wire5085;
wire wire5089;
wire wire5092;
wire wire5098;
wire wire5103;
wire wire5107;
wire wire5120;
wire wire5123;
wire wire5128;
wire wire5132;
wire wire5136;
wire wire5142;
wire wire5145;
wire wire5148;
wire wire5149;
wire wire5156;
wire wire5164;
wire wire5165;
wire wire5176;
wire wire5177;
wire wire5183;
wire wire5196;
wire wire5201;
wire wire5202;
wire wire5203;
wire wire5204;
wire wire5205;
wire wire5206;
wire wire5207;
wire wire5208;
wire wire5209;
wire wire5210;
wire wire5214;
wire wire5217;
wire wire5231;
wire wire5251;
wire wire5258;
wire wire5259;
wire wire5273;
wire wire5276;
wire wire5279;
wire wire5289;
wire wire5294;
wire wire5299;
wire wire5302;
wire wire5304;
wire wire5308;
wire wire5309;
wire wire5310;
wire wire5315;
wire wire5316;
wire wire5319;
wire wire5322;
wire wire5338;
wire wire5342;
wire wire5357;
wire wire5358;
wire wire5361;
wire wire5362;
wire wire5365;
wire wire5366;
wire wire5370;
wire wire5372;
wire wire5373;
wire wire5376;
wire wire5390;
wire wire5391;
wire wire5394;
wire wire5397;
wire wire5406;
wire wire5407;
wire wire5412;
wire wire5419;
wire wire5427;
wire wire5428;
wire wire5430;
wire wire5431;
wire wire5438;
wire wire5451;
wire wire5456;
wire wire5462;
wire wire5463;
wire wire5464;
wire wire5465;
wire wire5466;
wire wire5469;
wire wire5475;
wire wire5476;
wire wire5483;
wire wire5487;
wire wire5490;
wire wire5491;
wire wire5502;
wire wire5503;
wire wire5505;
wire wire5512;
wire wire5513;
wire wire5523;
wire wire5524;
wire wire5525;
wire wire5533;
wire wire5534;
wire wire5542;
wire wire5551;
wire wire5552;
wire wire5553;
wire wire5555;
wire wire5557;
wire wire5573;
wire wire5574;
wire wire5576;
wire wire5580;
wire wire5586;
wire wire5589;
wire wire5593;
wire wire5595;
wire wire5597;
wire wire5600;
wire wire5601;
wire wire5603;
wire wire5619;
wire wire5623;
wire wire5627;
wire wire5628;
wire wire5632;
wire wire5633;
wire wire5638;
wire wire5641;
wire wire5642;
wire wire5643;
wire wire5644;
wire wire5645;
wire wire5648;
wire wire5649;
wire wire5650;
wire wire5651;
wire wire5653;
wire wire5654;
wire wire5661;
wire wire5663;
wire wire5664;
wire wire5669;
wire wire5671;
wire wire5672;
wire wire5690;
wire wire5691;
wire wire5693;
wire wire5694;
wire wire5697;
wire wire5698;
wire wire5702;
wire wire5705;
wire wire5712;
wire wire5713;
wire wire5718;
wire wire5719;
wire wire5727;
wire wire5730;
wire wire5734;
wire wire5737;
wire wire5740;
wire wire5747;
wire wire5748;
wire wire5755;
wire wire5759;
wire wire5766;
wire wire5769;
wire wire5773;
wire wire5774;
wire wire5775;
wire wire5776;
wire wire5782;
wire wire5783;
wire wire5785;
wire wire5788;
wire wire5797;
wire wire5800;
wire wire5803;
wire wire5804;
wire wire5809;
wire wire5811;
wire wire5814;
wire wire5819;
wire wire5821;
wire wire5822;
wire wire5827;
wire wire5831;
wire wire5834;
wire wire5835;
wire wire5836;
wire wire5837;
wire wire5838;
wire wire5847;
wire wire5848;
wire wire5856;
wire wire5859;
wire wire5866;
wire wire5868;
wire wire5869;
wire wire5878;
wire wire5883;
wire wire5884;
wire wire5887;
wire wire5888;
wire wire5889;
wire wire5925;
wire wire5926;
wire wire5927;
wire wire5928;
wire wire5929;
wire wire5931;
wire wire5941;
wire wire5942;
wire wire5943;
wire wire5948;
wire wire5952;
wire wire5955;
wire wire5959;
wire wire5963;
wire wire5964;
wire wire5968;
wire wire5969;
wire wire5979;
wire wire5980;
wire wire5981;
wire wire5982;
wire wire6009;
wire wire6010;
wire wire6011;
wire wire6012;
wire wire6015;
wire wire6028;
wire wire6029;
wire wire6033;
wire wire6036;
wire wire6042;
wire wire6047;
wire wire6048;
wire wire6049;
wire wire6055;
wire wire6057;
wire wire6064;
wire wire6067;
wire wire6068;
wire wire6069;
wire wire6093;
wire wire6094;
wire wire6095;
wire wire6096;
wire wire6125;
wire wire6126;
wire wire6127;
wire wire6128;
wire wire6133;
wire wire6148;
wire wire6151;
wire wire6157;
wire wire6160;
wire wire6163;
wire wire6167;
wire wire6172;
wire wire6173;
wire wire6174;
wire wire6175;
wire wire6178;
wire wire6179;
wire wire6180;
wire wire6181;
wire wire6182;
wire wire6183;
wire wire6197;
wire wire6205;
wire wire6208;
wire wire6211;
wire wire6217;
wire wire6223;
wire wire6236;
wire wire6237;
wire wire6238;
wire wire6239;
wire wire6240;
wire wire6245;
wire wire6248;
wire wire6251;
wire wire6254;
wire wire6260;
wire wire6269;
wire wire6270;
wire wire6271;
wire wire6273;
wire wire6274;
wire wire6276;
wire wire6277;
wire wire6278;
wire wire6281;
wire wire6282;
wire wire6283;
wire wire6293;
wire wire6294;
wire wire6295;
wire wire6300;
wire wire6301;
wire wire6302;
wire wire6304;
wire wire6305;
wire wire6306;
wire wire6307;
wire wire6317;
wire wire6319;
wire wire6323;
wire wire6324;
wire wire6325;
wire wire6329;
wire wire6330;
wire wire6331;
wire wire6332;
wire wire6333;
wire wire6335;
wire wire6336;
wire wire6341;
wire wire6348;
wire wire6361;
wire wire6362;
wire wire6363;
wire wire6364;
wire wire6368;
wire wire6373;
wire wire6389;
wire wire6390;
wire wire6395;
wire wire6396;
wire wire6398;
wire wire6407;
wire wire6408;
wire wire6415;
wire wire6421;
wire wire6424;
wire wire6436;
wire wire6442;
wire wire6443;
wire wire6450;
wire wire6451;
wire wire6474;
wire wire6475;
wire wire6476;
wire wire6482;
wire wire6486;
wire wire6491;
wire wire6494;
wire wire6500;
wire wire6503;
wire wire6504;
wire wire6514;
wire wire6515;
wire wire6516;
wire wire6520;
wire wire6524;
wire wire6527;
wire wire6532;
wire wire6539;
wire wire6542;
wire wire6544;
wire wire6545;
wire wire6548;
wire wire6549;
wire wire6552;
wire wire6553;
wire wire6561;
wire wire6565;
wire wire6571;
wire wire6572;
wire wire6576;
wire wire6588;
wire wire6592;
wire wire6595;
wire wire6598;
wire wire6604;
wire wire6612;
wire wire6614;
wire wire6615;
wire wire6619;
wire wire6620;
wire wire6622;
wire wire6653;
wire wire6655;
wire wire6660;
wire wire6663;
wire wire6665;
wire wire6666;
wire wire6669;
wire wire6674;
wire wire6675;
wire wire6678;
wire wire6686;
wire wire6687;
wire wire6690;
wire wire6691;
wire wire6694;
wire wire6695;
wire wire6696;
wire wire6697;
wire wire6698;
wire wire6699;
wire wire6700;
wire wire6701;
wire wire6702;
wire wire6703;
wire wire6704;
wire wire6705;
wire wire6706;
wire wire6709;
wire wire6714;
wire wire6715;
wire wire6716;
wire wire6743;
wire wire6763;
wire wire6764;
wire wire6770;
wire wire6777;
wire wire6781;
wire wire6784;
wire wire6789;
wire wire6790;
wire wire6804;
wire wire6805;
wire wire6808;
wire wire6809;
wire wire6816;
wire wire6817;
wire wire6823;
wire wire6825;
wire wire6826;
wire wire6827;
wire wire6828;
wire wire6829;
wire wire6832;
wire wire6833;
wire wire6838;
wire wire6842;
wire wire6843;
wire wire6844;
wire wire6847;
wire wire6849;
wire wire6852;
wire wire6872;
wire wire6890;
wire wire6899;
wire wire6904;
wire wire6905;
wire wire6906;
wire wire6912;
wire wire6915;
wire wire6916;
wire wire6925;
wire wire6933;
wire wire6946;
wire wire6947;
wire wire6948;
wire wire6949;
wire wire6950;
wire wire6951;
wire wire6952;
wire wire6953;
wire wire6956;
wire wire6959;
wire wire6960;
wire wire6965;
wire wire6966;
wire wire6967;
wire wire6985;
wire wire6988;
wire wire6992;
wire wire7004;
wire wire7005;
wire wire7006;
wire wire7007;
wire wire7008;
wire wire7009;
wire wire7010;
wire wire7011;
wire wire7024;
wire wire7028;
wire wire7030;
wire wire7034;
wire wire7041;
wire wire7046;
wire wire7047;
wire wire7049;
wire wire7050;
wire wire7058;
wire wire7059;
wire wire7065;
wire wire7069;
wire wire7077;
wire wire7078;
wire wire7083;
wire wire7096;
wire wire7097;
wire wire7100;
wire wire7102;
wire wire7114;
wire wire7116;
wire wire7117;
wire wire7126;
wire wire7131;
wire wire7132;
wire wire7133;
wire wire7134;
wire wire7137;
wire wire7138;
wire wire7167;
wire wire7170;
wire wire7175;
wire wire7180;
wire wire7181;
wire wire7186;
wire wire7187;
wire wire7190;
wire wire7193;
wire wire7199;
wire wire7200;
wire wire7201;
wire wire7202;
wire wire7204;
wire wire7205;
wire wire7221;
wire wire7225;
wire wire7232;
wire wire7233;
wire wire7236;
wire wire7237;
wire wire7248;
wire wire7249;
wire wire7255;
wire wire7257;
wire wire7259;
wire wire7260;
wire wire7269;
wire wire7283;
wire wire7284;
wire wire7286;
wire wire7287;
wire wire7291;
wire wire7298;
wire wire7299;
wire wire7300;
wire wire7301;
wire wire7306;
wire wire7308;
wire wire7309;
wire wire7310;
wire wire7321;
wire wire7322;
wire wire7323;
wire wire7324;
wire wire7325;
wire wire7326;
wire wire7331;
wire wire7332;
wire wire7346;
wire wire7351;
wire wire7352;
wire wire7371;
wire wire7372;
wire wire7373;
wire wire7374;
wire wire7375;
wire wire7376;
wire wire7377;
wire wire7378;
wire wire7382;
wire wire7390;
wire wire7391;
wire wire7392;
wire wire7398;
wire wire7399;
wire wire7400;
wire wire7409;
wire wire7410;
wire wire7411;
wire wire7412;
wire wire7414;
wire wire7424;
wire wire7426;
wire wire7436;
wire wire7437;
wire wire7438;
wire wire7445;
wire wire7446;
wire wire7447;
wire wire7452;
wire wire7462;
wire wire7463;
wire wire7464;
wire wire7466;
wire wire7467;
wire wire7468;
wire wire7469;
wire wire7470;
wire wire7471;
wire wire7472;
wire wire7473;
wire wire7474;
wire wire7475;
wire wire7485;
wire wire7486;
wire wire7487;
wire wire7489;
wire wire7490;
wire wire7491;
wire wire7492;
wire wire7493;
wire wire7494;
wire wire7495;
wire wire7498;
wire wire7499;
wire wire7500;
wire wire7501;
wire wire7502;
wire wire7503;
wire wire7504;
wire wire7505;
wire wire7506;
wire wire7507;
wire wire7509;
wire wire7518;
wire wire7521;
wire wire7531;
wire wire7532;
wire wire7533;
wire wire7540;
wire wire7541;
wire wire7542;
wire wire7543;
wire wire7544;
wire wire7545;
wire wire7546;
wire wire7547;
wire wire7559;
wire wire7565;
wire wire7567;
wire wire7568;
wire wire7581;
wire wire7582;
wire wire7583;
wire wire7595;
wire wire7596;
wire wire7606;
wire wire7608;
wire wire7609;
wire wire7623;
wire wire7624;
wire wire7625;
wire wire7634;
wire wire7639;
wire wire7640;
wire wire7641;
wire wire7642;
wire wire7643;
wire wire7644;
wire wire7645;
wire wire7646;
wire wire7647;
wire wire7649;
wire wire7650;
wire wire7652;
wire wire7662;
wire wire7663;
wire wire7664;
wire wire7665;
wire wire7666;
wire wire7667;
wire wire7668;
wire wire7671;
wire wire7677;
wire wire7681;
wire wire7685;
wire wire7686;
wire wire7690;
wire wire7691;
wire wire7692;
wire wire7693;
wire wire7694;
wire wire7695;
wire wire7703;
wire wire7709;
wire wire7720;
wire wire7721;
wire wire7725;
wire wire7734;
wire wire7735;
wire wire28470;
wire wire28473;
wire wire28475;
wire wire28476;
wire wire28478;
wire wire28482;
wire wire28483;
wire wire28484;
wire wire28485;
wire wire28488;
wire wire28490;
wire wire28491;
wire wire28503;
wire wire28505;
wire wire28507;
wire wire28514;
wire wire28515;
wire wire28519;
wire wire28521;
wire wire28522;
wire wire28525;
wire wire28526;
wire wire28530;
wire wire28532;
wire wire28534;
wire wire28536;
wire wire28538;
wire wire28540;
wire wire28543;
wire wire28544;
wire wire28548;
wire wire28549;
wire wire28551;
wire wire28555;
wire wire28556;
wire wire28558;
wire wire28561;
wire wire28562;
wire wire28563;
wire wire28567;
wire wire28568;
wire wire28569;
wire wire28571;
wire wire28572;
wire wire28573;
wire wire28574;
wire wire28575;
wire wire28577;
wire wire28581;
wire wire28583;
wire wire28584;
wire wire28587;
wire wire28588;
wire wire28606;
wire wire28607;
wire wire28609;
wire wire28611;
wire wire28612;
wire wire28614;
wire wire28617;
wire wire28622;
wire wire28625;
wire wire28629;
wire wire28632;
wire wire28637;
wire wire28638;
wire wire28640;
wire wire28643;
wire wire28645;
wire wire28646;
wire wire28651;
wire wire28655;
wire wire28657;
wire wire28659;
wire wire28661;
wire wire28670;
wire wire28673;
wire wire28687;
wire wire28689;
wire wire28694;
wire wire28706;
wire wire28707;
wire wire28708;
wire wire28711;
wire wire28712;
wire wire28713;
wire wire28715;
wire wire28716;
wire wire28718;
wire wire28719;
wire wire28720;
wire wire28722;
wire wire28723;
wire wire28731;
wire wire28732;
wire wire28733;
wire wire28734;
wire wire28741;
wire wire28742;
wire wire28743;
wire wire28746;
wire wire28747;
wire wire28751;
wire wire28754;
wire wire28757;
wire wire28758;
wire wire28765;
wire wire28766;
wire wire28769;
wire wire28770;
wire wire28775;
wire wire28776;
wire wire28779;
wire wire28783;
wire wire28786;
wire wire28787;
wire wire28788;
wire wire28792;
wire wire28793;
wire wire28794;
wire wire28795;
wire wire28796;
wire wire28798;
wire wire28799;
wire wire28800;
wire wire28801;
wire wire28802;
wire wire28803;
wire wire28804;
wire wire28806;
wire wire28807;
wire wire28809;
wire wire28810;
wire wire28811;
wire wire28812;
wire wire28813;
wire wire28814;
wire wire28815;
wire wire28816;
wire wire28818;
wire wire28819;
wire wire28820;
wire wire28821;
wire wire28822;
wire wire28823;
wire wire28824;
wire wire28827;
wire wire28829;
wire wire28830;
wire wire28831;
wire wire28834;
wire wire28836;
wire wire28837;
wire wire28841;
wire wire28843;
wire wire28848;
wire wire28849;
wire wire28850;
wire wire28853;
wire wire28854;
wire wire28856;
wire wire28858;
wire wire28860;
wire wire28861;
wire wire28862;
wire wire28863;
wire wire28864;
wire wire28865;
wire wire28866;
wire wire28867;
wire wire28874;
wire wire28878;
wire wire28881;
wire wire28883;
wire wire28884;
wire wire28885;
wire wire28886;
wire wire28887;
wire wire28891;
wire wire28892;
wire wire28896;
wire wire28898;
wire wire28903;
wire wire28905;
wire wire28907;
wire wire28915;
wire wire28916;
wire wire28919;
wire wire28920;
wire wire28921;
wire wire28924;
wire wire28925;
wire wire28927;
wire wire28928;
wire wire28931;
wire wire28932;
wire wire28933;
wire wire28935;
wire wire28937;
wire wire28938;
wire wire28940;
wire wire28941;
wire wire28942;
wire wire28943;
wire wire28944;
wire wire28945;
wire wire28946;
wire wire28947;
wire wire28949;
wire wire28952;
wire wire28953;
wire wire28954;
wire wire28955;
wire wire28956;
wire wire28958;
wire wire28959;
wire wire28961;
wire wire28963;
wire wire28964;
wire wire28965;
wire wire28966;
wire wire28967;
wire wire28968;
wire wire28971;
wire wire28972;
wire wire28973;
wire wire28975;
wire wire28978;
wire wire28979;
wire wire28980;
wire wire28982;
wire wire28983;
wire wire28984;
wire wire28986;
wire wire28987;
wire wire28988;
wire wire28989;
wire wire28990;
wire wire28991;
wire wire28992;
wire wire28995;
wire wire28996;
wire wire29000;
wire wire29002;
wire wire29003;
wire wire29009;
wire wire29011;
wire wire29012;
wire wire29013;
wire wire29015;
wire wire29016;
wire wire29023;
wire wire29025;
wire wire29026;
wire wire29027;
wire wire29028;
wire wire29029;
wire wire29030;
wire wire29039;
wire wire29040;
wire wire29043;
wire wire29044;
wire wire29047;
wire wire29048;
wire wire29049;
wire wire29050;
wire wire29051;
wire wire29054;
wire wire29055;
wire wire29058;
wire wire29061;
wire wire29063;
wire wire29068;
wire wire29070;
wire wire29071;
wire wire29072;
wire wire29073;
wire wire29076;
wire wire29077;
wire wire29081;
wire wire29084;
wire wire29087;
wire wire29088;
wire wire29091;
wire wire29097;
wire wire29099;
wire wire29103;
wire wire29104;
wire wire29105;
wire wire29106;
wire wire29107;
wire wire29108;
wire wire29111;
wire wire29113;
wire wire29115;
wire wire29117;
wire wire29119;
wire wire29120;
wire wire29121;
wire wire29124;
wire wire29126;
wire wire29128;
wire wire29129;
wire wire29130;
wire wire29131;
wire wire29138;
wire wire29143;
wire wire29148;
wire wire29153;
wire wire29159;
wire wire29161;
wire wire29162;
wire wire29168;
wire wire29171;
wire wire29175;
wire wire29178;
wire wire29180;
wire wire29183;
wire wire29184;
wire wire29185;
wire wire29186;
wire wire29192;
wire wire29195;
wire wire29196;
wire wire29198;
wire wire29199;
wire wire29202;
wire wire29209;
wire wire29210;
wire wire29216;
wire wire29220;
wire wire29221;
wire wire29223;
wire wire29224;
wire wire29225;
wire wire29227;
wire wire29228;
wire wire29232;
wire wire29233;
wire wire29234;
wire wire29235;
wire wire29236;
wire wire29237;
wire wire29238;
wire wire29239;
wire wire29240;
wire wire29245;
wire wire29246;
wire wire29247;
wire wire29248;
wire wire29250;
wire wire29251;
wire wire29253;
wire wire29254;
wire wire29255;
wire wire29256;
wire wire29257;
wire wire29258;
wire wire29259;
wire wire29260;
wire wire29263;
wire wire29265;
wire wire29266;
wire wire29269;
wire wire29272;
wire wire29277;
wire wire29278;
wire wire29280;
wire wire29281;
wire wire29283;
wire wire29284;
wire wire29285;
wire wire29290;
wire wire29292;
wire wire29293;
wire wire29300;
wire wire29303;
wire wire29304;
wire wire29305;
wire wire29308;
wire wire29309;
wire wire29312;
wire wire29313;
wire wire29315;
wire wire29316;
wire wire29317;
wire wire29320;
wire wire29322;
wire wire29323;
wire wire29324;
wire wire29325;
wire wire29326;
wire wire29328;
wire wire29329;
wire wire29330;
wire wire29335;
wire wire29336;
wire wire29340;
wire wire29346;
wire wire29348;
wire wire29350;
wire wire29352;
wire wire29355;
wire wire29359;
wire wire29361;
wire wire29362;
wire wire29363;
wire wire29366;
wire wire29367;
wire wire29371;
wire wire29374;
wire wire29377;
wire wire29378;
wire wire29383;
wire wire29391;
wire wire29393;
wire wire29397;
wire wire29402;
wire wire29403;
wire wire29405;
wire wire29408;
wire wire29414;
wire wire29415;
wire wire29416;
wire wire29417;
wire wire29418;
wire wire29419;
wire wire29420;
wire wire29422;
wire wire29423;
wire wire29424;
wire wire29425;
wire wire29426;
wire wire29428;
wire wire29429;
wire wire29430;
wire wire29431;
wire wire29432;
wire wire29433;
wire wire29434;
wire wire29436;
wire wire29437;
wire wire29438;
wire wire29439;
wire wire29440;
wire wire29441;
wire wire29442;
wire wire29443;
wire wire29444;
wire wire29445;
wire wire29446;
wire wire29447;
wire wire29448;
wire wire29451;
wire wire29452;
wire wire29453;
wire wire29454;
wire wire29456;
wire wire29457;
wire wire29458;
wire wire29459;
wire wire29460;
wire wire29461;
wire wire29462;
wire wire29464;
wire wire29466;
wire wire29467;
wire wire29468;
wire wire29469;
wire wire29470;
wire wire29471;
wire wire29472;
wire wire29475;
wire wire29476;
wire wire29477;
wire wire29480;
wire wire29481;
wire wire29482;
wire wire29484;
wire wire29486;
wire wire29489;
wire wire29491;
wire wire29493;
wire wire29495;
wire wire29496;
wire wire29497;
wire wire29499;
wire wire29500;
wire wire29502;
wire wire29507;
wire wire29508;
wire wire29510;
wire wire29511;
wire wire29512;
wire wire29516;
wire wire29517;
wire wire29518;
wire wire29520;
wire wire29521;
wire wire29522;
wire wire29523;
wire wire29524;
wire wire29526;
wire wire29527;
wire wire29532;
wire wire29534;
wire wire29535;
wire wire29536;
wire wire29537;
wire wire29538;
wire wire29539;
wire wire29541;
wire wire29542;
wire wire29545;
wire wire29546;
wire wire29548;
wire wire29549;
wire wire29550;
wire wire29551;
wire wire29553;
wire wire29555;
wire wire29556;
wire wire29557;
wire wire29559;
wire wire29560;
wire wire29561;
wire wire29563;
wire wire29564;
wire wire29567;
wire wire29568;
wire wire29571;
wire wire29573;
wire wire29575;
wire wire29577;
wire wire29579;
wire wire29581;
wire wire29582;
wire wire29583;
wire wire29584;
wire wire29585;
wire wire29586;
wire wire29587;
wire wire29589;
wire wire29590;
wire wire29591;
wire wire29592;
wire wire29593;
wire wire29595;
wire wire29596;
wire wire29597;
wire wire29598;
wire wire29599;
wire wire29601;
wire wire29602;
wire wire29604;
wire wire29606;
wire wire29607;
wire wire29608;
wire wire29609;
wire wire29610;
wire wire29611;
wire wire29614;
wire wire29615;
wire wire29617;
wire wire29618;
wire wire29619;
wire wire29620;
wire wire29621;
wire wire29623;
wire wire29624;
wire wire29625;
wire wire29626;
wire wire29627;
wire wire29629;
wire wire29630;
wire wire29631;
wire wire29632;
wire wire29633;
wire wire29634;
wire wire29635;
wire wire29638;
wire wire29639;
wire wire29640;
wire wire29641;
wire wire29642;
wire wire29643;
wire wire29644;
wire wire29646;
wire wire29647;
wire wire29648;
wire wire29652;
wire wire29653;
wire wire29657;
wire wire29658;
wire wire29663;
wire wire29665;
wire wire29669;
wire wire29670;
wire wire29671;
wire wire29672;
wire wire29674;
wire wire29675;
wire wire29676;
wire wire29679;
wire wire29683;
wire wire29688;
wire wire29689;
wire wire29693;
wire wire29694;
wire wire29702;
wire wire29703;
wire wire29706;
wire wire29708;
wire wire29709;
wire wire29711;
wire wire29712;
wire wire29714;
wire wire29715;
wire wire29716;
wire wire29718;
wire wire29720;
wire wire29721;
wire wire29723;
wire wire29724;
wire wire29725;
wire wire29727;
wire wire29728;
wire wire29730;
wire wire29731;
wire wire29733;
wire wire29735;
wire wire29737;
wire wire29738;
wire wire29742;
wire wire29743;
wire wire29747;
wire wire29749;
wire wire29752;
wire wire29753;
wire wire29755;
wire wire29757;
wire wire29758;
wire wire29761;
wire wire29762;
wire wire29764;
wire wire29770;
wire wire29771;
wire wire29775;
wire wire29776;
wire wire29780;
wire wire29785;
wire wire29787;
wire wire29789;
wire wire29791;
wire wire29792;
wire wire29797;
wire wire29798;
wire wire29800;
wire wire29801;
wire wire29804;
wire wire29805;
wire wire29806;
wire wire29807;
wire wire29809;
wire wire29810;
wire wire29811;
wire wire29812;
wire wire29816;
wire wire29820;
wire wire29824;
wire wire29827;
wire wire29828;
wire wire29830;
wire wire29831;
wire wire29834;
wire wire29835;
wire wire29836;
wire wire29841;
wire wire29843;
wire wire29848;
wire wire29849;
wire wire29850;
wire wire29851;
wire wire29852;
wire wire29853;
wire wire29855;
wire wire29856;
wire wire29858;
wire wire29859;
wire wire29862;
wire wire29863;
wire wire29867;
wire wire29870;
wire wire29873;
wire wire29874;
wire wire29883;
wire wire29884;
wire wire29885;
wire wire29887;
wire wire29888;
wire wire29889;
wire wire29890;
wire wire29894;
wire wire29899;
wire wire29900;
wire wire29901;
wire wire29902;
wire wire29903;
wire wire29904;
wire wire29905;
wire wire29907;
wire wire29908;
wire wire29912;
wire wire29914;
wire wire29917;
wire wire29918;
wire wire29919;
wire wire29920;
wire wire29921;
wire wire29922;
wire wire29923;
wire wire29925;
wire wire29926;
wire wire29928;
wire wire29930;
wire wire29932;
wire wire29934;
wire wire29936;
wire wire29937;
wire wire29939;
wire wire29941;
wire wire29942;
wire wire29944;
wire wire29946;
wire wire29948;
wire wire29949;
wire wire29950;
wire wire29952;
wire wire29953;
wire wire29954;
wire wire29955;
wire wire29956;
wire wire29957;
wire wire29959;
wire wire29961;
wire wire29962;
wire wire29963;
wire wire29965;
wire wire29966;
wire wire29968;
wire wire29971;
wire wire29972;
wire wire29974;
wire wire29976;
wire wire29978;
wire wire29980;
wire wire29982;
wire wire29984;
wire wire29985;
wire wire29986;
wire wire29987;
wire wire29988;
wire wire29989;
wire wire29990;
wire wire29991;
wire wire29992;
wire wire29993;
wire wire29994;
wire wire29996;
wire wire29997;
wire wire29999;
wire wire30000;
wire wire30002;
wire wire30003;
wire wire30004;
wire wire30006;
wire wire30008;
wire wire30009;
wire wire30010;
wire wire30011;
wire wire30013;
wire wire30014;
wire wire30016;
wire wire30017;
wire wire30018;
wire wire30019;
wire wire30020;
wire wire30021;
wire wire30022;
wire wire30023;
wire wire30024;
wire wire30025;
wire wire30026;
wire wire30028;
wire wire30029;
wire wire30030;
wire wire30031;
wire wire30033;
wire wire30034;
wire wire30035;
wire wire30036;
wire wire30037;
wire wire30038;
wire wire30039;
wire wire30041;
wire wire30042;
wire wire30044;
wire wire30045;
wire wire30048;
wire wire30052;
wire wire30053;
wire wire30055;
wire wire30056;
wire wire30057;
wire wire30059;
wire wire30061;
wire wire30062;
wire wire30063;
wire wire30064;
wire wire30065;
wire wire30066;
wire wire30067;
wire wire30068;
wire wire30069;
wire wire30070;
wire wire30071;
wire wire30072;
wire wire30074;
wire wire30076;
wire wire30077;
wire wire30078;
wire wire30079;
wire wire30081;
wire wire30082;
wire wire30084;
wire wire30085;
wire wire30086;
wire wire30087;
wire wire30088;
wire wire30089;
wire wire30091;
wire wire30095;
wire wire30096;
wire wire30097;
wire wire30098;
wire wire30099;
wire wire30100;
wire wire30101;
wire wire30102;
wire wire30103;
wire wire30104;
wire wire30105;
wire wire30106;
wire wire30108;
wire wire30110;
wire wire30111;
wire wire30112;
wire wire30113;
wire wire30115;
wire wire30116;
wire wire30118;
wire wire30119;
wire wire30120;
wire wire30121;
wire wire30122;
wire wire30123;
wire wire30124;
wire wire30125;
wire wire30126;
wire wire30127;
wire wire30128;
wire wire30130;
wire wire30131;
wire wire30132;
wire wire30133;
wire wire30135;
wire wire30136;
wire wire30137;
wire wire30138;
wire wire30139;
wire wire30140;
wire wire30141;
wire wire30144;
wire wire30146;
wire wire30147;
wire wire30148;
wire wire30150;
wire wire30151;
wire wire30152;
wire wire30153;
wire wire30154;
wire wire30155;
wire wire30157;
wire wire30158;
wire wire30159;
wire wire30160;
wire wire30162;
wire wire30163;
wire wire30164;
wire wire30165;
wire wire30166;
wire wire30167;
wire wire30168;
wire wire30169;
wire wire30170;
wire wire30171;
wire wire30173;
wire wire30175;
wire wire30176;
wire wire30177;
wire wire30178;
wire wire30180;
wire wire30181;
wire wire30182;
wire wire30183;
wire wire30184;
wire wire30185;
wire wire30186;
wire wire30187;
wire wire30188;
wire wire30189;
wire wire30190;
wire wire30193;
wire wire30194;
wire wire30195;
wire wire30199;
wire wire30201;
wire wire30202;
wire wire30203;
wire wire30204;
wire wire30205;
wire wire30208;
wire wire30209;
wire wire30210;
wire wire30211;
wire wire30213;
wire wire30215;
wire wire30216;
wire wire30217;
wire wire30218;
wire wire30219;
wire wire30220;
wire wire30221;
wire wire30222;
wire wire30223;
wire wire30224;
wire wire30226;
wire wire30228;
wire wire30229;
wire wire30230;
wire wire30231;
wire wire30232;
wire wire30236;
wire wire30237;
wire wire30238;
wire wire30241;
wire wire30245;
wire wire30249;
wire wire30250;
wire wire30251;
wire wire30254;
wire wire30255;
wire wire30257;
wire wire30258;
wire wire30260;
wire wire30261;
wire wire30263;
wire wire30264;
wire wire30265;
wire wire30267;
wire wire30268;
wire wire30269;
wire wire30272;
wire wire30273;
wire wire30274;
wire wire30276;
wire wire30281;
wire wire30283;
wire wire30286;
wire wire30293;
wire wire30295;
wire wire30300;
wire wire30301;
wire wire30304;
wire wire30307;
wire wire30310;
wire wire30312;
wire wire30313;
wire wire30314;
wire wire30315;
wire wire30316;
wire wire30320;
wire wire30321;
wire wire30324;
wire wire30325;
wire wire30327;
wire wire30328;
wire wire30329;
wire wire30330;
wire wire30331;
wire wire30332;
wire wire30334;
wire wire30335;
wire wire30337;
wire wire30339;
wire wire30341;
wire wire30342;
wire wire30343;
wire wire30344;
wire wire30348;
wire wire30349;
wire wire30356;
wire wire30359;
wire wire30361;
wire wire30362;
wire wire30365;
wire wire30367;
wire wire30369;
wire wire30372;
wire wire30373;
wire wire30375;
wire wire30377;
wire wire30382;
wire wire30383;
wire wire30384;
wire wire30386;
wire wire30388;
wire wire30390;
wire wire30391;
wire wire30392;
wire wire30394;
wire wire30395;
wire wire30399;
wire wire30402;
wire wire30404;
wire wire30405;
wire wire30406;
wire wire30407;
wire wire30411;
wire wire30412;
wire wire30417;
wire wire30420;
wire wire30421;
wire wire30422;
wire wire30427;
wire wire30428;
wire wire30430;
wire wire30431;
wire wire30433;
wire wire30434;
wire wire30436;
wire wire30437;
wire wire30441;
wire wire30443;
wire wire30444;
wire wire30447;
wire wire30448;
wire wire30453;
wire wire30457;
wire wire30458;
wire wire30464;
wire wire30465;
wire wire30466;
wire wire30467;
wire wire30471;
wire wire30472;
wire wire30474;
wire wire30475;
wire wire30477;
wire wire30478;
wire wire30480;
wire wire30484;
wire wire30487;
wire wire30488;
wire wire30497;
wire wire30498;
wire wire30499;
wire wire30505;
wire wire30506;
wire wire30512;
wire wire30513;
wire wire30515;
wire wire30516;
wire wire30517;
wire wire30518;
wire wire30521;
wire wire30523;
wire wire30527;
wire wire30529;
wire wire30534;
wire wire30535;
wire wire30539;
wire wire30547;
wire wire30550;
wire wire30551;
wire wire30552;
wire wire30555;
wire wire30557;
wire wire30562;
wire wire30564;
wire wire30566;
wire wire30567;
wire wire30568;
wire wire30570;
wire wire30572;
wire wire30573;
wire wire30574;
wire wire30575;
wire wire30576;
wire wire30578;
wire wire30581;
wire wire30583;
wire wire30585;
wire wire30586;
wire wire30592;
wire wire30593;
wire wire30595;
wire wire30596;
wire wire30598;
wire wire30599;
wire wire30601;
wire wire30602;
wire wire30604;
wire wire30605;
wire wire30607;
wire wire30608;
wire wire30609;
wire wire30611;
wire wire30612;
wire wire30613;
wire wire30616;
wire wire30619;
wire wire30621;
wire wire30622;
wire wire30628;
wire wire30629;
wire wire30630;
wire wire30631;
wire wire30632;
wire wire30634;
wire wire30635;
wire wire30636;
wire wire30637;
wire wire30638;
wire wire30639;
wire wire30640;
wire wire30642;
wire wire30643;
wire wire30644;
wire wire30645;
wire wire30646;
wire wire30647;
wire wire30648;
wire wire30649;
wire wire30650;
wire wire30651;
wire wire30652;
wire wire30653;
wire wire30654;
wire wire30655;
wire wire30656;
wire wire30659;
wire wire30660;
wire wire30661;
wire wire30662;
wire wire30663;
wire wire30664;
wire wire30665;
wire wire30666;
wire wire30668;
wire wire30670;
wire wire30671;
wire wire30672;
wire wire30674;
wire wire30675;
wire wire30676;
wire wire30677;
wire wire30678;
wire wire30679;
wire wire30680;
wire wire30683;
wire wire30685;
wire wire30687;
wire wire30688;
wire wire30692;
wire wire30694;
wire wire30695;
wire wire30696;
wire wire30697;
wire wire30698;
wire wire30699;
wire wire30702;
wire wire30703;
wire wire30704;
wire wire30705;
wire wire30708;
wire wire30709;
wire wire30710;
wire wire30712;
wire wire30713;
wire wire30716;
wire wire30717;
wire wire30719;
wire wire30720;
wire wire30722;
wire wire30723;
wire wire30725;
wire wire30726;
wire wire30728;
wire wire30729;
wire wire30730;
wire wire30731;
wire wire30733;
wire wire30734;
wire wire30735;
wire wire30737;
wire wire30740;
wire wire30742;
wire wire30743;
wire wire30746;
wire wire30748;
wire wire30750;
wire wire30752;
wire wire30754;
wire wire30759;
wire wire30760;
wire wire30763;
wire wire30765;
wire wire30768;
wire wire30769;
wire wire30770;
wire wire30776;
wire wire30782;
wire wire30783;
wire wire30788;
wire wire30789;
wire wire30794;
wire wire30795;
wire wire30800;
wire wire30801;
wire wire30802;
wire wire30803;
wire wire30805;
wire wire30807;
wire wire30809;
wire wire30810;
wire wire30811;
wire wire30817;
wire wire30819;
wire wire30821;
wire wire30823;
wire wire30824;
wire wire30825;
wire wire30826;
wire wire30827;
wire wire30828;
wire wire30829;
wire wire30830;
wire wire30831;
wire wire30832;
wire wire30833;
wire wire30834;
wire wire30835;
wire wire30836;
wire wire30837;
wire wire30838;
wire wire30839;
wire wire30840;
wire wire30841;
wire wire30842;
wire wire30843;
wire wire30844;
wire wire30845;
wire wire30848;
wire wire30849;
wire wire30851;
wire wire30853;
wire wire30855;
wire wire30856;
wire wire30857;
wire wire30858;
wire wire30859;
wire wire30860;
wire wire30861;
wire wire30862;
wire wire30863;
wire wire30864;
wire wire30865;
wire wire30866;
wire wire30867;
wire wire30868;
wire wire30869;
wire wire30872;
wire wire30874;
wire wire30876;
wire wire30877;
wire wire30880;
wire wire30881;
wire wire30888;
wire wire30893;
wire wire30895;
wire wire30898;
wire wire30899;
wire wire30900;
wire wire30901;
wire wire30902;
wire wire30906;
wire wire30908;
wire wire30910;
wire wire30912;
wire wire30914;
wire wire30915;
wire wire30918;
wire wire30920;
wire wire30923;
wire wire30926;
wire wire30929;
wire wire30931;
wire wire30932;
wire wire30933;
wire wire30934;
wire wire30938;
wire wire30939;
wire wire30945;
wire wire30946;
wire wire30948;
wire wire30949;
wire wire30950;
wire wire30951;
wire wire30952;
wire wire30954;
wire wire30956;
wire wire30957;
wire wire30958;
wire wire30959;
wire wire30960;
wire wire30961;
wire wire30962;
wire wire30963;
wire wire30964;
wire wire30965;
wire wire30966;
wire wire30967;
wire wire30968;
wire wire30969;
wire wire30970;
wire wire30971;
wire wire30972;
wire wire30973;
wire wire30974;
wire wire30977;
wire wire30978;
wire wire30980;
wire wire30981;
wire wire30982;
wire wire30984;
wire wire30986;
wire wire30987;
wire wire30988;
wire wire30989;
wire wire30990;
wire wire30991;
wire wire30992;
wire wire30993;
wire wire30994;
wire wire30995;
wire wire30996;
wire wire30997;
wire wire30998;
wire wire31001;
wire wire31002;
wire wire31003;
wire wire31005;
wire wire31007;
wire wire31008;
wire wire31010;
wire wire31015;
wire wire31017;
wire wire31020;
wire wire31022;
wire wire31023;
wire wire31025;
wire wire31026;
wire wire31027;
wire wire31030;
wire wire31031;
wire wire31033;
wire wire31034;
wire wire31036;
wire wire31040;
wire wire31041;
wire wire31043;
wire wire31045;
wire wire31050;
wire wire31052;
wire wire31053;
wire wire31056;
wire wire31057;
wire wire31060;
wire wire31061;
wire wire31063;
wire wire31064;
wire wire31065;
wire wire31067;
wire wire31069;
wire wire31070;
wire wire31073;
wire wire31074;
wire wire31076;
wire wire31077;
wire wire31079;
wire wire31080;
wire wire31082;
wire wire31083;
wire wire31084;
wire wire31086;
wire wire31087;
wire wire31088;
wire wire31090;
wire wire31091;
wire wire31093;
wire wire31095;
wire wire31098;
wire wire31100;
wire wire31102;
wire wire31105;
wire wire31107;
wire wire31109;
wire wire31111;
wire wire31112;
wire wire31114;
wire wire31115;
wire wire31120;
wire wire31121;
wire wire31122;
wire wire31123;
wire wire31124;
wire wire31126;
wire wire31127;
wire wire31131;
wire wire31133;
wire wire31134;
wire wire31140;
wire wire31141;
wire wire31143;
wire wire31144;
wire wire31146;
wire wire31148;
wire wire31149;
wire wire31150;
wire wire31151;
wire wire31152;
wire wire31153;
wire wire31155;
wire wire31156;
wire wire31158;
wire wire31159;
wire wire31161;
wire wire31162;
wire wire31165;
wire wire31167;
wire wire31170;
wire wire31171;
wire wire31173;
wire wire31174;
wire wire31175;
wire wire31177;
wire wire31178;
wire wire31182;
wire wire31183;
wire wire31184;
wire wire31189;
wire wire31190;
wire wire31191;
wire wire31194;
wire wire31195;
wire wire31196;
wire wire31198;
wire wire31201;
wire wire31202;
wire wire31204;
wire wire31205;
wire wire31206;
wire wire31210;
wire wire31211;
wire wire31213;
wire wire31214;
wire wire31215;
wire wire31217;
wire wire31220;
wire wire31226;
wire wire31229;
wire wire31230;
wire wire31232;
wire wire31233;
wire wire31237;
wire wire31240;
wire wire31241;
wire wire31242;
wire wire31244;
wire wire31245;
wire wire31246;
wire wire31250;
wire wire31254;
wire wire31255;
wire wire31256;
wire wire31259;
wire wire31268;
wire wire31271;
wire wire31275;
wire wire31281;
wire wire31282;
wire wire31283;
wire wire31287;
wire wire31288;
wire wire31289;
wire wire31290;
wire wire31291;
wire wire31292;
wire wire31295;
wire wire31297;
wire wire31298;
wire wire31301;
wire wire31304;
wire wire31308;
wire wire31311;
wire wire31313;
wire wire31316;
wire wire31317;
wire wire31318;
wire wire31319;
wire wire31322;
wire wire31324;
wire wire31326;
wire wire31327;
wire wire31328;
wire wire31332;
wire wire31333;
wire wire31334;
wire wire31337;
wire wire31338;
wire wire31339;
wire wire31342;
wire wire31344;
wire wire31346;
wire wire31347;
wire wire31348;
wire wire31351;
wire wire31353;
wire wire31354;
wire wire31356;
wire wire31357;
wire wire31359;
wire wire31361;
wire wire31362;
wire wire31363;
wire wire31364;
wire wire31366;
wire wire31367;
wire wire31368;
wire wire31369;
wire wire31372;
wire wire31373;
wire wire31374;
wire wire31377;
wire wire31378;
wire wire31379;
wire wire31380;
wire wire31385;
wire wire31387;
wire wire31388;
wire wire31390;
wire wire31391;
wire wire31392;
wire wire31395;
wire wire31397;
wire wire31398;
wire wire31399;
wire wire31400;
wire wire31402;
wire wire31403;
wire wire31404;
wire wire31406;
wire wire31414;
wire wire31415;
wire wire31424;
wire wire31425;
wire wire31429;
wire wire31431;
wire wire31433;
wire wire31434;
wire wire31435;
wire wire31437;
wire wire31439;
wire wire31445;
wire wire31446;
wire wire31447;
wire wire31449;
wire wire31450;
wire wire31452;
wire wire31454;
wire wire31456;
wire wire31460;
wire wire31462;
wire wire31463;
wire wire31464;
wire wire31466;
wire wire31468;
wire wire31470;
wire wire31472;
wire wire31474;
wire wire31477;
wire wire31478;
wire wire31479;
wire wire31484;
wire wire31485;
wire wire31488;
wire wire31490;
wire wire31491;
wire wire31494;
wire wire31495;
wire wire31498;
wire wire31499;
wire wire31501;
wire wire31502;
wire wire31505;
wire wire31508;
wire wire31509;
wire wire31510;
wire wire31512;
wire wire31513;
wire wire31514;
wire wire31515;
wire wire31521;
wire wire31522;
wire wire31527;
wire wire31528;
wire wire31530;
wire wire31533;
wire wire31534;
wire wire31536;
wire wire31537;
wire wire31540;
wire wire31542;
wire wire31543;
wire wire31544;
wire wire31546;
wire wire31550;
wire wire31553;
wire wire31555;
wire wire31556;
wire wire31557;
wire wire31559;
wire wire31560;
wire wire31563;
wire wire31564;
wire wire31565;
wire wire31570;
wire wire31571;
wire wire31572;
wire wire31574;
wire wire31575;
wire wire31578;
wire wire31581;
wire wire31587;
wire wire31589;
wire wire31591;
wire wire31593;
wire wire31595;
wire wire31596;
wire wire31597;
wire wire31600;
wire wire31604;
wire wire31608;
wire wire31609;
wire wire31610;
wire wire31612;
wire wire31613;
wire wire31615;
wire wire31616;
wire wire31617;
wire wire31621;
wire wire31622;
wire wire31623;
wire wire31629;
wire wire31631;
wire wire31634;
wire wire31637;
wire wire31638;
wire wire31640;
wire wire31642;
wire wire31645;
wire wire31646;
wire wire31650;
wire wire31652;
wire wire31653;
wire wire31655;
wire wire31658;
wire wire31659;
wire wire31660;
wire wire31661;
wire wire31662;
wire wire31664;
wire wire31665;
wire wire31667;
wire wire31668;
wire wire31671;
wire wire31672;
wire wire31677;
wire wire31678;
wire wire31679;
wire wire31681;
wire wire31686;
wire wire31688;
wire wire31689;
wire wire31690;
wire wire31696;
wire wire31697;
wire wire31701;
wire wire31702;
wire wire31703;
wire wire31711;
wire wire31712;
wire wire31713;
wire wire31714;
wire wire31715;
wire wire31716;
wire wire31717;
wire wire31719;
wire wire31720;
wire wire31726;
wire wire31727;
wire wire31729;
wire wire31731;
wire wire31733;
wire wire31734;
wire wire31736;
wire wire31737;
wire wire31739;
wire wire31740;
wire wire31742;
wire wire31743;
wire wire31744;
wire wire31746;
wire wire31747;
wire wire31748;
wire wire31754;
wire wire31755;
wire wire31756;
wire wire31757;
wire wire31759;
wire wire31761;
wire wire31770;
wire wire31771;
wire wire31772;
wire wire31779;
wire wire31780;
wire wire31783;
wire wire31784;
wire wire31788;
wire wire31789;
wire wire31791;
wire wire31792;
wire wire31794;
wire wire31795;
wire wire31796;
wire wire31797;
wire wire31798;
wire wire31799;
wire wire31800;
wire wire31801;
wire wire31802;
wire wire31803;
wire wire31806;
wire wire31808;
wire wire31811;
wire wire31812;
wire wire31813;
wire wire31815;
wire wire31816;
wire wire31818;
wire wire31819;
wire wire31821;
wire wire31822;
wire wire31823;
wire wire31825;
wire wire31827;
wire wire31828;
wire wire31829;
wire wire31830;
wire wire31831;
wire wire31832;
wire wire31834;
wire wire31835;
wire wire31838;
wire wire31839;
wire wire31840;
wire wire31842;
wire wire31844;
wire wire31847;
wire wire31848;
wire wire31849;
wire wire31851;
wire wire31852;
wire wire31854;
wire wire31855;
wire wire31858;
wire wire31859;
wire wire31861;
wire wire31862;
wire wire31864;
wire wire31865;
wire wire31867;
wire wire31868;
wire wire31870;
wire wire31871;
wire wire31872;
wire wire31873;
wire wire31875;
wire wire31876;
wire wire31877;
wire wire31878;
wire wire31879;
wire wire31881;
wire wire31883;
wire wire31885;
wire wire31886;
wire wire31890;
wire wire31891;
wire wire31892;
wire wire31893;
wire wire31896;
wire wire31897;
wire wire31898;
wire wire31899;
wire wire31902;
wire wire31906;
wire wire31908;
wire wire31910;
wire wire31913;
wire wire31915;
wire wire31917;
wire wire31919;
wire wire31920;
wire wire31921;
wire wire31922;
wire wire31923;
wire wire31926;
wire wire31928;
wire wire31929;
wire wire31930;
wire wire31932;
wire wire31933;
wire wire31935;
wire wire31936;
wire wire31938;
wire wire31939;
wire wire31940;
wire wire31942;
wire wire31943;
wire wire31945;
wire wire31947;
wire wire31949;
wire wire31950;
wire wire31951;
wire wire31952;
wire wire31954;
wire wire31955;
wire wire31956;
wire wire31958;
wire wire31960;
wire wire31962;
wire wire31965;
wire wire31966;
wire wire31967;
wire wire31968;
wire wire31970;
wire wire31971;
wire wire31972;
wire wire31973;
wire wire31974;
wire wire31975;
wire wire31978;
wire wire31984;
wire wire31985;
wire wire31986;
wire wire31989;
wire wire31991;
wire wire31993;
wire wire31994;
wire wire31996;
wire wire31997;
wire wire31998;
wire wire32002;
wire wire32003;
wire wire32005;
wire wire32007;
wire wire32011;
wire wire32012;
wire wire32013;
wire wire32015;
wire wire32016;
wire wire32017;
wire wire32018;
wire wire32019;
wire wire32020;
wire wire32022;
wire wire32024;
wire wire32031;
wire wire32032;
wire wire32035;
wire wire32039;
wire wire32043;
wire wire32047;
wire wire32051;
wire wire32052;
wire wire32056;
wire wire32057;
wire wire32058;
wire wire32061;
wire wire32063;
wire wire32066;
wire wire32068;
wire wire32070;
wire wire32072;
wire wire32074;
wire wire32077;
wire wire32078;
wire wire32079;
wire wire32080;
wire wire32082;
wire wire32083;
wire wire32085;
wire wire32086;
wire wire32087;
wire wire32091;
wire wire32093;
wire wire32095;
wire wire32096;
wire wire32097;
wire wire32101;
wire wire32102;
wire wire32103;
wire wire32105;
wire wire32107;
wire wire32109;
wire wire32110;
wire wire32111;
wire wire32112;
wire wire32117;
wire wire32118;
wire wire32120;
wire wire32121;
wire wire32123;
wire wire32124;
wire wire32125;
wire wire32126;
wire wire32127;
wire wire32129;
wire wire32130;
wire wire32133;
wire wire32135;
wire wire32136;
wire wire32137;
wire wire32138;
wire wire32139;
wire wire32141;
wire wire32145;
wire wire32146;
wire wire32151;
wire wire32154;
wire wire32155;
wire wire32158;
wire wire32166;
wire wire32167;
wire wire32170;
wire wire32171;
wire wire32172;
wire wire32173;
wire wire32175;
wire wire32176;
wire wire32177;
wire wire32179;
wire wire32180;
wire wire32181;
wire wire32182;
wire wire32183;
wire wire32185;
wire wire32186;
wire wire32187;
wire wire32188;
wire wire32189;
wire wire32190;
wire wire32191;
wire wire32192;
wire wire32193;
wire wire32194;
wire wire32195;
wire wire32196;
wire wire32197;
wire wire32198;
wire wire32199;
wire wire32202;
wire wire32203;
wire wire32204;
wire wire32205;
wire wire32206;
wire wire32207;
wire wire32208;
wire wire32209;
wire wire32211;
wire wire32212;
wire wire32213;
wire wire32215;
wire wire32217;
wire wire32218;
wire wire32219;
wire wire32220;
wire wire32221;
wire wire32222;
wire wire32223;
wire wire32226;
wire wire32228;
wire wire32230;
wire wire32231;
wire wire32234;
wire wire32235;
wire wire32239;
wire wire32242;
wire wire32243;
wire wire32244;
wire wire32251;
wire wire32252;
wire wire32253;
wire wire32259;
wire wire32260;
wire wire32266;
wire wire32267;
wire wire32269;
wire wire32270;
wire wire32271;
wire wire32272;
wire wire32275;
wire wire32277;
wire wire32281;
wire wire32283;
wire wire32288;
wire wire32289;
wire wire32293;
wire wire32301;
wire wire32304;
wire wire32305;
wire wire32306;
wire wire32313;
wire wire32314;
wire wire32316;
wire wire32317;
wire wire32323;
wire wire32325;
wire wire32327;
wire wire32328;
wire wire32329;
wire wire32331;
wire wire32333;
wire wire32336;
wire wire32338;
wire wire32340;
wire wire32341;
wire wire32344;
wire wire32345;
wire wire32348;
wire wire32350;
wire wire32352;
wire wire32353;
wire wire32354;
wire wire32355;
wire wire32357;
wire wire32358;
wire wire32363;
wire wire32364;
wire wire32367;
wire wire32368;
wire wire32377;
wire wire32378;
wire wire32379;
wire wire32382;
wire wire32383;
wire wire32385;
wire wire32386;
wire wire32387;
wire wire32388;
wire wire32389;
wire wire32391;
wire wire32392;
wire wire32395;
wire wire32396;
wire wire32398;
wire wire32399;
wire wire32401;
wire wire32404;
wire wire32405;
wire wire32406;
wire wire32408;
wire wire32409;
wire wire32412;
wire wire32413;
wire wire32417;
wire wire32420;
wire wire32423;
wire wire32424;
wire wire32431;
wire wire32432;
wire wire32434;
wire wire32438;
wire wire32443;
wire wire32445;
wire wire32447;
wire wire32448;
wire wire32450;
wire wire32451;
wire wire32452;
wire wire32453;
wire wire32454;
wire wire32455;
wire wire32458;
wire wire32459;
wire wire32460;
wire wire32462;
wire wire32463;
wire wire32464;
wire wire32466;
wire wire32468;
wire wire32470;
wire wire32472;
wire wire32473;
wire wire32475;
wire wire32476;
wire wire32478;
wire wire32479;
wire wire32481;
wire wire32482;
wire wire32484;
wire wire32485;
wire wire32486;
wire wire32487;
wire wire32488;
wire wire32489;
wire wire32493;
wire wire32495;
wire wire32498;
wire wire32500;
wire wire32501;
wire wire32503;
wire wire32504;
wire wire32506;
wire wire32507;
wire wire32509;
wire wire32510;
wire wire32511;
wire wire32513;
wire wire32514;
wire wire32515;
wire wire32517;
wire wire32521;
wire wire32522;
wire wire32523;
wire wire32526;
wire wire32527;
wire wire32529;
wire wire32531;
wire wire32533;
wire wire32534;
wire wire32535;
wire wire32536;
wire wire32538;
wire wire32539;
wire wire32540;
wire wire32541;
wire wire32542;
wire wire32543;
wire wire32544;
wire wire32545;
wire wire32550;
wire wire32551;
wire wire32554;
wire wire32555;
wire wire32556;
wire wire32560;
wire wire32562;
wire wire32563;
wire wire32565;
wire wire32567;
wire wire32568;
wire wire32571;
wire wire32572;
wire wire32574;
wire wire32575;
wire wire32578;
wire wire32580;
wire wire32582;
wire wire32583;
wire wire32584;
wire wire32586;
wire wire32589;
wire wire32590;
wire wire32591;
wire wire32592;
wire wire32594;
wire wire32595;
wire wire32596;
wire wire32599;
wire wire32600;
wire wire32601;
wire wire32602;
wire wire32604;
wire wire32606;
wire wire32609;
wire wire32610;
wire wire32612;
wire wire32613;
wire wire32616;
wire wire32617;
wire wire32619;
wire wire32621;
wire wire32623;
wire wire32624;
wire wire32625;
wire wire32626;
wire wire32628;
wire wire32629;
wire wire32630;
wire wire32632;
wire wire32633;
wire wire32634;
wire wire32636;
wire wire32638;
wire wire32639;
wire wire32642;
wire wire32644;
wire wire32647;
wire wire32651;
wire wire32652;
wire wire32653;
wire wire32654;
wire wire32655;
wire wire32656;
wire wire32661;
wire wire32662;
wire wire32664;
wire wire32665;
wire wire32667;
wire wire32668;
wire wire32669;
wire wire32670;
wire wire32672;
wire wire32675;
wire wire32677;
wire wire32683;
wire wire32689;
wire wire32694;
wire wire32695;
wire wire32699;
wire wire32700;
wire wire32702;
wire wire32703;
wire wire32706;
wire wire32707;
wire wire32708;
wire wire32710;
wire wire32711;
wire wire32717;
wire wire32718;
wire wire32719;
wire wire32720;
wire wire32721;
wire wire32722;
wire wire32723;
wire wire32724;
wire wire32728;
wire wire32731;
wire wire32733;
wire wire32734;
wire wire32735;
wire wire32736;
wire wire32740;
wire wire32741;
wire wire32745;
wire wire32747;
wire wire32749;
wire wire32750;
wire wire32751;
wire wire32753;
wire wire32754;
wire wire32757;
wire wire32758;
wire wire32760;
wire wire32762;
wire wire32764;
wire wire32766;
wire wire32767;
wire wire32769;
wire wire32770;
wire wire32775;
wire wire32777;
wire wire32779;
wire wire32780;
wire wire32781;
wire wire32782;
wire wire32784;
wire wire32785;
wire wire32787;
wire wire32795;
wire wire32798;
wire wire32802;
wire wire32804;
wire wire32808;
wire wire32810;
wire wire32811;
wire wire32817;
wire wire32818;
wire wire32823;
wire wire32825;
wire wire32826;
wire wire32830;
wire wire32832;
wire wire32834;
wire wire32836;
wire wire32837;
wire wire32841;
wire wire32842;
wire wire32843;
wire wire32846;
wire wire32851;
wire wire32853;
wire wire32855;
wire wire32856;
wire wire32858;
wire wire32860;
wire wire32861;
wire wire32862;
wire wire32863;
wire wire32865;
wire wire32866;
wire wire32867;
wire wire32869;
wire wire32870;
wire wire32871;
wire wire32873;
wire wire32874;
wire wire32875;
wire wire32878;
wire wire32879;
wire wire32881;
wire wire32884;
wire wire32885;
wire wire32887;
wire wire32891;
wire wire32893;
wire wire32894;
wire wire32898;
wire wire32899;
wire wire32902;
wire wire32903;
wire wire32907;
wire wire32910;
wire wire32913;
wire wire32914;
wire wire32917;
wire wire32919;
wire wire32921;
wire wire32922;
wire wire32927;
wire wire32928;
wire wire32929;
wire wire32933;
wire wire32934;
wire wire32936;
wire wire32937;
wire wire32938;
wire wire32939;
wire wire32940;
wire wire32941;
wire wire32943;
wire wire32944;
wire wire32948;
wire wire32949;
wire wire32953;
wire wire32955;
wire wire32957;
wire wire32961;
wire wire32963;
wire wire32965;
wire wire32966;
wire wire32969;
wire wire32971;
wire wire32972;
wire wire32975;
wire wire32976;
wire wire32978;
wire wire32979;
wire wire32981;
wire wire32983;
wire wire32985;
wire wire32987;
wire wire32989;
wire wire32991;
wire wire32992;
wire wire32993;
wire wire32994;
wire wire32995;
wire wire32997;
wire wire32999;
wire wire33000;
wire wire33001;
wire wire33002;
wire wire33003;
wire wire33005;
wire wire33007;
wire wire33008;
wire wire33009;
wire wire33010;
wire wire33011;
wire wire33012;
wire wire33013;
wire wire33014;
wire wire33015;
wire wire33016;
wire wire33017;
wire wire33018;
wire wire33019;
wire wire33020;
wire wire33021;
wire wire33024;
wire wire33025;
wire wire33026;
wire wire33027;
wire wire33029;
wire wire33030;
wire wire33031;
wire wire33033;
wire wire33034;
wire wire33035;
wire wire33037;
wire wire33038;
wire wire33039;
wire wire33040;
wire wire33041;
wire wire33042;
wire wire33043;
wire wire33044;
wire wire33045;
wire wire33048;
wire wire33049;
wire wire33054;
wire wire33055;
wire wire33061;
wire wire33062;
wire wire33063;
wire wire33065;
wire wire33066;
wire wire33067;
wire wire33069;
wire wire33070;
wire wire33072;
wire wire33073;
wire wire33075;
wire wire33076;
wire wire33081;
wire wire33083;
wire wire33085;
wire wire33087;
wire wire33088;
wire wire33090;
wire wire33091;
wire wire33096;
wire wire33098;
wire wire33099;
wire wire33102;
wire wire33104;
wire wire33105;
wire wire33106;
wire wire33107;
wire wire33109;
wire wire33111;
wire wire33112;
wire wire33113;
wire wire33115;
wire wire33116;
wire wire33118;
wire wire33119;
wire wire33120;
wire wire33121;
wire wire33122;
wire wire33123;
wire wire33124;
wire wire33126;
wire wire33127;
wire wire33128;
wire wire33129;
wire wire33131;
wire wire33133;
wire wire33136;
wire wire33137;
wire wire33138;
wire wire33139;
wire wire33140;
wire wire33143;
wire wire33145;
wire wire33146;
wire wire33150;
wire wire33152;
wire wire33155;
wire wire33156;
wire wire33157;
wire wire33158;
wire wire33160;
wire wire33161;
wire wire33165;
wire wire33166;
wire wire33168;
wire wire33169;
wire wire33172;
wire wire33174;
wire wire33176;
wire wire33177;
wire wire33180;
wire wire33181;
wire wire33183;
wire wire33184;
wire wire33189;
wire wire33194;
wire wire33199;
wire wire33200;
wire wire33204;
wire wire33208;
wire wire33209;
wire wire33211;
wire wire33212;
wire wire33213;
wire wire33215;
wire wire33216;
wire wire33218;
wire wire33219;
wire wire33222;
wire wire33223;
wire wire33225;
wire wire33227;
wire wire33230;
wire wire33231;
wire wire33233;
wire wire33234;
wire wire33238;
wire wire33239;
wire wire33241;
wire wire33242;
wire wire33244;
wire wire33245;
wire wire33246;
wire wire33248;
wire wire33249;
wire wire33250;
wire wire33251;
wire wire33252;
wire wire33254;
wire wire33255;
wire wire33257;
wire wire33259;
wire wire33261;
wire wire33262;
wire wire33263;
wire wire33264;
wire wire33265;
wire wire33266;
wire wire33267;
wire wire33268;
wire wire33269;
wire wire33270;
wire wire33273;
wire wire33275;
wire wire33276;
wire wire33280;
wire wire33282;
wire wire33284;
wire wire33285;
wire wire33286;
wire wire33287;
wire wire33288;
wire wire33289;
wire wire33291;
wire wire33293;
wire wire33296;
wire wire33299;
wire wire33302;
wire wire33303;
wire wire33304;
wire wire33306;
wire wire33307;
wire wire33308;
wire wire33312;
wire wire33316;
wire wire33317;
wire wire33319;
wire wire33320;
wire wire33325;
wire wire33327;
wire wire33330;
wire wire33331;
wire wire33332;
wire wire33334;
wire wire33335;
wire wire33336;
wire wire33343;
wire wire33344;
wire wire33345;
wire wire33349;
wire wire33350;
wire wire33351;
wire wire33353;
wire wire33354;
wire wire33355;
wire wire33357;
wire wire33362;
wire wire33364;
wire wire33366;
wire wire33370;
wire wire33372;
wire wire33373;
wire wire33374;
wire wire33377;
wire wire33378;
wire wire33379;
wire wire33382;
wire wire33383;
wire wire33384;
wire wire33385;
wire wire33386;
wire wire33392;
wire wire33393;
wire wire33397;
wire wire33398;
wire wire33399;
wire wire33401;
wire wire33403;
wire wire33405;
wire wire33406;
wire wire33407;
wire wire33408;
wire wire33410;
wire wire33412;
wire wire33413;
wire wire33416;
wire wire33417;
wire wire33421;
wire wire33424;
wire wire33426;
wire wire33427;
wire wire33428;
wire wire33429;
wire wire33432;
wire wire33433;
wire wire33437;
wire wire33440;
wire wire33443;
wire wire33444;
wire wire33450;
wire wire33452;
wire wire33453;
wire wire33455;
wire wire33456;
wire wire33457;
wire wire33459;
wire wire33460;
wire wire33463;
wire wire33464;
wire wire33472;
wire wire33473;
wire wire33475;
wire wire33476;
wire wire33480;
wire wire33485;
wire wire33486;
wire wire33489;
wire wire33492;
wire wire33494;
wire wire33495;
wire wire33497;
wire wire33499;
wire wire33501;
wire wire33503;
wire wire33505;
wire wire33507;
wire wire33509;
wire wire33510;
wire wire33512;
wire wire33515;
wire wire33517;
wire wire33519;
wire wire33520;
wire wire33522;
wire wire33523;
wire wire33524;
wire wire33525;
wire wire33526;
wire wire33527;
wire wire33528;
wire wire33533;
wire wire33534;
wire wire33536;
wire wire33537;
wire wire33538;
wire wire33544;
wire wire33545;
wire wire33551;
wire wire33552;
wire wire33553;
wire wire33554;
wire wire33555;
wire wire33558;
wire wire33560;
wire wire33561;
wire wire33562;
wire wire33563;
wire wire33564;
wire wire33566;
wire wire33571;
wire wire33572;
wire wire33579;
wire wire33580;
wire wire33585;
wire wire33590;
wire wire33591;
wire wire33592;
wire wire33593;
wire wire33594;
wire wire33595;
wire wire33600;
wire wire33601;
wire wire33606;
wire wire33608;
wire wire33609;
wire wire33610;
wire wire33613;
wire wire33615;
wire wire33617;
wire wire33620;
wire wire33623;
wire wire33625;
wire wire33626;
wire wire33627;
wire wire33628;
wire wire33632;
wire wire33633;
wire wire33635;
wire wire33637;
wire wire33639;
wire wire33640;
wire wire33641;
wire wire33642;
wire wire33643;
wire wire33644;
wire wire33648;
wire wire33649;
wire wire33650;
wire wire33651;
wire wire33652;
wire wire33653;
wire wire33654;
wire wire33656;
wire wire33657;
wire wire33659;
wire wire33660;
wire wire33661;
wire wire33665;
wire wire33666;
wire wire33667;
wire wire33668;
wire wire33670;
wire wire33672;
wire wire33673;
wire wire33676;
wire wire33678;
wire wire33680;
wire wire33681;
wire wire33682;
wire wire33684;
wire wire33685;
wire wire33688;
wire wire33690;
wire wire33693;
wire wire33694;
wire wire33695;
wire wire33696;
wire wire33699;
wire wire33700;
wire wire33703;
wire wire33706;
wire wire33708;
wire wire33709;
wire wire33710;
wire wire33711;
wire wire33715;
wire wire33716;
wire wire33720;
wire wire33721;
wire wire33726;
wire wire33728;
wire wire33729;
wire wire33735;
wire wire33736;
wire wire33738;
wire wire33739;
wire wire33743;
wire wire33745;
wire wire33747;
wire wire33749;
wire wire33750;
wire wire33751;
wire wire33752;
wire wire33754;
wire wire33755;
wire wire33756;
wire wire33758;
wire wire33759;
wire wire33760;
wire wire33765;
wire wire33767;
wire wire33770;
wire wire33771;
wire wire33773;
wire wire33775;
wire wire33777;
wire wire33778;
wire wire33779;
wire wire33780;
wire wire33781;
wire wire33784;
wire wire33786;
wire wire33789;
wire wire33794;
wire wire33795;
wire wire33798;
wire wire33800;
wire wire33803;
wire wire33804;
wire wire33805;
wire wire33812;
wire wire33813;
wire wire33814;
wire wire33817;
wire wire33818;
wire wire33820;
wire wire33821;
wire wire33823;
wire wire33824;
wire wire33826;
wire wire33827;
wire wire33830;
wire wire33832;
wire wire33834;
wire wire33836;
wire wire33837;
wire wire33838;
wire wire33839;
wire wire33842;
wire wire33846;
wire wire33847;
wire wire33850;
wire wire33851;
wire wire33854;
wire wire33857;
wire wire33860;
wire wire33862;
wire wire33865;
wire wire33866;
wire wire33869;
wire wire33870;
wire wire33871;
wire wire33873;
wire wire33875;
wire wire33877;
wire wire33879;
wire wire33886;
wire wire33887;
wire wire33888;
wire wire33889;
wire wire33895;
wire wire33896;
wire wire33898;
wire wire33902;
wire wire33903;
wire wire33908;
wire wire33909;
wire wire33912;
wire wire33913;
wire wire33916;
wire wire33917;
wire wire33918;
wire wire33919;
wire wire33920;
wire wire33922;
wire wire33924;
wire wire33925;
wire wire33926;
wire wire33927;
wire wire33931;
wire wire33934;
wire wire33936;
wire wire33937;
wire wire33938;
wire wire33939;
wire wire33943;
wire wire33944;
wire wire33949;
wire wire33950;
wire wire33954;
wire wire33955;
wire wire33956;
wire wire33960;
wire wire33961;
wire wire33962;
wire wire33963;
wire wire33964;
wire wire33970;
wire wire33971;
wire wire33973;
wire wire33974;
wire wire33975;
wire wire33976;
wire wire33977;
wire wire33979;
wire wire33980;
wire wire33983;
wire wire33985;
wire wire33988;
wire wire33990;
wire wire33993;
wire wire33996;
wire wire33997;
wire wire33998;
wire wire34000;
wire wire34001;
wire wire34004;
wire wire34005;
wire wire34007;
wire wire34008;
wire wire34009;
wire wire34010;
wire wire34016;
wire wire34017;
wire wire34022;
wire wire34023;
wire wire34028;
wire wire34029;
wire wire34034;
wire wire34035;
wire wire34038;
wire wire34041;
wire wire34044;
wire wire34047;
wire wire34050;
wire wire34051;
wire wire34052;
wire wire34053;
wire wire34054;
wire wire34057;
wire wire34059;
wire wire34061;
wire wire34062;
wire wire34063;
wire wire34064;
wire wire34065;
wire wire34066;
wire wire34067;
wire wire34070;
wire wire34071;
wire wire34072;
wire wire34073;
wire wire34074;
wire wire34076;
wire wire34078;
wire wire34079;
wire wire34082;
wire wire34083;
wire wire34085;
wire wire34086;
wire wire34088;
wire wire34089;
wire wire34091;
wire wire34092;
wire wire34094;
wire wire34095;
wire wire34096;
wire wire34099;
wire wire34101;
wire wire34104;
wire wire34105;
wire wire34106;
wire wire34109;
wire wire34111;
wire wire34112;
wire wire34113;
wire wire34116;
wire wire34118;
wire wire34120;
wire wire34121;
wire wire34124;
wire wire34126;
wire wire34127;
wire wire34130;
wire wire34132;
wire wire34133;
wire wire34136;
wire wire34138;
wire wire34139;
wire wire34142;
wire wire34144;
wire wire34145;
wire wire34149;
wire wire34150;
wire wire34151;
wire wire34154;
wire wire34156;
wire wire34159;
wire wire34160;
wire wire34161;
wire wire34166;
wire wire34167;
wire wire34169;
wire wire34170;
wire wire34173;
wire wire34174;
wire wire34177;
wire wire34178;
wire wire34181;
wire wire34182;
wire wire34185;
wire wire34186;
wire wire34188;
wire wire34189;
wire wire34193;
wire wire34198;
wire wire34199;
wire wire34201;
wire wire34202;
wire wire34203;
wire wire34204;
wire wire34206;
wire wire34207;
wire wire34208;
wire wire34211;
wire wire34212;
wire wire34215;
wire wire34216;
wire wire34219;
wire wire34220;
wire wire34225;
wire wire34226;
wire wire34229;
wire wire34230;
wire wire34231;
wire wire34232;
wire wire34234;
wire wire34235;
wire wire34236;
wire wire34239;
wire wire34241;
wire wire34242;
wire wire34244;
wire wire34248;
wire wire34256;
wire wire34258;
wire wire34259;
wire wire34262;
wire wire34263;
wire wire34265;
wire wire34266;
wire wire34267;
wire wire34271;
wire wire34275;
wire wire34278;
wire wire34279;
wire wire34280;
wire wire34281;
wire wire34290;
wire wire34292;
wire wire34294;
wire wire34296;
reg ng6215;

reg ng4332;

reg ng2837;

reg ng1135;

reg ng2485;

reg ng4375;

reg pg9251;

reg ng1171;

reg ng3235;

reg ng2852;

reg ng222;

reg pg8719;

reg ng2815;

reg ng4888;

reg ng433;

reg ng246;

reg ng102;

reg ng1030;

reg ng110;

reg pg13966;

reg ng4801;

reg ng4045;

reg ng2145;

reg ng5138;

reg ng3873;

reg ng3752;

reg ng136;

reg ng1772;

reg ng990;

reg ng3171;

reg ng168;

reg ng441;

reg ng160;

reg pg17577;

reg ng1361;

reg ng6621;

reg ng5689;

reg ng6593;

reg ng5827;

reg pg17316;

reg ng74;

reg ng4443;

reg ng979;

reg ng1484;

reg ng6044;

reg ng3817;

reg ng316;

reg pg14167;

reg ng499;

reg pg17739;

reg pg8279;

reg ng2269;

reg ng2927;

reg ng577;

reg ng599;

reg pg8870;

reg ng781;

reg ng2759;

reg ng2715;

reg ng1870;

reg ng1768;

reg ng4031;

reg ng6181;

reg ng2173;

reg ng1783;

reg ng106;

reg ng2803;

reg ng6303;

reg ng3462;

reg ng482;

reg ng1811;

reg ng2890;

reg ng1542;

reg ng111;

reg ng2161;

reg ng947;

reg ng546;

reg ng3913;

reg pg12923;

reg pg8915;

reg ng5599;

reg ng3893;

reg ng4141;

reg ng3106;

reg ng3841;

reg ng2004;

reg ng3586;

reg ng939;

reg ng6195;

reg ng925;

reg ng6255;

reg ng2177;

reg ng5835;

reg ng4543;

reg ng5802;

reg ng5092;

reg ng3933;

reg pg17715;

reg ng911;

reg ng3901;

reg ng4297;

reg pg8475;

reg ng4049;

reg ng3139;

reg pg13881;

reg ng6649;

reg ng2599;

reg ng4087;

reg ng1467;

reg ng6519;

reg ng1700;

reg ng1950;

reg pg13926;

reg ng2417;

reg ng475;

reg ng333;

reg pg9553;

reg pg12422;

reg ng1779;

reg ng2834;

reg ng3470;

reg ng5188;

reg pg13259;

reg ng504;

reg ng6541;

reg ng6209;

reg ng5685;

reg pg7916;

reg ng3466;

reg ng3333;

reg ng4922;

reg ng6613;

reg ng93;

reg pg12368;

reg pg17787;

reg ng1478;

reg ng63;

reg ng2643;

reg ng191;

reg ng1620;

reg pg16924;

reg ng2495;

reg ng5583;

reg ng2138;

reg ng5244;

reg ng936;

reg ng429;

reg ng4854;

reg ng37;

reg ng6381;

reg ng347;

reg pg9019;

reg ng2767;

reg pg8788;

reg ng5921;

reg pg14673;

reg ng85;

reg ng5069;

reg ng1061;

reg ng4401;

reg pg14421;

reg ng3610;

reg ng4975;

reg ng4427;

reg ng4145;

reg ng1834;

reg ng5703;

reg pg10306;

reg ng1141;

reg ng4512;

reg ng4253;

reg ng4570;

reg ng1548;

reg ng4284;

reg ng385;

reg ng291;

reg pg17711;

reg ng3111;

reg ng718;

reg ng6267;

reg ng2399;

reg ng2898;

reg pg7257;

reg ng4831;

reg ng5889;

reg ng822;

reg ng43;

reg pg17649;

reg ng2112;

reg ng5543;

reg pg7260;

reg ng142;

reg ng5022;

reg ng6148;

reg ng1448;

reg ng3961;

reg ng1018;

reg ng5029;

reg ng513;

reg ng5109;

reg ng2016;

reg ng5575;

reg ng5052;

reg ng1992;

reg ng2902;

reg ng3808;

reg ng1608;

reg ng5535;

reg ng405;

reg pg8291;

reg pg9555;

reg ng3203;

reg ng655;

reg ng4423;

reg ng4633;

reg ng4116;

reg ng298;

reg pg17291;

reg ng4501;

reg ng6513;

reg ng5240;

reg ng1002;

reg ng896;

reg ng3451;

reg ng2712;

reg ng5929;

reg pg9743;

reg ng837;

reg ng2437;

reg pg17743;

reg pg16744;

reg ng785;

reg ng2575;

reg pg17871;

reg ng3925;

reg wire1457;

reg ng4765;

reg ng1266;

reg ng6605;

reg ng2868;

reg ng6573;

reg ng5485;

reg ng1211;

reg ng1821;

reg ng5124;

reg pg12470;

reg ng790;

reg ng5142;

reg ng3594;

reg ng5953;

reg pg14635;

reg ng6561;

reg ng2775;

reg ng4366;

reg ng5016;

reg pg13049;

reg ng5128;

reg ng5456;

reg ng4674;

reg ng4153;

reg ng117;

reg ng3239;

reg ng1437;

reg wire1421;

reg ng4269;

reg ng3343;

reg ng2819;

reg ng3050;

reg ng4495;

reg ng1070;

reg pg16775;

reg ng6251;

reg ng1283;

reg ng6537;

reg ng2932;

reg ng4584;

reg pg16955;

reg pg9680;

reg pg14125;

reg ng2984;

reg pg17320;

reg ng1256;

reg ng2841;

reg ng2307;

reg pg9615;

reg ng31;

reg ng4455;

reg ng9;

reg pg8785;

reg ng4950;

reg ng5216;

reg ng1936;

reg ng1668;

reg pg14662;

reg ng3689;

reg ng4146;

reg ng4681;

reg ng827;

reg ng287;

reg ng1277;

reg ng2799;

reg ng1945;

reg ng776;

reg ng358;

reg ng626;

reg ng4340;

reg ng2036;

reg ng1249;

reg ng2102;

reg ng6173;

reg ng2338;

reg ng6741;

reg ng65;

reg pg17845;

reg ng6509;

reg ng2070;

reg ng5563;

reg ng4473;

reg ng2445;

reg ng2407;

reg ng1677;

reg ng86;

reg ng2827;

reg pg17400;

reg ng1306;

reg ng1514;

reg ng4727;

reg ng3219;

reg ng6597;

reg ng5913;

reg ng3259;

reg ng2999;

reg ng2472;

reg ng3195;

reg ng4417;

reg ng2922;

reg ng3401;

reg ng3119;

reg ng3211;

reg ng3821;

reg ng3191;

reg ng2527;

reg ng3243;

reg ng5204;

reg ng1862;

reg ng1178;

reg pg14779;

reg ng3530;

reg ng4273;

reg ng4572;

reg ng2259;

reg ng6191;

reg ng6307;

reg ng4281;

reg ng4639;

reg ng5037;

reg ng6279;

reg ng5297;

reg pg8916;

reg ng232;

reg ng3498;

reg ng6555;

reg ng1472;

reg ng4760;

reg ng2204;

reg ng862;

reg ng6736;

reg ng6500;

reg ng2724;

reg ng2882;

reg ng2541;

reg ng6653;

reg ng4894;

reg ng2476;

reg ng2729;

reg pg16874;

reg ng930;

reg ng6682;

reg ng2873;

reg ng4899;

reg pg8919;

reg ng3484;

reg ng604;

reg ng1825;

reg ng4392;

reg ng4520;

reg ng1395;

reg ng714;

reg ng79;

reg ng6505;

reg ng5462;

reg ng5073;

reg ng1636;

reg ng5849;

reg ng2197;

reg ng1858;

reg ng6581;

reg ng1902;

reg ng2126;

reg pg8786;

reg ng582;

reg ng3845;

reg ng2079;

reg ng5841;

reg ng4239;

reg ng5148;

reg pg17604;

reg pg17607;

reg pg17685;

reg ng128;

reg ng2610;

reg ng6727;

reg ng3143;

reg ng4927;

reg ng5077;

reg ng2342;

reg ng3574;

reg ng2319;

reg ng5752;

reg ng1041;

reg ng4467;

reg ng2279;

reg pg14189;

reg ng2606;

reg ng262;

reg ng3502;

reg ng5817;

reg ng4944;

reg ng3827;

reg ng4704;

reg ng336;

reg ng2153;

reg ng3480;

reg pg17678;

reg ng4646;

reg ng5357;

reg ng4907;

reg ng3937;

reg ng5949;

reg ng1854;

reg ng4064;

reg ng6247;

reg ng1259;

reg ng6589;

reg ng1322;

reg ng1913;

reg ng5489;

reg ng182;

reg ng1592;

reg ng2689;

reg pg14217;

reg ng2509;

reg ng3921;

reg ng1756;

reg ng2950;

reg ng446;

reg ng4349;

reg ng6163;

reg ng5248;

reg pg7245;

reg pg11447;

reg ng2116;

reg ng2697;

reg pg16722;

reg ng2453;

reg ng4420;

reg ng3606;

reg ng843;

reg ng3506;

reg ng1036;

reg ng4104;

reg ng1706;

reg ng5523;

reg ng6159;

reg ng2960;

reg ng5495;

reg ng2975;

reg ng6549;

reg ng2315;

reg ng2595;

reg ng6545;

reg ng2652;

reg ng6235;

reg ng542;

reg ng1840;

reg ng703;

reg pg9497;

reg ng4072;

reg ng3133;

reg ng22;

reg ng1906;

reg ng4912;

reg ng1959;

reg ng3857;

reg ng2375;

reg ng4991;

reg ng2946;

reg ng2831;

reg ng739;

reg ng5084;

reg ng4785;

reg ng2791;

reg ng6609;

reg ng2098;

reg ng3546;

reg ng2185;

reg ng2491;

reg ng1312;

reg ng1129;

reg ng1221;

reg ng1624;

reg ng1848;

reg ng4859;

reg wire1411;

reg ng2994;

reg ng956;

reg ng2421;

reg ng6533;

reg ng370;

reg ng1874;

reg ng4125;

reg ng5481;

reg ng7;

reg ng2361;

reg ng2327;

reg ng723;

reg ng94;

reg ng3703;

reg ng4549;

reg ng4180;

reg ng1926;

reg ng676;

reg ng4558;

reg ng4864;

reg ng1532;

reg ng1389;

reg pg16627;

reg ng3802;

reg ng2255;

reg ng5499;

reg pg11770;

reg ng5917;

reg ng6167;

reg ng3917;

reg ng2537;

reg ng5268;

reg ng3881;

reg ng5256;

reg ng4732;

reg pg7540;

reg pg17813;

reg ng2878;

reg ng933;

reg ng4157;

reg ng3863;

reg pg16693;

reg ng1657;

reg pg17819;

reg ng4035;

reg ng667;

reg ng5475;

reg ng5603;

reg ng2719;

reg ng3949;

reg ng209;

reg ng4462;

reg ng4249;

reg ng5236;

reg pg8917;

reg ng4849;

reg pg16718;

reg ng2227;

reg ng5062;

reg ng34;

reg ng424;

reg ng1280;

reg ng650;

reg ng2181;

reg ng1046;

reg ng1345;

reg ng5694;

reg ng2441;

reg ng4821;

reg ng3694;

reg ng2779;

reg ng376;

reg ng907;

reg ng699;

reg ng3129;

reg ng4698;

reg ng6035;

reg ng4507;

reg ng4040;

reg ng5555;

reg ng590;

reg ng1752;

reg ng4477;

reg ng1296;

reg ng4382;

reg ng1052;

reg ng1728;

reg ng969;

reg ng355;

reg pg17639;

reg pg9817;

reg ng225;

reg ng5869;

reg ng153;

reg ng2811;

reg ng1585;

reg ng4108;

reg ng5881;

reg ng1146;

reg ng518;

reg ng4531;

reg ng5041;

reg ng2988;

reg ng1526;

reg ng568;

reg pg10122;

reg ng4546;

reg ng6098;

reg ng6283;

reg ng5120;

reg pg19357;

reg ng4322;

reg ng5252;

reg ng1274;

reg ng112;

reg ng5033;

reg ng4939;

reg ng5097;

reg ng5112;

reg ng3329;

reg ng943;

reg ng5200;

reg ng2912;

reg ng3352;

reg ng3125;

reg ng1988;

reg ng5348;

reg pg12832;

reg ng1878;

reg ng2547;

reg ng5343;

reg pg13099;

reg ng5567;

reg pg10500;

reg ng753;

reg ng351;

reg ng3179;

reg ng2807;

reg ng1682;

reg ng5831;

reg ng3231;

reg ng4486;

reg ng5579;

reg ng6625;

reg pg8398;

reg ng4388;

reg ng4564;

reg ng4308;

reg ng2625;

reg ng3897;

reg ng2860;

reg ng6641;

reg ng3538;

reg ng6523;

reg ng3263;

reg ng3562;

reg pg14828;

reg ng5937;

reg ng1242;

reg ng4771;

reg pg14705;

reg ng4966;

reg pg17674;

reg ng1199;

reg ng5941;

reg ng1152;

reg pg13085;

reg ng2856;

reg ng4818;

reg pg19334;

reg ng1964;

reg ng19;

reg ng5170;

reg ng1559;

reg ng4843;

reg pg14694;

reg ng6657;

reg ng2894;

reg ng4311;

reg ng3223;

reg ng3251;

reg ng5619;

reg ng559;

reg ng554;

reg ng1798;

reg ng4871;

reg ng1579;

reg ng4643;

reg ng2980;

reg ng5901;

reg ng479;

reg ng4653;

reg ng1105;

reg ng3889;

reg ng4098;

reg ng4504;

reg ng1589;

reg ng5990;

reg ng6275;

reg ng6239;

reg ng4571;

reg ng5406;

reg ng150;

reg ng538;

reg ng4743;

reg ng5571;

reg ng5196;

reg ng2351;

reg ng4434;

reg ng301;

reg ng854;

reg ng2518;

reg pg17646;

reg pg17764;

reg ng1236;

reg ng4616;

reg ng2523;

reg ng2551;

reg pg14749;

reg ng2579;

reg pg17519;

reg ng3929;

reg ng2012;

reg ng4836;

reg ng2108;

reg ng2571;

reg ng2093;

reg ng1554;

reg ng3207;

reg pg16748;

reg ng1720;

reg ng1193;

reg ng3255;

reg ng5893;

reg ng4456;

reg pg9682;

reg ng1300;

reg ng4552;

reg ng3187;

reg ng1996;

reg pg11388;

reg ng496;

reg pg14096;

reg ng4722;

reg ng6154;

reg ng5264;

reg ng3151;

reg ng2886;

reg ng6386;

reg ng4054;

reg ng1087;

reg ng3476;

reg ng4575;

reg ng5873;

reg ng4578;

reg ng4459;

reg ng6311;

reg ng4826;

reg pg13895;

reg ng3338;

reg ng1696;

reg ng6;

reg ng3578;

reg ng2380;

reg ng2648;

reg ng341;

reg ng4601;

reg ng2567;

reg ng890;

reg ng2864;

reg ng28;

reg ng4561;

reg ng5156;

reg ng2273;

reg ng904;

reg ng6227;

reg ng6203;

reg ng66;

reg pg13068;

reg ng2165;

reg ng4112;

reg ng1982;

reg ng4717;

reg ng4483;

reg ng3215;

reg ng1367;

reg ng2051;

reg ng1691;

reg ng1111;

reg ng5821;

reg ng411;

reg ng4057;

reg pg16686;

reg ng2661;

reg ng2970;

reg ng4628;

reg ng2771;

reg ng3570;

reg ng622;

reg ng3853;

reg ng2941;

reg ng3100;

reg ng4737;

reg ng4754;

reg ng4983;

reg ng4961;

reg ng3494;

reg ng4749;

reg ng2465;

reg ng4917;

reg ng3680;

reg ng1748;

reg pg8215;

reg ng758;

reg pg12919;

reg ng1664;

reg ng528;

reg ng2848;

reg ng1564;

reg ng962;

reg ng3831;

reg ng4793;

reg ng5808;

reg pg17760;

reg ng1890;

reg pg12184;

reg ng5897;

reg pg14597;

reg ng4093;

reg ng2619;

reg ng661;

reg ng6494;

reg ng1413;

reg ng2311;

reg ng794;

reg ng2667;

reg ng2555;

reg ng4581;

reg ng1616;

reg ng305;

reg ng255;

reg ng613;

reg ng817;

reg ng686;

reg ng4489;

reg ng4955;

reg ng2675;

reg ng25;

reg ng329;

reg pg17722;

reg pg17778;

reg ng2533;

reg ng2936;

reg pg16603;

reg ng6299;

reg ng319;

reg ng1351;

reg pg16624;

reg ng728;

reg ng2084;

reg ng691;

reg ng5698;

reg ng4515;

reg ng1882;

reg pg9048;

reg ng6336;

reg ng5134;

reg ng4076;

reg ng1495;

reg pg16659;

reg ng5160;

reg ng1189;

reg ng437;

reg ng5511;

reg ng3965;

reg ng6187;

reg ng914;

reg ng5551;

reg ng1373;

reg ng632;

reg ng1246;

reg ng4498;

reg ng2241;

reg ng2370;

reg ng2756;

reg ng2514;

reg ng2763;

reg ng6645;

reg ng3869;

reg ng2629;

reg ng3639;

reg ng269;

reg ng3957;

reg ng1183;

reg ng4669;

reg ng4411;

reg ng3602;

reg ng4688;

reg ng3227;

reg pg13906;

reg ng2040;

reg ng5857;

reg ng8;

reg ng550;

reg ng283;

reg ng2795;

reg pg8358;

reg ng6049;

reg ng4082;

reg ng1252;

reg ng5527;

reg ng5224;

reg ng1287;

reg ng1644;

reg ng5176;

reg ng1536;

reg ng5228;

reg ng3849;

reg ng2303;

reg pg8277;

reg ng324;

reg ng6527;

reg ng5644;

reg pg8416;

reg ng3953;

reg ng164;

reg ng1648;

reg ng6295;

reg ng1792;

reg ng2583;

reg pg8342;

reg ng278;

reg ng6395;

reg pg17404;

reg ng763;

reg ng1632;

reg ng744;

reg ng1442;

reg ng1454;

reg ng2287;

reg ng3566;

reg ng681;

reg ng3518;

reg ng736;

reg pg17580;

reg ng3835;

reg ng5339;

reg ng174;

reg ng2783;

reg pg14738;

reg ng6243;

reg ng16;

reg ng239;

reg ng4452;

reg pg14147;

reg ng5164;

reg pg8918;

reg ng2461;

reg ng4369;

reg ng3288;

reg ng1263;

reg ng4664;

reg ng2047;

reg ng4430;

reg ng572;

reg ng3990;

reg ng812;

reg ng3684;

reg ng401;

reg ng586;

reg ng2393;

reg pg13039;

reg ng2587;

reg ng6271;

reg ng2020;

reg ng460;

reg ng3247;

reg pg8789;

reg ng199;

reg ng5080;

reg ng2965;

reg ng1404;

reg ng617;

reg ng3161;

reg ng1844;

reg ng1955;

reg ng671;

reg ng1270;

reg ng5925;

reg ng2787;

reg ng6601;

reg ng4119;

reg ng5845;

reg pg17688;

reg ng3550;

reg ng1687;

reg ng1710;

reg ng5152;

reg ng2060;

reg ng5046;

reg pg8920;

reg ng4519;

reg ng3614;

reg ng5272;

reg ng4358;

reg ng3003;

reg ng5260;

reg ng4300;

reg ng71;

reg ng2299;

reg ng4492;

reg pg8344;

reg ng3905;

reg pg12238;

reg ng1917;

reg ng5965;

reg ng5933;

reg ng5611;

reg ng4534;

reg ng417;

reg ng1604;

reg ng2008;

reg ng2122;

reg ng2433;

reg ng4164;

reg ng6637;

reg ng3558;

reg ng157;

reg pg13272;

reg ng5961;

reg ng6629;

reg ng1216;

reg ng1430;

reg ng5208;

reg ng1333;

reg ng101;

reg ng1816;

reg ng2403;

reg ng952;

reg ng2223;

reg ng5957;

reg pg8783;

reg ng2130;

reg ng832;

reg ng2823;

reg ng6040;

reg ng1760;

reg pg14201;

reg ng2193;

reg ng996;

reg ng4474;

reg ng4480;

reg ng3582;

reg pg14518;

reg ng5467;

reg ng4608;

reg ng1894;

reg ng5011;

reg ng5863;

reg ng6444;

reg ng5220;

reg ng2384;

reg ng4527;

reg ng1489;

reg pg8839;

reg ng3347;

reg ng2265;

reg ng1974;

reg ng1124;

reg ng2429;

reg ng1978;

reg ng6390;

reg ng3199;

reg ng1740;

reg ng2681;

reg ng2413;

reg ng5352;

reg ng6617;

reg ng2704;

reg ng2250;

reg ng2357;

reg ng5115;

reg ng5595;

reg ng2735;

reg ng4659;

reg ng1094;

reg ng534;

reg ng1521;

reg pg8787;

reg ng59;

reg ng772;

reg ng2563;

reg ng3598;

reg ng294;

reg ng921;

reg ng3522;

reg ng1379;

reg ng5587;

reg pg7946;

reg ng4264;

reg ng6291;

reg ng2955;

reg ng3115;

reg ng1724;

reg ng6177;

reg ng4593;

reg ng1024;

reg pg16656;

reg ng203;

reg ng5057;

reg ng6377;

reg ng4776;

reg ng5591;

reg ng5507;

reg ng452;

reg ng807;

reg ng1600;

reg ng4621;

reg ng1099;

reg ng2024;

reg ng4242;

reg ng2741;

reg ng2217;

reg ng6219;

reg ng1714;

reg ng1968;

reg ng4878;

reg pg11349;

reg pg8784;

reg ng5503;

reg pg11678;

reg ng595;

reg ng3542;

reg ng847;

reg pg12350;

reg ng1736;

reg ng2389;

reg ng2638;

reg ng2066;

reg ng4258;

reg ng5232;

reg ng6031;

reg ng4235;

reg ng3147;

reg ng4438;

reg ng5547;

reg ng4122;

reg ng1319;

reg ng1612;

reg ng5813;

reg ng4172;

reg ng490;

reg ng3457;

reg ng2844;

reg ng4709;

reg ng1291;

reg ng2449;

reg ng5212;

reg ng1830;

reg pg7243;

reg ng2907;

reg ng976;

reg ng2236;

reg pg12300;

reg ng6287;

reg ng5180;

reg ng918;

reg ng5945;

reg ng5517;

reg ng4245;

reg ng2246;

reg ng1932;

reg pg10527;

reg ng3941;

reg ng1744;

reg ng3512;

reg pg14451;

reg ng2657;

reg ng4933;

reg ng608;

reg ng1886;

reg ng1008;

reg ng645;

reg ng392;

reg ng146;

reg ng2671;

reg ng6565;

reg ng5909;

reg ng4372;

reg ng3155;

reg ng5607;

reg ng4521;

reg ng562;

reg ng4291;

reg ng3590;

reg ng218;

reg ng2028;

reg ng2685;

reg ng1802;

reg ng3490;

reg ng3167;

reg ng2295;

reg pg13865;

reg ng3813;

reg ng1205;

reg ng2208;

reg ng732;

reg ng4176;

reg ng6263;

reg ng4540;

reg ng121;

reg ng6732;

reg ng3554;

reg ng749;

reg ng5615;

reg ng6199;

reg ng2089;

reg pg9741;

reg ng3909;

reg ng2917;

reg ng2504;

reg pg11418;

reg ng2331;

reg ng6723;

reg ng6585;

reg ng6633;

reg ng4555;

reg ng4567;

reg ng1339;

reg ng767;

reg pg9617;

reg ng6259;

reg ng4405;

reg ng3945;

reg ng2748;

reg ng2283;

reg pg17423;

reg ng3698;

reg ng311;

reg ng1384;

reg ng5853;

reg ng5559;

reg ng5905;

reg ng872;

reg ng5471;

reg ng2169;

always  @(posedge pclk)
	ng6215<=ng33063;

 always  @(posedge pclk)
	ng4332<=ng34455;

 always  @(posedge pclk)
	ng2837<=ng24264;

 always  @(posedge pclk)
	ng1135<=ng26917;

 always  @(posedge pclk)
	ng2485<=ng33013;

 always  @(posedge pclk)
	ng4375<=ng26951;

 always  @(posedge pclk)
	pg9251<=ng24281;

 always  @(posedge pclk)
	ng1171<=ng30338;

 always  @(posedge pclk)
	ng3235<=ng30403;

 always  @(posedge pclk)
	ng2852<=ng34610;

 always  @(posedge pclk)
	ng222<=ng33537;

 always  @(posedge pclk)
	pg8719<=ng25595;

 always  @(posedge pclk)
	ng2815<=ng34446;

 always  @(posedge pclk)
	ng4888<=ng34266;

 always  @(posedge pclk)
	ng433<=ng24205;

 always  @(posedge pclk)
	ng246<=ng26907;

 always  @(posedge pclk)
	ng102<=ng33962;

 always  @(posedge pclk)
	ng1030<=ng32983;

 always  @(posedge pclk)
	ng110<=ng30286;

 always  @(posedge pclk)
	pg13966<=pg11418;

 always  @(posedge pclk)
	ng4801<=ng34030;

 always  @(posedge pclk)
	ng4045<=ng24277;

 always  @(posedge pclk)
	ng2145<=ng34605;

 always  @(posedge pclk)
	ng5138<=ng29283;

 always  @(posedge pclk)
	ng3873<=ng33033;

 always  @(posedge pclk)
	ng3752<=ng25678;

 always  @(posedge pclk)
	ng136<=ng34598;

 always  @(posedge pclk)
	ng1772<=ng33553;

 always  @(posedge pclk)
	ng990<=pg8416;

 always  @(posedge pclk)
	ng3171<=ng33023;

 always  @(posedge pclk)
	ng168<=ng25600;

 always  @(posedge pclk)
	ng441<=ng24207;

 always  @(posedge pclk)
	ng160<=ng34249;

 always  @(posedge pclk)
	pg17577<=pg17519;

 always  @(posedge pclk)
	ng1361<=ng30343;

 always  @(posedge pclk)
	ng6621<=ng30551;

 always  @(posedge pclk)
	ng5689<=ng24341;

 always  @(posedge pclk)
	ng6593<=ng30546;

 always  @(posedge pclk)
	ng5827<=ng29294;

 always  @(posedge pclk)
	pg17316<=pg17291;

 always  @(posedge pclk)
	ng74<=ng26893;

 always  @(posedge pclk)
	ng4443<=pg7260;

 always  @(posedge pclk)
	ng979<=pg13259;

 always  @(posedge pclk)
	ng1484<=ng29238;

 always  @(posedge pclk)
	ng6044<=ng24347;

 always  @(posedge pclk)
	ng3817<=ng29270;

 always  @(posedge pclk)
	ng316<=ng26883;

 always  @(posedge pclk)
	pg14167<=pg14147;

 always  @(posedge pclk)
	ng499<=ng25609;

 always  @(posedge pclk)
	pg17739<=pg14738;

 always  @(posedge pclk)
	pg8279<=ng25662;

 always  @(posedge pclk)
	ng2269<=ng33581;

 always  @(posedge pclk)
	ng2927<=ng34803;

 always  @(posedge pclk)
	ng577<=ng30334;

 always  @(posedge pclk)
	ng599<=ng33964;

 always  @(posedge pclk)
	pg8870<=pg8917;

 always  @(posedge pclk)
	ng781<=ng34600;

 always  @(posedge pclk)
	ng2759<=ng33608;

 always  @(posedge pclk)
	ng2715<=ng24263;

 always  @(posedge pclk)
	ng1870<=ng33980;

 always  @(posedge pclk)
	ng1768<=ng30353;

 always  @(posedge pclk)
	ng4031<=pg16748;

 always  @(posedge pclk)
	ng6181<=ng29302;

 always  @(posedge pclk)
	ng2173<=ng33996;

 always  @(posedge pclk)
	ng1783<=ng32992;

 always  @(posedge pclk)
	ng106<=ng26889;

 always  @(posedge pclk)
	ng2803<=ng34445;

 always  @(posedge pclk)
	ng6303<=ng30537;

 always  @(posedge pclk)
	ng3462<=ng25670;

 always  @(posedge pclk)
	ng482<=ng28044;

 always  @(posedge pclk)
	ng1811<=ng29242;

 always  @(posedge pclk)
	ng2890<=ng34799;

 always  @(posedge pclk)
	ng1542<=ng30346;

 always  @(posedge pclk)
	ng111<=pg33079;

 always  @(posedge pclk)
	ng2161<=ng33994;

 always  @(posedge pclk)
	ng947<=ng34601;

 always  @(posedge pclk)
	ng546<=ng34722;

 always  @(posedge pclk)
	ng3913<=ng30454;

 always  @(posedge pclk)
	pg12923<=ng24258;

 always  @(posedge pclk)
	pg8915<=pg11770;

 always  @(posedge pclk)
	ng5599<=ng30492;

 always  @(posedge pclk)
	ng3893<=ng30437;

 always  @(posedge pclk)
	ng4141<=ng25687;

 always  @(posedge pclk)
	ng3106<=ng29257;

 always  @(posedge pclk)
	ng3841<=ng25682;

 always  @(posedge pclk)
	ng2004<=ng33987;

 always  @(posedge pclk)
	ng3586<=ng30424;

 always  @(posedge pclk)
	ng939<=ng34727;

 always  @(posedge pclk)
	ng6195<=ng29303;

 always  @(posedge pclk)
	ng925<=ng32981;

 always  @(posedge pclk)
	ng6255<=ng30526;

 always  @(posedge pclk)
	ng2177<=ng33997;

 always  @(posedge pclk)
	ng5835<=ng29296;

 always  @(posedge pclk)
	ng4543<=ng33042;

 always  @(posedge pclk)
	ng5802<=pg9617;

 always  @(posedge pclk)
	ng5092<=ng25697;

 always  @(posedge pclk)
	ng3933<=ng30444;

 always  @(posedge pclk)
	pg17715<=pg14673;

 always  @(posedge pclk)
	ng911<=ng29230;

 always  @(posedge pclk)
	ng3901<=ng30438;

 always  @(posedge pclk)
	ng4297<=pg10122;

 always  @(posedge pclk)
	pg8475<=pg7946;

 always  @(posedge pclk)
	ng4049<=ng24278;

 always  @(posedge pclk)
	ng3139<=ng25654;

 always  @(posedge pclk)
	pg13881<=pg16924;

 always  @(posedge pclk)
	ng6649<=ng30558;

 always  @(posedge pclk)
	ng2599<=ng33601;

 always  @(posedge pclk)
	ng4087<=ng29275;

 always  @(posedge pclk)
	ng1467<=ng29237;

 always  @(posedge pclk)
	ng6519<=ng29306;

 always  @(posedge pclk)
	ng1700<=ng30350;

 always  @(posedge pclk)
	ng1950<=ng33985;

 always  @(posedge pclk)
	pg13926<=pg11388;

 always  @(posedge pclk)
	ng2417<=ng30377;

 always  @(posedge pclk)
	ng475<=ng24208;

 always  @(posedge pclk)
	ng333<=ng26884;

 always  @(posedge pclk)
	pg9553<=ng25701;

 always  @(posedge pclk)
	pg12422<=ng24348;

 always  @(posedge pclk)
	ng1779<=ng33559;

 always  @(posedge pclk)
	ng2834<=ng30392;

 always  @(posedge pclk)
	ng3470<=ng25667;

 always  @(posedge pclk)
	ng5188<=ng33050;

 always  @(posedge pclk)
	pg13259<=pg19334;

 always  @(posedge pclk)
	ng504<=ng25610;

 always  @(posedge pclk)
	ng6541<=ng29309;

 always  @(posedge pclk)
	ng6209<=ng33062;

 always  @(posedge pclk)
	ng5685<=pg17678;

 always  @(posedge pclk)
	pg7916<=ng24240;

 always  @(posedge pclk)
	ng3466<=ng29264;

 always  @(posedge pclk)
	ng3333<=ng28063;

 always  @(posedge pclk)
	ng4922<=ng34639;

 always  @(posedge pclk)
	ng6613<=ng30549;

 always  @(posedge pclk)
	ng93<=ng31783;

 always  @(posedge pclk)
	pg12368<=ng23280;

 always  @(posedge pclk)
	pg17787<=pg13039;

 always  @(posedge pclk)
	ng1478<=ng26924;

 always  @(posedge pclk)
	ng63<=ng29730;

 always  @(posedge pclk)
	ng2643<=ng34020;

 always  @(posedge pclk)
	ng191<=pg8358;

 always  @(posedge pclk)
	ng1620<=ng33970;

 always  @(posedge pclk)
	pg16924<=pg14451;

 always  @(posedge pclk)
	ng2495<=ng33594;

 always  @(posedge pclk)
	ng5583<=ng30488;

 always  @(posedge pclk)
	ng2138<=ng34604;

 always  @(posedge pclk)
	ng5244<=ng30469;

 always  @(posedge pclk)
	ng936<=ng26912;

 always  @(posedge pclk)
	ng429<=ng24204;

 always  @(posedge pclk)
	ng4854<=ng34467;

 always  @(posedge pclk)
	ng37<=ng34613;

 always  @(posedge pclk)
	ng6381<=ng24349;

 always  @(posedge pclk)
	ng347<=pg7540;

 always  @(posedge pclk)
	pg9019<=ng21898;

 always  @(posedge pclk)
	ng2767<=ng26927;

 always  @(posedge pclk)
	pg8788<=pg8787;

 always  @(posedge pclk)
	ng5921<=ng30507;

 always  @(posedge pclk)
	pg14673<=pg17819;

 always  @(posedge pclk)
	ng85<=pg33435;

 always  @(posedge pclk)
	ng5069<=ng28092;

 always  @(posedge pclk)
	ng1061<=ng26914;

 always  @(posedge pclk)
	ng4401<=ng26948;

 always  @(posedge pclk)
	pg14421<=pg16624;

 always  @(posedge pclk)
	ng3610<=ng30430;

 always  @(posedge pclk)
	ng4975<=ng34037;

 always  @(posedge pclk)
	ng4427<=ng26952;

 always  @(posedge pclk)
	ng4145<=ng26939;

 always  @(posedge pclk)
	ng1834<=ng30355;

 always  @(posedge pclk)
	ng5703<=ng33620;

 always  @(posedge pclk)
	pg10306<=ng34024;

 always  @(posedge pclk)
	ng1141<=ng29233;

 always  @(posedge pclk)
	ng4512<=ng33040;

 always  @(posedge pclk)
	ng4253<=ng34630;

 always  @(posedge pclk)
	ng4570<=ng33617;

 always  @(posedge pclk)
	ng1548<=ng24260;

 always  @(posedge pclk)
	ng4284<=ng21897;

 always  @(posedge pclk)
	ng385<=ng25598;

 always  @(posedge pclk)
	ng291<=ng32977;

 always  @(posedge pclk)
	pg17711<=pg14694;

 always  @(posedge pclk)
	ng3111<=ng25656;

 always  @(posedge pclk)
	ng718<=ng28051;

 always  @(posedge pclk)
	ng6267<=ng30528;

 always  @(posedge pclk)
	ng2399<=ng33588;

 always  @(posedge pclk)
	ng2898<=ng34795;

 always  @(posedge pclk)
	pg7257<=ng26946;

 always  @(posedge pclk)
	ng4831<=ng28099;

 always  @(posedge pclk)
	ng5889<=ng30502;

 always  @(posedge pclk)
	ng822<=ng26899;

 always  @(posedge pclk)
	ng43<=ng28140;

 always  @(posedge pclk)
	pg17649<=pg17760;

 always  @(posedge pclk)
	ng2112<=ng33573;

 always  @(posedge pclk)
	ng5543<=ng30481;

 always  @(posedge pclk)
	pg7260<=ng26955;

 always  @(posedge pclk)
	ng142<=ng34250;

 always  @(posedge pclk)
	ng5022<=ng25703;

 always  @(posedge pclk)
	ng6148<=pg9682;

 always  @(posedge pclk)
	ng1448<=ng26922;

 always  @(posedge pclk)
	ng3961<=ng30451;

 always  @(posedge pclk)
	ng1018<=ng30337;

 always  @(posedge pclk)
	ng5029<=ng31902;

 always  @(posedge pclk)
	ng513<=ng25611;

 always  @(posedge pclk)
	ng5109<=pg9497;

 always  @(posedge pclk)
	ng2016<=ng33989;

 always  @(posedge pclk)
	ng5575<=ng30486;

 always  @(posedge pclk)
	ng5052<=ng31903;

 always  @(posedge pclk)
	ng1992<=ng30362;

 always  @(posedge pclk)
	ng2902<=ng34801;

 always  @(posedge pclk)
	ng3808<=ng29269;

 always  @(posedge pclk)
	ng1608<=ng33967;

 always  @(posedge pclk)
	ng5535<=ng33055;

 always  @(posedge pclk)
	ng405<=ng24201;

 always  @(posedge pclk)
	pg8291<=ng25591;

 always  @(posedge pclk)
	pg9555<=ng25714;

 always  @(posedge pclk)
	ng3203<=ng30411;

 always  @(posedge pclk)
	ng655<=ng28050;

 always  @(posedge pclk)
	ng4423<=pg10306;

 always  @(posedge pclk)
	ng4633<=ng34458;

 always  @(posedge pclk)
	ng4116<=ng28072;

 always  @(posedge pclk)
	ng298<=ng33961;

 always  @(posedge pclk)
	pg17291<=ng24238;

 always  @(posedge pclk)
	ng4501<=ng33038;

 always  @(posedge pclk)
	ng6513<=ng25761;

 always  @(posedge pclk)
	ng5240<=ng30468;

 always  @(posedge pclk)
	ng1002<=ng28057;

 always  @(posedge pclk)
	ng896<=ng26910;

 always  @(posedge pclk)
	ng3451<=pg8279;

 always  @(posedge pclk)
	ng2712<=ng24266;

 always  @(posedge pclk)
	ng5929<=ng30509;

 always  @(posedge pclk)
	pg9743<=ng25756;

 always  @(posedge pclk)
	ng837<=ng24215;

 always  @(posedge pclk)
	ng2437<=ng34009;

 always  @(posedge pclk)
	pg17743<=pg14705;

 always  @(posedge pclk)
	pg16744<=pg13926;

 always  @(posedge pclk)
	ng785<=ng34725;

 always  @(posedge pclk)
	ng2575<=ng34017;

 always  @(posedge pclk)
	pg17871<=pg13099;

 always  @(posedge pclk)
	ng3925<=ng30442;

 always  @(posedge pclk)
	wire1457<=wire1421;

 always  @(posedge pclk)
	ng4765<=ng34264;

 always  @(posedge pclk)
	ng1266<=ng25630;

 always  @(posedge pclk)
	ng6605<=ng30562;

 always  @(posedge pclk)
	ng2868<=ng34616;

 always  @(posedge pclk)
	ng6573<=ng33070;

 always  @(posedge pclk)
	ng5485<=ng29289;

 always  @(posedge pclk)
	ng1211<=ng25628;

 always  @(posedge pclk)
	ng1821<=ng33555;

 always  @(posedge pclk)
	ng5124<=ng29281;

 always  @(posedge pclk)
	pg12470<=ng24352;

 always  @(posedge pclk)
	ng790<=ng34791;

 always  @(posedge pclk)
	ng5142<=ng29284;

 always  @(posedge pclk)
	ng3594<=ng30426;

 always  @(posedge pclk)
	ng5953<=ng30515;

 always  @(posedge pclk)
	pg14635<=pg17813;

 always  @(posedge pclk)
	ng6561<=ng33068;

 always  @(posedge pclk)
	ng2775<=ng34443;

 always  @(posedge pclk)
	ng4366<=ng26944;

 always  @(posedge pclk)
	ng5016<=ng31898;

 always  @(posedge pclk)
	pg13049<=pg17604;

 always  @(posedge pclk)
	ng5128<=ng25705;

 always  @(posedge pclk)
	ng5456<=pg9555;

 always  @(posedge pclk)
	ng4674<=ng34026;

 always  @(posedge pclk)
	ng4153<=ng30457;

 always  @(posedge pclk)
	ng117<=ng30390;

 always  @(posedge pclk)
	ng3239<=ng30404;

 always  @(posedge pclk)
	ng1437<=ng29236;

 always  @(posedge pclk)
	wire1421<=ng24627;

 always  @(posedge pclk)
	ng4269<=ng21895;

 always  @(posedge pclk)
	ng3343<=ng24269;

 always  @(posedge pclk)
	ng2819<=ng34448;

 always  @(posedge pclk)
	ng3050<=ng25650;

 always  @(posedge pclk)
	ng4495<=ng33036;

 always  @(posedge pclk)
	ng1070<=ng30341;

 always  @(posedge pclk)
	pg16775<=pg13966;

 always  @(posedge pclk)
	ng6251<=ng30540;

 always  @(posedge pclk)
	ng1283<=ng34730;

 always  @(posedge pclk)
	ng6537<=ng25763;

 always  @(posedge pclk)
	ng2932<=ng24282;

 always  @(posedge pclk)
	ng4584<=ng34451;

 always  @(posedge pclk)
	pg16955<=pg14518;

 always  @(posedge pclk)
	pg9680<=ng25729;

 always  @(posedge pclk)
	pg14125<=pg14096;

 always  @(posedge pclk)
	ng2984<=ng34980;

 always  @(posedge pclk)
	pg17320<=ng24254;

 always  @(posedge pclk)
	ng1256<=ng29235;

 always  @(posedge pclk)
	ng2841<=ng2837;

 always  @(posedge pclk)
	ng2307<=ng34003;

 always  @(posedge pclk)
	pg9615<=ng25715;

 always  @(posedge pclk)
	ng31<=ng33149;

 always  @(posedge pclk)
	ng4455<=ng4456;

 always  @(posedge pclk)
	ng9<=ng33197;

 always  @(posedge pclk)
	pg8785<=pg8784;

 always  @(posedge pclk)
	ng4950<=ng28089;

 always  @(posedge pclk)
	ng5216<=ng30463;

 always  @(posedge pclk)
	ng1936<=ng33562;

 always  @(posedge pclk)
	ng1668<=ng33546;

 always  @(posedge pclk)
	pg14662<=pg12238;

 always  @(posedge pclk)
	ng3689<=ng24272;

 always  @(posedge pclk)
	ng4146<=ng34628;

 always  @(posedge pclk)
	ng4681<=ng34027;

 always  @(posedge pclk)
	ng827<=ng28055;

 always  @(posedge pclk)
	ng287<=ng31865;

 always  @(posedge pclk)
	ng1277<=ng32985;

 always  @(posedge pclk)
	ng2799<=ng26931;

 always  @(posedge pclk)
	ng1945<=ng29244;

 always  @(posedge pclk)
	ng776<=ng34439;

 always  @(posedge pclk)
	ng358<=pg8719;

 always  @(posedge pclk)
	ng626<=ng34849;

 always  @(posedge pclk)
	ng4340<=ng34459;

 always  @(posedge pclk)
	ng2036<=ng30363;

 always  @(posedge pclk)
	ng1249<=ng24247;

 always  @(posedge pclk)
	ng2102<=ng30365;

 always  @(posedge pclk)
	ng6173<=ng29300;

 always  @(posedge pclk)
	ng2338<=ng33591;

 always  @(posedge pclk)
	ng6741<=ng33626;

 always  @(posedge pclk)
	ng65<=ng66;

 always  @(posedge pclk)
	pg17845<=pg13085;

 always  @(posedge pclk)
	ng6509<=ng29305;

 always  @(posedge pclk)
	ng2070<=ng33570;

 always  @(posedge pclk)
	ng5563<=ng30484;

 always  @(posedge pclk)
	ng4473<=ng34256;

 always  @(posedge pclk)
	ng2445<=ng34011;

 always  @(posedge pclk)
	ng2407<=ng33590;

 always  @(posedge pclk)
	ng1677<=ng29240;

 always  @(posedge pclk)
	ng86<=ng25699;

 always  @(posedge pclk)
	ng2827<=ng26934;

 always  @(posedge pclk)
	pg17400<=pg17316;

 always  @(posedge pclk)
	ng1306<=ng25636;

 always  @(posedge pclk)
	ng1514<=ng30344;

 always  @(posedge pclk)
	ng4727<=ng34633;

 always  @(posedge pclk)
	ng3219<=ng30399;

 always  @(posedge pclk)
	ng6597<=ng30561;

 always  @(posedge pclk)
	ng5913<=ng30520;

 always  @(posedge pclk)
	ng3259<=ng30409;

 always  @(posedge pclk)
	ng2999<=ng34805;

 always  @(posedge pclk)
	ng2472<=ng33599;

 always  @(posedge pclk)
	ng3195<=ng30410;

 always  @(posedge pclk)
	ng4417<=ng31895;

 always  @(posedge pclk)
	ng2922<=ng34619;

 always  @(posedge pclk)
	ng3401<=ng25664;

 always  @(posedge pclk)
	ng3119<=ng25653;

 always  @(posedge pclk)
	ng3211<=ng30412;

 always  @(posedge pclk)
	ng3821<=ng25681;

 always  @(posedge pclk)
	ng3191<=ng30395;

 always  @(posedge pclk)
	ng2527<=ng30380;

 always  @(posedge pclk)
	ng3243<=ng30405;

 always  @(posedge pclk)
	ng5204<=ng30476;

 always  @(posedge pclk)
	ng1862<=ng33560;

 always  @(posedge pclk)
	ng1178<=ng24236;

 always  @(posedge pclk)
	pg14779<=pg12422;

 always  @(posedge pclk)
	ng3530<=ng33029;

 always  @(posedge pclk)
	ng4273<=ng24280;

 always  @(posedge pclk)
	ng4572<=ng28626;

 always  @(posedge pclk)
	ng2259<=ng30370;

 always  @(posedge pclk)
	ng6191<=ng25749;

 always  @(posedge pclk)
	ng6307<=ng30538;

 always  @(posedge pclk)
	ng4281<=pg8839;

 always  @(posedge pclk)
	ng4639<=ng34025;

 always  @(posedge pclk)
	ng5037<=ng31899;

 always  @(posedge pclk)
	ng6279<=ng30531;

 always  @(posedge pclk)
	ng5297<=ng33619;

 always  @(posedge pclk)
	pg8916<=pg8915;

 always  @(posedge pclk)
	ng232<=ng26903;

 always  @(posedge pclk)
	ng3498<=ng29268;

 always  @(posedge pclk)
	ng6555<=ng33067;

 always  @(posedge pclk)
	ng1472<=ng26923;

 always  @(posedge pclk)
	ng4760<=ng28085;

 always  @(posedge pclk)
	ng2204<=ng33583;

 always  @(posedge pclk)
	ng862<=ng26909;

 always  @(posedge pclk)
	ng6736<=ng24355;

 always  @(posedge pclk)
	ng6500<=ng29304;

 always  @(posedge pclk)
	ng2724<=ng26926;

 always  @(posedge pclk)
	ng2882<=ng34796;

 always  @(posedge pclk)
	ng2541<=ng33598;

 always  @(posedge pclk)
	ng6653<=ng30559;

 always  @(posedge pclk)
	ng4894<=ng28087;

 always  @(posedge pclk)
	ng2476<=ng33012;

 always  @(posedge pclk)
	ng2729<=ng28060;

 always  @(posedge pclk)
	pg16874<=pg14421;

 always  @(posedge pclk)
	ng930<=ng33540;

 always  @(posedge pclk)
	ng6682<=ng33627;

 always  @(posedge pclk)
	ng2873<=ng34615;

 always  @(posedge pclk)
	ng4899<=ng34040;

 always  @(posedge pclk)
	pg8919<=pg8918;

 always  @(posedge pclk)
	ng3484<=ng29267;

 always  @(posedge pclk)
	ng604<=ng34251;

 always  @(posedge pclk)
	ng1825<=ng29243;

 always  @(posedge pclk)
	ng4392<=ng26950;

 always  @(posedge pclk)
	ng4520<=ng4519;

 always  @(posedge pclk)
	ng1395<=ng25634;

 always  @(posedge pclk)
	ng714<=ng29227;

 always  @(posedge pclk)
	ng79<=ng26896;

 always  @(posedge pclk)
	ng6505<=ng25764;

 always  @(posedge pclk)
	ng5462<=ng29286;

 always  @(posedge pclk)
	ng5073<=ng28091;

 always  @(posedge pclk)
	ng1636<=ng33545;

 always  @(posedge pclk)
	ng5849<=ng29297;

 always  @(posedge pclk)
	ng2197<=ng33577;

 always  @(posedge pclk)
	ng1858<=ng30357;

 always  @(posedge pclk)
	ng6581<=ng30544;

 always  @(posedge pclk)
	ng1902<=ng30358;

 always  @(posedge pclk)
	ng2126<=ng30367;

 always  @(posedge pclk)
	pg8786<=pg8785;

 always  @(posedge pclk)
	ng582<=ng31866;

 always  @(posedge pclk)
	ng3845<=ng25683;

 always  @(posedge pclk)
	ng2079<=ng29246;

 always  @(posedge pclk)
	ng5841<=ng25734;

 always  @(posedge pclk)
	ng4239<=ng21892;

 always  @(posedge pclk)
	ng5148<=ng25706;

 always  @(posedge pclk)
	pg17604<=pg17580;

 always  @(posedge pclk)
	pg17607<=pg17739;

 always  @(posedge pclk)
	pg17685<=pg17649;

 always  @(posedge pclk)
	ng128<=ng28093;

 always  @(posedge pclk)
	ng2610<=ng33016;

 always  @(posedge pclk)
	ng6727<=ng24353;

 always  @(posedge pclk)
	ng3143<=ng25655;

 always  @(posedge pclk)
	ng4927<=ng34642;

 always  @(posedge pclk)
	ng5077<=ng25704;

 always  @(posedge pclk)
	ng2342<=ng33008;

 always  @(posedge pclk)
	ng3574<=ng30421;

 always  @(posedge pclk)
	ng2319<=ng33007;

 always  @(posedge pclk)
	ng5752<=ng25730;

 always  @(posedge pclk)
	ng1041<=ng25624;

 always  @(posedge pclk)
	ng4467<=ng34255;

 always  @(posedge pclk)
	ng2279<=ng30371;

 always  @(posedge pclk)
	pg14189<=ng26900;

 always  @(posedge pclk)
	ng2606<=ng33607;

 always  @(posedge pclk)
	ng262<=ng26904;

 always  @(posedge pclk)
	ng3502<=ng34626;

 always  @(posedge pclk)
	ng5817<=ng29293;

 always  @(posedge pclk)
	ng4944<=ng34268;

 always  @(posedge pclk)
	ng3827<=ng29271;

 always  @(posedge pclk)
	ng4704<=ng28083;

 always  @(posedge pclk)
	ng336<=ng26886;

 always  @(posedge pclk)
	ng2153<=ng33576;

 always  @(posedge pclk)
	ng3480<=ng29266;

 always  @(posedge pclk)
	pg17678<=pg14635;

 always  @(posedge pclk)
	ng4646<=ng34260;

 always  @(posedge pclk)
	ng5357<=ng33618;

 always  @(posedge pclk)
	ng4907<=ng34640;

 always  @(posedge pclk)
	ng3937<=ng30445;

 always  @(posedge pclk)
	ng5949<=ng30514;

 always  @(posedge pclk)
	ng1854<=ng30356;

 always  @(posedge pclk)
	ng4064<=ng25685;

 always  @(posedge pclk)
	ng6247<=ng30525;

 always  @(posedge pclk)
	ng1259<=ng30342;

 always  @(posedge pclk)
	ng6589<=ng30560;

 always  @(posedge pclk)
	ng1322<=pg13272;

 always  @(posedge pclk)
	ng1913<=ng33567;

 always  @(posedge pclk)
	ng5489<=ng29290;

 always  @(posedge pclk)
	ng182<=ng25602;

 always  @(posedge pclk)
	ng1592<=ng33544;

 always  @(posedge pclk)
	ng2689<=ng34606;

 always  @(posedge pclk)
	pg14217<=pg14201;

 always  @(posedge pclk)
	ng2509<=ng34013;

 always  @(posedge pclk)
	ng3921<=ng30441;

 always  @(posedge pclk)
	ng1756<=ng33977;

 always  @(posedge pclk)
	ng2950<=ng34621;

 always  @(posedge pclk)
	ng446<=ng26908;

 always  @(posedge pclk)
	ng4349<=ng34257;

 always  @(posedge pclk)
	ng6163<=ng29299;

 always  @(posedge pclk)
	ng5248<=ng30470;

 always  @(posedge pclk)
	pg7245<=ng26954;

 always  @(posedge pclk)
	pg11447<=ng21901;

 always  @(posedge pclk)
	ng2116<=ng33574;

 always  @(posedge pclk)
	ng2697<=ng34607;

 always  @(posedge pclk)
	pg16722<=pg13881;

 always  @(posedge pclk)
	ng2453<=ng33011;

 always  @(posedge pclk)
	ng4420<=ng26965;

 always  @(posedge pclk)
	ng3606<=ng30429;

 always  @(posedge pclk)
	ng843<=ng25619;

 always  @(posedge pclk)
	ng3506<=ng30414;

 always  @(posedge pclk)
	ng1036<=ng33541;

 always  @(posedge pclk)
	ng4104<=ng33615;

 always  @(posedge pclk)
	ng1706<=ng33548;

 always  @(posedge pclk)
	ng5523<=ng33053;

 always  @(posedge pclk)
	ng6159<=ng25750;

 always  @(posedge pclk)
	ng2960<=ng34622;

 always  @(posedge pclk)
	ng5495<=ng25720;

 always  @(posedge pclk)
	ng2975<=ng34804;

 always  @(posedge pclk)
	ng6549<=ng30543;

 always  @(posedge pclk)
	ng2315<=ng34005;

 always  @(posedge pclk)
	ng2595<=ng30383;

 always  @(posedge pclk)
	ng6545<=ng34647;

 always  @(posedge pclk)
	ng2652<=ng29255;

 always  @(posedge pclk)
	ng6235<=ng30523;

 always  @(posedge pclk)
	ng542<=ng24211;

 always  @(posedge pclk)
	ng1840<=ng33556;

 always  @(posedge pclk)
	ng703<=ng24214;

 always  @(posedge pclk)
	pg9497<=ng25700;

 always  @(posedge pclk)
	ng4072<=ng25691;

 always  @(posedge pclk)
	ng3133<=ng29261;

 always  @(posedge pclk)
	ng22<=ng27511;

 always  @(posedge pclk)
	ng1906<=ng33561;

 always  @(posedge pclk)
	ng4912<=ng34641;

 always  @(posedge pclk)
	ng1959<=ng29245;

 always  @(posedge pclk)
	ng3857<=ng30435;

 always  @(posedge pclk)
	ng2375<=ng34006;

 always  @(posedge pclk)
	ng4991<=ng34038;

 always  @(posedge pclk)
	ng2946<=ng21899;

 always  @(posedge pclk)
	ng2831<=ng30391;

 always  @(posedge pclk)
	ng739<=ng29228;

 always  @(posedge pclk)
	ng5084<=ng25696;

 always  @(posedge pclk)
	ng4785<=ng34029;

 always  @(posedge pclk)
	ng2791<=ng26929;

 always  @(posedge pclk)
	ng6609<=ng30548;

 always  @(posedge pclk)
	ng2098<=ng30364;

 always  @(posedge pclk)
	ng3546<=ng30431;

 always  @(posedge pclk)
	ng2185<=ng33003;

 always  @(posedge pclk)
	ng2491<=ng33014;

 always  @(posedge pclk)
	ng1312<=ng25631;

 always  @(posedge pclk)
	ng1129<=ng26916;

 always  @(posedge pclk)
	ng1221<=ng24246;

 always  @(posedge pclk)
	ng1624<=ng32987;

 always  @(posedge pclk)
	ng1848<=ng33558;

 always  @(posedge pclk)
	ng4859<=ng34468;

 always  @(posedge pclk)
	wire1411<=wire1457;

 always  @(posedge pclk)
	ng2994<=ng34732;

 always  @(posedge pclk)
	ng956<=ng25626;

 always  @(posedge pclk)
	ng2421<=ng33592;

 always  @(posedge pclk)
	ng6533<=ng25762;

 always  @(posedge pclk)
	ng370<=ng25597;

 always  @(posedge pclk)
	ng1874<=ng33986;

 always  @(posedge pclk)
	ng4125<=ng25690;

 always  @(posedge pclk)
	ng5481<=ng29288;

 always  @(posedge pclk)
	ng7<=ng33212;

 always  @(posedge pclk)
	ng2361<=ng33586;

 always  @(posedge pclk)
	ng2327<=ng30373;

 always  @(posedge pclk)
	ng723<=ng29229;

 always  @(posedge pclk)
	ng94<=ng34614;

 always  @(posedge pclk)
	ng3703<=ng33611;

 always  @(posedge pclk)
	ng4549<=ng33041;

 always  @(posedge pclk)
	ng4180<=pg8789;

 always  @(posedge pclk)
	ng1926<=ng32997;

 always  @(posedge pclk)
	ng676<=ng29226;

 always  @(posedge pclk)
	ng4558<=ng26966;

 always  @(posedge pclk)
	ng4864<=ng34034;

 always  @(posedge pclk)
	ng1532<=ng24253;

 always  @(posedge pclk)
	ng1389<=ng26920;

 always  @(posedge pclk)
	pg16627<=pg16744;

 always  @(posedge pclk)
	ng3802<=pg8344;

 always  @(posedge pclk)
	ng2255<=ng30369;

 always  @(posedge pclk)
	ng5499<=ng25721;

 always  @(posedge pclk)
	pg11770<=ng21891;

 always  @(posedge pclk)
	ng5917<=ng30506;

 always  @(posedge pclk)
	ng6167<=ng25747;

 always  @(posedge pclk)
	ng3917<=ng30440;

 always  @(posedge pclk)
	ng2537<=ng33597;

 always  @(posedge pclk)
	ng5268<=ng30475;

 always  @(posedge pclk)
	ng3881<=ng33034;

 always  @(posedge pclk)
	ng5256<=ng30472;

 always  @(posedge pclk)
	ng4732<=ng34634;

 always  @(posedge pclk)
	pg7540<=ng26890;

 always  @(posedge pclk)
	pg17813<=pg13049;

 always  @(posedge pclk)
	ng2878<=ng34797;

 always  @(posedge pclk)
	ng933<=ng32982;

 always  @(posedge pclk)
	ng4157<=ng34629;

 always  @(posedge pclk)
	ng3863<=ng33031;

 always  @(posedge pclk)
	pg16693<=pg16659;

 always  @(posedge pclk)
	ng1657<=ng32989;

 always  @(posedge pclk)
	pg17819<=pg13068;

 always  @(posedge pclk)
	ng4035<=ng28069;

 always  @(posedge pclk)
	ng667<=ng25615;

 always  @(posedge pclk)
	ng5475<=ng25719;

 always  @(posedge pclk)
	ng5603<=ng30493;

 always  @(posedge pclk)
	ng2719<=ng25639;

 always  @(posedge pclk)
	ng3949<=ng30448;

 always  @(posedge pclk)
	ng209<=ng25593;

 always  @(posedge pclk)
	ng4462<=ng34254;

 always  @(posedge pclk)
	ng4249<=ng34631;

 always  @(posedge pclk)
	ng5236<=ng30467;

 always  @(posedge pclk)
	pg8917<=pg8916;

 always  @(posedge pclk)
	ng4849<=ng34465;

 always  @(posedge pclk)
	pg16718<=pg13895;

 always  @(posedge pclk)
	ng2227<=ng33578;

 always  @(posedge pclk)
	ng5062<=ng25702;

 always  @(posedge pclk)
	ng34<=ng34650;

 always  @(posedge pclk)
	ng424<=ng24202;

 always  @(posedge pclk)
	ng1280<=ng26919;

 always  @(posedge pclk)
	ng650<=ng28049;

 always  @(posedge pclk)
	ng2181<=ng33998;

 always  @(posedge pclk)
	ng1046<=ng26913;

 always  @(posedge pclk)
	ng1345<=ng28059;

 always  @(posedge pclk)
	ng5694<=ng24342;

 always  @(posedge pclk)
	ng2441<=ng34010;

 always  @(posedge pclk)
	ng4821<=ng28096;

 always  @(posedge pclk)
	ng3694<=ng24273;

 always  @(posedge pclk)
	ng2779<=ng26928;

 always  @(posedge pclk)
	ng376<=ng25596;

 always  @(posedge pclk)
	ng907<=ng28056;

 always  @(posedge pclk)
	ng699<=ng28053;

 always  @(posedge pclk)
	ng3129<=ng29260;

 always  @(posedge pclk)
	ng4698<=ng34261;

 always  @(posedge pclk)
	ng6035<=ng24345;

 always  @(posedge pclk)
	ng4507<=ng30458;

 always  @(posedge pclk)
	ng4040<=ng24276;

 always  @(posedge pclk)
	ng5555<=ng30483;

 always  @(posedge pclk)
	ng590<=ng32978;

 always  @(posedge pclk)
	ng1752<=ng33976;

 always  @(posedge pclk)
	ng4477<=ng4474;

 always  @(posedge pclk)
	ng1296<=ng34729;

 always  @(posedge pclk)
	ng4382<=ng26947;

 always  @(posedge pclk)
	ng1052<=ng25625;

 always  @(posedge pclk)
	ng1728<=ng33552;

 always  @(posedge pclk)
	ng969<=ng25622;

 always  @(posedge pclk)
	ng355<=ng26892;

 always  @(posedge pclk)
	pg17639<=pg14597;

 always  @(posedge pclk)
	pg9817<=ng25757;

 always  @(posedge pclk)
	ng225<=ng26901;

 always  @(posedge pclk)
	ng5869<=ng33058;

 always  @(posedge pclk)
	ng153<=ng33534;

 always  @(posedge pclk)
	ng2811<=ng26932;

 always  @(posedge pclk)
	ng1585<=pg12923;

 always  @(posedge pclk)
	ng4108<=ng33035;

 always  @(posedge pclk)
	ng5881<=ng33060;

 always  @(posedge pclk)
	ng1146<=ng24233;

 always  @(posedge pclk)
	ng518<=ng25612;

 always  @(posedge pclk)
	ng4531<=ng24335;

 always  @(posedge pclk)
	ng5041<=ng31900;

 always  @(posedge pclk)
	ng2988<=ng34624;

 always  @(posedge pclk)
	ng1526<=ng30345;

 always  @(posedge pclk)
	ng568<=ng26895;

 always  @(posedge pclk)
	pg10122<=ng21900;

 always  @(posedge pclk)
	ng4546<=ng33045;

 always  @(posedge pclk)
	ng6098<=ng25744;

 always  @(posedge pclk)
	ng6283<=ng30532;

 always  @(posedge pclk)
	ng5120<=ng25708;

 always  @(posedge pclk)
	pg19357<=ng24257;

 always  @(posedge pclk)
	ng4322<=ng34450;

 always  @(posedge pclk)
	ng5252<=ng30471;

 always  @(posedge pclk)
	ng1274<=ng33542;

 always  @(posedge pclk)
	ng112<=ng30605;

 always  @(posedge pclk)
	ng5033<=ng31904;

 always  @(posedge pclk)
	ng4939<=ng28088;

 always  @(posedge pclk)
	ng5097<=ng25698;

 always  @(posedge pclk)
	ng5112<=pg9553;

 always  @(posedge pclk)
	ng3329<=pg16686;

 always  @(posedge pclk)
	ng943<=ng34728;

 always  @(posedge pclk)
	ng5200<=ng30461;

 always  @(posedge pclk)
	ng2912<=ng34618;

 always  @(posedge pclk)
	ng3352<=ng33609;

 always  @(posedge pclk)
	ng3125<=ng29259;

 always  @(posedge pclk)
	ng1988<=ng30361;

 always  @(posedge pclk)
	ng5348<=ng24338;

 always  @(posedge pclk)
	pg12832<=ng26958;

 always  @(posedge pclk)
	ng1878<=ng33981;

 always  @(posedge pclk)
	ng2547<=ng30381;

 always  @(posedge pclk)
	ng5343<=ng24337;

 always  @(posedge pclk)
	pg13099<=pg17722;

 always  @(posedge pclk)
	ng5567<=ng30499;

 always  @(posedge pclk)
	pg10500<=ng24239;

 always  @(posedge pclk)
	ng753<=ng26897;

 always  @(posedge pclk)
	ng351<=ng26891;

 always  @(posedge pclk)
	ng3179<=ng33024;

 always  @(posedge pclk)
	ng2807<=ng34447;

 always  @(posedge pclk)
	ng1682<=ng33971;

 always  @(posedge pclk)
	ng5831<=ng29295;

 always  @(posedge pclk)
	ng3231<=ng30402;

 always  @(posedge pclk)
	ng4486<=ng26961;

 always  @(posedge pclk)
	ng5579<=ng30487;

 always  @(posedge pclk)
	ng6625<=ng30552;

 always  @(posedge pclk)
	pg8398<=ng25677;

 always  @(posedge pclk)
	ng4388<=ng26949;

 always  @(posedge pclk)
	ng4564<=ng26967;

 always  @(posedge pclk)
	ng4308<=pg9251;

 always  @(posedge pclk)
	ng2625<=ng33018;

 always  @(posedge pclk)
	ng3897<=ng30452;

 always  @(posedge pclk)
	ng2860<=ng34611;

 always  @(posedge pclk)
	ng6641<=ng30556;

 always  @(posedge pclk)
	ng3538<=ng30415;

 always  @(posedge pclk)
	ng6523<=ng29307;

 always  @(posedge pclk)
	ng3263<=ng30413;

 always  @(posedge pclk)
	ng3562<=ng30433;

 always  @(posedge pclk)
	pg14828<=pg12470;

 always  @(posedge pclk)
	ng5937<=ng30511;

 always  @(posedge pclk)
	ng1242<=pg12919;

 always  @(posedge pclk)
	ng4771<=ng28086;

 always  @(posedge pclk)
	pg14705<=pg17845;

 always  @(posedge pclk)
	ng4966<=ng34039;

 always  @(posedge pclk)
	pg17674<=pg14662;

 always  @(posedge pclk)
	ng1199<=ng30340;

 always  @(posedge pclk)
	ng5941<=ng30512;

 always  @(posedge pclk)
	ng1152<=ng24234;

 always  @(posedge pclk)
	pg13085<=pg17685;

 always  @(posedge pclk)
	ng2856<=ng34793;

 always  @(posedge pclk)
	ng4818<=wire1411;

 always  @(posedge pclk)
	pg19334<=ng24241;

 always  @(posedge pclk)
	ng1964<=ng30359;

 always  @(posedge pclk)
	ng19<=ng33176;

 always  @(posedge pclk)
	ng5170<=ng33047;

 always  @(posedge pclk)
	ng1559<=ng25638;

 always  @(posedge pclk)
	ng4843<=ng34466;

 always  @(posedge pclk)
	pg14694<=pg12300;

 always  @(posedge pclk)
	ng6657<=ng30563;

 always  @(posedge pclk)
	ng2894<=ng34612;

 always  @(posedge pclk)
	ng4311<=ng34449;

 always  @(posedge pclk)
	ng3223<=ng30400;

 always  @(posedge pclk)
	ng3251<=ng30407;

 always  @(posedge pclk)
	ng5619<=ng30500;

 always  @(posedge pclk)
	ng559<=pg9048;

 always  @(posedge pclk)
	ng554<=ng34911;

 always  @(posedge pclk)
	ng1798<=ng32994;

 always  @(posedge pclk)
	ng4871<=ng34035;

 always  @(posedge pclk)
	ng1579<=pg10527;

 always  @(posedge pclk)
	ng4643<=ng34259;

 always  @(posedge pclk)
	ng2980<=ng34800;

 always  @(posedge pclk)
	ng5901<=ng30504;

 always  @(posedge pclk)
	ng479<=ng24210;

 always  @(posedge pclk)
	ng4653<=ng34462;

 always  @(posedge pclk)
	ng1105<=ng26915;

 always  @(posedge pclk)
	ng3889<=ng30436;

 always  @(posedge pclk)
	ng4098<=ng31894;

 always  @(posedge pclk)
	ng4504<=ng33039;

 always  @(posedge pclk)
	ng1589<=ng24261;

 always  @(posedge pclk)
	ng5990<=ng33623;

 always  @(posedge pclk)
	ng6275<=ng30530;

 always  @(posedge pclk)
	ng6239<=ng30524;

 always  @(posedge pclk)
	ng4571<=ng4570;

 always  @(posedge pclk)
	ng5406<=ng25716;

 always  @(posedge pclk)
	ng150<=ng32976;

 always  @(posedge pclk)
	ng538<=ng34719;

 always  @(posedge pclk)
	ng4743<=ng34262;

 always  @(posedge pclk)
	ng5571<=ng30485;

 always  @(posedge pclk)
	ng5196<=ng30460;

 always  @(posedge pclk)
	ng2351<=ng33009;

 always  @(posedge pclk)
	ng4434<=ng26956;

 always  @(posedge pclk)
	ng301<=ng33536;

 always  @(posedge pclk)
	ng854<=ng32980;

 always  @(posedge pclk)
	ng2518<=ng29253;

 always  @(posedge pclk)
	pg17646<=pg17607;

 always  @(posedge pclk)
	pg17764<=pg14749;

 always  @(posedge pclk)
	ng1236<=pg10500;

 always  @(posedge pclk)
	ng4616<=ng34456;

 always  @(posedge pclk)
	ng2523<=ng30379;

 always  @(posedge pclk)
	ng2551<=ng30382;

 always  @(posedge pclk)
	pg14749<=pg17871;

 always  @(posedge pclk)
	ng2579<=ng34018;

 always  @(posedge pclk)
	pg17519<=pg17674;

 always  @(posedge pclk)
	ng3929<=ng30443;

 always  @(posedge pclk)
	ng2012<=ng33988;

 always  @(posedge pclk)
	ng4836<=ng34265;

 always  @(posedge pclk)
	ng2108<=ng33572;

 always  @(posedge pclk)
	ng2571<=ng34016;

 always  @(posedge pclk)
	ng2093<=ng29247;

 always  @(posedge pclk)
	ng1554<=ng25637;

 always  @(posedge pclk)
	ng3207<=ng30397;

 always  @(posedge pclk)
	pg16748<=pg13906;

 always  @(posedge pclk)
	ng1720<=ng30351;

 always  @(posedge pclk)
	ng1193<=ng26918;

 always  @(posedge pclk)
	ng3255<=ng30408;

 always  @(posedge pclk)
	ng5893<=ng30503;

 always  @(posedge pclk)
	ng4456<=ng24298;

 always  @(posedge pclk)
	pg9682<=ng25742;

 always  @(posedge pclk)
	ng1300<=ng25635;

 always  @(posedge pclk)
	ng4552<=ng33044;

 always  @(posedge pclk)
	ng3187<=ng30394;

 always  @(posedge pclk)
	ng1996<=ng33568;

 always  @(posedge pclk)
	pg11388<=ng24271;

 always  @(posedge pclk)
	ng496<=ng33963;

 always  @(posedge pclk)
	pg14096<=pg14217;

 always  @(posedge pclk)
	ng4722<=ng34636;

 always  @(posedge pclk)
	ng6154<=ng29298;

 always  @(posedge pclk)
	ng5264<=ng30474;

 always  @(posedge pclk)
	ng3151<=ng34625;

 always  @(posedge pclk)
	ng2886<=ng34798;

 always  @(posedge pclk)
	ng6386<=ng24350;

 always  @(posedge pclk)
	ng4054<=ng33613;

 always  @(posedge pclk)
	ng1087<=pg17400;

 always  @(posedge pclk)
	ng3476<=ng29265;

 always  @(posedge pclk)
	ng4575<=ng29276;

 always  @(posedge pclk)
	ng5873<=ng33059;

 always  @(posedge pclk)
	ng4578<=ng29278;

 always  @(posedge pclk)
	ng4459<=ng34253;

 always  @(posedge pclk)
	ng6311<=ng30542;

 always  @(posedge pclk)
	ng4826<=ng28102;

 always  @(posedge pclk)
	pg13895<=pg11349;

 always  @(posedge pclk)
	ng3338<=ng24268;

 always  @(posedge pclk)
	ng1696<=ng30349;

 always  @(posedge pclk)
	ng6<=ng33219;

 always  @(posedge pclk)
	ng3578<=ng30422;

 always  @(posedge pclk)
	ng2380<=ng33587;

 always  @(posedge pclk)
	ng2648<=ng33603;

 always  @(posedge pclk)
	ng341<=ng26888;

 always  @(posedge pclk)
	ng4601<=ng34453;

 always  @(posedge pclk)
	ng2567<=ng34021;

 always  @(posedge pclk)
	ng890<=ng34440;

 always  @(posedge pclk)
	ng2864<=ng34794;

 always  @(posedge pclk)
	ng28<=ng33164;

 always  @(posedge pclk)
	ng4561<=ng26968;

 always  @(posedge pclk)
	ng5156<=ng29285;

 always  @(posedge pclk)
	ng2273<=ng33582;

 always  @(posedge pclk)
	ng904<=ng24231;

 always  @(posedge pclk)
	ng6227<=ng33065;

 always  @(posedge pclk)
	ng6203<=ng30522;

 always  @(posedge pclk)
	ng66<=ng24334;

 always  @(posedge pclk)
	pg13068<=pg17646;

 always  @(posedge pclk)
	ng2165<=ng34000;

 always  @(posedge pclk)
	ng4112<=ng28071;

 always  @(posedge pclk)
	ng1982<=ng33566;

 always  @(posedge pclk)
	ng4717<=ng34635;

 always  @(posedge pclk)
	ng4483<=ng4520;

 always  @(posedge pclk)
	ng3215<=ng30398;

 always  @(posedge pclk)
	ng1367<=ng31871;

 always  @(posedge pclk)
	ng2051<=ng33000;

 always  @(posedge pclk)
	ng1691<=ng29241;

 always  @(posedge pclk)
	ng1111<=ng29234;

 always  @(posedge pclk)
	ng5821<=ng25733;

 always  @(posedge pclk)
	ng411<=ng29222;

 always  @(posedge pclk)
	ng4057<=ng25686;

 always  @(posedge pclk)
	pg16686<=pg13865;

 always  @(posedge pclk)
	ng2661<=ng30385;

 always  @(posedge pclk)
	ng2970<=ng34623;

 always  @(posedge pclk)
	ng4628<=ng34457;

 always  @(posedge pclk)
	ng2771<=ng34441;

 always  @(posedge pclk)
	ng3570<=ng30420;

 always  @(posedge pclk)
	ng622<=ng34790;

 always  @(posedge pclk)
	ng3853<=ng34627;

 always  @(posedge pclk)
	ng2941<=ng34806;

 always  @(posedge pclk)
	ng3100<=pg8215;

 always  @(posedge pclk)
	ng4737<=ng34637;

 always  @(posedge pclk)
	ng4754<=ng34263;

 always  @(posedge pclk)
	ng4983<=ng34041;

 always  @(posedge pclk)
	ng4961<=ng28090;

 always  @(posedge pclk)
	ng3494<=ng25669;

 always  @(posedge pclk)
	ng4749<=ng28084;

 always  @(posedge pclk)
	ng2465<=ng33593;

 always  @(posedge pclk)
	ng4917<=ng34638;

 always  @(posedge pclk)
	ng3680<=pg16722;

 always  @(posedge pclk)
	ng1748<=ng33975;

 always  @(posedge pclk)
	pg8215<=ng25648;

 always  @(posedge pclk)
	ng758<=ng32979;

 always  @(posedge pclk)
	pg12919<=ng24242;

 always  @(posedge pclk)
	ng1664<=ng32990;

 always  @(posedge pclk)
	ng528<=ng26894;

 always  @(posedge pclk)
	ng2848<=ng34792;

 always  @(posedge pclk)
	ng1564<=ng24262;

 always  @(posedge pclk)
	ng962<=ng25627;

 always  @(posedge pclk)
	ng3831<=ng29272;

 always  @(posedge pclk)
	ng4793<=ng34033;

 always  @(posedge pclk)
	ng5808<=ng29292;

 always  @(posedge pclk)
	pg17760<=pg14779;

 always  @(posedge pclk)
	ng1890<=ng33984;

 always  @(posedge pclk)
	pg12184<=ng24213;

 always  @(posedge pclk)
	ng5897<=ng30518;

 always  @(posedge pclk)
	pg14597<=pg17787;

 always  @(posedge pclk)
	ng4093<=ng30456;

 always  @(posedge pclk)
	ng2619<=ng33017;

 always  @(posedge pclk)
	ng661<=ng28052;

 always  @(posedge pclk)
	ng6494<=pg9743;

 always  @(posedge pclk)
	ng1413<=ng30347;

 always  @(posedge pclk)
	ng2311<=ng34004;

 always  @(posedge pclk)
	ng794<=ng34850;

 always  @(posedge pclk)
	ng2667<=ng33604;

 always  @(posedge pclk)
	ng2555<=ng33600;

 always  @(posedge pclk)
	ng4581<=ng26969;

 always  @(posedge pclk)
	ng1616<=ng33969;

 always  @(posedge pclk)
	ng305<=ng26880;

 always  @(posedge pclk)
	ng255<=ng26902;

 always  @(posedge pclk)
	ng613<=ng34599;

 always  @(posedge pclk)
	ng817<=ng25617;

 always  @(posedge pclk)
	ng686<=ng25614;

 always  @(posedge pclk)
	ng4489<=ng26962;

 always  @(posedge pclk)
	ng4955<=ng34269;

 always  @(posedge pclk)
	ng2675<=ng33606;

 always  @(posedge pclk)
	ng25<=ng25;

 always  @(posedge pclk)
	ng329<=ng319;

 always  @(posedge pclk)
	pg17722<=pg17688;

 always  @(posedge pclk)
	pg17778<=pg14828;

 always  @(posedge pclk)
	ng2533<=ng33596;

 always  @(posedge pclk)
	ng2936<=ng34620;

 always  @(posedge pclk)
	pg16603<=pg16718;

 always  @(posedge pclk)
	ng6299<=ng30536;

 always  @(posedge pclk)
	ng319<=ng26882;

 always  @(posedge pclk)
	ng1351<=ng25632;

 always  @(posedge pclk)
	pg16624<=pg16603;

 always  @(posedge pclk)
	ng728<=ng28054;

 always  @(posedge pclk)
	ng2084<=ng33992;

 always  @(posedge pclk)
	ng691<=ng28048;

 always  @(posedge pclk)
	ng5698<=ng24343;

 always  @(posedge pclk)
	ng4515<=ng26964;

 always  @(posedge pclk)
	ng1882<=ng33982;

 always  @(posedge pclk)
	pg9048<=pg12368;

 always  @(posedge pclk)
	ng6336<=ng33625;

 always  @(posedge pclk)
	ng5134<=ng29282;

 always  @(posedge pclk)
	ng4076<=ng28070;

 always  @(posedge pclk)
	ng1495<=ng24250;

 always  @(posedge pclk)
	pg16659<=pg16775;

 always  @(posedge pclk)
	ng5160<=ng34643;

 always  @(posedge pclk)
	ng1189<=ng24237;

 always  @(posedge pclk)
	ng437<=ng24206;

 always  @(posedge pclk)
	ng5511<=ng30480;

 always  @(posedge pclk)
	ng3965<=ng30455;

 always  @(posedge pclk)
	ng6187<=ng25748;

 always  @(posedge pclk)
	ng914<=ng30336;

 always  @(posedge pclk)
	ng5551<=ng30497;

 always  @(posedge pclk)
	ng1373<=ng32986;

 always  @(posedge pclk)
	ng632<=ng34880;

 always  @(posedge pclk)
	ng1246<=ng24245;

 always  @(posedge pclk)
	ng4498<=ng33037;

 always  @(posedge pclk)
	ng2241<=ng33999;

 always  @(posedge pclk)
	ng2370<=ng29250;

 always  @(posedge pclk)
	ng2756<=ng33019;

 always  @(posedge pclk)
	ng2514<=ng33595;

 always  @(posedge pclk)
	ng2763<=ng34022;

 always  @(posedge pclk)
	ng6645<=ng30557;

 always  @(posedge pclk)
	ng3869<=ng33032;

 always  @(posedge pclk)
	ng2629<=ng33602;

 always  @(posedge pclk)
	ng3639<=ng33612;

 always  @(posedge pclk)
	ng269<=ng26906;

 always  @(posedge pclk)
	ng3957<=ng30450;

 always  @(posedge pclk)
	ng1183<=ng30339;

 always  @(posedge pclk)
	ng4669<=ng34464;

 always  @(posedge pclk)
	ng4411<=pg7257;

 always  @(posedge pclk)
	ng3602<=ng30428;

 always  @(posedge pclk)
	ng4688<=ng34028;

 always  @(posedge pclk)
	ng3227<=ng30401;

 always  @(posedge pclk)
	pg13906<=pg16955;

 always  @(posedge pclk)
	ng2040<=ng33569;

 always  @(posedge pclk)
	ng5857<=ng30501;

 always  @(posedge pclk)
	ng8<=ng33204;

 always  @(posedge pclk)
	ng550<=ng34720;

 always  @(posedge pclk)
	ng283<=ng28043;

 always  @(posedge pclk)
	ng2795<=ng26930;

 always  @(posedge pclk)
	pg8358<=ng25592;

 always  @(posedge pclk)
	ng6049<=ng33622;

 always  @(posedge pclk)
	ng4082<=ng26938;

 always  @(posedge pclk)
	ng1252<=ng28058;

 always  @(posedge pclk)
	ng5527<=ng33054;

 always  @(posedge pclk)
	ng5224<=ng30464;

 always  @(posedge pclk)
	ng1287<=ng34731;

 always  @(posedge pclk)
	ng1644<=ng33551;

 always  @(posedge pclk)
	ng5176<=ng33048;

 always  @(posedge pclk)
	ng1536<=ng26925;

 always  @(posedge pclk)
	ng5228<=ng30465;

 always  @(posedge pclk)
	ng3849<=ng29274;

 always  @(posedge pclk)
	ng2303<=ng34002;

 always  @(posedge pclk)
	pg8277<=ng25649;

 always  @(posedge pclk)
	ng324<=ng26887;

 always  @(posedge pclk)
	ng6527<=ng29308;

 always  @(posedge pclk)
	ng5644<=ng33621;

 always  @(posedge pclk)
	pg8416<=pg7916;

 always  @(posedge pclk)
	ng3953<=ng30449;

 always  @(posedge pclk)
	ng164<=ng31864;

 always  @(posedge pclk)
	ng1648<=ng32988;

 always  @(posedge pclk)
	ng6295<=ng30535;

 always  @(posedge pclk)
	ng1792<=ng32993;

 always  @(posedge pclk)
	ng2583<=ng34019;

 always  @(posedge pclk)
	pg8342<=ng25663;

 always  @(posedge pclk)
	ng278<=ng25594;

 always  @(posedge pclk)
	ng6395<=ng33624;

 always  @(posedge pclk)
	pg17404<=pg17320;

 always  @(posedge pclk)
	ng763<=ng33539;

 always  @(posedge pclk)
	ng1632<=ng30348;

 always  @(posedge pclk)
	ng744<=ng30335;

 always  @(posedge pclk)
	ng1442<=ng24251;

 always  @(posedge pclk)
	ng1454<=ng29239;

 always  @(posedge pclk)
	ng2287<=ng33584;

 always  @(posedge pclk)
	ng3566<=ng30419;

 always  @(posedge pclk)
	ng681<=ng28047;

 always  @(posedge pclk)
	ng3518<=ng33027;

 always  @(posedge pclk)
	ng736<=pg11678;

 always  @(posedge pclk)
	pg17580<=pg17711;

 always  @(posedge pclk)
	ng3835<=ng29273;

 always  @(posedge pclk)
	ng5339<=pg17639;

 always  @(posedge pclk)
	ng174<=ng25601;

 always  @(posedge pclk)
	ng2783<=ng34442;

 always  @(posedge pclk)
	pg14738<=pg12350;

 always  @(posedge pclk)
	ng6243<=ng30539;

 always  @(posedge pclk)
	ng16<=ng33187;

 always  @(posedge pclk)
	ng239<=ng26905;

 always  @(posedge pclk)
	ng4452<=pg7245;

 always  @(posedge pclk)
	pg14147<=pg14125;

 always  @(posedge pclk)
	ng5164<=ng30459;

 always  @(posedge pclk)
	pg8918<=pg8870;

 always  @(posedge pclk)
	ng2461<=ng30378;

 always  @(posedge pclk)
	ng4369<=ng26970;

 always  @(posedge pclk)
	ng3288<=ng33610;

 always  @(posedge pclk)
	ng1263<=ng31870;

 always  @(posedge pclk)
	ng4664<=ng34463;

 always  @(posedge pclk)
	ng2047<=ng33575;

 always  @(posedge pclk)
	ng4430<=ng26957;

 always  @(posedge pclk)
	ng572<=ng28045;

 always  @(posedge pclk)
	ng3990<=ng33614;

 always  @(posedge pclk)
	ng812<=ng26898;

 always  @(posedge pclk)
	ng3684<=ng28066;

 always  @(posedge pclk)
	ng401<=ng24203;

 always  @(posedge pclk)
	ng586<=ng29224;

 always  @(posedge pclk)
	ng2393<=ng30375;

 always  @(posedge pclk)
	pg13039<=pg17577;

 always  @(posedge pclk)
	ng2587<=ng33015;

 always  @(posedge pclk)
	ng6271<=ng30529;

 always  @(posedge pclk)
	ng2020<=ng33990;

 always  @(posedge pclk)
	ng460<=ng25605;

 always  @(posedge pclk)
	ng3247<=ng30406;

 always  @(posedge pclk)
	pg8789<=pg8788;

 always  @(posedge pclk)
	ng199<=ng34721;

 always  @(posedge pclk)
	ng5080<=ng25695;

 always  @(posedge pclk)
	ng2965<=ng34808;

 always  @(posedge pclk)
	ng1404<=ng26921;

 always  @(posedge pclk)
	ng617<=ng34724;

 always  @(posedge pclk)
	ng3161<=ng33021;

 always  @(posedge pclk)
	ng1844<=ng33557;

 always  @(posedge pclk)
	ng1955<=ng33563;

 always  @(posedge pclk)
	ng671<=ng29225;

 always  @(posedge pclk)
	ng1270<=ng32984;

 always  @(posedge pclk)
	ng5925<=ng30508;

 always  @(posedge pclk)
	ng2787<=ng34444;

 always  @(posedge pclk)
	ng6601<=ng30547;

 always  @(posedge pclk)
	ng4119<=ng28073;

 always  @(posedge pclk)
	ng5845<=ng25735;

 always  @(posedge pclk)
	pg17688<=pg17778;

 always  @(posedge pclk)
	ng3550<=ng30417;

 always  @(posedge pclk)
	ng1687<=ng33547;

 always  @(posedge pclk)
	ng1710<=ng33549;

 always  @(posedge pclk)
	ng5152<=ng25707;

 always  @(posedge pclk)
	ng2060<=ng33001;

 always  @(posedge pclk)
	ng5046<=ng31901;

 always  @(posedge pclk)
	pg8920<=pg8919;

 always  @(posedge pclk)
	ng4519<=ng33616;

 always  @(posedge pclk)
	ng3614<=ng30434;

 always  @(posedge pclk)
	ng5272<=ng30479;

 always  @(posedge pclk)
	ng4358<=ng34258;

 always  @(posedge pclk)
	ng3003<=ng18597;

 always  @(posedge pclk)
	ng5260<=ng30473;

 always  @(posedge pclk)
	ng4300<=ng34735;

 always  @(posedge pclk)
	ng71<=ng16696;

 always  @(posedge pclk)
	ng2299<=ng34007;

 always  @(posedge pclk)
	ng4492<=ng26963;

 always  @(posedge pclk)
	pg8344<=ng25676;

 always  @(posedge pclk)
	ng3905<=ng30453;

 always  @(posedge pclk)
	pg12238<=ng24336;

 always  @(posedge pclk)
	ng1917<=ng32996;

 always  @(posedge pclk)
	ng5965<=ng30521;

 always  @(posedge pclk)
	ng5933<=ng30510;

 always  @(posedge pclk)
	ng5611<=ng30495;

 always  @(posedge pclk)
	ng4534<=ng34023;

 always  @(posedge pclk)
	ng417<=ng24209;

 always  @(posedge pclk)
	ng1604<=ng33972;

 always  @(posedge pclk)
	ng2008<=ng33993;

 always  @(posedge pclk)
	ng2122<=ng30366;

 always  @(posedge pclk)
	ng2433<=ng34014;

 always  @(posedge pclk)
	ng4164<=ng26940;

 always  @(posedge pclk)
	ng6637<=ng30555;

 always  @(posedge pclk)
	ng3558<=ng30418;

 always  @(posedge pclk)
	ng157<=ng33960;

 always  @(posedge pclk)
	pg13272<=pg19357;

 always  @(posedge pclk)
	ng5961<=ng30517;

 always  @(posedge pclk)
	ng6629<=ng30553;

 always  @(posedge pclk)
	ng1216<=ng25629;

 always  @(posedge pclk)
	ng1430<=pg17423;

 always  @(posedge pclk)
	ng5208<=ng30462;

 always  @(posedge pclk)
	ng1333<=pg8475;

 always  @(posedge pclk)
	ng101<=ng16663;

 always  @(posedge pclk)
	ng1816<=ng33978;

 always  @(posedge pclk)
	ng2403<=ng33589;

 always  @(posedge pclk)
	ng952<=ng34726;

 always  @(posedge pclk)
	ng2223<=ng33006;

 always  @(posedge pclk)
	ng5957<=ng30516;

 always  @(posedge pclk)
	pg8783<=pg11447;

 always  @(posedge pclk)
	ng2130<=ng34603;

 always  @(posedge pclk)
	ng832<=ng25618;

 always  @(posedge pclk)
	ng2823<=ng26933;

 always  @(posedge pclk)
	ng6040<=ng24346;

 always  @(posedge pclk)
	ng1760<=ng32991;

 always  @(posedge pclk)
	pg14201<=pg14189;

 always  @(posedge pclk)
	ng2193<=ng30368;

 always  @(posedge pclk)
	ng996<=ng24243;

 always  @(posedge pclk)
	ng4474<=ng4467;

 always  @(posedge pclk)
	ng4480<=ng31896;

 always  @(posedge pclk)
	ng3582<=ng30423;

 always  @(posedge pclk)
	pg14518<=pg16693;

 always  @(posedge pclk)
	ng5467<=ng25722;

 always  @(posedge pclk)
	ng4608<=ng34454;

 always  @(posedge pclk)
	ng1894<=ng32995;

 always  @(posedge pclk)
	ng5011<=ng28105;

 always  @(posedge pclk)
	ng5863<=ng33057;

 always  @(posedge pclk)
	ng6444<=ng25758;

 always  @(posedge pclk)
	ng5220<=ng30478;

 always  @(posedge pclk)
	ng2384<=ng29251;

 always  @(posedge pclk)
	ng4527<=ng28082;

 always  @(posedge pclk)
	ng1489<=ng24249;

 always  @(posedge pclk)
	pg8839<=ng21896;

 always  @(posedge pclk)
	ng3347<=ng24270;

 always  @(posedge pclk)
	ng2265<=ng33580;

 always  @(posedge pclk)
	ng1974<=ng33564;

 always  @(posedge pclk)
	ng1124<=ng29232;

 always  @(posedge pclk)
	ng2429<=ng34008;

 always  @(posedge pclk)
	ng1978<=ng33565;

 always  @(posedge pclk)
	ng6390<=ng24351;

 always  @(posedge pclk)
	ng3199<=ng30396;

 always  @(posedge pclk)
	ng1740<=ng33979;

 always  @(posedge pclk)
	ng2681<=ng30386;

 always  @(posedge pclk)
	ng2413<=ng30376;

 always  @(posedge pclk)
	ng5352<=ng24339;

 always  @(posedge pclk)
	ng6617<=ng30550;

 always  @(posedge pclk)
	ng2704<=ng34608;

 always  @(posedge pclk)
	ng2250<=ng29249;

 always  @(posedge pclk)
	ng2357<=ng33010;

 always  @(posedge pclk)
	ng5115<=ng29280;

 always  @(posedge pclk)
	ng5595<=ng30491;

 always  @(posedge pclk)
	ng2735<=ng29256;

 always  @(posedge pclk)
	ng4659<=ng34461;

 always  @(posedge pclk)
	ng1094<=ng29231;

 always  @(posedge pclk)
	ng534<=ng34723;

 always  @(posedge pclk)
	ng1521<=ng24252;

 always  @(posedge pclk)
	pg8787<=pg8786;

 always  @(posedge pclk)
	ng59<=ng28440;

 always  @(posedge pclk)
	ng772<=ng34252;

 always  @(posedge pclk)
	ng2563<=ng34015;

 always  @(posedge pclk)
	ng3598<=ng30427;

 always  @(posedge pclk)
	ng294<=ng33535;

 always  @(posedge pclk)
	ng921<=ng25621;

 always  @(posedge pclk)
	ng3522<=ng33028;

 always  @(posedge pclk)
	ng1379<=ng33543;

 always  @(posedge pclk)
	ng5587<=ng30489;

 always  @(posedge pclk)
	pg7946<=ng24256;

 always  @(posedge pclk)
	ng4264<=ng21894;

 always  @(posedge pclk)
	ng6291<=ng30534;

 always  @(posedge pclk)
	ng2955<=ng34807;

 always  @(posedge pclk)
	ng3115<=ng29258;

 always  @(posedge pclk)
	ng1724<=ng30352;

 always  @(posedge pclk)
	ng6177<=ng29301;

 always  @(posedge pclk)
	ng4593<=ng34452;

 always  @(posedge pclk)
	ng1024<=ng31869;

 always  @(posedge pclk)
	pg16656<=pg16627;

 always  @(posedge pclk)
	ng203<=ng25599;

 always  @(posedge pclk)
	ng5057<=ng33046;

 always  @(posedge pclk)
	ng6377<=pg17743;

 always  @(posedge pclk)
	ng4776<=ng34031;

 always  @(posedge pclk)
	ng5591<=ng30490;

 always  @(posedge pclk)
	ng5507<=ng34644;

 always  @(posedge pclk)
	ng452<=ng25604;

 always  @(posedge pclk)
	ng807<=ng34881;

 always  @(posedge pclk)
	ng1600<=ng33966;

 always  @(posedge pclk)
	ng4621<=ng34460;

 always  @(posedge pclk)
	ng1099<=ng24235;

 always  @(posedge pclk)
	ng2024<=ng33991;

 always  @(posedge pclk)
	ng4242<=ng24279;

 always  @(posedge pclk)
	ng2741<=ng30388;

 always  @(posedge pclk)
	ng2217<=ng33005;

 always  @(posedge pclk)
	ng6219<=ng33064;

 always  @(posedge pclk)
	ng1714<=ng33550;

 always  @(posedge pclk)
	ng1968<=ng30360;

 always  @(posedge pclk)
	ng4878<=ng34036;

 always  @(posedge pclk)
	pg11349<=ng24267;

 always  @(posedge pclk)
	pg8784<=pg8783;

 always  @(posedge pclk)
	ng5503<=ng29291;

 always  @(posedge pclk)
	pg11678<=pg12184;

 always  @(posedge pclk)
	ng595<=ng33538;

 always  @(posedge pclk)
	ng3542<=ng30416;

 always  @(posedge pclk)
	ng847<=ng24216;

 always  @(posedge pclk)
	pg12350<=ng24344;

 always  @(posedge pclk)
	ng1736<=ng33973;

 always  @(posedge pclk)
	ng2389<=ng30374;

 always  @(posedge pclk)
	ng2638<=ng29254;

 always  @(posedge pclk)
	ng2066<=ng33002;

 always  @(posedge pclk)
	ng4258<=ng21893;

 always  @(posedge pclk)
	ng5232<=ng30466;

 always  @(posedge pclk)
	ng6031<=pg17715;

 always  @(posedge pclk)
	ng4235<=pg8920;

 always  @(posedge pclk)
	ng3147<=ng29262;

 always  @(posedge pclk)
	ng4438<=ng26390;

 always  @(posedge pclk)
	ng5547<=ng30482;

 always  @(posedge pclk)
	ng4122<=ng28074;

 always  @(posedge pclk)
	ng1319<=ng24248;

 always  @(posedge pclk)
	ng1612<=ng33968;

 always  @(posedge pclk)
	ng5813<=ng25736;

 always  @(posedge pclk)
	ng4172<=ng34733;

 always  @(posedge pclk)
	ng490<=ng29223;

 always  @(posedge pclk)
	ng3457<=ng29263;

 always  @(posedge pclk)
	ng2844<=ng34609;

 always  @(posedge pclk)
	ng4709<=ng34032;

 always  @(posedge pclk)
	ng1291<=ng34602;

 always  @(posedge pclk)
	ng2449<=ng34012;

 always  @(posedge pclk)
	ng5212<=ng30477;

 always  @(posedge pclk)
	ng1830<=ng30354;

 always  @(posedge pclk)
	pg7243<=ng26945;

 always  @(posedge pclk)
	ng2907<=ng34617;

 always  @(posedge pclk)
	ng976<=ng24232;

 always  @(posedge pclk)
	ng2236<=ng29248;

 always  @(posedge pclk)
	pg12300<=ng24340;

 always  @(posedge pclk)
	ng6287<=ng30533;

 always  @(posedge pclk)
	ng5180<=ng33049;

 always  @(posedge pclk)
	ng918<=ng31868;

 always  @(posedge pclk)
	ng5945<=ng30513;

 always  @(posedge pclk)
	ng5517<=ng33052;

 always  @(posedge pclk)
	ng4245<=ng34632;

 always  @(posedge pclk)
	ng2246<=ng33579;

 always  @(posedge pclk)
	ng1932<=ng32998;

 always  @(posedge pclk)
	pg10527<=ng24255;

 always  @(posedge pclk)
	ng3941<=ng30446;

 always  @(posedge pclk)
	ng1744<=ng33974;

 always  @(posedge pclk)
	ng3512<=ng33026;

 always  @(posedge pclk)
	pg14451<=pg16656;

 always  @(posedge pclk)
	ng2657<=ng30384;

 always  @(posedge pclk)
	ng4933<=ng34267;

 always  @(posedge pclk)
	ng608<=ng34438;

 always  @(posedge pclk)
	ng1886<=ng33983;

 always  @(posedge pclk)
	ng1008<=ng25623;

 always  @(posedge pclk)
	ng645<=ng28046;

 always  @(posedge pclk)
	ng392<=ng24200;

 always  @(posedge pclk)
	ng146<=ng30333;

 always  @(posedge pclk)
	ng2671<=ng33605;

 always  @(posedge pclk)
	ng6565<=ng33069;

 always  @(posedge pclk)
	ng5909<=ng30505;

 always  @(posedge pclk)
	ng4372<=ng34882;

 always  @(posedge pclk)
	ng3155<=ng30393;

 always  @(posedge pclk)
	ng5607<=ng30494;

 always  @(posedge pclk)
	ng4521<=ng26971;

 always  @(posedge pclk)
	ng562<=ng25613;

 always  @(posedge pclk)
	ng4291<=pg9019;

 always  @(posedge pclk)
	ng3590<=ng30425;

 always  @(posedge pclk)
	ng218<=pg8291;

 always  @(posedge pclk)
	ng2028<=ng32999;

 always  @(posedge pclk)
	ng2685<=ng30387;

 always  @(posedge pclk)
	ng1802<=ng33554;

 always  @(posedge pclk)
	ng3490<=ng25668;

 always  @(posedge pclk)
	ng3167<=ng33022;

 always  @(posedge pclk)
	ng2295<=ng34001;

 always  @(posedge pclk)
	pg13865<=pg16874;

 always  @(posedge pclk)
	ng3813<=ng25684;

 always  @(posedge pclk)
	ng1205<=ng24244;

 always  @(posedge pclk)
	ng2208<=ng33004;

 always  @(posedge pclk)
	ng732<=ng25616;

 always  @(posedge pclk)
	ng4176<=ng34734;

 always  @(posedge pclk)
	ng6263<=ng30527;

 always  @(posedge pclk)
	ng4540<=ng31897;

 always  @(posedge pclk)
	ng121<=ng30389;

 always  @(posedge pclk)
	ng6732<=ng24354;

 always  @(posedge pclk)
	ng3554<=ng30432;

 always  @(posedge pclk)
	ng749<=ng31867;

 always  @(posedge pclk)
	ng5615<=ng30496;

 always  @(posedge pclk)
	ng6199<=ng34646;

 always  @(posedge pclk)
	ng2089<=ng33571;

 always  @(posedge pclk)
	pg9741<=ng25743;

 always  @(posedge pclk)
	ng3909<=ng30439;

 always  @(posedge pclk)
	ng2917<=ng34802;

 always  @(posedge pclk)
	ng2504<=ng29252;

 always  @(posedge pclk)
	pg11418<=ng24275;

 always  @(posedge pclk)
	ng2331<=ng33585;

 always  @(posedge pclk)
	ng6723<=pg17764;

 always  @(posedge pclk)
	ng6585<=ng30545;

 always  @(posedge pclk)
	ng6633<=ng30554;

 always  @(posedge pclk)
	ng4555<=ng4571;

 always  @(posedge pclk)
	ng4567<=ng33043;

 always  @(posedge pclk)
	ng1339<=ng24259;

 always  @(posedge pclk)
	ng767<=ng33965;

 always  @(posedge pclk)
	pg9617<=ng25728;

 always  @(posedge pclk)
	ng6259<=ng30541;

 always  @(posedge pclk)
	ng4405<=pg7243;

 always  @(posedge pclk)
	ng3945<=ng30447;

 always  @(posedge pclk)
	ng2748<=ng31872;

 always  @(posedge pclk)
	ng2283<=ng30372;

 always  @(posedge pclk)
	pg17423<=pg17404;

 always  @(posedge pclk)
	ng3698<=ng24274;

 always  @(posedge pclk)
	ng311<=ng26881;

 always  @(posedge pclk)
	ng1384<=ng25633;

 always  @(posedge pclk)
	ng5853<=ng34645;

 always  @(posedge pclk)
	ng5559<=ng30498;

 always  @(posedge pclk)
	ng5905<=ng30519;

 always  @(posedge pclk)
	ng872<=pg14167;

 always  @(posedge pclk)
	ng5471<=ng29287;

 always  @(posedge pclk)
	ng2169<=ng33995;

 assign pg28030 = ( wire34052 ) | ( wire34053 ) | ( wire34057 ) ;
 assign pg28041 = ( (~ ng19422) ) | ( (~ ng19402) ) ;
 assign pg33435 = ( (~ ng2729)  &  (~ ng23554) ) | ( (~ ng23554)  &  wire29308 ) | ( (~ ng23554)  &  wire29309 ) ;
 assign pg34425 = ( wire29245 ) | ( wire29246 ) | ( (~ wire3190)  &  (~ wire3191) ) ;
 assign pg30327 = ( (~ ng37) ) ;
 assign pg31793 = ( wire3189 ) | ( wire34096 ) | ( wire34099 ) | ( wire34101 ) ;
 assign pg21727 = ( (~ pg35)  &  ng3003 ) ;
 assign pg26876 = ( (~ ng17657) ) | ( (~ ng17700) ) ;
 assign pg30329 = ( (~ ng136) ) ;
 assign pg34239 = ( wire3176 ) | ( wire3177 ) | ( wire34166 ) | ( wire34167 ) ;
 assign pg26877 = ( (~ ng17694) ) | ( (~ ng17727) ) ;
 assign pg32454 = () ;
 assign pg34597 =((~ pg115) & pg115);
 assign pg23190 = ( (~ ng22)  &  (~ ng25) ) ;
 assign pg24151 = () ;
 assign pg33874 = ( ng66 ) | ( ng29186 ) ;
 assign pg28042 = ( (~ pg35) ) | ( ng1306 ) | ( ng962 ) ;
 assign pg12833 = ( (~ pg5) ) ;
 assign pg23652 = ( (~ ng2834) ) ;
 assign pg34201 = ( (~ ng25357) ) | ( wire28637 ) | ( wire28638 ) | ( wire34256 ) ;
 assign pg34236 = ( ni31843 ) | ( wire3140 ) | ( wire3141 ) | ( wire34275 ) ;
 assign pg34972 = ( (~ ng22) ) | ( ng34650 ) ;
 assign pg34956 = ( ng4369  &  (~ wire34278) ) | ( (~ pg72)  &  ng4322  &  ng4369 ) | ( pg72  &  (~ ng4322)  &  ng4369 ) ;
 assign pg23612 = ( (~ ng136) ) ;
 assign pg34232 = () ;
 assign pg30330 = ( (~ ng2834) ) ;
 assign pg30331 = ( (~ ng2831) ) ;
 assign pg34221 = ( ng29730 ) | ( (~ wire3190)  &  (~ wire3191) ) ;
 assign pg33948 = () ;
 assign pg34927 = ( (~ ng22) ) | ( ng33164 ) ;
 assign pg33949 = () ;
 assign pg34917 = ( (~ ng22) ) | ( ng33212 ) ;
 assign pg32185 = ( (~ wire3134)  &  (~ wire34279)  &  (~ wire34280)  &  (~ wire34281) ) ;
 assign pg33946 = () ;
 assign pg34839 = ( ng4369  &  (~ wire34278) ) | ( (~ pg72)  &  ng4322  &  ng4369 ) | ( pg72  &  (~ ng4322)  &  ng4369 ) ;
 assign pg33947 = () ;
 assign pg34919 = ( (~ ng22) ) | ( ni30751 ) | ( wire30180 ) | ( wire30181 ) ;
 assign pg34383 = ( (~ ng26314) ) | ( wire31726 ) | ( wire31727 ) | ( wire34290 ) ;
 assign pg34923 = ( (~ ng22) ) | ( ng33187 ) ;
 assign pg33079 = ( wire7186 ) | ( wire7187 ) | ( wire28915 ) | ( wire28916 ) ;
 assign pg33945 = () ;
 assign pg34913 = ( (~ ng22) ) | ( ng33219 ) ;
 assign pg33935 = ( (~ ng24374) ) | ( wire30515 ) | ( wire30516 ) | ( wire34292 ) ;
 assign pg34925 = ( (~ ng22) ) | ( ng33176 ) ;
 assign pg34915 = ( ng33149 ) | ( (~ ng22) ) ;
 assign pg33659 = ( (~ ng24688) ) | ( wire29507 ) | ( wire29508 ) | ( wire34294 ) ;
 assign pg33950 = () ;
 assign pg34921 = ( (~ ng22) ) | ( wire30135 ) | ( wire30136 ) | ( wire30150 ) ;
 assign pg26875 = ( (~ wire32542)  &  (~ wire32543) ) | ( (~ wire32544)  &  (~ wire32545) ) ;
 assign pg32429 = () ;
 assign pg23002 = ( (~ ng37) ) ;
 assign pg33636 = ( (~ ng24374) ) | ( wire32269 ) | ( wire32270 ) | ( wire34296 ) ;
 assign pg23759 = ( (~ ng2831) ) ;
 assign ng33063 = ( (~ pg35)  &  ng6209 ) | ( (~ ng26977)  &  wire28473 ) ;
 assign ng34455 = ( wire7734 ) | ( wire7735 ) | ( (~ pg35)  &  ng4322 ) ;
 assign ng24264 = ( pg125  &  pg35 ) ;
 assign ng26917 = ( wire28485 ) | ( ng10929  &  wire28483 ) | ( ng13846  &  wire28483 ) ;
 assign ng33013 = ( wire7720 ) | ( wire28507 ) | ( (~ pg35)  &  ng2491 ) ;
 assign ng26951 = ( (~ pg35)  &  ng4427 ) | ( pg35  &  ng4423 ) ;
 assign ng24281 = ( pg35  &  pg9251  &  (~ ng4308) ) | ( pg35  &  (~ pg9251)  &  (~ ng4308) ) ;
 assign ng30338 = ( pg35  &  ng24591 ) | ( pg35  &  (~ pg7916)  &  ng1171 ) | ( pg35  &  pg7916  &  (~ ng1171) ) ;
 assign ng30403 = ( wire7703 ) | ( (~ ng13977)  &  wire28521 ) | ( ng13977  &  wire28522 ) ;
 assign ng34610 = ( pg35  &  ng2852 ) | ( (~ pg35)  &  ng2844 ) ;
 assign ng33537 = ( wire7686 ) | ( (~ pg35)  &  ng301 ) ;
 assign ng25595 = ( pg35  &  (~ pg8719)  &  (~ ng358) ) ;
 assign ng34446 = ( wire28574 ) | ( pg35  &  ng29503  &  wire28571 ) ;
 assign ng34266 = ( wire7681 ) | ( wire28581 ) | ( ng29676  &  wire28577 ) ;
 assign ng24205 = ( wire7677 ) | ( (~ ng8806)  &  wire28583 ) | ( ng8806  &  wire28584 ) ;
 assign ng26907 = ( wire7671 ) | ( (~ ng10632)  &  wire28587 ) | ( ng10632  &  wire28588 ) ;
 assign ng33962 = ( wire7662 ) | ( wire7667 ) | ( wire7668 ) | ( wire28606 ) ;
 assign ng32983 = ( wire7647 ) | ( wire28612 ) ;
 assign ng34030 = ( wire28646 ) | ( ng28336  &  ng13464  &  wire28645 ) ;
 assign ng24277 = ( (~ pg35)  &  ng4040 ) | ( pg35  &  (~ ng4049)  &  (~ ng4040) ) | ( pg35  &  (~ ng4049)  &  ng8751 ) ;
 assign ng34605 = ( pg35  &  ng2145 ) | ( (~ pg35)  &  ng2138 ) ;
 assign ng29283 = ( wire7623 ) | ( wire28659 ) | ( (~ ng23590)  &  wire28655 ) ;
 assign ng33033 = ( (~ pg35)  &  ng3869 ) | ( (~ ng3873)  &  ng3869  &  (~ ng27635) ) | ( pg35  &  ng3873  &  (~ ng3869)  &  (~ ng27635) ) ;
 assign ng25678 = ( wire28670 ) | ( pg35  &  (~ pg8398)  &  ng3752 ) ;
 assign ng34598 = ( pg35  &  ng136 ) | ( (~ pg35)  &  ng550 ) ;
 assign ng33553 = ( wire7595 ) | ( wire7596 ) | ( (~ pg35)  &  ng1779 ) ;
 assign ng33023 = ( (~ pg35)  &  ng3167 ) | ( (~ ng3171)  &  ng3167  &  (~ ng27602) ) | ( pg35  &  ng3171  &  (~ ng3167)  &  (~ ng27602) ) ;
 assign ng25600 = ( (~ pg35)  &  ng174 ) | ( ng174  &  (~ ng11676) ) | ( pg35  &  ng168  &  ng11676 ) ;
 assign ng24207 = ( (~ pg35)  &  ng475 ) | ( ng475  &  (~ ng8806) ) | ( pg35  &  ng441  &  ng8806 ) ;
 assign ng34249 = ( wire28715 ) | ( pg35  &  (~ ng160)  &  ng31134 ) ;
 assign ng30343 = ( wire7567 ) | ( wire7568 ) | ( ng25917  &  wire28719 ) ;
 assign ng30551 = ( wire7565 ) | ( (~ ng14868)  &  wire28722 ) | ( ng14868  &  wire28723 ) ;
 assign ng24341 = ( (~ pg35)  &  ng5685 ) | ( pg35  &  ng5689  &  ng10160 ) | ( pg35  &  (~ ng5689)  &  (~ ng10160) ) ;
 assign ng30546 = ( wire28733 ) | ( (~ ng12632)  &  wire28732 ) | ( (~ ng12716)  &  wire28732 ) ;
 assign ng29294 = ( (~ pg35)  &  ng5821 ) | ( ng5821  &  (~ ng23666) ) | ( pg35  &  ng5827  &  ng23666 ) ;
 assign ng26893 = ( wire7346 ) | ( wire28741 ) ;
 assign ng29238 = ( wire7331 ) | ( wire7332 ) | ( wire28757 ) | ( wire28758 ) ;
 assign ng24347 = ( (~ pg35)  &  ng6040 ) | ( (~ ng6035)  &  ng6040 ) | ( ng6040  &  ng10185 ) ;
 assign ng29270 = ( wire7321 ) | ( wire7322 ) | ( wire7323 ) | ( wire7324 ) ;
 assign ng26883 = ( (~ pg35)  &  ng324 ) | ( pg35  &  ng305  &  ng324 ) | ( pg35  &  (~ ng324)  &  ng311 ) ;
 assign ng25609 = ( wire7310 ) | ( wire28779 ) | ( (~ ng11607)  &  wire28775 ) ;
 assign ng25662 = ( pg35  &  ng3530 ) ;
 assign ng33581 = ( wire7298 ) | ( wire7299 ) | ( wire7300 ) | ( wire7301 ) ;
 assign ng34803 = ( wire28792 ) | ( pg35  &  ng2932 ) | ( (~ pg35)  &  ng2917 ) ;
 assign ng30334 = ( wire28800 ) | ( (~ ng23978)  &  wire28796  &  wire28799 ) ;
 assign ng33964 = ( wire7286 ) | ( wire7287 ) | ( (~ pg35)  &  ng595 ) ;
 assign ng34600 = ( wire28820 ) | ( ng32212  &  (~ wire28816)  &  wire28819 ) ;
 assign ng33608 = ( wire28824 ) | ( (~ ng2756)  &  wire28822 ) | ( (~ ng25317)  &  wire28822 ) ;
 assign ng24263 = ( pg35  &  (~ ng2715) ) | ( (~ pg35)  &  ng2712 ) | ( pg35  &  (~ ng2841) ) ;
 assign ng33980 = ( wire7259 ) | ( wire7260 ) | ( ng30304  &  wire28830 ) ;
 assign ng30353 = ( wire7255 ) | ( wire28841 ) | ( (~ ng25385)  &  wire28837 ) ;
 assign ng29302 = ( (~ pg35)  &  ng6177 ) | ( pg35  &  ng6181  &  ng23699 ) | ( pg35  &  (~ ng6181)  &  (~ ng23699) ) ;
 assign ng33996 = ( wire7236 ) | ( wire7237 ) | ( ng30300  &  wire28849 ) ;
 assign ng32992 = ( wire7232 ) | ( wire28856 ) | ( (~ pg35)  &  ng1760 ) ;
 assign ng26889 = ( (~ pg35)  &  ng74 ) | ( (~ ng13385)  &  wire28858 ) ;
 assign ng34445 = ( wire28865 ) | ( pg35  &  ng29503  &  wire28860 ) ;
 assign ng30537 = ( wire7221 ) | ( (~ ng15036)  &  wire28866 ) | ( ng15036  &  wire28867 ) ;
 assign ng25670 = ( (~ pg35)  &  ng3498 ) | ( ng3498  &  ng12692 ) | ( pg35  &  ng3462  &  (~ ng12692) ) ;
 assign ng28044 = ( wire28874 ) | ( pg35  &  (~ ng482)  &  ng20000 ) | ( pg35  &  ng482  &  (~ ng20000) ) ;
 assign ng29242 = ( wire7202 ) | ( wire7204 ) | ( wire28891 ) | ( wire28892 ) ;
 assign ng34799 = ( pg35  &  (~ pg44) ) | ( pg35  &  ng2890 ) | ( (~ pg35)  &  ng2873 ) ;
 assign ng30346 = ( wire7190 ) | ( (~ ng24609)  &  wire28905 ) | ( (~ ng24609)  &  wire28907 ) ;
 assign ng33994 = ( wire7180 ) | ( wire7181 ) | ( ng30300  &  wire28920 ) ;
 assign ng34601 = ( pg35  &  ng947 ) ;
 assign ng34722 = ( pg35  &  ng546 ) | ( (~ pg35)  &  ng538 ) | ( pg35  &  (~ ng691) ) ;
 assign ng30454 = ( wire7175 ) | ( (~ ng14058)  &  wire28924 ) | ( ng14058  &  wire28925 ) ;
 assign ng24258 = ( (~ pg35)  &  ng1554 ) | ( pg35  &  ng496 ) ;
 assign ng30492 = ( wire7170 ) | ( (~ ng14885)  &  wire28927 ) | ( ng14885  &  wire28928 ) ;
 assign ng30437 = ( wire28933 ) | ( (~ ng11626)  &  wire28932 ) | ( (~ ng11763)  &  wire28932 ) ;
 assign ng25687 = ( wire28938 ) | ( pg35  &  ng2841  &  wire28937 ) ;
 assign ng29257 = ( wire7131 ) | ( wire7132 ) | ( wire7133 ) | ( wire7134 ) ;
 assign ng25682 = ( (~ pg35)  &  ng3835 ) | ( ng3835  &  ng12735 ) | ( pg35  &  ng3841  &  (~ ng12735) ) ;
 assign ng33987 = ( wire7116 ) | ( wire7117 ) | ( ng30311  &  wire29012 ) ;
 assign ng30424 = ( wire7114 ) | ( (~ ng14015)  &  wire29015 ) | ( ng14015  &  wire29016 ) ;
 assign ng34727 = ( pg35  &  ng939 ) | ( pg35  &  ng933 ) | ( (~ pg35)  &  ng952 ) ;
 assign ng29303 = ( pg35  &  ng4284  &  (~ ng14271) ) | ( pg35  &  (~ ng4180)  &  (~ ng14271) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng14271 ) ;
 assign ng32981 = ( wire7102 ) | ( wire29023 ) ;
 assign ng30526 = ( wire29027 ) | ( (~ ng12622)  &  wire29026 ) | ( (~ ng12667)  &  wire29026 ) ;
 assign ng33997 = ( wire7096 ) | ( wire7097 ) | ( ng30300  &  wire29029 ) ;
 assign ng29296 = ( (~ pg35)  &  ng5831 ) | ( pg35  &  ng5835  &  ng23666 ) | ( pg35  &  (~ ng5835)  &  (~ ng23666) ) ;
 assign ng33042 = ( wire29039 ) | ( wire29040 ) ;
 assign ng25697 = ( (~ pg35)  &  ng5084 ) | ( (~ ng5092)  &  ng5084 ) | ( pg35  &  ng5092  &  (~ ng5084) ) ;
 assign ng30444 = ( wire7083 ) | ( (~ ng14021)  &  wire29043 ) | ( ng14021  &  wire29044 ) ;
 assign ng29230 = ( wire7078 ) | ( wire29048 ) ;
 assign ng30438 = ( wire29051 ) | ( (~ ng11626)  &  wire29050 ) | ( (~ ng11537)  &  wire29050 ) ;
 assign ng24278 = ( (~ pg35)  &  ng4045 ) | ( ng4045  &  (~ ng4040) ) | ( ng4045  &  ng8751 ) ;
 assign ng25654 = ( (~ pg35)  &  ng3133 ) | ( ng3133  &  ng12641 ) | ( pg35  &  ng3139  &  (~ ng12641) ) ;
 assign ng30558 = ( wire7069 ) | ( (~ ng12915)  &  wire29054 ) | ( ng12915  &  wire29055 ) ;
 assign ng33601 = ( wire7058 ) | ( wire7059 ) | ( (~ pg35)  &  ng2606 ) ;
 assign ng29275 = ( wire29071 ) | ( ng4076  &  (~ ng13217)  &  wire29070 ) ;
 assign ng29237 = ( wire7049 ) | ( wire7050 ) | ( wire29087 ) | ( wire29088 ) ;
 assign ng29306 = ( (~ pg35)  &  ng6513 ) | ( ng6513  &  (~ ng23733) ) | ( pg35  &  ng6519  &  ng23733 ) ;
 assign ng30350 = ( (~ pg35)  &  ng1696 ) | ( pg35  &  ng1700  &  ng25275 ) | ( pg35  &  (~ ng1700)  &  (~ ng25275) ) ;
 assign ng33985 = ( wire29108 ) | ( ng29488  &  wire29104 ) | ( (~ ng29488)  &  wire29106 ) ;
 assign ng30377 = ( wire7028 ) | ( wire29119 ) | ( (~ ng25349)  &  wire29115 ) ;
 assign ng24208 = ( wire7024 ) | ( (~ ng8806)  &  wire29120 ) | ( ng8806  &  wire29121 ) ;
 assign ng26884 = ( wire29130 ) | ( wire29131 ) | ( ng13385  &  wire29129 ) ;
 assign ng25701 = ( (~ pg35)  &  ng5062 ) | ( pg35  &  ng5343 ) ;
 assign ng24348 = ( wire7008 ) | ( wire7009 ) | ( wire7010 ) | ( wire7011 ) ;
 assign ng33559 = ( wire7004 ) | ( wire7005 ) | ( wire7006 ) | ( wire7007 ) ;
 assign ng30392 = ( wire6992 ) | ( wire29184 ) | ( wire29185 ) | ( wire29186 ) ;
 assign ng25667 = ( (~ pg35)  &  ng3466 ) | ( pg35  &  (~ ng3470)  &  ng12692 ) | ( pg35  &  ng3470  &  (~ ng12692) ) ;
 assign ng33050 = ( wire6988 ) | ( (~ ng27999)  &  wire29195 ) | ( (~ ng27999)  &  wire29196 ) ;
 assign ng25610 = ( wire6985 ) | ( wire29202 ) | ( (~ ng11607)  &  wire29198 ) ;
 assign ng29309 = ( pg35  &  ng4284  &  (~ ng14306) ) | ( pg35  &  (~ ng4180)  &  (~ ng14306) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng14306 ) ;
 assign ng33062 = ( (~ pg35)  &  ng6203 ) | ( (~ ng6209)  &  ng6203  &  (~ ng26977) ) | ( pg35  &  ng6209  &  (~ ng6203)  &  (~ ng26977) ) ;
 assign ng24240 = ( (~ pg35)  &  ng996 ) | ( pg35  &  ng8417  &  ng16246 ) | ( pg35  &  (~ ng8417)  &  (~ ng16246) ) ;
 assign ng29264 = ( wire6965 ) | ( wire29223 ) | ( (~ ng23112)  &  wire29220 ) ;
 assign ng28063 = ( wire6959 ) | ( wire6960 ) | ( (~ pg35)  &  ng3263 ) ;
 assign ng34639 = ( pg35  &  ng4922 ) | ( (~ pg35)  &  ng4917 ) ;
 assign ng30549 = ( wire6956 ) | ( (~ ng14782)  &  wire29227 ) | ( ng14782  &  wire29228 ) ;
 assign ng26924 = ( wire29251 ) | ( (~ ng10961)  &  (~ ng13861)  &  wire29248 ) ;
 assign ng34020 = ( wire29260 ) | ( (~ ng29501)  &  wire29256 ) | ( ng29501  &  wire29258 ) ;
 assign ng33970 = ( wire6915 ) | ( wire6916 ) | ( ng30293  &  wire29265 ) ;
 assign ng33594 = ( wire6905 ) | ( wire6906 ) | ( (~ pg35)  &  ng2465 ) ;
 assign ng30488 = ( wire6904 ) | ( (~ ng14727)  &  wire29277 ) | ( ng14727  &  wire29278 ) ;
 assign ng34604 = ( pg35  &  ng2138 ) | ( (~ pg35)  &  ng2130 ) ;
 assign ng30469 = ( wire6899 ) | ( (~ ng14755)  &  wire29280 ) | ( ng14755  &  wire29281 ) ;
 assign ng26912 = ( wire29285 ) | ( (~ ng19063)  &  wire29283 ) ;
 assign ng24204 = ( (~ pg35)  &  ng433 ) | ( ng433  &  (~ ng8806) ) | ( pg35  &  ng429  &  ng8806 ) ;
 assign ng34467 = ( wire29293 ) | ( ng31009  &  (~ ng10862)  &  wire29292 ) ;
 assign ng34613 = ( pg35  &  ng37 ) | ( (~ pg35)  &  ng2894 ) ;
 assign ng24349 = ( (~ pg35)  &  ng6377 ) | ( pg35  &  ng6381  &  ng10207 ) | ( pg35  &  (~ ng6381)  &  (~ ng10207) ) ;
 assign ng21898 = ( (~ pg35)  &  ng4284 ) | ( pg35  &  pg9019  &  (~ ng4291) ) | ( pg35  &  (~ pg9019)  &  (~ ng4291) ) ;
 assign ng26927 = ( wire29303 ) | ( ng17625  &  (~ ng12377)  &  wire29300 ) ;
 assign ng30507 = ( wire6872 ) | ( (~ ng14697)  &  wire29304 ) | ( ng14697  &  wire29305 ) ;
 assign ng28092 = ( (~ pg35)  &  ng5057 ) | ( (~ ng25290)  &  wire29317 ) ;
 assign ng26914 = ( wire29323 ) | ( ng1052  &  (~ ng13121)  &  wire29322 ) ;
 assign ng26948 = ( ng4405 ) | ( (~ ng4405)  &  wire29324  &  wire29325  &  wire29328 ) ;
 assign ng30430 = ( wire6852 ) | ( (~ ng13923)  &  wire29329 ) | ( ng13923  &  wire29330 ) ;
 assign ng34037 = ( wire6847 ) | ( wire29336 ) ;
 assign ng26952 = ( wire6842 ) | ( wire6843 ) | ( wire6844 ) | ( wire29340 ) ;
 assign ng26939 = ( wire6838 ) | ( (~ pg35)  &  ng4104 ) ;
 assign ng30355 = ( (~ pg35)  &  ng1830 ) | ( pg35  &  ng1834  &  ng25300 ) | ( pg35  &  (~ ng1834)  &  (~ ng25300) ) ;
 assign ng33620 = ( wire6828 ) | ( wire6829 ) | ( (~ pg35)  &  ng5698 ) ;
 assign ng34024 = ( wire29361 ) | ( (~ wire6826)  &  (~ wire6827)  &  wire29355 ) ;
 assign ng29233 = ( wire6816 ) | ( wire6817 ) | ( wire29377 ) | ( wire29378 ) ;
 assign ng33040 = ( wire6808 ) | ( wire6809 ) | ( wire29383 ) ;
 assign ng34630 = ( pg35  &  ng4253 ) | ( (~ pg35)  &  ng4300 ) ;
 assign ng33617 = ( (~ pg35)  &  ng4552 ) | ( pg35  &  ng4552  &  (~ wire6804) ) | ( pg35  &  ng4581  &  (~ wire6804) ) ;
 assign ng24260 = ( (~ pg35)  &  ng1430 ) | ( (~ ng1548)  &  ng1430 ) | ( pg35  &  ng1548  &  (~ ng1430) ) ;
 assign ng21897 = ( (~ pg35)  &  ng4281 ) | ( pg35  &  (~ pg8839)  &  ng4281 ) | ( pg35  &  pg8839  &  (~ ng4281) ) ;
 assign ng25598 = ( (~ pg35)  &  ng376 ) | ( pg35  &  ng385  &  (~ ng358) ) | ( pg35  &  ng385  &  (~ ng376) ) | ( pg35  &  (~ ng385)  &  ng358  &  ng376 ) ;
 assign ng32977 = ( wire6789 ) | ( wire6790 ) | ( (~ pg35)  &  ng287 ) ;
 assign ng25656 = ( (~ pg35)  &  ng3147 ) | ( ng3147  &  ng12641 ) | ( pg35  &  ng3111  &  (~ ng12641) ) ;
 assign ng28051 = ( (~ pg35)  &  ng655 ) | ( ng655  &  (~ ng20248) ) | ( pg35  &  ng718  &  ng20248 ) ;
 assign ng30528 = ( wire6777 ) | ( (~ ng14741)  &  wire29402 ) | ( ng14741  &  wire29403 ) ;
 assign ng33588 = ( wire6763 ) | ( wire6764 ) | ( (~ pg35)  &  ng2393 ) ;
 assign ng34795 = ( wire29415 ) | ( pg35  &  (~ ni24685) ) | ( pg35  &  wire29414 ) ;
 assign ng26946 = ( wire29418 ) | ( (~ wire29325)  &  wire29417 ) | ( (~ wire29326)  &  wire29417 ) ;
 assign ng28099 = ( wire6715 ) | ( wire6716 ) | ( (~ pg35)  &  ng5965 ) ;
 assign ng30502 = ( wire29482 ) | ( (~ ng10312)  &  wire29481 ) | ( (~ ng12609)  &  wire29481 ) ;
 assign ng26899 = ( wire6709 ) | ( (~ ng17264)  &  wire29484 ) | ( ng17264  &  wire29486 ) ;
 assign ng33573 = ( wire6695 ) | ( wire6696 ) | ( wire6697 ) | ( wire6698 ) ;
 assign ng30481 = ( wire29518 ) | ( (~ ng10281)  &  wire29517 ) | ( (~ ng12558)  &  wire29517 ) ;
 assign ng26955 = ( wire29524 ) | ( wire29520  &  wire29521  &  wire29523 ) ;
 assign ng34250 = ( wire6686 ) | ( wire6687 ) | ( (~ pg35)  &  ng298 ) ;
 assign ng25703 = ( wire29532 ) | ( pg35  &  (~ pg9497)  &  ng5022 ) ;
 assign ng26922 = ( wire29537 ) | ( ng13273  &  wire29535 ) | ( ng10961  &  wire29535 ) ;
 assign ng30451 = ( wire6678 ) | ( (~ ng13963)  &  wire29538 ) | ( ng13963  &  wire29539 ) ;
 assign ng30337 = ( wire6674 ) | ( wire6675 ) | ( ng25911  &  wire29541 ) ;
 assign ng31902 = ( wire29555 ) | ( (~ wire29550)  &  (~ wire29551)  &  wire29553 ) ;
 assign ng25611 = ( wire6669 ) | ( (~ ng11607)  &  wire29556 ) | ( ng11607  &  wire29557 ) ;
 assign ng33989 = ( wire6665 ) | ( wire6666 ) | ( ng30311  &  wire29560 ) ;
 assign ng30486 = ( wire6663 ) | ( (~ ng14665)  &  wire29563 ) | ( ng14665  &  wire29564 ) ;
 assign ng31903 = ( wire6660 ) | ( ng26625  &  wire29567 ) | ( (~ ng26625)  &  wire29568 ) ;
 assign ng30362 = ( wire6653 ) | ( wire29579 ) | ( (~ ng25341)  &  wire29575 ) ;
 assign ng34801 = ( wire29581 ) | ( pg35  &  ng301 ) | ( (~ pg35)  &  ng2970 ) ;
 assign ng29269 = ( wire6619 ) | ( wire6620 ) | ( wire29644 ) ;
 assign ng33967 = ( wire6614 ) | ( wire6615 ) | ( ng30293  &  wire29647 ) ;
 assign ng33055 = ( wire6612 ) | ( (~ ng28010)  &  wire29652 ) | ( (~ ng28010)  &  wire29653 ) ;
 assign ng24201 = ( (~ pg35)  &  ng392 ) | ( ng392  &  (~ ng8806) ) | ( pg35  &  ng405  &  ng8806 ) ;
 assign ng25591 = ( (~ pg35)  &  ng209 ) | ( pg35  &  (~ ng218) ) ;
 assign ng25714 = ( pg35  &  ng5535 ) ;
 assign ng30411 = ( wire6604 ) | ( (~ ng13951)  &  wire29657 ) | ( ng13951  &  wire29658 ) ;
 assign ng28050 = ( (~ pg35)  &  ng650 ) | ( ng650  &  (~ ng20248) ) | ( pg35  &  ng655  &  ng20248 ) ;
 assign ng34458 = ( wire6598 ) | ( (~ ng31950)  &  wire29663 ) | ( (~ ng31950)  &  wire29665 ) ;
 assign ng28072 = ( wire29672 ) | ( (~ ng13806)  &  wire29671 ) | ( wire29669  &  wire29671 ) ;
 assign ng33961 = ( wire29676 ) | ( ng28444  &  (~ wire28561)  &  wire29675 ) ;
 assign ng24238 = ( wire6588 ) | ( (~ ng11148)  &  wire29683 ) ;
 assign ng33038 = ( wire29688 ) | ( wire29689 ) ;
 assign ng25761 = ( (~ pg35)  &  ng6509 ) | ( pg35  &  (~ ng6513)  &  ng10887 ) | ( pg35  &  ng6513  &  (~ ng10887) ) ;
 assign ng30468 = ( wire6576 ) | ( (~ ng14720)  &  wire29693 ) | ( ng14720  &  wire29694 ) ;
 assign ng28057 = ( wire6571 ) | ( wire6572 ) | ( (~ pg35)  &  ng1008 ) ;
 assign ng26910 = ( (~ pg35)  &  ng862 ) | ( ng862  &  ng890 ) | ( pg35  &  (~ ng862)  &  (~ ng890) ) ;
 assign ng24266 = ( (~ pg35)  &  ng2841 ) | ( pg35  &  ng2837  &  (~ ng2712) ) ;
 assign ng30509 = ( wire6565 ) | ( (~ ng14768)  &  wire29702 ) | ( ng14768  &  wire29703 ) ;
 assign ng25756 = ( pg35  &  ng6573 ) ;
 assign ng24215 = ( wire6561 ) | ( wire29711 ) | ( wire29712 ) ;
 assign ng34009 = ( wire6552 ) | ( wire6553 ) | ( ng30314  &  wire29715 ) ;
 assign ng34725 = ( wire6548 ) | ( wire6549 ) | ( (~ pg35)  &  ng781 ) ;
 assign ng34017 = ( wire6544 ) | ( wire6545 ) | ( ng29313  &  wire29724 ) ;
 assign ng30442 = ( wire6542 ) | ( (~ ng13960)  &  wire29727 ) | ( ng13960  &  wire29728 ) ;
 assign ng34264 = ( wire6539 ) | ( wire29735 ) | ( ng29719  &  wire29731 ) ;
 assign ng25630 = ( (~ pg35)  &  ng1249 ) | ( pg12923  &  (~ ng1266)  &  ng1249 ) | ( pg35  &  pg12923  &  ng1266  &  (~ ng1249) ) ;
 assign ng30562 = ( wire6532 ) | ( (~ ng14950)  &  wire29737 ) | ( ng14950  &  wire29738 ) ;
 assign ng34616 = ( pg35  &  ng2868 ) | ( (~ pg35)  &  ng2988 ) ;
 assign ng33070 = ( wire6527 ) | ( (~ ng26994)  &  wire29742 ) | ( (~ ng26994)  &  wire29743 ) ;
 assign ng29289 = ( wire6524 ) | ( wire29752 ) | ( (~ ng23630)  &  wire29747 ) ;
 assign ng25628 = ( wire29757 ) | ( (~ ng11148)  &  ng13570  &  wire29755 ) ;
 assign ng33555 = ( wire6515 ) | ( wire6516 ) | ( (~ pg35)  &  ng1816 ) ;
 assign ng29281 = ( wire6514 ) | ( wire29764 ) | ( (~ ng23590)  &  wire29761 ) ;
 assign ng24352 = ( wire6503 ) | ( wire6504 ) | ( wire29787 ) ;
 assign ng34791 = ( wire6500 ) | ( ng34162  &  wire29791 ) | ( (~ ng34162)  &  wire29792 ) ;
 assign ng29284 = ( (~ pg35)  &  ng5138 ) | ( pg35  &  ng5142  &  ng23590 ) | ( pg35  &  (~ ng5142)  &  (~ ng23590) ) ;
 assign ng30426 = ( wire6494 ) | ( (~ ng14075)  &  wire29797 ) | ( ng14075  &  wire29798 ) ;
 assign ng30515 = ( wire6491 ) | ( (~ ng14999)  &  wire29800 ) | ( ng14999  &  wire29801 ) ;
 assign ng33068 = ( (~ pg35)  &  ng6555 ) | ( (~ ng26994)  &  wire29804 ) ;
 assign ng34443 = ( wire29812 ) | ( pg35  &  ng29503  &  wire29809 ) ;
 assign ng26944 = ( wire6474 ) | ( wire6475 ) | ( wire6476 ) ;
 assign ng31898 = ( wire29843 ) | ( (~ wire29550)  &  (~ wire29551)  &  wire29841 ) ;
 assign ng25705 = ( (~ pg35)  &  ng5124 ) | ( pg35  &  (~ ng5128)  &  ng10823 ) | ( pg35  &  ng5128  &  (~ ng10823) ) ;
 assign ng34026 = ( (~ pg35)  &  ng4646 ) | ( ng4646  &  ng31003 ) ;
 assign ng30457 = ( wire29852 ) | ( wire29853 ) | ( ng26256  &  wire29851 ) ;
 assign ng30390 = ( wire6451 ) | ( wire29184 ) | ( wire29185 ) | ( wire29186 ) ;
 assign ng30404 = ( wire6450 ) | ( (~ ng14008)  &  wire29855 ) | ( ng14008  &  wire29856 ) ;
 assign ng29236 = ( wire6442 ) | ( wire6443 ) | ( wire29873 ) | ( wire29874 ) ;
 assign ng21895 = ( (~ pg35)  &  ng4264 ) | ( pg35  &  ng4269  &  (~ ng4264) ) | ( pg35  &  ng4269  &  (~ ng4258) ) | ( pg35  &  (~ ng4269)  &  ng4264  &  ng4258 ) ;
 assign ng24269 = ( (~ pg35)  &  ng3338 ) | ( pg35  &  (~ ng3338)  &  (~ ng3347) ) | ( pg35  &  (~ ng3347)  &  ng8691 ) ;
 assign ng34448 = ( wire29890 ) | ( pg35  &  ng29503  &  wire29887 ) ;
 assign ng25650 = ( wire29894 ) | ( pg35  &  (~ pg8277)  &  ng3050 ) ;
 assign ng33036 = ( wire29899 ) | ( wire29900 ) ;
 assign ng30341 = ( wire6424 ) | ( (~ ng24591)  &  wire29903 ) | ( (~ ng24591)  &  wire29905 ) ;
 assign ng30540 = ( wire6421 ) | ( (~ ng14864)  &  wire29907 ) | ( ng14864  &  wire29908 ) ;
 assign ng34730 = ( pg35  &  ng1283 ) | ( pg35  &  ng1277 ) | ( (~ pg35)  &  ng1296 ) ;
 assign ng25763 = ( wire6415 ) | ( wire29917 ) | ( ng10887  &  wire29912 ) ;
 assign ng24282 = ( (~ pg35)  &  ng4308 ) | ( pg35  &  (~ pg9251)  &  ng4308 ) | ( pg35  &  pg9251  &  (~ ng4308) ) ;
 assign ng34451 = ( wire29923 ) | ( (~ ng30583)  &  (~ wire6408)  &  wire29922 ) ;
 assign ng25729 = ( (~ pg35)  &  ng5752 ) | ( pg35  &  ng6035 ) ;
 assign ng34980 = ( wire30237 ) | ( ng34650  &  wire30236 ) ;
 assign ng24254 = ( wire6398 ) | ( (~ ng11171)  &  wire30245 ) ;
 assign ng29235 = ( wire6395 ) | ( wire6396 ) | ( (~ pg35)  &  ng1252 ) ;
 assign ng34003 = ( wire6389 ) | ( wire6390 ) | ( ng30307  &  wire30250 ) ;
 assign ng25715 = ( pg35  &  ng5689 ) | ( (~ pg35)  &  ng5406 ) ;
 assign ng33149 = ( wire30061 ) | ( wire30062 ) | ( wire30081 ) | ( wire30082 ) ;
 assign ng33197 = ( wire30131 ) | ( wire30132 ) | ( wire30136 ) | ( wire30150 ) ;
 assign ng28089 = ( wire30267 ) | ( wire30268 ) | ( wire30269 ) ;
 assign ng30463 = ( wire30274 ) | ( (~ ng12443)  &  wire30273 ) | ( (~ ng12492)  &  wire30273 ) ;
 assign ng33562 = ( wire6363 ) | ( wire6364 ) | ( (~ pg35)  &  ng1906 ) ;
 assign ng33546 = ( wire6361 ) | ( wire30286 ) ;
 assign ng24272 = ( (~ pg35)  &  ng3680 ) | ( pg35  &  ng3689  &  ng8728 ) | ( pg35  &  (~ ng3689)  &  (~ ng8728) ) ;
 assign ng34628 = ( pg35  &  ng4146 ) | ( (~ pg35)  &  ng4176 ) ;
 assign ng34027 = ( (~ pg35)  &  ng4674 ) | ( ng4674  &  ng31003 ) ;
 assign ng28055 = ( wire6348 ) | ( (~ ng20905)  &  wire30293 ) | ( ng20905  &  wire30295 ) ;
 assign ng31865 = ( (~ pg35)  &  ng283 ) | ( (~ ng287)  &  ng283  &  ng23204 ) | ( pg35  &  ng287  &  (~ ng283)  &  ng23204 ) ;
 assign ng32985 = ( wire6341 ) | ( (~ pg35)  &  ng1274 ) ;
 assign ng26931 = ( wire30304 ) | ( ng17625  &  (~ ng12377)  &  wire30301 ) ;
 assign ng29244 = ( wire6333 ) | ( wire6335 ) | ( wire30320 ) | ( wire30321 ) ;
 assign ng34439 = ( wire6329 ) | ( (~ ng32212)  &  wire30324 ) | ( ng32212  &  wire30325 ) ;
 assign ng34849 = ( wire6324 ) | ( wire6325 ) | ( (~ pg35)  &  ng622 ) ;
 assign ng34459 = ( wire6323 ) | ( wire30341 ) | ( ng31971  &  wire30337 ) ;
 assign ng30363 = ( wire6317 ) | ( wire30348 ) | ( (~ ng25470)  &  wire30344 ) ;
 assign ng24247 = ( pg35  &  pg12923  &  (~ ng1249) ) ;
 assign ng30365 = ( (~ pg35)  &  ng2098 ) | ( pg35  &  ng2102  &  ng25389 ) | ( pg35  &  (~ ng2102)  &  (~ ng25389) ) ;
 assign ng29300 = ( (~ pg35)  &  ng6167 ) | ( ng6167  &  (~ ng23699) ) | ( pg35  &  ng6173  &  ng23699 ) ;
 assign ng33591 = ( wire6304 ) | ( wire6305 ) | ( wire6306 ) | ( wire6307 ) ;
 assign ng33626 = ( wire6301 ) | ( wire6302 ) | ( (~ pg35)  &  ng6736 ) ;
 assign ng29305 = ( wire6300 ) | ( wire30375 ) | ( (~ ng23733)  &  wire30372 ) ;
 assign ng33570 = ( wire6294 ) | ( wire6295 ) | ( (~ pg35)  &  ng2040 ) ;
 assign ng30484 = ( wire30384 ) | ( (~ ng12505)  &  wire30383 ) | ( (~ ng12558)  &  wire30383 ) ;
 assign ng34256 = ( wire6283 ) | ( wire30388 ) | ( pg35  &  (~ ng33394) ) ;
 assign ng34011 = ( wire6281 ) | ( wire6282 ) | ( ng30314  &  wire30391 ) ;
 assign ng33590 = ( wire6277 ) | ( wire6278 ) | ( (~ pg35)  &  ng2403 ) ;
 assign ng29240 = ( wire6273 ) | ( wire6274 ) | ( wire30411 ) | ( wire30412 ) ;
 assign ng25699 = ( (~ pg35)  &  ng5097 ) | ( pg35  &  ng86  &  (~ ng5097) ) | ( pg35  &  ng86  &  ng9724 ) | ( pg35  &  (~ ng86)  &  ng5097  &  (~ ng9724) ) ;
 assign ng26934 = ( wire30420 ) | ( ng17625  &  (~ ng12377)  &  wire30417 ) ;
 assign ng25636 = ( wire6260 ) | ( (~ ng13291)  &  wire30421 ) | ( ng13291  &  wire30422 ) ;
 assign ng30344 = ( pg35  &  ng24609 ) | ( pg35  &  (~ pg7946)  &  ng1514 ) | ( pg35  &  pg7946  &  (~ ng1514) ) ;
 assign ng34633 = ( pg35  &  ng4727 ) ;
 assign ng30399 = ( wire6254 ) | ( (~ ng13873)  &  wire30427 ) | ( ng13873  &  wire30428 ) ;
 assign ng30561 = ( wire6251 ) | ( (~ ng14908)  &  wire30430 ) | ( ng14908  &  wire30431 ) ;
 assign ng30520 = ( wire6248 ) | ( (~ ng14858)  &  wire30433 ) | ( ng14858  &  wire30434 ) ;
 assign ng30409 = ( wire6245 ) | ( (~ ng13892)  &  wire30436 ) | ( ng13892  &  wire30437 ) ;
 assign ng34805 = ( pg35  &  ng2932 ) | ( pg35  &  ng2999 ) ;
 assign ng33599 = ( wire6237 ) | ( wire6238 ) | ( wire6239 ) | ( wire6240 ) ;
 assign ng30410 = ( wire6236 ) | ( (~ ng11432)  &  wire30447 ) | ( ng11432  &  wire30448 ) ;
 assign ng31895 = ( (~ pg35)  &  ng4382 ) | ( pg35  &  ng29503 ) ;
 assign ng34619 = ( pg35  &  ng2922 ) | ( (~ pg35)  &  ng2912 ) ;
 assign ng25664 = ( wire30453 ) | ( pg35  &  (~ pg8342)  &  ng3401 ) ;
 assign ng25653 = ( (~ pg35)  &  ng3115 ) | ( pg35  &  (~ ng3119)  &  ng12641 ) | ( pg35  &  ng3119  &  (~ ng12641) ) ;
 assign ng30412 = ( wire6223 ) | ( (~ ng13980)  &  wire30457 ) | ( ng13980  &  wire30458 ) ;
 assign ng25681 = ( (~ pg35)  &  ng3817 ) | ( pg35  &  (~ ng3821)  &  ng12735 ) | ( pg35  &  ng3821  &  (~ ng12735) ) ;
 assign ng30395 = ( wire30466 ) | ( (~ ng11514)  &  wire30465 ) | ( (~ ng11729)  &  wire30465 ) ;
 assign ng30380 = ( (~ pg35)  &  ng2523 ) | ( pg35  &  ng2527  &  ng25400 ) | ( pg35  &  (~ ng2527)  &  (~ ng25400) ) ;
 assign ng30405 = ( wire6211 ) | ( (~ ng14041)  &  wire30471 ) | ( ng14041  &  wire30472 ) ;
 assign ng30476 = ( wire6208 ) | ( (~ ng12402)  &  wire30474 ) | ( ng12402  &  wire30475 ) ;
 assign ng33560 = ( wire6205 ) | ( ng28927  &  wire30480 ) ;
 assign ng24236 = ( wire30484 ) | ( pg35  &  pg7916  &  ng996 ) ;
 assign ng33029 = ( wire6197 ) | ( (~ ng27617)  &  wire30487 ) | ( (~ ng27617)  &  wire30488 ) ;
 assign ng24280 = ( (~ pg35)  &  ng4269 ) | ( pg35  &  (~ ng4269)  &  ng4273 ) | ( pg35  &  ng4273  &  ng8967 ) | ( pg35  &  ng4269  &  (~ ng4273)  &  (~ ng8967) ) ;
 assign ng30370 = ( (~ pg35)  &  ng2255 ) | ( pg35  &  ng2259  &  ng25309 ) | ( pg35  &  (~ ng2259)  &  (~ ng25309) ) ;
 assign ng25749 = ( wire6167 ) | ( wire30566 ) | ( ng10874  &  wire30562 ) ;
 assign ng30538 = ( wire6163 ) | ( (~ ng14776)  &  wire30567 ) | ( ng14776  &  wire30568 ) ;
 assign ng34025 = ( pg35  &  (~ ng4639)  &  (~ ng31950) ) ;
 assign ng31899 = ( wire30574 ) | ( (~ wire29550)  &  (~ wire29551)  &  wire30572 ) ;
 assign ng30531 = ( wire6157 ) | ( (~ ng14861)  &  wire30575 ) | ( ng14861  &  wire30576 ) ;
 assign ng33619 = ( wire6151 ) | ( (~ ng28982)  &  wire30581 ) | ( (~ ng28982)  &  wire30583 ) ;
 assign ng26903 = ( wire6148 ) | ( (~ ng10632)  &  wire30585 ) | ( ng10632  &  wire30586 ) ;
 assign ng29268 = ( pg35  &  ng4284  &  (~ ng13517) ) | ( pg35  &  (~ ng4180)  &  (~ ng13517) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng13517 ) ;
 assign ng33067 = ( (~ pg35)  &  ng6549 ) | ( (~ ng6555)  &  ng6549  &  (~ ng26994) ) | ( pg35  &  ng6555  &  (~ ng6549)  &  (~ ng26994) ) ;
 assign ng26923 = ( wire30596 ) | ( ng13315  &  wire30593 ) | ( ng10961  &  wire30593 ) ;
 assign ng28085 = ( wire30611 ) | ( wire30612 ) | ( wire30613 ) ;
 assign ng33583 = ( wire6125 ) | ( wire6126 ) | ( wire6127 ) | ( wire6128 ) ;
 assign ng26909 = ( (~ pg35)  &  ng890 ) | ( pg35  &  (~ ng896)  &  ng862 ) | ( pg35  &  ng896  &  (~ ng890) ) ;
 assign ng24355 = ( (~ pg35)  &  ng6732 ) | ( (~ ng6727)  &  ng6732 ) | ( ng6732  &  ng10224 ) ;
 assign ng29304 = ( wire6093 ) | ( wire6094 ) | ( wire6095 ) | ( wire6096 ) ;
 assign ng26926 = ( wire30695 ) | ( pg35  &  ng2841  &  wire30694 ) ;
 assign ng34796 = ( wire30708 ) | ( pg35  &  ng17694 ) | ( pg35  &  ng17727 ) ;
 assign ng33598 = ( wire6068 ) | ( wire6069 ) | ( (~ pg35)  &  ng2537 ) ;
 assign ng30559 = ( wire6067 ) | ( (~ ng14825)  &  wire30712 ) | ( ng14825  &  wire30713 ) ;
 assign ng28087 = ( wire30729 ) | ( wire30730 ) | ( wire30731 ) ;
 assign ng33012 = ( wire6055 ) | ( wire30737 ) | ( (~ pg35)  &  ng2453 ) ;
 assign ng28060 = ( wire30740 ) | ( pg35  &  (~ ng2729)  &  ng14291 ) | ( pg35  &  ng2729  &  (~ ng14291) ) ;
 assign ng33540 = ( wire6048 ) | ( wire6049 ) | ( (~ pg35)  &  ng925 ) ;
 assign ng33627 = ( wire6047 ) | ( (~ ng29110)  &  wire30746 ) | ( (~ ng29110)  &  wire30748 ) ;
 assign ng34615 = ( (~ pg35)  &  ng2868 ) | ( pg35  &  ng2873 ) ;
 assign ng34040 = ( wire30754 ) | ( ng16187  &  ng28349  &  wire30752 ) ;
 assign ng29267 = ( (~ pg35)  &  ng3480 ) | ( pg35  &  ng3484  &  ng23112 ) | ( pg35  &  (~ ng3484)  &  (~ ng23112) ) ;
 assign ng34251 = ( wire6036 ) | ( ng31509  &  wire30759 ) | ( (~ ng31509)  &  wire30760 ) ;
 assign ng29243 = ( wire6033 ) | ( wire30768 ) | ( ng22369  &  wire30763 ) ;
 assign ng26950 = ( wire6028 ) | ( wire6029 ) | ( (~ pg35)  &  ng4417 ) ;
 assign ng25634 = ( pg35  &  ng1395  &  (~ ng1322)  &  ng13134 ) | ( pg35  &  (~ ng1395)  &  (~ ng1322)  &  (~ ng13134) ) ;
 assign ng29227 = ( wire6015 ) | ( (~ ng23324)  &  wire30805 ) | ( (~ ng23324)  &  wire30807 ) ;
 assign ng26896 = ( wire6009 ) | ( wire6010 ) | ( wire6011 ) | ( wire6012 ) ;
 assign ng25764 = ( (~ pg35)  &  ng6541 ) | ( ng6541  &  ng10887 ) | ( pg35  &  ng6505  &  (~ ng10887) ) ;
 assign ng29286 = ( wire5979 ) | ( wire5980 ) | ( wire5981 ) | ( wire5982 ) ;
 assign ng28091 = ( (~ pg35)  &  ng5069 ) | ( (~ ng25371)  &  wire30880 ) ;
 assign ng33545 = ( wire5968 ) | ( wire5969 ) | ( (~ pg35)  &  ng1644 ) ;
 assign ng29297 = ( pg35  &  ng4284  &  (~ ng14247) ) | ( pg35  &  (~ ng4180)  &  (~ ng14247) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng14247 ) ;
 assign ng33577 = ( wire5963 ) | ( wire5964 ) | ( (~ pg35)  &  ng2204 ) ;
 assign ng30357 = ( wire5959 ) | ( wire30898 ) | ( (~ ng25300)  &  wire30893 ) ;
 assign ng30544 = ( wire30901 ) | ( (~ ng7142)  &  wire30900 ) | ( (~ ng12716)  &  wire30900 ) ;
 assign ng30358 = ( wire5952 ) | ( wire30906 ) | ( (~ ng25429)  &  wire30902 ) ;
 assign ng30367 = ( wire5948 ) | ( wire30912 ) | ( (~ ng25389)  &  wire30908 ) ;
 assign ng31866 = ( wire5942 ) | ( wire5943 ) | ( (~ pg35)  &  ng577 ) ;
 assign ng25683 = ( wire5941 ) | ( wire30923 ) | ( ng12735  &  wire30918 ) ;
 assign ng29246 = ( wire5928 ) | ( wire5929 ) | ( wire30938 ) | ( wire30939 ) ;
 assign ng25734 = ( (~ pg35)  &  ng5835 ) | ( ng5835  &  ng10869 ) | ( pg35  &  ng5841  &  (~ ng10869) ) ;
 assign ng21892 = ( (~ pg35)  &  ng4273 ) | ( pg35  &  (~ ng4239) ) ;
 assign ng25706 = ( (~ pg35)  &  ng5142 ) | ( ng5142  &  ng10823 ) | ( pg35  &  ng5148  &  (~ ng10823) ) ;
 assign ng28093 = ( wire5888 ) | ( wire5889 ) | ( (~ pg35)  &  ng5272 ) ;
 assign ng33016 = ( wire5883 ) | ( wire31010 ) | ( (~ pg35)  &  ng2587 ) ;
 assign ng24353 = ( (~ pg35)  &  ng6723 ) | ( pg35  &  ng6727  &  ng10224 ) | ( pg35  &  (~ ng6727)  &  (~ ng10224) ) ;
 assign ng25655 = ( wire5878 ) | ( wire31020 ) | ( ng12641  &  wire31015 ) ;
 assign ng34642 = ( pg35  &  ng4927 ) | ( (~ pg35)  &  ng4912 ) ;
 assign ng25704 = ( (~ pg35)  &  ng5073 ) | ( ng5069  &  ng5073 ) ;
 assign ng33008 = ( wire5868 ) | ( wire31025 ) | ( (~ pg35)  &  ng2319 ) ;
 assign ng30421 = ( wire5866 ) | ( (~ ng13920)  &  wire31026 ) | ( ng13920  &  wire31027 ) ;
 assign ng33007 = ( wire5856 ) | ( wire31034 ) | ( wire31036 ) ;
 assign ng25730 = ( wire31040 ) | ( pg35  &  (~ pg9680)  &  ng5752 ) ;
 assign ng25624 = ( wire31043 ) | ( pg35  &  (~ ng13211)  &  wire5848 ) ;
 assign ng34255 = ( (~ ng33394) ) | ( wire31045 ) ;
 assign ng30371 = ( (~ pg35)  &  ng2273 ) | ( ng2273  &  (~ ng25309) ) | ( pg35  &  ng2279  &  ng25309 ) ;
 assign ng26900 = ( pg35  &  ng106 ) ;
 assign ng33607 = ( wire5835 ) | ( wire5836 ) | ( wire5837 ) | ( wire5838 ) ;
 assign ng26904 = ( wire5834 ) | ( (~ ng10632)  &  wire31056 ) | ( ng10632  &  wire31057 ) ;
 assign ng34626 = ( pg35  &  ng3502 ) ;
 assign ng29293 = ( wire5831 ) | ( wire31063 ) | ( (~ ng23666)  &  wire31060 ) ;
 assign ng34268 = ( wire5827 ) | ( wire31069 ) | ( ng29722  &  wire31065 ) ;
 assign ng29271 = ( wire5821 ) | ( wire5822 ) | ( (~ pg35)  &  ng3821 ) ;
 assign ng28083 = ( wire31086 ) | ( wire31087 ) | ( wire31088 ) ;
 assign ng26886 = ( wire5814 ) | ( (~ ng13385)  &  wire31090 ) | ( ng13385  &  wire31091 ) ;
 assign ng33576 = ( wire5811 ) | ( ng28903  &  wire31095 ) ;
 assign ng29266 = ( wire5809 ) | ( wire31102 ) | ( (~ ng23112)  &  wire31098 ) ;
 assign ng34260 = ( ng31003  &  (~ ng10831)  &  wire31105 ) ;
 assign ng33618 = ( wire5803 ) | ( wire5804 ) | ( (~ pg35)  &  ng5352 ) ;
 assign ng34640 = ( (~ pg35)  &  ng4922 ) | ( pg35  &  ng4907 ) ;
 assign ng30445 = ( wire5800 ) | ( (~ ng14055)  &  wire31111 ) | ( ng14055  &  wire31112 ) ;
 assign ng30514 = ( wire5797 ) | ( (~ ng14968)  &  wire31114 ) | ( ng14968  &  wire31115 ) ;
 assign ng30356 = ( (~ pg35)  &  ng1848 ) | ( ng1848  &  (~ ng25300) ) | ( pg35  &  ng1854  &  ng25300 ) ;
 assign ng25685 = ( pg35  &  (~ ng2841) ) | ( pg35  &  (~ ng4064) ) | ( (~ pg35)  &  ng4072 ) ;
 assign ng30525 = ( wire31122 ) | ( (~ ng12581)  &  wire31121 ) | ( (~ ng12667)  &  wire31121 ) ;
 assign ng30342 = ( wire5783 ) | ( wire5785 ) | ( ng25895  &  wire31124 ) ;
 assign ng30560 = ( wire5782 ) | ( (~ ng12629)  &  wire31126 ) | ( ng12629  &  wire31127 ) ;
 assign ng33567 = ( wire5773 ) | ( wire5774 ) | ( wire5775 ) | ( wire5776 ) ;
 assign ng29290 = ( (~ pg35)  &  ng5485 ) | ( pg35  &  ng5489  &  ng23630 ) | ( pg35  &  (~ ng5489)  &  (~ ng23630) ) ;
 assign ng25602 = ( wire5769 ) | ( (~ ng11676)  &  wire31140 ) | ( ng11676  &  wire31141 ) ;
 assign ng33544 = ( wire5766 ) | ( ng28853  &  wire31146 ) ;
 assign ng34606 = ( pg35  &  ng2689 ) ;
 assign ng34013 = ( wire31153 ) | ( (~ ng29496)  &  wire31149 ) | ( ng29496  &  wire31151 ) ;
 assign ng30441 = ( wire5755 ) | ( (~ ng13929)  &  wire31155 ) | ( ng13929  &  wire31156 ) ;
 assign ng33977 = ( wire5747 ) | ( wire5748 ) | ( ng30298  &  wire31158 ) ;
 assign ng34621 = ( pg35  &  ng2950 ) | ( (~ pg35)  &  ng2936 ) ;
 assign ng26908 = ( wire5740 ) | ( ng10632  &  wire31161 ) | ( (~ ng10632)  &  wire31162 ) ;
 assign ng34257 = ( wire5737 ) | ( (~ ng30583)  &  wire31165 ) | ( (~ ng30583)  &  wire31167 ) ;
 assign ng29299 = ( wire5734 ) | ( wire31173 ) | ( (~ ng23699)  &  wire31170 ) ;
 assign ng30470 = ( wire5730 ) | ( (~ ng14797)  &  wire31174 ) | ( ng14797  &  wire31175 ) ;
 assign ng26954 = ( wire31178 ) | ( ng4438  &  (~ wire6690)  &  (~ wire29524) ) ;
 assign ng21901 = ( wire31189 ) | ( wire31182  &  wire31183  &  wire31184 ) ;
 assign ng33574 = ( wire5718 ) | ( wire5719 ) | ( (~ pg35)  &  ng2112 ) ;
 assign ng34607 = ( (~ pg35)  &  ng2689 ) | ( pg35  &  ng2697 ) ;
 assign ng33011 = ( wire5712 ) | ( wire31198 ) | ( (~ pg35)  &  ng2461 ) ;
 assign ng26965 = ( (~ pg35)  &  ng4534 ) | ( (~ pg10306)  &  ng4534 ) | ( pg35  &  pg10306  &  (~ ng4534) ) ;
 assign ng30429 = ( wire5705 ) | ( (~ ng14151)  &  wire31201 ) | ( ng14151  &  wire31202 ) ;
 assign ng25619 = ( wire31206 ) | ( (~ ng847)  &  wire31205 ) | ( ng8806  &  wire31205 ) ;
 assign ng30414 = ( pg35  &  (~ ng3506)  &  (~ ng3518)  &  (~ ng27617) ) ;
 assign ng33541 = ( wire5697 ) | ( wire5698 ) | ( (~ pg35)  &  ng1030 ) ;
 assign ng33615 = ( wire5693 ) | ( wire5694 ) | ( wire31215 ) ;
 assign ng33548 = ( wire5690 ) | ( wire5691 ) | ( (~ pg35)  &  ng1700 ) ;
 assign ng33053 = ( (~ pg35)  &  ng5517 ) | ( (~ ng28010)  &  wire31220 ) ;
 assign ng25750 = ( (~ pg35)  &  ng6195 ) | ( ng6195  &  ng10874 ) | ( pg35  &  ng6159  &  (~ ng10874) ) ;
 assign ng34622 = ( (~ pg35)  &  ng2950 ) | ( pg35  &  ng2960 ) ;
 assign ng25720 = ( (~ pg35)  &  ng5489 ) | ( ng5489  &  ng10838 ) | ( pg35  &  ng5495  &  (~ ng10838) ) ;
 assign ng34804 = ( wire31226 ) | ( pg35  &  ng2975 ) | ( (~ pg35)  &  ng2965 ) ;
 assign ng30543 = ( pg35  &  (~ ng6561)  &  (~ ng6549)  &  (~ ng26994) ) ;
 assign ng34005 = ( wire5671 ) | ( wire5672 ) | ( ng30307  &  wire31229 ) ;
 assign ng30383 = ( wire5669 ) | ( wire31237 ) | ( (~ ng25498)  &  wire31233 ) ;
 assign ng34647 = ( pg35  &  ng6545 ) ;
 assign ng29255 = ( wire5663 ) | ( wire5664 ) | ( wire31242 ) ;
 assign ng30523 = ( wire31246 ) | ( (~ ng10341)  &  wire31245 ) | ( (~ ng12667)  &  wire31245 ) ;
 assign ng24211 = ( wire5653 ) | ( wire5654 ) | ( (~ pg35)  &  ng546 ) ;
 assign ng33556 = ( wire5650 ) | ( wire5651 ) | ( (~ pg35)  &  ng1834 ) ;
 assign ng24214 = ( wire5645 ) | ( wire5648 ) | ( wire31259 ) ;
 assign ng25700 = ( pg35  &  ng5188 ) ;
 assign ng25691 = ( wire5638 ) | ( wire5643 ) | ( wire5644 ) | ( wire31271 ) ;
 assign ng29261 = ( (~ pg35)  &  ng3129 ) | ( pg35  &  ng3133  &  ng23067 ) | ( pg35  &  (~ ng3133)  &  (~ ng23067) ) ;
 assign ng27511 = ( pg54  &  (~ pg53)  &  wire29926 ) ;
 assign ng33561 = ( wire5632 ) | ( wire5633 ) | ( (~ pg35)  &  ng1913 ) ;
 assign ng34641 = ( (~ pg35)  &  ng4907 ) | ( pg35  &  ng4912 ) ;
 assign ng29245 = ( wire5627 ) | ( wire5628 ) | ( wire31283 ) ;
 assign ng30435 = ( pg35  &  (~ ng3857)  &  (~ ng3869)  &  (~ ng27635) ) ;
 assign ng34006 = ( wire31292 ) | ( (~ ng29489)  &  wire31288 ) | ( ng29489  &  wire31290 ) ;
 assign ng34038 = ( wire31298 ) | ( ng28349  &  ng13486  &  wire31297 ) ;
 assign ng21899 = ( (~ pg35)  &  ng4291 ) | ( pg35  &  (~ pg9019)  &  ng4291 ) | ( pg35  &  pg9019  &  (~ ng4291) ) ;
 assign ng30391 = ( wire5603 ) | ( wire31317 ) | ( wire31318 ) | ( wire31319 ) ;
 assign ng29228 = ( wire5600 ) | ( wire5601 ) | ( (~ pg35)  &  ng736 ) ;
 assign ng25696 = ( wire5597 ) | ( wire31328 ) | ( wire31326  &  wire31327 ) ;
 assign ng34029 = ( wire5593 ) | ( wire31333 ) ;
 assign ng26929 = ( wire31337 ) | ( ng17625  &  (~ ng12377)  &  wire31334 ) ;
 assign ng30548 = ( wire5589 ) | ( (~ ng15039)  &  wire31338 ) | ( ng15039  &  wire31339 ) ;
 assign ng30364 = ( wire5586 ) | ( wire31346 ) | ( (~ ng25492)  &  wire31342 ) ;
 assign ng30431 = ( wire5580 ) | ( (~ ng11480)  &  wire31347 ) | ( ng11480  &  wire31348 ) ;
 assign ng33003 = ( wire5574 ) | ( wire31356 ) | ( (~ pg35)  &  ng2193 ) ;
 assign ng33014 = ( wire31363 ) | ( wire31364 ) ;
 assign ng25631 = ( wire31374 ) | ( (~ ng15748)  &  wire31367 ) | ( ng15748  &  wire31372 ) ;
 assign ng26916 = ( wire31380 ) | ( ng13307  &  wire31378 ) | ( ng10929  &  wire31378 ) ;
 assign ng24246 = ( (~ pg35)  &  ng1205 ) | ( pg35  &  ng1221  &  (~ ng1087) ) | ( pg35  &  ng1221  &  (~ ng1205) ) | ( pg35  &  (~ ng1221)  &  ng1087  &  ng1205 ) ;
 assign ng32987 = ( wire5555 ) | ( wire31390 ) | ( (~ pg35)  &  ng1632 ) ;
 assign ng33558 = ( wire5552 ) | ( wire5553 ) | ( (~ pg35)  &  ng1844 ) ;
 assign ng34468 = ( wire31398 ) | ( ng31009  &  (~ ng10862)  &  wire31397 ) ;
 assign ng34732 = ( (~ pg35)  &  ng2999 ) | ( pg35  &  ng2994 ) ;
 assign ng25626 = ( wire31403 ) | ( (~ ng10929)  &  (~ ng10909)  &  wire31400 ) ;
 assign ng33592 = ( wire5542 ) | ( ng28973  &  wire31406 ) ;
 assign ng25762 = ( (~ pg35)  &  ng6527 ) | ( ng6527  &  ng10887 ) | ( pg35  &  ng6533  &  (~ ng10887) ) ;
 assign ng25597 = ( (~ pg35)  &  ng358 ) | ( pg35  &  (~ ng370)  &  ng8721 ) | ( pg35  &  ng370  &  (~ ng8721) ) ;
 assign ng33986 = ( wire5533 ) | ( wire5534 ) | ( ng30304  &  wire31414 ) ;
 assign ng25690 = ( (~ pg35)  &  ng2841 ) | ( pg35  &  ng2837  &  (~ ng4125) ) ;
 assign ng29288 = ( (~ pg35)  &  ng5475 ) | ( ng5475  &  (~ ng23630) ) | ( pg35  &  ng5481  &  ng23630 ) ;
 assign ng33212 = ( wire30202 ) | ( wire30203 ) | ( wire30204 ) | ( wire30205 ) ;
 assign ng33586 = ( wire5524 ) | ( wire5525 ) | ( (~ pg35)  &  ng2331 ) ;
 assign ng30373 = ( wire5523 ) | ( wire31429 ) | ( (~ ng25435)  &  wire31425 ) ;
 assign ng29229 = ( wire31434 ) | ( (~ ng827)  &  wire31433 ) | ( ng20905  &  wire31433 ) ;
 assign ng34614 = ( (~ pg35)  &  ng37 ) | ( pg35  &  ng94 ) ;
 assign ng33611 = ( wire5512 ) | ( wire5513 ) | ( (~ pg35)  &  ng3698 ) ;
 assign ng33041 = ( wire31445 ) | ( wire31446 ) ;
 assign ng32997 = ( wire5503 ) | ( wire31452 ) | ( (~ pg35)  &  ng1932 ) ;
 assign ng29226 = ( wire5502 ) | ( (~ ng23324)  &  wire31454 ) | ( (~ ng23324)  &  wire31456 ) ;
 assign ng26966 = ( pg6748  &  pg35 ) | ( (~ pg35)  &  ng4555 ) ;
 assign ng34034 = ( (~ pg35)  &  ng4836 ) | ( ng4836  &  ng31009 ) ;
 assign ng24253 = ( wire31460 ) | ( pg35  &  pg7946  &  ng1521 ) ;
 assign ng26920 = ( wire31464 ) | ( ng13242  &  wire31463 ) | ( wire5491  &  wire31463 ) ;
 assign ng30369 = ( wire5487 ) | ( wire31470 ) | ( (~ ng25432)  &  wire31466 ) ;
 assign ng25721 = ( wire5483 ) | ( wire31477 ) | ( ng10838  &  wire31472 ) ;
 assign ng21891 = ( wire5476 ) | ( (~ pg35)  &  ng4180 ) ;
 assign ng30506 = ( wire5475 ) | ( (~ ng14996)  &  wire31478 ) | ( ng14996  &  wire31479 ) ;
 assign ng25747 = ( (~ pg35)  &  ng6163 ) | ( pg35  &  (~ ng6167)  &  ng10874 ) | ( pg35  &  ng6167  &  (~ ng10874) ) ;
 assign ng30440 = ( wire5469 ) | ( (~ ng14154)  &  wire31484 ) | ( ng14154  &  wire31485 ) ;
 assign ng33597 = ( wire5463 ) | ( wire5464 ) | ( wire5465 ) | ( wire5466 ) ;
 assign ng30475 = ( wire5462 ) | ( (~ ng14659)  &  wire31494 ) | ( ng14659  &  wire31495 ) ;
 assign ng33034 = ( wire5456 ) | ( (~ ng27635)  &  wire31498 ) | ( (~ ng27635)  &  wire31499 ) ;
 assign ng30472 = ( wire5451 ) | ( (~ ng14879)  &  wire31501 ) | ( ng14879  &  wire31502 ) ;
 assign ng34634 = ( (~ pg35)  &  ng4727 ) | ( pg35  &  ng4732 ) ;
 assign ng26890 = ( (~ pg35)  &  ng333 ) | ( pg35  &  (~ ng347) ) ;
 assign ng34797 = ( (~ pg91)  &  pg35 ) | ( (~ pg35)  &  ng2882 ) | ( pg35  &  ng2878 ) ;
 assign ng32982 = ( wire5438 ) | ( (~ pg35)  &  ng930 ) ;
 assign ng34629 = ( (~ pg35)  &  ng4146 ) | ( pg35  &  ng4157 ) ;
 assign ng33031 = ( (~ pg35)  &  ng3857 ) | ( ng3857  &  (~ ng3863)  &  (~ ng27635) ) | ( pg35  &  (~ ng3857)  &  ng3863  &  (~ ng27635) ) ;
 assign ng32989 = ( wire5430 ) | ( wire31512 ) | ( (~ pg35)  &  ng1664 ) ;
 assign ng28069 = ( wire5427 ) | ( wire31515 ) ;
 assign ng25615 = ( (~ pg35)  &  ng686 ) | ( ng686  &  ng11607 ) | ( pg35  &  ng667  &  (~ ng11607) ) ;
 assign ng25719 = ( (~ pg35)  &  ng5471 ) | ( pg35  &  (~ ng5475)  &  ng10838 ) | ( pg35  &  ng5475  &  (~ ng10838) ) ;
 assign ng30493 = ( wire5419 ) | ( (~ ng14927)  &  wire31521 ) | ( ng14927  &  wire31522 ) ;
 assign ng25639 = ( (~ pg35)  &  ng2715 ) | ( pg35  &  (~ ng2841) ) | ( ng2715  &  (~ ng2719) ) | ( pg35  &  (~ ng2715)  &  ng2719 ) ;
 assign ng30448 = ( wire5412 ) | ( (~ ng14142)  &  wire31527 ) | ( ng14142  &  wire31528 ) ;
 assign ng25593 = ( wire5406 ) | ( wire5407 ) | ( ng8359  &  wire31530 ) ;
 assign ng34254 = ( wire31533 ) | ( wire31534 ) | ( pg35  &  (~ ng33394) ) ;
 assign ng34631 = ( (~ pg35)  &  ng4253 ) | ( pg35  &  ng4249 ) ;
 assign ng30467 = ( wire5397 ) | ( (~ ng14683)  &  wire31536 ) | ( ng14683  &  wire31537 ) ;
 assign ng34465 = ( wire31543 ) | ( ng31009  &  (~ ng10862)  &  wire31542 ) ;
 assign ng33578 = ( wire5390 ) | ( wire31546 ) ;
 assign ng25702 = ( wire31550 ) | ( pg35  &  (~ pg9553)  &  ng5062 ) ;
 assign ng34650 = ( (~ ng25779)  &  ng34056  &  ng34051  &  ng34424 ) | ( ng25779  &  (~ ng34056)  &  ng34051  &  ng34424 ) | ( ng25779  &  ng34056  &  (~ ng34051)  &  ng34424 ) | ( (~ ng25779)  &  (~ ng34056)  &  (~ ng34051)  &  ng34424 ) | ( ng25779  &  ng34056  &  ng34051  &  (~ ng34424) ) | ( (~ ng25779)  &  (~ ng34056)  &  ng34051  &  (~ ng34424) ) | ( (~ ng25779)  &  ng34056  &  (~ ng34051)  &  (~ ng34424) ) | ( ng25779  &  (~ ng34056)  &  (~ ng34051)  &  (~ ng34424) ) ;
 assign ng24202 = ( (~ pg35)  &  ng411 ) | ( ng411  &  (~ ng8806) ) | ( pg35  &  ng424  &  ng8806 ) ;
 assign ng26919 = ( wire31555 ) | ( (~ ng19140)  &  wire31553 ) ;
 assign ng28049 = ( wire5376 ) | ( (~ ng20248)  &  wire31556 ) | ( ng20248  &  wire31557 ) ;
 assign ng33998 = ( wire5372 ) | ( wire5373 ) | ( ng30300  &  wire31559 ) ;
 assign ng26913 = ( wire31565 ) | ( ng13211  &  wire31564 ) | ( wire5848  &  wire31564 ) ;
 assign ng28059 = ( wire5365 ) | ( wire5366 ) | ( (~ pg35)  &  ng1351 ) ;
 assign ng24342 = ( (~ pg35)  &  ng5689 ) | ( pg35  &  (~ ng5689)  &  (~ ng5698) ) | ( pg35  &  (~ ng5698)  &  ng10160 ) ;
 assign ng34010 = ( wire5361 ) | ( wire5362 ) | ( ng30314  &  wire31571 ) ;
 assign ng28096 = ( wire5357 ) | ( wire5358 ) | ( (~ pg35)  &  ng5619 ) ;
 assign ng24273 = ( (~ pg35)  &  ng3689 ) | ( pg35  &  (~ ng3689)  &  (~ ng3698) ) | ( pg35  &  (~ ng3698)  &  ng8728 ) ;
 assign ng26928 = ( wire31581 ) | ( ng17625  &  (~ ng12377)  &  wire31578 ) ;
 assign ng25596 = ( (~ pg35)  &  ng370 ) | ( pg35  &  (~ ng358)  &  ng376 ) | ( pg35  &  ng358  &  (~ ng376) ) ;
 assign ng28056 = ( wire31587 ) | ( ng907  &  ng22992  &  (~ ng19063) ) ;
 assign ng28053 = ( wire31589 ) | ( pg35  &  (~ ng20248) ) ;
 assign ng29260 = ( wire5342 ) | ( wire31595 ) | ( (~ ng23067)  &  wire31591 ) ;
 assign ng34261 = ( wire5338 ) | ( wire31600 ) | ( (~ ng29657)  &  wire31596 ) ;
 assign ng24345 = ( (~ pg35)  &  ng6031 ) | ( pg35  &  ng6035  &  ng10185 ) | ( pg35  &  (~ ng6035)  &  (~ ng10185) ) ;
 assign ng30458 = ( wire31604 ) | ( pg113  &  ng4473  &  (~ ng4459) ) ;
 assign ng24276 = ( (~ pg35)  &  ng4031 ) | ( pg35  &  ng4040  &  ng8751 ) | ( pg35  &  (~ ng4040)  &  (~ ng8751) ) ;
 assign ng30483 = ( wire31610 ) | ( (~ ng12453)  &  wire31609 ) | ( (~ ng12558)  &  wire31609 ) ;
 assign ng32978 = ( wire5319 ) | ( (~ ng27629)  &  wire31612 ) | ( ng27629  &  wire31613 ) ;
 assign ng33976 = ( wire5315 ) | ( wire5316 ) | ( ng30298  &  wire31616 ) ;
 assign ng34729 = ( pg35  &  (~ ng1306) ) | ( pg35  &  ng1296 ) | ( (~ pg35)  &  ng1291 ) ;
 assign ng26947 = ( wire5308 ) | ( wire5309 ) | ( wire31623 ) ;
 assign ng25625 = ( pg35  &  (~ ng979)  &  ng1052  &  ng13121 ) | ( pg35  &  (~ ng979)  &  (~ ng1052)  &  (~ ng13121) ) ;
 assign ng33552 = ( wire5304 ) | ( ng28892  &  wire31631 ) ;
 assign ng25622 = ( wire5299 ) | ( wire31642 ) | ( ng15737  &  wire31640 ) ;
 assign ng26892 = ( (~ pg35)  &  ng351 ) | ( pg35  &  ng333  &  (~ ng351) ) | ( pg35  &  ng355  &  (~ ng351) ) ;
 assign ng25757 = ( pg35  &  ng6727 ) | ( (~ pg35)  &  ng6444 ) ;
 assign ng26901 = ( wire5294 ) | ( (~ ng10632)  &  wire31645 ) | ( ng10632  &  wire31646 ) ;
 assign ng33058 = ( (~ pg35)  &  ng5863 ) | ( (~ ng28020)  &  wire31650 ) ;
 assign ng33534 = ( wire5289 ) | ( (~ ng28353)  &  wire31652 ) | ( ng28353  &  wire31653 ) ;
 assign ng26932 = ( wire31658 ) | ( ng17625  &  (~ ng12377)  &  wire31655 ) ;
 assign ng33035 = ( wire31662 ) | ( (~ ng4098)  &  wire31660 ) | ( (~ ng22654)  &  wire31660 ) ;
 assign ng33060 = ( wire5279 ) | ( (~ ng28020)  &  wire31664 ) | ( (~ ng28020)  &  wire31665 ) ;
 assign ng24233 = ( wire5276 ) | ( (~ ng10909)  &  wire31667 ) | ( ng10909  &  wire31668 ) ;
 assign ng25612 = ( wire5273 ) | ( ng11607  &  wire31671 ) | ( (~ ng11607)  &  wire31672 ) ;
 assign ng24335 = ( (~ pg35)  &  ng66 ) | ( wire31677  &  wire31678 ) ;
 assign ng31900 = ( wire5258 ) | ( wire5259 ) | ( (~ pg35)  &  ng5037 ) ;
 assign ng34624 = ( (~ pg35)  &  ng2994 ) | ( pg35  &  ng2988 ) ;
 assign ng30345 = ( wire31686 ) | ( pg35  &  ng24609 ) ;
 assign ng26895 = ( wire31690 ) | ( ng14708  &  (~ wire28793)  &  wire31689 ) ;
 assign ng21900 = ( (~ pg35)  &  ng4239 ) | ( pg35  &  (~ pg10122)  &  (~ ng4297) ) ;
 assign ng33045 = ( wire31696 ) | ( wire31697 ) ;
 assign ng25744 = ( wire31701 ) | ( pg35  &  (~ pg9741)  &  ng6098 ) ;
 assign ng30532 = ( wire5231 ) | ( (~ ng14899)  &  wire31702 ) | ( ng14899  &  wire31703 ) ;
 assign ng25708 = ( (~ pg35)  &  ng5156 ) | ( ng5156  &  ng10823 ) | ( pg35  &  ng5120  &  (~ ng10823) ) ;
 assign ng24257 = ( (~ pg35)  &  ng1333 ) | ( ng1333  &  (~ ng16272) ) | ( pg35  &  (~ ng1333)  &  ng16272 ) ;
 assign ng34450 = ( wire31715 ) | ( (~ ng30583)  &  ng15591  &  wire31714 ) ;
 assign ng30471 = ( wire5214 ) | ( (~ ng14841)  &  wire31716 ) | ( ng14841  &  wire31717 ) ;
 assign ng33542 = ( wire5209 ) | ( wire5210 ) | ( (~ pg35)  &  ng1270 ) ;
 assign ng31904 = ( wire31731 ) | ( (~ wire29550)  &  (~ wire29551)  &  wire31729 ) ;
 assign ng28088 = ( wire31746 ) | ( wire31747 ) | ( wire31748 ) ;
 assign ng25698 = ( (~ pg35)  &  ng5092 ) | ( pg35  &  (~ ng5092)  &  ng5097 ) | ( pg35  &  (~ ng5084)  &  ng5097 ) | ( pg35  &  ng5092  &  ng5084  &  (~ ng5097) ) ;
 assign ng34728 = ( ng19402 ) | ( (~ pg35)  &  ng939 ) | ( pg35  &  ng943 ) ;
 assign ng30461 = ( wire31756 ) | ( (~ ng12772)  &  wire31755 ) | ( (~ ng12492)  &  wire31755 ) ;
 assign ng34618 = ( pg35  &  ng2912 ) | ( (~ pg35)  &  ng2907 ) ;
 assign ng33609 = ( wire5176 ) | ( wire5177 ) | ( (~ pg35)  &  ng3347 ) ;
 assign ng29259 = ( (~ pg35)  &  ng3119 ) | ( ng3119  &  (~ ng23067) ) | ( pg35  &  ng3125  &  ng23067 ) ;
 assign ng30361 = ( (~ pg35)  &  ng1982 ) | ( ng1982  &  (~ ng25341) ) | ( pg35  &  ng1988  &  ng25341 ) ;
 assign ng24338 = ( (~ pg35)  &  ng5343 ) | ( pg35  &  (~ ng5343)  &  (~ ng5352) ) | ( pg35  &  (~ ng5352)  &  ng10124 ) ;
 assign ng26958 = ( wire6028 ) | ( wire6029 ) | ( (~ pg35)  &  ng4455 ) ;
 assign ng33981 = ( wire5164 ) | ( wire5165 ) | ( ng30304  &  wire31771 ) ;
 assign ng30381 = ( (~ pg35)  &  ng2541 ) | ( ng2541  &  (~ ng25400) ) | ( pg35  &  ng2547  &  ng25400 ) ;
 assign ng24337 = ( (~ pg35)  &  ng5339 ) | ( pg35  &  ng5343  &  ng10124 ) | ( pg35  &  (~ ng5343)  &  (~ ng10124) ) ;
 assign ng30499 = ( wire5156 ) | ( (~ ng14807)  &  wire31779 ) | ( ng14807  &  wire31780 ) ;
 assign ng24239 = ( wire31783 ) | ( pg35  &  pg12919  &  pg17400 ) ;
 assign ng26897 = ( wire5148 ) | ( wire5149 ) | ( (~ pg35)  &  ng732 ) ;
 assign ng26891 = ( (~ pg35)  &  ng347 ) | ( pg35  &  pg7540  &  (~ ng347) ) ;
 assign ng33024 = ( wire5145 ) | ( (~ ng27602)  &  wire31788 ) | ( (~ ng27602)  &  wire31789 ) ;
 assign ng34447 = ( wire31797 ) | ( pg35  &  ng29503  &  wire31794 ) ;
 assign ng33971 = ( wire31803 ) | ( (~ ng29482)  &  wire31799 ) | ( ng29482  &  wire31801 ) ;
 assign ng29295 = ( wire5132 ) | ( wire31811 ) | ( (~ ng23666)  &  wire31806 ) ;
 assign ng30402 = ( wire5128 ) | ( (~ ng13948)  &  wire31812 ) | ( ng13948  &  wire31813 ) ;
 assign ng26961 = ( pg6748  &  pg35 ) | ( (~ pg35)  &  ng4483 ) ;
 assign ng30487 = ( wire5123 ) | ( (~ ng14688)  &  wire31815 ) | ( ng14688  &  wire31816 ) ;
 assign ng30552 = ( wire5120 ) | ( (~ ng14905)  &  wire31818 ) | ( ng14905  &  wire31819 ) ;
 assign ng25677 = ( (~ pg35)  &  ng3752 ) | ( pg35  &  ng4040 ) ;
 assign ng26949 = ( wire31822 ) | ( wire29325  &  wire29326  &  wire31821 ) ;
 assign ng26967 = ( pg6750  &  pg35 ) | ( (~ pg35)  &  ng4561 ) ;
 assign ng33018 = ( wire31829 ) | ( wire31830 ) ;
 assign ng30452 = ( wire5103 ) | ( (~ ng11534)  &  wire31831 ) | ( ng11534  &  wire31832 ) ;
 assign ng34611 = ( (~ pg35)  &  ng2852 ) | ( pg35  &  ng2860 ) ;
 assign ng30556 = ( wire5098 ) | ( (~ ng15033)  &  wire31834 ) | ( ng15033  &  wire31835 ) ;
 assign ng30415 = ( wire31840 ) | ( (~ ng8906)  &  wire31839 ) | ( (~ ng11571)  &  wire31839 ) ;
 assign ng29307 = ( wire5089 ) | ( wire31847 ) | ( (~ ng23733)  &  wire31842 ) ;
 assign ng30413 = ( wire5085 ) | ( (~ ng14011)  &  wire31848 ) | ( ng14011  &  wire31849 ) ;
 assign ng30433 = ( wire5082 ) | ( (~ ng14018)  &  wire31851 ) | ( ng14018  &  wire31852 ) ;
 assign ng30511 = ( wire5079 ) | ( (~ ng14855)  &  wire31854 ) | ( ng14855  &  wire31855 ) ;
 assign ng28086 = ( wire31871 ) | ( wire31872 ) | ( wire31873 ) ;
 assign ng34039 = ( wire31879 ) | ( ng28349  &  ng13486  &  wire31878 ) ;
 assign ng30340 = ( wire5067 ) | ( (~ ng24591)  &  wire31881 ) | ( (~ ng24591)  &  wire31883 ) ;
 assign ng30512 = ( wire5064 ) | ( (~ ng14892)  &  wire31885 ) | ( ng14892  &  wire31886 ) ;
 assign ng24234 = ( (~ pg35)  &  ng1146 ) | ( ng1146  &  (~ ng10909) ) | ( pg35  &  ng1152  &  ng10909 ) ;
 assign ng34793 = ( wire31902 ) | ( pg35  &  ng17657 ) | ( pg35  &  ng17700 ) ;
 assign ng24241 = ( (~ pg35)  &  ng990 ) | ( ng990  &  (~ ng16246) ) | ( pg35  &  (~ ng990)  &  ng16246 ) ;
 assign ng30359 = ( wire5036 ) | ( wire31910 ) | ( (~ ng25467)  &  wire31906 ) ;
 assign ng33176 = ( wire29971 ) | ( wire29972 ) | ( wire30013 ) | ( wire30014 ) ;
 assign ng33047 = ( (~ pg35)  &  ng5164 ) | ( (~ ng5170)  &  ng5164  &  (~ ng27999) ) | ( pg35  &  ng5170  &  (~ ng5164)  &  (~ ng27999) ) ;
 assign ng25638 = ( wire31917 ) | ( (~ ng11171)  &  ng11149  &  wire31915 ) ;
 assign ng34466 = ( wire31921 ) | ( ng31009  &  (~ ng10862)  &  wire31920 ) ;
 assign ng30563 = ( wire5018 ) | ( (~ ng14984)  &  wire31922 ) | ( ng14984  &  wire31923 ) ;
 assign ng34612 = ( (~ pg35)  &  ng2860 ) | ( pg35  &  ng2894 ) ;
 assign ng34449 = ( (~ ng30583)  &  ng15591  &  wire31926 ) | ( (~ ng30583)  &  ng15591  &  wire31928 ) ;
 assign ng30400 = ( wire5011 ) | ( (~ ng13889)  &  wire31929 ) | ( ng13889  &  wire31930 ) ;
 assign ng30407 = ( wire5008 ) | ( (~ ng14101)  &  wire31932 ) | ( ng14101  &  wire31933 ) ;
 assign ng30500 = ( wire5005 ) | ( (~ ng14851)  &  wire31935 ) | ( ng14851  &  wire31936 ) ;
 assign ng34911 = ( wire5002 ) | ( (~ ng34703)  &  wire31942 ) | ( ng34703  &  wire31943 ) ;
 assign ng32994 = ( wire31951 ) | ( wire31952 ) ;
 assign ng34035 = ( (~ pg35)  &  ng4864 ) | ( ng4864  &  ng31009 ) ;
 assign ng34259 = ( wire4993 ) | ( (~ ng11320)  &  (~ ng31950)  &  wire30570 ) ;
 assign ng34800 = ( pg35  &  ng34 ) | ( pg35  &  ng2980 ) | ( (~ pg35)  &  ng2886 ) ;
 assign ng30504 = ( wire31956 ) | ( (~ ng12609)  &  wire31955 ) | ( (~ ng12515)  &  wire31955 ) ;
 assign ng24210 = ( (~ ng13756)  &  wire31958 ) | ( (~ ng13756)  &  wire31960 ) | ( (~ ng13756)  &  wire31962 ) ;
 assign ng34462 = ( wire31967 ) | ( ng31003  &  (~ ng10831)  &  wire31966 ) ;
 assign ng26915 = ( wire31972 ) | ( ng10929  &  wire31970 ) | ( ng13260  &  wire31970 ) ;
 assign ng30436 = ( wire31975 ) | ( ng11626  &  ng8958  &  wire31974 ) ;
 assign ng31894 = ( wire31978 ) | ( pg35  &  (~ ng4098)  &  ng22654 ) | ( pg35  &  ng4098  &  (~ ng22654) ) ;
 assign ng33039 = ( wire31984 ) | ( wire31985 ) ;
 assign ng24261 = ( pg35  &  pg12923 ) | ( (~ pg35)  &  ng1585 ) ;
 assign ng33623 = ( wire4958 ) | ( (~ ng29036)  &  wire31989 ) | ( (~ ng29036)  &  wire31991 ) ;
 assign ng30530 = ( wire4955 ) | ( (~ ng14817)  &  wire31993 ) | ( ng14817  &  wire31994 ) ;
 assign ng30524 = ( wire31998 ) | ( (~ ng10421)  &  wire31997 ) | ( (~ ng12667)  &  wire31997 ) ;
 assign ng25716 = ( wire32002 ) | ( pg35  &  (~ pg9615)  &  ng5406 ) ;
 assign ng32976 = ( wire4944 ) | ( wire4945 ) | ( (~ pg35)  &  ng164 ) ;
 assign ng34719 = ( pg35  &  ng209 ) | ( pg35  &  ng538 ) ;
 assign ng34262 = ( wire4941 ) | ( wire32011 ) | ( ng29672  &  wire32007 ) ;
 assign ng30485 = ( wire4937 ) | ( (~ ng14956)  &  wire32012 ) | ( ng14956  &  wire32013 ) ;
 assign ng30460 = ( wire32017 ) | ( (~ ng10266)  &  wire32016 ) | ( (~ ng12492)  &  wire32016 ) ;
 assign ng33009 = ( wire4929 ) | ( wire32022 ) | ( (~ pg35)  &  ng2357 ) ;
 assign ng26956 = ( ng4452 ) | ( (~ ng4443)  &  (~ ng4452)  &  wire29521  &  wire32024 ) ;
 assign ng33536 = ( wire7582 ) | ( (~ pg35)  &  ng160 ) ;
 assign ng32980 = ( wire4912 ) | ( (~ ng23975)  &  wire32052 ) | ( wire32051  &  wire32052 ) ;
 assign ng29253 = ( wire4908 ) | ( wire4909 ) | ( wire32058 ) ;
 assign ng34456 = ( wire4906 ) | ( ng28144  &  wire32061 ) | ( (~ ng28144)  &  wire32063 ) ;
 assign ng30379 = ( wire4903 ) | ( wire32070 ) | ( (~ ng25495)  &  wire32066 ) ;
 assign ng30382 = ( wire4899 ) | ( wire32077 ) | ( (~ ng25400)  &  wire32072 ) ;
 assign ng34018 = ( wire4893 ) | ( wire4895 ) | ( ng29313  &  wire32080 ) ;
 assign ng30443 = ( wire4892 ) | ( (~ ng13990)  &  wire32082 ) | ( ng13990  &  wire32083 ) ;
 assign ng33988 = ( wire4888 ) | ( wire4889 ) | ( ng30311  &  wire32086 ) ;
 assign ng34265 = ( ng31009  &  (~ ng10862)  &  wire32091 ) ;
 assign ng33572 = ( wire4884 ) | ( wire4885 ) | ( (~ pg35)  &  ng2102 ) ;
 assign ng34016 = ( wire4882 ) | ( wire4883 ) | ( ng29313  &  wire32096 ) ;
 assign ng29247 = ( wire4878 ) | ( wire4879 ) | ( wire32103 ) ;
 assign ng25637 = ( wire32109 ) | ( (~ ng11171)  &  ng13597  &  wire32107 ) ;
 assign ng30397 = ( wire32112 ) | ( ng11473  &  ng11514  &  wire32111 ) ;
 assign ng30351 = ( (~ pg35)  &  ng1714 ) | ( ng1714  &  (~ ng25275) ) | ( pg35  &  ng1720  &  ng25275 ) ;
 assign ng26918 = ( wire4861 ) | ( wire4863 ) | ( wire32118 ) ;
 assign ng30408 = ( wire4860 ) | ( (~ ng14127)  &  wire32120 ) | ( ng14127  &  wire32121 ) ;
 assign ng30503 = ( wire32125 ) | ( (~ ng12609)  &  wire32124 ) | ( (~ ng12824)  &  wire32124 ) ;
 assign ng24298 = ( (~ pg35)  &  ng4392 ) ;
 assign ng25742 = ( pg35  &  ng6227 ) ;
 assign ng25635 = ( wire32130 ) | ( ng10939  &  wire32127 ) | ( ng10961  &  wire32127 ) ;
 assign ng33044 = ( wire4842 ) | ( wire4843 ) | ( wire32133 ) ;
 assign ng30394 = ( wire32137 ) | ( (~ ng8864)  &  wire32136 ) | ( (~ ng11514)  &  wire32136 ) ;
 assign ng33568 = ( wire4836 ) | ( ng28962  &  wire32141 ) ;
 assign ng24271 = ( wire4834 ) | ( ng8728  &  wire32145  &  wire32146 ) ;
 assign ng33963 = ( wire4827 ) | ( wire4828 ) | ( wire32166 ) | ( wire32167 ) ;
 assign ng34636 = ( pg35  &  ng4722 ) | ( (~ pg35)  &  ng4717 ) ;
 assign ng29298 = ( wire4795 ) | ( wire4796 ) | ( wire4797 ) | ( wire4798 ) ;
 assign ng30474 = ( wire4794 ) | ( ng14953  &  wire32234 ) | ( (~ ng14953)  &  wire32235 ) ;
 assign ng34625 = ( pg35  &  ng3151 ) ;
 assign ng34798 = ( pg35  &  ng2946 ) | ( (~ pg35)  &  ng2878 ) | ( pg35  &  ng2886 ) ;
 assign ng24350 = ( (~ pg35)  &  ng6381 ) | ( pg35  &  (~ ng6381)  &  (~ ng6390) ) | ( pg35  &  (~ ng6390)  &  ng10207 ) ;
 assign ng33613 = ( wire32244 ) | ( (~ ng28484)  &  wire32242 ) ;
 assign ng29265 = ( (~ pg35)  &  ng3470 ) | ( ng3470  &  (~ ng23112) ) | ( pg35  &  ng3476  &  ng23112 ) ;
 assign ng29276 = ( wire4757 ) | ( wire32304 ) | ( wire32305 ) | ( wire32306 ) ;
 assign ng33059 = ( (~ pg35)  &  ng5869 ) | ( ng5869  &  (~ ng5873)  &  (~ ng28020) ) | ( pg35  &  (~ ng5869)  &  ng5873  &  (~ ng28020) ) ;
 assign ng29278 = ( wire4749 ) | ( wire30550 ) | ( wire30551 ) | ( wire30552 ) ;
 assign ng34253 = ( pg35  &  (~ ng4467) ) | ( pg35  &  (~ ng4462) ) | ( pg35  &  (~ ng33394) ) ;
 assign ng30542 = ( wire4745 ) | ( (~ ng14943)  &  wire32313 ) | ( ng14943  &  wire32314 ) ;
 assign ng28102 = ( wire4740 ) | ( wire4741 ) | ( (~ pg35)  &  ng6311 ) ;
 assign ng24268 = ( (~ pg35)  &  ng3329 ) | ( pg35  &  ng3338  &  ng8691 ) | ( pg35  &  (~ ng3338)  &  (~ ng8691) ) ;
 assign ng30349 = ( wire4736 ) | ( wire32327 ) | ( (~ ng25382)  &  wire32323 ) ;
 assign ng33219 = ( wire30215 ) | ( wire30216 ) | ( wire30231 ) | ( wire30232 ) ;
 assign ng30422 = ( wire4729 ) | ( ng13955  &  wire32328 ) | ( (~ ng13955)  &  wire32329 ) ;
 assign ng33587 = ( wire4724 ) | ( wire4725 ) | ( (~ pg35)  &  ng2375 ) ;
 assign ng33603 = ( wire4721 ) | ( wire4722 ) | ( (~ pg35)  &  ng2643 ) ;
 assign ng26888 = ( pg35  &  ng316 ) | ( (~ pg35)  &  ng106 ) ;
 assign ng34453 = ( wire4715 ) | ( (~ ng31997)  &  wire32336 ) | ( (~ ng31997)  &  wire32338 ) ;
 assign ng34021 = ( wire4711 ) | ( wire4712 ) | ( ng29313  &  wire32340 ) ;
 assign ng34440 = ( wire32353 ) | ( ng23975  &  (~ wire32051)  &  wire32344 ) ;
 assign ng34794 = ( (~ pg35)  &  ng2856 ) | ( pg35  &  ng2864 ) | ( pg35  &  ng28220 ) ;
 assign ng33164 = ( wire30095 ) | ( wire30096 ) | ( wire30115 ) | ( wire30116 ) ;
 assign ng26968 = ( pg6749  &  pg35 ) | ( (~ pg35)  &  ng4558 ) ;
 assign ng29285 = ( pg35  &  ng4284  &  (~ ng14211) ) | ( pg35  &  (~ ng4180)  &  (~ ng14211) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng14211 ) ;
 assign ng33582 = ( wire4692 ) | ( wire4693 ) | ( (~ pg35)  &  ng2269 ) ;
 assign ng24231 = ( pg35  &  pg12919  &  (~ ng904) ) ;
 assign ng33065 = ( wire4689 ) | ( (~ ng26977)  &  wire32367 ) | ( (~ ng26977)  &  wire32368 ) ;
 assign ng30522 = ( pg35  &  (~ ng6215)  &  (~ ng6203)  &  (~ ng26977) ) ;
 assign ng24334 = ( wire4685 ) | ( (~ pg35)  &  ng4358 ) ;
 assign ng34000 = ( wire4683 ) | ( wire4684 ) | ( ng30300  &  wire32382 ) ;
 assign ng28071 = ( wire32387 ) | ( ng4145  &  ng13806  &  (~ wire32385) ) ;
 assign ng33566 = ( wire4676 ) | ( wire4677 ) | ( (~ pg35)  &  ng1978 ) ;
 assign ng34635 = ( (~ pg35)  &  ng4732 ) | ( pg35  &  ng4717 ) ;
 assign ng30398 = ( wire4673 ) | ( ng14098  &  wire32391 ) | ( (~ ng14098)  &  wire32392 ) ;
 assign ng31871 = ( wire32396 ) | ( ng25917  &  wire32395 ) | ( wire4669  &  wire32395 ) ;
 assign ng33000 = ( wire4663 ) | ( wire32401 ) | ( (~ pg35)  &  ng2028 ) ;
 assign ng29241 = ( wire4659 ) | ( wire4660 ) | ( wire32406 ) ;
 assign ng29234 = ( wire4652 ) | ( wire4653 ) | ( wire32423 ) | ( wire32424 ) ;
 assign ng25733 = ( (~ pg35)  &  ng5817 ) | ( pg35  &  (~ ng5821)  &  ng10869 ) | ( pg35  &  ng5821  &  (~ ng10869) ) ;
 assign ng29222 = ( wire32434 ) | ( (~ ng23975)  &  wire32431 ) | ( ng23975  &  wire32432 ) ;
 assign ng25686 = ( (~ pg35)  &  ng4064 ) | ( pg35  &  ng2841  &  (~ ng4064)  &  ng4057 ) | ( pg35  &  ng2841  &  ng4064  &  (~ ng4057) ) ;
 assign ng30385 = ( (~ pg35)  &  ng2657 ) | ( pg35  &  ng2661  &  ng25439 ) | ( pg35  &  (~ ng2661)  &  (~ ng25439) ) ;
 assign ng34623 = ( (~ pg35)  &  ng2960 ) | ( pg35  &  ng2970 ) ;
 assign ng34457 = ( wire4633 ) | ( (~ ng31950)  &  wire32443 ) | ( (~ ng31950)  &  wire32445 ) ;
 assign ng34441 = ( wire32453 ) | ( pg35  &  ng29503  &  wire32450 ) ;
 assign ng30420 = ( wire4626 ) | ( ng13898  &  wire32454 ) | ( (~ ng13898)  &  wire32455 ) ;
 assign ng34790 = ( wire32460 ) | ( ng33851  &  (~ wire30331)  &  wire32459 ) ;
 assign ng34627 = ( pg35  &  ng3853 ) ;
 assign ng34806 = ( wire32462 ) | ( pg35  &  ng4072 ) | ( pg35  &  ng2941 ) ;
 assign ng34637 = ( (~ pg35)  &  ng4722 ) | ( pg35  &  ng4737 ) ;
 assign ng34263 = ( wire4608 ) | ( wire32468 ) | ( ng29694  &  wire32464 ) ;
 assign ng34041 = ( wire32473 ) | ( ng28349  &  ng13486  &  wire32472 ) ;
 assign ng28090 = ( wire4596 ) | ( wire4598 ) | ( wire32488 ) | ( wire32489 ) ;
 assign ng25669 = ( wire4595 ) | ( wire32498 ) | ( ng12692  &  wire32493 ) ;
 assign ng28084 = ( wire32513 ) | ( wire32514 ) | ( wire32515 ) ;
 assign ng33593 = ( wire4583 ) | ( wire4584 ) | ( (~ pg35)  &  ng2472 ) ;
 assign ng34638 = ( pg35  &  ng4917 ) ;
 assign ng33975 = ( wire4581 ) | ( wire4582 ) | ( ng30298  &  wire32522 ) ;
 assign ng25648 = ( pg35  &  ng3179 ) ;
 assign ng32979 = ( wire4577 ) | ( wire4578 ) | ( (~ pg35)  &  ng749 ) ;
 assign ng24242 = ( pg35  &  ng102 ) | ( (~ pg35)  &  ng1211 ) ;
 assign ng32990 = ( wire32535 ) | ( wire32536 ) ;
 assign ng26894 = ( wire32541 ) | ( (~ ng20000)  &  wire32540 ) ;
 assign ng34792 = ( (~ pg35)  &  ng94 ) | ( pg35  &  ng2848 ) | ( pg35  &  ng22585 ) ;
 assign ng24262 = ( (~ pg35)  &  ng1548 ) | ( pg35  &  (~ ng1548)  &  ng1564 ) | ( pg35  &  ng1564  &  (~ ng1430) ) | ( pg35  &  ng1548  &  (~ ng1564)  &  ng1430 ) ;
 assign ng25627 = ( wire4550 ) | ( ng13284  &  wire32550 ) | ( (~ ng13284)  &  wire32551 ) ;
 assign ng29272 = ( wire4538 ) | ( wire4539 ) | ( wire4540 ) | ( wire4541 ) ;
 assign ng34033 = ( wire32563 ) | ( ng28336  &  ng13464  &  wire32562 ) ;
 assign ng29292 = ( wire4531 ) | ( wire4532 ) | ( wire4533 ) | ( wire4534 ) ;
 assign ng33984 = ( wire4528 ) | ( wire4530 ) | ( ng30304  &  wire32572 ) ;
 assign ng24213 = ( pg64  &  pg35 ) | ( (~ pg35)  &  ng753 ) ;
 assign ng30518 = ( wire4525 ) | ( (~ ng12512)  &  wire32574 ) | ( ng12512  &  wire32575 ) ;
 assign ng30456 = ( wire4517 ) | ( wire4518 ) | ( (~ pg35)  &  ng4087 ) ;
 assign ng33017 = ( wire4514 ) | ( wire32586 ) | ( (~ pg35)  &  ng2625 ) ;
 assign ng28052 = ( (~ pg35)  &  ng718 ) | ( ng718  &  (~ ng20248) ) | ( pg35  &  ng661  &  ng20248 ) ;
 assign ng30347 = ( wire4509 ) | ( (~ ng24609)  &  wire32590 ) | ( (~ ng24609)  &  wire32592 ) ;
 assign ng34004 = ( wire4505 ) | ( wire4506 ) | ( ng30307  &  wire32595 ) ;
 assign ng34850 = ( wire32601 ) | ( (~ ng34162)  &  wire31938  &  wire32600 ) ;
 assign ng33604 = ( wire4494 ) | ( wire4495 ) | ( (~ pg35)  &  ng2661 ) ;
 assign ng33600 = ( wire4493 ) | ( ng29001  &  wire32606 ) ;
 assign ng26969 = ( (~ pg35)  &  ng4462 ) | ( pg35  &  (~ ng4473)  &  (~ ng4467) ) ;
 assign ng33969 = ( wire4488 ) | ( wire4489 ) | ( ng30293  &  wire32609 ) ;
 assign ng26880 = ( pg6745  &  pg35 ) ;
 assign ng26902 = ( wire4486 ) | ( (~ ng10632)  &  wire32612 ) | ( ng10632  &  wire32613 ) ;
 assign ng34599 = ( wire4477 ) | ( wire4478 ) | ( (~ pg35)  &  ng608 ) ;
 assign ng25617 = ( wire32623 ) | ( ng8806  &  (~ ng14279)  &  wire32621 ) ;
 assign ng25614 = ( wire4466 ) | ( wire4467 ) | ( (~ ng11607)  &  wire32624 ) ;
 assign ng26962 = ( pg6749  &  pg35 ) | ( (~ pg35)  &  ng4486 ) ;
 assign ng34269 = ( wire4462 ) | ( wire32632 ) | ( (~ ng29737)  &  wire32628 ) ;
 assign ng33606 = ( wire4456 ) | ( wire4457 ) | ( (~ pg35)  &  ng2671 ) ;
 assign ng33596 = ( wire4445 ) | ( wire4446 ) | ( (~ pg35)  &  ng2527 ) ;
 assign ng34620 = ( (~ pg35)  &  ng2922 ) | ( pg35  &  ng2936 ) ;
 assign ng30536 = ( wire4439 ) | ( ng15024  &  wire32638 ) | ( (~ ng15024)  &  wire32639 ) ;
 assign ng26882 = ( (~ pg35)  &  ng316 ) | ( pg35  &  ng305 ) | ( pg35  &  ng311 ) ;
 assign ng25632 = ( wire4430 ) | ( wire32647 ) | ( (~ ng15748)  &  wire32642 ) ;
 assign ng28054 = ( (~ pg35)  &  ng661 ) | ( ng661  &  (~ ng20248) ) | ( pg35  &  ng728  &  ng20248 ) ;
 assign ng33992 = ( wire32656 ) | ( (~ ng29495)  &  wire32652 ) | ( ng29495  &  wire32654 ) ;
 assign ng28048 = ( wire4415 ) | ( wire32664 ) ;
 assign ng24343 = ( (~ pg35)  &  ng5694 ) | ( (~ ng5689)  &  ng5694 ) | ( ng5694  &  ng10160 ) ;
 assign ng26964 = ( wire32667 ) | ( (~ ng4527)  &  ng12228  &  wire32665 ) | ( ng4527  &  (~ ng12228)  &  wire32665 ) ;
 assign ng33982 = ( wire4404 ) | ( wire4406 ) | ( ng30304  &  wire32670 ) ;
 assign ng33625 = ( wire4403 ) | ( (~ ng29073)  &  wire32675 ) | ( (~ ng29073)  &  wire32677 ) ;
 assign ng29282 = ( (~ pg35)  &  ng5128 ) | ( ng5128  &  (~ ng23590) ) | ( pg35  &  ng5134  &  ng23590 ) ;
 assign ng28070 = ( wire32683 ) | ( pg35  &  ng4076  &  ng13217 ) | ( pg35  &  (~ ng4076)  &  (~ ng13217) ) ;
 assign ng24250 = ( (~ pg35)  &  ng1489 ) | ( ng1489  &  (~ ng10939) ) | ( pg35  &  ng1495  &  ng10939 ) ;
 assign ng34643 = ( pg35  &  ng5160 ) ;
 assign ng24237 = ( wire32689 ) | ( pg35  &  (~ pg7916)  &  ng1189 ) ;
 assign ng24206 = ( (~ pg35)  &  ng441 ) | ( ng441  &  (~ ng8806) ) | ( pg35  &  ng437  &  ng8806 ) ;
 assign ng30480 = ( pg35  &  (~ ng5523)  &  (~ ng5511)  &  (~ ng28010) ) ;
 assign ng30455 = ( wire4378 ) | ( ng14085  &  wire32694 ) | ( (~ ng14085)  &  wire32695 ) ;
 assign ng25748 = ( (~ pg35)  &  ng6181 ) | ( ng6181  &  ng10874 ) | ( pg35  &  ng6187  &  (~ ng10874) ) ;
 assign ng30336 = ( wire4367 ) | ( wire4368 ) | ( (~ pg35)  &  ng911 ) ;
 assign ng30497 = ( wire4366 ) | ( (~ ng12450)  &  wire32702 ) | ( ng12450  &  wire32703 ) ;
 assign ng32986 = ( wire4359 ) | ( wire32707 ) ;
 assign ng34880 = ( wire4355 ) | ( ng34550  &  wire32710 ) | ( (~ ng34550)  &  wire32711 ) ;
 assign ng24245 = ( pg35  &  pg12919 ) | ( (~ pg35)  &  ng1242 ) ;
 assign ng33037 = ( wire32717 ) | ( wire32718 ) ;
 assign ng33999 = ( wire32724 ) | ( ng29486  &  wire32720 ) | ( (~ ng29486)  &  wire32722 ) ;
 assign ng29250 = ( wire4335 ) | ( wire4336 ) | ( wire32740 ) | ( wire32741 ) ;
 assign ng33019 = ( wire32745 ) | ( pg35  &  (~ ng2756)  &  ng25317 ) | ( pg35  &  ng2756  &  (~ ng25317) ) ;
 assign ng33595 = ( wire4319 ) | ( wire4320 ) | ( (~ pg35)  &  ng2509 ) ;
 assign ng34022 = ( wire4315 ) | ( wire4316 ) | ( wire32751 ) ;
 assign ng30557 = ( wire4314 ) | ( (~ ng15042)  &  wire32753 ) | ( ng15042  &  wire32754 ) ;
 assign ng33032 = ( (~ pg35)  &  ng3863 ) | ( (~ ng27635)  &  wire32757 ) ;
 assign ng33602 = ( wire4308 ) | ( wire32760 ) ;
 assign ng33612 = ( wire4306 ) | ( (~ ng28471)  &  wire32762 ) | ( (~ ng28471)  &  wire32764 ) ;
 assign ng26906 = ( wire4303 ) | ( (~ ng10632)  &  wire32766 ) | ( ng10632  &  wire32767 ) ;
 assign ng30450 = ( wire4300 ) | ( (~ ng14170)  &  wire32769 ) | ( ng14170  &  wire32770 ) ;
 assign ng30339 = ( wire32775 ) | ( pg35  &  ng24591 ) ;
 assign ng34464 = ( wire32780 ) | ( ng31003  &  (~ ng10831)  &  wire32779 ) ;
 assign ng30428 = ( wire4288 ) | ( (~ ng14133)  &  wire32781 ) | ( ng14133  &  wire32782 ) ;
 assign ng34028 = ( (~ pg35)  &  ng4681 ) | ( ng4681  &  ng31003 ) ;
 assign ng30401 = ( wire4283 ) | ( ng13915  &  wire32784 ) | ( (~ ng13915)  &  wire32785 ) ;
 assign ng33569 = ( wire4278 ) | ( wire4279 ) | ( (~ pg35)  &  ng2047 ) ;
 assign ng30501 = ( pg35  &  (~ ng5869)  &  (~ ng5857)  &  (~ ng28020) ) ;
 assign ng33204 = ( ni30751 ) | ( wire30176 ) | ( wire30177 ) | ( wire30181 ) ;
 assign ng34720 = ( pg35  &  (~ ng79) ) | ( pg35  &  ng550 ) | ( (~ pg35)  &  ng534 ) ;
 assign ng28043 = ( (~ pg35)  &  ng278 ) | ( pg35  &  (~ ng283)  &  ng23204 ) ;
 assign ng26930 = ( wire32798 ) | ( ng17625  &  (~ ng12377)  &  wire32795 ) ;
 assign ng25592 = ( (~ pg35)  &  ng222 ) | ( pg35  &  pg8358  &  ng11737 ) | ( pg35  &  (~ pg8358)  &  (~ ng11737) ) ;
 assign ng33622 = ( wire4253 ) | ( wire4254 ) | ( (~ pg35)  &  ng6044 ) ;
 assign ng26938 = ( wire32808 ) | ( pg35  &  (~ ng4082)  &  ng10808 ) | ( pg35  &  ng4082  &  (~ ng10808) ) ;
 assign ng28058 = ( wire4248 ) | ( (~ ng19140)  &  wire32810 ) | ( ng19140  &  wire32811 ) ;
 assign ng33054 = ( (~ pg35)  &  ng5523 ) | ( ng5523  &  (~ ng5527)  &  (~ ng28010) ) | ( pg35  &  (~ ng5523)  &  ng5527  &  (~ ng28010) ) ;
 assign ng30464 = ( wire4242 ) | ( ng14915  &  wire32817 ) | ( (~ ng14915)  &  wire32818 ) ;
 assign ng34731 = ( ng19422 ) | ( (~ pg35)  &  ng1283 ) | ( pg35  &  ng1287 ) ;
 assign ng33551 = ( wire4233 ) | ( wire4234 ) | ( wire4235 ) | ( wire4236 ) ;
 assign ng33048 = ( (~ pg35)  &  ng5170 ) | ( (~ ng27999)  &  wire32830 ) ;
 assign ng26925 = ( wire4227 ) | ( wire4228 ) | ( wire32834 ) ;
 assign ng30465 = ( wire4226 ) | ( ng14627  &  wire32836 ) | ( (~ ng14627)  &  wire32837 ) ;
 assign ng29274 = ( pg35  &  ng4284  &  (~ ng13539) ) | ( pg35  &  (~ ng4180)  &  (~ ng13539) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng13539 ) ;
 assign ng34002 = ( wire4220 ) | ( wire4221 ) | ( ng30307  &  wire32842 ) ;
 assign ng25649 = ( (~ pg35)  &  ng3050 ) | ( pg35  &  ng3338 ) ;
 assign ng26887 = ( wire32846 ) | ( pg35  &  ng324  &  (~ ng311) ) ;
 assign ng29308 = ( (~ pg35)  &  ng6523 ) | ( pg35  &  ng6527  &  ng23733 ) | ( pg35  &  (~ ng6527)  &  (~ ng23733) ) ;
 assign ng33621 = ( wire4210 ) | ( (~ ng29008)  &  wire32851 ) | ( (~ ng29008)  &  wire32853 ) ;
 assign ng30449 = ( wire4207 ) | ( (~ ng14157)  &  wire32855 ) | ( ng14157  &  wire32856 ) ;
 assign ng31864 = ( wire32861 ) | ( ng23042  &  wire28708  &  wire32860 ) ;
 assign ng32988 = ( wire4199 ) | ( wire32865 ) | ( (~ pg35)  &  ng1624 ) ;
 assign ng30535 = ( wire4197 ) | ( (~ ng15008)  &  wire32866 ) | ( ng15008  &  wire32867 ) ;
 assign ng32993 = ( wire4191 ) | ( wire32873 ) | ( (~ pg35)  &  ng1798 ) ;
 assign ng34019 = ( wire4189 ) | ( wire4190 ) | ( ng29313  &  wire32874 ) ;
 assign ng25663 = ( pg35  &  ng3689 ) | ( (~ pg35)  &  ng3401 ) ;
 assign ng25594 = ( (~ ng11144)  &  wire32878 ) | ( pg35  &  ng278  &  (~ ng11144) ) ;
 assign ng33624 = ( wire4176 ) | ( wire4177 ) | ( (~ pg35)  &  ng6390 ) ;
 assign ng33539 = ( wire4175 ) | ( ng28504  &  wire32884 ) | ( (~ ng28504)  &  wire32885 ) ;
 assign ng30348 = ( wire4172 ) | ( wire32891 ) | ( (~ ng25337)  &  wire32887 ) ;
 assign ng30335 = ( wire4168 ) | ( (~ ng24875)  &  wire32893 ) | ( ng24875  &  wire32894 ) ;
 assign ng24251 = ( (~ pg35)  &  ng1495 ) | ( ng1495  &  (~ ng10939) ) | ( pg35  &  ng1442  &  ng10939 ) ;
 assign ng29239 = ( wire4157 ) | ( wire4158 ) | ( wire32913 ) | ( wire32914 ) ;
 assign ng33584 = ( wire4156 ) | ( ng28942  &  wire32919 ) ;
 assign ng30419 = ( wire4154 ) | ( ng14130  &  wire32921 ) | ( (~ ng14130)  &  wire32922 ) ;
 assign ng28047 = ( (~ pg35)  &  ng645 ) | ( ng645  &  (~ ng20248) ) | ( pg35  &  ng681  &  ng20248 ) ;
 assign ng33027 = ( (~ pg35)  &  ng3512 ) | ( (~ ng27617)  &  wire32927 ) ;
 assign ng29273 = ( wire4144 ) | ( wire4145 ) | ( (~ pg35)  &  ng3831 ) ;
 assign ng25601 = ( (~ pg35)  &  ng182 ) | ( ng182  &  (~ ng11676) ) | ( pg35  &  ng174  &  ng11676 ) ;
 assign ng34442 = ( wire32939 ) | ( pg35  &  ng29503  &  wire32936 ) ;
 assign ng30539 = ( wire4133 ) | ( (~ ng12578)  &  wire32940 ) | ( ng12578  &  wire32941 ) ;
 assign ng33187 = ( wire30033 ) | ( wire30034 ) | ( wire30052 ) | ( wire30053 ) ;
 assign ng26905 = ( wire4127 ) | ( (~ ng10632)  &  wire32943 ) | ( ng10632  &  wire32944 ) ;
 assign ng30459 = ( pg35  &  (~ ng5176)  &  (~ ng5164)  &  (~ ng27999) ) ;
 assign ng30378 = ( wire4124 ) | ( wire32953 ) | ( (~ ng25476)  &  wire32949 ) ;
 assign ng26970 = ( pg35  &  ng4473 ) | ( (~ pg35)  &  ng4459 ) ;
 assign ng33610 = ( wire4118 ) | ( (~ ng28458)  &  wire32955 ) | ( (~ ng28458)  &  wire32957 ) ;
 assign ng31870 = ( wire32961 ) | ( pg35  &  (~ ng1263)  &  (~ ng25895) ) ;
 assign ng34463 = ( wire32966 ) | ( ng31003  &  (~ ng10831)  &  wire32965 ) ;
 assign ng33575 = ( wire4106 ) | ( wire4107 ) | ( wire4108 ) | ( wire4109 ) ;
 assign ng26957 = ( wire32976 ) | ( wire29520  &  wire29521  &  wire32975 ) ;
 assign ng28045 = ( wire4100 ) | ( wire4101 ) | ( (~ pg35)  &  ng568 ) ;
 assign ng33614 = ( wire32985 ) | ( (~ ng28484)  &  ng23342  &  wire32983 ) ;
 assign ng26898 = ( wire4094 ) | ( wire4095 ) | ( (~ pg35)  &  ng843 ) ;
 assign ng28066 = ( wire4068 ) | ( wire4069 ) | ( (~ pg35)  &  ng3614 ) ;
 assign ng24203 = ( (~ pg35)  &  ng429 ) | ( ng429  &  (~ ng8806) ) | ( pg35  &  ng401  &  ng8806 ) ;
 assign ng29224 = ( wire4064 ) | ( ng23978  &  wire33054 ) | ( (~ ng23978)  &  wire33055 ) ;
 assign ng30375 = ( (~ pg35)  &  ng2389 ) | ( pg35  &  ng2393  &  ng25349 ) | ( pg35  &  (~ ng2393)  &  (~ ng25349) ) ;
 assign ng33015 = ( wire4051 ) | ( wire33065 ) | ( (~ pg35)  &  ng2595 ) ;
 assign ng30529 = ( wire4050 ) | ( (~ ng14773)  &  wire33066 ) | ( ng14773  &  wire33067 ) ;
 assign ng33990 = ( wire4045 ) | ( wire4047 ) | ( ng30311  &  wire33070 ) ;
 assign ng25605 = ( wire4044 ) | ( (~ ng11676)  &  wire33072 ) | ( ng11676  &  wire33073 ) ;
 assign ng30406 = ( wire4041 ) | ( ng14069  &  wire33075 ) | ( (~ ng14069)  &  wire33076 ) ;
 assign ng34721 = ( pg35  &  ng222 ) | ( (~ pg35)  &  ng136 ) | ( pg35  &  ng199 ) ;
 assign ng25695 = ( wire4034 ) | ( wire33081 ) ;
 assign ng34808 = ( wire33083 ) | ( pg35  &  ng17694 ) | ( pg35  &  ng17727 ) ;
 assign ng26921 = ( wire33088 ) | ( (~ ng1395)  &  wire33087 ) | ( ng13134  &  wire33087 ) ;
 assign ng34724 = ( wire4025 ) | ( (~ ng33851)  &  wire33090 ) | ( ng33851  &  wire33091 ) ;
 assign ng33021 = ( (~ pg35)  &  ng3155 ) | ( (~ ng3161)  &  ng3155  &  (~ ng27602) ) | ( pg35  &  ng3161  &  (~ ng3155)  &  (~ ng27602) ) ;
 assign ng33557 = ( wire4016 ) | ( wire4017 ) | ( wire4018 ) | ( wire4019 ) ;
 assign ng33563 = ( wire4011 ) | ( wire4012 ) | ( (~ pg35)  &  ng1950 ) ;
 assign ng29225 = ( wire4007 ) | ( (~ ng23324)  &  wire33105 ) | ( (~ ng23324)  &  wire33107 ) ;
 assign ng32984 = ( wire4003 ) | ( wire33111 ) ;
 assign ng30508 = ( wire4001 ) | ( ng14732  &  wire33112 ) | ( (~ ng14732)  &  wire33113 ) ;
 assign ng34444 = ( wire33121 ) | ( pg35  &  ng29503  &  wire33118 ) ;
 assign ng30547 = ( wire33124 ) | ( (~ ng12716)  &  wire33123 ) | ( (~ ng12680)  &  wire33123 ) ;
 assign ng28073 = ( wire33129 ) | ( (~ ng13806)  &  wire33128 ) | ( wire33126  &  wire33128 ) ;
 assign ng25735 = ( wire3988 ) | ( wire33136 ) | ( ng10869  &  wire33131 ) ;
 assign ng30417 = ( wire33139 ) | ( ng11483  &  ng11571  &  wire33138 ) ;
 assign ng33547 = ( wire3979 ) | ( wire3980 ) | ( (~ pg35)  &  ng1682 ) ;
 assign ng33549 = ( wire3975 ) | ( wire3976 ) | ( wire3977 ) | ( wire3978 ) ;
 assign ng25707 = ( wire3974 ) | ( wire33155 ) | ( ng10823  &  wire33150 ) ;
 assign ng33001 = ( wire3967 ) | ( wire33160 ) | ( (~ pg35)  &  ng2066 ) ;
 assign ng31901 = ( wire3961 ) | ( wire3962 ) | ( (~ pg35)  &  ng5041 ) ;
 assign ng33616 = ( (~ pg35)  &  ng4515 ) | ( pg35  &  (~ wire6826)  &  (~ wire6827) ) ;
 assign ng30434 = ( wire3958 ) | ( (~ ng14051)  &  wire33165 ) | ( ng14051  &  wire33166 ) ;
 assign ng30479 = ( wire3955 ) | ( ng14800  &  wire33168 ) | ( (~ ng14800)  &  wire33169 ) ;
 assign ng34258 = ( wire3952 ) | ( (~ ng30583)  &  wire33172 ) | ( (~ ng30583)  &  wire33174 ) ;
 assign ng18597 = ( (~ pg35)  &  ng2975 ) ;
 assign ng30473 = ( wire3946 ) | ( ng14918  &  wire33176 ) | ( (~ ng14918)  &  wire33177 ) ;
 assign ng34735 = ( (~ pg35)  &  ng4297 ) | ( pg35  &  ng4300 ) | ( pg35  &  ng4242 ) ;
 assign ng34007 = ( wire3939 ) | ( wire3940 ) | ( ng30307  &  wire33180 ) ;
 assign ng26963 = ( pg6750  &  pg35 ) | ( (~ pg35)  &  ng4489 ) ;
 assign ng25676 = ( pg35  &  ng3881 ) ;
 assign ng30453 = ( wire3932 ) | ( (~ ng14024)  &  wire33183 ) | ( ng14024  &  wire33184 ) ;
 assign ng24336 = ( wire3926 ) | ( wire3927 ) | ( wire3928 ) | ( wire3929 ) ;
 assign ng32996 = ( wire3922 ) | ( wire33211 ) | ( (~ pg35)  &  ng1894 ) ;
 assign ng30521 = ( wire3921 ) | ( (~ ng14895)  &  wire33212 ) | ( ng14895  &  wire33213 ) ;
 assign ng30510 = ( wire3918 ) | ( ng14810  &  wire33215 ) | ( (~ ng14810)  &  wire33216 ) ;
 assign ng30495 = ( wire3915 ) | ( (~ ng14993)  &  wire33218 ) | ( ng14993  &  wire33219 ) ;
 assign ng34023 = ( wire33227 ) | ( (~ wire6804)  &  (~ wire6805)  &  wire33225 ) ;
 assign ng24209 = ( pg35  &  ng417  &  ng8806 ) | ( pg35  &  ng446  &  (~ ng8806) ) ;
 assign ng33972 = ( wire3905 ) | ( wire3906 ) | ( ng30293  &  wire33230 ) ;
 assign ng33993 = ( wire3902 ) | ( wire3903 ) | ( ng30311  &  wire33233 ) ;
 assign ng30366 = ( (~ pg35)  &  ng2116 ) | ( ng2116  &  (~ ng25389) ) | ( pg35  &  ng2122  &  ng25389 ) ;
 assign ng34014 = ( wire3895 ) | ( wire3897 ) | ( ng30314  &  wire33239 ) ;
 assign ng26940 = ( wire3894 ) | ( (~ pg35)  &  ng4153 ) ;
 assign ng30555 = ( wire3892 ) | ( ng15014  &  wire33241 ) | ( (~ ng15014)  &  wire33242 ) ;
 assign ng30418 = ( wire33246 ) | ( ng11527  &  ng11571  &  wire33245 ) ;
 assign ng33960 = ( wire33250 ) | ( ng28353  &  (~ wire28711)  &  wire33249 ) ;
 assign ng30517 = ( wire3883 ) | ( (~ ng14735)  &  wire33251 ) | ( ng14735  &  wire33252 ) ;
 assign ng30553 = ( wire3880 ) | ( (~ ng14947)  &  wire33254 ) | ( ng14947  &  wire33255 ) ;
 assign ng25629 = ( wire33261 ) | ( ng11130  &  (~ ng11148)  &  wire33259 ) ;
 assign ng30462 = ( wire33264 ) | ( (~ ng12405)  &  wire33263 ) | ( (~ ng12492)  &  wire33263 ) ;
 assign ng33978 = ( wire33270 ) | ( ng29485  &  wire33266 ) | ( (~ ng29485)  &  wire33268 ) ;
 assign ng33589 = ( wire3853 ) | ( wire3854 ) | ( wire3855 ) | ( wire3856 ) ;
 assign ng34726 = ( (~ pg35)  &  ng947 ) | ( pg35  &  (~ ng962) ) | ( pg35  &  ng952 ) ;
 assign ng33006 = ( wire33286 ) | ( wire33287 ) ;
 assign ng30516 = ( wire3845 ) | ( (~ ng15018)  &  wire33288 ) | ( ng15018  &  wire33289 ) ;
 assign ng34603 = ( pg35  &  ng2130 ) ;
 assign ng25618 = ( wire3837 ) | ( wire3838 ) | ( (~ pg35)  &  ng817 ) ;
 assign ng26933 = ( wire33299 ) | ( ng17625  &  (~ ng12377)  &  wire33296 ) ;
 assign ng24346 = ( (~ pg35)  &  ng6035 ) | ( pg35  &  (~ ng6044)  &  (~ ng6035) ) | ( pg35  &  (~ ng6044)  &  ng10185 ) ;
 assign ng32991 = ( wire3828 ) | ( wire33306 ) | ( (~ pg35)  &  ng1768 ) ;
 assign ng30368 = ( wire3827 ) | ( wire33312 ) | ( ng25396  &  wire33308 ) ;
 assign ng24243 = ( pg35  &  pg12919 ) | ( (~ pg35)  &  ng1236 ) ;
 assign ng31896 = ( wire3821 ) | ( wire33316 ) | ( wire33317 ) ;
 assign ng30423 = ( wire3816 ) | ( (~ ng13983)  &  wire33319 ) | ( ng13983  &  wire33320 ) ;
 assign ng25722 = ( (~ pg35)  &  ng5503 ) | ( ng5503  &  ng10838 ) | ( pg35  &  ng5467  &  (~ ng10838) ) ;
 assign ng34454 = ( wire3810 ) | ( ng27020  &  wire33325 ) | ( (~ ng27020)  &  wire33327 ) ;
 assign ng32995 = ( wire3804 ) | ( wire33334 ) | ( (~ pg35)  &  ng1902 ) ;
 assign ng28105 = ( wire3801 ) | ( wire3802 ) | ( (~ pg35)  &  ng6657 ) ;
 assign ng33057 = ( (~ pg35)  &  ng5857 ) | ( ng5857  &  (~ ng5863)  &  (~ ng28020) ) | ( pg35  &  (~ ng5857)  &  ng5863  &  (~ ng28020) ) ;
 assign ng25758 = ( wire33343 ) | ( pg35  &  (~ pg9817)  &  ng6444 ) ;
 assign ng30478 = ( wire3791 ) | ( (~ ng14758)  &  wire33344 ) | ( ng14758  &  wire33345 ) ;
 assign ng29251 = ( wire3786 ) | ( wire3787 ) | ( wire33351 ) ;
 assign ng28082 = ( wire3782 ) | ( wire33354 ) ;
 assign ng24249 = ( wire3780 ) | ( ng10939  &  wire33355 ) | ( (~ ng10939)  &  wire33357 ) ;
 assign ng21896 = ( (~ pg35)  &  ng4245 ) | ( pg35  &  pg8839  &  (~ ng4281) ) | ( pg35  &  (~ pg8839)  &  (~ ng4281) ) ;
 assign ng24270 = ( (~ pg35)  &  ng3343 ) | ( ng3343  &  (~ ng3338) ) | ( ng3343  &  ng8691 ) ;
 assign ng33580 = ( wire3771 ) | ( wire3772 ) | ( (~ pg35)  &  ng2259 ) ;
 assign ng33564 = ( wire3768 ) | ( wire3769 ) | ( (~ pg35)  &  ng1968 ) ;
 assign ng29232 = ( wire3762 ) | ( wire3763 ) | ( wire33370 ) ;
 assign ng34008 = ( wire3760 ) | ( wire3761 ) | ( ng30314  &  wire33373 ) ;
 assign ng33565 = ( wire3755 ) | ( wire3756 ) | ( wire3757 ) | ( wire3758 ) ;
 assign ng24351 = ( (~ pg35)  &  ng6386 ) | ( (~ ng6381)  &  ng6386 ) | ( ng6386  &  ng10207 ) ;
 assign ng30396 = ( wire33384 ) | ( ng11514  &  ng11435  &  wire33383 ) ;
 assign ng33979 = ( wire3746 ) | ( wire3747 ) | ( ng30298  &  wire33385 ) ;
 assign ng30386 = ( (~ pg35)  &  ng2675 ) | ( ng2675  &  (~ ng25439) ) | ( pg35  &  ng2681  &  ng25439 ) ;
 assign ng30376 = ( (~ pg35)  &  ng2407 ) | ( ng2407  &  (~ ng25349) ) | ( pg35  &  ng2413  &  ng25349 ) ;
 assign ng24339 = ( (~ pg35)  &  ng5348 ) | ( ng5348  &  (~ ng5343) ) | ( ng5348  &  ng10124 ) ;
 assign ng30550 = ( wire3736 ) | ( (~ ng14822)  &  wire33392 ) | ( ng14822  &  wire33393 ) ;
 assign ng34608 = ( (~ pg35)  &  ng2697 ) | ( pg35  &  ng2704 ) ;
 assign ng29249 = ( wire3729 ) | ( wire3730 ) | ( wire33399 ) ;
 assign ng33010 = ( wire33407 ) | ( wire33408 ) ;
 assign ng29280 = ( wire3720 ) | ( wire3721 ) | ( wire3722 ) | ( wire3723 ) ;
 assign ng30491 = ( wire3719 ) | ( (~ ng14848)  &  wire33416 ) | ( ng14848  &  wire33417 ) ;
 assign ng29256 = ( wire33421 ) | ( pg35  &  ng2735  &  ng17297 ) | ( pg35  &  (~ ng2735)  &  (~ ng17297) ) ;
 assign ng34461 = ( wire33427 ) | ( ng31003  &  (~ ng10831)  &  wire33426 ) ;
 assign ng29231 = ( wire3704 ) | ( wire3705 ) | ( wire33443 ) | ( wire33444 ) ;
 assign ng34723 = ( (~ pg35)  &  ng542 ) | ( pg35  &  ng301 ) | ( pg35  &  ng534 ) ;
 assign ng24252 = ( wire33450 ) | ( pg35  &  pg7946  &  ng1339 ) ;
 assign ng34252 = ( wire3695 ) | ( wire3696 ) | ( (~ pg35)  &  ng767 ) ;
 assign ng34015 = ( wire3693 ) | ( wire3694 ) | ( ng29313  &  wire33456 ) ;
 assign ng30427 = ( wire3691 ) | ( (~ ng14110)  &  wire33459 ) | ( ng14110  &  wire33460 ) ;
 assign ng33535 = ( wire3688 ) | ( (~ ng28444)  &  wire33463 ) | ( ng28444  &  wire33464 ) ;
 assign ng25621 = ( (~ pg35)  &  ng904 ) | ( pg12919  &  ng904  &  (~ ng921) ) | ( pg35  &  pg12919  &  (~ ng904)  &  ng921 ) ;
 assign ng33028 = ( (~ pg35)  &  ng3518 ) | ( ng3518  &  (~ ng3522)  &  (~ ng27617) ) | ( pg35  &  (~ ng3518)  &  ng3522  &  (~ ng27617) ) ;
 assign ng33543 = ( wire3677 ) | ( wire3678 ) | ( (~ pg35)  &  ng1373 ) ;
 assign ng30489 = ( wire3676 ) | ( (~ ng14761)  &  wire33475 ) | ( ng14761  &  wire33476 ) ;
 assign ng24256 = ( (~ pg35)  &  ng1339 ) | ( pg35  &  ng16272  &  ng8476 ) | ( pg35  &  (~ ng16272)  &  (~ ng8476) ) ;
 assign ng21894 = ( (~ pg35)  &  ng4258 ) | ( (~ ng4264)  &  ng4258 ) | ( pg35  &  ng4264  &  (~ ng4258) ) ;
 assign ng30534 = ( wire3667 ) | ( ng14974  &  wire33485 ) | ( (~ ng14974)  &  wire33486 ) ;
 assign ng34807 = ( wire3658 ) | ( wire3659 ) | ( wire33492 ) ;
 assign ng29258 = ( wire3657 ) | ( wire33497 ) | ( (~ ng23067)  &  wire33494 ) ;
 assign ng30352 = ( wire3653 ) | ( wire33503 ) | ( (~ ng25275)  &  wire33499 ) ;
 assign ng29301 = ( wire3649 ) | ( wire33509 ) | ( (~ ng23699)  &  wire33505 ) ;
 assign ng34452 = ( wire3643 ) | ( wire3644 ) | ( (~ pg35)  &  ng4584 ) ;
 assign ng31869 = ( wire33517 ) | ( pg35  &  (~ ng25911)  &  wire7652 ) ;
 assign ng25599 = ( (~ pg35)  &  ng385 ) | ( pg35  &  pg8719  &  ng385  &  ng376 ) ;
 assign ng33046 = ( wire3635 ) | ( (~ ng27670)  &  wire33519 ) | ( ng27670  &  wire33520 ) ;
 assign ng34031 = ( wire33526 ) | ( ng28336  &  ng13464  &  wire33525 ) ;
 assign ng30490 = ( wire3629 ) | ( ng14804  &  wire33527 ) | ( (~ ng14804)  &  wire33528 ) ;
 assign ng34644 = ( pg35  &  ng5507 ) ;
 assign ng25604 = ( (~ pg35)  &  ng460 ) | ( ng460  &  (~ ng11676) ) | ( pg35  &  ng452  &  ng11676 ) ;
 assign ng34881 = ( wire3618 ) | ( wire3619 ) | ( (~ pg35)  &  ng794 ) ;
 assign ng33966 = ( wire3616 ) | ( wire3617 ) | ( ng30293  &  wire33537 ) ;
 assign ng34460 = ( (~ pg35)  &  ng4639 ) | ( ng4639  &  (~ ng4621)  &  (~ ng31950) ) | ( pg35  &  (~ ng4639)  &  ng4621  &  (~ ng31950) ) ;
 assign ng24235 = ( (~ pg35)  &  ng1152 ) | ( ng1152  &  (~ ng10909) ) | ( pg35  &  ng1099  &  ng10909 ) ;
 assign ng33991 = ( wire3607 ) | ( wire3608 ) | ( ng30311  &  wire33544 ) ;
 assign ng24279 = ( wire3600 ) | ( wire3601 ) | ( (~ pg35)  &  ng4235 ) ;
 assign ng30388 = ( wire33561 ) | ( (~ ng2735)  &  wire33560 ) | ( ng17297  &  wire33560 ) ;
 assign ng33005 = ( wire3594 ) | ( wire33566 ) | ( (~ pg35)  &  ng2223 ) ;
 assign ng33064 = ( (~ pg35)  &  ng6215 ) | ( ng6215  &  (~ ng6219)  &  (~ ng26977) ) | ( pg35  &  (~ ng6215)  &  ng6219  &  (~ ng26977) ) ;
 assign ng33550 = ( wire3584 ) | ( wire3585 ) | ( (~ pg35)  &  ng1710 ) ;
 assign ng30360 = ( (~ pg35)  &  ng1964 ) | ( pg35  &  ng1968  &  ng25341 ) | ( pg35  &  (~ ng1968)  &  (~ ng25341) ) ;
 assign ng34036 = ( (~ pg35)  &  ng4871 ) | ( ng4871  &  ng31009 ) ;
 assign ng24267 = ( wire3578 ) | ( ng8691  &  wire33579  &  wire33580 ) ;
 assign ng29291 = ( pg35  &  ng4284  &  (~ ng14227) ) | ( pg35  &  (~ ng4180)  &  (~ ng14227) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng14227 ) ;
 assign ng33538 = ( wire33592 ) | ( ng27629  &  (~ wire28803)  &  wire33591 ) ;
 assign ng30416 = ( wire33595 ) | ( (~ ng11747)  &  wire33594 ) | ( (~ ng11571)  &  wire33594 ) ;
 assign ng24216 = ( (~ pg35)  &  ng854 ) | ( ng854  &  (~ ng8806) ) | ( pg35  &  ng847  &  ng8806 ) ;
 assign ng24344 = ( wire3565 ) | ( ng10185  &  wire33600  &  wire33601 ) ;
 assign ng33973 = ( wire3562 ) | ( wire3563 ) | ( ng30298  &  wire33609 ) ;
 assign ng30374 = ( wire3560 ) | ( wire33617 ) | ( (~ ng25473)  &  wire33613 ) ;
 assign ng29254 = ( wire3549 ) | ( wire3551 ) | ( wire33632 ) | ( wire33633 ) ;
 assign ng33002 = ( wire33641 ) | ( wire33642 ) ;
 assign ng21893 = ( pg35  &  (~ ng4258) ) ;
 assign ng30466 = ( wire3541 ) | ( (~ ng14656)  &  wire33643 ) | ( ng14656  &  wire33644 ) ;
 assign ng29262 = ( pg35  &  ng4284  &  (~ ng13500) ) | ( pg35  &  (~ ng4180)  &  (~ ng13500) ) | ( pg35  &  (~ ng4284)  &  ng4180  &  ng13500 ) ;
 assign ng30482 = ( wire33650 ) | ( (~ ng12798)  &  wire33649 ) | ( (~ ng12558)  &  wire33649 ) ;
 assign ng28074 = ( wire33654 ) | ( ng13806  &  (~ wire33651)  &  wire33653 ) ;
 assign ng24248 = ( wire3526 ) | ( wire33656 ) | ( wire33657 ) ;
 assign ng33968 = ( wire3521 ) | ( wire3522 ) | ( ng30293  &  wire33660 ) ;
 assign ng25736 = ( (~ pg35)  &  ng5849 ) | ( ng5849  &  ng10869 ) | ( pg35  &  ng5813  &  (~ ng10869) ) ;
 assign ng34733 = ( pg35  &  ng4153 ) | ( pg35  &  ng4172 ) ;
 assign ng29223 = ( wire33668 ) | ( (~ ng482)  &  wire33666 ) | ( (~ ng20000)  &  wire33666 ) ;
 assign ng29263 = ( wire3504 ) | ( wire3505 ) | ( wire3506 ) | ( wire3507 ) ;
 assign ng34609 = ( (~ pg35)  &  ng2890 ) | ( pg35  &  ng2844 ) ;
 assign ng34032 = ( wire33680 ) | ( ng28336  &  ng16173  &  wire33678 ) ;
 assign ng34602 = ( pg35  &  ng1291 ) ;
 assign ng34012 = ( wire3497 ) | ( wire3498 ) | ( ng30314  &  wire33681 ) ;
 assign ng30477 = ( wire3495 ) | ( ng14723  &  wire33684 ) | ( (~ ng14723)  &  wire33685 ) ;
 assign ng30354 = ( wire3492 ) | ( wire33693 ) | ( (~ ng25426)  &  wire33688 ) ;
 assign ng26945 = ( wire33696 ) | ( wire29325  &  wire29326  &  wire33695 ) ;
 assign ng34617 = ( (~ pg35)  &  ng2984 ) | ( pg35  &  ng2907 ) ;
 assign ng24232 = ( wire33699 ) | ( wire33700 ) ;
 assign ng29248 = ( wire3468 ) | ( wire3470 ) | ( wire33715 ) | ( wire33716 ) ;
 assign ng24340 = ( wire3464 ) | ( ng10160  &  wire33720  &  wire33721 ) ;
 assign ng30533 = ( wire3462 ) | ( (~ ng14940)  &  wire33728 ) | ( ng14940  &  wire33729 ) ;
 assign ng33049 = ( (~ pg35)  &  ng5176 ) | ( ng5176  &  (~ ng5180)  &  (~ ng27999) ) | ( pg35  &  (~ ng5176)  &  ng5180  &  (~ ng27999) ) ;
 assign ng31868 = ( wire3456 ) | ( (~ ng25888)  &  wire33735 ) | ( ng25888  &  wire33736 ) ;
 assign ng30513 = ( wire3453 ) | ( (~ ng14933)  &  wire33738 ) | ( ng14933  &  wire33739 ) ;
 assign ng33052 = ( (~ pg35)  &  ng5511 ) | ( ng5511  &  (~ ng5517)  &  (~ ng28010) ) | ( pg35  &  (~ ng5511)  &  ng5517  &  (~ ng28010) ) ;
 assign ng34632 = ( (~ pg35)  &  ng4249 ) | ( pg35  &  ng4245 ) ;
 assign ng33579 = ( wire3443 ) | ( wire3444 ) | ( (~ pg35)  &  ng2241 ) ;
 assign ng32998 = ( wire33751 ) | ( wire33752 ) ;
 assign ng24255 = ( wire33754 ) | ( pg35  &  pg17423  &  pg12923 ) ;
 assign ng30446 = ( wire3435 ) | ( ng14082  &  wire33755 ) | ( (~ ng14082)  &  wire33756 ) ;
 assign ng33974 = ( wire3431 ) | ( wire3432 ) | ( ng30298  &  wire33759 ) ;
 assign ng33026 = ( (~ pg35)  &  ng3506 ) | ( ng3506  &  (~ ng3512)  &  (~ ng27617) ) | ( pg35  &  (~ ng3506)  &  ng3512  &  (~ ng27617) ) ;
 assign ng30384 = ( wire3426 ) | ( wire33770 ) | ( (~ ng25514)  &  wire33765 ) ;
 assign ng34267 = ( wire3422 ) | ( wire33775 ) | ( ng29702  &  wire33771 ) ;
 assign ng34438 = ( wire33779 ) | ( (~ ng31509)  &  wire30328  &  wire33778 ) ;
 assign ng33983 = ( wire3411 ) | ( wire3412 ) | ( ng30304  &  wire33780 ) ;
 assign ng25623 = ( wire3408 ) | ( wire33789 ) | ( (~ ng15737)  &  wire33786 ) ;
 assign ng28046 = ( pg35  &  ng645  &  ng20248 ) | ( pg35  &  ng446  &  (~ ng20248) ) ;
 assign ng24200 = ( wire3402 ) | ( (~ ng8806)  &  wire33794 ) | ( ng8806  &  wire33795 ) ;
 assign ng30333 = ( wire3399 ) | ( ng23042  &  wire33798 ) | ( ng23042  &  wire33800 ) ;
 assign ng33605 = ( wire3393 ) | ( wire3394 ) | ( wire3395 ) | ( wire3396 ) ;
 assign ng33069 = ( (~ pg35)  &  ng6561 ) | ( ng6561  &  (~ ng6565)  &  (~ ng26994) ) | ( pg35  &  (~ ng6561)  &  ng6565  &  (~ ng26994) ) ;
 assign ng30505 = ( wire33814 ) | ( ng12609  &  ng12571  &  wire33813 ) ;
 assign ng34882 = ( wire3382 ) | ( wire3383 ) | ( wire33842 ) ;
 assign ng30393 = ( pg35  &  (~ ng3155)  &  (~ ng3167)  &  (~ ng27602) ) ;
 assign ng30494 = ( wire3376 ) | ( (~ ng14959)  &  wire33846 ) | ( ng14959  &  wire33847 ) ;
 assign ng26971 = ( (~ pg35)  &  ng4512 ) | ( pg35  &  (~ ng4531) ) | ( pg35  &  (~ ng4581) ) ;
 assign ng25613 = ( wire3367 ) | ( wire3368 ) | ( wire3369 ) | ( wire33862 ) ;
 assign ng30425 = ( wire3356 ) | ( (~ ng14048)  &  wire33865 ) | ( ng14048  &  wire33866 ) ;
 assign ng32999 = ( wire3350 ) | ( wire33873 ) | ( (~ pg35)  &  ng2036 ) ;
 assign ng30387 = ( wire3349 ) | ( wire33879 ) | ( (~ ng25439)  &  wire33875 ) ;
 assign ng33554 = ( wire3343 ) | ( wire3344 ) | ( (~ pg35)  &  ng1772 ) ;
 assign ng25668 = ( (~ pg35)  &  ng3484 ) | ( ng3484  &  ng12692 ) | ( pg35  &  ng3490  &  (~ ng12692) ) ;
 assign ng33022 = ( (~ pg35)  &  ng3161 ) | ( (~ ng27602)  &  wire33886 ) ;
 assign ng34001 = ( wire3336 ) | ( wire3337 ) | ( ng30307  &  wire33888 ) ;
 assign ng25684 = ( (~ pg35)  &  ng3849 ) | ( ng3849  &  ng12735 ) | ( pg35  &  ng3813  &  (~ ng12735) ) ;
 assign ng24244 = ( (~ pg35)  &  ng1087 ) | ( ng1087  &  (~ ng1205) ) | ( pg35  &  (~ ng1087)  &  ng1205 ) ;
 assign ng33004 = ( wire3326 ) | ( wire33898 ) | ( (~ pg35)  &  ng2185 ) ;
 assign ng25616 = ( pg35  &  ng11292  &  ng21284  &  ng12332 ) | ( pg35  &  (~ ng11292)  &  (~ ng21284)  &  ng12332 ) | ( pg35  &  (~ ng11292)  &  ng21284  &  (~ ng12332) ) | ( pg35  &  ng11292  &  (~ ng21284)  &  (~ ng12332) ) ;
 assign ng34734 = ( pg35  &  ng4072 ) | ( (~ pg35)  &  ng4172 ) | ( pg35  &  ng4176 ) ;
 assign ng30527 = ( wire3307 ) | ( ng15021  &  wire33902 ) | ( (~ ng15021)  &  wire33903 ) ;
 assign ng31897 = ( wire3304 ) | ( wire33908 ) | ( wire33909 ) ;
 assign ng30389 = ( wire3298 ) | ( wire31317 ) | ( wire31318 ) | ( wire31319 ) ;
 assign ng24354 = ( (~ pg35)  &  ng6727 ) | ( pg35  &  (~ ng6736)  &  (~ ng6727) ) | ( pg35  &  (~ ng6736)  &  ng10224 ) ;
 assign ng30432 = ( wire3295 ) | ( ng13986  &  wire33912 ) | ( (~ ng13986)  &  wire33913 ) ;
 assign ng31867 = ( wire33918 ) | ( ng24875  &  (~ wire28810)  &  wire33917 ) ;
 assign ng30496 = ( wire3289 ) | ( ng14691  &  wire33919 ) | ( (~ ng14691)  &  wire33920 ) ;
 assign ng34646 = ( pg35  &  ng6199 ) ;
 assign ng33571 = ( wire3284 ) | ( wire3285 ) | ( (~ pg35)  &  ng2084 ) ;
 assign ng25743 = ( pg35  &  ng6381 ) | ( (~ pg35)  &  ng6098 ) ;
 assign ng30439 = ( wire33926 ) | ( (~ ng11626)  &  wire33925 ) | ( (~ ng11584)  &  wire33925 ) ;
 assign ng34802 = ( wire3276 ) | ( wire3278 ) | ( wire33927 ) ;
 assign ng29252 = ( wire3271 ) | ( wire3272 ) | ( wire33943 ) | ( wire33944 ) ;
 assign ng24275 = ( wire33949  &  wire33950 ) | ( wire33954  &  wire33955 ) ;
 assign ng33585 = ( wire3257 ) | ( wire3258 ) | ( (~ pg35)  &  ng2338 ) ;
 assign ng30545 = ( wire33962 ) | ( (~ ng10491)  &  wire33961 ) | ( (~ ng12716)  &  wire33961 ) ;
 assign ng30554 = ( wire3253 ) | ( (~ ng14981)  &  wire33963 ) | ( ng14981  &  wire33964 ) ;
 assign ng33043 = ( wire33970 ) | ( wire33971 ) ;
 assign ng24259 = ( pg35  &  pg12923 ) | ( (~ pg35)  &  ng1579 ) ;
 assign ng33965 = ( wire33975 ) | ( (~ ng28504)  &  wire28813  &  wire33974 ) ;
 assign ng25728 = ( pg35  &  ng5881 ) ;
 assign ng30541 = ( wire3237 ) | ( ng14902  &  wire33976 ) | ( (~ ng14902)  &  wire33977 ) ;
 assign ng30447 = ( wire3234 ) | ( (~ ng14116)  &  wire33979 ) | ( ng14116  &  wire33980 ) ;
 assign ng31872 = ( wire3229 ) | ( wire3230 ) | ( (~ pg35)  &  ng2741 ) ;
 assign ng30372 = ( wire3228 ) | ( wire33993 ) | ( (~ ng25309)  &  wire33988 ) ;
 assign ng24274 = ( (~ pg35)  &  ng3694 ) | ( (~ ng3689)  &  ng3694 ) | ( ng3694  &  ng8728 ) ;
 assign ng26881 = ( pg6744  &  pg35 ) | ( (~ pg35)  &  ng305 ) ;
 assign ng25633 = ( wire33996 ) | ( pg35  &  (~ ng13242)  &  wire5491 ) ;
 assign ng34645 = ( pg35  &  ng5853 ) ;
 assign ng30498 = ( wire3215 ) | ( (~ ng14764)  &  wire33997 ) | ( ng14764  &  wire33998 ) ;
 assign ng30519 = ( wire3212 ) | ( (~ ng14813)  &  wire34000 ) | ( ng14813  &  wire34001 ) ;
 assign ng29287 = ( wire3209 ) | ( wire34007 ) | ( (~ ng23630)  &  wire34004 ) ;
 assign ng33995 = ( wire3203 ) | ( wire3205 ) | ( ng30300  &  wire34010 ) ;
 assign ng20841 = ( pg35  &  ng5138 ) | ( pg35  &  ng5152 ) ;
 assign ng21193 = ( pg35  &  ng6191 ) | ( pg35  &  ng6177 ) ;
 assign ng20982 = ( pg35  &  ng5485 ) | ( pg35  &  ng5499 ) ;
 assign ni24685 = ( (~ ng21193)  &  (~ ng20982)  &  (~ ng21127)  &  (~ ng21256) ) ;
 assign ng19968 = ( pg35  &  ng3480 ) | ( pg35  &  ng3494 ) ;
 assign ng20014 = ( pg35  &  ng3845 ) | ( pg35  &  ng3831 ) ;
 assign ng19919 = ( pg35  &  ng3143 ) | ( pg35  &  ng3129 ) ;
 assign ng21127 = ( pg35  &  ng5831 ) | ( pg35  &  ng5845 ) ;
 assign ng21256 = ( pg35  &  ng6537 ) | ( pg35  &  ng6523 ) ;
 assign ng19422 = ( pg35  &  (~ ng1536) ) | ( pg35  &  (~ ng1312)  &  (~ ng1351) ) ;
 assign ng19402 = ( pg35  &  (~ ng1193) ) | ( pg35  &  (~ ng969)  &  (~ ng1008) ) ;
 assign ng19984 = ( pg35  &  ng3817 ) ;
 assign ng26365 = ( pg35  &  ng4427 ) | ( pg35  &  ng4420 ) ;
 assign ng17657 = ( wire31890 ) | ( wire31891 ) | ( wire31892 ) | ( wire31893 ) ;
 assign ng17700 = ( wire31896 ) | ( wire31897 ) | ( wire31898 ) | ( wire31899 ) ;
 assign ni31106 = ( (~ ng30735)  &  (~ wire29984)  &  (~ wire29985)  &  wire34142 ) ;
 assign ng30937 = ( pg54  &  (~ pg53)  &  ng17653  &  wire29926 ) ;
 assign ng31021 = ( wire29948 ) | ( wire29949 ) | ( wire29950 ) ;
 assign ng31376 = ( wire29985 ) | ( ng27511  &  ng17613 ) | ( ng27511  &  ng17747 ) ;
 assign ng30673 = ( (~ ng31)  &  ng28  &  ng13156  &  wire30042 ) ;
 assign ng30614 = ( (~ ng31)  &  (~ ng28)  &  ng13156  &  wire30045 ) ;
 assign ni31271 = ( (~ ng30735)  &  (~ wire29984)  &  (~ wire29985)  &  wire34136 ) ;
 assign ng30735 = ( (~ ng31)  &  ng28  &  ng13156  &  wire30000 ) ;
 assign ng28180 = ( pg53 ) | ( pg54  &  (~ pg53)  &  wire29926 ) ;
 assign ni31191 = ( ng30735  &  (~ wire29984)  &  (~ wire29985)  &  wire34130 ) ;
 assign ni31121 = ( (~ ng30735)  &  (~ wire29984)  &  (~ wire29985)  &  wire34154 ) ;
 assign ni31141 = ( (~ ng30735)  &  wire29984  &  wire34124 ) | ( (~ ng30735)  &  wire29985  &  wire34124 ) ;
 assign ni30330 = ( ng30735 ) | ( wire29984 ) | ( wire29985 ) | ( wire34118 ) ;
 assign ni31221 = ( (~ wire29984)  &  (~ wire29985)  &  wire34149 ) ;
 assign ng31327 = ( (~ ng31)  &  ng28  &  ng13156  &  wire29997 ) ;
 assign ng17694 = ( wire30696 ) | ( wire30697 ) | ( wire30698 ) | ( wire30699 ) ;
 assign ng17727 = ( wire30702 ) | ( wire30703 ) | ( wire30704 ) | ( wire30705 ) ;
 assign ng31566 = ( (~ ng31)  &  (~ ng28)  &  ng13156  &  wire29962 ) ;
 assign ng31710 = ( ng31  &  (~ ng28)  &  ng13156  &  wire29966 ) ;
 assign ng34237 = ( wire3165 ) | ( wire3166 ) | ( wire34198 ) | ( wire34199 ) ;
 assign ng33496 = ( (~ ng30614)  &  (~ ng31070)  &  wire34201  &  wire34206 ) ;
 assign ni31171 = ( ng31566  &  (~ wire29984)  &  (~ wire29985)  &  wire34239 ) ;
 assign ng31070 = ( ng30937 ) | ( wire29948 ) | ( wire29949 ) | ( wire29950 ) ;
 assign ni31843 = ( wire3155 ) | ( wire3156 ) | ( wire3157 ) | ( wire3158 ) ;
 assign ng34235 = ( ni31843 ) | ( wire3151 ) | ( wire3152 ) | ( wire34248 ) ;
 assign ng25590 = () ;
 assign ng26977 = ( ng43  &  ng29503  &  ng24688  &  wire28470 ) ;
 assign ng18935 = ( ng4322  &  ng4311  &  (~ ng10511)  &  (~ ng8347) ) ;
 assign ng27903 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28503) ) ;
 assign ng22472 = ( wire7725 ) | ( ng14367  &  wire28488 ) ;
 assign ng26390 = ( pg35  &  ng4423 ) ;
 assign ng24591 = ( (~ ng1193)  &  wire7709 ) | ( ng10666  &  wire7709 ) | ( (~ ng1193)  &  wire28519 ) | ( ng10666  &  wire28519 ) ;
 assign ng13977 = ( (~ ng3171) ) | ( ng3179 ) | ( (~ ng3161) ) | ( ng3155 ) ;
 assign ng29503 = ( pg134  &  (~ pg113) ) | ( pg99  &  (~ pg113)  &  ng37 ) ;
 assign ng29676 = ( ng11834  &  ng11283 ) | ( ng24374  &  (~ wire28575) ) ;
 assign ng30590 = ( (~ wire1421)  &  (~ ng4818)  &  ng71  &  ng24374 ) ;
 assign ng8806 = ( (~ ng385) ) | ( (~ ng358) ) | ( (~ ng376) ) | ( ng385  &  ng358  &  (~ ng370)  &  ng376 ) ;
 assign ng10632 = ( (~ ng896)  &  (~ ng862)  &  ng890 ) ;
 assign ng23590 = ( (~ ng11111) ) | ( (~ wire7624)  &  (~ wire7625)  &  (~ wire28651) ) ;
 assign ng27635 = ( ng43  &  ng29503  &  ng24688  &  wire28661 ) ;
 assign ng28761 = ( ng112  &  ng29503  &  ng26314  &  wire28687 ) ;
 assign ng27602 = ( ng43  &  ng29503  &  ng24688  &  wire28694 ) ;
 assign ng11676 = ( (~ ng385) ) | ( (~ ng358) ) | ( ng370 ) | ( (~ ng376) ) ;
 assign ng31134 = ( ng153  &  ng157  &  ng23042  &  ng28353 ) ;
 assign ng23042 = ( (~ wire28543)  &  (~ wire28544)  &  wire28706 ) | ( (~ wire28543)  &  (~ wire28544)  &  wire28707 ) ;
 assign ng25917 = ( ng7601 ) | ( (~ ng1361)  &  (~ ng15748) ) | ( (~ ng1345)  &  (~ ng15748) ) ;
 assign ng14868 = ( (~ ng6573) ) | ( ng6555 ) | ( (~ ng6549) ) | ( (~ ng6565) ) ;
 assign ng10160 = ( (~ pg14694) ) | ( (~ pg17580) ) | ( (~ pg17711) ) | ( (~ pg12300) ) ;
 assign ng23666 = ( (~ ng11139) ) | ( (~ wire7351)  &  (~ wire7352)  &  (~ wire28734) ) ;
 assign ng10939 = ( (~ pg13272) ) | ( ng1514 ) | ( ng1526 ) ;
 assign ng13378 = ( ng1312  &  ng1536  &  (~ ng1319) ) | ( ng1351  &  ng1536  &  (~ ng1319) ) ;
 assign ng13385 = ( ng305  &  ng324 ) | ( (~ ng324)  &  ng311 ) ;
 assign ng11607 = ( ng385  &  ng358  &  (~ ng376) ) ;
 assign ng30304 = ( ng24457 ) | ( (~ ng4180)  &  wire7269 ) | ( ng1242  &  (~ ng24457)  &  (~ wire7269) ) ;
 assign ng25385 = ( wire28836 ) | ( (~ ng14367)  &  (~ wire7257) ) | ( (~ wire7257)  &  (~ wire28834) ) ;
 assign ng23699 = ( (~ ng11160) ) | ( (~ wire7248)  &  (~ wire7249)  &  (~ wire28843) ) ;
 assign ng30300 = ( ng24447 ) | ( (~ ng4180)  &  wire7306 ) | ( ng1585  &  (~ ng24447)  &  (~ wire7306) ) ;
 assign ng22369 = ( wire7257 ) | ( ng14367  &  wire28834 ) ;
 assign ng27775 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng12377) ) | ( (~ ng25357) ) ;
 assign ng15036 = ( (~ ng6209) ) | ( (~ ng6227) ) | ( (~ ng6203) ) | ( ng6219 ) ;
 assign ng12692 = ( ng3530  &  ng3518  &  ng3522 ) ;
 assign ng20000 = ( ng528  &  ng11607  &  ng12812 ) | ( ng11607  &  ng11185  &  ng12812 ) ;
 assign ng25300 = ( wire28887 ) | ( (~ ng14367)  &  (~ wire7257) ) | ( (~ wire7257)  &  (~ wire28834) ) ;
 assign ng12371 = ( ng1783  &  (~ ng1760) ) ;
 assign ng24609 = ( (~ ng1536)  &  wire7193 ) | ( ng10699  &  wire7193 ) | ( (~ ng1536)  &  wire28903 ) | ( ng10699  &  wire28903 ) ;
 assign ng14058 = ( ng3873 ) | ( (~ ng3881) ) | ( (~ ng3869) ) ;
 assign ng14885 = ( (~ ng5535) ) | ( ng5511 ) | ( (~ ng5527) ) | ( (~ ng5517) ) ;
 assign ng20887 = ( wire7137 ) | ( wire7138 ) | ( wire28996 ) ;
 assign ng12735 = ( ng3873  &  ng3881  &  ng3869 ) ;
 assign ng30311 = ( ng24468 ) | ( (~ ng4180)  &  wire7126 ) | ( (~ ng1242)  &  (~ ng24468)  &  (~ wire7126) ) ;
 assign ng17625 = ( ng2756  &  (~ ng2735) ) | ( ng2756  &  (~ ng2741) ) | ( (~ ng2756)  &  ng2748 ) | ( (~ ng2735)  &  ng2748 ) | ( (~ ng2741)  &  ng2748 ) | ( ng2756  &  (~ ng2748) ) ;
 assign ng12377 = ( (~ ng2756)  &  ng2741  &  (~ ng2748) ) ;
 assign ng31003 = ( (~ ng63) ) | ( (~ ng29503) ) | ( ng24380 ) | ( (~ wire28640) ) ;
 assign ng28336 = ( (~ ng63) ) | ( (~ ng29503) ) | ( ng24380 ) | ( (~ wire28640) ) ;
 assign ng16173 = ( (~ ng4785) ) | ( (~ ng4793) ) | ( (~ ng4776) ) | ( (~ ng10831) ) ;
 assign ng28010 = ( ng43  &  ng29503  &  ng24688  &  wire29495 ) ;
 assign ng13307 = ( (~ pg13259) ) | ( (~ ng1171) ) | ( (~ ng1183) ) ;
 assign ng15039 = ( ng6573 ) | ( ng6555 ) | ( (~ ng6549) ) | ( ng6565 ) ;
 assign ng14683 = ( (~ ng5188) ) | ( ng5170 ) | ( (~ ng5164) ) | ( (~ ng5180) ) ;
 assign ng25371 = ( ng5041  &  ng5046  &  wire29549 ) ;
 assign ng14858 = ( (~ ng5869) ) | ( (~ ng5881) ) | ( ng5873 ) ;
 assign ng11626 = ( (~ ng3857)  &  (~ ng3863)  &  (~ ng3869) ) ;
 assign ng11537 = ( (~ ng3873)  &  ng3881 ) ;
 assign ng7142 = ( (~ ng6573)  &  (~ ng6565) ) ;
 assign ng14905 = ( ng6573 ) | ( (~ ng6555) ) | ( ng6549 ) | ( ng6565 ) ;
 assign ng10925 = ( (~ ng947)  &  ng956 ) ;
 assign ng24468 = ( wire7608 ) | ( wire7609 ) | ( (~ ng947)  &  ng956 ) ;
 assign ng26759 = ( ng10925 ) | ( wire7126 ) | ( wire7608 ) | ( wire7609 ) ;
 assign ng34162 = ( (~ ng32212) ) | ( wire28816 ) | ( (~ wire29718) ) | ( wire29789 ) ;
 assign ng10312 = ( (~ ng5881)  &  (~ ng5873) ) ;
 assign ng12609 = ( (~ ng5869)  &  (~ ng5857)  &  (~ ng5863) ) ;
 assign ng12515 = ( ng5881  &  (~ ng5873) ) ;
 assign ng8958 = ( (~ ng3873)  &  (~ ng3881) ) ;
 assign ng11534 = ( ng3873 ) | ( ng3881 ) | ( (~ ng3869) ) ;
 assign ng10715 = ( ng1514  &  ng1526 ) ;
 assign ng13315 = ( (~ pg13272) ) | ( (~ ng1514) ) | ( (~ ng1526) ) ;
 assign ng12824 = ( (~ ng5881)  &  ng5873 ) ;
 assign ng14697 = ( ng5881 ) | ( (~ ng5873) ) | ( (~ ng5857) ) | ( ng5863 ) ;
 assign ng28140 = ( wire29507 ) | ( wire29508 ) ;
 assign ng27972 = ( pg73 ) | ( pg72 ) ;
 assign ng22432 = ( wire7030 ) | ( ng14367  &  wire29111 ) ;
 assign ng12437 = ( ng2342  &  (~ ng2319) ) ;
 assign ng25473 = ( (~ ng12437) ) | ( (~ ng14367)  &  (~ wire7030) ) | ( (~ wire7030)  &  (~ wire29111) ) ;
 assign ng10491 = ( (~ ng6573)  &  ng6565 ) ;
 assign ng14947 = ( ng6573 ) | ( (~ ng6555) ) | ( ng6549 ) | ( (~ ng6565) ) ;
 assign ng17766 = ( ng31  &  (~ ng28)  &  ng13156  &  wire29982 ) ;
 assign ng17613 = ( (~ ng31)  &  (~ ng28)  &  ng13156  &  wire29980 ) ;
 assign ng17747 = ( (~ ng31)  &  (~ ng28)  &  ng13156  &  wire29978 ) ;
 assign ng17724 = ( ng31  &  ng28  &  ng13156  &  wire29976 ) ;
 assign ng17690 = ( (~ ng31)  &  ng28  &  ng13156  &  wire29974 ) ;
 assign ng24374 = ( pg134 ) | ( pg99  &  ng37 ) ;
 assign ng20875 = ( wire7351 ) | ( wire7352 ) | ( wire28734 ) ;
 assign ng23932 = ( (~ ng6049) ) | ( (~ wire7351)  &  (~ wire7352)  &  (~ wire28734) ) ;
 assign ng31509 = ( (~ ng27629) ) | ( wire28803 ) | ( (~ wire28804) ) | ( wire30327 ) ;
 assign ng12571 = ( ng5881  &  ng5873 ) ;
 assign ng14735 = ( (~ ng5881) ) | ( (~ ng5873) ) | ( (~ ng5857) ) | ( (~ ng5863) ) ;
 assign ng9694 = ( (~ ng1936)  &  (~ ng1862) ) ;
 assign ng26314 = ( pg73  &  pg72  &  ng482  &  ng490 ) | ( pg73  &  (~ pg72)  &  (~ ng482)  &  ng490 ) | ( (~ pg73)  &  pg72  &  ng482  &  (~ ng490) ) | ( (~ pg73)  &  (~ pg72)  &  (~ ng482)  &  (~ ng490) ) ;
 assign ng27494 = ( (~ ng504)  &  ng518  &  ng528  &  ng26314 ) ;
 assign ni18740 = ( (~ ng31)  &  (~ ng28)  &  ng13156 ) ;
 assign ng10967 = ( ng1448  &  (~ ng1291) ) ;
 assign ng12512 = ( (~ ng5869) ) | ( ng5881 ) | ( ng5873 ) ;
 assign ng12632 = ( ng6573  &  (~ ng6565) ) ;
 assign ng14950 = ( (~ ng6573) ) | ( (~ ng6561) ) | ( ng6565 ) ;
 assign ng26770 = ( ng10999 ) | ( wire6912 ) | ( wire7308 ) | ( wire7309 ) ;
 assign ng17424 = ( wire29269 ) | ( pg17423  &  (~ ng10715) ) | ( pg17423  &  (~ ng7675) ) ;
 assign ng11012 = ( ng4849  &  ng4843  &  ng4878 ) ;
 assign ng11797 = ( ng4785  &  ng4709 ) ;
 assign ng11261 = ( (~ ng4801)  &  ng4793  &  ng4776 ) ;
 assign ng10831 = ( ng4653  &  ng4669  &  ng4688  &  ng4659 ) ;
 assign ng29737 = ( ng11804  &  ng11283 ) | ( ng24374  &  (~ wire28575) ) ;
 assign ng11194 = ( (~ ng3352)  &  (~ ng3288) ) ;
 assign ng11350 = ( (~ pg11349)  &  ng3338 ) | ( pg11349  &  (~ ng3338) ) ;
 assign ng13700 = ( ng3352  &  (~ ng3288) ) ;
 assign ng13765 = ( ng3352  &  ng3288 ) ;
 assign ng24457 = ( wire7608 ) | ( wire7609 ) | ( (~ ng947)  &  ng1129 ) ;
 assign ng26725 = ( ng10902 ) | ( wire7269 ) | ( wire7608 ) | ( wire7609 ) ;
 assign ng12026 = ( (~ ng2724)  &  (~ ng2729) ) ;
 assign ng14367 = ( (~ ng2756)  &  ng2735  &  (~ ng2741)  &  (~ ng2748) ) ;
 assign ng11960 = ( ng2495  &  (~ ng2465) ) ;
 assign ng11804 = ( (~ ng4975)  &  ng4899 ) ;
 assign ng11173 = ( ng4991 ) | ( (~ ng4966) ) | ( ng4983 ) ;
 assign ng21024 = ( wire6966 ) | ( wire6967 ) | ( wire29216 ) ;
 assign ng11389 = ( (~ pg11388)  &  ng3689 ) | ( pg11388  &  (~ ng3689) ) ;
 assign ng13806 = ( (~ ng4087)  &  (~ ng4098)  &  (~ ng4093)  &  (~ ng4076) ) ;
 assign ng29672 = ( ng11261  &  ng8933 ) | ( ng24374  &  (~ wire29730) ) ;
 assign ng14708 = ( pg9048  &  ng74 ) | ( (~ pg12368)  &  ng74 ) ;
 assign ng17653 = ( (~ ng31)  &  (~ ng28)  &  ng13156  &  wire29959 ) ;
 assign ng24688 = ( pg73  &  pg72  &  ng4104  &  ng4108 ) | ( (~ pg73)  &  pg72  &  (~ ng4104)  &  ng4108 ) | ( pg73  &  (~ pg72)  &  ng4104  &  (~ ng4108) ) | ( (~ pg73)  &  (~ pg72)  &  (~ ng4104)  &  (~ ng4108) ) ;
 assign ng30583 = ( pg73  &  ng65 ) | ( pg72  &  ng65 ) | ( ng65  &  ng29503 ) ;
 assign ng11780 = ( ng4975  &  (~ ng4899) ) ;
 assign ng22342 = ( wire7041 ) | ( ng14367  &  wire29097 ) ;
 assign ng25275 = ( wire29099 ) | ( (~ ng14367)  &  (~ wire7041) ) | ( (~ wire7041)  &  (~ wire29097) ) ;
 assign ng10511 = ( ng4639 ) | ( (~ ng4628) ) | ( (~ ng4621) ) ;
 assign ng10902 = ( (~ ng947)  &  ng1129 ) ;
 assign ng16244 = ( (~ ng31)  &  (~ ng28)  &  ng14988  &  wire29946 ) ;
 assign ng16194 = ( (~ ng31)  &  ng28  &  ng13156  &  wire29941 ) ;
 assign ng17725 = ( (~ ng31)  &  ng28  &  ng13156  &  wire29939 ) ;
 assign ng16283 = ( (~ ng31)  &  ng28  &  ng14988  &  wire29936 ) ;
 assign ng16205 = ( ng31  &  ng28  &  ng13156  &  wire29934 ) ;
 assign ng12333 = ( (~ ng1624)  &  ng1648 ) ;
 assign ng25776 = ( pg72  &  ng4322  &  wire29233 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233 ) ;
 assign ng31009 = ( (~ ng63) ) | ( (~ ng29503) ) | ( ng24380 ) | ( (~ wire29233) ) ;
 assign ng22457 = ( wire6319 ) | ( ng14367  &  wire30342 ) ;
 assign ng25470 = ( wire30343 ) | ( (~ ng14367)  &  (~ wire6319) ) | ( (~ wire6319)  &  (~ wire30342) ) ;
 assign ng13273 = ( (~ pg13272) ) | ( ng1514 ) | ( (~ ng1526) ) ;
 assign ng10961 = ( ng1495 ) | ( (~ ng1442) ) ;
 assign ng16539 = ( (~ ng31)  &  (~ ng28)  &  ng14988  &  wire29944 ) ;
 assign ng16486 = ( (~ ng31)  &  ng28  &  ng14988  &  wire29930 ) ;
 assign ng25317 = ( ng2735  &  ng2741  &  ng2748  &  (~ ng17297) ) ;
 assign ng11473 = ( ng3171  &  ng3179 ) ;
 assign ng13892 = ( (~ ng3171) ) | ( (~ ng3179) ) | ( (~ ng3161) ) | ( (~ ng3155) ) ;
 assign ng10671 = ( ng1514  &  (~ ng1526) ) ;
 assign ng13861 = ( (~ pg13272) ) | ( (~ ng1514) ) | ( ng1526 ) ;
 assign ng12581 = ( ng6227  &  (~ ng6219) ) ;
 assign ng11185 = ( ng482  &  (~ ng528)  &  ng490 ) ;
 assign ng14822 = ( (~ ng6573) ) | ( ng6555 ) | ( (~ ng6549) ) | ( ng6565 ) ;
 assign ng25382 = ( (~ ng12333) ) | ( (~ ng14367)  &  (~ wire7041) ) | ( (~ wire7041)  &  (~ wire29097) ) ;
 assign ng14291 = ( ng2715  &  ng2724  &  ng2719 ) ;
 assign ng17297 = ( (~ ng2715) ) | ( (~ ng2724) ) | ( (~ ng2729) ) | ( (~ ng2719) ) ;
 assign ng8864 = ( (~ ng3171)  &  (~ ng3179) ) ;
 assign ng11514 = ( (~ ng3161)  &  (~ ng3155)  &  (~ ng3167) ) ;
 assign ng11155 = ( ng4801 ) | ( ng4793 ) | ( (~ ng4776) ) ;
 assign ng11755 = ( ng4785  &  (~ ng4709) ) ;
 assign ng20739 = ( wire6832 ) | ( wire6833 ) | ( wire29346 ) ;
 assign ng10808 = ( ng4141  &  ng4064  &  ng4057 ) ;
 assign ng13217 = ( (~ ng4141) ) | ( (~ ng4064) ) | ( (~ ng4057) ) | ( (~ ng4082) ) ;
 assign ng24875 = ( (~ wire7284)  &  wire28543  &  wire28809 ) | ( (~ wire7284)  &  wire28544  &  wire28809 ) ;
 assign ng12716 = ( (~ ng6561)  &  (~ ng6555)  &  (~ ng6549) ) ;
 assign ng8906 = ( (~ ng3530)  &  (~ ng3522) ) ;
 assign ng11480 = ( ng3530 ) | ( (~ ng3518) ) | ( ng3522 ) ;
 assign ng15737 = ( ng969 ) | ( wire28609 ) | ( (~ ng7598)  &  wire28607 ) ;
 assign ng25911 = ( ng7567 ) | ( (~ ng1018)  &  (~ ng15737) ) | ( (~ ng1002)  &  (~ ng15737) ) ;
 assign ng34703 = ( (~ ng34162)  &  wire31938  &  (~ wire31939)  &  wire31940 ) ;
 assign ng8967 = ( (~ ng4264) ) | ( (~ ng4258) ) ;
 assign ng14996 = ( ng5881 ) | ( ng5873 ) | ( (~ ng5857) ) | ( ng5863 ) ;
 assign ng29186 = ( (~ ng4507) ) | ( (~ pg99)  &  (~ pg134) ) | ( (~ pg134)  &  (~ ng37) ) ;
 assign ng22417 = ( wire6655 ) | ( ng14367  &  wire29571 ) ;
 assign ng10421 = ( (~ ng6227)  &  ng6219 ) ;
 assign ng14741 = ( ng6209 ) | ( ng6227 ) | ( (~ ng6203) ) | ( (~ ng6219) ) ;
 assign ng12911 = ( (~ ng4639) ) | ( (~ ng4628) ) | ( (~ ng4621) ) ;
 assign ng13242 = ( (~ ng1322)  &  (~ ng1333) ) | ( ng1322  &  ng1339 ) | ( (~ ng1322)  &  (~ ng1339) ) ;
 assign ng27440 = ( ng504  &  ng518  &  (~ ng528)  &  ng26314 ) ;
 assign ng17401 = ( wire28827 ) | ( pg17400  &  (~ ng7661) ) | ( pg17400  &  (~ ng10695) ) ;
 assign ng10341 = ( (~ ng6227)  &  (~ ng6219) ) ;
 assign ng14861 = ( (~ ng6209) ) | ( ng6227 ) | ( ng6203 ) | ( ng6219 ) ;
 assign ni18785 = ( ng31  &  (~ ng28)  &  ng13156 ) ;
 assign ng12289 = ( ng2756 ) | ( ng2741 ) | ( ng2748 ) ;
 assign ng21277 = ( (~ ng2724)  &  (~ ng2729)  &  (~ ng2735)  &  (~ ng12289) ) ;
 assign ng10929 = ( ng1152 ) | ( (~ ng1099) ) ;
 assign ng14015 = ( ng3530 ) | ( ng3506 ) | ( (~ ng3522) ) | ( (~ ng3512) ) ;
 assign ng14271 = ( (~ ng6215)  &  ng6195 ) | ( ng6195  &  (~ ng6227) ) | ( ng6195  &  (~ ng6219) ) ;
 assign ng22992 = ( pg35  &  pg12919 ) ;
 assign ng28903 = ( (~ ng2197) ) | ( ng2153 ) | ( (~ ng26703)  &  (~ ng17321) ) ;
 assign ng14021 = ( ng3873 ) | ( ng3857 ) | ( ng3881 ) | ( (~ ng3863) ) ;
 assign ng12641 = ( ng3171  &  ng3179  &  ng3167 ) ;
 assign ng12915 = ( (~ ng6573) ) | ( (~ ng6555) ) | ( (~ ng6549) ) | ( ng6565 ) ;
 assign ng28880 = ( ng112  &  ng29503  &  ng26314  &  wire29061 ) ;
 assign ng23733 = ( (~ ng11178) ) | ( (~ wire7046)  &  (~ wire7047)  &  (~ wire29091) ) ;
 assign ng29488 = ( ng24457 ) | ( (~ ng4180)  &  wire7269 ) | ( ng1246  &  (~ ng24457)  &  (~ wire7269) ) ;
 assign ng25349 = ( wire29113 ) | ( (~ ng14367)  &  (~ wire7030) ) | ( (~ wire7030)  &  (~ wire29111) ) ;
 assign ng10207 = ( (~ pg17760) ) | ( (~ pg14779) ) | ( (~ pg17649) ) | ( (~ pg12422) ) ;
 assign ng11915 = ( (~ ng1772)  &  ng1802 ) ;
 assign ng27999 = ( ng43  &  ng29503  &  ng24688  &  wire29192 ) ;
 assign ng14306 = ( ng6541  &  (~ ng6573) ) | ( ng6541  &  (~ ng6561) ) | ( ng6541  &  (~ ng6565) ) ;
 assign ng8417 = ( pg13259 ) | ( pg8416 ) | ( wire29209 ) ;
 assign ng16246 = ( (~ ng979)  &  ng1236  &  (~ ng13211)  &  (~ wire29210) ) | ( ng979  &  (~ ng1236)  &  (~ ng13211)  &  (~ wire29210) ) ;
 assign ng23112 = ( (~ ng10733) ) | ( (~ wire6966)  &  (~ wire6967)  &  (~ wire29216) ) ;
 assign ng14782 = ( ng6573 ) | ( ng6555 ) | ( (~ ng6549) ) | ( (~ ng6565) ) ;
 assign ng23280 = ( pg64  &  pg35 ) ;
 assign ng29501 = ( ng24478 ) | ( (~ ng4180)  &  wire7065 ) | ( (~ ng1589)  &  (~ ng24478)  &  (~ wire7065) ) ;
 assign ng30293 = ( ng24433 ) | ( (~ ng4180)  &  wire6925 ) | ( ng1242  &  (~ ng24433)  &  (~ wire6925) ) ;
 assign ng28846 = ( ng112  &  ng29503  &  ng26314  &  wire29272 ) ;
 assign ng14727 = ( (~ ng5535) ) | ( (~ ng5511) ) | ( (~ ng5527) ) | ( ng5517 ) ;
 assign ng14755 = ( ng5188 ) | ( (~ ng5170) ) | ( ng5164 ) | ( (~ ng5180) ) ;
 assign ng19063 = ( pg12919  &  ng936  &  ng904  &  ng921 ) ;
 assign ng15674 = ( (~ pg12919) ) | ( (~ ng904) ) | ( (~ ng921) ) ;
 assign ng25290 = ( (~ ng5041)  &  (~ ng5046)  &  wire29316 ) ;
 assign ng13923 = ( (~ ng3530) ) | ( (~ ng3506) ) | ( (~ ng3522) ) | ( (~ ng3512) ) ;
 assign ng16187 = ( (~ ng4975) ) | ( (~ ng4966) ) | ( (~ ng4983) ) | ( (~ ng10862) ) ;
 assign ng28349 = ( (~ ng63) ) | ( (~ ng29503) ) | ( ng24380 ) | ( (~ wire29233) ) ;
 assign ng29008 = ( ng20739  &  (~ ng24380)  &  wire28640  &  wire29348 ) ;
 assign ng12228 = ( ng4486  &  ng4483  &  ng4489  &  ng4492 ) ;
 assign ng10909 = ( (~ pg13259) ) | ( ng1171 ) | ( ng1183 ) ;
 assign ng13336 = ( ng969  &  ng1193  &  (~ ng976) ) | ( ng1193  &  (~ ng976)  &  ng1008 ) ;
 assign ng27833 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28614) ) ;
 assign ng12432 = ( ng1917  &  (~ ng1894) ) ;
 assign ng14678 = ( ng1959  &  (~ ng1917) ) | ( ng1959  &  ng1894 ) ;
 assign ng32212 = ( (~ ng28504)  &  wire28813  &  (~ wire28814)  &  wire28815 ) ;
 assign ng22862 = ( pg35  &  pg12923 ) ;
 assign ng14142 = ( ng3873 ) | ( (~ ng3857) ) | ( ng3881 ) | ( (~ ng3863) ) ;
 assign ng8359 = ( (~ pg8358)  &  ng191 ) | ( pg8358  &  (~ ng191) ) ;
 assign ng8751 = ( (~ pg11418) ) | ( (~ pg16659) ) | ( (~ pg16775) ) | ( (~ pg13966) ) ;
 assign ng11893 = ( ng1668  &  (~ ng1636) ) ;
 assign ng15695 = ( (~ pg12923) ) | ( (~ ng1266) ) | ( (~ ng1249) ) ;
 assign ng19140 = ( pg12923  &  ng1266  &  ng1249  &  ng1280 ) ;
 assign ng25429 = ( wire30314 ) | ( (~ ng14367)  &  (~ wire6655) ) | ( (~ wire6655)  &  (~ wire29571) ) ;
 assign ng25389 = ( wire30349 ) | ( (~ ng14367)  &  (~ wire6319) ) | ( (~ wire6319)  &  (~ wire30342) ) ;
 assign ng7661 = ( (~ ng1211)  &  (~ ng1221)  &  (~ ng1216)  &  (~ ng1205) ) ;
 assign ng10695 = ( ng1171  &  ng1183 ) ;
 assign ng14908 = ( ng6573 ) | ( (~ ng6561) ) | ( (~ ng6565) ) ;
 assign ng24478 = ( wire7308 ) | ( wire7309 ) | ( ng1300  &  (~ ng1291) ) ;
 assign ng26793 = ( ng11003 ) | ( wire7065 ) | ( wire7308 ) | ( wire7309 ) ;
 assign ng29313 = ( ng24478 ) | ( (~ ng4180)  &  wire7065 ) | ( (~ ng1585)  &  (~ ng24478)  &  (~ wire7065) ) ;
 assign ng12405 = ( ng5188  &  (~ ng5180) ) ;
 assign ng14656 = ( (~ ng5188) ) | ( ng5170 ) | ( (~ ng5164) ) | ( ng5180 ) ;
 assign ng25233 = ( (~ ng5037)  &  (~ ng5041)  &  (~ ng17217) ) | ( ng5037  &  ng5041  &  (~ ng14317) ) ;
 assign ng27020 = ( ng4601  &  ng4593  &  ng24411 ) ;
 assign ng28144 = ( ng4601  &  ng4608  &  ng4593  &  ng24411 ) ;
 assign ng13156 = ( (~ ng7)  &  (~ ng6)  &  (~ ng8) ) ;
 assign ng25357 = ( pg73  &  pg72  &  ng2759  &  ng2763 ) | ( pg73  &  (~ pg72)  &  (~ ng2759)  &  ng2763 ) | ( (~ pg73)  &  pg72  &  ng2759  &  (~ ng2763) ) | ( (~ pg73)  &  (~ pg72)  &  (~ ng2759)  &  (~ ng2763) ) ;
 assign ng12812 = ( (~ ng513)  &  ng518 ) ;
 assign ng14855 = ( ng5881 ) | ( (~ ng5873) ) | ( ng5857 ) | ( (~ ng5863) ) ;
 assign ng11729 = ( ng3171  &  (~ ng3179) ) ;
 assign ng13951 = ( (~ ng3171) ) | ( ng3179 ) | ( (~ ng3167) ) ;
 assign ng10999 = ( ng1472  &  (~ ng1291) ) ;
 assign ng24471 = ( wire7308 ) | ( wire7309 ) | ( ng1472  &  (~ ng1291) ) ;
 assign ng31971 = ( (~ ng10511) ) | ( ng65  &  ng29503 ) | ( ng65  &  ng27972 ) ;
 assign ng13983 = ( ng3530 ) | ( ng3506 ) | ( ng3522 ) | ( (~ ng3512) ) ;
 assign ng11747 = ( (~ ng3530)  &  ng3522 ) ;
 assign ng14101 = ( (~ ng3171) ) | ( ng3179 ) | ( (~ ng3161) ) | ( (~ ng3155) ) ;
 assign ng25779 = ( (~ ng34) ) | ( (~ pg56)  &  pg54 ) ;
 assign ng10281 = ( (~ ng5535)  &  (~ ng5527) ) ;
 assign ng14927 = ( ng5535 ) | ( (~ ng5511) ) | ( ng5527 ) | ( (~ ng5517) ) ;
 assign ng12772 = ( (~ ng5188)  &  ng5180 ) ;
 assign ng14723 = ( ng5188 ) | ( (~ ng5176) ) | ( (~ ng5180) ) ;
 assign ng23309 = ( (~ ng3703) ) | ( (~ wire6966)  &  (~ wire6967)  &  (~ wire29216) ) ;
 assign ng14768 = ( (~ ng5881) ) | ( (~ ng5873) ) | ( (~ ng5857) ) | ( ng5863 ) ;
 assign ng29657 = ( ng11797  &  ng11261 ) | ( ng24374  &  (~ wire29730) ) ;
 assign ng28973 = ( ng2421 ) | ( (~ ng2465) ) | ( (~ ng26770)  &  (~ ng17424) ) ;
 assign ng23204 = ( (~ wire28543)  &  (~ wire28544)  &  wire28551 ) | ( (~ wire28543)  &  (~ wire28544)  &  wire28558 ) ;
 assign ng7675 = ( (~ ng1548)  &  (~ ng1559)  &  (~ ng1554)  &  (~ ng1564) ) ;
 assign ng7352 = ( (~ ng1514)  &  (~ ng1526) ) ;
 assign ng14506 = ( wire29058 ) | ( ng1430  &  (~ ng7675) ) | ( ng1430  &  (~ ng7352) ) ;
 assign ng11160 = ( pg17685  &  ng6381  &  ng6336  &  ng6395 ) ;
 assign ng21012 = ( wire7248 ) | ( wire7249 ) | ( wire28843 ) ;
 assign ng11405 = ( (~ ng2756) ) | ( (~ ng2735) ) | ( (~ ng2741) ) | ( (~ ng2748) ) ;
 assign ng14133 = ( ng3530 ) | ( (~ ng3506) ) | ( (~ ng3522) ) | ( (~ ng3512) ) ;
 assign ng23978 = ( (~ ng14708) ) | ( wire28793 ) | ( (~ wire28794) ) | ( wire28795 ) ;
 assign ng27395 = ( (~ ng504)  &  (~ ng518)  &  (~ ng528)  &  ng26314 ) ;
 assign ng28739 = ( ng112  &  ng29503  &  ng26314  &  wire30283 ) ;
 assign ng22498 = ( wire5887 ) | ( ng14367  &  wire31005 ) ;
 assign ng12629 = ( ng6573 ) | ( (~ ng6561) ) | ( ng6565 ) ;
 assign ng25341 = ( wire29573 ) | ( (~ ng14367)  &  (~ wire6655) ) | ( (~ wire6655)  &  (~ wire29571) ) ;
 assign ng27629 = ( (~ ng23978)  &  wire28796  &  (~ wire28801)  &  wire28802 ) ;
 assign ng14438 = ( wire29009 ) | ( ng1087  &  (~ ng7661) ) | ( ng1087  &  (~ ng7304) ) ;
 assign ng11432 = ( ng3171 ) | ( ng3179 ) | ( (~ ng3167) ) ;
 assign ng30576 = ( (~ wire1421)  &  (~ ng4818)  &  ng101  &  ng24374 ) ;
 assign ng12301 = ( (~ pg12300)  &  ng5689 ) | ( pg12300  &  (~ ng5689) ) ;
 assign ng27474 = ( ng504  &  ng518  &  ng528  &  ng26314 ) ;
 assign ng27445 = ( ng504  &  (~ ng518)  &  ng528  &  ng26314 ) ;
 assign ng17405 = ( wire29405 ) | ( pg17404  &  (~ ng7675) ) | ( pg17404  &  (~ ng10699) ) ;
 assign ng10721 = ( pg16624  &  ng3352  &  ng3338  &  ng3288 ) ;
 assign ng23067 = ( (~ ng10721) ) | ( (~ wire7137)  &  (~ wire7138)  &  (~ wire28996) ) ;
 assign ng12798 = ( (~ ng5535)  &  ng5527 ) ;
 assign ng14764 = ( ng5535 ) | ( (~ ng5523) ) | ( (~ ng5527) ) ;
 assign ng24460 = ( wire7308 ) | ( wire7309 ) | ( ng1448  &  (~ ng1291) ) ;
 assign ng26737 = ( ng10967 ) | ( wire6770 ) | ( wire7308 ) | ( wire7309 ) ;
 assign ni17529 = ( (~ ng31)  &  ng28  &  ng13156 ) ;
 assign ng12483 = ( ng2476  &  (~ ng2453) ) ;
 assign ng9649 = ( (~ ng2153)  &  (~ ng2227) ) ;
 assign ng11320 = ( (~ ng4633) ) | ( ng4639 ) | ( (~ ng4621) ) ;
 assign ng26218 = ( ng2756  &  (~ ng2741)  &  ng2748  &  ng25357 ) ;
 assign ng11773 = ( (~ ng4785)  &  ng4709 ) ;
 assign ng11834 = ( ng4975  &  ng4899 ) ;
 assign ng11283 = ( (~ ng4991)  &  ng4966  &  ng4983 ) ;
 assign ng11527 = ( ng3530  &  ng3522 ) ;
 assign ng13955 = ( (~ ng3530) ) | ( (~ ng3506) ) | ( (~ ng3522) ) | ( ng3512 ) ;
 assign ng14902 = ( (~ ng6215) ) | ( (~ ng6227) ) | ( ng6219 ) ;
 assign ng24447 = ( wire7308 ) | ( wire7309 ) | ( ng1478  &  (~ ng1291) ) ;
 assign ng26703 = ( ng10948 ) | ( wire7306 ) | ( wire7308 ) | ( wire7309 ) ;
 assign ng13134 = ( (~ pg12923) ) | ( (~ pg19357)  &  (~ pg7946)  &  (~ ng1333) ) ;
 assign ng26195 = ( ng2756  &  ng2741  &  (~ ng2748)  &  ng25357 ) ;
 assign ng11130 = ( (~ ng1221) ) | ( (~ ng1087) ) | ( (~ ng1205) ) ;
 assign ng34550 = ( (~ ng33851) ) | ( wire30331 ) | ( (~ wire30332) ) | ( wire32708 ) ;
 assign ng13948 = ( ng3171 ) | ( ng3179 ) | ( (~ ng3161) ) | ( ng3155 ) ;
 assign ng25498 = ( wire31232 ) | ( (~ ng14367)  &  (~ wire5887) ) | ( (~ wire5887)  &  (~ wire31005) ) ;
 assign ng25439 = ( wire32438 ) | ( (~ ng14367)  &  (~ wire5887) ) | ( (~ wire5887)  &  (~ wire31005) ) ;
 assign ng13986 = ( ng3530 ) | ( (~ ng3518) ) | ( (~ ng3522) ) ;
 assign ng12453 = ( ng5535  &  (~ ng5527) ) ;
 assign ng14807 = ( (~ ng5535) ) | ( (~ ng5523) ) | ( ng5527 ) ;
 assign ng28652 = ( (~ ng479)  &  ng890 ) | ( ng890  &  ng528 ) | ( ng890  &  (~ ng26314) ) ;
 assign ng13960 = ( ng3873 ) | ( (~ ng3857) ) | ( (~ ng3881) ) | ( ng3863 ) ;
 assign ng11435 = ( (~ ng3171)  &  ng3179 ) ;
 assign ng14008 = ( ng3171 ) | ( (~ ng3179) ) | ( (~ ng3161) ) | ( ng3155 ) ;
 assign ng27421 = ( (~ ng504)  &  (~ ng518)  &  ng528  &  ng26314 ) ;
 assign ng17321 = ( wire28783 ) | ( pg17320  &  (~ ng10671) ) | ( pg17320  &  (~ ng7675) ) ;
 assign ng12680 = ( ng6573  &  ng6565 ) ;
 assign ng15014 = ( (~ ng6573) ) | ( (~ ng6555) ) | ( ng6549 ) | ( (~ ng6565) ) ;
 assign ng25467 = ( (~ ng12432) ) | ( (~ ng14367)  &  (~ wire6655) ) | ( (~ wire6655)  &  (~ wire29571) ) ;
 assign ng25495 = ( (~ ng12483) ) | ( (~ ng14367)  &  (~ wire7725) ) | ( (~ wire7725)  &  (~ wire28488) ) ;
 assign ng25144 = ( (~ ng5037)  &  (~ ng5041)  &  (~ ng5046)  &  (~ ng17217) ) ;
 assign ng23560 = ( ng5037  &  ng5041  &  ng5046  &  (~ ng14317) ) ;
 assign ng27670 = ( (~ ng5052)  &  ng25144 ) | ( ng5052  &  ng23560 ) ;
 assign ng30286 = ( wire28637 ) | ( wire28638 ) ;
 assign ng25435 = ( wire31424 ) | ( (~ ng14367)  &  (~ wire7030) ) | ( (~ wire7030)  &  (~ wire29111) ) ;
 assign ng10266 = ( (~ ng5188)  &  (~ ng5180) ) ;
 assign ng12402 = ( ng5188 ) | ( (~ ng5176) ) | ( ng5180 ) ;
 assign ng13284 = ( (~ pg7916) ) | ( (~ ng1171) ) | ( (~ ng1183) ) ;
 assign ng14981 = ( (~ ng6573) ) | ( (~ ng6555) ) | ( ng6549 ) | ( ng6565 ) ;
 assign ng20248 = ( ng11676 ) | ( wire6781 ) | ( wire6784 ) | ( wire29397 ) ;
 assign ng17264 = ( (~ ng817) ) | ( (~ ng832) ) | ( ng8806 ) ;
 assign ng14279 = ( (~ ng837)  &  ng847 ) | ( ng812  &  ng847 ) ;
 assign ng13963 = ( (~ ng3873) ) | ( (~ ng3857) ) | ( (~ ng3881) ) | ( (~ ng3863) ) ;
 assign ng12933 = ( ng5022  &  (~ ng5016) ) | ( ng5016  &  ng5062 ) ;
 assign ng14665 = ( ng5535 ) | ( (~ ng5511) ) | ( (~ ng5527) ) | ( ng5517 ) ;
 assign ng26625 = ( (~ ng25144)  &  (~ ng23560) ) ;
 assign ng31950 = ( ng4643 ) | ( ng65  &  ng29503 ) | ( ng65  &  ng27972 ) ;
 assign ng11148 = ( ng1211  &  ng1221  &  ng1087  &  ng1205 ) ;
 assign ng10887 = ( ng6573  &  ng6561  &  ng6565 ) ;
 assign ng14720 = ( ng5188 ) | ( (~ ng5170) ) | ( ng5164 ) | ( ng5180 ) ;
 assign ng7567 = ( (~ ng990)  &  (~ ng979) ) ;
 assign ng30314 = ( ng24471 ) | ( (~ ng4180)  &  wire6912 ) | ( ng1585  &  (~ ng24471)  &  (~ wire6912) ) ;
 assign ng29719 = ( ng11261  &  ng11773 ) | ( ng24374  &  (~ wire29730) ) ;
 assign ng26994 = ( ng43  &  ng29503  &  ng24688  &  wire29502 ) ;
 assign ng23630 = ( (~ ng11123) ) | ( (~ wire6832)  &  (~ wire6833)  &  (~ wire29346) ) ;
 assign ng13570 = ( (~ ng1221) ) | ( (~ ng1087) ) | ( (~ ng1216) ) | ( (~ ng1205) ) ;
 assign ng10224 = ( (~ pg14828) ) | ( (~ pg12470) ) | ( (~ pg17778) ) | ( (~ pg17688) ) ;
 assign ng14075 = ( (~ ng3530) ) | ( ng3506 ) | ( (~ ng3522) ) | ( (~ ng3512) ) ;
 assign ng14999 = ( ng5881 ) | ( (~ ng5873) ) | ( (~ ng5857) ) | ( (~ ng5863) ) ;
 assign ng8347 = ( (~ ng4340) ) | ( (~ ng4349) ) | ( (~ ng4358) ) ;
 assign ng10823 = ( ng5188  &  ng5176  &  ng5180 ) ;
 assign ng12374 = ( (~ ng2185)  &  ng2208 ) ;
 assign ng22384 = ( wire6172 ) | ( ng14367  &  wire30555 ) ;
 assign ng25309 = ( wire30557 ) | ( (~ ng14367)  &  (~ wire6172) ) | ( (~ wire6172)  &  (~ wire30555) ) ;
 assign ng25396 = ( wire33307 ) | ( (~ ng14367)  &  (~ wire6172) ) | ( (~ wire6172)  &  (~ wire30555) ) ;
 assign ng14713 = ( (~ ng2476)  &  ng2518 ) | ( ng2453  &  ng2518 ) ;
 assign ng20682 = ( wire7624 ) | ( wire7625 ) | ( wire28651 ) ;
 assign ng28982 = ( ng20682  &  (~ ng24380)  &  wire28640  &  wire30578 ) ;
 assign ng14915 = ( ng5188 ) | ( ng5170 ) | ( (~ ng5164) ) | ( ng5180 ) ;
 assign ng11939 = ( ng2361  &  (~ ng2331) ) ;
 assign ng28833 = ( ng112  &  ng29503  &  ng26314  &  wire30377 ) ;
 assign ng7601 = ( (~ ng1322)  &  (~ ng1333) ) ;
 assign ng15748 = ( ng1312 ) | ( wire28718 ) | ( (~ ng7620)  &  wire28716 ) ;
 assign ng11869 = ( ng1345  &  ng1367  &  ng1379 ) ;
 assign ng14048 = ( (~ ng3530) ) | ( ng3506 ) | ( ng3522 ) | ( (~ ng3512) ) ;
 assign ng12505 = ( ng5535  &  ng5527 ) ;
 assign ng10838 = ( ng5535  &  ng5523  &  ng5527 ) ;
 assign ng14758 = ( (~ ng5188) ) | ( (~ ng5176) ) | ( ng5180 ) ;
 assign ng13889 = ( ng3171 ) | ( (~ ng3179) ) | ( ng3161 ) | ( (~ ng3155) ) ;
 assign ng12622 = ( ng6227  &  ng6219 ) ;
 assign ng10874 = ( ng6215  &  ng6227  &  ng6219 ) ;
 assign ng24411 = ( ng4584  &  (~ ng10511)  &  (~ ng8347)  &  (~ wire28475) ) ;
 assign ng26166 = ( (~ ng2756)  &  ng2741  &  (~ ng2748)  &  ng25357 ) ;
 assign ng13846 = ( (~ pg13259) ) | ( (~ ng1171) ) | ( ng1183 ) ;
 assign ng14899 = ( (~ ng6209) ) | ( ng6227 ) | ( ng6203 ) | ( (~ ng6219) ) ;
 assign ng12471 = ( (~ pg12470)  &  ng6727 ) | ( pg12470  &  (~ ng6727) ) ;
 assign ng14170 = ( ng3873 ) | ( (~ ng3857) ) | ( (~ ng3881) ) | ( (~ ng3863) ) ;
 assign ng8691 = ( (~ pg16718) ) | ( (~ pg16603) ) | ( (~ pg13895) ) | ( (~ pg11349) ) ;
 assign ng23618 = ( (~ ng2715)  &  (~ ng1945)  &  ng2719 ) | ( ng2715  &  (~ ng2079)  &  ng2719 ) ;
 assign ng14988 = ( ng7  &  ng6  &  ng8 ) ;
 assign ng10733 = ( pg16656  &  ng3689  &  ng3703  &  ng3639 ) ;
 assign ng10756 = ( pg16693  &  ng4040  &  ng4054  &  ng3990 ) ;
 assign ng15018 = ( (~ ng5881) ) | ( ng5873 ) | ( (~ ng5857) ) | ( (~ ng5863) ) ;
 assign ng28768 = ( ng112  &  ng29503  &  ng26314  &  wire30616 ) ;
 assign ng11483 = ( ng3530  &  (~ ng3522) ) ;
 assign ng10666 = ( (~ ng1171)  &  ng1183 ) ;
 assign ng10893 = ( ng1178  &  (~ ng1189)  &  ng996 ) ;
 assign ng14848 = ( (~ ng5535) ) | ( ng5511 ) | ( ng5527 ) | ( (~ ng5517) ) ;
 assign ng11292 = ( ng232  &  ng225  &  ng255 ) | ( (~ ng232)  &  (~ ng225)  &  ng255 ) | ( (~ ng232)  &  ng225  &  (~ ng255) ) | ( ng232  &  (~ ng225)  &  (~ ng255) ) ;
 assign ni27429 = ( ng93  &  ng29503 ) ;
 assign ng25851 = ( pg72  &  ng4322  &  wire28640 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640 ) ;
 assign ng29073 = ( ng21012  &  (~ ng24380)  &  wire28640  &  wire32672 ) ;
 assign ng28353 = ( ng150  &  ng164  &  ng23042  &  wire28708 ) ;
 assign ng25888 = ( (~ ng911) ) | ( (~ ng907) ) | ( (~ ng914) ) | ( (~ ng19063) ) ;
 assign ng23890 = ( (~ ng5357) ) | ( (~ wire7624)  &  (~ wire7625)  &  (~ wire28651) ) ;
 assign ng13346 = ( (~ ng4854) ) | ( (~ ng4849) ) | ( (~ ng4843) ) | ( (~ ng4878) ) ;
 assign ng9762 = ( (~ ng2495)  &  (~ ng2421) ) ;
 assign ng28927 = ( ng1862 ) | ( (~ ng1906) ) | ( (~ ng26725)  &  (~ ng17401) ) ;
 assign ng15033 = ( ng6573 ) | ( (~ ng6555) ) | ( (~ ng6549) ) | ( ng6565 ) ;
 assign ng12667 = ( (~ ng6215)  &  (~ ng6209)  &  (~ ng6203) ) ;
 assign ng20375 = ( ng671  &  (~ ng8806)  &  ng11185  &  wire30776 ) ;
 assign ng26256 = ( pg116  &  ng4157 ) | ( (~ pg115)  &  (~ ng4157) ) ;
 assign ng26212 = ( pg124  &  ng4146 ) | ( (~ pg126)  &  (~ ng4146) ) ;
 assign ng24627 = ( pg113  &  pg35 ) ;
 assign ng14864 = ( (~ ng6215) ) | ( ng6227 ) | ( (~ ng6219) ) ;
 assign ng31997 = ( wire6408 ) | ( ng65  &  ng29503 ) | ( ng65  &  ng27972 ) ;
 assign ng11171 = ( ng1548  &  ng1554  &  ng1564  &  ng1430 ) ;
 assign ng30307 = ( ng24460 ) | ( (~ ng4180)  &  wire6770 ) | ( (~ ng1585)  &  (~ ng24460)  &  (~ wire6770) ) ;
 assign ng28789 = ( ng112  &  ng29503  &  ng26314  &  wire30276 ) ;
 assign ng8728 = ( (~ pg13926) ) | ( (~ pg11388) ) | ( (~ pg16627) ) | ( (~ pg16744) ) ;
 assign ng20905 = ( (~ ng822) ) | ( (~ ng817) ) | ( (~ ng832) ) | ( ng8806 ) ;
 assign ng20751 = ( wire7046 ) | ( wire7047 ) | ( wire29091 ) ;
 assign ng29110 = ( ng93  &  ng29503  &  ng20751  &  wire30365 ) ;
 assign ng33394 = ( wire30386 ) | ( (~ ng27972)  &  (~ ng24374) ) | ( ng4507  &  (~ ng27972)  &  ng24374 ) ;
 assign ng25337 = ( (~ ng12729) ) | ( (~ ng14367)  &  (~ wire7041) ) | ( (~ wire7041)  &  (~ wire29097) ) ;
 assign ng13291 = ( (~ pg7946) ) | ( (~ ng1514) ) | ( (~ ng1526) ) ;
 assign ng13873 = ( (~ ng3171) ) | ( ng3179 ) | ( ng3161 ) | ( (~ ng3155) ) ;
 assign ng13980 = ( ng3171 ) | ( (~ ng3179) ) | ( (~ ng3167) ) ;
 assign ng25400 = ( wire30467 ) | ( (~ ng14367)  &  (~ wire7725) ) | ( (~ wire7725)  &  (~ wire28488) ) ;
 assign ng23553 = ( ng2815  &  (~ ng2715)  &  ng2719 ) | ( ng2715  &  ng2819  &  ng2719 ) ;
 assign ng23657 = ( ng2715  &  ng2719  &  (~ ng2638) ) | ( (~ ng2715)  &  ng2719  &  (~ ng2504) ) ;
 assign ng29036 = ( ng20875  &  (~ ng24380)  &  wire28640  &  wire31986 ) ;
 assign ng25895 = ( (~ ng1256) ) | ( (~ ng1259) ) | ( (~ ng1252) ) | ( (~ ng19140) ) ;
 assign ng25426 = ( (~ ng12371) ) | ( (~ ng14367)  &  (~ wire7257) ) | ( (~ wire7257)  &  (~ wire28834) ) ;
 assign ng13756 = ( ng513 ) | ( (~ ng518) ) | ( (~ ng203) ) ;
 assign ng27796 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28625) ) ;
 assign ng29496 = ( ng24471 ) | ( (~ ng4180)  &  wire6912 ) | ( ng1589  &  (~ ng24471)  &  (~ wire6912) ) ;
 assign ng11003 = ( ng1300  &  (~ ng1291) ) ;
 assign ng10862 = ( ng4859  &  ng4849  &  ng4843  &  ng4878 ) ;
 assign ng11245 = ( ng4087 ) | ( ng4098 ) | ( ng4093 ) ;
 assign ng25448 = ( wire3192 ) | ( (~ ng4064)  &  (~ ng4057)  &  wire34061 ) ;
 assign ng14069 = ( ng3171 ) | ( ng3179 ) | ( (~ ng3161) ) | ( (~ ng3155) ) ;
 assign ng14959 = ( ng5535 ) | ( (~ ng5511) ) | ( (~ ng5527) ) | ( (~ ng5517) ) ;
 assign ng12925 = ( (~ ng4340) ) | ( ng4639 ) | ( (~ ng4628) ) | ( (~ ng4621) ) ;
 assign ng25432 = ( (~ ng12374) ) | ( (~ ng14367)  &  (~ wire6172) ) | ( (~ wire6172)  &  (~ wire30555) ) ;
 assign ng11123 = ( pg17604  &  ng5689  &  ng5703  &  ng5644 ) ;
 assign ng12443 = ( ng5188  &  ng5180 ) ;
 assign ng14659 = ( (~ ng5188) ) | ( (~ ng5170) ) | ( (~ ng5164) ) | ( (~ ng5180) ) ;
 assign ng27469 = ( (~ ng504)  &  ng518  &  (~ ng528)  &  ng26314 ) ;
 assign ng28444 = ( ng291  &  ng287  &  ng283  &  ng23204 ) ;
 assign ng29001 = ( (~ ng2599) ) | ( ng2555 ) | ( (~ ng26793)  &  (~ ng14506) ) ;
 assign ng29486 = ( ng24447 ) | ( (~ ng4180)  &  wire7306 ) | ( ng1589  &  (~ ng24447)  &  (~ wire7306) ) ;
 assign ng11178 = ( pg17722  &  ng6741  &  ng6682  &  ng6727 ) ;
 assign ng11584 = ( ng3873  &  ng3881 ) ;
 assign ng13920 = ( (~ ng3530) ) | ( (~ ng3506) ) | ( ng3522 ) | ( ng3512 ) ;
 assign ng14688 = ( (~ ng5535) ) | ( (~ ng5511) ) | ( ng5527 ) | ( ng5517 ) ;
 assign ng12578 = ( (~ ng6215) ) | ( ng6227 ) | ( ng6219 ) ;
 assign ng11571 = ( (~ ng3506)  &  (~ ng3518)  &  (~ ng3512) ) ;
 assign ng25531 = ( (~ pg113) ) | ( (~ ng2868) ) ;
 assign ng10588 = ( ng5297  &  ng5357 ) ;
 assign ng31783 = ( wire29245 ) | ( wire29246 ) ;
 assign ng11006 = ( ng4653  &  ng4688  &  ng4659 ) ;
 assign ng13330 = ( (~ ng4653) ) | ( (~ ng4688) ) | ( (~ ng4664) ) | ( (~ ng4659) ) ;
 assign ng14627 = ( ng5188 ) | ( ng5170 ) | ( (~ ng5164) ) | ( (~ ng5180) ) ;
 assign ng14974 = ( (~ ng6209) ) | ( (~ ng6227) ) | ( ng6203 ) | ( (~ ng6219) ) ;
 assign ng14041 = ( (~ ng3171) ) | ( (~ ng3179) ) | ( (~ ng3161) ) | ( ng3155 ) ;
 assign ng27617 = ( ng43  &  ng29503  &  ng24688  &  wire29499 ) ;
 assign ng28626 = ( wire6178 ) | ( wire30547 ) | ( wire30551 ) | ( wire30552 ) ;
 assign ng14776 = ( (~ ng6209) ) | ( (~ ng6227) ) | ( (~ ng6203) ) | ( (~ ng6219) ) ;
 assign ng13517 = ( (~ ng3530)  &  ng3498 ) | ( ng3498  &  (~ ng3518) ) | ( ng3498  &  (~ ng3522) ) ;
 assign ng11916 = ( (~ ng2197)  &  ng2227 ) ;
 assign ng14825 = ( (~ ng6573) ) | ( (~ ng6555) ) | ( (~ ng6549) ) | ( (~ ng6565) ) ;
 assign ng23972 = ( (~ ng6741) ) | ( (~ wire7046)  &  (~ wire7047)  &  (~ wire29091) ) ;
 assign ng14640 = ( (~ ng1783)  &  ng1825 ) | ( ng1825  &  ng1760 ) ;
 assign ng23324 = ( (~ ng703) ) | ( ng16846  &  wire30802 ) | ( ng16846  &  wire30803 ) ;
 assign ng16846 = ( ng499  &  (~ ng504)  &  (~ ng8806)  &  ng11185 ) ;
 assign ng14247 = ( ng5849  &  (~ ng5869) ) | ( ng5849  &  (~ ng5881) ) | ( ng5849  &  (~ ng5873) ) ;
 assign ng12479 = ( ng2051  &  (~ ng2028) ) ;
 assign ng10869 = ( ng5869  &  ng5881  &  ng5873 ) ;
 assign ng14761 = ( ng5535 ) | ( ng5511 ) | ( ng5527 ) | ( (~ ng5517) ) ;
 assign ng28220 = ( wire32354 ) | ( wire32355 ) | ( wire32357 ) | ( wire32358 ) ;
 assign ng23286 = ( (~ ng3352) ) | ( (~ wire7137)  &  (~ wire7138)  &  (~ wire28996) ) ;
 assign ng14098 = ( ng3171 ) | ( ng3179 ) | ( ng3161 ) | ( (~ ng3155) ) ;
 assign ng27738 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28632) ) ;
 assign ng7598 = ( (~ ng979)  &  ng996 ) | ( ng979  &  (~ ng996) ) ;
 assign ng13211 = ( (~ ng990)  &  (~ ng979) ) | ( ng979  &  ng996 ) | ( (~ ng979)  &  (~ ng996) ) ;
 assign ng22654 = ( ng4087  &  ng4093  &  ng4076  &  (~ ng13217) ) ;
 assign ng26171 = ( ng2756  &  (~ ng2741)  &  (~ ng2748)  &  ng25357 ) ;
 assign ng15591 = ( (~ ng4332) ) | ( (~ ng4322) ) | ( ng10511 ) | ( ng8347 ) ;
 assign ng14085 = ( (~ ng3873) ) | ( (~ ng3881) ) | ( (~ ng3869) ) ;
 assign ng28853 = ( (~ ng1636) ) | ( ng1592 ) | ( (~ ng26673)  &  (~ ng17292) ) ;
 assign ng11419 = ( (~ pg11418)  &  ng4040 ) | ( pg11418  &  (~ ng4040) ) ;
 assign ng11255 = ( (~ ng4054)  &  ng3990 ) ;
 assign ng14018 = ( (~ ng3530) ) | ( (~ ng3518) ) | ( ng3522 ) ;
 assign ng11139 = ( pg17646  &  ng6035  &  ng5990  &  ng6049 ) ;
 assign ng14051 = ( (~ ng3530) ) | ( (~ ng3518) ) | ( (~ ng3522) ) ;
 assign ng24433 = ( wire7608 ) | ( wire7609 ) | ( ng1135  &  (~ ng947) ) ;
 assign ng26673 = ( ng10878 ) | ( wire6925 ) | ( wire7608 ) | ( wire7609 ) ;
 assign ng14813 = ( (~ ng5869) ) | ( ng5881 ) | ( (~ ng5873) ) ;
 assign ng11111 = ( pg17577  &  ng5297  &  ng5357  &  ng5343 ) ;
 assign ng12239 = ( (~ pg12238)  &  ng5343 ) | ( pg12238  &  (~ ng5343) ) ;
 assign ng12423 = ( (~ pg12422)  &  ng6381 ) | ( pg12422  &  (~ ng6381) ) ;
 assign ng9586 = ( (~ ng1668)  &  (~ ng1592) ) ;
 assign ng15042 = ( ng6573 ) | ( (~ ng6555) ) | ( (~ ng6549) ) | ( (~ ng6565) ) ;
 assign ng12492 = ( (~ ng5170)  &  (~ ng5176)  &  (~ ng5164) ) ;
 assign ng14127 = ( ng3171 ) | ( (~ ng3179) ) | ( (~ ng3161) ) | ( (~ ng3155) ) ;
 assign ng7620 = ( (~ ng1322)  &  ng1339 ) | ( ng1322  &  (~ ng1339) ) ;
 assign ng14879 = ( ng5188 ) | ( (~ ng5170) ) | ( (~ ng5164) ) | ( ng5180 ) ;
 assign ng28962 = ( ng1996 ) | ( (~ ng2040) ) | ( (~ ng26759)  &  (~ ng14438) ) ;
 assign ng14953 = ( (~ ng5188) ) | ( (~ ng5170) ) | ( (~ ng5164) ) | ( ng5180 ) ;
 assign ng27933 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28622) ) ;
 assign ng27854 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28629) ) ;
 assign ng11978 = ( (~ ng2599)  &  ng2629 ) ;
 assign ng29722 = ( ng11780  &  ng11283 ) | ( ng24374  &  (~ wire28575) ) ;
 assign ng14055 = ( (~ ng3873) ) | ( ng3857 ) | ( ng3881 ) | ( (~ ng3863) ) ;
 assign ng14968 = ( ng5881 ) | ( ng5873 ) | ( (~ ng5857) ) | ( (~ ng5863) ) ;
 assign ng11937 = ( ng1936  &  (~ ng1906) ) ;
 assign ng13929 = ( (~ ng3873) ) | ( (~ ng3857) ) | ( ng3881 ) | ( ng3863 ) ;
 assign ng30298 = ( ng24444 ) | ( (~ ng4180)  &  wire7606 ) | ( (~ ng1242)  &  (~ ng24444)  &  (~ wire7606) ) ;
 assign ng14797 = ( (~ ng5188) ) | ( (~ ng5170) ) | ( ng5164 ) | ( ng5180 ) ;
 assign ng28020 = ( ng43  &  ng29503  &  ng24688  &  wire29491 ) ;
 assign ng29489 = ( ng24460 ) | ( (~ ng4180)  &  wire6770 ) | ( (~ ng1589)  &  (~ ng24460)  &  (~ wire6770) ) ;
 assign ng14679 = ( (~ ng2342)  &  ng2384 ) | ( ng2319  &  ng2384 ) ;
 assign ng9724 = ( (~ ng5092) ) | ( (~ ng5084) ) ;
 assign ng27882 = ( (~ ng110) ) | ( (~ ng29503) ) | ( (~ ng25357) ) | ( (~ wire28617) ) ;
 assign ng10185 = ( (~ pg14738) ) | ( (~ pg17607) ) | ( (~ pg17739) ) | ( (~ pg12350) ) ;
 assign ng13260 = ( (~ pg13259) ) | ( ng1171 ) | ( (~ ng1183) ) ;
 assign ng8933 = ( (~ ng4785)  &  (~ ng4709) ) ;
 assign ng23554 = ( ng2775  &  ng2724  &  (~ ng2729) ) | ( (~ ng2724)  &  (~ ng2729)  &  ng2771 ) ;
 assign ng10878 = ( ng1135  &  (~ ng947) ) ;
 assign ng15585 = ( (~ ng5022)  &  (~ ng5029) ) | ( (~ ng5029)  &  ng5016 ) | ( (~ ng5022)  &  (~ ng5016) ) | ( ng5029  &  (~ ng5016) ) | ( (~ ng5022)  &  (~ ng5062) ) | ( ng5029  &  (~ ng5062) ) | ( ng5016  &  (~ ng5062) ) ;
 assign ng27416 = ( ng504  &  (~ ng518)  &  (~ ng528)  &  ng26314 ) ;
 assign ng26148 = ( (~ ng2756)  &  (~ ng2741)  &  (~ ng2748)  &  ng25357 ) ;
 assign ng26213 = ( (~ ng2756)  &  ng2741  &  ng2748  &  ng25357 ) ;
 assign ng11763 = ( ng3873  &  (~ ng3881) ) ;
 assign ng23909 = ( (~ ng5703) ) | ( (~ wire6832)  &  (~ wire6833)  &  (~ wire29346) ) ;
 assign ng7304 = ( (~ ng1171)  &  (~ ng1183) ) ;
 assign ng14956 = ( ng5535 ) | ( (~ ng5511) ) | ( ng5527 ) | ( ng5517 ) ;
 assign ng29702 = ( ng11283  &  ng8984 ) | ( ng24374  &  (~ wire28575) ) ;
 assign ng13121 = ( (~ pg12919) ) | ( (~ pg19334)  &  (~ pg7916)  &  (~ ng990) ) ;
 assign ng12540 = ( ng2610  &  (~ ng2587) ) ;
 assign ng25514 = ( (~ ng12540) ) | ( (~ ng14367)  &  (~ wire5887) ) | ( (~ wire5887)  &  (~ wire31005) ) ;
 assign ng14984 = ( (~ ng6573) ) | ( (~ ng6561) ) | ( (~ ng6565) ) ;
 assign ng14130 = ( ng3530 ) | ( (~ ng3506) ) | ( ng3522 ) | ( ng3512 ) ;
 assign ng14151 = ( (~ ng3530) ) | ( (~ ng3506) ) | ( ng3522 ) | ( (~ ng3512) ) ;
 assign ng14752 = ( (~ ng2610)  &  ng2652 ) | ( ng2652  &  ng2587 ) ;
 assign ng25492 = ( (~ ng12479) ) | ( (~ ng14367)  &  (~ wire6319) ) | ( (~ wire6319)  &  (~ wire30342) ) ;
 assign ng8721 = ( pg8719  &  ng385  &  ng376 ) ;
 assign ng28799 = ( ng112  &  ng29503  &  ng26314  &  wire30356 ) ;
 assign ng28471 = ( ng93  &  ng29503  &  ng21024  &  wire31435 ) ;
 assign ng28892 = ( (~ ng1772) ) | ( ng1728 ) | ( (~ ng17317)  &  (~ ng26694) ) ;
 assign ng23586 = ( (~ ng5037)  &  ng17217 ) | ( ng5037  &  ng14317 ) | ( ng17217  &  ng14317 ) ;
 assign ng14211 = ( (~ ng5188)  &  ng5156 ) | ( ng5156  &  (~ ng5176) ) | ( ng5156  &  (~ ng5180) ) ;
 assign ng29730 = ( ng25851  &  wire29253 ) | ( ng25776  &  wire29254 ) ;
 assign ng24380 = ( (~ pg72)  &  ng4322 ) | ( pg72  &  (~ ng4322) ) ;
 assign ng10699 = ( (~ ng1514)  &  ng1526 ) ;
 assign ng10918 = ( (~ ng1532)  &  ng1521  &  ng1339 ) ;
 assign ng14892 = ( (~ ng5881) ) | ( ng5873 ) | ( ng5857 ) | ( (~ ng5863) ) ;
 assign ng11956 = ( ng2070  &  (~ ng2040) ) ;
 assign ng25537 = ( (~ pg113) ) | ( (~ ng2873) ) ;
 assign ng12450 = ( ng5535 ) | ( (~ ng5523) ) | ( ng5527 ) ;
 assign ng8984 = ( (~ ng4975)  &  (~ ng4899) ) ;
 assign ng14943 = ( (~ ng6215) ) | ( (~ ng6227) ) | ( (~ ng6219) ) ;
 assign ng17317 = ( wire28673 ) | ( pg17316  &  (~ ng7661) ) | ( pg17316  &  (~ ng10666) ) ;
 assign ng12558 = ( (~ ng5523)  &  (~ ng5511)  &  (~ ng5517) ) ;
 assign ng13486 = ( (~ ng4966) ) | ( (~ ng4983) ) | ( (~ ng10862) ) ;
 assign ng28484 = ( ni27429  &  wire28765  &  wire32239 ) | ( ni27429  &  wire28766  &  wire32239 ) ;
 assign ng10890 = ( (~ ng947)  &  ng1105 ) ;
 assign ni30751 = ( wire30158 ) | ( wire30159 ) | ( wire30160 ) ;
 assign ng14157 = ( (~ ng3873) ) | ( (~ ng3857) ) | ( ng3881 ) | ( (~ ng3863) ) ;
 assign ng14918 = ( ng5188 ) | ( (~ ng5170) ) | ( (~ ng5164) ) | ( (~ ng5180) ) ;
 assign ng14154 = ( ng3873 ) | ( (~ ng3857) ) | ( ng3881 ) | ( ng3863 ) ;
 assign ng13500 = ( (~ ng3171)  &  ng3147 ) | ( (~ ng3179)  &  ng3147 ) | ( ng3147  &  (~ ng3167) ) ;
 assign ng14732 = ( (~ ng5881) ) | ( ng5873 ) | ( (~ ng5857) ) | ( ng5863 ) ;
 assign ng10649 = ( ng1171  &  (~ ng1183) ) ;
 assign ng17292 = ( wire29263 ) | ( pg17291  &  (~ ng7661) ) | ( pg17291  &  (~ ng10649) ) ;
 assign ng16696 = ( wire30515 ) | ( wire30516 ) ;
 assign ng14800 = ( (~ ng5188) ) | ( (~ ng5176) ) | ( (~ ng5180) ) ;
 assign ng11737 = ( (~ pg8291) ) | ( (~ ng218) ) | ( (~ pg8358)  &  ng191 ) | ( pg8358  &  (~ ng191) ) ;
 assign ng9755 = ( (~ ng2070)  &  (~ ng1996) ) ;
 assign ng14841 = ( (~ ng5188) ) | ( (~ ng5170) ) | ( ng5164 ) | ( (~ ng5180) ) ;
 assign ng14024 = ( (~ ng3873) ) | ( ng3881 ) | ( (~ ng3869) ) ;
 assign ng22585 = ( wire32542 ) | ( wire32543 ) | ( wire32544 ) | ( wire32545 ) ;
 assign ng12351 = ( (~ pg12350)  &  ng6035 ) | ( pg12350  &  (~ ng6035) ) ;
 assign ng11846 = ( ng1002  &  ng1036  &  ng1024 ) ;
 assign ng16272 = ( (~ ng1322)  &  ng1579  &  (~ ng13242)  &  (~ wire30238) ) | ( ng1322  &  (~ ng1579)  &  (~ ng13242)  &  (~ wire30238) ) ;
 assign ng28458 = ( ng93  &  ng29503  &  ng20887  &  wire31757 ) ;
 assign ng11144 = ( ng246  &  ng232  &  ng239  &  wire28549 ) ;
 assign ng14773 = ( ng6209 ) | ( (~ ng6227) ) | ( (~ ng6203) ) | ( ng6219 ) ;
 assign ng14227 = ( (~ ng5535)  &  ng5503 ) | ( (~ ng5523)  &  ng5503 ) | ( (~ ng5527)  &  ng5503 ) ;
 assign ng23532 = ( (~ ng2715)  &  ng2719  &  ng2783 ) | ( ng2715  &  ng2719  &  ng2787 ) ;
 assign ng10948 = ( ng1478  &  (~ ng1291) ) ;
 assign ng14082 = ( ng3873 ) | ( ng3857 ) | ( (~ ng3881) ) | ( (~ ng3863) ) ;
 assign ng14895 = ( (~ ng5869) ) | ( (~ ng5881) ) | ( (~ ng5873) ) ;
 assign ng14933 = ( (~ ng5881) ) | ( (~ ng5873) ) | ( ng5857 ) | ( (~ ng5863) ) ;
 assign ng23342 = ( (~ ng4054) ) | ( (~ wire7325)  &  (~ wire7326)  &  (~ wire28766) ) ;
 assign ng24444 = ( wire7608 ) | ( wire7609 ) | ( (~ ng947)  &  ng1105 ) ;
 assign ng26694 = ( ng10890 ) | ( wire7606 ) | ( wire7608 ) | ( wire7609 ) ;
 assign ng11326 = ( (~ pg8719) ) | ( ng385 ) | ( (~ ng370) ) | ( (~ ng376) ) ;
 assign ng10124 = ( (~ pg17674) ) | ( (~ pg14662) ) | ( (~ pg17519) ) | ( (~ pg12238) ) ;
 assign ng11149 = ( (~ ng1548) ) | ( (~ ng1564) ) | ( (~ ng1430) ) ;
 assign ng13597 = ( (~ ng1548) ) | ( (~ ng1559) ) | ( (~ ng1564) ) | ( (~ ng1430) ) ;
 assign ng13898 = ( ng3530 ) | ( (~ ng3506) ) | ( (~ ng3522) ) | ( ng3512 ) ;
 assign ng14691 = ( (~ ng5535) ) | ( (~ ng5511) ) | ( (~ ng5527) ) | ( (~ ng5517) ) ;
 assign ng29482 = ( ng24433 ) | ( (~ ng4180)  &  wire6925 ) | ( ng1246  &  (~ ng24433)  &  (~ wire6925) ) ;
 assign ng14011 = ( (~ ng3171) ) | ( (~ ng3179) ) | ( (~ ng3167) ) ;
 assign ng23949 = ( (~ ng6395) ) | ( (~ wire7248)  &  (~ wire7249)  &  (~ wire28843) ) ;
 assign ng14851 = ( (~ ng5535) ) | ( (~ ng5523) ) | ( (~ ng5527) ) ;
 assign ng13990 = ( (~ ng3873) ) | ( (~ ng3857) ) | ( (~ ng3881) ) | ( ng3863 ) ;
 assign ng26236 = ( ng2756  &  ng2741  &  ng2748  &  ng25357 ) ;
 assign ng23975 = ( (~ ng417)  &  wire32031 ) | ( (~ ng417)  &  wire32032 ) | ( ng417  &  (~ wire32031)  &  (~ wire32032) ) ;
 assign ng13657 = ( ng452  &  ng392 ) | ( ng174  &  (~ ng392) ) ;
 assign ng14804 = ( ng5535 ) | ( ng5511 ) | ( (~ ng5527) ) | ( (~ ng5517) ) ;
 assign ng12729 = ( (~ ng1657)  &  ng1648 ) ;
 assign ng14817 = ( ng6209 ) | ( (~ ng6227) ) | ( (~ ng6203) ) | ( (~ ng6219) ) ;
 assign ng14712 = ( ng2093  &  (~ ng2051) ) | ( ng2093  &  ng2028 ) ;
 assign ng13539 = ( (~ ng3873)  &  ng3849 ) | ( (~ ng3881)  &  ng3849 ) | ( (~ ng3869)  &  ng3849 ) ;
 assign ng13464 = ( (~ ng4793) ) | ( (~ ng4776) ) | ( (~ ng10831) ) ;
 assign ng28504 = ( (~ ng24875) ) | ( wire28810 ) | ( (~ wire28811) ) | ( wire28812 ) ;
 assign ng29694 = ( ng11261  &  ng11755 ) | ( ng24374  &  (~ wire29730) ) ;
 assign ng28942 = ( ng2287 ) | ( (~ ng2331) ) | ( (~ ng17405)  &  (~ ng26737) ) ;
 assign ng28440 = ( wire4764 ) | ( wire32301 ) | ( wire32305 ) | ( wire32306 ) ;
 assign ng14611 = ( ng1624  &  ng1691 ) | ( ng1691  &  (~ ng1648) ) ;
 assign ng9640 = ( (~ ng1728)  &  (~ ng1802) ) ;
 assign ng8476 = ( pg7946 ) | ( pg8475 ) | ( wire33480 ) ;
 assign ng15021 = ( ng6209 ) | ( ng6227 ) | ( (~ ng6203) ) | ( ng6219 ) ;
 assign ng30605 = ( wire31726 ) | ( wire31727 ) ;
 assign ng15024 = ( (~ ng6209) ) | ( ng6227 ) | ( (~ ng6203) ) | ( (~ ng6219) ) ;
 assign ng29495 = ( ng24468 ) | ( (~ ng4180)  &  wire7126 ) | ( (~ ng1246)  &  (~ ng24468)  &  (~ wire7126) ) ;
 assign ng14116 = ( (~ ng3873) ) | ( ng3857 ) | ( (~ ng3881) ) | ( (~ ng3863) ) ;
 assign ng14110 = ( ng3530 ) | ( (~ ng3506) ) | ( ng3522 ) | ( (~ ng3512) ) ;
 assign ng9700 = ( (~ ng2361)  &  (~ ng2287) ) ;
 assign ng16757 = ( wire30517 ) | ( wire30518 ) ;
 assign ng17217 = ( (~ ng5022) ) | ( ng5029 ) | ( ng5016 ) | ( ng5033 ) ;
 assign ng14317 = ( (~ ng5029) ) | ( (~ ng5016) ) | ( (~ ng5062) ) | ( (~ ng5033) ) ;
 assign ng14993 = ( (~ ng5535) ) | ( (~ ng5511) ) | ( ng5527 ) | ( (~ ng5517) ) ;
 assign ng13915 = ( (~ ng3171) ) | ( (~ ng3179) ) | ( ng3161 ) | ( (~ ng3155) ) ;
 assign ng15008 = ( (~ ng6209) ) | ( ng6227 ) | ( (~ ng6203) ) | ( ng6219 ) ;
 assign ng14940 = ( (~ ng6209) ) | ( (~ ng6227) ) | ( ng6203 ) | ( ng6219 ) ;
 assign ng16663 = ( wire32269 ) | ( wire32270 ) ;
 assign ng25476 = ( wire32948 ) | ( (~ ng14367)  &  (~ wire7725) ) | ( (~ wire7725)  &  (~ wire28488) ) ;
 assign ng33851 = ( (~ ng31509)  &  wire30328  &  (~ wire30329)  &  wire30330 ) ;
 assign ng21284 = ( ng732  &  ng11676 ) | ( ng732  &  (~ wire28525) ) | ( ng732  &  (~ wire28526) ) ;
 assign ng14810 = ( ng5881 ) | ( ng5873 ) | ( ng5857 ) | ( (~ ng5863) ) ;
 assign ng29485 = ( ng24444 ) | ( (~ ng4180)  &  wire7606 ) | ( (~ ng1246)  &  (~ ng24444)  &  (~ wire7606) ) ;
 assign ng14642 = ( ng2185  &  ng2250 ) | ( ng2250  &  (~ ng2208) ) ;
 assign ng34056 = ( ni30751  &  (~ ni30745)  &  (~ wire30150) ) | ( (~ ni30745)  &  (~ wire30150)  &  wire30182 ) | ( (~ ni30751)  &  ni30745  &  (~ wire30182) ) | ( (~ ni30751)  &  wire30150  &  (~ wire30182) ) ;
 assign ng34051 = ( (~ ng33212)  &  ng33219 ) | ( ng33212  &  (~ ng33219) ) ;
 assign ng34424 = ( (~ ng33149)  &  ng33176  &  ng33164  &  ng33187 ) | ( ng33149  &  (~ ng33176)  &  ng33164  &  ng33187 ) | ( ng33149  &  ng33176  &  (~ ng33164)  &  ng33187 ) | ( (~ ng33149)  &  (~ ng33176)  &  (~ ng33164)  &  ng33187 ) | ( ng33149  &  ng33176  &  ng33164  &  (~ ng33187) ) | ( (~ ng33149)  &  (~ ng33176)  &  ng33164  &  (~ ng33187) ) | ( (~ ng33149)  &  ng33176  &  (~ ng33164)  &  (~ ng33187) ) | ( ng33149  &  (~ ng33176)  &  (~ ng33164)  &  (~ ng33187) ) ;
 assign ng16728 = ( wire32271 ) | ( wire32272 ) ;
 assign ng9835 = ( (~ ng2555)  &  (~ ng2629) ) ;
 assign ni30745 = ( wire30131 ) | ( wire30132 ) | ( wire30136 ) ;
 assign ng12332 = ( (~ ng246)  &  ng262  &  ng269  &  ng239 ) | ( ng246  &  (~ ng262)  &  ng269  &  ng239 ) | ( ng246  &  ng262  &  (~ ng269)  &  ng239 ) | ( (~ ng246)  &  (~ ng262)  &  (~ ng269)  &  ng239 ) | ( ng246  &  ng262  &  ng269  &  (~ ng239) ) | ( (~ ng246)  &  (~ ng262)  &  ng269  &  (~ ng239) ) | ( (~ ng246)  &  ng262  &  (~ ng269)  &  (~ ng239) ) | ( ng246  &  (~ ng262)  &  (~ ng269)  &  (~ ng239) ) ;
 assign pg8353 = ( wire1411 ) ;
 assign pg33533 = ( ng17292 ) ;
 assign pg34437 = ( ng25531 ) ;
 assign pg8132 = ( wire1421 ) ;
 assign pg31521 = ( ng25448 ) ;
 assign pg18101 = ( pg6746 ) ;
 assign pg34435 = ( ng25448 ) ;
 assign pg18100 = ( pg6751 ) ;
 assign pg20899 = ( ng79 ) ;
 assign pg34436 = ( ng25537 ) ;
 assign pg20557 = ( ng86 ) ;
 assign pg20654 = ( ng121 ) ;
 assign pg24171 = ( pg92 ) ;
 assign pg24182 = ( pg127 ) ;
 assign pg33894 = ( ng28652 ) ;
 assign pg8235 = ( wire1457 ) ;
 assign pg24172 = ( pg99 ) ;
 assign pg24181 = ( pg126 ) ;
 assign pg8403 = ( wire1411 ) ;
 assign pg24162 = ( pg54 ) ;
 assign pg24180 = ( pg125 ) ;
 assign pg26801 = ( ng10823 ) ;
 assign pg34237 = ( ng34237 ) ;
 assign pg20763 = ( ng74 ) ;
 assign pg24161 = ( pg53 ) ;
 assign pg24170 = ( pg91 ) ;
 assign pg34238 = ( ng34237 ) ;
 assign pg18097 = ( pg6747 ) ;
 assign pg24164 = ( pg57 ) ;
 assign pg24175 = ( pg114 ) ;
 assign pg29211 = ( ng74 ) ;
 assign pg34235 = ( ng34235 ) ;
 assign pg18098 = ( pg6744 ) ;
 assign pg20901 = ( ng102 ) ;
 assign pg24163 = ( pg56 ) ;
 assign pg24176 = ( pg115 ) ;
 assign pg24185 = ( pg44 ) ;
 assign pg29210 = ( ng59 ) ;
 assign pg18099 = ( pg6745 ) ;
 assign pg20652 = ( ng94 ) ;
 assign pg24166 = ( pg72 ) ;
 assign pg24173 = ( pg100 ) ;
 assign pg24184 = ( pg135 ) ;
 assign pg29213 = ( ng86 ) ;
 assign pg29220 = ( ng128 ) ;
 assign pg34233 = ( ng34235 ) ;
 assign pg21292 = ( ng136 ) ;
 assign pg24165 = ( pg64 ) ;
 assign pg24174 = ( pg113 ) ;
 assign pg24183 = ( pg134 ) ;
 assign pg29212 = ( ng79 ) ;
 assign pg29221 = ( ng136 ) ;
 assign pg32975 = ( ng10823 ) ;
 assign pg34234 = ( ng34235 ) ;
 assign pg34788 = ( ng28652 ) ;
 assign pg24168 = ( pg84 ) ;
 assign pg24179 = ( pg124 ) ;
 assign pg25219 = ( ng5343 ) ;
 assign pg29215 = ( ng102 ) ;
 assign pg30332 = ( ng1242 ) ;
 assign pg24167 = ( pg73 ) ;
 assign pg29214 = ( ng94 ) ;
 assign pg24177 = ( pg116 ) ;
 assign pg25167 = ( ng12729 ) ;
 assign pg29217 = ( ng117 ) ;
 assign pg34240 = ( ng34237 ) ;
 assign pg24169 = ( pg90 ) ;
 assign pg24178 = ( pg120 ) ;
 assign pg29216 = ( ng106 ) ;
 assign pg20049 = ( ng59 ) ;
 assign pg25259 = ( ng11893 ) ;
 assign pg25583 = ( ng25590 ) ;
 assign pg29219 = ( ng121 ) ;
 assign pg33959 = ( ng20682 ) ;
 assign pg21245 = ( ng128 ) ;
 assign pg25584 = ( ng25590 ) ;
 assign pg29218 = ( ng66 ) ;
 assign pg25585 = ( ng25590 ) ;
 assign pg18092 = ( pg6753 ) ;
 assign pg25586 = ( ng25590 ) ;
 assign pg21176 = ( ng106 ) ;
 assign pg25114 = ( ng10588 ) ;
 assign pg25590 = ( ng25590 ) ;
 assign pg18094 = ( pg6748 ) ;
 assign pg18881 = ( ng66 ) ;
 assign pg23683 = ( ng1242 ) ;
 assign pg18095 = ( pg6749 ) ;
 assign pg18096 = ( pg6750 ) ;
 assign pg21270 = ( ng117 ) ;
 assign pg25582 = ( ng25590 ) ;
 assign pg31863 = ( ng12729 ) ;
 assign pg27831 = ( ng17292 ) ;
 assign pg31861 = ( ng5343 ) ;
 assign pg31862 = ( ng11893 ) ;
 assign pg8283 = ( wire1457 ) ;
 assign pg25587 = ( ng25590 ) ;
 assign pg31665 = ( ng25531 ) ;
 assign pg21698 = ( pg36 ) ;
 assign pg25588 = ( ng25590 ) ;
 assign pg31860 = ( ng10588 ) ;
 assign pg25589 = ( ng25590 ) ;
 assign pg28753 = ( ng20682 ) ;
 assign pg31656 = ( ng25537 ) ;
 assign pg8178 = ( wire1421 ) ;
 assign wire3134 = ( ng2927  &  ng2922 ) ;
 assign wire3137 = ( (~ ni30330)  &  (~ ng31070)  &  wire34258  &  wire34259 ) ;
 assign wire3138 = ( ng31070  &  wire34230  &  wire34265 ) ;
 assign wire3139 = ( ni31121  &  (~ ng31070)  &  wire34266  &  wire34267 ) ;
 assign wire3140 = ( ni31171  &  (~ ng31070)  &  wire34202  &  wire34242 ) ;
 assign wire3141 = ( (~ ng31710)  &  (~ ng31070)  &  wire34241  &  wire34271 ) ;
 assign wire3148 = ( (~ ni30330)  &  (~ ng31070)  &  wire34225  &  wire34226 ) ;
 assign wire3149 = ( ng31070  &  wire34230  &  wire34234 ) ;
 assign wire3150 = ( ni31121  &  (~ ng31070)  &  wire34235  &  wire34236 ) ;
 assign wire3151 = ( (~ ng30673)  &  ni31171  &  (~ ng31070)  &  wire34242 ) ;
 assign wire3152 = ( (~ ng31710)  &  (~ ng31070)  &  wire34241  &  wire34244 ) ;
 assign wire3155 = ( ni31141  &  (~ ng31070)  &  wire34207  &  wire34208 ) ;
 assign wire3156 = ( ni31191  &  (~ ng31070)  &  wire34211  &  wire34212 ) ;
 assign wire3157 = ( ni31271  &  (~ ng31070)  &  wire34215  &  wire34216 ) ;
 assign wire3158 = ( ni31106  &  (~ ng31070)  &  wire34219  &  wire34220 ) ;
 assign wire3159 = ( (~ ng31021)  &  ni31141  &  wire34169  &  wire34170 ) ;
 assign wire3160 = ( (~ ng31021)  &  ni31191  &  wire34173  &  wire34174 ) ;
 assign wire3161 = ( (~ ng31021)  &  ni31271  &  wire34177  &  wire34178 ) ;
 assign wire3162 = ( ni31106  &  (~ ng31021)  &  wire34181  &  wire34182 ) ;
 assign wire3163 = ( (~ ni30330)  &  wire34185  &  wire34186 ) ;
 assign wire3164 = ( (~ ng31021)  &  (~ ni30330)  &  (~ ng31327)  &  wire34189 ) ;
 assign wire3165 = ( (~ ni30330)  &  (~ ng31710)  &  (~ ng31070)  &  wire34156 ) ;
 assign wire3166 = ( (~ ni30330)  &  (~ ng31566)  &  (~ ng31070)  &  wire34156 ) ;
 assign wire3167 = ( (~ ng31021)  &  (~ ng31710)  &  wire34188  &  wire34193 ) ;
 assign wire3170 = ( (~ ng31021)  &  (~ ni30330)  &  wire34120  &  wire34121 ) ;
 assign wire3171 = ( (~ ng31021)  &  ni31141  &  wire34126  &  wire34127 ) ;
 assign wire3172 = ( (~ ng31021)  &  ni31191  &  wire34132  &  wire34133 ) ;
 assign wire3173 = ( (~ ng31021)  &  ni31271  &  wire34138  &  wire34139 ) ;
 assign wire3174 = ( ni31106  &  (~ ng31021)  &  wire34144  &  wire34145 ) ;
 assign wire3175 = ( (~ ng31021)  &  ni31221  &  wire34150  &  wire34151 ) ;
 assign wire3176 = ( (~ ng30673)  &  ni31121  &  (~ ng31070)  &  wire34156 ) ;
 assign wire3177 = ( (~ ng31070)  &  wire34156  &  wire34160 ) ;
 assign wire3183 = ( wire34071  &  wire34072  &  wire34078  &  wire34079 ) ;
 assign wire3184 = ( wire34071  &  wire34072  &  wire34082  &  wire34083 ) ;
 assign wire3185 = ( (~ wire32354)  &  (~ wire32355)  &  wire34085  &  wire34086 ) ;
 assign wire3186 = ( (~ wire32354)  &  (~ wire32355)  &  wire34088  &  wire34089 ) ;
 assign wire3187 = ( (~ wire32354)  &  (~ wire32355)  &  wire34091  &  wire34092 ) ;
 assign wire3189 = ( (~ wire32354)  &  (~ wire32355)  &  wire34095 ) ;
 assign wire3190 = ( pg72  &  ng4322  &  wire28640  &  wire34062 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640  &  wire34062 ) ;
 assign wire3191 = ( pg72  &  ng4322  &  wire29233  &  wire34063 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233  &  wire34063 ) ;
 assign wire3192 = ( (~ ng4125)  &  ng4112  &  (~ ng11245)  &  wire34059 ) ;
 assign wire3203 = ( wire34008  &  wire34009 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire34009 ) ;
 assign wire3205 = ( (~ pg35)  &  ng2161 ) ;
 assign wire3209 = ( (~ pg35)  &  ng5462 ) ;
 assign wire3212 = ( (~ pg35)  &  ng5953 ) ;
 assign wire3215 = ( (~ pg35)  &  ng5607 ) ;
 assign wire3228 = ( (~ pg35)  &  ng2279 ) ;
 assign wire3229 = ( ng2735  &  ng2741  &  (~ ng17297)  &  wire33983 ) ;
 assign wire3230 = ( (~ ng2735)  &  wire33985 ) | ( (~ ng2741)  &  wire33985 ) | ( ng17297  &  wire33985 ) ;
 assign wire3234 = ( (~ pg35)  &  ng3929 ) ;
 assign wire3237 = ( (~ pg35)  &  ng6303 ) ;
 assign wire3240 = ( (~ pg35)  &  ng763 ) ;
 assign wire3253 = ( (~ pg35)  &  ng6617 ) ;
 assign wire3256 = ( (~ pg35)  &  ng6589 ) ;
 assign wire3257 = ( ng17405  &  (~ ng28799)  &  wire33956 ) | ( ng26737  &  (~ ng28799)  &  wire33956 ) ;
 assign wire3258 = ( pg35  &  ng2331  &  (~ ng17405)  &  (~ ng26737) ) ;
 assign wire3267 = ( wire7725  &  wire33931 ) | ( ng14367  &  wire28488  &  wire33931 ) ;
 assign wire3268 = ( wire7725  &  wire33934 ) | ( ng14367  &  wire28488  &  wire33934 ) ;
 assign wire3269 = ( wire7725  &  wire33936 ) | ( ng14367  &  wire28488  &  wire33936 ) ;
 assign wire3271 = ( (~ ng14367)  &  (~ wire7725)  &  wire33938 ) | ( (~ wire7725)  &  (~ wire28488)  &  wire33938 ) ;
 assign wire3272 = ( wire7725  &  wire33939 ) | ( ng14367  &  wire28488  &  wire33939 ) ;
 assign wire3274 = ( (~ pg35)  &  ng2485 ) ;
 assign wire3276 = ( pg35  &  (~ ng1193) ) | ( pg35  &  (~ ng969)  &  (~ ng1008) ) ;
 assign wire3278 = ( pg35  &  (~ ng1536) ) | ( pg35  &  (~ ng1312)  &  (~ ng1351) ) ;
 assign wire3281 = ( (~ pg35)  &  ng3913 ) ;
 assign wire3284 = ( (~ ng9755)  &  wire33922 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire33922 ) ;
 assign wire3285 = ( ng2084  &  ng26759  &  ng9755 ) | ( ng2084  &  ng14438  &  ng9755 ) ;
 assign wire3289 = ( (~ pg35)  &  ng5599 ) ;
 assign wire3292 = ( (~ pg35)  &  ng744 ) ;
 assign wire3295 = ( (~ pg35)  &  ng3602 ) ;
 assign wire3298 = ( (~ pg35)  &  ng2831 ) ;
 assign wire3304 = ( pg35  &  (~ ng4581)  &  ng4372 ) ;
 assign wire3307 = ( (~ pg35)  &  ng6235 ) ;
 assign wire3326 = ( (~ ng14367)  &  (~ wire6172)  &  wire33896 ) | ( (~ wire6172)  &  (~ wire30555)  &  wire33896 ) ;
 assign wire3327 = ( ng2185  &  wire6172 ) | ( ng2185  &  ng14367  &  wire30555 ) ;
 assign wire3336 = ( wire33887  &  wire33889 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire33889 ) ;
 assign wire3337 = ( (~ pg35)  &  ng2299 ) ;
 assign wire3343 = ( ng1772  &  (~ ng28761)  &  ng17317 ) | ( ng1772  &  (~ ng28761)  &  ng26694 ) ;
 assign wire3344 = ( pg35  &  ng1802  &  (~ ng17317)  &  (~ ng26694) ) ;
 assign wire3349 = ( (~ pg35)  &  ng2681 ) ;
 assign wire3350 = ( wire6319  &  wire33869 ) | ( ng14367  &  wire30342  &  wire33869 ) ;
 assign wire3351 = ( (~ ng14367)  &  (~ wire6319)  &  wire33870 ) | ( (~ wire6319)  &  (~ wire30342)  &  wire33870 ) ;
 assign wire3356 = ( (~ pg35)  &  ng3574 ) ;
 assign wire3367 = ( pg35  &  (~ ng626)  &  ng14708  &  wire33854 ) ;
 assign wire3368 = ( pg35  &  (~ ng632)  &  (~ ng14708)  &  wire33857 ) ;
 assign wire3369 = ( pg35  &  (~ ng626)  &  (~ ng14708)  &  wire33860 ) ;
 assign wire3370 = ( (~ pg35)  &  ng559 ) ;
 assign wire3376 = ( (~ pg35)  &  ng5591 ) ;
 assign wire3382 = ( wire29834  &  wire33832 ) | ( wire29835  &  wire33832 ) | ( wire29836  &  wire33832 ) ;
 assign wire3383 = ( wire29834  &  wire33834 ) | ( wire29835  &  wire33834 ) | ( wire29836  &  wire33834 ) ;
 assign wire3384 = ( pg35  &  ng4340  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire3385 = ( pg35  &  ng4340  &  ng4349  &  ng4358 ) ;
 assign wire3389 = ( (~ pg35)  &  ng5913 ) ;
 assign wire3393 = ( ng26793  &  ng9835  &  wire33803 ) | ( ng14506  &  ng9835  &  wire33803 ) ;
 assign wire3394 = ( ng26793  &  ng9835  &  wire33804 ) | ( ng14506  &  ng9835  &  wire33804 ) ;
 assign wire3395 = ( (~ ng9835)  &  wire33805 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire33805 ) ;
 assign wire3396 = ( (~ pg35)  &  ng2667 ) ;
 assign wire3399 = ( (~ pg35)  &  ng142 ) ;
 assign wire3402 = ( (~ pg35)  &  ng401 ) ;
 assign wire3407 = ( pg35  &  (~ ng990)  &  (~ ng979)  &  ng1008 ) ;
 assign wire3408 = ( ng979  &  ng969  &  (~ ng996) ) | ( ng990  &  (~ ng979)  &  ng969  &  ng996 ) ;
 assign wire3409 = ( (~ pg35)  &  ng969 ) ;
 assign wire3411 = ( wire30477  &  wire33781 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire33781 ) ;
 assign wire3412 = ( (~ pg35)  &  ng1890 ) ;
 assign wire3418 = ( (~ pg35)  &  ng604 ) ;
 assign wire3422 = ( (~ pg35)  &  ng4939 ) ;
 assign wire3426 = ( (~ pg35)  &  ng2652 ) ;
 assign wire3431 = ( wire33758  &  wire33760 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire33760 ) ;
 assign wire3432 = ( (~ pg35)  &  ng1736 ) ;
 assign wire3435 = ( (~ pg35)  &  ng3925 ) ;
 assign wire3442 = ( (~ pg35)  &  ng1917 ) ;
 assign wire3443 = ( (~ ng9649)  &  wire33743 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire33743 ) ;
 assign wire3444 = ( ng2241  &  ng9649  &  ng26703 ) | ( ng2241  &  ng9649  &  ng17321 ) ;
 assign wire3453 = ( (~ pg35)  &  ng5929 ) ;
 assign wire3456 = ( (~ pg35)  &  ng914 ) ;
 assign wire3462 = ( (~ pg35)  &  ng6271 ) ;
 assign wire3464 = ( (~ pg17604)  &  (~ pg13049)  &  ng10160  &  wire33726 ) ;
 assign wire3465 = ( wire6172  &  wire33703 ) | ( ng14367  &  wire30555  &  wire33703 ) ;
 assign wire3466 = ( wire6172  &  wire33706 ) | ( ng14367  &  wire30555  &  wire33706 ) ;
 assign wire3467 = ( wire6172  &  wire33708 ) | ( ng14367  &  wire30555  &  wire33708 ) ;
 assign wire3468 = ( wire6172  &  wire33709 ) | ( ng14367  &  wire30555  &  wire33709 ) ;
 assign wire3470 = ( (~ ng14367)  &  (~ wire6172)  &  wire33711 ) | ( (~ wire6172)  &  (~ wire30555)  &  wire33711 ) ;
 assign wire3471 = ( (~ pg35)  &  ng2217 ) ;
 assign wire3485 = ( (~ pg35)  &  ng4411 ) ;
 assign wire3492 = ( (~ pg35)  &  ng1825 ) ;
 assign wire3495 = ( (~ pg35)  &  ng5260 ) ;
 assign wire3497 = ( (~ ng11960)  &  wire33682 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire33682 ) ;
 assign wire3498 = ( (~ pg35)  &  ng2437 ) ;
 assign wire3501 = ( (~ pg35)  &  ng4785 ) ;
 assign wire3504 = ( wire33024  &  wire33670 ) | ( wire33025  &  wire33670 ) | ( wire33048  &  wire33670 ) ;
 assign wire3505 = ( (~ wire33024)  &  (~ wire33025)  &  (~ wire33048)  &  wire33672 ) ;
 assign wire3506 = ( (~ wire6966)  &  (~ wire6967)  &  (~ wire29216)  &  wire33673 ) ;
 assign wire3507 = ( (~ pg35)  &  ng3462 ) ;
 assign wire3521 = ( wire33659  &  wire33661 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33661 ) ;
 assign wire3522 = ( (~ pg35)  &  ng1616 ) ;
 assign wire3526 = ( pg35  &  pg12923  &  ng1395 ) ;
 assign wire3530 = ( (~ pg35)  &  ng4119 ) ;
 assign wire3533 = ( (~ pg35)  &  ng5551 ) ;
 assign wire3541 = ( (~ pg35)  &  ng5208 ) ;
 assign wire3545 = ( (~ pg35)  &  ng2051 ) ;
 assign wire3546 = ( wire5887  &  wire33620 ) | ( ng14367  &  wire31005  &  wire33620 ) ;
 assign wire3547 = ( wire5887  &  wire33623 ) | ( ng14367  &  wire31005  &  wire33623 ) ;
 assign wire3548 = ( wire5887  &  wire33625 ) | ( ng14367  &  wire31005  &  wire33625 ) ;
 assign wire3549 = ( wire5887  &  wire33626 ) | ( ng14367  &  wire31005  &  wire33626 ) ;
 assign wire3551 = ( (~ ng14367)  &  (~ wire5887)  &  wire33628 ) | ( (~ wire5887)  &  (~ wire31005)  &  wire33628 ) ;
 assign wire3553 = ( (~ pg35)  &  ng2619 ) ;
 assign wire3560 = ( (~ pg35)  &  ng2384 ) ;
 assign wire3562 = ( wire33608  &  wire33610 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire33610 ) ;
 assign wire3563 = ( (~ pg35)  &  ng1740 ) ;
 assign wire3565 = ( (~ pg17646)  &  (~ pg17739)  &  ng10185  &  wire33606 ) ;
 assign wire3571 = ( (~ pg35)  &  ng3546 ) ;
 assign wire3574 = ( (~ pg35)  &  ng590 ) ;
 assign wire3578 = ( (~ pg13895)  &  (~ pg14421)  &  ng8691  &  wire33585 ) ;
 assign wire3584 = ( ng26673  &  ng9586  &  wire33571 ) | ( ng9586  &  ng17292  &  wire33571 ) ;
 assign wire3585 = ( (~ ng9586)  &  wire33572 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33572 ) ;
 assign wire3594 = ( (~ ng14367)  &  (~ wire6172)  &  wire33563 ) | ( (~ wire6172)  &  (~ wire30555)  &  wire33563 ) ;
 assign wire3595 = ( wire6172  &  wire33564 ) | ( ng14367  &  wire30555  &  wire33564 ) ;
 assign wire3600 = ( (~ wire33551)  &  (~ wire33553)  &  wire33554 ) | ( (~ wire33552)  &  (~ wire33553)  &  wire33554 ) ;
 assign wire3601 = ( wire33553  &  wire33555 ) | ( wire33551  &  wire33552  &  wire33555 ) ;
 assign wire3607 = ( (~ ng11956)  &  wire33545 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire33545 ) ;
 assign wire3608 = ( (~ pg35)  &  ng2012 ) ;
 assign wire3616 = ( wire33536  &  wire33538 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33538 ) ;
 assign wire3617 = ( (~ pg35)  &  ng1604 ) ;
 assign wire3618 = ( ng34162  &  wire33533 ) | ( (~ wire31938)  &  wire33533 ) | ( wire31939  &  wire33533 ) ;
 assign wire3619 = ( (~ ng34162)  &  wire31938  &  (~ wire31939)  &  wire33534 ) ;
 assign wire3629 = ( (~ pg35)  &  ng5575 ) ;
 assign wire3632 = ( (~ pg35)  &  ng4801 ) ;
 assign wire3635 = ( (~ pg35)  &  ng5052 ) ;
 assign wire3642 = ( (~ pg35)  &  ng1018 ) ;
 assign wire3643 = ( (~ ng30583)  &  ng24411  &  (~ wire6408)  &  wire33510 ) ;
 assign wire3644 = ( (~ ng30583)  &  (~ ng24411)  &  (~ wire6408)  &  wire33512 ) ;
 assign wire3649 = ( (~ pg35)  &  ng6173 ) ;
 assign wire3653 = ( (~ pg35)  &  ng1720 ) ;
 assign wire3657 = ( (~ pg35)  &  ng3106 ) ;
 assign wire3658 = ( pg35  &  (~ ni24685) ) | ( pg35  &  wire29414 ) ;
 assign wire3659 = ( pg35  &  ng17657 ) | ( pg35  &  ng17700 ) ;
 assign wire3667 = ( (~ pg35)  &  ng6275 ) ;
 assign wire3676 = ( (~ pg35)  &  ng5571 ) ;
 assign wire3677 = ( (~ ng25917)  &  (~ wire4362)  &  (~ wire4669)  &  wire33472 ) ;
 assign wire3678 = ( ng25917  &  wire33473 ) | ( wire4362  &  wire33473 ) | ( wire4669  &  wire33473 ) ;
 assign wire3688 = ( (~ pg35)  &  ng291 ) ;
 assign wire3691 = ( (~ pg35)  &  ng3582 ) ;
 assign wire3693 = ( wire33455  &  wire33457 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire33457 ) ;
 assign wire3694 = ( (~ pg35)  &  ng2567 ) ;
 assign wire3695 = ( ng28504  &  wire33452 ) | ( (~ wire28813)  &  wire33452 ) | ( wire28814  &  wire33452 ) ;
 assign wire3696 = ( (~ ng28504)  &  wire28813  &  (~ wire28814)  &  wire33453 ) ;
 assign wire3704 = ( (~ ng13336)  &  (~ ng13846)  &  wire33428  &  wire33429 ) ;
 assign wire3705 = ( ng13336  &  (~ ng13846)  &  wire33432  &  wire33433 ) ;
 assign wire3712 = ( (~ pg35)  &  ng4653 ) ;
 assign wire3719 = ( (~ pg35)  &  ng5579 ) ;
 assign wire3720 = ( wire30977  &  wire33410 ) | ( wire30978  &  wire33410 ) | ( wire31001  &  wire33410 ) ;
 assign wire3721 = ( (~ wire30977)  &  (~ wire30978)  &  (~ wire31001)  &  wire33412 ) ;
 assign wire3722 = ( (~ wire7624)  &  (~ wire7625)  &  (~ wire28651)  &  wire33413 ) ;
 assign wire3723 = ( (~ pg35)  &  ng5120 ) ;
 assign wire3727 = ( (~ pg35)  &  ng2342 ) ;
 assign wire3729 = ( wire6172  &  wire33397 ) | ( ng14367  &  wire30555  &  wire33397 ) ;
 assign wire3730 = ( (~ ng14367)  &  (~ wire6172)  &  wire33398 ) | ( (~ wire6172)  &  (~ wire30555)  &  wire33398 ) ;
 assign wire3736 = ( (~ pg35)  &  ng6593 ) ;
 assign wire3746 = ( (~ ng9640)  &  wire33386 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire33386 ) ;
 assign wire3747 = ( (~ pg35)  &  ng1821 ) ;
 assign wire3752 = ( (~ pg35)  &  ng3203 ) ;
 assign wire3755 = ( ng9694  &  ng26725  &  wire33377 ) | ( ng9694  &  ng17401  &  wire33377 ) ;
 assign wire3756 = ( ng9694  &  ng26725  &  wire33378 ) | ( ng9694  &  ng17401  &  wire33378 ) ;
 assign wire3757 = ( (~ ng9694)  &  wire33379 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire33379 ) ;
 assign wire3758 = ( (~ pg35)  &  ng1974 ) ;
 assign wire3760 = ( wire33372  &  wire33374 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire33374 ) ;
 assign wire3761 = ( (~ pg35)  &  ng2433 ) ;
 assign wire3762 = ( (~ ng1129)  &  (~ ng13307)  &  ng13336  &  wire33366 ) | ( ng1129  &  (~ ng13307)  &  (~ ng13336)  &  wire33366 ) ;
 assign wire3763 = ( pg35  &  (~ ng1129)  &  ng1124  &  ng13336 ) | ( pg35  &  ng1129  &  ng1124  &  (~ ng13336) ) ;
 assign wire3768 = ( (~ ng9694)  &  wire33364 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire33364 ) ;
 assign wire3769 = ( ng1968  &  ng9694  &  ng26725 ) | ( ng1968  &  ng9694  &  ng17401 ) ;
 assign wire3771 = ( (~ ng9649)  &  wire33362 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire33362 ) ;
 assign wire3772 = ( ng2259  &  ng9649  &  ng26703 ) | ( ng2259  &  ng9649  &  ng17321 ) ;
 assign wire3780 = ( pg35  &  (~ ng1495)  &  ng1489 ) ;
 assign wire3782 = ( wire29834  &  wire33353 ) | ( wire29835  &  wire33353 ) | ( wire29836  &  wire33353 ) ;
 assign wire3786 = ( wire7030  &  wire33349 ) | ( ng14367  &  wire29111  &  wire33349 ) ;
 assign wire3787 = ( (~ ng14367)  &  (~ wire7030)  &  wire33350 ) | ( (~ wire7030)  &  (~ wire29111)  &  wire33350 ) ;
 assign wire3791 = ( (~ pg35)  &  ng5264 ) ;
 assign wire3801 = ( (~ wire7046)  &  (~ wire7047)  &  (~ wire29091)  &  wire33335 ) ;
 assign wire3802 = ( wire30659  &  wire33336 ) | ( wire30660  &  wire33336 ) | ( wire30683  &  wire33336 ) ;
 assign wire3804 = ( wire6655  &  wire33330 ) | ( ng14367  &  wire29571  &  wire33330 ) ;
 assign wire3805 = ( (~ ng14367)  &  (~ wire6655)  &  wire33331 ) | ( (~ wire6655)  &  (~ wire29571)  &  wire33331 ) ;
 assign wire3810 = ( (~ pg35)  &  ng4601 ) ;
 assign wire3816 = ( (~ pg35)  &  ng3566 ) ;
 assign wire3821 = ( pg35  &  (~ ng4581)  &  ng4372 ) ;
 assign wire3827 = ( (~ pg35)  &  ng2173 ) ;
 assign wire3828 = ( wire7257  &  wire33302 ) | ( ng14367  &  wire28834  &  wire33302 ) ;
 assign wire3829 = ( (~ ng14367)  &  (~ wire7257)  &  wire33303 ) | ( (~ wire7257)  &  (~ wire28834)  &  wire33303 ) ;
 assign wire3837 = ( ng817  &  (~ ng8806)  &  (~ ng14279)  &  wire33291 ) ;
 assign wire3838 = ( (~ ng817)  &  (~ ng14279)  &  wire33293 ) | ( ng8806  &  (~ ng14279)  &  wire33293 ) ;
 assign wire3845 = ( (~ pg35)  &  ng5941 ) ;
 assign wire3849 = ( (~ pg35)  &  ng2208 ) ;
 assign wire3853 = ( ng17405  &  ng9700  &  wire33273 ) | ( ng26737  &  ng9700  &  wire33273 ) ;
 assign wire3854 = ( ng17405  &  ng9700  &  wire33275 ) | ( ng26737  &  ng9700  &  wire33275 ) ;
 assign wire3855 = ( (~ ng9700)  &  wire33276 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire33276 ) ;
 assign wire3856 = ( (~ pg35)  &  ng2399 ) ;
 assign wire3860 = ( (~ pg35)  &  ng1802 ) ;
 assign wire3868 = ( (~ pg35)  &  ng5212 ) ;
 assign wire3874 = ( (~ pg35)  &  ng1221 ) ;
 assign wire3880 = ( (~ pg35)  &  ng6613 ) ;
 assign wire3883 = ( (~ pg35)  &  ng5945 ) ;
 assign wire3886 = ( (~ pg35)  &  ng153 ) ;
 assign wire3889 = ( (~ pg35)  &  ng3562 ) ;
 assign wire3892 = ( (~ pg35)  &  ng6621 ) ;
 assign wire3894 = ( pg116  &  pg35  &  ng4157 ) | ( pg114  &  pg35  &  (~ ng4157) ) ;
 assign wire3895 = ( (~ ng9762)  &  wire33238 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire33238 ) ;
 assign wire3897 = ( (~ pg35)  &  ng2514 ) ;
 assign wire3902 = ( (~ ng9755)  &  wire33234 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire33234 ) ;
 assign wire3903 = ( (~ pg35)  &  ng2089 ) ;
 assign wire3905 = ( (~ ng9586)  &  wire33231 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33231 ) ;
 assign wire3906 = ( (~ pg35)  &  ng1687 ) ;
 assign wire3910 = ( (~ pg73)  &  (~ pg72)  &  pg35  &  ng2988 ) ;
 assign wire3912 = ( (~ pg35)  &  ng4564 ) ;
 assign wire3915 = ( (~ pg35)  &  ng5595 ) ;
 assign wire3918 = ( (~ pg35)  &  ng5917 ) ;
 assign wire3921 = ( (~ pg35)  &  ng5961 ) ;
 assign wire3922 = ( (~ ng14367)  &  (~ wire6655)  &  wire33208 ) | ( (~ wire6655)  &  (~ wire29571)  &  wire33208 ) ;
 assign wire3924 = ( ng1894  &  wire6655 ) | ( ng1894  &  ng14367  &  wire29571 ) ;
 assign wire3926 = ( (~ pg17519)  &  (~ pg13039)  &  ng10124  &  wire33189 ) ;
 assign wire3927 = ( pg12238  &  (~ pg13039)  &  ng10124  &  wire33194 ) ;
 assign wire3928 = ( wire33199  &  wire33200 ) ;
 assign wire3929 = ( pg12238  &  (~ pg13039)  &  ng10124  &  wire33204 ) ;
 assign wire3932 = ( (~ pg35)  &  ng3953 ) ;
 assign wire3939 = ( (~ ng9700)  &  wire33181 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire33181 ) ;
 assign wire3940 = ( (~ pg35)  &  ng2380 ) ;
 assign wire3946 = ( (~ pg35)  &  ng5244 ) ;
 assign wire3952 = ( (~ pg35)  &  ng4349 ) ;
 assign wire3955 = ( (~ pg35)  &  ng5268 ) ;
 assign wire3958 = ( (~ pg35)  &  ng3610 ) ;
 assign wire3961 = ( (~ ng25233)  &  (~ wire29550)  &  (~ wire29551)  &  wire33161 ) ;
 assign wire3962 = ( pg35  &  (~ ng5046)  &  ng25233 ) ;
 assign wire3967 = ( (~ ng14367)  &  (~ wire6319)  &  wire33156 ) | ( (~ wire6319)  &  (~ wire30342)  &  wire33156 ) ;
 assign wire3969 = ( wire6319  &  wire33158 ) | ( ng14367  &  wire30342  &  wire33158 ) ;
 assign wire3974 = ( (~ pg35)  &  ng5148 ) ;
 assign wire3975 = ( ng26673  &  ng9586  &  wire33143 ) | ( ng9586  &  ng17292  &  wire33143 ) ;
 assign wire3976 = ( ng26673  &  ng9586  &  wire33145 ) | ( ng9586  &  ng17292  &  wire33145 ) ;
 assign wire3977 = ( (~ ng9586)  &  wire33146 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33146 ) ;
 assign wire3978 = ( (~ pg35)  &  ng1706 ) ;
 assign wire3979 = ( (~ ng9586)  &  wire33140 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire33140 ) ;
 assign wire3980 = ( ng1682  &  ng26673  &  ng9586 ) | ( ng1682  &  ng9586  &  ng17292 ) ;
 assign wire3984 = ( (~ pg35)  &  ng3554 ) ;
 assign wire3988 = ( (~ pg35)  &  ng5841 ) ;
 assign wire3991 = ( (~ pg35)  &  ng4116 ) ;
 assign wire3994 = ( (~ pg35)  &  ng6605 ) ;
 assign wire3998 = ( (~ pg35)  &  ng2795 ) ;
 assign wire4001 = ( (~ pg35)  &  ng5901 ) ;
 assign wire4003 = ( pg35  &  ng1263  &  (~ ng1270)  &  (~ ng25895) ) ;
 assign wire4007 = ( (~ pg35)  &  ng667 ) ;
 assign wire4011 = ( (~ ng9694)  &  wire33102 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire33102 ) ;
 assign wire4012 = ( ng1950  &  ng9694  &  ng26725 ) | ( ng1950  &  ng9694  &  ng17401 ) ;
 assign wire4016 = ( ng17317  &  ng9640  &  wire33096 ) | ( ng26694  &  ng9640  &  wire33096 ) ;
 assign wire4017 = ( ng17317  &  ng9640  &  wire33098 ) | ( ng26694  &  ng9640  &  wire33098 ) ;
 assign wire4018 = ( (~ ng9640)  &  wire33099 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire33099 ) ;
 assign wire4019 = ( (~ pg35)  &  ng1840 ) ;
 assign wire4025 = ( (~ pg35)  &  ng613 ) ;
 assign wire4034 = ( pg35  &  (~ ng5069)  &  ng5077  &  ng5084 ) ;
 assign wire4041 = ( (~ pg35)  &  ng3231 ) ;
 assign wire4044 = ( (~ pg35)  &  ng168 ) ;
 assign wire4045 = ( wire32138  &  wire33069 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire33069 ) ;
 assign wire4047 = ( (~ pg35)  &  ng2024 ) ;
 assign wire4050 = ( (~ pg35)  &  ng6247 ) ;
 assign wire4051 = ( wire5887  &  wire33061 ) | ( ng14367  &  wire31005  &  wire33061 ) ;
 assign wire4053 = ( (~ ng14367)  &  (~ wire5887)  &  wire33063 ) | ( (~ wire5887)  &  (~ wire31005)  &  wire33063 ) ;
 assign wire4064 = ( (~ pg35)  &  ng572 ) ;
 assign wire4068 = ( (~ wire6966)  &  (~ wire6967)  &  (~ wire29216)  &  wire32991 ) ;
 assign wire4069 = ( wire33024  &  wire33049 ) | ( wire33025  &  wire33049 ) | ( wire33048  &  wire33049 ) ;
 assign wire4094 = ( ng843  &  ng847  &  (~ ng8806)  &  wire32987 ) ;
 assign wire4095 = ( (~ ng843)  &  wire32989 ) | ( (~ ng847)  &  wire32989 ) | ( ng8806  &  wire32989 ) ;
 assign wire4099 = ( (~ pg35)  &  ng4054 ) ;
 assign wire4100 = ( (~ ng14708)  &  wire32978 ) | ( wire28793  &  wire32978 ) | ( (~ wire28794)  &  wire32978 ) ;
 assign wire4101 = ( ng14708  &  (~ wire28793)  &  wire28794  &  wire32979 ) ;
 assign wire4106 = ( ng29503  &  ng14438  &  ng27469  &  wire32969 ) ;
 assign wire4107 = ( ng29503  &  ng14438  &  ng27469  &  wire32971 ) ;
 assign wire4108 = ( (~ ng29503)  &  wire32972 ) | ( (~ ng14438)  &  wire32972 ) | ( (~ ng27469)  &  wire32972 ) ;
 assign wire4109 = ( (~ pg35)  &  ng1996 ) ;
 assign wire4112 = ( (~ pg35)  &  ng4659 ) ;
 assign wire4115 = ( (~ pg35)  &  ng1259 ) ;
 assign wire4118 = ( (~ pg35)  &  ng3352 ) ;
 assign wire4124 = ( (~ pg35)  &  ng2441 ) ;
 assign wire4127 = ( (~ pg35)  &  ng262 ) ;
 assign wire4133 = ( (~ pg35)  &  ng6295 ) ;
 assign wire4137 = ( (~ pg35)  &  ng2787 ) ;
 assign wire4144 = ( ng10756  &  wire28765  &  wire32928 ) | ( ng10756  &  wire28766  &  wire32928 ) ;
 assign wire4145 = ( (~ ng10756)  &  wire32929 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire32929 ) ;
 assign wire4154 = ( (~ pg35)  &  ng3538 ) ;
 assign wire4156 = ( pg35  &  ng2287  &  (~ ng17405)  &  (~ ng26737) ) ;
 assign wire4157 = ( (~ ng13378)  &  (~ ng13273)  &  wire32898  &  wire32899 ) ;
 assign wire4158 = ( ng13378  &  (~ ng13273)  &  wire32902  &  wire32903 ) ;
 assign wire4168 = ( (~ pg35)  &  ng739 ) ;
 assign wire4172 = ( (~ pg35)  &  ng1612 ) ;
 assign wire4175 = ( (~ pg35)  &  ng758 ) ;
 assign wire4176 = ( ng21012  &  (~ ng25851)  &  wire32879 ) | ( ng21012  &  (~ wire32672)  &  wire32879 ) ;
 assign wire4177 = ( (~ wire7248)  &  (~ wire7249)  &  (~ wire28843)  &  wire32881 ) ;
 assign wire4189 = ( (~ ng11978)  &  wire32875 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32875 ) ;
 assign wire4190 = ( (~ pg35)  &  ng2571 ) ;
 assign wire4191 = ( (~ ng14367)  &  (~ wire7257)  &  wire32869 ) | ( (~ wire7257)  &  (~ wire28834)  &  wire32869 ) ;
 assign wire4193 = ( wire7257  &  wire32871 ) | ( ng14367  &  wire28834  &  wire32871 ) ;
 assign wire4197 = ( (~ pg35)  &  ng6279 ) ;
 assign wire4199 = ( (~ ng14367)  &  (~ wire7041)  &  wire32863 ) | ( (~ wire7041)  &  (~ wire29097)  &  wire32863 ) ;
 assign wire4200 = ( ng1624  &  wire7041 ) | ( ng1624  &  ng14367  &  wire29097 ) ;
 assign wire4204 = ( (~ pg35)  &  ng146 ) ;
 assign wire4207 = ( (~ pg35)  &  ng3937 ) ;
 assign wire4210 = ( (~ pg35)  &  ng5703 ) ;
 assign wire4220 = ( wire32841  &  wire32843 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire32843 ) ;
 assign wire4221 = ( (~ pg35)  &  ng2295 ) ;
 assign wire4226 = ( (~ pg35)  &  ng5200 ) ;
 assign wire4227 = ( pg35  &  (~ ng1536)  &  wire7193 ) | ( pg35  &  (~ ng1536)  &  wire28903 ) ;
 assign wire4228 = ( (~ ng1542)  &  wire32832 ) | ( ng10918  &  wire32832 ) | ( (~ wire28896)  &  wire32832 ) ;
 assign wire4233 = ( ng29503  &  ng27395  &  ng17292  &  wire32823 ) ;
 assign wire4234 = ( ng29503  &  ng27395  &  ng17292  &  wire32825 ) ;
 assign wire4235 = ( (~ ng29503)  &  wire32826 ) | ( (~ ng27395)  &  wire32826 ) | ( (~ ng17292)  &  wire32826 ) ;
 assign wire4236 = ( (~ pg35)  &  ng1592 ) ;
 assign wire4242 = ( (~ pg35)  &  ng5196 ) ;
 assign wire4248 = ( (~ pg35)  &  ng1280 ) ;
 assign wire4253 = ( ng20875  &  (~ ng25851)  &  wire32802 ) | ( ng20875  &  (~ wire31986)  &  wire32802 ) ;
 assign wire4254 = ( (~ wire7351)  &  (~ wire7352)  &  (~ wire28734)  &  wire32804 ) ;
 assign wire4278 = ( ng26759  &  (~ ng28833)  &  wire32787 ) | ( ng14438  &  (~ ng28833)  &  wire32787 ) ;
 assign wire4279 = ( pg35  &  ng2040  &  (~ ng26759)  &  (~ ng14438) ) ;
 assign wire4283 = ( (~ pg35)  &  ng3207 ) ;
 assign wire4288 = ( (~ pg35)  &  ng3586 ) ;
 assign wire4291 = ( (~ pg35)  &  ng4664 ) ;
 assign wire4300 = ( (~ pg35)  &  ng3941 ) ;
 assign wire4303 = ( (~ pg35)  &  ng239 ) ;
 assign wire4306 = ( (~ pg35)  &  ng3703 ) ;
 assign wire4308 = ( ng2599  &  (~ ng28880)  &  ng26793 ) | ( ng2599  &  (~ ng28880)  &  ng14506 ) ;
 assign wire4309 = ( (~ pg35)  &  ng2599 ) ;
 assign wire4314 = ( (~ pg35)  &  ng6629 ) ;
 assign wire4315 = ( ng2759  &  ng2756  &  ng25317  &  wire32749 ) ;
 assign wire4316 = ( (~ ng2759)  &  wire32750 ) | ( (~ ng2756)  &  wire32750 ) | ( (~ ng25317)  &  wire32750 ) ;
 assign wire4319 = ( (~ ng9762)  &  wire32747 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire32747 ) ;
 assign wire4320 = ( ng2509  &  ng26770  &  ng9762 ) | ( ng2509  &  ng17424  &  ng9762 ) ;
 assign wire4332 = ( wire7030  &  wire32728 ) | ( ng14367  &  wire29111  &  wire32728 ) ;
 assign wire4333 = ( wire7030  &  wire32731 ) | ( ng14367  &  wire29111  &  wire32731 ) ;
 assign wire4334 = ( wire7030  &  wire32733 ) | ( ng14367  &  wire29111  &  wire32733 ) ;
 assign wire4335 = ( wire7030  &  wire32734 ) | ( ng14367  &  wire29111  &  wire32734 ) ;
 assign wire4336 = ( (~ ng14367)  &  (~ wire7030)  &  wire32735 ) | ( (~ wire7030)  &  (~ wire29111)  &  wire32735 ) ;
 assign wire4339 = ( (~ pg35)  &  ng2351 ) ;
 assign wire4343 = ( (~ pg35)  &  ng2227 ) ;
 assign wire4355 = ( (~ pg35)  &  ng626 ) ;
 assign wire4359 = ( pg35  &  (~ ng25917)  &  wire4362  &  (~ wire4669) ) ;
 assign wire4361 = ( (~ pg35)  &  ng1367 ) ;
 assign wire4362 = ( (~ ng1373)  &  (~ ng15748) ) ;
 assign wire4366 = ( (~ pg35)  &  ng5603 ) ;
 assign wire4367 = ( ng911  &  ng907  &  ng19063  &  wire32699 ) ;
 assign wire4368 = ( (~ ng911)  &  wire32700 ) | ( (~ ng907)  &  wire32700 ) | ( (~ ng19063)  &  wire32700 ) ;
 assign wire4378 = ( (~ pg35)  &  ng3961 ) ;
 assign wire4403 = ( (~ pg35)  &  ng6395 ) ;
 assign wire4404 = ( wire32668  &  wire32669 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire32669 ) ;
 assign wire4406 = ( (~ pg35)  &  ng1886 ) ;
 assign wire4414 = ( pg35  &  (~ ng714)  &  ng703  &  ng691 ) ;
 assign wire4415 = ( wire30802  &  (~ wire32625)  &  wire32661 ) | ( wire30803  &  (~ wire32625)  &  wire32661 ) ;
 assign wire4417 = ( (~ pg35)  &  ng79 ) ;
 assign wire4421 = ( (~ pg35)  &  ng2070 ) ;
 assign wire4429 = ( pg35  &  (~ ng1322)  &  ng1351  &  (~ ng1333) ) ;
 assign wire4430 = ( ng1322  &  ng1312  &  (~ ng1339) ) | ( (~ ng1322)  &  ng1312  &  ng1333  &  ng1339 ) ;
 assign wire4431 = ( (~ pg35)  &  ng1312 ) ;
 assign wire4439 = ( (~ pg35)  &  ng6283 ) ;
 assign wire4445 = ( (~ ng9762)  &  wire32636 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire32636 ) ;
 assign wire4446 = ( ng2527  &  ng26770  &  ng9762 ) | ( ng2527  &  ng17424  &  ng9762 ) ;
 assign wire4456 = ( ng26793  &  ng9835  &  wire32633 ) | ( ng14506  &  ng9835  &  wire32633 ) ;
 assign wire4457 = ( (~ ng9835)  &  wire32634 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32634 ) ;
 assign wire4462 = ( (~ pg35)  &  ng4961 ) ;
 assign wire4466 = ( wire32625  &  wire32626 ) | ( (~ wire30802)  &  (~ wire30803)  &  wire32626 ) ;
 assign wire4467 = ( (~ pg35)  &  ng691 ) ;
 assign wire4470 = ( (~ pg35)  &  ng812 ) ;
 assign wire4477 = ( ng31509  &  wire32616 ) | ( (~ wire30328)  &  wire32616 ) | ( wire30329  &  wire32616 ) ;
 assign wire4478 = ( (~ ng31509)  &  wire30328  &  (~ wire30329)  &  wire32617 ) ;
 assign wire4486 = ( (~ pg35)  &  ng225 ) ;
 assign wire4488 = ( wire31143  &  wire32610 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire32610 ) ;
 assign wire4489 = ( (~ pg35)  &  ng1620 ) ;
 assign wire4493 = ( pg35  &  ng2555  &  (~ ng26793)  &  (~ ng14506) ) ;
 assign wire4494 = ( (~ ng9835)  &  wire32602 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32602 ) ;
 assign wire4495 = ( ng2661  &  ng26793  &  ng9835 ) | ( ng2661  &  ng14506  &  ng9835 ) ;
 assign wire4499 = ( (~ pg35)  &  ng790 ) ;
 assign wire4505 = ( wire32594  &  wire32596 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire32596 ) ;
 assign wire4506 = ( (~ pg35)  &  ng2315 ) ;
 assign wire4509 = ( (~ pg35)  &  ng1542 ) ;
 assign wire4514 = ( (~ ng14367)  &  (~ wire5887)  &  wire32583 ) | ( (~ wire5887)  &  (~ wire31005)  &  wire32583 ) ;
 assign wire4515 = ( wire5887  &  wire32584 ) | ( ng14367  &  wire31005  &  wire32584 ) ;
 assign wire4517 = ( ng4087  &  ng4076  &  (~ ng13217)  &  wire32578 ) ;
 assign wire4518 = ( (~ ng4087)  &  wire32580 ) | ( (~ ng4076)  &  wire32580 ) | ( ng13217  &  wire32580 ) ;
 assign wire4525 = ( (~ pg35)  &  ng5949 ) ;
 assign wire4528 = ( (~ ng11937)  &  wire32571 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire32571 ) ;
 assign wire4530 = ( (~ pg35)  &  ng1878 ) ;
 assign wire4531 = ( wire29451  &  wire32565 ) | ( wire29452  &  wire32565 ) | ( wire29475  &  wire32565 ) ;
 assign wire4532 = ( (~ wire29451)  &  (~ wire29452)  &  (~ wire29475)  &  wire32567 ) ;
 assign wire4533 = ( (~ wire7351)  &  (~ wire7352)  &  (~ wire28734)  &  wire32568 ) ;
 assign wire4534 = ( (~ pg35)  &  ng5813 ) ;
 assign wire4537 = ( (~ pg35)  &  ng4818 ) ;
 assign wire4538 = ( ng10756  &  wire28765  &  wire32554 ) | ( ng10756  &  wire28766  &  wire32554 ) ;
 assign wire4539 = ( (~ ng10756)  &  wire32555 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire32555 ) ;
 assign wire4540 = ( ng10756  &  wire28765  &  wire32556 ) | ( ng10756  &  wire28766  &  wire32556 ) ;
 assign wire4541 = ( (~ pg35)  &  ng3827 ) ;
 assign wire4550 = ( (~ pg35)  &  ng1178 ) ;
 assign wire4570 = ( (~ pg35)  &  ng518 ) ;
 assign wire4574 = ( (~ pg35)  &  ng1648 ) ;
 assign wire4577 = ( (~ ng24875)  &  wire32526 ) | ( wire28810  &  wire32526 ) | ( (~ wire28811)  &  wire32526 ) ;
 assign wire4578 = ( ng24875  &  (~ wire28810)  &  wire28811  &  wire32527 ) ;
 assign wire4581 = ( wire32521  &  wire32523 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire32523 ) ;
 assign wire4582 = ( (~ pg35)  &  ng1752 ) ;
 assign wire4583 = ( ng26770  &  (~ ng28846)  &  wire32517 ) | ( ng17424  &  (~ ng28846)  &  wire32517 ) ;
 assign wire4584 = ( pg35  &  ng2465  &  (~ ng26770)  &  (~ ng17424) ) ;
 assign wire4590 = ( (~ ng4785)  &  (~ ng4709)  &  ng11261  &  wire32511 ) ;
 assign wire4595 = ( (~ pg35)  &  ng3490 ) ;
 assign wire4596 = ( ng4054  &  wire28765  &  wire32476 ) | ( ng4054  &  wire28766  &  wire32476 ) ;
 assign wire4598 = ( ng4054  &  wire28765  &  wire32482 ) | ( ng4054  &  wire28766  &  wire32482 ) ;
 assign wire4600 = ( (~ ng4975)  &  ng4899  &  ng11283  &  wire32486 ) ;
 assign wire4604 = ( (~ pg35)  &  ng4818 ) ;
 assign wire4608 = ( (~ pg35)  &  ng4760 ) ;
 assign wire4623 = ( (~ pg35)  &  ng617 ) ;
 assign wire4626 = ( (~ pg35)  &  ng3542 ) ;
 assign wire4630 = ( (~ pg35)  &  ng2775 ) ;
 assign wire4633 = ( (~ pg35)  &  ng4621 ) ;
 assign wire4652 = ( (~ ng13336)  &  (~ ng13260)  &  wire32408  &  wire32409 ) ;
 assign wire4653 = ( ng13336  &  (~ ng13260)  &  wire32412  &  wire32413 ) ;
 assign wire4659 = ( wire7041  &  wire32404 ) | ( ng14367  &  wire29097  &  wire32404 ) ;
 assign wire4660 = ( (~ ng14367)  &  (~ wire7041)  &  wire32405 ) | ( (~ wire7041)  &  (~ wire29097)  &  wire32405 ) ;
 assign wire4663 = ( (~ ng14367)  &  (~ wire6319)  &  wire32399 ) | ( (~ wire6319)  &  (~ wire30342)  &  wire32399 ) ;
 assign wire4664 = ( ng2028  &  wire6319 ) | ( ng2028  &  ng14367  &  wire30342 ) ;
 assign wire4669 = ( (~ ng1367)  &  (~ ng15748) ) ;
 assign wire4673 = ( (~ pg35)  &  ng3187 ) ;
 assign wire4676 = ( ng9694  &  ng26725  &  wire32388 ) | ( ng9694  &  ng17401  &  wire32388 ) ;
 assign wire4677 = ( (~ ng9694)  &  wire32389 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire32389 ) ;
 assign wire4681 = ( (~ pg35)  &  ng4145 ) ;
 assign wire4683 = ( (~ ng9649)  &  wire32383 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire32383 ) ;
 assign wire4684 = ( (~ pg35)  &  ng2246 ) ;
 assign wire4685 = ( (~ ng11320)  &  wire32377  &  wire32378  &  wire32379 ) ;
 assign wire4689 = ( (~ pg35)  &  ng6219 ) ;
 assign wire4692 = ( ng9649  &  ng26703  &  wire32363 ) | ( ng9649  &  ng17321  &  wire32363 ) ;
 assign wire4693 = ( (~ ng9649)  &  wire32364 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire32364 ) ;
 assign wire4708 = ( pg35  &  (~ ng896)  &  ng862 ) ;
 assign wire4711 = ( (~ ng9835)  &  wire32341 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32341 ) ;
 assign wire4712 = ( (~ pg35)  &  ng2648 ) ;
 assign wire4715 = ( (~ pg35)  &  ng4593 ) ;
 assign wire4721 = ( (~ ng9835)  &  wire32333 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32333 ) ;
 assign wire4722 = ( ng2643  &  ng26793  &  ng9835 ) | ( ng2643  &  ng14506  &  ng9835 ) ;
 assign wire4724 = ( (~ ng9700)  &  wire32331 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire32331 ) ;
 assign wire4725 = ( ng2375  &  ng17405  &  ng9700 ) | ( ng2375  &  ng26737  &  ng9700 ) ;
 assign wire4729 = ( (~ pg35)  &  ng3558 ) ;
 assign wire4736 = ( (~ pg35)  &  ng1691 ) ;
 assign wire4740 = ( (~ wire7248)  &  (~ wire7249)  &  (~ wire28843)  &  wire32316 ) ;
 assign wire4741 = ( wire32202  &  wire32317 ) | ( wire32203  &  wire32317 ) | ( wire32226  &  wire32317 ) ;
 assign wire4745 = ( (~ pg35)  &  ng6307 ) ;
 assign wire4749 = ( (~ pg35)  &  ng4572 ) ;
 assign wire4757 = ( (~ pg35)  &  ng59 ) ;
 assign wire4759 = ( wire32251  &  wire32252  &  wire32253 ) ;
 assign wire4760 = ( (~ ng4688)  &  (~ ng4776)  &  wire32259  &  wire32260 ) ;
 assign wire4761 = ( (~ ng4688)  &  (~ ng4776)  &  wire32266  &  wire32267 ) ;
 assign wire4764 = ( wire32269  &  wire32288  &  wire32289 ) | ( wire32270  &  wire32288  &  wire32289 ) ;
 assign wire4765 = ( (~ ng4681)  &  (~ ng4646)  &  ng11261  &  wire32293 ) ;
 assign wire4766 = ( pg35  &  (~ ng4826)  &  ng4688 ) ;
 assign wire4767 = ( pg35  &  ng4674  &  (~ ng4821) ) ;
 assign wire4768 = ( pg35  &  ng128  &  ng4646 ) ;
 assign wire4769 = ( pg35  &  ng4831  &  ng4681 ) ;
 assign wire4783 = ( (~ pg35)  &  ng4049 ) ;
 assign wire4794 = ( (~ pg35)  &  ng5248 ) ;
 assign wire4795 = ( wire32202  &  wire32228 ) | ( wire32203  &  wire32228 ) | ( wire32226  &  wire32228 ) ;
 assign wire4796 = ( (~ wire32202)  &  (~ wire32203)  &  (~ wire32226)  &  wire32230 ) ;
 assign wire4797 = ( (~ wire7248)  &  (~ wire7249)  &  (~ wire28843)  &  wire32231 ) ;
 assign wire4798 = ( (~ pg35)  &  ng6159 ) ;
 assign wire4826 = ( pg73  &  (~ pg72)  &  pg35  &  ng255 ) ;
 assign wire4827 = ( (~ pg73)  &  (~ pg72)  &  pg35  &  ng269 ) ;
 assign wire4828 = ( (~ pg73)  &  pg72  &  pg35  &  ng262 ) ;
 assign wire4834 = ( (~ pg16627)  &  (~ pg16656)  &  ng8728  &  wire32151 ) ;
 assign wire4836 = ( pg35  &  ng1996  &  (~ ng26759)  &  (~ ng14438) ) ;
 assign wire4839 = ( (~ pg35)  &  ng3179 ) ;
 assign wire4842 = ( pg73  &  pg35  &  ng4581 ) | ( pg72  &  pg35  &  ng4581 ) ;
 assign wire4843 = ( pg35  &  ng4578  &  ng4581 ) ;
 assign wire4857 = ( (~ pg35)  &  ng5897 ) ;
 assign wire4860 = ( (~ pg35)  &  ng3239 ) ;
 assign wire4861 = ( pg35  &  (~ ng1193)  &  wire7709 ) | ( pg35  &  (~ ng1193)  &  wire28519 ) ;
 assign wire4863 = ( (~ ng1199)  &  wire32117 ) | ( ng10893  &  wire32117 ) | ( (~ wire29901)  &  wire32117 ) ;
 assign wire4870 = ( (~ pg35)  &  ng3211 ) ;
 assign wire4873 = ( (~ pg35)  &  ng1559 ) ;
 assign wire4878 = ( wire6319  &  wire32101 ) | ( ng14367  &  wire30342  &  wire32101 ) ;
 assign wire4879 = ( (~ ng14367)  &  (~ wire6319)  &  wire32102 ) | ( (~ wire6319)  &  (~ wire30342)  &  wire32102 ) ;
 assign wire4882 = ( wire32095  &  wire32097 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32097 ) ;
 assign wire4883 = ( (~ pg35)  &  ng2563 ) ;
 assign wire4884 = ( (~ ng9755)  &  wire32093 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire32093 ) ;
 assign wire4885 = ( ng2102  &  ng26759  &  ng9755 ) | ( ng2102  &  ng14438  &  ng9755 ) ;
 assign wire4888 = ( wire32085  &  wire32087 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire32087 ) ;
 assign wire4889 = ( (~ pg35)  &  ng2004 ) ;
 assign wire4892 = ( (~ pg35)  &  ng3909 ) ;
 assign wire4893 = ( wire32078  &  wire32079 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32079 ) ;
 assign wire4895 = ( (~ pg35)  &  ng2583 ) ;
 assign wire4899 = ( (~ pg35)  &  ng2547 ) ;
 assign wire4903 = ( (~ pg35)  &  ng2518 ) ;
 assign wire4906 = ( (~ pg35)  &  ng4608 ) ;
 assign wire4908 = ( wire7725  &  wire32056 ) | ( ng14367  &  wire28488  &  wire32056 ) ;
 assign wire4909 = ( (~ ng14367)  &  (~ wire7725)  &  wire32057 ) | ( (~ wire7725)  &  (~ wire28488)  &  wire32057 ) ;
 assign wire4912 = ( pg35  &  ng854  &  ng11326 ) ;
 assign wire4913 = ( (~ ng691)  &  (~ ng417)  &  (~ ng13657)  &  wire32035 ) ;
 assign wire4914 = ( (~ ng691)  &  (~ ng417)  &  (~ ng13657)  &  wire32039 ) ;
 assign wire4915 = ( (~ ng691)  &  (~ ng417)  &  ng13657  &  wire32043 ) ;
 assign wire4916 = ( (~ ng691)  &  (~ ng417)  &  ng13657  &  wire32047 ) ;
 assign wire4929 = ( (~ ng14367)  &  (~ wire7030)  &  wire32019 ) | ( (~ wire7030)  &  (~ wire29111)  &  wire32019 ) ;
 assign wire4930 = ( wire7030  &  wire32020 ) | ( ng14367  &  wire29111  &  wire32020 ) ;
 assign wire4934 = ( (~ pg35)  &  ng5188 ) ;
 assign wire4937 = ( (~ pg35)  &  ng5543 ) ;
 assign wire4941 = ( (~ pg35)  &  ng4749 ) ;
 assign wire4944 = ( (~ ng164)  &  ng23042  &  wire32003 ) | ( ng23042  &  (~ wire28708)  &  wire32003 ) ;
 assign wire4945 = ( ng164  &  ng23042  &  wire28708  &  wire32005 ) ;
 assign wire4952 = ( (~ pg35)  &  ng6243 ) ;
 assign wire4955 = ( (~ pg35)  &  ng6255 ) ;
 assign wire4958 = ( (~ pg35)  &  ng6049 ) ;
 assign wire4972 = ( (~ pg35)  &  ng3881 ) ;
 assign wire4982 = ( (~ pg35)  &  ng4688 ) ;
 assign wire4988 = ( (~ pg35)  &  ng5905 ) ;
 assign wire4993 = ( (~ pg35)  &  ng4633 ) ;
 assign wire4999 = ( (~ pg35)  &  ng1783 ) ;
 assign wire5002 = ( (~ pg35)  &  ng807 ) ;
 assign wire5005 = ( (~ pg35)  &  ng5615 ) ;
 assign wire5008 = ( (~ pg35)  &  ng3235 ) ;
 assign wire5011 = ( (~ pg35)  &  ng3199 ) ;
 assign wire5018 = ( (~ pg35)  &  ng6653 ) ;
 assign wire5021 = ( (~ pg35)  &  ng4878 ) ;
 assign wire5024 = ( (~ pg35)  &  ng1564 ) ;
 assign wire5036 = ( (~ pg35)  &  ng1959 ) ;
 assign wire5064 = ( (~ pg35)  &  ng5925 ) ;
 assign wire5067 = ( (~ pg35)  &  ng1193 ) ;
 assign wire5070 = ( (~ pg35)  &  ng4991 ) ;
 assign wire5076 = ( (~ ng4785)  &  ng4709  &  ng11261  &  wire31870 ) ;
 assign wire5079 = ( (~ pg35)  &  ng5921 ) ;
 assign wire5082 = ( (~ pg35)  &  ng3606 ) ;
 assign wire5085 = ( (~ pg35)  &  ng3259 ) ;
 assign wire5089 = ( (~ pg35)  &  ng6519 ) ;
 assign wire5092 = ( (~ pg35)  &  ng3530 ) ;
 assign wire5098 = ( (~ pg35)  &  ng6625 ) ;
 assign wire5103 = ( (~ pg35)  &  ng3949 ) ;
 assign wire5107 = ( (~ pg35)  &  ng2610 ) ;
 assign wire5120 = ( (~ pg35)  &  ng6609 ) ;
 assign wire5123 = ( (~ pg35)  &  ng5555 ) ;
 assign wire5128 = ( (~ pg35)  &  ng3215 ) ;
 assign wire5132 = ( (~ pg35)  &  ng5827 ) ;
 assign wire5136 = ( (~ pg35)  &  ng1668 ) ;
 assign wire5142 = ( (~ pg35)  &  ng2815 ) ;
 assign wire5145 = ( (~ pg35)  &  ng3171 ) ;
 assign wire5148 = ( ng11676  &  wire31784 ) | ( (~ wire28525)  &  wire31784 ) | ( (~ wire28526)  &  wire31784 ) ;
 assign wire5149 = ( ng732  &  (~ ng11676)  &  wire28525  &  wire28526 ) ;
 assign wire5156 = ( (~ pg35)  &  ng5611 ) ;
 assign wire5164 = ( wire31770  &  wire31772 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire31772 ) ;
 assign wire5165 = ( (~ pg35)  &  ng1870 ) ;
 assign wire5176 = ( ng20887  &  (~ ni27429)  &  wire31759 ) | ( ng20887  &  (~ wire31757)  &  wire31759 ) ;
 assign wire5177 = ( (~ wire7137)  &  (~ wire7138)  &  (~ wire28996)  &  wire31761 ) ;
 assign wire5183 = ( (~ pg35)  &  ng5204 ) ;
 assign wire5196 = ( (~ ng4975)  &  (~ ng4899)  &  ng11283  &  wire31744 ) ;
 assign wire5201 = ( ng2070  &  (~ ng2040)  &  ng26314  &  wire30377 ) ;
 assign wire5202 = ( (~ ng2599)  &  ng2629  &  ng26314  &  wire29061 ) ;
 assign wire5203 = ( ng1668  &  (~ ng1636)  &  ng26314  &  wire30283 ) ;
 assign wire5204 = ( ng2495  &  (~ ng2465)  &  ng26314  &  wire29272 ) ;
 assign wire5205 = ( ng1936  &  (~ ng1906)  &  ng26314  &  wire30276 ) ;
 assign wire5206 = ( (~ ng1772)  &  ng1802  &  ng26314  &  wire28687 ) ;
 assign wire5207 = ( (~ ng2197)  &  ng2227  &  ng26314  &  wire30616 ) ;
 assign wire5208 = ( ng2361  &  (~ ng2331)  &  ng26314  &  wire30356 ) ;
 assign wire5209 = ( ng1263  &  ng1270  &  (~ ng25895)  &  wire31719 ) ;
 assign wire5210 = ( (~ ng1263)  &  wire31720 ) | ( (~ ng1270)  &  wire31720 ) | ( ng25895  &  wire31720 ) ;
 assign wire5214 = ( (~ pg35)  &  ng5236 ) ;
 assign wire5217 = ( (~ pg35)  &  ng4311 ) ;
 assign wire5231 = ( (~ pg35)  &  ng6267 ) ;
 assign wire5251 = ( (~ pg35)  &  ng562 ) ;
 assign wire5258 = ( ng23586  &  (~ wire29550)  &  (~ wire29551)  &  wire31679 ) ;
 assign wire5259 = ( (~ ng5037)  &  (~ ng17217)  &  wire31681 ) | ( ng5037  &  (~ ng14317)  &  wire31681 ) ;
 assign wire5273 = ( (~ pg35)  &  ng513 ) ;
 assign wire5276 = ( pg35  &  ng1146  &  (~ ng1152) ) ;
 assign wire5279 = ( (~ pg35)  &  ng5873 ) ;
 assign wire5289 = ( (~ pg35)  &  ng150 ) ;
 assign wire5294 = ( (~ pg35)  &  ng872 ) ;
 assign wire5299 = ( ng979  &  ng996  &  ng11846  &  wire31634 ) | ( (~ ng979)  &  (~ ng996)  &  ng11846  &  wire31634 ) ;
 assign wire5302 = ( pg35  &  (~ ng990)  &  (~ ng979)  &  ng969 ) ;
 assign wire5304 = ( pg35  &  ng1728  &  (~ ng17317)  &  (~ ng26694) ) ;
 assign wire5308 = ( ng4375  &  wire31622 ) | ( ng4411  &  wire31622 ) | ( (~ wire29326)  &  wire31622 ) ;
 assign wire5309 = ( pg35  &  wire29325  &  wire29326  &  wire30770 ) ;
 assign wire5310 = ( (~ pg35)  &  ng4388 ) ;
 assign wire5315 = ( wire31615  &  wire31617 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire31617 ) ;
 assign wire5316 = ( (~ pg35)  &  ng1756 ) ;
 assign wire5319 = ( (~ pg35)  &  ng582 ) ;
 assign wire5322 = ( (~ pg35)  &  ng5559 ) ;
 assign wire5338 = ( (~ pg35)  &  ng4704 ) ;
 assign wire5342 = ( (~ pg35)  &  ng3125 ) ;
 assign wire5357 = ( (~ wire6832)  &  (~ wire6833)  &  (~ wire29346)  &  wire31574 ) ;
 assign wire5358 = ( wire30848  &  wire31575 ) | ( wire30849  &  wire31575 ) | ( wire30872  &  wire31575 ) ;
 assign wire5361 = ( wire31570  &  wire31572 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire31572 ) ;
 assign wire5362 = ( (~ pg35)  &  ng2445 ) ;
 assign wire5365 = ( pg35  &  (~ ng1322)  &  ng1345  &  (~ ng1333) ) ;
 assign wire5366 = ( pg35  &  (~ ng1345)  &  (~ ng7601)  &  (~ ng15748) ) ;
 assign wire5370 = ( (~ pg35)  &  ng1041 ) ;
 assign wire5372 = ( (~ ng11916)  &  wire31560 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire31560 ) ;
 assign wire5373 = ( (~ pg35)  &  ng2169 ) ;
 assign wire5376 = ( (~ pg35)  &  ng699 ) ;
 assign wire5390 = ( ng2197  &  ng26703  &  (~ ng28768) ) | ( ng2197  &  ng17321  &  (~ ng28768) ) ;
 assign wire5391 = ( (~ pg35)  &  ng2197 ) ;
 assign wire5394 = ( (~ pg35)  &  ng4843 ) ;
 assign wire5397 = ( (~ pg35)  &  ng5216 ) ;
 assign wire5406 = ( pg35  &  (~ pg8291)  &  ng209 ) | ( pg35  &  ng209  &  (~ ng218) ) ;
 assign wire5407 = ( (~ pg35)  &  ng191 ) ;
 assign wire5412 = ( (~ pg35)  &  ng3933 ) ;
 assign wire5419 = ( (~ pg35)  &  ng5587 ) ;
 assign wire5427 = ( wire29614  &  wire31514 ) | ( wire29615  &  wire31514 ) | ( wire29638  &  wire31514 ) ;
 assign wire5428 = ( (~ pg35)  &  ng3965 ) ;
 assign wire5430 = ( wire7041  &  wire31509 ) | ( ng14367  &  wire29097  &  wire31509 ) ;
 assign wire5431 = ( (~ ng14367)  &  (~ wire7041)  &  wire31510 ) | ( (~ wire7041)  &  (~ wire29097)  &  wire31510 ) ;
 assign wire5438 = ( ng925  &  ng918  &  (~ ng25888)  &  wire31505 ) ;
 assign wire5451 = ( (~ pg35)  &  ng5240 ) ;
 assign wire5456 = ( (~ pg35)  &  ng3873 ) ;
 assign wire5462 = ( (~ pg35)  &  ng5252 ) ;
 assign wire5463 = ( ng26770  &  ng9762  &  wire31488 ) | ( ng17424  &  ng9762  &  wire31488 ) ;
 assign wire5464 = ( ng26770  &  ng9762  &  wire31490 ) | ( ng17424  &  ng9762  &  wire31490 ) ;
 assign wire5465 = ( (~ ng9762)  &  wire31491 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire31491 ) ;
 assign wire5466 = ( (~ pg35)  &  ng2533 ) ;
 assign wire5469 = ( (~ pg35)  &  ng3889 ) ;
 assign wire5475 = ( (~ pg35)  &  ng5889 ) ;
 assign wire5476 = ( pg35  &  (~ ng4145)  &  (~ ng4253) ) | ( pg35  &  ng4253  &  (~ ng4164) ) ;
 assign wire5483 = ( (~ pg35)  &  ng5495 ) ;
 assign wire5487 = ( (~ pg35)  &  ng2250 ) ;
 assign wire5490 = ( (~ pg35)  &  ng1384 ) ;
 assign wire5491 = ( ng1351  &  (~ ng1384) ) ;
 assign wire5502 = ( (~ pg35)  &  ng671 ) ;
 assign wire5503 = ( wire6655  &  wire31447 ) | ( ng14367  &  wire29571  &  wire31447 ) ;
 assign wire5505 = ( (~ ng14367)  &  (~ wire6655)  &  wire31450 ) | ( (~ wire6655)  &  (~ wire29571)  &  wire31450 ) ;
 assign wire5512 = ( ng21024  &  (~ ni27429)  &  wire31437 ) | ( ng21024  &  (~ wire31435)  &  wire31437 ) ;
 assign wire5513 = ( (~ wire6966)  &  (~ wire6967)  &  (~ wire29216)  &  wire31439 ) ;
 assign wire5523 = ( (~ pg35)  &  ng2307 ) ;
 assign wire5524 = ( ng2331  &  ng17405  &  (~ ng28799) ) | ( ng2331  &  ng26737  &  (~ ng28799) ) ;
 assign wire5525 = ( pg35  &  ng2361  &  (~ ng17405)  &  (~ ng26737) ) ;
 assign wire5533 = ( (~ ng9694)  &  wire31415 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire31415 ) ;
 assign wire5534 = ( (~ pg35)  &  ng1955 ) ;
 assign wire5542 = ( pg35  &  ng2421  &  (~ ng26770)  &  (~ ng17424) ) ;
 assign wire5551 = ( (~ pg35)  &  ng4854 ) ;
 assign wire5552 = ( ng17317  &  ng9640  &  wire31391 ) | ( ng26694  &  ng9640  &  wire31391 ) ;
 assign wire5553 = ( (~ ng9640)  &  wire31392 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire31392 ) ;
 assign wire5555 = ( wire7041  &  wire31385 ) | ( ng14367  &  wire29097  &  wire31385 ) ;
 assign wire5557 = ( (~ ng14367)  &  (~ wire7041)  &  wire31388 ) | ( (~ wire7041)  &  (~ wire29097)  &  wire31388 ) ;
 assign wire5573 = ( (~ pg35)  &  ng2476 ) ;
 assign wire5574 = ( wire6172  &  wire31351 ) | ( ng14367  &  wire30555  &  wire31351 ) ;
 assign wire5576 = ( (~ ng14367)  &  (~ wire6172)  &  wire31354 ) | ( (~ wire6172)  &  (~ wire30555)  &  wire31354 ) ;
 assign wire5580 = ( (~ pg35)  &  ng3598 ) ;
 assign wire5586 = ( (~ pg35)  &  ng2093 ) ;
 assign wire5589 = ( (~ pg35)  &  ng6581 ) ;
 assign wire5593 = ( pg35  &  (~ ng4785)  &  ng28336  &  (~ ng13464) ) ;
 assign wire5595 = ( (~ pg35)  &  ng4776 ) ;
 assign wire5597 = ( pg35  &  (~ ng5073)  &  ng5077 ) ;
 assign wire5600 = ( (~ wire7284)  &  wire28543  &  wire31322 ) | ( (~ wire7284)  &  wire28544  &  wire31322 ) ;
 assign wire5601 = ( wire7284  &  wire31324 ) | ( (~ wire28543)  &  (~ wire28544)  &  wire31324 ) ;
 assign wire5603 = ( (~ pg35)  &  ng2771 ) ;
 assign wire5619 = ( (~ pg35)  &  ng4983 ) ;
 assign wire5623 = ( (~ pg35)  &  ng2361 ) ;
 assign wire5627 = ( wire6655  &  wire31281 ) | ( ng14367  &  wire29571  &  wire31281 ) ;
 assign wire5628 = ( (~ ng14367)  &  (~ wire6655)  &  wire31282 ) | ( (~ wire6655)  &  (~ wire29571)  &  wire31282 ) ;
 assign wire5632 = ( ng26725  &  (~ ng28789)  &  wire31275 ) | ( ng17401  &  (~ ng28789)  &  wire31275 ) ;
 assign wire5633 = ( pg35  &  ng1906  &  (~ ng26725)  &  (~ ng17401) ) ;
 assign wire5638 = ( pg35  &  ng4141  &  (~ ng2841) ) | ( pg35  &  (~ ng2841)  &  ng4082 ) ;
 assign wire5641 = ( pg35  &  (~ ng2841)  &  ng4093 ) ;
 assign wire5642 = ( pg35  &  (~ ng2841)  &  ng4064 ) | ( pg35  &  (~ ng2841)  &  ng4057 ) ;
 assign wire5643 = ( pg35  &  (~ ng4087)  &  (~ ng2841) ) ;
 assign wire5644 = ( (~ pg35)  &  ng4125 ) ;
 assign wire5645 = ( ng817  &  (~ ng8806)  &  wire31254 ) ;
 assign wire5648 = ( pg35  &  ng703  &  (~ ng847) ) | ( pg35  &  ng703  &  ng8806 ) ;
 assign wire5649 = ( (~ pg35)  &  ng847 ) ;
 assign wire5650 = ( (~ ng9640)  &  wire31250 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire31250 ) ;
 assign wire5651 = ( ng1834  &  ng17317  &  ng9640 ) | ( ng1834  &  ng26694  &  ng9640 ) ;
 assign wire5653 = ( pg35  &  (~ pg11678)  &  ng542 ) | ( pg35  &  ng542  &  ng736 ) ;
 assign wire5654 = ( pg35  &  (~ pg11678)  &  (~ ng691) ) | ( pg35  &  (~ ng691)  &  ng736 ) ;
 assign wire5661 = ( (~ pg35)  &  ng6227 ) ;
 assign wire5663 = ( wire5887  &  wire31240 ) | ( ng14367  &  wire31005  &  wire31240 ) ;
 assign wire5664 = ( (~ ng14367)  &  (~ wire5887)  &  wire31241 ) | ( (~ wire5887)  &  (~ wire31005)  &  wire31241 ) ;
 assign wire5669 = ( (~ pg35)  &  ng2575 ) ;
 assign wire5671 = ( (~ ng11939)  &  wire31230 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire31230 ) ;
 assign wire5672 = ( (~ pg35)  &  ng2303 ) ;
 assign wire5690 = ( (~ ng9586)  &  wire31217 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire31217 ) ;
 assign wire5691 = ( ng1700  &  ng26673  &  ng9586 ) | ( ng1700  &  ng9586  &  ng17292 ) ;
 assign wire5693 = ( (~ ng4108)  &  wire31213 ) | ( (~ ng4098)  &  wire31213 ) | ( (~ ng22654)  &  wire31213 ) ;
 assign wire5694 = ( ng4108  &  ng4098  &  ng22654  &  wire31214 ) ;
 assign wire5697 = ( (~ ng25911)  &  (~ wire7650)  &  (~ wire7652)  &  wire31210 ) ;
 assign wire5698 = ( ng25911  &  wire31211 ) | ( wire7650  &  wire31211 ) | ( wire7652  &  wire31211 ) ;
 assign wire5702 = ( (~ pg35)  &  ng837 ) ;
 assign wire5705 = ( (~ pg35)  &  ng3590 ) ;
 assign wire5712 = ( wire7725  &  wire31194 ) | ( ng14367  &  wire28488  &  wire31194 ) ;
 assign wire5713 = ( (~ ng14367)  &  (~ wire7725)  &  wire31195 ) | ( (~ wire7725)  &  (~ wire28488)  &  wire31195 ) ;
 assign wire5718 = ( ng26759  &  ng9755  &  wire31190 ) | ( ng14438  &  ng9755  &  wire31190 ) ;
 assign wire5719 = ( (~ ng9755)  &  wire31191 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire31191 ) ;
 assign wire5727 = ( (~ pg35)  &  ng4443 ) ;
 assign wire5730 = ( (~ pg35)  &  ng5232 ) ;
 assign wire5734 = ( (~ pg35)  &  ng6154 ) ;
 assign wire5737 = ( (~ pg35)  &  ng4340 ) ;
 assign wire5740 = ( (~ pg35)  &  ng246 ) ;
 assign wire5747 = ( (~ ng11915)  &  wire31159 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire31159 ) ;
 assign wire5748 = ( (~ pg35)  &  ng1744 ) ;
 assign wire5755 = ( (~ pg35)  &  ng3893 ) ;
 assign wire5759 = ( (~ pg35)  &  ng2495 ) ;
 assign wire5766 = ( pg35  &  ng1592  &  (~ ng26673)  &  (~ ng17292) ) ;
 assign wire5769 = ( (~ pg35)  &  ng405 ) ;
 assign wire5773 = ( ng29503  &  ng27440  &  ng17401  &  wire31131 ) ;
 assign wire5774 = ( ng29503  &  ng27440  &  ng17401  &  wire31133 ) ;
 assign wire5775 = ( (~ ng29503)  &  wire31134 ) | ( (~ ng27440)  &  wire31134 ) | ( (~ ng17401)  &  wire31134 ) ;
 assign wire5776 = ( (~ pg35)  &  ng1862 ) ;
 assign wire5782 = ( (~ pg35)  &  ng6641 ) ;
 assign wire5783 = ( (~ ng1256)  &  wire31123 ) | ( (~ ng1252)  &  wire31123 ) | ( (~ ng19140)  &  wire31123 ) ;
 assign wire5785 = ( (~ pg35)  &  ng1256 ) ;
 assign wire5788 = ( (~ pg35)  &  ng6251 ) ;
 assign wire5797 = ( (~ pg35)  &  ng5933 ) ;
 assign wire5800 = ( (~ pg35)  &  ng3921 ) ;
 assign wire5803 = ( ng20682  &  (~ ng25851)  &  wire31107 ) | ( ng20682  &  (~ wire30578)  &  wire31107 ) ;
 assign wire5804 = ( (~ wire7624)  &  (~ wire7625)  &  (~ wire28651)  &  wire31109 ) ;
 assign wire5809 = ( (~ pg35)  &  ng3476 ) ;
 assign wire5811 = ( pg35  &  ng2153  &  (~ ng26703)  &  (~ ng17321) ) ;
 assign wire5814 = ( (~ pg35)  &  ng311 ) ;
 assign wire5819 = ( ng4785  &  ng4709  &  ng11261  &  wire31084 ) ;
 assign wire5821 = ( (~ ng10756)  &  wire31070 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire31070 ) ;
 assign wire5822 = ( ng3821  &  ng10756  &  wire28765 ) | ( ng3821  &  ng10756  &  wire28766 ) ;
 assign wire5827 = ( (~ pg35)  &  ng4950 ) ;
 assign wire5831 = ( (~ pg35)  &  ng5808 ) ;
 assign wire5834 = ( (~ pg35)  &  ng232 ) ;
 assign wire5835 = ( ng29503  &  ng27494  &  ng14506  &  wire31050 ) ;
 assign wire5836 = ( ng29503  &  ng27494  &  ng14506  &  wire31052 ) ;
 assign wire5837 = ( (~ ng29503)  &  wire31053 ) | ( (~ ng27494)  &  wire31053 ) | ( (~ ng14506)  &  wire31053 ) ;
 assign wire5838 = ( (~ pg35)  &  ng2555 ) ;
 assign wire5847 = ( (~ pg35)  &  ng1036 ) ;
 assign wire5848 = ( (~ ng1041)  &  ng1008 ) ;
 assign wire5856 = ( wire7030  &  wire31030 ) | ( ng14367  &  wire29111  &  wire31030 ) ;
 assign wire5859 = ( (~ ng14367)  &  (~ wire7030)  &  wire31033 ) | ( (~ wire7030)  &  (~ wire29111)  &  wire31033 ) ;
 assign wire5866 = ( (~ pg35)  &  ng3550 ) ;
 assign wire5868 = ( (~ ng14367)  &  (~ wire7030)  &  wire31023 ) | ( (~ wire7030)  &  (~ wire29111)  &  wire31023 ) ;
 assign wire5869 = ( ng2319  &  wire7030 ) | ( ng2319  &  ng14367  &  wire29111 ) ;
 assign wire5878 = ( (~ pg35)  &  ng3139 ) ;
 assign wire5883 = ( (~ ng14367)  &  (~ wire5887)  &  wire31008 ) | ( (~ wire5887)  &  (~ wire31005)  &  wire31008 ) ;
 assign wire5884 = ( ng2587  &  wire5887 ) | ( ng2587  &  ng14367  &  wire31005 ) ;
 assign wire5887 = ( ng2715  &  ng2724  &  ng2719 ) | ( ng2715  &  ng2729  &  ng2719 ) ;
 assign wire5888 = ( wire30977  &  wire31002 ) | ( wire30978  &  wire31002 ) | ( wire31001  &  wire31002 ) ;
 assign wire5889 = ( (~ wire7624)  &  (~ wire7625)  &  (~ wire28651)  &  wire31003 ) ;
 assign wire5925 = ( wire6319  &  wire30926 ) | ( ng14367  &  wire30342  &  wire30926 ) ;
 assign wire5926 = ( wire6319  &  wire30929 ) | ( ng14367  &  wire30342  &  wire30929 ) ;
 assign wire5927 = ( wire6319  &  wire30931 ) | ( ng14367  &  wire30342  &  wire30931 ) ;
 assign wire5928 = ( wire6319  &  wire30932 ) | ( ng14367  &  wire30342  &  wire30932 ) ;
 assign wire5929 = ( (~ ng14367)  &  (~ wire6319)  &  wire30933 ) | ( (~ wire6319)  &  (~ wire30342)  &  wire30933 ) ;
 assign wire5931 = ( (~ pg35)  &  ng2060 ) ;
 assign wire5941 = ( (~ pg35)  &  ng3841 ) ;
 assign wire5942 = ( ng23978  &  wire30914 ) | ( (~ wire28796)  &  wire30914 ) | ( wire28801  &  wire30914 ) ;
 assign wire5943 = ( (~ ng23978)  &  wire28796  &  (~ wire28801)  &  wire30915 ) ;
 assign wire5948 = ( (~ pg35)  &  ng2122 ) ;
 assign wire5952 = ( (~ pg35)  &  ng1882 ) ;
 assign wire5955 = ( (~ pg35)  &  ng6573 ) ;
 assign wire5959 = ( (~ pg35)  &  ng1854 ) ;
 assign wire5963 = ( ng26703  &  (~ ng28768)  &  wire30888 ) | ( ng17321  &  (~ ng28768)  &  wire30888 ) ;
 assign wire5964 = ( pg35  &  ng2197  &  (~ ng26703)  &  (~ ng17321) ) ;
 assign wire5968 = ( (~ ng28739)  &  ng26673  &  wire30881 ) | ( (~ ng28739)  &  ng17292  &  wire30881 ) ;
 assign wire5969 = ( pg35  &  ng1636  &  (~ ng26673)  &  (~ ng17292) ) ;
 assign wire5979 = ( wire30848  &  wire30874 ) | ( wire30849  &  wire30874 ) | ( wire30872  &  wire30874 ) ;
 assign wire5980 = ( (~ wire30848)  &  (~ wire30849)  &  (~ wire30872)  &  wire30876 ) ;
 assign wire5981 = ( (~ wire6832)  &  (~ wire6833)  &  (~ wire29346)  &  wire30877 ) ;
 assign wire5982 = ( (~ pg35)  &  ng5467 ) ;
 assign wire6009 = ( ng8806  &  wire30809 ) | ( (~ ng11185)  &  wire30809 ) | ( (~ wire30776)  &  wire30809 ) ;
 assign wire6010 = ( (~ ng8806)  &  ng11185  &  wire30776  &  wire30810 ) ;
 assign wire6011 = ( (~ ng8806)  &  ng11185  &  wire30776  &  wire30811 ) ;
 assign wire6012 = ( (~ pg35)  &  ng728 ) ;
 assign wire6015 = ( (~ pg35)  &  ng676 ) ;
 assign wire6028 = ( ng4375  &  wire30769 ) | ( ng4411  &  wire30769 ) | ( (~ wire29326)  &  wire30769 ) ;
 assign wire6029 = ( pg35  &  wire29325  &  wire29326  &  wire30770 ) ;
 assign wire6033 = ( (~ pg35)  &  ng1811 ) ;
 assign wire6036 = ( (~ pg35)  &  ng599 ) ;
 assign wire6042 = ( (~ pg35)  &  ng4975 ) ;
 assign wire6047 = ( (~ pg35)  &  ng6741 ) ;
 assign wire6048 = ( ng925  &  ng918  &  (~ ng25888)  &  wire30742 ) ;
 assign wire6049 = ( (~ ng925)  &  wire30743 ) | ( (~ ng918)  &  wire30743 ) | ( ng25888  &  wire30743 ) ;
 assign wire6055 = ( (~ ng14367)  &  (~ wire7725)  &  wire30733 ) | ( (~ wire7725)  &  (~ wire28488)  &  wire30733 ) ;
 assign wire6057 = ( wire7725  &  wire30735 ) | ( ng14367  &  wire28488  &  wire30735 ) ;
 assign wire6064 = ( ng4975  &  ng4899  &  ng11283  &  wire30728 ) ;
 assign wire6067 = ( (~ pg35)  &  ng6637 ) ;
 assign wire6068 = ( ng26770  &  ng9762  &  wire30709 ) | ( ng17424  &  ng9762  &  wire30709 ) ;
 assign wire6069 = ( (~ ng9762)  &  wire30710 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire30710 ) ;
 assign wire6093 = ( (~ wire30659)  &  (~ wire30660)  &  (~ wire30683)  &  wire30685 ) ;
 assign wire6094 = ( wire30659  &  wire30687 ) | ( wire30660  &  wire30687 ) | ( wire30683  &  wire30687 ) ;
 assign wire6095 = ( (~ wire7046)  &  (~ wire7047)  &  (~ wire29091)  &  wire30688 ) ;
 assign wire6096 = ( (~ pg35)  &  ng6505 ) ;
 assign wire6125 = ( ng29503  &  ng27421  &  ng17321  &  wire30619 ) ;
 assign wire6126 = ( ng29503  &  ng27421  &  ng17321  &  wire30621 ) ;
 assign wire6127 = ( (~ ng29503)  &  wire30622 ) | ( (~ ng27421)  &  wire30622 ) | ( (~ ng17321)  &  wire30622 ) ;
 assign wire6128 = ( (~ pg35)  &  ng2153 ) ;
 assign wire6133 = ( ng4785  &  (~ ng4709)  &  ng11261  &  wire30609 ) ;
 assign wire6148 = ( (~ pg35)  &  ng255 ) ;
 assign wire6151 = ( (~ pg35)  &  ng5357 ) ;
 assign wire6157 = ( (~ pg35)  &  ng6263 ) ;
 assign wire6160 = ( (~ pg35)  &  ng5033 ) ;
 assign wire6163 = ( (~ pg35)  &  ng6291 ) ;
 assign wire6167 = ( (~ pg35)  &  ng6187 ) ;
 assign wire6172 = ( (~ ng2715)  &  ng2724  &  (~ ng2719) ) | ( (~ ng2715)  &  ng2729  &  (~ ng2719) ) ;
 assign wire6173 = ( wire30497  &  wire30498  &  wire30499 ) ;
 assign wire6174 = ( (~ ng4983)  &  (~ ng4878)  &  wire30505  &  wire30506 ) ;
 assign wire6175 = ( (~ ng4983)  &  (~ ng4878)  &  wire30512  &  wire30513 ) ;
 assign wire6178 = ( wire30515  &  wire30534  &  wire30535 ) | ( wire30516  &  wire30534  &  wire30535 ) ;
 assign wire6179 = ( (~ ng4871)  &  (~ ng4836)  &  ng11283  &  wire30539 ) ;
 assign wire6180 = ( pg35  &  ng4836  &  ng5011 ) ;
 assign wire6181 = ( pg35  &  ng4871  &  ng3684 ) ;
 assign wire6182 = ( pg35  &  (~ ng4035)  &  ng4878 ) ;
 assign wire6183 = ( pg35  &  (~ ng3333)  &  ng4864 ) ;
 assign wire6197 = ( (~ pg35)  &  ng3522 ) ;
 assign wire6205 = ( pg35  &  ng1862  &  (~ ng26725)  &  (~ ng17401) ) ;
 assign wire6208 = ( (~ pg35)  &  ng5256 ) ;
 assign wire6211 = ( (~ pg35)  &  ng3227 ) ;
 assign wire6217 = ( (~ pg35)  &  ng3195 ) ;
 assign wire6223 = ( (~ pg35)  &  ng3255 ) ;
 assign wire6236 = ( (~ pg35)  &  ng3247 ) ;
 assign wire6237 = ( ng29503  &  ng17424  &  ng27474  &  wire30441 ) ;
 assign wire6238 = ( ng29503  &  ng17424  &  ng27474  &  wire30443 ) ;
 assign wire6239 = ( (~ ng29503)  &  wire30444 ) | ( (~ ng17424)  &  wire30444 ) | ( (~ ng27474)  &  wire30444 ) ;
 assign wire6240 = ( (~ pg35)  &  ng2421 ) ;
 assign wire6245 = ( (~ pg35)  &  ng3243 ) ;
 assign wire6248 = ( (~ pg35)  &  ng5957 ) ;
 assign wire6251 = ( (~ pg35)  &  ng6645 ) ;
 assign wire6254 = ( (~ pg35)  &  ng3191 ) ;
 assign wire6260 = ( (~ pg35)  &  ng1521 ) ;
 assign wire6269 = ( wire7041  &  wire30399 ) | ( ng14367  &  wire29097  &  wire30399 ) ;
 assign wire6270 = ( wire7041  &  wire30402 ) | ( ng14367  &  wire29097  &  wire30402 ) ;
 assign wire6271 = ( wire7041  &  wire30404 ) | ( ng14367  &  wire29097  &  wire30404 ) ;
 assign wire6273 = ( wire7041  &  wire30406 ) | ( ng14367  &  wire29097  &  wire30406 ) ;
 assign wire6274 = ( (~ ng14367)  &  (~ wire7041)  &  wire30407 ) | ( (~ wire7041)  &  (~ wire29097)  &  wire30407 ) ;
 assign wire6276 = ( (~ pg35)  &  ng1657 ) ;
 assign wire6277 = ( ng17405  &  ng9700  &  wire30394 ) | ( ng26737  &  ng9700  &  wire30394 ) ;
 assign wire6278 = ( (~ ng9700)  &  wire30395 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire30395 ) ;
 assign wire6281 = ( wire30390  &  wire30392 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire30392 ) ;
 assign wire6282 = ( (~ pg35)  &  ng2449 ) ;
 assign wire6283 = ( pg35  &  ng4473  &  (~ ng4462) ) ;
 assign wire6293 = ( (~ pg35)  &  ng5567 ) ;
 assign wire6294 = ( ng2040  &  ng26759  &  (~ ng28833) ) | ( ng2040  &  ng14438  &  (~ ng28833) ) ;
 assign wire6295 = ( pg35  &  ng2070  &  (~ ng26759)  &  (~ ng14438) ) ;
 assign wire6300 = ( (~ pg35)  &  ng6500 ) ;
 assign wire6301 = ( (~ ni27429)  &  ng20751  &  wire30367 ) | ( ng20751  &  (~ wire30365)  &  wire30367 ) ;
 assign wire6302 = ( (~ wire7046)  &  (~ wire7047)  &  (~ wire29091)  &  wire30369 ) ;
 assign wire6304 = ( ng29503  &  ng27445  &  ng17405  &  wire30359 ) ;
 assign wire6305 = ( ng29503  &  ng27445  &  ng17405  &  wire30361 ) ;
 assign wire6306 = ( (~ ng29503)  &  wire30362 ) | ( (~ ng27445)  &  wire30362 ) | ( (~ ng17405)  &  wire30362 ) ;
 assign wire6307 = ( (~ pg35)  &  ng2287 ) ;
 assign wire6317 = ( (~ pg35)  &  ng2016 ) ;
 assign wire6319 = ( ng2715  &  ng2724  &  ng2719 ) | ( ng2715  &  ng2729  &  ng2719 ) ;
 assign wire6323 = ( (~ pg35)  &  ng4643 ) ;
 assign wire6324 = ( (~ ng33851)  &  wire30334 ) | ( wire30331  &  wire30334 ) | ( (~ wire30332)  &  wire30334 ) ;
 assign wire6325 = ( ng33851  &  (~ wire30331)  &  wire30332  &  wire30335 ) ;
 assign wire6329 = ( (~ pg35)  &  ng772 ) ;
 assign wire6330 = ( wire6655  &  wire30307 ) | ( ng14367  &  wire29571  &  wire30307 ) ;
 assign wire6331 = ( wire6655  &  wire30310 ) | ( ng14367  &  wire29571  &  wire30310 ) ;
 assign wire6332 = ( wire6655  &  wire30312 ) | ( ng14367  &  wire29571  &  wire30312 ) ;
 assign wire6333 = ( wire6655  &  wire30313 ) | ( ng14367  &  wire29571  &  wire30313 ) ;
 assign wire6335 = ( (~ ng14367)  &  (~ wire6655)  &  wire30316 ) | ( (~ wire6655)  &  (~ wire29571)  &  wire30316 ) ;
 assign wire6336 = ( (~ pg35)  &  ng1926 ) ;
 assign wire6341 = ( ng1263  &  ng1270  &  (~ ng25895)  &  wire30300 ) ;
 assign wire6348 = ( (~ pg35)  &  ng822 ) ;
 assign wire6361 = ( ng1636  &  (~ ng28739)  &  ng26673 ) | ( ng1636  &  (~ ng28739)  &  ng17292 ) ;
 assign wire6362 = ( (~ pg35)  &  ng1636 ) ;
 assign wire6363 = ( ng1906  &  ng26725  &  (~ ng28789) ) | ( ng1906  &  ng17401  &  (~ ng28789) ) ;
 assign wire6364 = ( pg35  &  ng1936  &  (~ ng26725)  &  (~ ng17401) ) ;
 assign wire6368 = ( (~ pg35)  &  ng5220 ) ;
 assign wire6373 = ( ng4975  &  (~ ng4899)  &  ng11283  &  wire30265 ) ;
 assign wire6389 = ( wire30249  &  wire30251 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire30251 ) ;
 assign wire6390 = ( (~ pg35)  &  ng2311 ) ;
 assign wire6395 = ( ng1256  &  (~ ng1252)  &  ng22862 ) | ( ng1256  &  ng22862  &  (~ ng19140) ) ;
 assign wire6396 = ( pg35  &  (~ ng1256)  &  ng1252  &  ng19140 ) ;
 assign wire6398 = ( (~ ng1312)  &  (~ ng1351)  &  (~ ng13242)  &  wire30241 ) ;
 assign wire6407 = ( (~ pg35)  &  ng4332 ) ;
 assign wire6408 = ( (~ ng10511)  &  (~ ng8347)  &  (~ wire28475)  &  wire29918 ) ;
 assign wire6415 = ( (~ pg35)  &  ng6533 ) ;
 assign wire6421 = ( (~ pg35)  &  ng6299 ) ;
 assign wire6424 = ( (~ pg35)  &  ng1199 ) ;
 assign wire6436 = ( (~ pg35)  &  ng2827 ) ;
 assign wire6442 = ( (~ ng13378)  &  (~ ng13861)  &  wire29858  &  wire29859 ) ;
 assign wire6443 = ( ng13378  &  (~ ng13861)  &  wire29862  &  wire29863 ) ;
 assign wire6450 = ( (~ pg35)  &  ng3223 ) ;
 assign wire6451 = ( (~ pg35)  &  ng2834 ) ;
 assign wire6474 = ( pg35  &  (~ ng4340) ) | ( pg35  &  (~ ng4349) ) | ( pg35  &  (~ ng4358) ) ;
 assign wire6475 = ( pg35  &  (~ wire29834)  &  (~ wire29835)  &  (~ wire29836) ) ;
 assign wire6476 = ( pg35  &  (~ ng4633) ) | ( pg35  &  ng4639 ) | ( pg35  &  (~ ng4621) ) ;
 assign wire6482 = ( (~ pg135)  &  (~ ng4584)  &  ng4608  &  (~ ng4593) ) ;
 assign wire6486 = ( (~ pg35)  &  ng2783 ) ;
 assign wire6491 = ( (~ pg35)  &  ng5937 ) ;
 assign wire6494 = ( (~ pg35)  &  ng3578 ) ;
 assign wire6500 = ( (~ pg35)  &  ng785 ) ;
 assign wire6503 = ( (~ pg17722)  &  pg17778  &  ng10224  &  wire29780 ) ;
 assign wire6504 = ( (~ pg17722)  &  (~ pg17688)  &  ng10224  &  wire29785 ) ;
 assign wire6514 = ( (~ pg35)  &  ng5115 ) ;
 assign wire6515 = ( (~ ng9640)  &  wire29758 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire29758 ) ;
 assign wire6516 = ( ng1816  &  ng17317  &  ng9640 ) | ( ng1816  &  ng26694  &  ng9640 ) ;
 assign wire6520 = ( (~ pg35)  &  ng1216 ) ;
 assign wire6524 = ( (~ pg35)  &  ng5481 ) ;
 assign wire6527 = ( (~ pg35)  &  ng6565 ) ;
 assign wire6532 = ( (~ pg35)  &  ng6649 ) ;
 assign wire6539 = ( (~ pg35)  &  ng4771 ) ;
 assign wire6542 = ( (~ pg35)  &  ng3901 ) ;
 assign wire6544 = ( wire29723  &  wire29725 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire29725 ) ;
 assign wire6545 = ( (~ pg35)  &  ng2579 ) ;
 assign wire6548 = ( (~ ng32212)  &  wire29720 ) | ( wire28816  &  wire29720 ) | ( (~ wire29718)  &  wire29720 ) ;
 assign wire6549 = ( ng32212  &  (~ wire28816)  &  wire29718  &  wire29721 ) ;
 assign wire6552 = ( wire29714  &  wire29716 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire29716 ) ;
 assign wire6553 = ( (~ pg35)  &  ng2429 ) ;
 assign wire6561 = ( (~ ng837)  &  ng703  &  ng847  &  (~ ng8806) ) ;
 assign wire6565 = ( (~ pg35)  &  ng5909 ) ;
 assign wire6571 = ( pg35  &  (~ ng1002)  &  (~ ng15737)  &  (~ ng7567) ) ;
 assign wire6572 = ( pg35  &  (~ ng990)  &  (~ ng979)  &  ng1002 ) ;
 assign wire6576 = ( (~ pg35)  &  ng5224 ) ;
 assign wire6588 = ( (~ ng969)  &  (~ ng1008)  &  (~ ng13211)  &  wire29679 ) ;
 assign wire6592 = ( (~ pg35)  &  ng294 ) ;
 assign wire6595 = ( (~ pg35)  &  ng4112 ) ;
 assign wire6598 = ( (~ pg35)  &  ng4628 ) ;
 assign wire6604 = ( (~ pg35)  &  ng3251 ) ;
 assign wire6612 = ( (~ pg35)  &  ng5527 ) ;
 assign wire6614 = ( wire29646  &  wire29648 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire29648 ) ;
 assign wire6615 = ( (~ pg35)  &  ng1600 ) ;
 assign wire6619 = ( (~ wire29614)  &  (~ wire29615)  &  (~ wire29638)  &  wire29640 ) ;
 assign wire6620 = ( wire29614  &  wire29642 ) | ( wire29615  &  wire29642 ) | ( wire29638  &  wire29642 ) ;
 assign wire6622 = ( (~ pg35)  &  ng3813 ) ;
 assign wire6653 = ( (~ pg35)  &  ng1988 ) ;
 assign wire6655 = ( (~ ng2715)  &  ng2724  &  ng2719 ) | ( (~ ng2715)  &  ng2729  &  ng2719 ) ;
 assign wire6660 = ( (~ pg35)  &  ng5046 ) ;
 assign wire6663 = ( (~ pg35)  &  ng5547 ) ;
 assign wire6665 = ( wire29559  &  wire29561 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire29561 ) ;
 assign wire6666 = ( (~ pg35)  &  ng2020 ) ;
 assign wire6669 = ( (~ pg35)  &  ng504 ) ;
 assign wire6674 = ( ng7567  &  wire29542 ) | ( (~ ng1002)  &  (~ ng15737)  &  wire29542 ) ;
 assign wire6675 = ( (~ pg35)  &  ng1002 ) ;
 assign wire6678 = ( (~ pg35)  &  ng3945 ) ;
 assign wire6686 = ( (~ ng28444)  &  wire29526 ) | ( wire28561  &  wire29526 ) | ( (~ wire28562)  &  wire29526 ) ;
 assign wire6687 = ( ng28444  &  (~ wire28561)  &  wire28562  &  wire29527 ) ;
 assign wire6690 = ( (~ ng4443)  &  (~ ng4452)  &  wire29521  &  wire29523 ) ;
 assign wire6691 = ( (~ pg35)  &  ng4438 ) ;
 assign wire6694 = ( (~ pg35)  &  ng5535 ) ;
 assign wire6695 = ( ng26759  &  ng9755  &  wire29510 ) | ( ng14438  &  ng9755  &  wire29510 ) ;
 assign wire6696 = ( ng26759  &  ng9755  &  wire29511 ) | ( ng14438  &  ng9755  &  wire29511 ) ;
 assign wire6697 = ( (~ ng9755)  &  wire29512 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire29512 ) ;
 assign wire6698 = ( (~ pg35)  &  ng2108 ) ;
 assign wire6699 = ( ng24688  &  wire28661  &  wire29489 ) ;
 assign wire6700 = ( ng24688  &  wire29491  &  wire29493 ) ;
 assign wire6701 = ( ng24688  &  wire29495  &  wire29496 ) ;
 assign wire6702 = ( ng24688  &  wire28694  &  wire29497 ) ;
 assign wire6703 = ( ng24688  &  wire29499  &  wire29500 ) ;
 assign wire6704 = ( ng24688  &  ng10887  &  wire29502 ) ;
 assign wire6705 = ( ng24688  &  ng10823  &  wire29192 ) ;
 assign wire6706 = ( ng24688  &  ng10874  &  wire28470 ) ;
 assign wire6709 = ( (~ pg35)  &  ng832 ) ;
 assign wire6714 = ( (~ pg35)  &  ng5881 ) ;
 assign wire6715 = ( wire29451  &  wire29476 ) | ( wire29452  &  wire29476 ) | ( wire29475  &  wire29476 ) ;
 assign wire6716 = ( (~ wire7351)  &  (~ wire7352)  &  (~ wire28734)  &  wire29477 ) ;
 assign wire6743 = ( (~ pg35)  &  ng4375 ) ;
 assign wire6763 = ( (~ ng9700)  &  wire29408 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire29408 ) ;
 assign wire6764 = ( ng2393  &  ng17405  &  ng9700 ) | ( ng2393  &  ng26737  &  ng9700 ) ;
 assign wire6770 = ( ng2689  &  (~ ng2697)  &  ng2704 ) ;
 assign wire6777 = ( (~ pg35)  &  ng6239 ) ;
 assign wire6781 = ( ng499  &  ng691 ) | ( ng518  &  ng691 ) ;
 assign wire6784 = ( ng411  &  (~ ng691) ) ;
 assign wire6789 = ( (~ ng287)  &  ng23204  &  wire29391 ) | ( (~ ng283)  &  ng23204  &  wire29391 ) ;
 assign wire6790 = ( ng287  &  ng283  &  ng23204  &  wire29393 ) ;
 assign wire6804 = ( (~ pg73)  &  (~ pg72)  &  (~ ng4575)  &  ng4581 ) ;
 assign wire6805 = ( (~ ng4552)  &  (~ ng4581) ) ;
 assign wire6808 = ( pg73  &  pg35  &  ng4581 ) | ( pg72  &  pg35  &  ng4581 ) ;
 assign wire6809 = ( pg35  &  ng4572  &  ng4581 ) ;
 assign wire6816 = ( (~ ng10909)  &  (~ ng13336)  &  wire29362  &  wire29363 ) ;
 assign wire6817 = ( (~ ng10909)  &  ng13336  &  wire29366  &  wire29367 ) ;
 assign wire6823 = ( (~ pg73)  &  (~ pg72)  &  pg35  &  ng2988 ) ;
 assign wire6825 = ( (~ pg35)  &  ng4492 ) ;
 assign wire6826 = ( (~ pg73)  &  (~ pg72)  &  ng4581  &  (~ ng59) ) ;
 assign wire6827 = ( (~ ng4512)  &  (~ ng4581) ) ;
 assign wire6828 = ( ng20739  &  (~ ng25851)  &  wire29350 ) | ( ng20739  &  (~ wire29348)  &  wire29350 ) ;
 assign wire6829 = ( (~ wire6832)  &  (~ wire6833)  &  (~ wire29346)  &  wire29352 ) ;
 assign wire6832 = ( ng4801  &  ng4674 ) | ( ng4674  &  ng4793 ) | ( ng4674  &  (~ ng4776) ) ;
 assign wire6833 = ( ng4674  &  (~ ng4653) ) | ( ng4674  &  (~ ng4669) ) | ( ng4674  &  (~ ng4659) ) ;
 assign wire6838 = ( pg124  &  pg35  &  ng4146 ) | ( pg120  &  pg35  &  (~ ng4146) ) ;
 assign wire6842 = ( pg35  &  ng4388  &  (~ ng4430) ) ;
 assign wire6843 = ( pg35  &  ng4401  &  (~ ng4434) ) ;
 assign wire6844 = ( pg35  &  (~ ng4401)  &  ng4434 ) ;
 assign wire6847 = ( pg35  &  (~ ng4975)  &  ng28349  &  (~ ng13486) ) ;
 assign wire6849 = ( (~ pg35)  &  ng4966 ) ;
 assign wire6852 = ( (~ pg35)  &  ng3594 ) ;
 assign wire6872 = ( (~ pg35)  &  ng5893 ) ;
 assign wire6890 = ( (~ pg35)  &  ng4849 ) ;
 assign wire6899 = ( (~ pg35)  &  ng5228 ) ;
 assign wire6904 = ( (~ pg35)  &  ng5563 ) ;
 assign wire6905 = ( ng2465  &  ng26770  &  (~ ng28846) ) | ( ng2465  &  ng17424  &  (~ ng28846) ) ;
 assign wire6906 = ( pg35  &  ng2495  &  (~ ng26770)  &  (~ ng17424) ) ;
 assign wire6912 = ( ng2689  &  ng2697  &  (~ ng2704) ) ;
 assign wire6915 = ( (~ ng11893)  &  wire29266 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire29266 ) ;
 assign wire6916 = ( (~ pg35)  &  ng1608 ) ;
 assign wire6925 = ( (~ ng2145)  &  (~ ng2138)  &  ng2130 ) ;
 assign wire6933 = ( (~ pg35)  &  ng2629 ) ;
 assign wire6946 = ( pg72  &  ng4322  &  wire28640  &  wire29232 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640  &  wire29232 ) ;
 assign wire6947 = ( pg72  &  ng4322  &  wire29233  &  wire29234 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233  &  wire29234 ) ;
 assign wire6948 = ( pg72  &  ng4322  &  wire29233  &  wire29235 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233  &  wire29235 ) ;
 assign wire6949 = ( pg72  &  ng4322  &  wire28640  &  wire29236 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640  &  wire29236 ) ;
 assign wire6950 = ( pg72  &  ng4322  &  wire29233  &  wire29237 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233  &  wire29237 ) ;
 assign wire6951 = ( pg72  &  ng4322  &  wire28640  &  wire29238 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640  &  wire29238 ) ;
 assign wire6952 = ( pg72  &  ng4322  &  wire28640  &  wire29239 ) | ( (~ pg72)  &  (~ ng4322)  &  wire28640  &  wire29239 ) ;
 assign wire6953 = ( pg72  &  ng4322  &  wire29233  &  wire29240 ) | ( (~ pg72)  &  (~ ng4322)  &  wire29233  &  wire29240 ) ;
 assign wire6956 = ( (~ pg35)  &  ng6585 ) ;
 assign wire6959 = ( (~ wire7137)  &  (~ wire7138)  &  (~ wire28996)  &  wire29224 ) ;
 assign wire6960 = ( wire28971  &  wire29225 ) | ( wire28972  &  wire29225 ) | ( wire28995  &  wire29225 ) ;
 assign wire6965 = ( (~ pg35)  &  ng3457 ) ;
 assign wire6966 = ( ng4991  &  ng4871 ) | ( (~ ng4966)  &  ng4871 ) | ( ng4871  &  ng4983 ) ;
 assign wire6967 = ( (~ ng4859)  &  ng4871 ) | ( (~ ng4849)  &  ng4871 ) | ( (~ ng4843)  &  ng4871 ) ;
 assign wire6985 = ( (~ pg35)  &  ng499 ) ;
 assign wire6988 = ( (~ pg35)  &  ng5180 ) ;
 assign wire6992 = ( (~ pg35)  &  ng2803 ) ;
 assign wire7004 = ( ng29503  &  ng27416  &  ng17317  &  wire29159 ) ;
 assign wire7005 = ( ng29503  &  ng27416  &  ng17317  &  wire29161 ) ;
 assign wire7006 = ( (~ ng29503)  &  wire29162 ) | ( (~ ng27416)  &  wire29162 ) | ( (~ ng17317)  &  wire29162 ) ;
 assign wire7007 = ( (~ pg35)  &  ng1728 ) ;
 assign wire7008 = ( (~ pg17685)  &  (~ pg13085)  &  ng10207  &  wire29138 ) ;
 assign wire7009 = ( pg12422  &  (~ pg13085)  &  ng10207  &  wire29143 ) ;
 assign wire7010 = ( pg12422  &  (~ pg13085)  &  ng10207  &  wire29148 ) ;
 assign wire7011 = ( pg17685  &  pg12422  &  ng10207  &  wire29153 ) ;
 assign wire7024 = ( (~ pg35)  &  ng424 ) ;
 assign wire7028 = ( (~ pg35)  &  ng2413 ) ;
 assign wire7030 = ( ng2715  &  ng2724  &  (~ ng2719) ) | ( ng2715  &  ng2729  &  (~ ng2719) ) ;
 assign wire7034 = ( (~ pg35)  &  ng1936 ) ;
 assign wire7041 = ( (~ ng2715)  &  ng2724  &  (~ ng2719) ) | ( (~ ng2715)  &  ng2729  &  (~ ng2719) ) ;
 assign wire7046 = ( ng4991  &  ng4836 ) | ( (~ ng4966)  &  ng4836 ) | ( ng4836  &  ng4983 ) ;
 assign wire7047 = ( (~ ng4859)  &  ng4836 ) | ( (~ ng4849)  &  ng4836 ) | ( (~ ng4843)  &  ng4836 ) ;
 assign wire7049 = ( (~ ng13378)  &  (~ ng13315)  &  wire29072  &  wire29073 ) ;
 assign wire7050 = ( ng13378  &  (~ ng13315)  &  wire29076  &  wire29077 ) ;
 assign wire7058 = ( (~ ng28880)  &  ng26793  &  wire29063 ) | ( (~ ng28880)  &  ng14506  &  wire29063 ) ;
 assign wire7059 = ( pg35  &  ng2599  &  (~ ng26793)  &  (~ ng14506) ) ;
 assign wire7065 = ( ng2689  &  ng2697  &  ng2704 ) ;
 assign wire7069 = ( (~ pg35)  &  ng6633 ) ;
 assign wire7077 = ( (~ pg35)  &  ng3905 ) ;
 assign wire7078 = ( pg35  &  (~ ng911)  &  ng907  &  ng19063 ) ;
 assign wire7083 = ( (~ pg35)  &  ng3917 ) ;
 assign wire7096 = ( wire29028  &  wire29030 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire29030 ) ;
 assign wire7097 = ( (~ pg35)  &  ng2181 ) ;
 assign wire7100 = ( (~ pg35)  &  ng6259 ) ;
 assign wire7102 = ( ng925  &  (~ ng918)  &  ng22992 ) | ( ng925  &  ng22992  &  ng25888 ) ;
 assign wire7114 = ( (~ pg35)  &  ng3570 ) ;
 assign wire7116 = ( wire29011  &  wire29013 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire29013 ) ;
 assign wire7117 = ( (~ pg35)  &  ng2008 ) ;
 assign wire7126 = ( ng2145  &  ng2138  &  ng2130 ) ;
 assign wire7131 = ( wire28971  &  wire29000 ) | ( wire28972  &  wire29000 ) | ( wire28995  &  wire29000 ) ;
 assign wire7132 = ( (~ wire28971)  &  (~ wire28972)  &  (~ wire28995)  &  wire29002 ) ;
 assign wire7133 = ( (~ wire7137)  &  (~ wire7138)  &  (~ wire28996)  &  wire29003 ) ;
 assign wire7134 = ( (~ pg35)  &  ng3111 ) ;
 assign wire7137 = ( ng4991  &  ng4864 ) | ( ng4864  &  (~ ng4966) ) | ( ng4864  &  ng4983 ) ;
 assign wire7138 = ( (~ ng4859)  &  ng4864 ) | ( ng4864  &  (~ ng4849) ) | ( ng4864  &  (~ ng4843) ) ;
 assign wire7167 = ( (~ pg35)  &  ng3897 ) ;
 assign wire7170 = ( (~ pg35)  &  ng5583 ) ;
 assign wire7175 = ( (~ pg35)  &  ng3957 ) ;
 assign wire7180 = ( wire28919  &  wire28921 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire28921 ) ;
 assign wire7181 = ( (~ pg35)  &  ng2165 ) ;
 assign wire7186 = ( (~ ng2815)  &  (~ ng2803)  &  (~ ng2724) ) ;
 assign wire7187 = ( (~ ng2819)  &  ng2724  &  ng2729 ) ;
 assign wire7190 = ( (~ pg35)  &  ng1536 ) ;
 assign wire7193 = ( ng11869  &  (~ ng7620)  &  ng10918  &  wire28898 ) ;
 assign wire7199 = ( wire7257  &  wire28878 ) | ( ng14367  &  wire28834  &  wire28878 ) ;
 assign wire7200 = ( wire7257  &  wire28881 ) | ( ng14367  &  wire28834  &  wire28881 ) ;
 assign wire7201 = ( wire7257  &  wire28883 ) | ( ng14367  &  wire28834  &  wire28883 ) ;
 assign wire7202 = ( wire7257  &  wire28884 ) | ( ng14367  &  wire28834  &  wire28884 ) ;
 assign wire7204 = ( (~ ng14367)  &  (~ wire7257)  &  wire28886 ) | ( (~ wire7257)  &  (~ wire28834)  &  wire28886 ) ;
 assign wire7205 = ( (~ pg35)  &  ng1792 ) ;
 assign wire7221 = ( (~ pg35)  &  ng6287 ) ;
 assign wire7225 = ( (~ pg35)  &  ng2807 ) ;
 assign wire7232 = ( (~ ng14367)  &  (~ wire7257)  &  wire28854 ) | ( (~ wire7257)  &  (~ wire28834)  &  wire28854 ) ;
 assign wire7233 = ( ng1760  &  wire7257 ) | ( ng1760  &  ng14367  &  wire28834 ) ;
 assign wire7236 = ( wire28848  &  wire28850 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire28850 ) ;
 assign wire7237 = ( (~ pg35)  &  ng2177 ) ;
 assign wire7248 = ( ng4801  &  ng4688 ) | ( ng4793  &  ng4688 ) | ( ng4688  &  (~ ng4776) ) ;
 assign wire7249 = ( (~ ng4653)  &  ng4688 ) | ( (~ ng4669)  &  ng4688 ) | ( ng4688  &  (~ ng4659) ) ;
 assign wire7255 = ( (~ pg35)  &  ng1748 ) ;
 assign wire7257 = ( ng2715  &  ng2724  &  (~ ng2719) ) | ( ng2715  &  ng2729  &  (~ ng2719) ) ;
 assign wire7259 = ( wire28829  &  wire28831 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire28831 ) ;
 assign wire7260 = ( (~ pg35)  &  ng1874 ) ;
 assign wire7269 = ( (~ ng2145)  &  ng2138  &  ng2130 ) ;
 assign wire7283 = ( (~ pg35)  &  ng776 ) ;
 assign wire7284 = ( pg12184  &  (~ pg11678) ) ;
 assign wire7286 = ( (~ ng27629)  &  wire28806 ) | ( wire28803  &  wire28806 ) | ( (~ wire28804)  &  wire28806 ) ;
 assign wire7287 = ( ng27629  &  (~ wire28803)  &  wire28804  &  wire28807 ) ;
 assign wire7291 = ( (~ pg35)  &  ng586 ) ;
 assign wire7298 = ( ng9649  &  ng26703  &  wire28786 ) | ( ng9649  &  ng17321  &  wire28786 ) ;
 assign wire7299 = ( ng9649  &  ng26703  &  wire28787 ) | ( ng9649  &  ng17321  &  wire28787 ) ;
 assign wire7300 = ( (~ ng9649)  &  wire28788 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire28788 ) ;
 assign wire7301 = ( (~ pg35)  &  ng2265 ) ;
 assign wire7306 = ( ng2689  &  (~ ng2697)  &  (~ ng2704) ) ;
 assign wire7308 = ( (~ pg134)  &  ng209 ) | ( (~ pg134)  &  (~ ng691) ) ;
 assign wire7309 = ( (~ pg134)  &  (~ ng1536) ) | ( (~ pg134)  &  (~ ng1312)  &  (~ ng1351) ) ;
 assign wire7310 = ( pg35  &  ng499  &  (~ ng513) ) ;
 assign wire7321 = ( ng10756  &  wire28765  &  wire28769 ) | ( ng10756  &  wire28766  &  wire28769 ) ;
 assign wire7322 = ( ng10756  &  wire28765  &  wire28770 ) | ( ng10756  &  wire28766  &  wire28770 ) ;
 assign wire7323 = ( ng19984  &  (~ ng10756) ) | ( ng19984  &  (~ wire28765)  &  (~ wire28766) ) ;
 assign wire7324 = ( (~ pg35)  &  ng3808 ) ;
 assign wire7325 = ( (~ ng4955)  &  ng4878 ) ;
 assign wire7326 = ( (~ ng4859)  &  ng4878 ) | ( (~ ng4849)  &  ng4878 ) | ( (~ ng4843)  &  ng4878 ) ;
 assign wire7331 = ( (~ ng10939)  &  (~ ng13378)  &  wire28742  &  wire28743 ) ;
 assign wire7332 = ( (~ ng10939)  &  ng13378  &  wire28746  &  wire28747 ) ;
 assign wire7346 = ( pg35  &  ng333  &  ng351 ) | ( pg35  &  ng355  &  ng351 ) ;
 assign wire7351 = ( ng4801  &  ng4681 ) | ( ng4681  &  ng4793 ) | ( ng4681  &  (~ ng4776) ) ;
 assign wire7352 = ( ng4681  &  (~ ng4653) ) | ( ng4681  &  (~ ng4669) ) | ( ng4681  &  (~ ng4659) ) ;
 assign wire7371 = ( wire29984  &  (~ wire30193)  &  (~ wire30194) ) | ( wire29985  &  (~ wire30193)  &  (~ wire30194) ) ;
 assign wire7372 = ( (~ pg54)  &  (~ pg53)  &  ng7 ) | ( (~ pg53)  &  ng7  &  (~ wire29926) ) ;
 assign wire7373 = ( (~ ng947)  &  ng1129  &  ni17529  &  wire30000 ) ;
 assign wire7374 = ( ng4732  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire7375 = ( ng1472  &  (~ ng1291)  &  ni18740  &  wire30003 ) ;
 assign wire7376 = ( ng4922  &  ng13156  &  wire29937  &  wire30042 ) ;
 assign wire7377 = ( ng5853  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7378 = ( (~ ng13156)  &  wire30190 ) | ( (~ wire29957)  &  wire30190 ) | ( (~ wire29978)  &  wire30190 ) ;
 assign wire7382 = ( wire29984  &  wire30217 ) | ( wire29985  &  wire30217 ) ;
 assign wire7390 = ( ng6199  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7391 = ( (~ pg54)  &  (~ pg53)  &  ng6 ) | ( (~ pg53)  &  ng6  &  (~ wire29926) ) ;
 assign wire7392 = ( ng1300  &  (~ ng1291)  &  ni18740  &  wire30003 ) ;
 assign wire7398 = ( ng4917  &  ng13156  &  wire29937  &  wire30042 ) ;
 assign wire7399 = ( ng3853  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7400 = ( ng4727  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire7409 = ( ng5160  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7410 = ( ng6545  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7411 = ( ng4912  &  ng13156  &  wire29937  &  wire30042 ) ;
 assign wire7412 = ( ng4722  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire7414 = ( wire29984  &  wire30118 ) | ( wire29985  &  wire30118 ) ;
 assign wire7424 = ( (~ pg54)  &  (~ pg53)  &  ng9 ) | ( (~ pg53)  &  ng9  &  (~ wire29926) ) ;
 assign wire7426 = ( wire29984  &  wire30162 ) | ( wire29985  &  wire30162 ) ;
 assign wire7436 = ( (~ pg54)  &  (~ pg53)  &  ng8 ) | ( (~ pg53)  &  ng8  &  (~ wire29926) ) ;
 assign wire7437 = ( ng5507  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7438 = ( ng1448  &  (~ ng1291)  &  ni18740  &  wire30003 ) ;
 assign wire7445 = ( ng3151  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7446 = ( ng4907  &  ng13156  &  wire29937  &  wire30042 ) ;
 assign wire7447 = ( ng4717  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire7452 = ( wire29984  &  wire30097 ) | ( wire29985  &  wire30097 ) ;
 assign wire7462 = ( (~ pg54)  &  (~ pg53)  &  ng28 ) | ( (~ pg53)  &  ng28  &  (~ wire29926) ) ;
 assign wire7463 = ( ng939  &  ng13156  &  wire29937  &  wire30000 ) ;
 assign wire7464 = ( ng1283  &  ng13156  &  wire29957  &  wire30003 ) ;
 assign wire7466 = ( wire29948  &  wire30084 ) | ( wire29949  &  wire30084 ) | ( wire29950  &  wire30084 ) ;
 assign wire7467 = ( wire29948  &  wire30085 ) | ( wire29949  &  wire30085 ) | ( wire29950  &  wire30085 ) ;
 assign wire7468 = ( wire29948  &  wire30086 ) | ( wire29949  &  wire30086 ) | ( wire29950  &  wire30086 ) ;
 assign wire7469 = ( wire29948  &  wire30087 ) | ( wire29949  &  wire30087 ) | ( wire29950  &  wire30087 ) ;
 assign wire7470 = ( wire29948  &  wire30088 ) | ( wire29949  &  wire30088 ) | ( wire29950  &  wire30088 ) ;
 assign wire7471 = ( wire29948  &  wire30089 ) | ( wire29949  &  wire30089 ) | ( wire29950  &  wire30089 ) ;
 assign wire7472 = ( ng2697  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7473 = ( ng4146  &  ng17653  &  wire29925  &  wire29926 ) ;
 assign wire7474 = ( ng2138  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7475 = ( wire29984  &  wire30063 ) | ( wire29985  &  wire30063 ) ;
 assign wire7485 = ( ng943  &  ng13156  &  wire29937  &  wire30000 ) ;
 assign wire7486 = ( (~ pg54)  &  (~ pg53)  &  ng31 ) | ( (~ pg53)  &  ng31  &  (~ wire29926) ) ;
 assign wire7487 = ( ng1287  &  ng13156  &  wire29957  &  wire30003 ) ;
 assign wire7489 = ( wire29948  &  wire30055 ) | ( wire29949  &  wire30055 ) | ( wire29950  &  wire30055 ) ;
 assign wire7490 = ( wire29948  &  wire30056 ) | ( wire29949  &  wire30056 ) | ( wire29950  &  wire30056 ) ;
 assign wire7491 = ( wire29948  &  wire30057 ) | ( wire29949  &  wire30057 ) | ( wire29950  &  wire30057 ) ;
 assign wire7492 = ( ng16486  &  wire29948 ) | ( ng16486  &  wire29949 ) | ( ng16486  &  wire29950 ) ;
 assign wire7493 = ( ng2704  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7494 = ( ng4157  &  ng17653  &  wire29925  &  wire29926 ) ;
 assign wire7495 = ( ng2145  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7498 = ( wire29948  &  wire30035 ) | ( wire29949  &  wire30035 ) | ( wire29950  &  wire30035 ) ;
 assign wire7499 = ( wire29948  &  wire30036 ) | ( wire29949  &  wire30036 ) | ( wire29950  &  wire30036 ) ;
 assign wire7500 = ( wire29948  &  wire30037 ) | ( wire29949  &  wire30037 ) | ( wire29950  &  wire30037 ) ;
 assign wire7501 = ( wire29948  &  wire30038 ) | ( wire29949  &  wire30038 ) | ( wire29950  &  wire30038 ) ;
 assign wire7502 = ( wire29948  &  wire30039 ) | ( wire29949  &  wire30039 ) | ( wire29950  &  wire30039 ) ;
 assign wire7503 = ( ng4300  &  ng13156  &  wire29937  &  wire29997 ) ;
 assign wire7504 = ( ng16486  &  wire29948 ) | ( ng16486  &  wire29949 ) | ( ng16486  &  wire29950 ) ;
 assign wire7505 = ( (~ ng4927)  &  ng13156  &  wire29937  &  wire30042 ) ;
 assign wire7506 = ( (~ ng4737)  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire7507 = ( ng4172  &  ng17653  &  wire29925  &  wire29926 ) ;
 assign wire7509 = ( wire29984  &  wire30016 ) | ( wire29985  &  wire30016 ) ;
 assign wire7518 = ( (~ pg54)  &  (~ pg53)  &  ng16 ) | ( (~ pg53)  &  ng16  &  (~ wire29926) ) ;
 assign wire7521 = ( wire29984  &  wire29986 ) | ( wire29985  &  wire29986 ) ;
 assign wire7531 = ( (~ pg54)  &  (~ pg53)  &  ng19 ) | ( (~ pg53)  &  ng19  &  (~ wire29926) ) ;
 assign wire7532 = ( (~ ng952)  &  ng13156  &  wire29937  &  wire30000 ) ;
 assign wire7533 = ( (~ ng1296)  &  ng13156  &  wire29957  &  wire30003 ) ;
 assign wire7540 = ( wire29948  &  wire29952 ) | ( wire29949  &  wire29952 ) | ( wire29950  &  wire29952 ) ;
 assign wire7541 = ( wire29948  &  wire29953 ) | ( wire29949  &  wire29953 ) | ( wire29950  &  wire29953 ) ;
 assign wire7542 = ( wire29948  &  wire29954 ) | ( wire29949  &  wire29954 ) | ( wire29950  &  wire29954 ) ;
 assign wire7543 = ( wire29948  &  wire29955 ) | ( wire29949  &  wire29955 ) | ( wire29950  &  wire29955 ) ;
 assign wire7544 = ( wire29948  &  wire29956 ) | ( wire29949  &  wire29956 ) | ( wire29950  &  wire29956 ) ;
 assign wire7545 = ( ng4176  &  ng17653  &  wire29925  &  wire29926 ) ;
 assign wire7546 = ( ng2130  &  ng13156  &  wire29957  &  wire29962 ) ;
 assign wire7547 = ( ng2689  &  ng13156  &  wire29963  &  wire29966 ) ;
 assign wire7559 = ( (~ pg35)  &  ng6597 ) ;
 assign wire7565 = ( (~ pg35)  &  ng6601 ) ;
 assign wire7567 = ( ng7601  &  wire28720 ) | ( (~ ng1345)  &  (~ ng15748)  &  wire28720 ) ;
 assign wire7568 = ( (~ pg35)  &  ng1345 ) ;
 assign wire7581 = ( (~ pg35)  &  ng157 ) ;
 assign wire7582 = ( ng160  &  ng28353  &  (~ wire28711)  &  wire28712 ) ;
 assign wire7583 = ( (~ pg35)  &  ng160 ) ;
 assign wire7595 = ( (~ ng28761)  &  ng17317  &  wire28689 ) | ( (~ ng28761)  &  ng26694  &  wire28689 ) ;
 assign wire7596 = ( pg35  &  ng1772  &  (~ ng17317)  &  (~ ng26694) ) ;
 assign wire7606 = ( ng2145  &  (~ ng2138)  &  ng2130 ) ;
 assign wire7608 = ( (~ pg134)  &  ng209 ) | ( (~ pg134)  &  (~ ng691) ) ;
 assign wire7609 = ( (~ pg134)  &  (~ ng1193) ) | ( (~ pg134)  &  (~ ng969)  &  (~ ng1008) ) ;
 assign wire7623 = ( (~ pg35)  &  ng5134 ) ;
 assign wire7624 = ( ng4801  &  ng4646 ) | ( ng4646  &  ng4793 ) | ( ng4646  &  (~ ng4776) ) ;
 assign wire7625 = ( ng4646  &  (~ ng4653) ) | ( ng4646  &  (~ ng4669) ) | ( ng4646  &  (~ ng4659) ) ;
 assign wire7634 = ( (~ pg35)  &  ng4793 ) ;
 assign wire7639 = ( (~ ng1926)  &  ng1917  &  ng25357  &  wire28614 ) ;
 assign wire7640 = ( ng2051  &  (~ ng2060)  &  ng25357  &  wire28617 ) ;
 assign wire7641 = ( ng1783  &  (~ ng1792)  &  ng12377  &  ng25357 ) ;
 assign wire7642 = ( ng2610  &  (~ ng2619)  &  ng25357  &  wire28622 ) ;
 assign wire7643 = ( (~ ng2217)  &  ng2208  &  ng25357  &  wire28625 ) ;
 assign wire7644 = ( (~ ng2485)  &  ng2476  &  ng25357  &  wire28503 ) ;
 assign wire7645 = ( ng2342  &  (~ ng2351)  &  ng25357  &  wire28629 ) ;
 assign wire7646 = ( (~ ng1657)  &  ng1648  &  ng25357  &  wire28632 ) ;
 assign wire7647 = ( pg35  &  (~ ng25911)  &  wire7650  &  (~ wire7652) ) ;
 assign wire7649 = ( (~ pg35)  &  ng1024 ) ;
 assign wire7650 = ( (~ ng1030)  &  (~ ng15737) ) ;
 assign wire7652 = ( (~ ng1024)  &  (~ ng15737) ) ;
 assign wire7662 = ( pg72  &  pg35  &  ng225  &  ng239 ) ;
 assign wire7663 = ( pg73  &  pg72  &  pg35  &  ng225 ) ;
 assign wire7664 = ( (~ pg72)  &  pg35  &  ng246  &  ng232 ) ;
 assign wire7665 = ( pg73  &  (~ pg72)  &  pg35  &  ng232 ) ;
 assign wire7666 = ( (~ pg73)  &  pg72  &  pg35  &  ng239 ) ;
 assign wire7667 = ( (~ pg73)  &  (~ pg72)  &  pg35  &  ng246 ) ;
 assign wire7668 = ( (~ pg35)  &  ng479 ) ;
 assign wire7671 = ( (~ pg35)  &  ng269 ) ;
 assign wire7677 = ( (~ pg35)  &  ng437 ) ;
 assign wire7681 = ( (~ pg35)  &  ng4894 ) ;
 assign wire7685 = ( (~ pg35)  &  ng2819 ) ;
 assign wire7686 = ( ng28444  &  (~ wire28561)  &  wire28562  &  wire28563 ) ;
 assign wire7690 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28530 ) ;
 assign wire7691 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28532 ) ;
 assign wire7692 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28534 ) ;
 assign wire7693 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28536 ) ;
 assign wire7694 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28538 ) ;
 assign wire7695 = ( (~ ng11676)  &  wire28525  &  wire28526  &  wire28540 ) ;
 assign wire7703 = ( (~ pg35)  &  ng3219 ) ;
 assign wire7709 = ( ng11846  &  wire28514  &  wire28515 ) ;
 assign wire7720 = ( (~ ng14367)  &  (~ wire7725)  &  wire28490 ) | ( (~ wire7725)  &  (~ wire28488)  &  wire28490 ) ;
 assign wire7721 = ( wire7725  &  wire28491 ) | ( ng14367  &  wire28488  &  wire28491 ) ;
 assign wire7725 = ( (~ ng2715)  &  ng2724  &  ng2719 ) | ( (~ ng2715)  &  ng2729  &  ng2719 ) ;
 assign wire7734 = ( (~ ng18935)  &  (~ ng30583)  &  ng15591  &  wire28476 ) ;
 assign wire7735 = ( ng18935  &  (~ ng30583)  &  ng15591  &  wire28478 ) ;
 assign wire28470 = ( ng4087  &  (~ ng4098)  &  ng4093 ) ;
 assign wire28473 = ( pg35  &  (~ ng6215)  &  ng6209  &  ng6203 ) ;
 assign wire28475 = ( (~ ng4322) ) | ( (~ ng4332) ) ;
 assign wire28476 = ( ng4332  &  pg35 ) ;
 assign wire28478 = ( (~ ng4332)  &  pg35 ) ;
 assign wire28482 = ( ng1094  &  (~ ng1135) ) ;
 assign wire28483 = ( ng1135  &  pg35 ) ;
 assign wire28484 = ( (~ pg35)  &  ng1094 ) | ( pg35  &  ng1135  &  (~ ng1094) ) ;
 assign wire28485 = ( wire28484 ) | ( (~ ng10929)  &  (~ ng13846)  &  wire28482 ) ;
 assign wire28488 = ( (~ ng2815)  &  (~ ng2715)  &  ng2719 ) ;
 assign wire28490 = ( ng2485  &  pg35 ) ;
 assign wire28491 = ( ng2476  &  pg35 ) ;
 assign wire28503 = ( ng2756  &  (~ ng2741)  &  ng2748 ) ;
 assign wire28505 = ( pg35  &  wire7725 ) | ( pg35  &  ng14367  &  wire28488 ) ;
 assign wire28507 = ( wire7721 ) | ( (~ ng27903)  &  wire28505 ) ;
 assign wire28514 = ( pg7916  &  ng990 ) | ( pg7916  &  ng979 ) ;
 assign wire28515 = ( ng979  &  ng1178  &  (~ ng1189)  &  ng996 ) ;
 assign wire28519 = ( pg7916  &  ng969  &  ng10893 ) | ( pg7916  &  ng1008  &  ng10893 ) ;
 assign wire28521 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28522 = ( ng3235  &  pg35 ) ;
 assign wire28525 = ( (~ ng528)  &  (~ ng482) ) ;
 assign wire28526 = ( (~ ng499)  &  (~ ng518)  &  (~ ng490) ) ;
 assign wire28530 = ( ng718  &  (~ ng753)  &  (~ ng554) ) | ( ng655  &  (~ ng753)  &  (~ ng554) ) ;
 assign wire28532 = ( ng718  &  (~ ng753)  &  (~ ng807) ) | ( ng655  &  (~ ng753)  &  (~ ng807) ) ;
 assign wire28534 = ( ng718  &  (~ ng655)  &  (~ ng554) ) | ( (~ ng655)  &  ng753  &  (~ ng554) ) ;
 assign wire28536 = ( (~ ng718)  &  ng655  &  (~ ng554) ) | ( (~ ng718)  &  ng753  &  (~ ng554) ) ;
 assign wire28538 = ( ng718  &  (~ ng655)  &  (~ ng807) ) | ( (~ ng655)  &  ng753  &  (~ ng807) ) ;
 assign wire28540 = ( (~ ng718)  &  ng655  &  (~ ng807) ) | ( (~ ng718)  &  ng753  &  (~ ng807) ) ;
 assign wire28543 = ( wire7695 ) | ( wire7694 ) ;
 assign wire28544 = ( wire7690 ) | ( wire7691 ) | ( wire7692 ) | ( wire7693 ) ;
 assign wire28548 = ( ng246  &  ng232  &  ng239 ) ;
 assign wire28549 = ( (~ ng262)  &  ng225  &  (~ ng255)  &  (~ ng269) ) ;
 assign wire28551 = ( ng691  &  ng278  &  wire28548  &  wire28549 ) ;
 assign wire28555 = ( (~ ng246)  &  (~ ng232)  &  (~ ng239) ) ;
 assign wire28556 = ( ng262  &  (~ ng225)  &  ng255  &  ng269 ) ;
 assign wire28558 = ( ng691  &  (~ ng278)  &  wire28555  &  wire28556 ) ;
 assign wire28561 = ( (~ ng23204) ) | ( (~ ng294) ) ;
 assign wire28562 = ( ng23204  &  ng298 ) ;
 assign wire28563 = ( ng142  &  pg35 ) ;
 assign wire28567 = ( (~ ng2729) ) | ( ng2724 ) ;
 assign wire28568 = ( (~ ng2823)  &  pg35 ) ;
 assign wire28569 = ( (~ ng2724)  &  ng2729  &  (~ ng11405)  &  wire28568 ) ;
 assign wire28571 = ( (~ ng111)  &  (~ ng11405)  &  (~ wire28567) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire28567) ) ;
 assign wire28572 = ( ng2815  &  pg35 ) ;
 assign wire28573 = ( wire7685 ) | ( ng11405  &  wire28572 ) | ( wire28567  &  wire28572 ) ;
 assign wire28574 = ( wire28573 ) | ( (~ ng111)  &  wire28569 ) | ( (~ ng29503)  &  wire28569 ) ;
 assign wire28575 = ( ng4818 ) | ( wire1421 ) ;
 assign wire28577 = ( wire1421  &  ng4894 ) | ( ng4894  &  ng4818 ) | ( ng4894  &  (~ ng24374) ) ;
 assign wire28581 = ( pg35  &  ng4888  &  (~ ng29676) ) | ( pg35  &  ng29676  &  ng30590 ) ;
 assign wire28583 = ( ng269  &  pg35 ) ;
 assign wire28584 = ( ng433  &  pg35 ) ;
 assign wire28587 = ( ng246  &  pg35 ) ;
 assign wire28588 = ( pg14167  &  pg35 ) ;
 assign wire28606 = ( wire7663 ) | ( wire7664 ) | ( wire7665 ) | ( wire7666 ) ;
 assign wire28607 = ( ng1030  &  ng1018  &  ng1008 ) ;
 assign wire28609 = ( (~ ng979)  &  ng1046  &  ng996 ) | ( ng979  &  ng1046  &  (~ ng996) ) | ( (~ ng979)  &  ng996  &  (~ ng1008) ) | ( ng979  &  (~ ng996)  &  (~ ng1008) ) ;
 assign wire28611 = ( ng1030  &  pg35 ) ;
 assign wire28612 = ( wire7649 ) | ( ng25911  &  wire28611 ) | ( wire7652  &  wire28611 ) ;
 assign wire28614 = ( (~ ng2756)  &  (~ ng2741)  &  ng2748 ) ;
 assign wire28617 = ( (~ ng2756)  &  ng2741  &  ng2748 ) ;
 assign wire28622 = ( ng2756  &  ng2741  &  ng2748 ) ;
 assign wire28625 = ( ng2756  &  (~ ng2741)  &  (~ ng2748) ) ;
 assign wire28629 = ( ng2756  &  ng2741  &  (~ ng2748) ) ;
 assign wire28632 = ( (~ ng2756)  &  (~ ng2741)  &  (~ ng2748) ) ;
 assign wire28637 = ( wire7639 ) | ( wire7640 ) | ( wire7641 ) | ( wire7642 ) ;
 assign wire28638 = ( wire7643 ) | ( wire7644 ) | ( wire7645 ) | ( wire7646 ) ;
 assign wire28640 = ( pg73  &  ng4332  &  (~ ng4311) ) | ( (~ pg73)  &  (~ ng4332)  &  (~ ng4311) ) ;
 assign wire28643 = ( pg35  &  (~ ng4801)  &  ng4793  &  ng10831 ) ;
 assign wire28645 = ( pg35  &  ng4801  &  (~ ng4793) ) | ( pg35  &  ng4801  &  (~ ng10831) ) ;
 assign wire28646 = ( wire7634 ) | ( ng28336  &  ng13464  &  wire28643 ) ;
 assign wire28651 = ( ng4646  &  ng4785 ) | ( ng4646  &  (~ ng4698) ) | ( ng4646  &  ng4709 ) ;
 assign wire28655 = ( pg35  &  (~ ng5128)  &  (~ ng5134) ) ;
 assign wire28657 = ( ng5138  &  pg35 ) ;
 assign wire28659 = ( ng23590  &  wire28657 ) | ( ng5128  &  ng5134  &  (~ ng23590) ) ;
 assign wire28661 = ( ng4087  &  ng4098  &  ng4093 ) ;
 assign wire28670 = ( (~ pg35)  &  ng3802 ) | ( pg35  &  pg8344  &  (~ pg8398)  &  (~ ng3802) ) ;
 assign wire28673 = ( pg17316  &  (~ ng979) ) | ( pg17316  &  (~ ng1061) ) ;
 assign wire28687 = ( ng504  &  (~ ng518)  &  (~ ng528) ) ;
 assign wire28689 = ( ng1728  &  pg35 ) ;
 assign wire28694 = ( ng4087  &  ng4098  &  (~ ng4093) ) ;
 assign wire28706 = ( (~ ng168)  &  (~ ng182)  &  ng691  &  (~ ng174) ) ;
 assign wire28707 = ( ng513  &  ng691 ) | ( (~ ng518)  &  ng691 ) | ( ng691  &  (~ ng203) ) ;
 assign wire28708 = ( (~ ng513)  &  ng518  &  ng203  &  ng146 ) ;
 assign wire28711 = ( (~ ng23042) ) | ( (~ ng153) ) ;
 assign wire28712 = ( ng23042  &  ng157 ) ;
 assign wire28713 = ( ng23042  &  ng160 ) ;
 assign wire28715 = ( wire7581 ) | ( (~ wire7582)  &  (~ wire7583)  &  wire28713 ) ;
 assign wire28716 = ( ng1361  &  ng1351  &  ng1373 ) ;
 assign wire28718 = ( (~ ng1322)  &  ng1389  &  ng1339 ) | ( (~ ng1322)  &  (~ ng1351)  &  ng1339 ) | ( ng1322  &  ng1389  &  (~ ng1339) ) | ( ng1322  &  (~ ng1351)  &  (~ ng1339) ) ;
 assign wire28719 = ( pg35  &  ng1345  &  (~ ng7601) ) | ( pg35  &  (~ ng7601)  &  ng15748 ) ;
 assign wire28720 = ( ng1361  &  pg35 ) ;
 assign wire28722 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28723 = ( ng6621  &  pg35 ) ;
 assign wire28731 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28732 = ( ng6593  &  pg35 ) ;
 assign wire28733 = ( wire7559 ) | ( ng12632  &  ng12716  &  wire28731 ) ;
 assign wire28734 = ( ng4681  &  ng4785 ) | ( ng4681  &  (~ ng4754) ) | ( ng4681  &  (~ ng4709) ) ;
 assign wire28741 = ( (~ pg35)  &  ng355 ) | ( pg35  &  ng74  &  (~ ng351) ) ;
 assign wire28742 = ( ng1484  &  pg35 ) ;
 assign wire28743 = ( ng1300  &  ng1442 ) | ( ng1300  &  ng1489 ) ;
 assign wire28746 = ( ng1484  &  pg35 ) ;
 assign wire28747 = ( (~ ng1300)  &  ng1442 ) | ( (~ ng1300)  &  ng1489 ) ;
 assign wire28751 = ( pg35  &  ng1300  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire28754 = ( pg35  &  (~ ng1300)  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire28757 = ( (~ pg35)  &  ng1472 ) | ( pg35  &  ng1484  &  ng10939 ) ;
 assign wire28758 = ( (~ ng10939)  &  (~ ng13378)  &  wire28751 ) | ( (~ ng10939)  &  ng13378  &  wire28754 ) ;
 assign wire28765 = ( wire7326 ) | ( (~ ng4955)  &  ng4878 ) ;
 assign wire28766 = ( (~ ng4975)  &  ng10862 ) | ( (~ ng4899)  &  ng10862 ) | ( ng11173  &  ng10862 ) ;
 assign wire28769 = ( pg35  &  (~ ng3808)  &  ng3813 ) ;
 assign wire28770 = ( (~ ng3813)  &  ng3808 ) ;
 assign wire28775 = ( ng499  &  pg35 ) ;
 assign wire28776 = ( pg35  &  ng667  &  (~ ng686) ) ;
 assign wire28779 = ( ng11607  &  wire28776 ) | ( pg35  &  (~ ng518)  &  ng11607 ) ;
 assign wire28783 = ( pg17320  &  (~ ng1322) ) | ( pg17320  &  (~ ng1404) ) ;
 assign wire28786 = ( pg35  &  (~ ng2259)  &  (~ ng2265) ) ;
 assign wire28787 = ( ng2265  &  ng2259 ) ;
 assign wire28788 = ( ng2269  &  pg35 ) ;
 assign wire28792 = ( pg35  &  (~ pg44) ) | ( pg35  &  ng2927 ) ;
 assign wire28793 = ( (~ ng562) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire28794 = ( (~ pg9048)  &  ng568 ) | ( ng568  &  ng559 ) ;
 assign wire28795 = ( (~ ng572) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire28796 = ( (~ pg9048)  &  ng586 ) | ( ng559  &  ng586 ) ;
 assign wire28798 = ( pg35  &  (~ pg9048)  &  ng577 ) | ( pg35  &  ng577  &  ng559 ) ;
 assign wire28799 = ( (~ ng577)  &  pg35 ) ;
 assign wire28800 = ( wire7291 ) | ( ng23978  &  wire28798 ) | ( (~ wire28796)  &  wire28798 ) ;
 assign wire28801 = ( (~ ng577) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire28802 = ( (~ pg9048)  &  ng582 ) | ( ng582  &  ng559 ) ;
 assign wire28803 = ( (~ ng590) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire28804 = ( (~ pg9048)  &  ng595 ) | ( ng559  &  ng595 ) ;
 assign wire28806 = ( pg35  &  (~ pg9048)  &  ng599 ) | ( pg35  &  ng599  &  ng559 ) ;
 assign wire28807 = ( (~ ng599)  &  pg35 ) ;
 assign wire28809 = ( (~ pg11678)  &  ng739 ) | ( ng739  &  ng736 ) ;
 assign wire28810 = ( (~ ng744) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire28811 = ( (~ pg11678)  &  ng749 ) | ( ng736  &  ng749 ) ;
 assign wire28812 = ( (~ ng758) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire28813 = ( (~ pg11678)  &  ng763 ) | ( ng763  &  ng736 ) ;
 assign wire28814 = ( (~ ng767) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire28815 = ( (~ pg11678)  &  ng772 ) | ( ng736  &  ng772 ) ;
 assign wire28816 = ( (~ ng776) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire28818 = ( pg35  &  (~ pg11678)  &  ng781 ) | ( pg35  &  ng781  &  ng736 ) ;
 assign wire28819 = ( (~ ng781)  &  pg35 ) ;
 assign wire28820 = ( wire7283 ) | ( (~ ng32212)  &  wire28818 ) | ( wire28816  &  wire28818 ) ;
 assign wire28821 = ( (~ ng2759)  &  pg35 ) ;
 assign wire28822 = ( ng2759  &  pg35 ) ;
 assign wire28823 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng2756 ) ;
 assign wire28824 = ( wire28823 ) | ( ng2756  &  ng25317  &  wire28821 ) ;
 assign wire28827 = ( pg17400  &  (~ ng979) ) | ( pg17400  &  (~ ng1061) ) ;
 assign wire28829 = ( ng1906 ) | ( (~ ng1862) ) ;
 assign wire28830 = ( pg35  &  ng26725  &  (~ wire28829) ) | ( pg35  &  ng17401  &  (~ wire28829) ) ;
 assign wire28831 = ( ng1870  &  pg35 ) ;
 assign wire28834 = ( ng2715  &  (~ ng2775)  &  (~ ng2719) ) ;
 assign wire28836 = ( ng1792 ) | ( (~ ng1783) ) ;
 assign wire28837 = ( ng1728  &  pg35 ) ;
 assign wire28841 = ( pg35  &  ng1768  &  ng25385 ) | ( pg35  &  (~ ng1772)  &  (~ ng25385) ) ;
 assign wire28843 = ( (~ ng4765)  &  ng4688 ) | ( (~ ng4785)  &  ng4688 ) | ( ng4688  &  (~ ng4709) ) ;
 assign wire28848 = ( (~ ng2227) ) | ( (~ ng2153) ) ;
 assign wire28849 = ( pg35  &  ng26703  &  (~ wire28848) ) | ( pg35  &  ng17321  &  (~ wire28848) ) ;
 assign wire28850 = ( ng2173  &  pg35 ) ;
 assign wire28853 = ( pg35  &  wire7257 ) | ( pg35  &  ng14367  &  wire28834 ) ;
 assign wire28854 = ( ng1783  &  pg35 ) ;
 assign wire28856 = ( wire7233 ) | ( (~ ng27775)  &  wire28853 ) ;
 assign wire28858 = ( pg35  &  (~ ng341)  &  ng329 ) ;
 assign wire28860 = ( (~ ng111)  &  ng12026  &  (~ ng11405) ) | ( (~ ng29503)  &  ng12026  &  (~ ng11405) ) ;
 assign wire28861 = ( (~ ng2799)  &  pg35 ) ;
 assign wire28862 = ( (~ ng2724)  &  (~ ng2729)  &  (~ ng11405)  &  wire28861 ) ;
 assign wire28863 = ( ng2803  &  pg35 ) ;
 assign wire28864 = ( wire7225 ) | ( (~ ng12026)  &  wire28863 ) | ( ng11405  &  wire28863 ) ;
 assign wire28865 = ( wire28864 ) | ( (~ ng111)  &  wire28862 ) | ( (~ ng29503)  &  wire28862 ) ;
 assign wire28866 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28867 = ( ng6303  &  pg35 ) ;
 assign wire28874 = ( (~ pg35)  &  ng528 ) | ( pg35  &  ng667  &  (~ ng686) ) ;
 assign wire28878 = ( pg35  &  ng1748  &  (~ ng1792)  &  (~ ng1760) ) ;
 assign wire28881 = ( pg35  &  (~ ng1783)  &  ng1752  &  ng1760 ) ;
 assign wire28883 = ( pg35  &  ng1783  &  (~ ng1760)  &  ng1736 ) ;
 assign wire28884 = ( (~ ng1783)  &  ng1792  &  ng1744 ) ;
 assign wire28885 = ( ng1756  &  pg35 ) ;
 assign wire28886 = ( ng1811  &  pg35 ) ;
 assign wire28887 = ( (~ ng1760) ) | ( (~ ng1792) ) ;
 assign wire28891 = ( ng1740  &  (~ ng25300) ) | ( (~ ng25385)  &  wire28885 ) ;
 assign wire28892 = ( wire7199 ) | ( wire7200 ) | ( wire7201 ) | ( wire7205 ) ;
 assign wire28896 = ( pg7946  &  (~ ng1514)  &  ng1526 ) ;
 assign wire28898 = ( pg7946  &  ng1322 ) | ( pg7946  &  ng1333 ) ;
 assign wire28903 = ( pg7946  &  ng1312  &  ng10918 ) | ( pg7946  &  ng1351  &  ng10918 ) ;
 assign wire28905 = ( pg35  &  ng1542  &  ng10918 ) | ( pg35  &  ng1542  &  (~ wire28896) ) ;
 assign wire28907 = ( pg35  &  (~ ng1542)  &  (~ ng10918)  &  wire28896 ) ;
 assign wire28915 = ( (~ ng2819)  &  ng2724  &  (~ ng2807) ) | ( ng2724  &  (~ ng2729)  &  (~ ng2807) ) ;
 assign wire28916 = ( (~ ng2815)  &  (~ ng2724)  &  ng2729 ) | ( (~ ng2803)  &  (~ ng2724)  &  (~ ng2729) ) ;
 assign wire28919 = ( (~ ng2153) ) | ( ng2197 ) ;
 assign wire28920 = ( pg35  &  ng26703  &  (~ wire28919) ) | ( pg35  &  ng17321  &  (~ wire28919) ) ;
 assign wire28921 = ( ng2161  &  pg35 ) ;
 assign wire28924 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28925 = ( ng3913  &  pg35 ) ;
 assign wire28927 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28928 = ( ng5599  &  pg35 ) ;
 assign wire28931 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire28932 = ( ng3893  &  pg35 ) ;
 assign wire28933 = ( wire7167 ) | ( ng11626  &  ng11763  &  wire28931 ) ;
 assign wire28935 = ( (~ ng4141)  &  ng4064  &  ng4057 ) ;
 assign wire28937 = ( ng4141  &  (~ ng4064) ) | ( ng4141  &  (~ ng4057) ) ;
 assign wire28938 = ( (~ pg35)  &  ng4057 ) | ( pg35  &  ng2841  &  wire28935 ) ;
 assign wire28940 = ( pg16718  &  ng3235  &  ng3352  &  ng3288 ) ;
 assign wire28941 = ( ng3338  &  pg16686 ) ;
 assign wire28942 = ( ng3352  &  ng3288  &  ng3247 ) ;
 assign wire28943 = ( ng3223  &  pg16874 ) ;
 assign wire28944 = ( ng3352  &  (~ ng3338)  &  ng3288 ) ;
 assign wire28945 = ( ng3338  &  pg16874 ) ;
 assign wire28946 = ( ng3352  &  ng3215  &  (~ ng3288) ) ;
 assign wire28947 = ( ng3191  &  pg11349 ) ;
 assign wire28949 = ( ng3203  &  pg16624 ) ;
 assign wire28952 = ( pg13895  &  ng3219  &  (~ ng3352)  &  ng3288 ) ;
 assign wire28953 = ( ng3231  &  pg13865 ) ;
 assign wire28954 = ( (~ ng3352)  &  ng3338  &  ng3288 ) ;
 assign wire28955 = ( (~ ng3338)  &  pg14421 ) ;
 assign wire28956 = ( (~ ng3352)  &  ng3288  &  ng3199 ) ;
 assign wire28958 = ( pg16603  &  (~ ng3352)  &  ng3251  &  (~ ng3288) ) ;
 assign wire28959 = ( ng3329  &  ng3195 ) ;
 assign wire28961 = ( ng3187  &  pg14421 ) ;
 assign wire28963 = ( (~ ng11350)  &  wire28940 ) | ( wire28941  &  wire28942 ) ;
 assign wire28964 = ( wire28943  &  wire28944 ) | ( wire28945  &  wire28946 ) ;
 assign wire28965 = ( ng3338  &  ng13700  &  wire28947 ) | ( (~ ng3338)  &  ng13700  &  wire28949 ) ;
 assign wire28966 = ( (~ ng11350)  &  wire28952 ) | ( wire28953  &  wire28954 ) ;
 assign wire28967 = ( wire28955  &  wire28956 ) | ( (~ ng11350)  &  wire28958 ) ;
 assign wire28968 = ( ng3338  &  ng11194  &  wire28959 ) | ( ng3338  &  ng11194  &  wire28961 ) ;
 assign wire28971 = ( wire28968 ) | ( wire28967 ) ;
 assign wire28972 = ( wire28963 ) | ( wire28964 ) | ( wire28965 ) | ( wire28966 ) ;
 assign wire28973 = ( ng3207  &  pg11349 ) ;
 assign wire28975 = ( ng3263  &  pg16624 ) ;
 assign wire28978 = ( pg16718  &  ng3243  &  ng3352  &  (~ ng3288) ) ;
 assign wire28979 = ( ng3255  &  pg16686 ) ;
 assign wire28980 = ( ng3352  &  (~ ng3338)  &  (~ ng3288) ) ;
 assign wire28982 = ( pg16603  &  ng3259  &  (~ ng3352)  &  ng3288 ) ;
 assign wire28983 = ( ng3329  &  ng3211 ) ;
 assign wire28984 = ( (~ ng3352)  &  (~ ng3338)  &  ng3288 ) ;
 assign wire28986 = ( pg13895  &  (~ ng3352)  &  ng3227  &  (~ ng3288) ) ;
 assign wire28987 = ( ng3239  &  pg13865 ) ;
 assign wire28988 = ( (~ ng3352)  &  (~ ng3338)  &  (~ ng3288) ) ;
 assign wire28989 = ( (~ ng3338)  &  ng13765  &  wire28973 ) | ( ng3338  &  ng13765  &  wire28975 ) ;
 assign wire28990 = ( ng11350  &  wire28978 ) | ( wire28979  &  wire28980 ) ;
 assign wire28991 = ( ng11350  &  wire28982 ) | ( wire28983  &  wire28984 ) ;
 assign wire28992 = ( ng11350  &  wire28986 ) | ( wire28987  &  wire28988 ) ;
 assign wire28995 = ( wire28989 ) | ( wire28990 ) | ( wire28991 ) | ( wire28992 ) ;
 assign wire28996 = ( (~ ng4975)  &  ng4864 ) | ( ng4899  &  ng4864 ) | ( ng4864  &  (~ ng4933) ) ;
 assign wire29000 = ( pg35  &  (~ ng3106)  &  ng20887 ) | ( pg35  &  ng20887  &  ng10721 ) ;
 assign wire29002 = ( pg35  &  ng3106  &  ng20887  &  (~ ng10721) ) ;
 assign wire29003 = ( ng3106  &  pg35 ) ;
 assign wire29009 = ( (~ ng979)  &  ng1087 ) | ( (~ ng1061)  &  ng1087 ) ;
 assign wire29011 = ( ng2040 ) | ( (~ ng1996) ) ;
 assign wire29012 = ( pg35  &  ng26759  &  (~ wire29011) ) | ( pg35  &  ng14438  &  (~ wire29011) ) ;
 assign wire29013 = ( ng2004  &  pg35 ) ;
 assign wire29015 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29016 = ( ng3586  &  pg35 ) ;
 assign wire29023 = ( (~ pg35)  &  ng918 ) | ( pg35  &  (~ ng925)  &  ng918  &  (~ ng25888) ) ;
 assign wire29025 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29026 = ( ng6255  &  pg35 ) ;
 assign wire29027 = ( wire7100 ) | ( ng12622  &  ng12667  &  wire29025 ) ;
 assign wire29028 = ( ng2153 ) | ( (~ ng2197) ) ;
 assign wire29029 = ( pg35  &  ng26703  &  (~ wire29028) ) | ( pg35  &  ng17321  &  (~ wire29028) ) ;
 assign wire29030 = ( ng2177  &  pg35 ) ;
 assign wire29039 = ( pg72  &  pg35  &  ng4581 ) | ( pg35  &  ng4578  &  ng4581 ) ;
 assign wire29040 = ( (~ pg35)  &  ng4540 ) | ( (~ ng4581)  &  ng4540 ) | ( (~ pg73)  &  pg35  &  ng4581 ) ;
 assign wire29043 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29044 = ( ng3933  &  pg35 ) ;
 assign wire29047 = ( pg35  &  pg12919  &  ng911 ) ;
 assign wire29048 = ( (~ pg35)  &  ng907 ) | ( (~ ng907)  &  wire29047 ) | ( (~ ng19063)  &  wire29047 ) ;
 assign wire29049 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29050 = ( ng3901  &  pg35 ) ;
 assign wire29051 = ( wire7077 ) | ( ng11626  &  ng11537  &  wire29049 ) ;
 assign wire29054 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29055 = ( ng6649  &  pg35 ) ;
 assign wire29058 = ( (~ ng1322)  &  ng1430 ) | ( (~ ng1404)  &  ng1430 ) ;
 assign wire29061 = ( (~ ng504)  &  ng518  &  ng528 ) ;
 assign wire29063 = ( ng2555  &  pg35 ) ;
 assign wire29068 = ( pg35  &  ng4087  &  ng2841 ) ;
 assign wire29070 = ( pg35  &  (~ ng4087)  &  ng2841 ) ;
 assign wire29071 = ( (~ pg35)  &  ng4076 ) | ( (~ ng4076)  &  wire29068 ) | ( ng13217  &  wire29068 ) ;
 assign wire29072 = ( ng1467  &  pg35 ) ;
 assign wire29073 = ( ng1472  &  ng1442 ) | ( ng1472  &  ng1489 ) ;
 assign wire29076 = ( ng1467  &  pg35 ) ;
 assign wire29077 = ( (~ ng1472)  &  ng1442 ) | ( (~ ng1472)  &  ng1489 ) ;
 assign wire29081 = ( pg35  &  ng1472  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire29084 = ( pg35  &  (~ ng1472)  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire29087 = ( (~ pg35)  &  ng1448 ) | ( pg35  &  ng1467  &  ng13315 ) ;
 assign wire29088 = ( (~ ng13378)  &  (~ ng13315)  &  wire29081 ) | ( ng13378  &  (~ ng13315)  &  wire29084 ) ;
 assign wire29091 = ( (~ ng4888)  &  ng4836 ) | ( ng4975  &  ng4836 ) | ( ng4899  &  ng4836 ) ;
 assign wire29097 = ( (~ ng2715)  &  (~ ng2719)  &  (~ ng2771) ) ;
 assign wire29099 = ( (~ ng1657) ) | ( (~ ng1624) ) ;
 assign wire29103 = ( pg35  &  (~ ng1950) ) | ( pg35  &  (~ ng1936)  &  (~ ng1862) ) ;
 assign wire29104 = ( ng26725  &  wire29103 ) | ( ng17401  &  wire29103 ) ;
 assign wire29105 = ( pg35  &  ng1950  &  ng1936 ) | ( pg35  &  ng1950  &  ng1862 ) ;
 assign wire29106 = ( ng26725  &  wire29105 ) | ( ng17401  &  wire29105 ) ;
 assign wire29107 = ( ng1950  &  pg35 ) ;
 assign wire29108 = ( wire7034 ) | ( (~ ng26725)  &  (~ ng17401)  &  wire29107 ) ;
 assign wire29111 = ( ng2715  &  (~ ng2719)  &  (~ ng2807) ) ;
 assign wire29113 = ( (~ ng2351) ) | ( (~ ng2319) ) ;
 assign wire29115 = ( pg35  &  (~ ng2407)  &  (~ ng2413) ) ;
 assign wire29117 = ( ng2417  &  pg35 ) ;
 assign wire29119 = ( ng25349  &  wire29117 ) | ( ng2407  &  ng2413  &  (~ ng25349) ) ;
 assign wire29120 = ( ng246  &  pg35 ) ;
 assign wire29121 = ( ng475  &  pg35 ) ;
 assign wire29124 = ( (~ ng305)  &  (~ ng319)  &  (~ ng311) ) ;
 assign wire29126 = ( pg35  &  (~ ng336)  &  ng311 ) ;
 assign wire29128 = ( pg35  &  ng336  &  ng305 ) ;
 assign wire29129 = ( ng319  &  pg35 ) ;
 assign wire29130 = ( (~ pg35)  &  ng329 ) | ( pg35  &  (~ ng329)  &  wire29124 ) ;
 assign wire29131 = ( ng13385  &  wire29126 ) | ( ng13385  &  wire29128 ) ;
 assign wire29138 = ( pg35  &  (~ pg17760)  &  (~ pg14779)  &  (~ pg17649) ) ;
 assign wire29143 = ( pg35  &  pg17760  &  pg14779  &  (~ pg17685) ) ;
 assign wire29148 = ( pg35  &  (~ pg17760)  &  (~ pg17649)  &  (~ pg17685) ) ;
 assign wire29153 = ( pg35  &  pg17760  &  pg14779  &  pg17649 ) ;
 assign wire29159 = ( pg35  &  (~ ng1772)  &  (~ ng112)  &  ng1802 ) ;
 assign wire29161 = ( pg35  &  ng1772  &  ng112 ) | ( pg35  &  ng112  &  (~ ng1802) ) ;
 assign wire29162 = ( ng1779  &  pg35 ) ;
 assign wire29168 = ( pg35  &  ng2715  &  ng2370 ) ;
 assign wire29171 = ( pg35  &  (~ ng2715)  &  ng2236 ) ;
 assign wire29175 = ( pg35  &  ng2715  &  (~ ng2807) ) ;
 assign wire29178 = ( pg35  &  (~ ng2715)  &  (~ ng2803) ) ;
 assign wire29180 = ( ng2719  &  pg35 ) ;
 assign wire29183 = ( pg35  &  ng2719  &  (~ ng23553) ) ;
 assign wire29184 = ( (~ ng21277)  &  (~ ng23657)  &  wire29168 ) | ( (~ ng21277)  &  (~ ng23657)  &  wire29171 ) ;
 assign wire29185 = ( ng21277  &  (~ ng23553)  &  wire29175 ) | ( ng21277  &  (~ ng23553)  &  wire29178 ) ;
 assign wire29186 = ( ng21277  &  wire29183 ) | ( (~ ng21277)  &  (~ ng23657)  &  wire29180 ) ;
 assign wire29192 = ( (~ ng4087)  &  (~ ng4098)  &  (~ ng4093) ) ;
 assign wire29195 = ( pg35  &  (~ ng5188)  &  ng5176  &  ng5180 ) ;
 assign wire29196 = ( pg35  &  ng5188  &  (~ ng5176) ) | ( pg35  &  ng5188  &  (~ ng5180) ) ;
 assign wire29198 = ( ng504  &  pg35 ) ;
 assign wire29199 = ( pg35  &  ng667  &  (~ ng686) ) ;
 assign wire29202 = ( ng11607  &  wire29199 ) | ( pg35  &  ng499  &  ng11607 ) ;
 assign wire29209 = ( pg19334 ) | ( pg7916 ) | ( ng990 ) ;
 assign wire29210 = ( ng1008 ) | ( ng969 ) ;
 assign wire29216 = ( ng4975  &  ng4871 ) | ( (~ ng4899)  &  ng4871 ) | ( (~ ng4944)  &  ng4871 ) ;
 assign wire29220 = ( pg35  &  ng3462  &  (~ ng3457) ) ;
 assign wire29221 = ( ng3457  &  (~ ng3462) ) ;
 assign wire29223 = ( (~ ng23112)  &  wire29221 ) | ( pg35  &  ng3466  &  ng23112 ) ;
 assign wire29224 = ( ng3333  &  pg35 ) ;
 assign wire29225 = ( pg35  &  wire7137 ) | ( pg35  &  wire7138 ) | ( pg35  &  wire28996 ) ;
 assign wire29227 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29228 = ( ng6613  &  pg35 ) ;
 assign wire29232 = ( ng5703  &  ng4349  &  ng5644  &  (~ ng4358) ) ;
 assign wire29233 = ( pg73  &  ng4332  &  ng4311 ) | ( (~ pg73)  &  (~ ng4332)  &  ng4311 ) ;
 assign wire29234 = ( ng4349  &  ng3352  &  ng3288  &  (~ ng4358) ) ;
 assign wire29235 = ( ng6741  &  ng6682  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire29236 = ( ng4349  &  ng6336  &  ng6395  &  ng4358 ) ;
 assign wire29237 = ( ng4349  &  ng4054  &  ng3990  &  ng4358 ) ;
 assign wire29238 = ( (~ ng4349)  &  ng5990  &  ng6049  &  ng4358 ) ;
 assign wire29239 = ( ng5297  &  ng5357  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire29240 = ( (~ ng4349)  &  ng3703  &  ng3639  &  ng4358 ) ;
 assign wire29245 = ( wire6946 ) | ( wire6947 ) | ( wire6948 ) | ( wire6949 ) ;
 assign wire29246 = ( wire6950 ) | ( wire6951 ) | ( wire6952 ) | ( wire6953 ) ;
 assign wire29247 = ( ng1478  &  pg35 ) ;
 assign wire29248 = ( ng1437  &  (~ ng1478) ) ;
 assign wire29250 = ( (~ pg35)  &  ng1437 ) | ( pg35  &  ng1478  &  (~ ng1437) ) ;
 assign wire29251 = ( wire29250 ) | ( ng10961  &  wire29247 ) | ( ng13861  &  wire29247 ) ;
 assign wire29253 = ( ng4785  &  ng4709  &  ng11261  &  ng10831 ) ;
 assign wire29254 = ( ng4975  &  ng4899  &  ng11283  &  ng10862 ) ;
 assign wire29255 = ( pg35  &  ng2643  &  ng2555 ) | ( pg35  &  ng2643  &  ng2629 ) ;
 assign wire29256 = ( ng26793  &  wire29255 ) | ( ng14506  &  wire29255 ) ;
 assign wire29257 = ( pg35  &  (~ ng2643) ) | ( pg35  &  (~ ng2555)  &  (~ ng2629) ) ;
 assign wire29258 = ( ng26793  &  wire29257 ) | ( ng14506  &  wire29257 ) ;
 assign wire29259 = ( ng2643  &  pg35 ) ;
 assign wire29260 = ( wire6933 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire29259 ) ;
 assign wire29263 = ( pg17291  &  (~ ng979) ) | ( pg17291  &  (~ ng1061) ) ;
 assign wire29265 = ( pg35  &  ng11893  &  ng26673 ) | ( pg35  &  ng11893  &  ng17292 ) ;
 assign wire29266 = ( ng1620  &  pg35 ) ;
 assign wire29269 = ( pg17423  &  (~ ng1322) ) | ( pg17423  &  (~ ng1404) ) ;
 assign wire29272 = ( ng504  &  ng518  &  ng528 ) ;
 assign wire29277 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29278 = ( ng5583  &  pg35 ) ;
 assign wire29280 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29281 = ( ng5244  &  pg35 ) ;
 assign wire29283 = ( pg35  &  pg12919  &  ng904  &  ng921 ) ;
 assign wire29284 = ( pg35  &  pg12919  &  ng936 ) ;
 assign wire29285 = ( (~ pg35)  &  ng921 ) | ( ng15674  &  wire29284 ) ;
 assign wire29290 = ( pg35  &  (~ ng4854)  &  ng11012 ) ;
 assign wire29292 = ( pg35  &  ng4854  &  (~ ng11012) ) ;
 assign wire29293 = ( wire6890 ) | ( ng31009  &  (~ ng10862)  &  wire29290 ) ;
 assign wire29300 = ( (~ ng1632)  &  pg35 ) ;
 assign wire29303 = ( (~ pg35)  &  ng2763 ) | ( pg35  &  ng2767  &  (~ ng12377) ) ;
 assign wire29304 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29305 = ( ng5921  &  pg35 ) ;
 assign wire29308 = ( (~ ng2783)  &  (~ ng2724) ) ;
 assign wire29309 = ( (~ ng2787)  &  ng2724 ) ;
 assign wire29312 = ( (~ ng5046)  &  (~ ng5052) ) ;
 assign wire29313 = ( (~ pg84)  &  ng5022  &  ng5057 ) ;
 assign wire29315 = ( (~ ng5046)  &  (~ ng5041) ) ;
 assign wire29316 = ( pg84  &  ng5022  &  ng5057 ) ;
 assign wire29317 = ( pg35  &  ng5052 ) | ( pg35  &  ng5046 ) | ( pg35  &  (~ wire29313) ) ;
 assign wire29320 = ( pg35  &  (~ ng979)  &  ng1061 ) ;
 assign wire29322 = ( pg35  &  (~ ng979)  &  (~ ng1061) ) ;
 assign wire29323 = ( (~ pg35)  &  ng1052 ) | ( (~ ng1052)  &  wire29320 ) | ( ng13121  &  wire29320 ) ;
 assign wire29324 = ( (~ pg7257)  &  (~ pg7243) ) ;
 assign wire29325 = ( (~ ng4411)  &  (~ ng4375) ) ;
 assign wire29326 = ( (~ pg7243)  &  (~ pg7257)  &  (~ ng4405) ) ;
 assign wire29328 = ( pg35  &  (~ ng4392)  &  ng4388 ) ;
 assign wire29329 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29330 = ( ng3610  &  pg35 ) ;
 assign wire29335 = ( ng4975  &  pg35 ) ;
 assign wire29336 = ( wire6849 ) | ( ng28349  &  ng13486  &  wire29335 ) ;
 assign wire29340 = ( (~ pg35)  &  ng4430 ) | ( (~ ng4388)  &  ng4430 ) ;
 assign wire29346 = ( ng4674  &  (~ ng4785) ) | ( ng4674  &  (~ ng4743) ) | ( ng4674  &  ng4709 ) ;
 assign wire29348 = ( ng93  &  ng4349  &  (~ ng4358)  &  ng29503 ) ;
 assign wire29350 = ( (~ ng5703)  &  pg35 ) ;
 assign wire29352 = ( ng5703  &  pg35 ) ;
 assign wire29355 = ( pg73  &  pg35 ) | ( pg72  &  pg35 ) ;
 assign wire29359 = ( (~ pg73)  &  (~ pg72)  &  pg35 ) ;
 assign wire29361 = ( wire6823 ) | ( wire6825 ) | ( ng12228  &  wire29359 ) ;
 assign wire29362 = ( ng1141  &  pg35 ) ;
 assign wire29363 = ( ng956  &  ng1146 ) | ( ng956  &  ng1099 ) ;
 assign wire29366 = ( ng1141  &  pg35 ) ;
 assign wire29367 = ( (~ ng956)  &  ng1146 ) | ( (~ ng956)  &  ng1099 ) ;
 assign wire29371 = ( pg35  &  ng956  &  (~ ng1146)  &  (~ ng1099) ) ;
 assign wire29374 = ( pg35  &  (~ ng956)  &  (~ ng1146)  &  (~ ng1099) ) ;
 assign wire29377 = ( (~ pg35)  &  ng1129 ) | ( pg35  &  ng1141  &  ng10909 ) ;
 assign wire29378 = ( (~ ng10909)  &  (~ ng13336)  &  wire29371 ) | ( (~ ng10909)  &  ng13336  &  wire29374 ) ;
 assign wire29383 = ( (~ pg35)  &  ng4504 ) | ( ng4504  &  (~ ng4581) ) ;
 assign wire29391 = ( ng291  &  pg35 ) ;
 assign wire29393 = ( (~ ng291)  &  pg35 ) ;
 assign wire29397 = ( ng424  &  (~ ng691) ) | ( (~ ng691)  &  (~ ng417) ) ;
 assign wire29402 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29403 = ( ng6267  &  pg35 ) ;
 assign wire29405 = ( pg17404  &  (~ ng1322) ) | ( pg17404  &  (~ ng1404) ) ;
 assign wire29408 = ( ng2399  &  pg35 ) ;
 assign wire29414 = ( ng20841 ) | ( ng19968 ) | ( ng20014 ) | ( ng19919 ) ;
 assign wire29415 = ( pg35  &  ng2898 ) | ( (~ pg35)  &  ng2864 ) ;
 assign wire29416 = ( ng4392  &  pg35 ) ;
 assign wire29417 = ( ng4382  &  ng4375 ) ;
 assign wire29418 = ( wire6743 ) | ( wire29325  &  wire29326  &  wire29416 ) ;
 assign wire29419 = ( ng5897  &  ng6035 ) ;
 assign wire29420 = ( (~ ng5990)  &  (~ ng6049)  &  ng6031 ) ;
 assign wire29422 = ( pg17607  &  ng5953  &  (~ ng5990)  &  (~ ng6049) ) ;
 assign wire29423 = ( ng5889  &  pg13068 ) ;
 assign wire29424 = ( ng6035  &  (~ ng5990)  &  (~ ng6049) ) ;
 assign wire29425 = ( (~ ng6035)  &  pg17819 ) ;
 assign wire29426 = ( ng5990  &  ng6049  &  ng5925 ) ;
 assign wire29428 = ( pg17739  &  ng5937  &  ng5990  &  ng6049 ) ;
 assign wire29429 = ( ng5949  &  pg17715 ) ;
 assign wire29430 = ( ng6035  &  ng5990  &  ng6049 ) ;
 assign wire29431 = ( ng6035  &  pg14673 ) ;
 assign wire29432 = ( ng5990  &  (~ ng6049)  &  ng5933 ) ;
 assign wire29433 = ( ng6035  &  pg12350 ) ;
 assign wire29434 = ( (~ ng5990)  &  ng5893  &  ng6049 ) ;
 assign wire29436 = ( pg14738  &  ng5921  &  ng5990  &  (~ ng6049) ) ;
 assign wire29437 = ( (~ ng6035)  &  pg13068 ) ;
 assign wire29438 = ( ng5901  &  ng5990  &  (~ ng6049) ) ;
 assign wire29439 = ( (~ ng6035)  &  pg17646 ) ;
 assign wire29440 = ( (~ ng5990)  &  ng6049  &  ng5905 ) ;
 assign wire29441 = ( ng5917  &  pg17819 ) ;
 assign wire29442 = ( ng6035  &  (~ ng5990)  &  ng6049 ) ;
 assign wire29443 = ( wire29419  &  wire29420 ) | ( (~ ng12351)  &  wire29422 ) ;
 assign wire29444 = ( wire29423  &  wire29424 ) | ( wire29425  &  wire29426 ) ;
 assign wire29445 = ( (~ ng12351)  &  wire29428 ) | ( wire29429  &  wire29430 ) ;
 assign wire29446 = ( wire29431  &  wire29432 ) | ( wire29433  &  wire29434 ) ;
 assign wire29447 = ( (~ ng12351)  &  wire29436 ) | ( wire29437  &  wire29438 ) ;
 assign wire29448 = ( wire29439  &  wire29440 ) | ( wire29441  &  wire29442 ) ;
 assign wire29451 = ( wire29448 ) | ( wire29447 ) ;
 assign wire29452 = ( wire29443 ) | ( wire29444 ) | ( wire29445 ) | ( wire29446 ) ;
 assign wire29453 = ( (~ ng6035)  &  pg14673 ) ;
 assign wire29454 = ( ng5941  &  (~ ng5990)  &  (~ ng6049) ) ;
 assign wire29456 = ( pg14738  &  ng5929  &  (~ ng5990)  &  (~ ng6049) ) ;
 assign wire29457 = ( (~ ng6035)  &  pg12350 ) ;
 assign wire29458 = ( ng5990  &  ng6049  &  ng5909 ) ;
 assign wire29459 = ( ng6035  &  pg17646 ) ;
 assign wire29460 = ( ng5990  &  ng6049  &  ng5965 ) ;
 assign wire29461 = ( (~ ng6035)  &  ng5913 ) ;
 assign wire29462 = ( ng5990  &  (~ ng6049)  &  ng6031 ) ;
 assign wire29464 = ( pg17607  &  ng5990  &  (~ ng6049)  &  ng5961 ) ;
 assign wire29466 = ( pg17739  &  (~ ng5990)  &  ng6049  &  ng5945 ) ;
 assign wire29467 = ( (~ ng6035)  &  pg17715 ) ;
 assign wire29468 = ( (~ ng5990)  &  ng6049  &  ng5957 ) ;
 assign wire29469 = ( wire29453  &  wire29454 ) | ( ng12351  &  wire29456 ) ;
 assign wire29470 = ( wire29457  &  wire29458 ) | ( wire29459  &  wire29460 ) ;
 assign wire29471 = ( wire29461  &  wire29462 ) | ( ng12351  &  wire29464 ) ;
 assign wire29472 = ( ng12351  &  wire29466 ) | ( wire29467  &  wire29468 ) ;
 assign wire29475 = ( wire29469 ) | ( wire29470 ) | ( wire29471 ) | ( wire29472 ) ;
 assign wire29476 = ( pg35  &  wire7351 ) | ( pg35  &  wire7352 ) | ( pg35  &  wire28734 ) ;
 assign wire29477 = ( ng4831  &  pg35 ) ;
 assign wire29480 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29481 = ( ng5889  &  pg35 ) ;
 assign wire29482 = ( wire6714 ) | ( ng10312  &  ng12609  &  wire29480 ) ;
 assign wire29484 = ( pg35  &  (~ ng822)  &  (~ ng14279) ) ;
 assign wire29486 = ( pg35  &  ng822  &  (~ ng14279) ) ;
 assign wire29489 = ( ng3873  &  ng3881  &  ng3869 ) ;
 assign wire29491 = ( (~ ng4087)  &  (~ ng4098)  &  ng4093 ) ;
 assign wire29493 = ( ng5869  &  ng5881  &  ng5873 ) ;
 assign wire29495 = ( ng4087  &  (~ ng4098)  &  (~ ng4093) ) ;
 assign wire29496 = ( ng5535  &  ng5523  &  ng5527 ) ;
 assign wire29497 = ( ng3171  &  ng3179  &  ng3167 ) ;
 assign wire29499 = ( (~ ng4087)  &  ng4098  &  ng4093 ) ;
 assign wire29500 = ( ng3530  &  ng3518  &  ng3522 ) ;
 assign wire29502 = ( (~ ng4087)  &  ng4098  &  (~ ng4093) ) ;
 assign wire29507 = ( wire6699 ) | ( wire6700 ) | ( wire6701 ) | ( wire6702 ) ;
 assign wire29508 = ( wire6703 ) | ( wire6704 ) | ( wire6705 ) | ( wire6706 ) ;
 assign wire29510 = ( pg35  &  (~ ng2102)  &  (~ ng2108) ) ;
 assign wire29511 = ( ng2108  &  ng2102 ) ;
 assign wire29512 = ( ng2112  &  pg35 ) ;
 assign wire29516 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29517 = ( ng5543  &  pg35 ) ;
 assign wire29518 = ( wire6694 ) | ( ng10281  &  ng12558  &  wire29516 ) ;
 assign wire29520 = ( (~ ng4452)  &  (~ ng4443) ) ;
 assign wire29521 = ( (~ pg7260)  &  (~ pg7245)  &  (~ ng4438) ) ;
 assign wire29522 = ( ng4438  &  ng4382 ) ;
 assign wire29523 = ( ng4392  &  pg35 ) ;
 assign wire29524 = ( wire6691 ) | ( (~ wire29520)  &  wire29522 ) | ( (~ wire29521)  &  wire29522 ) ;
 assign wire29526 = ( pg35  &  ng142  &  ng23204 ) ;
 assign wire29527 = ( (~ ng142)  &  pg35 ) ;
 assign wire29532 = ( (~ pg35)  &  ng5112 ) | ( pg35  &  (~ pg9497)  &  pg9553  &  (~ ng5112) ) ;
 assign wire29534 = ( ng1454  &  (~ ng1448) ) ;
 assign wire29535 = ( ng1448  &  pg35 ) ;
 assign wire29536 = ( (~ pg35)  &  ng1454 ) | ( pg35  &  ng1448  &  (~ ng1454) ) ;
 assign wire29537 = ( wire29536 ) | ( (~ ng13273)  &  (~ ng10961)  &  wire29534 ) ;
 assign wire29538 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29539 = ( ng3961  &  pg35 ) ;
 assign wire29541 = ( pg35  &  ng1002  &  (~ ng7567) ) | ( pg35  &  ng15737  &  (~ ng7567) ) ;
 assign wire29542 = ( ng1018  &  pg35 ) ;
 assign wire29545 = ( ng5046  &  ng5062 ) ;
 assign wire29546 = ( (~ pg84)  &  ng5052  &  (~ ng5057) ) ;
 assign wire29548 = ( ng5046  &  ng5041 ) ;
 assign wire29549 = ( pg84  &  ng5062  &  (~ ng5057) ) ;
 assign wire29550 = ( wire29545  &  wire29546 ) | ( wire29548  &  wire29549 ) ;
 assign wire29551 = ( wire29312  &  wire29313 ) | ( wire29315  &  wire29316 ) ;
 assign wire29553 = ( pg35  &  ng5029  &  (~ ng12933) ) ;
 assign wire29555 = ( (~ pg35)  &  ng5016 ) | ( pg35  &  (~ ng5029)  &  ng12933 ) ;
 assign wire29556 = ( ng513  &  pg35 ) ;
 assign wire29557 = ( ng504  &  (~ ng667) ) | ( ng504  &  ng686 ) ;
 assign wire29559 = ( (~ ng1996) ) | ( (~ ng2070) ) ;
 assign wire29560 = ( pg35  &  ng26759  &  (~ wire29559) ) | ( pg35  &  ng14438  &  (~ wire29559) ) ;
 assign wire29561 = ( ng2016  &  pg35 ) ;
 assign wire29563 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29564 = ( ng5575  &  pg35 ) ;
 assign wire29567 = ( pg35  &  ng5052  &  (~ wire29550)  &  (~ wire29551) ) ;
 assign wire29568 = ( (~ ng5052)  &  pg35 ) ;
 assign wire29571 = ( (~ ng2715)  &  ng2719  &  (~ ng2783) ) ;
 assign wire29573 = ( (~ ng1894) ) | ( (~ ng1926) ) ;
 assign wire29575 = ( pg35  &  (~ ng1988)  &  (~ ng1982) ) ;
 assign wire29577 = ( ng1992  &  pg35 ) ;
 assign wire29579 = ( ng25341  &  wire29577 ) | ( ng1988  &  ng1982  &  (~ ng25341) ) ;
 assign wire29581 = ( pg35  &  ng2902 ) | ( pg35  &  ng209 ) | ( pg35  &  (~ ng691) ) ;
 assign wire29582 = ( (~ ng4040)  &  pg16693 ) ;
 assign wire29583 = ( ng4054  &  (~ ng3990)  &  ng3905 ) ;
 assign wire29584 = ( ng3917  &  pg16955 ) ;
 assign wire29585 = ( ng4040  &  ng4054  &  (~ ng3990) ) ;
 assign wire29586 = ( ng3893  &  pg11418 ) ;
 assign wire29587 = ( ng4040  &  ng4054  &  (~ ng3990) ) ;
 assign wire29589 = ( pg16659  &  (~ ng4054)  &  ng3953  &  (~ ng3990) ) ;
 assign wire29590 = ( ng4040  &  pg14518 ) ;
 assign wire29591 = ( ng3889  &  (~ ng4054)  &  (~ ng3990) ) ;
 assign wire29592 = ( ng4040  &  ng4031 ) ;
 assign wire29593 = ( ng3897  &  (~ ng4054)  &  (~ ng3990) ) ;
 assign wire29595 = ( pg16775  &  ng3937  &  ng4054  &  ng3990 ) ;
 assign wire29596 = ( ng3925  &  pg16955 ) ;
 assign wire29597 = ( (~ ng4040)  &  ng4054  &  ng3990 ) ;
 assign wire29598 = ( ng3949  &  pg16748 ) ;
 assign wire29599 = ( ng4040  &  ng4054  &  ng3990 ) ;
 assign wire29601 = ( pg13966  &  ng3921  &  (~ ng4054)  &  ng3990 ) ;
 assign wire29602 = ( ng3933  &  pg13906 ) ;
 assign wire29604 = ( ng3901  &  pg14518 ) ;
 assign wire29606 = ( wire29582  &  wire29583 ) | ( wire29584  &  wire29585 ) ;
 assign wire29607 = ( wire29586  &  wire29587 ) | ( (~ ng11419)  &  wire29589 ) ;
 assign wire29608 = ( wire29590  &  wire29591 ) | ( wire29592  &  wire29593 ) ;
 assign wire29609 = ( (~ ng11419)  &  wire29595 ) | ( wire29596  &  wire29597 ) ;
 assign wire29610 = ( wire29598  &  wire29599 ) | ( (~ ng11419)  &  wire29601 ) ;
 assign wire29611 = ( ng4040  &  ng11255  &  wire29602 ) | ( (~ ng4040)  &  ng11255  &  wire29604 ) ;
 assign wire29614 = ( wire29611 ) | ( wire29610 ) ;
 assign wire29615 = ( wire29606 ) | ( wire29607 ) | ( wire29608 ) | ( wire29609 ) ;
 assign wire29617 = ( pg16775  &  ng4054  &  (~ ng3990)  &  ng3945 ) ;
 assign wire29618 = ( (~ ng4040)  &  pg16748 ) ;
 assign wire29619 = ( ng4054  &  ng3957  &  (~ ng3990) ) ;
 assign wire29620 = ( (~ ng4040)  &  pg13906 ) ;
 assign wire29621 = ( (~ ng4054)  &  (~ ng3990)  &  ng3941 ) ;
 assign wire29623 = ( pg13966  &  ng3929  &  (~ ng4054)  &  (~ ng3990) ) ;
 assign wire29624 = ( ng4040  &  pg16693 ) ;
 assign wire29625 = ( ng4054  &  ng3965  &  ng3990 ) ;
 assign wire29626 = ( (~ ng4040)  &  pg11418 ) ;
 assign wire29627 = ( ng4054  &  ng3990  &  ng3909 ) ;
 assign wire29629 = ( pg16659  &  ng3961  &  (~ ng4054)  &  ng3990 ) ;
 assign wire29630 = ( ng3913  &  ng4031 ) ;
 assign wire29631 = ( (~ ng4040)  &  (~ ng4054)  &  ng3990 ) ;
 assign wire29632 = ( ng11419  &  wire29617 ) | ( wire29618  &  wire29619 ) ;
 assign wire29633 = ( wire29620  &  wire29621 ) | ( ng11419  &  wire29623 ) ;
 assign wire29634 = ( wire29624  &  wire29625 ) | ( wire29626  &  wire29627 ) ;
 assign wire29635 = ( ng11419  &  wire29629 ) | ( wire29630  &  wire29631 ) ;
 assign wire29638 = ( wire29632 ) | ( wire29633 ) | ( wire29634 ) | ( wire29635 ) ;
 assign wire29639 = ( pg35  &  ng3808  &  (~ ng10756) ) ;
 assign wire29640 = ( wire7325  &  wire29639 ) | ( wire7326  &  wire29639 ) | ( wire28766  &  wire29639 ) ;
 assign wire29641 = ( pg35  &  (~ ng3808) ) | ( pg35  &  ng10756 ) ;
 assign wire29642 = ( wire7325  &  wire29641 ) | ( wire7326  &  wire29641 ) | ( wire28766  &  wire29641 ) ;
 assign wire29643 = ( ng3808  &  pg35 ) ;
 assign wire29644 = ( wire6622 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire29643 ) ;
 assign wire29646 = ( (~ ng1636) ) | ( ng1668 ) ;
 assign wire29647 = ( pg35  &  ng26673  &  (~ wire29646) ) | ( pg35  &  ng17292  &  (~ wire29646) ) ;
 assign wire29648 = ( ng1608  &  pg35 ) ;
 assign wire29652 = ( pg35  &  (~ ng5535)  &  ng5523  &  ng5527 ) ;
 assign wire29653 = ( pg35  &  ng5535  &  (~ ng5523) ) | ( pg35  &  ng5535  &  (~ ng5527) ) ;
 assign wire29657 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29658 = ( ng3203  &  pg35 ) ;
 assign wire29663 = ( pg35  &  (~ ng4633)  &  (~ ng12911) ) ;
 assign wire29665 = ( pg35  &  ng4633  &  ng12911 ) ;
 assign wire29669 = ( ng4141 ) | ( (~ ng4064) ) | ( ng4057 ) | ( ng4082 ) ;
 assign wire29670 = ( ng4145  &  pg35 ) ;
 assign wire29671 = ( ng4116  &  pg35 ) ;
 assign wire29672 = ( wire6595 ) | ( ng13806  &  (~ wire29669)  &  wire29670 ) ;
 assign wire29674 = ( pg35  &  ng298  &  ng23204 ) ;
 assign wire29675 = ( (~ ng298)  &  pg35 ) ;
 assign wire29676 = ( wire6592 ) | ( (~ ng28444)  &  wire29674 ) | ( wire28561  &  wire29674 ) ;
 assign wire29679 = ( pg35  &  (~ pg17291)  &  (~ pg17316)  &  (~ pg17400) ) ;
 assign wire29683 = ( pg35  &  (~ pg17291)  &  (~ pg17316)  &  (~ pg17400) ) ;
 assign wire29688 = ( (~ pg72)  &  pg35  &  ng4581 ) | ( pg35  &  ng4572  &  ng4581 ) ;
 assign wire29689 = ( (~ pg35)  &  ng4498 ) | ( (~ ng4581)  &  ng4498 ) | ( pg73  &  pg35  &  ng4581 ) ;
 assign wire29693 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29694 = ( ng5240  &  pg35 ) ;
 assign wire29702 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29703 = ( ng5929  &  pg35 ) ;
 assign wire29706 = ( pg35  &  ng837  &  (~ ng832) ) ;
 assign wire29708 = ( pg35  &  ng837  &  (~ ng827) ) ;
 assign wire29709 = ( ng837  &  pg35 ) ;
 assign wire29711 = ( (~ pg35)  &  ng703 ) | ( (~ ng14279)  &  wire29706 ) ;
 assign wire29712 = ( (~ ng14279)  &  wire29708 ) | ( ng8806  &  wire29709 ) ;
 assign wire29714 = ( (~ ng2465) ) | ( ng2495 ) ;
 assign wire29715 = ( pg35  &  ng26770  &  (~ wire29714) ) | ( pg35  &  ng17424  &  (~ wire29714) ) ;
 assign wire29716 = ( ng2437  &  pg35 ) ;
 assign wire29718 = ( (~ pg11678)  &  ng781 ) | ( ng781  &  ng736 ) ;
 assign wire29720 = ( pg35  &  (~ pg11678)  &  ng785 ) | ( pg35  &  ng785  &  ng736 ) ;
 assign wire29721 = ( (~ ng785)  &  pg35 ) ;
 assign wire29723 = ( (~ ng2629) ) | ( (~ ng2555) ) ;
 assign wire29724 = ( pg35  &  ng26793  &  (~ wire29723) ) | ( pg35  &  ng14506  &  (~ wire29723) ) ;
 assign wire29725 = ( ng2575  &  pg35 ) ;
 assign wire29727 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29728 = ( ng3925  &  pg35 ) ;
 assign wire29730 = ( ng4818 ) | ( wire1421 ) ;
 assign wire29731 = ( wire1421  &  ng4771 ) | ( ng4771  &  ng4818 ) | ( ng4771  &  (~ ng24374) ) ;
 assign wire29733 = ( pg35  &  ng101  &  ng24374  &  (~ wire29730) ) ;
 assign wire29735 = ( ng29719  &  wire29733 ) | ( pg35  &  ng4765  &  (~ ng29719) ) ;
 assign wire29737 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29738 = ( ng6605  &  pg35 ) ;
 assign wire29742 = ( pg35  &  (~ ng6573)  &  ng6561  &  ng6565 ) ;
 assign wire29743 = ( pg35  &  ng6573  &  (~ ng6561) ) | ( pg35  &  ng6573  &  (~ ng6565) ) ;
 assign wire29747 = ( pg35  &  (~ ng5481)  &  (~ ng5475) ) ;
 assign wire29749 = ( pg35  &  ng5481  &  ng5475 ) ;
 assign wire29752 = ( (~ ng23630)  &  wire29749 ) | ( pg35  &  ng5485  &  ng23630 ) ;
 assign wire29753 = ( (~ ng1211)  &  pg35 ) ;
 assign wire29755 = ( ng1211  &  pg35 ) ;
 assign wire29757 = ( wire6520 ) | ( (~ ng11148)  &  (~ ng13570)  &  wire29753 ) ;
 assign wire29758 = ( ng1821  &  pg35 ) ;
 assign wire29761 = ( pg35  &  ng5120  &  (~ ng5115) ) ;
 assign wire29762 = ( ng5115  &  (~ ng5120) ) ;
 assign wire29764 = ( (~ ng23590)  &  wire29762 ) | ( pg35  &  ng5124  &  ng23590 ) ;
 assign wire29770 = ( pg35  &  (~ pg13099)  &  (~ pg14828)  &  (~ pg17722) ) ;
 assign wire29771 = ( (~ pg17778)  &  (~ pg17688) ) ;
 assign wire29775 = ( pg35  &  pg14828  &  pg12470  &  pg17722 ) ;
 assign wire29776 = ( (~ pg14828)  &  pg17778  &  pg17688 ) | ( (~ pg12470)  &  pg17778  &  pg17688 ) ;
 assign wire29780 = ( pg35  &  (~ pg13099)  &  pg14828  &  pg12470 ) ;
 assign wire29785 = ( pg35  &  (~ pg13099)  &  pg14828  &  pg12470 ) ;
 assign wire29787 = ( wire29770  &  wire29771 ) | ( wire29775  &  wire29776 ) ;
 assign wire29789 = ( (~ ng785) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire29791 = ( pg35  &  (~ pg11678)  &  ng790 ) | ( pg35  &  ng790  &  ng736 ) ;
 assign wire29792 = ( (~ ng790)  &  pg35 ) ;
 assign wire29797 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29798 = ( ng3594  &  pg35 ) ;
 assign wire29800 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29801 = ( ng5953  &  pg35 ) ;
 assign wire29804 = ( pg35  &  (~ ng6561)  &  ng6555  &  ng6549 ) ;
 assign wire29805 = ( ng2729 ) | ( (~ ng2724) ) ;
 assign wire29806 = ( (~ ng2779)  &  pg35 ) ;
 assign wire29807 = ( ng2724  &  (~ ng2729)  &  (~ ng11405)  &  wire29806 ) ;
 assign wire29809 = ( (~ ng85)  &  (~ ng11405)  &  (~ wire29805) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire29805) ) ;
 assign wire29810 = ( ng2775  &  pg35 ) ;
 assign wire29811 = ( wire6486 ) | ( ng11405  &  wire29810 ) | ( wire29805  &  wire29810 ) ;
 assign wire29812 = ( wire29811 ) | ( (~ ng85)  &  wire29807 ) | ( (~ ng29503)  &  wire29807 ) ;
 assign wire29816 = ( (~ pg135)  &  (~ ng4584)  &  (~ ng4616)  &  (~ ng4601) ) ;
 assign wire29820 = ( (~ pg135)  &  ng4584  &  (~ ng4616)  &  (~ ng4601) ) ;
 assign wire29824 = ( (~ pg135)  &  (~ ng4584)  &  (~ ng4616)  &  ng4601 ) ;
 assign wire29827 = ( ng4593  &  ng4608 ) ;
 assign wire29828 = ( (~ pg135)  &  ng4584  &  (~ ng4616)  &  ng4601 ) ;
 assign wire29830 = ( (~ ng4608)  &  (~ ng4601) ) ;
 assign wire29831 = ( (~ pg135)  &  ng4584  &  ng4593 ) ;
 assign wire29834 = ( wire6482 ) | ( (~ ng4608)  &  (~ ng4593)  &  wire29816 ) ;
 assign wire29835 = ( ng4608  &  (~ ng4593)  &  wire29820 ) | ( (~ ng4608)  &  ng4593  &  wire29824 ) ;
 assign wire29836 = ( wire29827  &  wire29828 ) | ( wire29830  &  wire29831 ) ;
 assign wire29841 = ( pg35  &  ng5022  &  (~ ng5016) ) | ( pg35  &  (~ ng5016)  &  ng5062 ) ;
 assign wire29843 = ( (~ pg35)  &  ng5022 ) | ( pg35  &  (~ ng5022)  &  ng5016  &  (~ ng5062) ) ;
 assign wire29848 = ( pg124  &  pg35  &  ng4146 ) | ( pg120  &  pg35  &  (~ ng4146) ) ;
 assign wire29849 = ( (~ pg120)  &  (~ pg124)  &  pg35 ) | ( (~ pg124)  &  pg35  &  ng4146 ) | ( (~ pg120)  &  pg35  &  (~ ng4146) ) ;
 assign wire29850 = ( pg116  &  pg35  &  ng4157 ) | ( pg114  &  pg35  &  (~ ng4157) ) ;
 assign wire29851 = ( (~ pg116)  &  (~ pg114)  &  pg35 ) | ( (~ pg116)  &  pg35  &  ng4157 ) | ( (~ pg114)  &  pg35  &  (~ ng4157) ) ;
 assign wire29852 = ( (~ pg35)  &  ng4122 ) | ( (~ ng26212)  &  wire29848 ) ;
 assign wire29853 = ( ng26212  &  wire29849 ) | ( (~ ng26256)  &  wire29850 ) ;
 assign wire29855 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29856 = ( ng3239  &  pg35 ) ;
 assign wire29858 = ( ng1478  &  pg35 ) ;
 assign wire29859 = ( ng1437  &  ng1442 ) | ( ng1437  &  ng1489 ) ;
 assign wire29862 = ( (~ ng1478)  &  pg35 ) ;
 assign wire29863 = ( ng1437  &  ng1442 ) | ( ng1437  &  ng1489 ) ;
 assign wire29867 = ( pg35  &  ng1478  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire29870 = ( pg35  &  (~ ng1478)  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire29873 = ( (~ pg35)  &  ng1442 ) | ( pg35  &  ng1437  &  ng13861 ) ;
 assign wire29874 = ( (~ ng13378)  &  (~ ng13861)  &  wire29867 ) | ( ng13378  &  (~ ng13861)  &  wire29870 ) ;
 assign wire29883 = ( (~ ng2729) ) | ( (~ ng2724) ) ;
 assign wire29884 = ( (~ ng2827)  &  pg35 ) ;
 assign wire29885 = ( ng2724  &  ng2729  &  (~ ng11405)  &  wire29884 ) ;
 assign wire29887 = ( (~ ng111)  &  (~ ng11405)  &  (~ wire29883) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire29883) ) ;
 assign wire29888 = ( ng2819  &  pg35 ) ;
 assign wire29889 = ( wire6436 ) | ( ng11405  &  wire29888 ) | ( wire29883  &  wire29888 ) ;
 assign wire29890 = ( wire29889 ) | ( (~ ng111)  &  wire29885 ) | ( (~ ng29503)  &  wire29885 ) ;
 assign wire29894 = ( (~ pg35)  &  ng3100 ) | ( pg35  &  pg8215  &  (~ pg8277)  &  (~ ng3100) ) ;
 assign wire29899 = ( pg72  &  pg35  &  ng4581 ) | ( pg35  &  ng4572  &  ng4581 ) ;
 assign wire29900 = ( (~ pg35)  &  ng4480 ) | ( (~ ng4581)  &  ng4480 ) | ( (~ pg73)  &  pg35  &  ng4581 ) ;
 assign wire29901 = ( pg7916  &  (~ ng1171)  &  ng1183 ) ;
 assign wire29902 = ( (~ ng1070)  &  pg35 ) ;
 assign wire29903 = ( ng1199  &  (~ ng10893)  &  wire29901  &  wire29902 ) ;
 assign wire29904 = ( ng1070  &  pg35 ) ;
 assign wire29905 = ( (~ ng1199)  &  wire29904 ) | ( ng10893  &  wire29904 ) | ( (~ wire29901)  &  wire29904 ) ;
 assign wire29907 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire29908 = ( ng6251  &  pg35 ) ;
 assign wire29912 = ( pg35  &  (~ ng6533)  &  (~ ng6527) ) ;
 assign wire29914 = ( pg35  &  ng6533  &  ng6527 ) ;
 assign wire29917 = ( ng10887  &  wire29914 ) | ( pg35  &  ng6537  &  (~ ng10887) ) ;
 assign wire29918 = ( ng4616  &  ng4584 ) ;
 assign wire29919 = ( ng4584  &  pg35 ) ;
 assign wire29920 = ( ng10511  &  wire29919 ) | ( ng8347  &  wire29919 ) | ( wire28475  &  wire29919 ) ;
 assign wire29921 = ( (~ ng4584)  &  pg35 ) ;
 assign wire29922 = ( (~ ng10511)  &  (~ ng8347)  &  (~ wire28475)  &  wire29921 ) ;
 assign wire29923 = ( wire6407 ) | ( (~ ng30583)  &  (~ wire6408)  &  wire29920 ) ;
 assign wire29925 = ( (~ pg53)  &  pg54 ) ;
 assign wire29926 = ( (~ pg56)  &  (~ pg57)  &  (~ ng34) ) ;
 assign wire29928 = ( ng28  &  (~ ng31) ) ;
 assign wire29930 = ( ng9  &  ng19  &  (~ ng16) ) ;
 assign wire29932 = ( ng28  &  ng31 ) ;
 assign wire29934 = ( (~ ng9)  &  (~ ng19)  &  ng16 ) ;
 assign wire29936 = ( ng9  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29937 = ( ng28  &  (~ ng31) ) ;
 assign wire29939 = ( ng9  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29941 = ( (~ ng9)  &  (~ ng19)  &  ng16 ) ;
 assign wire29942 = ( (~ ng28)  &  (~ ng31) ) ;
 assign wire29944 = ( ng9  &  (~ ng19)  &  ng16 ) ;
 assign wire29946 = ( ng9  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29948 = ( ng17725  &  wire29925  &  wire29926 ) | ( ng16283  &  wire29925  &  wire29926 ) ;
 assign wire29949 = ( ng16194  &  wire29925  &  wire29926 ) | ( ng16539  &  wire29925  &  wire29926 ) ;
 assign wire29950 = ( ng27511  &  ng16244 ) | ( ng27511  &  ng16205 ) | ( ng27511  &  ng16486 ) ;
 assign wire29952 = ( ng94  &  ng13156  &  wire29932  &  wire29934 ) ;
 assign wire29953 = ( ng2965  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire29954 = ( ng2960  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire29955 = ( ng2878  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire29956 = ( ng2873  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire29957 = ( (~ ng28)  &  (~ ng31) ) ;
 assign wire29959 = ( ng9  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29961 = ( ng9  &  ng19  &  (~ ng16) ) ;
 assign wire29962 = ( pg54  &  (~ pg53)  &  wire29926  &  wire29961 ) ;
 assign wire29963 = ( (~ ng28)  &  ng31 ) ;
 assign wire29965 = ( ng9  &  ng19  &  (~ ng16) ) ;
 assign wire29966 = ( pg54  &  (~ pg53)  &  wire29926  &  wire29965 ) ;
 assign wire29968 = ( wire7545 ) | ( wire7546 ) | ( wire7547 ) ;
 assign wire29971 = ( wire7544 ) | ( wire7543 ) ;
 assign wire29972 = ( wire7540 ) | ( wire7541 ) | ( wire7542 ) | ( wire29968 ) ;
 assign wire29974 = ( (~ ng9)  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29976 = ( (~ ng9)  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29978 = ( (~ ng9)  &  ng19  &  (~ ng16) ) ;
 assign wire29980 = ( (~ ng9)  &  (~ ng19)  &  (~ ng16) ) ;
 assign wire29982 = ( (~ ng9)  &  ng19  &  (~ ng16) ) ;
 assign wire29984 = ( ng17613  &  wire29925  &  wire29926 ) | ( ng17747  &  wire29925  &  wire29926 ) ;
 assign wire29985 = ( ng27511  &  ng17766 ) | ( ng27511  &  ng17724 ) | ( ng27511  &  ng17690 ) ;
 assign wire29986 = ( ng790  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire29987 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire29988 = ( ng572  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire29989 = ( ng749  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire29990 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire29991 = ( (~ ng550)  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire29992 = ( ng608  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire29993 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire29994 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire29996 = ( ng9  &  ng19  &  (~ ng16) ) ;
 assign wire29997 = ( pg54  &  (~ pg53)  &  wire29926  &  wire29996 ) ;
 assign wire29999 = ( (~ ng9)  &  ng19  &  (~ ng16) ) ;
 assign wire30000 = ( pg54  &  (~ pg53)  &  wire29926  &  wire29999 ) ;
 assign wire30002 = ( (~ ng9)  &  (~ ng19)  &  ng16 ) ;
 assign wire30003 = ( pg54  &  (~ pg53)  &  wire29926  &  wire30002 ) ;
 assign wire30004 = ( wire7531 ) | ( ng4253  &  ni17529  &  wire29997 ) ;
 assign wire30006 = ( wire7532 ) | ( wire7533 ) | ( wire30004 ) ;
 assign wire30008 = ( wire29984  &  wire29987 ) | ( wire29985  &  wire29987 ) | ( wire29984  &  wire29988 ) | ( wire29985  &  wire29988 ) ;
 assign wire30009 = ( wire29984  &  wire29989 ) | ( wire29985  &  wire29989 ) | ( wire29984  &  wire29990 ) | ( wire29985  &  wire29990 ) ;
 assign wire30010 = ( wire29984  &  wire29991 ) | ( wire29985  &  wire29991 ) | ( wire29984  &  wire29992 ) | ( wire29985  &  wire29992 ) ;
 assign wire30011 = ( wire29984  &  wire29993 ) | ( wire29985  &  wire29993 ) | ( wire29984  &  wire29994 ) | ( wire29985  &  wire29994 ) ;
 assign wire30013 = ( wire30010 ) | ( wire30009 ) ;
 assign wire30014 = ( wire7521 ) | ( wire30006 ) | ( wire30008 ) | ( wire30011 ) ;
 assign wire30016 = ( ng794  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30017 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30018 = ( ng534  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30019 = ( ng758  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30020 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30021 = ( ng586  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30022 = ( ng613  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30023 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30024 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30025 = ( wire7518 ) | ( ng947  &  ni17529  &  wire30000 ) ;
 assign wire30026 = ( wire30025 ) | ( ng1291  &  ni18740  &  wire30003 ) ;
 assign wire30028 = ( wire29984  &  wire30017 ) | ( wire29985  &  wire30017 ) | ( wire29984  &  wire30018 ) | ( wire29985  &  wire30018 ) ;
 assign wire30029 = ( wire29984  &  wire30019 ) | ( wire29985  &  wire30019 ) | ( wire29984  &  wire30020 ) | ( wire29985  &  wire30020 ) ;
 assign wire30030 = ( wire29984  &  wire30021 ) | ( wire29985  &  wire30021 ) | ( wire29984  &  wire30022 ) | ( wire29985  &  wire30022 ) ;
 assign wire30031 = ( wire29984  &  wire30023 ) | ( wire29985  &  wire30023 ) | ( wire29984  &  wire30024 ) | ( wire29985  &  wire30024 ) ;
 assign wire30033 = ( wire30030 ) | ( wire30029 ) ;
 assign wire30034 = ( wire7509 ) | ( wire30026 ) | ( wire30028 ) | ( wire30031 ) ;
 assign wire30035 = ( ng37  &  ng13156  &  wire29932  &  wire29934 ) ;
 assign wire30036 = ( ng2950  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30037 = ( ng2882  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30038 = ( ng2868  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30039 = ( ng2955  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30041 = ( (~ ng9)  &  ng19  &  ng16 ) ;
 assign wire30042 = ( pg54  &  (~ pg53)  &  wire29926  &  wire30041 ) ;
 assign wire30044 = ( (~ ng9)  &  ng19  &  ng16 ) ;
 assign wire30045 = ( pg54  &  (~ pg53)  &  wire29926  &  wire30044 ) ;
 assign wire30048 = ( wire7503 ) | ( wire7505 ) | ( wire7506 ) | ( wire7507 ) ;
 assign wire30052 = ( wire7498 ) | ( wire7504 ) | ( wire30048 ) ;
 assign wire30053 = ( wire7499 ) | ( wire7500 ) | ( wire7501 ) | ( wire7502 ) ;
 assign wire30055 = ( pg100  &  ng13156  &  wire29932  &  wire29934 ) ;
 assign wire30056 = ( ng2890  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30057 = ( ng2984  &  ng14988  &  wire29942  &  wire29944 ) ;
 assign wire30059 = ( wire7493 ) | ( wire7494 ) | ( wire7495 ) ;
 assign wire30061 = ( wire7491 ) | ( wire7490 ) ;
 assign wire30062 = ( wire7489 ) | ( wire7492 ) | ( wire30059 ) ;
 assign wire30063 = ( ng781  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30064 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30065 = ( ng562  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30066 = ( ng739  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30067 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30068 = ( ng199  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30069 = ( ng599  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30070 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30071 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30072 = ( wire7486 ) | ( ng4245  &  ni17529  &  wire29997 ) ;
 assign wire30074 = ( wire7485 ) | ( wire7487 ) | ( wire30072 ) ;
 assign wire30076 = ( wire29984  &  wire30064 ) | ( wire29985  &  wire30064 ) | ( wire29984  &  wire30065 ) | ( wire29985  &  wire30065 ) ;
 assign wire30077 = ( wire29984  &  wire30066 ) | ( wire29985  &  wire30066 ) | ( wire29984  &  wire30067 ) | ( wire29985  &  wire30067 ) ;
 assign wire30078 = ( wire29984  &  wire30068 ) | ( wire29985  &  wire30068 ) | ( wire29984  &  wire30069 ) | ( wire29985  &  wire30069 ) ;
 assign wire30079 = ( wire29984  &  wire30070 ) | ( wire29985  &  wire30070 ) | ( wire29984  &  wire30071 ) | ( wire29985  &  wire30071 ) ;
 assign wire30081 = ( wire30078 ) | ( wire30077 ) ;
 assign wire30082 = ( wire7475 ) | ( wire30074 ) | ( wire30076 ) | ( wire30079 ) ;
 assign wire30084 = ( ng2886  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30085 = ( pg92  &  ng13156  &  wire29932  &  wire29934 ) ;
 assign wire30086 = ( ng2970  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30087 = ( pg127  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30088 = ( ng2980  &  ng14988  &  wire29942  &  wire29944 ) ;
 assign wire30089 = ( ng2975  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30091 = ( wire7472 ) | ( wire7473 ) | ( wire7474 ) ;
 assign wire30095 = ( wire7466 ) | ( wire7471 ) | ( wire30091 ) ;
 assign wire30096 = ( wire7467 ) | ( wire7468 ) | ( wire7469 ) | ( wire7470 ) ;
 assign wire30097 = ( ng785  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30098 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30099 = ( ng744  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30100 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30101 = ( ng568  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30102 = ( ng604  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30103 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30104 = ( ng136  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30105 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30106 = ( wire7462 ) | ( ng4249  &  ni17529  &  wire29997 ) ;
 assign wire30108 = ( wire7463 ) | ( wire7464 ) | ( wire30106 ) ;
 assign wire30110 = ( wire29984  &  wire30098 ) | ( wire29985  &  wire30098 ) | ( wire29984  &  wire30099 ) | ( wire29985  &  wire30099 ) ;
 assign wire30111 = ( wire29984  &  wire30100 ) | ( wire29985  &  wire30100 ) | ( wire29984  &  wire30101 ) | ( wire29985  &  wire30101 ) ;
 assign wire30112 = ( wire29984  &  wire30102 ) | ( wire29985  &  wire30102 ) | ( wire29984  &  wire30103 ) | ( wire29985  &  wire30103 ) ;
 assign wire30113 = ( wire29984  &  wire30104 ) | ( wire29985  &  wire30104 ) | ( wire29984  &  wire30105 ) | ( wire29985  &  wire30105 ) ;
 assign wire30115 = ( wire30112 ) | ( wire30111 ) ;
 assign wire30116 = ( wire7452 ) | ( wire30108 ) | ( wire30110 ) | ( wire30113 ) ;
 assign wire30118 = ( ng807  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30119 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30120 = ( ng763  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30121 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30122 = ( ng542  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30123 = ( ng617  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30124 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30125 = ( ng577  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30126 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30127 = ( wire7424 ) | ( ni18740  &  ng10948  &  wire30003 ) ;
 assign wire30128 = ( wire30127 ) | ( ni17529  &  ng10878  &  wire30000 ) ;
 assign wire30130 = ( wire29984  &  wire30119 ) | ( wire29985  &  wire30119 ) | ( wire29984  &  wire30120 ) | ( wire29985  &  wire30120 ) ;
 assign wire30131 = ( wire29984  &  wire30121 ) | ( wire29985  &  wire30121 ) | ( wire29984  &  wire30122 ) | ( wire29985  &  wire30122 ) ;
 assign wire30132 = ( wire29984  &  wire30123 ) | ( wire29985  &  wire30123 ) | ( wire29984  &  wire30124 ) | ( wire29985  &  wire30124 ) ;
 assign wire30133 = ( wire29984  &  wire30125 ) | ( wire29985  &  wire30125 ) | ( wire29984  &  wire30126 ) | ( wire29985  &  wire30126 ) ;
 assign wire30135 = ( wire30132 ) | ( wire30131 ) ;
 assign wire30136 = ( wire7414 ) | ( wire30128 ) | ( wire30130 ) | ( wire30133 ) ;
 assign wire30137 = ( ng2936  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30138 = ( ng2894  &  ng13156  &  wire29957  &  wire29959 ) ;
 assign wire30139 = ( ng2988  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30140 = ( ng2898  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30141 = ( ng2941  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30144 = ( wire7409 ) | ( wire7410 ) | ( wire7411 ) | ( wire7412 ) ;
 assign wire30146 = ( ng31070  &  wire30138 ) | ( ng31070  &  wire30139 ) ;
 assign wire30147 = ( ng31070  &  wire30140 ) | ( ng31070  &  wire30141 ) ;
 assign wire30148 = ( wire30144 ) | ( ng31070  &  ng16486 ) | ( ng31070  &  wire30137 ) ;
 assign wire30150 = ( wire30146 ) | ( wire30147 ) | ( wire30148 ) ;
 assign wire30151 = ( ng2860  &  ng13156  &  wire29957  &  wire29959 ) ;
 assign wire30152 = ( ng2864  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30153 = ( ng2922  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30154 = ( (~ ng2994)  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30155 = ( ng2927  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30157 = ( wire7445 ) | ( wire7446 ) | ( wire7447 ) ;
 assign wire30158 = ( wire30157 ) | ( ng31070  &  wire30151 ) ;
 assign wire30159 = ( ng31070  &  wire30152 ) | ( ng31070  &  wire30153 ) ;
 assign wire30160 = ( ng31070  &  wire30154 ) | ( ng31070  &  wire30155 ) ;
 assign wire30162 = ( ng554  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30163 = ( (~ pg35)  &  ng13156  &  wire29937  &  wire29974 ) ;
 assign wire30164 = ( ng767  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30165 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30166 = ( ng622  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30167 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30168 = ( ng582  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30169 = ( ng546  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30170 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30171 = ( wire7436 ) | ( ni17529  &  ng10890  &  wire30000 ) ;
 assign wire30173 = ( wire7437 ) | ( wire7438 ) | ( wire30171 ) ;
 assign wire30175 = ( wire29984  &  wire30163 ) | ( wire29985  &  wire30163 ) | ( wire29984  &  wire30164 ) | ( wire29985  &  wire30164 ) ;
 assign wire30176 = ( wire29984  &  wire30165 ) | ( wire29985  &  wire30165 ) | ( wire29984  &  wire30166 ) | ( wire29985  &  wire30166 ) ;
 assign wire30177 = ( wire29984  &  wire30167 ) | ( wire29985  &  wire30167 ) | ( wire29984  &  wire30168 ) | ( wire29985  &  wire30168 ) ;
 assign wire30178 = ( wire29984  &  wire30169 ) | ( wire29985  &  wire30169 ) | ( wire29984  &  wire30170 ) | ( wire29985  &  wire30170 ) ;
 assign wire30180 = ( wire30177 ) | ( wire30176 ) ;
 assign wire30181 = ( wire7426 ) | ( wire30173 ) | ( wire30175 ) | ( wire30178 ) ;
 assign wire30182 = ( wire30176 ) | ( wire30177 ) | ( wire30181 ) ;
 assign wire30183 = ( ng2917  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30184 = ( ng772  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30185 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30186 = ( ng2852  &  ng13156  &  wire29957  &  wire29959 ) ;
 assign wire30187 = ( ng2912  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30188 = ( ng2856  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30189 = ( ng2999  &  ng13156  &  wire29937  &  wire29941 ) ;
 assign wire30190 = ( (~ ng590)  &  pg35 ) ;
 assign wire30193 = ( wire7378 ) | ( pg35  &  (~ ng626)  &  (~ ng590) ) ;
 assign wire30194 = ( (~ ng17766)  &  (~ ng17747) ) | ( pg35  &  (~ ng626)  &  (~ ng17766) ) ;
 assign wire30195 = ( wire7372 ) | ( ng3502  &  ni18785  &  wire29966 ) ;
 assign wire30199 = ( wire7373 ) | ( wire7374 ) | ( wire7375 ) | ( wire7376 ) ;
 assign wire30201 = ( wire29984  &  wire30184 ) | ( wire29985  &  wire30184 ) | ( wire29984  &  wire30185 ) | ( wire29985  &  wire30185 ) ;
 assign wire30202 = ( wire7371 ) | ( wire7377 ) | ( wire30195 ) | ( wire30199 ) ;
 assign wire30203 = ( ng31070  &  wire30183 ) | ( ng31070  &  wire30186 ) ;
 assign wire30204 = ( ng31070  &  wire30187 ) | ( ng31070  &  wire30188 ) ;
 assign wire30205 = ( wire30201 ) | ( ng31070  &  wire30189 ) ;
 assign wire30208 = ( ng2848  &  ng13156  &  wire29937  &  wire29939 ) ;
 assign wire30209 = ( ng2844  &  ng13156  &  wire29957  &  wire29959 ) ;
 assign wire30210 = ( ng2907  &  ng14988  &  wire29928  &  wire29936 ) ;
 assign wire30211 = ( ng2902  &  ng14988  &  wire29942  &  wire29946 ) ;
 assign wire30213 = ( wire7398 ) | ( wire7399 ) | ( wire7400 ) ;
 assign wire30215 = ( ng31070  &  wire30209 ) | ( ng31070  &  wire30210 ) ;
 assign wire30216 = ( wire30213 ) | ( ng31070  &  wire30208 ) | ( ng31070  &  wire30211 ) ;
 assign wire30217 = ( ng776  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30218 = ( (~ pg35)  &  ng13156  &  wire29932  &  wire29976 ) ;
 assign wire30219 = ( ng632  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30220 = ( ng595  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30221 = ( ng538  &  ng13156  &  wire29957  &  wire29980 ) ;
 assign wire30222 = ( (~ pg35)  &  ng13156  &  wire29957  &  wire29978 ) ;
 assign wire30223 = ( (~ pg35)  &  ng13156  &  wire29963  &  wire29982 ) ;
 assign wire30224 = ( wire7391 ) | ( ng10925  &  ni17529  &  wire30000 ) ;
 assign wire30226 = ( wire7390 ) | ( wire7392 ) | ( wire30224 ) ;
 assign wire30228 = ( wire29984  &  wire30218 ) | ( wire29985  &  wire30218 ) | ( wire29984  &  wire30219 ) | ( wire29985  &  wire30219 ) ;
 assign wire30229 = ( wire29984  &  wire30220 ) | ( wire29985  &  wire30220 ) | ( wire29984  &  wire30221 ) | ( wire29985  &  wire30221 ) ;
 assign wire30230 = ( wire29984  &  wire30222 ) | ( wire29985  &  wire30222 ) | ( wire29984  &  wire30223 ) | ( wire29985  &  wire30223 ) ;
 assign wire30231 = ( wire7382 ) | ( wire30226 ) | ( wire30228 ) ;
 assign wire30232 = ( wire30230 ) | ( wire30229 ) ;
 assign wire30236 = ( (~ pg56)  &  (~ pg54)  &  pg35  &  (~ pg53) ) ;
 assign wire30237 = ( pg35  &  ng2984 ) | ( (~ pg35)  &  ng2980 ) ;
 assign wire30238 = ( ng1351 ) | ( ng1312 ) ;
 assign wire30241 = ( pg35  &  (~ pg17320)  &  (~ pg17423)  &  (~ pg17404) ) ;
 assign wire30245 = ( pg35  &  (~ pg17320)  &  (~ pg17423)  &  (~ pg17404) ) ;
 assign wire30249 = ( (~ ng2287) ) | ( (~ ng2361) ) ;
 assign wire30250 = ( pg35  &  ng17405  &  (~ wire30249) ) | ( pg35  &  ng26737  &  (~ wire30249) ) ;
 assign wire30251 = ( ng2307  &  pg35 ) ;
 assign wire30254 = ( pg35  &  ng3703  &  (~ ng3639)  &  (~ ng3698) ) ;
 assign wire30255 = ( ng4975  &  (~ ng4899)  &  ng11283  &  wire30254 ) ;
 assign wire30257 = ( pg35  &  (~ ng3703)  &  (~ ng3694)  &  (~ ng3639) ) ;
 assign wire30258 = ( ng4975  &  (~ ng4899)  &  ng11283  &  wire30257 ) ;
 assign wire30260 = ( pg35  &  ng3703  &  ng3639  &  ng3698 ) ;
 assign wire30261 = ( ng4975  &  (~ ng4899)  &  ng11283  &  wire30260 ) ;
 assign wire30263 = ( pg35  &  (~ ng3703)  &  ng3694  &  ng3639 ) ;
 assign wire30264 = ( ng4975  &  (~ ng4899)  &  ng11283  &  wire30263 ) ;
 assign wire30265 = ( ng4950  &  pg35 ) ;
 assign wire30267 = ( wire6373 ) | ( ng21024  &  wire30258 ) ;
 assign wire30268 = ( ng21024  &  wire30264 ) | ( pg35  &  ng4950  &  (~ ng21024) ) ;
 assign wire30269 = ( (~ ng23309)  &  wire30255 ) | ( (~ ng23309)  &  wire30261 ) ;
 assign wire30272 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30273 = ( ng5216  &  pg35 ) ;
 assign wire30274 = ( wire6368 ) | ( ng12443  &  ng12492  &  wire30272 ) ;
 assign wire30276 = ( ng504  &  ng518  &  (~ ng528) ) ;
 assign wire30281 = ( ng1668  &  pg35 ) ;
 assign wire30283 = ( (~ ng504)  &  (~ ng518)  &  (~ ng528) ) ;
 assign wire30286 = ( wire6362 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire30281 ) ;
 assign wire30293 = ( pg35  &  (~ ng827)  &  (~ ng14279) ) ;
 assign wire30295 = ( pg35  &  ng827  &  (~ ng14279) ) ;
 assign wire30300 = ( ng1274  &  (~ ng1536) ) | ( (~ ng1312)  &  ng1274  &  (~ ng1351) ) ;
 assign wire30301 = ( (~ ng2193)  &  pg35 ) ;
 assign wire30304 = ( (~ pg35)  &  ng121 ) | ( pg35  &  ng2799  &  (~ ng12377) ) ;
 assign wire30307 = ( pg35  &  (~ ng1926)  &  ng1882  &  (~ ng1894) ) ;
 assign wire30310 = ( pg35  &  (~ ng1917)  &  ng1894  &  ng1886 ) ;
 assign wire30312 = ( pg35  &  ng1870  &  ng1917  &  (~ ng1894) ) ;
 assign wire30313 = ( ng1926  &  ng1878  &  (~ ng1917) ) ;
 assign wire30314 = ( (~ ng1917) ) | ( ng1926 ) ;
 assign wire30315 = ( ng1890  &  pg35 ) ;
 assign wire30316 = ( ng1945  &  pg35 ) ;
 assign wire30320 = ( ng1874  &  (~ ng25341) ) | ( (~ ng25429)  &  wire30315 ) ;
 assign wire30321 = ( wire6330 ) | ( wire6331 ) | ( wire6332 ) | ( wire6336 ) ;
 assign wire30324 = ( pg35  &  (~ pg11678)  &  ng776 ) | ( pg35  &  ng776  &  ng736 ) ;
 assign wire30325 = ( (~ ng776)  &  pg35 ) ;
 assign wire30327 = ( (~ ng599) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire30328 = ( (~ pg9048)  &  ng604 ) | ( ng604  &  ng559 ) ;
 assign wire30329 = ( (~ ng608) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire30330 = ( (~ pg9048)  &  ng613 ) | ( ng559  &  ng613 ) ;
 assign wire30331 = ( (~ ng617) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire30332 = ( (~ pg9048)  &  ng622 ) | ( ng559  &  ng622 ) ;
 assign wire30334 = ( pg35  &  (~ pg9048)  &  ng626 ) | ( pg35  &  ng626  &  ng559 ) ;
 assign wire30335 = ( (~ ng626)  &  pg35 ) ;
 assign wire30337 = ( (~ ng4340)  &  pg35 ) ;
 assign wire30339 = ( pg35  &  ng65  &  ng29503 ) | ( pg35  &  ng65  &  ng27972 ) ;
 assign wire30341 = ( ng31971  &  wire30339 ) | ( pg35  &  ng4340  &  (~ ng31971) ) ;
 assign wire30342 = ( ng2715  &  ng2719  &  (~ ng2787) ) ;
 assign wire30343 = ( ng2060 ) | ( (~ ng2051) ) ;
 assign wire30344 = ( (~ ng2040)  &  pg35 ) ;
 assign wire30348 = ( pg35  &  ng2036  &  ng25470 ) | ( pg35  &  ng1996  &  (~ ng25470) ) ;
 assign wire30349 = ( (~ ng2028) ) | ( (~ ng2060) ) ;
 assign wire30356 = ( ng504  &  (~ ng518)  &  ng528 ) ;
 assign wire30359 = ( pg35  &  ng2361  &  (~ ng112)  &  (~ ng2331) ) ;
 assign wire30361 = ( pg35  &  (~ ng2361)  &  ng112 ) | ( pg35  &  ng112  &  ng2331 ) ;
 assign wire30362 = ( ng2338  &  pg35 ) ;
 assign wire30365 = ( (~ ng4349)  &  (~ ng4358)  &  (~ ng24380)  &  wire29233 ) ;
 assign wire30367 = ( (~ ng6741)  &  pg35 ) ;
 assign wire30369 = ( ng6741  &  pg35 ) ;
 assign wire30372 = ( pg35  &  (~ ng6500)  &  ng6505 ) ;
 assign wire30373 = ( (~ ng6505)  &  ng6500 ) ;
 assign wire30375 = ( (~ ng23733)  &  wire30373 ) | ( pg35  &  ng6509  &  ng23733 ) ;
 assign wire30377 = ( (~ ng504)  &  ng518  &  (~ ng528) ) ;
 assign wire30382 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30383 = ( ng5563  &  pg35 ) ;
 assign wire30384 = ( wire6293 ) | ( ng12505  &  ng12558  &  wire30382 ) ;
 assign wire30386 = ( (~ ng4474) ) | ( ng4477 ) ;
 assign wire30388 = ( pg35  &  ng4459 ) | ( (~ pg35)  &  ng4369 ) ;
 assign wire30390 = ( (~ ng2465) ) | ( ng2421 ) ;
 assign wire30391 = ( pg35  &  ng26770  &  (~ wire30390) ) | ( pg35  &  ng17424  &  (~ wire30390) ) ;
 assign wire30392 = ( ng2445  &  pg35 ) ;
 assign wire30394 = ( (~ ng2407)  &  pg35 ) ;
 assign wire30395 = ( ng2407  &  pg35 ) ;
 assign wire30399 = ( pg35  &  (~ ng1624)  &  (~ ng1657)  &  ng1612 ) ;
 assign wire30402 = ( pg35  &  ng1624  &  ng1616  &  (~ ng1648) ) ;
 assign wire30404 = ( pg35  &  (~ ng1624)  &  ng1648  &  ng1600 ) ;
 assign wire30405 = ( ng1620  &  pg35 ) ;
 assign wire30406 = ( ng1608  &  ng1657  &  (~ ng1648) ) ;
 assign wire30407 = ( ng1677  &  pg35 ) ;
 assign wire30411 = ( ng1604  &  (~ ng25275) ) | ( (~ ng25337)  &  wire30405 ) ;
 assign wire30412 = ( wire6269 ) | ( wire6270 ) | ( wire6271 ) | ( wire6276 ) ;
 assign wire30417 = ( (~ ng2595)  &  pg35 ) ;
 assign wire30420 = ( (~ pg35)  &  ng2823 ) | ( pg35  &  ng2827  &  (~ ng12377) ) ;
 assign wire30421 = ( ng1339  &  pg35 ) ;
 assign wire30422 = ( ng1306  &  pg35 ) ;
 assign wire30427 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30428 = ( ng3219  &  pg35 ) ;
 assign wire30430 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30431 = ( ng6597  &  pg35 ) ;
 assign wire30433 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30434 = ( ng5913  &  pg35 ) ;
 assign wire30436 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30437 = ( ng3259  &  pg35 ) ;
 assign wire30441 = ( pg35  &  ng2495  &  (~ ng112)  &  (~ ng2465) ) ;
 assign wire30443 = ( pg35  &  (~ ng2495)  &  ng112 ) | ( pg35  &  ng112  &  ng2465 ) ;
 assign wire30444 = ( ng2472  &  pg35 ) ;
 assign wire30447 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30448 = ( ng3195  &  pg35 ) ;
 assign wire30453 = ( (~ pg35)  &  ng3451 ) | ( pg35  &  (~ pg8342)  &  pg8279  &  (~ ng3451) ) ;
 assign wire30457 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30458 = ( ng3211  &  pg35 ) ;
 assign wire30464 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30465 = ( ng3191  &  pg35 ) ;
 assign wire30466 = ( wire6217 ) | ( ng11514  &  ng11729  &  wire30464 ) ;
 assign wire30467 = ( (~ ng2453) ) | ( (~ ng2485) ) ;
 assign wire30471 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30472 = ( ng3243  &  pg35 ) ;
 assign wire30474 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30475 = ( ng5204  &  pg35 ) ;
 assign wire30477 = ( (~ ng1906) ) | ( ng1862 ) ;
 assign wire30478 = ( (~ ng1936)  &  pg35 ) ;
 assign wire30480 = ( ng26725  &  (~ ng28789)  &  wire30478 ) | ( ng17401  &  (~ ng28789)  &  wire30478 ) ;
 assign wire30484 = ( (~ pg35)  &  ng1183 ) | ( pg35  &  (~ pg7916)  &  ng1178 ) ;
 assign wire30487 = ( pg35  &  (~ ng3530)  &  ng3518  &  ng3522 ) ;
 assign wire30488 = ( pg35  &  ng3530  &  (~ ng3518) ) | ( pg35  &  ng3530  &  (~ ng3522) ) ;
 assign wire30497 = ( ng4975  &  ng4899  &  (~ ng4878) ) ;
 assign wire30498 = ( pg35  &  (~ ng4927)  &  (~ ng4991)  &  (~ ng4864) ) ;
 assign wire30499 = ( (~ ng4966)  &  (~ ng4871)  &  (~ ng4836)  &  (~ ng4983) ) ;
 assign wire30505 = ( pg35  &  ng4975  &  (~ ng4899)  &  (~ ng4991) ) ;
 assign wire30506 = ( (~ ng4864)  &  (~ ng4966)  &  (~ ng4871)  &  (~ ng4836) ) ;
 assign wire30512 = ( pg35  &  (~ ng4975)  &  ng4899  &  (~ ng4991) ) ;
 assign wire30513 = ( (~ ng4864)  &  (~ ng4966)  &  (~ ng4871)  &  (~ ng4836) ) ;
 assign wire30515 = ( ng4975  &  ng4899  &  ng4955 ) | ( ng4975  &  (~ ng4899)  &  ng4933 ) ;
 assign wire30516 = ( ng4888  &  (~ ng4975)  &  (~ ng4899) ) | ( (~ ng4975)  &  ng4899  &  ng4944 ) ;
 assign wire30517 = ( ng4975  &  (~ ng4899)  &  ng4907 ) | ( ng4975  &  ng4899  &  ng4917 ) ;
 assign wire30518 = ( ng4922  &  (~ ng4975)  &  ng4899 ) | ( (~ ng4975)  &  (~ ng4899)  &  ng4912 ) ;
 assign wire30521 = ( pg35  &  (~ ng4864)  &  (~ ng4878) ) ;
 assign wire30523 = ( (~ ng4871)  &  (~ ng4836)  &  (~ ng11173)  &  wire30521 ) ;
 assign wire30527 = ( pg35  &  (~ ng4864)  &  (~ ng4878) ) ;
 assign wire30529 = ( (~ ng4871)  &  (~ ng4836)  &  (~ ng11173)  &  wire30527 ) ;
 assign wire30534 = ( pg35  &  (~ ng4864)  &  (~ ng4878) ) ;
 assign wire30535 = ( (~ ng4966)  &  (~ ng4871)  &  (~ ng4836)  &  ng4983 ) ;
 assign wire30539 = ( pg35  &  (~ ng4864)  &  (~ ng4878) ) ;
 assign wire30547 = ( wire6180 ) | ( wire6181 ) | ( wire6182 ) | ( wire6183 ) ;
 assign wire30550 = ( wire6178 ) | ( wire30547 ) ;
 assign wire30551 = ( wire6173 ) | ( wire6174 ) | ( wire6175 ) | ( wire6179 ) ;
 assign wire30552 = ( ng16696  &  (~ ng16757)  &  wire30523 ) | ( (~ ng16696)  &  ng16757  &  wire30529 ) ;
 assign wire30555 = ( (~ ng2715)  &  (~ ng2803)  &  (~ ng2719) ) ;
 assign wire30557 = ( (~ ng2217) ) | ( (~ ng2185) ) ;
 assign wire30562 = ( pg35  &  (~ ng6181)  &  (~ ng6187) ) ;
 assign wire30564 = ( ng6191  &  pg35 ) ;
 assign wire30566 = ( (~ ng10874)  &  wire30564 ) | ( ng6181  &  ng6187  &  ng10874 ) ;
 assign wire30567 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30568 = ( ng6307  &  pg35 ) ;
 assign wire30570 = ( (~ ng4639)  &  pg35 ) ;
 assign wire30572 = ( pg35  &  ng5037  &  ng17217  &  ng14317 ) ;
 assign wire30573 = ( (~ ng5037)  &  pg35 ) ;
 assign wire30574 = ( wire6160 ) | ( (~ ng17217)  &  wire30573 ) | ( (~ ng14317)  &  wire30573 ) ;
 assign wire30575 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30576 = ( ng6279  &  pg35 ) ;
 assign wire30578 = ( ng93  &  (~ ng4349)  &  (~ ng4358)  &  ng29503 ) ;
 assign wire30581 = ( pg35  &  (~ ng5297)  &  (~ ng23890) ) ;
 assign wire30583 = ( pg35  &  ng5297  &  ng23890 ) ;
 assign wire30585 = ( ng232  &  pg35 ) ;
 assign wire30586 = ( pg14217  &  pg35 ) ;
 assign wire30592 = ( (~ ng1472)  &  ng1467 ) ;
 assign wire30593 = ( ng1472  &  pg35 ) ;
 assign wire30595 = ( (~ pg35)  &  ng1467 ) | ( pg35  &  (~ ng1467)  &  ng1472 ) ;
 assign wire30596 = ( wire30595 ) | ( (~ ng13315)  &  (~ ng10961)  &  wire30592 ) ;
 assign wire30598 = ( pg35  &  (~ ng5990)  &  (~ ng6049)  &  (~ ng6040) ) ;
 assign wire30599 = ( ng4785  &  (~ ng4709)  &  ng11261  &  wire30598 ) ;
 assign wire30601 = ( pg35  &  ng6044  &  ng5990  &  ng6049 ) ;
 assign wire30602 = ( ng4785  &  (~ ng4709)  &  ng11261  &  wire30601 ) ;
 assign wire30604 = ( pg35  &  ng5990  &  (~ ng6049)  &  ng6040 ) ;
 assign wire30605 = ( ng4785  &  (~ ng4709)  &  ng11261  &  wire30604 ) ;
 assign wire30607 = ( pg35  &  (~ ng6044)  &  (~ ng5990)  &  ng6049 ) ;
 assign wire30608 = ( ng4785  &  (~ ng4709)  &  ng11261  &  wire30607 ) ;
 assign wire30609 = ( ng4760  &  pg35 ) ;
 assign wire30611 = ( wire6133 ) | ( ng20875  &  wire30599 ) ;
 assign wire30612 = ( ng20875  &  wire30605 ) | ( pg35  &  ng4760  &  (~ ng20875) ) ;
 assign wire30613 = ( (~ ng23932)  &  wire30602 ) | ( (~ ng23932)  &  wire30608 ) ;
 assign wire30616 = ( (~ ng504)  &  (~ ng518)  &  ng528 ) ;
 assign wire30619 = ( pg35  &  (~ ng2197)  &  ng2227  &  (~ ng112) ) ;
 assign wire30621 = ( pg35  &  ng2197  &  ng112 ) | ( pg35  &  (~ ng2227)  &  ng112 ) ;
 assign wire30622 = ( ng2204  &  pg35 ) ;
 assign wire30628 = ( pg17778  &  ng6741  &  ng6682  &  ng6629 ) ;
 assign wire30629 = ( ng6727  &  pg17764 ) ;
 assign wire30630 = ( ng6741  &  ng6682  &  ng6641 ) ;
 assign wire30631 = ( (~ ng6727)  &  pg17871 ) ;
 assign wire30632 = ( ng6741  &  ng6682  &  ng6617 ) ;
 assign wire30634 = ( pg17688  &  (~ ng6741)  &  (~ ng6682)  &  ng6645 ) ;
 assign wire30635 = ( ng6581  &  pg13099 ) ;
 assign wire30636 = ( (~ ng6741)  &  (~ ng6682)  &  ng6727 ) ;
 assign wire30637 = ( ng6589  &  ng6727 ) ;
 assign wire30638 = ( (~ ng6741)  &  (~ ng6682)  &  ng6723 ) ;
 assign wire30639 = ( ng6727  &  pg14749 ) ;
 assign wire30640 = ( (~ ng6741)  &  ng6682  &  ng6625 ) ;
 assign wire30642 = ( pg14828  &  ng6613  &  (~ ng6741)  &  ng6682 ) ;
 assign wire30643 = ( ng6593  &  pg13099 ) ;
 assign wire30644 = ( (~ ng6741)  &  ng6682  &  (~ ng6727) ) ;
 assign wire30645 = ( ng6597  &  pg17722 ) ;
 assign wire30646 = ( ng6741  &  (~ ng6682)  &  (~ ng6727) ) ;
 assign wire30647 = ( ng6727  &  pg12470 ) ;
 assign wire30648 = ( ng6741  &  (~ ng6682)  &  ng6585 ) ;
 assign wire30649 = ( ng6727  &  pg17871 ) ;
 assign wire30650 = ( ng6741  &  (~ ng6682)  &  ng6609 ) ;
 assign wire30651 = ( (~ ng12471)  &  wire30628 ) | ( wire30629  &  wire30630 ) ;
 assign wire30652 = ( wire30631  &  wire30632 ) | ( (~ ng12471)  &  wire30634 ) ;
 assign wire30653 = ( wire30635  &  wire30636 ) | ( wire30637  &  wire30638 ) ;
 assign wire30654 = ( wire30639  &  wire30640 ) | ( (~ ng12471)  &  wire30642 ) ;
 assign wire30655 = ( wire30643  &  wire30644 ) | ( wire30645  &  wire30646 ) ;
 assign wire30656 = ( wire30647  &  wire30648 ) | ( wire30649  &  wire30650 ) ;
 assign wire30659 = ( wire30656 ) | ( wire30655 ) ;
 assign wire30660 = ( wire30651 ) | ( wire30652 ) | ( wire30653 ) | ( wire30654 ) ;
 assign wire30661 = ( ng6727  &  pg17722 ) ;
 assign wire30662 = ( ng6741  &  ng6682  &  ng6657 ) ;
 assign wire30663 = ( (~ ng6727)  &  pg12470 ) ;
 assign wire30664 = ( ng6741  &  ng6682  &  ng6601 ) ;
 assign wire30665 = ( (~ ng6727)  &  pg14749 ) ;
 assign wire30666 = ( (~ ng6741)  &  (~ ng6682)  &  ng6633 ) ;
 assign wire30668 = ( pg14828  &  ng6621  &  (~ ng6741)  &  (~ ng6682) ) ;
 assign wire30670 = ( pg17688  &  (~ ng6741)  &  ng6653  &  ng6682 ) ;
 assign wire30671 = ( (~ ng6727)  &  ng6605 ) ;
 assign wire30672 = ( (~ ng6741)  &  ng6682  &  ng6723 ) ;
 assign wire30674 = ( pg17778  &  ng6741  &  (~ ng6682)  &  ng6637 ) ;
 assign wire30675 = ( ng6649  &  pg17764 ) ;
 assign wire30676 = ( ng6741  &  (~ ng6682)  &  (~ ng6727) ) ;
 assign wire30677 = ( wire30661  &  wire30662 ) | ( wire30663  &  wire30664 ) ;
 assign wire30678 = ( wire30665  &  wire30666 ) | ( ng12471  &  wire30668 ) ;
 assign wire30679 = ( ng12471  &  wire30670 ) | ( wire30671  &  wire30672 ) ;
 assign wire30680 = ( ng12471  &  wire30674 ) | ( wire30675  &  wire30676 ) ;
 assign wire30683 = ( wire30677 ) | ( wire30678 ) | ( wire30679 ) | ( wire30680 ) ;
 assign wire30685 = ( pg35  &  ng6500  &  ng20751  &  (~ ng11178) ) ;
 assign wire30687 = ( pg35  &  (~ ng6500)  &  ng20751 ) | ( pg35  &  ng20751  &  ng11178 ) ;
 assign wire30688 = ( ng6500  &  pg35 ) ;
 assign wire30692 = ( ng2715  &  (~ ng2724)  &  ng2719 ) ;
 assign wire30694 = ( (~ ng2715)  &  ng2724 ) | ( ng2724  &  (~ ng2719) ) ;
 assign wire30695 = ( (~ pg35)  &  ng2719 ) | ( pg35  &  ng2841  &  wire30692 ) ;
 assign wire30696 = ( pg35  &  ng1644 ) | ( pg35  &  ng2047 ) ;
 assign wire30697 = ( pg35  &  ng2066 ) | ( pg35  &  ng1932 ) ;
 assign wire30698 = ( pg35  &  ng1913 ) | ( pg35  &  ng1664 ) ;
 assign wire30699 = ( pg35  &  ng1779 ) | ( pg35  &  ng1798 ) ;
 assign wire30702 = ( pg35  &  ng2223 ) | ( pg35  &  ng2357 ) ;
 assign wire30703 = ( pg35  &  ng2491 ) | ( pg35  &  ng2625 ) ;
 assign wire30704 = ( pg35  &  ng2472 ) | ( pg35  &  ng2606 ) ;
 assign wire30705 = ( pg35  &  ng2338 ) | ( pg35  &  ng2204 ) ;
 assign wire30708 = ( (~ pg35)  &  ng2898 ) | ( pg35  &  ng2882 ) ;
 assign wire30709 = ( (~ ng2541)  &  pg35 ) ;
 assign wire30710 = ( ng2541  &  pg35 ) ;
 assign wire30712 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30713 = ( ng6653  &  pg35 ) ;
 assign wire30716 = ( pg35  &  ng6741  &  ng6736  &  ng6682 ) ;
 assign wire30717 = ( ng4975  &  ng4899  &  ng11283  &  wire30716 ) ;
 assign wire30719 = ( pg35  &  (~ ng6741)  &  (~ ng6682)  &  (~ ng6732) ) ;
 assign wire30720 = ( ng4975  &  ng4899  &  ng11283  &  wire30719 ) ;
 assign wire30722 = ( pg35  &  (~ ng6741)  &  ng6682  &  ng6732 ) ;
 assign wire30723 = ( ng4975  &  ng4899  &  ng11283  &  wire30722 ) ;
 assign wire30725 = ( pg35  &  ng6741  &  (~ ng6736)  &  (~ ng6682) ) ;
 assign wire30726 = ( ng4975  &  ng4899  &  ng11283  &  wire30725 ) ;
 assign wire30728 = ( ng4894  &  pg35 ) ;
 assign wire30729 = ( wire6064 ) | ( ng20751  &  wire30720 ) ;
 assign wire30730 = ( ng20751  &  wire30723 ) | ( pg35  &  ng4894  &  (~ ng20751) ) ;
 assign wire30731 = ( (~ ng23972)  &  wire30717 ) | ( (~ ng23972)  &  wire30726 ) ;
 assign wire30733 = ( ng2476  &  pg35 ) ;
 assign wire30734 = ( pg35  &  wire7725 ) | ( pg35  &  ng14367  &  wire28488 ) ;
 assign wire30735 = ( ng2453  &  pg35 ) ;
 assign wire30737 = ( wire6057 ) | ( (~ ng27903)  &  wire30734 ) ;
 assign wire30740 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng2724 ) ;
 assign wire30742 = ( (~ ng930)  &  pg35 ) ;
 assign wire30743 = ( pg35  &  pg12919  &  ng930 ) ;
 assign wire30746 = ( pg35  &  (~ ng6682)  &  (~ ng23972) ) ;
 assign wire30748 = ( pg35  &  ng6682  &  ng23972 ) ;
 assign wire30750 = ( (~ ng4899)  &  pg35 ) ;
 assign wire30752 = ( ng4899  &  pg35 ) ;
 assign wire30754 = ( wire6042 ) | ( (~ ng16187)  &  ng28349  &  wire30750 ) ;
 assign wire30759 = ( pg35  &  (~ pg9048)  &  ng604 ) | ( pg35  &  ng604  &  ng559 ) ;
 assign wire30760 = ( (~ ng604)  &  pg35 ) ;
 assign wire30763 = ( pg35  &  ng1811  &  (~ ng14640) ) ;
 assign wire30765 = ( pg35  &  (~ ng1811)  &  ng14640 ) ;
 assign wire30768 = ( ng22369  &  wire30765 ) | ( pg35  &  ng1825  &  (~ ng22369) ) ;
 assign wire30769 = ( ng4392  &  pg35 ) ;
 assign wire30770 = ( (~ ng4392)  &  (~ ng4417) ) ;
 assign wire30776 = ( (~ ng504)  &  ng499 ) ;
 assign wire30782 = ( (~ ng718)  &  (~ ng655)  &  (~ ng650)  &  ng699 ) ;
 assign wire30783 = ( (~ ng661)  &  (~ ng728)  &  ng681  &  (~ ng645) ) ;
 assign wire30788 = ( (~ ng718)  &  (~ ng655)  &  (~ ng650)  &  ng699 ) ;
 assign wire30789 = ( ng661  &  ng728  &  ng681  &  (~ ng645) ) ;
 assign wire30794 = ( ng718  &  ng655  &  (~ ng650)  &  ng699 ) ;
 assign wire30795 = ( (~ ng661)  &  (~ ng728)  &  ng681  &  (~ ng645) ) ;
 assign wire30800 = ( ng718  &  ng655  &  (~ ng650)  &  ng699 ) ;
 assign wire30801 = ( ng661  &  ng728  &  ng681  &  (~ ng645) ) ;
 assign wire30802 = ( wire30782  &  wire30783 ) | ( wire30788  &  wire30789 ) ;
 assign wire30803 = ( wire30794  &  wire30795 ) | ( wire30800  &  wire30801 ) ;
 assign wire30805 = ( pg35  &  (~ ng714)  &  ng676  &  ng20375 ) ;
 assign wire30807 = ( pg35  &  ng714  &  (~ ng676) ) | ( pg35  &  ng714  &  (~ ng20375) ) ;
 assign wire30809 = ( ng79  &  pg35 ) ;
 assign wire30810 = ( ng728  &  pg35 ) ;
 assign wire30811 = ( ng661  &  pg35 ) ;
 assign wire30817 = ( pg17711  &  ng5703  &  ng5644  &  ng5591 ) ;
 assign wire30819 = ( pg17580  &  (~ ng5703)  &  (~ ng5644)  &  ng5607 ) ;
 assign wire30821 = ( pg14694  &  (~ ng5703)  &  ng5575  &  ng5644 ) ;
 assign wire30823 = ( ng5703  &  (~ ng5644)  &  ng5547 ) ;
 assign wire30824 = ( (~ ng5689)  &  pg17604 ) ;
 assign wire30825 = ( ng5703  &  (~ ng5644)  &  ng5559 ) ;
 assign wire30826 = ( ng5689  &  pg17813 ) ;
 assign wire30827 = ( ng5703  &  ng5571  &  (~ ng5644) ) ;
 assign wire30828 = ( ng5685  &  ng5689 ) ;
 assign wire30829 = ( (~ ng5703)  &  ng5551  &  (~ ng5644) ) ;
 assign wire30830 = ( ng5689  &  pg13049 ) ;
 assign wire30831 = ( (~ ng5703)  &  ng5543  &  (~ ng5644) ) ;
 assign wire30832 = ( ng5689  &  pg14635 ) ;
 assign wire30833 = ( (~ ng5703)  &  ng5644  &  ng5587 ) ;
 assign wire30834 = ( (~ ng5689)  &  pg13049 ) ;
 assign wire30835 = ( (~ ng5703)  &  ng5555  &  ng5644 ) ;
 assign wire30836 = ( ng5689  &  pg17678 ) ;
 assign wire30837 = ( ng5703  &  ng5603  &  ng5644 ) ;
 assign wire30838 = ( (~ ng5689)  &  pg17813 ) ;
 assign wire30839 = ( ng5703  &  ng5579  &  ng5644 ) ;
 assign wire30840 = ( pg12300  &  ng5689  &  wire30817 ) | ( (~ pg12300)  &  (~ ng5689)  &  wire30817 ) | ( pg12300  &  ng5689  &  wire30819 ) | ( (~ pg12300)  &  (~ ng5689)  &  wire30819 ) ;
 assign wire30841 = ( pg12300  &  ng5689  &  wire30821 ) | ( (~ pg12300)  &  (~ ng5689)  &  wire30821 ) | ( pg12300  &  ng5689  &  wire30823 ) ;
 assign wire30842 = ( wire30824  &  wire30825 ) | ( wire30826  &  wire30827 ) ;
 assign wire30843 = ( wire30828  &  wire30829 ) | ( wire30830  &  wire30831 ) ;
 assign wire30844 = ( wire30832  &  wire30833 ) | ( wire30834  &  wire30835 ) ;
 assign wire30845 = ( wire30836  &  wire30837 ) | ( wire30838  &  wire30839 ) ;
 assign wire30848 = ( wire30845 ) | ( wire30844 ) ;
 assign wire30849 = ( wire30840 ) | ( wire30841 ) | ( wire30842 ) | ( wire30843 ) ;
 assign wire30851 = ( pg17711  &  ng5599  &  ng5703  &  (~ ng5644) ) ;
 assign wire30853 = ( pg17580  &  (~ ng5703)  &  ng5644  &  ng5615 ) ;
 assign wire30855 = ( pg14694  &  ng5583  &  (~ ng5703)  &  (~ ng5644) ) ;
 assign wire30856 = ( (~ ng5689)  &  pg17678 ) ;
 assign wire30857 = ( ng5703  &  (~ ng5644)  &  ng5611 ) ;
 assign wire30858 = ( (~ ng5689)  &  pg14635 ) ;
 assign wire30859 = ( (~ ng5703)  &  (~ ng5644)  &  ng5595 ) ;
 assign wire30860 = ( ng5685  &  (~ ng5689) ) ;
 assign wire30861 = ( (~ ng5703)  &  ng5567  &  ng5644 ) ;
 assign wire30862 = ( ng5689  &  pg17604 ) ;
 assign wire30863 = ( ng5703  &  ng5619  &  ng5644 ) ;
 assign wire30864 = ( (~ ng5689)  &  pg12300 ) ;
 assign wire30865 = ( ng5703  &  ng5563  &  ng5644 ) ;
 assign wire30866 = ( (~ pg12300)  &  ng5689  &  wire30851 ) | ( pg12300  &  (~ ng5689)  &  wire30851 ) | ( (~ pg12300)  &  ng5689  &  wire30853 ) | ( pg12300  &  (~ ng5689)  &  wire30853 ) ;
 assign wire30867 = ( ng12301  &  wire30855 ) | ( wire30856  &  wire30857 ) ;
 assign wire30868 = ( wire30858  &  wire30859 ) | ( wire30860  &  wire30861 ) ;
 assign wire30869 = ( wire30862  &  wire30863 ) | ( wire30864  &  wire30865 ) ;
 assign wire30872 = ( wire30866 ) | ( wire30867 ) | ( wire30868 ) | ( wire30869 ) ;
 assign wire30874 = ( pg35  &  (~ ng5462)  &  ng20739 ) | ( pg35  &  ng20739  &  ng11123 ) ;
 assign wire30876 = ( pg35  &  ng5462  &  ng20739  &  (~ ng11123) ) ;
 assign wire30877 = ( ng5462  &  pg35 ) ;
 assign wire30880 = ( pg35  &  (~ ng5062) ) | ( pg35  &  (~ ng5046) ) | ( pg35  &  (~ wire29546) ) ;
 assign wire30881 = ( ng1592  &  pg35 ) ;
 assign wire30888 = ( ng2153  &  pg35 ) ;
 assign wire30893 = ( pg35  &  (~ ng1854)  &  (~ ng1848) ) ;
 assign wire30895 = ( pg35  &  ng1854  &  ng1848 ) ;
 assign wire30898 = ( (~ ng25300)  &  wire30895 ) | ( pg35  &  ng1858  &  ng25300 ) ;
 assign wire30899 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire30900 = ( ng6581  &  pg35 ) ;
 assign wire30901 = ( wire5955 ) | ( ng7142  &  ng12716  &  wire30899 ) ;
 assign wire30902 = ( (~ ng1906)  &  pg35 ) ;
 assign wire30906 = ( pg35  &  ng1902  &  ng25429 ) | ( pg35  &  ng1862  &  (~ ng25429) ) ;
 assign wire30908 = ( pg35  &  (~ ng2116)  &  (~ ng2122) ) ;
 assign wire30910 = ( ng2126  &  pg35 ) ;
 assign wire30912 = ( ng25389  &  wire30910 ) | ( ng2116  &  ng2122  &  (~ ng25389) ) ;
 assign wire30914 = ( pg35  &  (~ pg9048)  &  ng582 ) | ( pg35  &  ng582  &  ng559 ) ;
 assign wire30915 = ( (~ ng582)  &  pg35 ) ;
 assign wire30918 = ( pg35  &  (~ ng3841)  &  (~ ng3835) ) ;
 assign wire30920 = ( pg35  &  ng3841  &  ng3835 ) ;
 assign wire30923 = ( ng12735  &  wire30920 ) | ( pg35  &  ng3845  &  (~ ng12735) ) ;
 assign wire30926 = ( pg35  &  ng2016  &  (~ ng2060)  &  (~ ng2028) ) ;
 assign wire30929 = ( pg35  &  (~ ng2051)  &  ng2020  &  ng2028 ) ;
 assign wire30931 = ( pg35  &  ng2004  &  ng2051  &  (~ ng2028) ) ;
 assign wire30932 = ( ng2012  &  (~ ng2051)  &  ng2060 ) ;
 assign wire30933 = ( ng2079  &  pg35 ) ;
 assign wire30934 = ( ng2024  &  pg35 ) ;
 assign wire30938 = ( ng2008  &  (~ ng25389) ) | ( (~ ng25470)  &  wire30934 ) ;
 assign wire30939 = ( wire5925 ) | ( wire5926 ) | ( wire5927 ) | ( wire5931 ) ;
 assign wire30945 = ( (~ ng5343)  &  pg17577 ) ;
 assign wire30946 = ( (~ ng5297)  &  ng5357  &  ng5212 ) ;
 assign wire30948 = ( pg17519  &  (~ ng5297)  &  (~ ng5357)  &  ng5260 ) ;
 assign wire30949 = ( ng5343  &  ng5204 ) ;
 assign wire30950 = ( (~ ng5297)  &  (~ ng5357)  &  ng5339 ) ;
 assign wire30951 = ( ng5343  &  pg13039 ) ;
 assign wire30952 = ( (~ ng5297)  &  (~ ng5357)  &  ng5196 ) ;
 assign wire30954 = ( pg14662  &  ng5297  &  (~ ng5357)  &  ng5228 ) ;
 assign wire30956 = ( pg17674  &  ng5244  &  ng5297  &  ng5357 ) ;
 assign wire30957 = ( (~ ng5343)  &  pg13039 ) ;
 assign wire30958 = ( ng5297  &  (~ ng5357)  &  ng5208 ) ;
 assign wire30959 = ( ng5240  &  pg14597 ) ;
 assign wire30960 = ( ng5297  &  (~ ng5357)  &  ng5343 ) ;
 assign wire30961 = ( ng5343  &  pg17787 ) ;
 assign wire30962 = ( (~ ng5297)  &  ng5357  &  ng5224 ) ;
 assign wire30963 = ( ng5200  &  pg12238 ) ;
 assign wire30964 = ( (~ ng5297)  &  ng5357  &  ng5343 ) ;
 assign wire30965 = ( (~ ng5343)  &  pg17787 ) ;
 assign wire30966 = ( ng5297  &  ng5357  &  ng5232 ) ;
 assign wire30967 = ( ng5256  &  pg17639 ) ;
 assign wire30968 = ( ng5297  &  ng5357  &  ng5343 ) ;
 assign wire30969 = ( wire30945  &  wire30946 ) | ( (~ ng12239)  &  wire30948 ) ;
 assign wire30970 = ( wire30949  &  wire30950 ) | ( wire30951  &  wire30952 ) ;
 assign wire30971 = ( pg12238  &  ng5343  &  wire30954 ) | ( (~ pg12238)  &  (~ ng5343)  &  wire30954 ) | ( pg12238  &  ng5343  &  wire30956 ) | ( (~ pg12238)  &  (~ ng5343)  &  wire30956 ) ;
 assign wire30972 = ( wire30957  &  wire30958 ) | ( wire30959  &  wire30960 ) ;
 assign wire30973 = ( wire30961  &  wire30962 ) | ( wire30963  &  wire30964 ) ;
 assign wire30974 = ( wire30965  &  wire30966 ) | ( wire30967  &  wire30968 ) ;
 assign wire30977 = ( wire30974 ) | ( wire30973 ) ;
 assign wire30978 = ( wire30969 ) | ( wire30970 ) | ( wire30971 ) | ( wire30972 ) ;
 assign wire30980 = ( pg14662  &  (~ ng5297)  &  (~ ng5357)  &  ng5236 ) ;
 assign wire30981 = ( ng5248  &  pg14597 ) ;
 assign wire30982 = ( (~ ng5297)  &  (~ ng5357)  &  (~ ng5343) ) ;
 assign wire30984 = ( pg17519  &  ng5297  &  (~ ng5357)  &  ng5268 ) ;
 assign wire30986 = ( pg17674  &  (~ ng5297)  &  ng5357  &  ng5252 ) ;
 assign wire30987 = ( ng5339  &  (~ ng5343) ) ;
 assign wire30988 = ( ng5297  &  (~ ng5357)  &  ng5220 ) ;
 assign wire30989 = ( (~ ng5343)  &  pg17639 ) ;
 assign wire30990 = ( (~ ng5297)  &  ng5357  &  ng5264 ) ;
 assign wire30991 = ( ng5343  &  pg17577 ) ;
 assign wire30992 = ( ng5297  &  ng5357  &  ng5272 ) ;
 assign wire30993 = ( ng5216  &  pg12238 ) ;
 assign wire30994 = ( ng5297  &  ng5357  &  (~ ng5343) ) ;
 assign wire30995 = ( ng12239  &  wire30980 ) | ( wire30981  &  wire30982 ) ;
 assign wire30996 = ( (~ pg12238)  &  ng5343  &  wire30984 ) | ( pg12238  &  (~ ng5343)  &  wire30984 ) | ( (~ pg12238)  &  ng5343  &  wire30986 ) | ( pg12238  &  (~ ng5343)  &  wire30986 ) ;
 assign wire30997 = ( wire30987  &  wire30988 ) | ( wire30989  &  wire30990 ) ;
 assign wire30998 = ( wire30991  &  wire30992 ) | ( wire30993  &  wire30994 ) ;
 assign wire31001 = ( wire30995 ) | ( wire30996 ) | ( wire30997 ) | ( wire30998 ) ;
 assign wire31002 = ( pg35  &  wire7624 ) | ( pg35  &  wire7625 ) | ( pg35  &  wire28651 ) ;
 assign wire31003 = ( ng128  &  pg35 ) ;
 assign wire31005 = ( ng2715  &  (~ ng2819)  &  ng2719 ) ;
 assign wire31007 = ( pg35  &  wire5887 ) | ( pg35  &  ng14367  &  wire31005 ) ;
 assign wire31008 = ( ng2610  &  pg35 ) ;
 assign wire31010 = ( wire5884 ) | ( (~ ng27933)  &  wire31007 ) ;
 assign wire31015 = ( pg35  &  (~ ng3139)  &  (~ ng3133) ) ;
 assign wire31017 = ( pg35  &  ng3139  &  ng3133 ) ;
 assign wire31020 = ( ng12641  &  wire31017 ) | ( pg35  &  ng3143  &  (~ ng12641) ) ;
 assign wire31022 = ( pg35  &  wire7030 ) | ( pg35  &  ng14367  &  wire29111 ) ;
 assign wire31023 = ( ng2342  &  pg35 ) ;
 assign wire31025 = ( wire5869 ) | ( (~ ng27854)  &  wire31022 ) ;
 assign wire31026 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31027 = ( ng3574  &  pg35 ) ;
 assign wire31030 = ( pg35  &  (~ ng2342)  &  (~ ng2351) ) ;
 assign wire31031 = ( pg35  &  wire7030 ) | ( pg35  &  ng14367  &  wire29111 ) ;
 assign wire31033 = ( ng2319  &  pg35 ) ;
 assign wire31034 = ( (~ pg35)  &  ng2327 ) | ( pg35  &  ng2319  &  (~ ng2351) ) ;
 assign wire31036 = ( wire5859 ) | ( (~ ng27854)  &  wire31031 ) ;
 assign wire31040 = ( (~ pg35)  &  ng5802 ) | ( pg35  &  pg9617  &  (~ pg9680)  &  (~ ng5802) ) ;
 assign wire31041 = ( ng1041  &  pg35 ) ;
 assign wire31043 = ( wire5847 ) | ( ng13211  &  wire31041 ) | ( wire5848  &  wire31041 ) ;
 assign wire31045 = ( (~ pg35) ) | ( ng4462 ) | ( ng4473  &  ng4467 ) ;
 assign wire31050 = ( pg35  &  ng2599  &  ng112 ) | ( pg35  &  ng112  &  (~ ng2629) ) ;
 assign wire31052 = ( pg35  &  (~ ng2599)  &  (~ ng112)  &  ng2629 ) ;
 assign wire31053 = ( ng2606  &  pg35 ) ;
 assign wire31056 = ( ng262  &  pg35 ) ;
 assign wire31057 = ( pg14096  &  pg35 ) ;
 assign wire31060 = ( pg35  &  (~ ng5808)  &  ng5813 ) ;
 assign wire31061 = ( (~ ng5813)  &  ng5808 ) ;
 assign wire31063 = ( (~ ng23666)  &  wire31061 ) | ( pg35  &  ng5817  &  ng23666 ) ;
 assign wire31064 = ( ng4950  &  pg35 ) ;
 assign wire31065 = ( wire1421  &  wire31064 ) | ( ng4818  &  wire31064 ) | ( (~ ng24374)  &  wire31064 ) ;
 assign wire31067 = ( pg35  &  ng71  &  ng24374  &  (~ wire28575) ) ;
 assign wire31069 = ( ng29722  &  wire31067 ) | ( pg35  &  ng4944  &  (~ ng29722) ) ;
 assign wire31070 = ( ng3827  &  pg35 ) ;
 assign wire31073 = ( pg35  &  (~ ng5297)  &  (~ ng5357)  &  (~ ng5348) ) ;
 assign wire31074 = ( ng4785  &  ng4709  &  ng11261  &  wire31073 ) ;
 assign wire31076 = ( pg35  &  ng5297  &  (~ ng5357)  &  ng5348 ) ;
 assign wire31077 = ( ng4785  &  ng4709  &  ng11261  &  wire31076 ) ;
 assign wire31079 = ( pg35  &  (~ ng5297)  &  ng5357  &  (~ ng5352) ) ;
 assign wire31080 = ( ng4785  &  ng4709  &  ng11261  &  wire31079 ) ;
 assign wire31082 = ( pg35  &  ng5297  &  ng5357  &  ng5352 ) ;
 assign wire31083 = ( ng4785  &  ng4709  &  ng11261  &  wire31082 ) ;
 assign wire31084 = ( ng4704  &  pg35 ) ;
 assign wire31086 = ( wire5819 ) | ( ng20682  &  wire31074 ) ;
 assign wire31087 = ( ng20682  &  wire31077 ) | ( pg35  &  ng4704  &  (~ ng20682) ) ;
 assign wire31088 = ( (~ ng23890)  &  wire31080 ) | ( (~ ng23890)  &  wire31083 ) ;
 assign wire31090 = ( ng336  &  pg35 ) ;
 assign wire31091 = ( ng305  &  pg35 ) ;
 assign wire31093 = ( (~ ng2227)  &  pg35 ) ;
 assign wire31095 = ( ng26703  &  (~ ng28768)  &  wire31093 ) | ( ng17321  &  (~ ng28768)  &  wire31093 ) ;
 assign wire31098 = ( pg35  &  (~ ng3470)  &  (~ ng3476) ) ;
 assign wire31100 = ( ng3480  &  pg35 ) ;
 assign wire31102 = ( ng23112  &  wire31100 ) | ( ng3470  &  ng3476  &  (~ ng23112) ) ;
 assign wire31105 = ( pg35  &  (~ ng4674)  &  (~ ng4681)  &  (~ ng4646) ) ;
 assign wire31107 = ( (~ ng5357)  &  pg35 ) ;
 assign wire31109 = ( ng5357  &  pg35 ) ;
 assign wire31111 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31112 = ( ng3937  &  pg35 ) ;
 assign wire31114 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31115 = ( ng5949  &  pg35 ) ;
 assign wire31120 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31121 = ( ng6247  &  pg35 ) ;
 assign wire31122 = ( wire5788 ) | ( ng12581  &  ng12667  &  wire31120 ) ;
 assign wire31123 = ( pg35  &  pg12923  &  ng1259 ) ;
 assign wire31124 = ( pg35  &  ng1256  &  ng1252  &  ng19140 ) ;
 assign wire31126 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31127 = ( ng6589  &  pg35 ) ;
 assign wire31131 = ( pg35  &  ng1936  &  (~ ng1906)  &  (~ ng112) ) ;
 assign wire31133 = ( pg35  &  (~ ng1936)  &  ng112 ) | ( pg35  &  ng1906  &  ng112 ) ;
 assign wire31134 = ( ng1913  &  pg35 ) ;
 assign wire31140 = ( ng446  &  pg35 ) ;
 assign wire31141 = ( ng182  &  pg35 ) ;
 assign wire31143 = ( ng1592 ) | ( (~ ng1636) ) ;
 assign wire31144 = ( (~ ng1668)  &  pg35 ) ;
 assign wire31146 = ( (~ ng28739)  &  ng26673  &  wire31144 ) | ( (~ ng28739)  &  ng17292  &  wire31144 ) ;
 assign wire31148 = ( pg35  &  ng2495  &  ng2509 ) | ( pg35  &  ng2509  &  ng2421 ) ;
 assign wire31149 = ( ng26770  &  wire31148 ) | ( ng17424  &  wire31148 ) ;
 assign wire31150 = ( pg35  &  (~ ng2509) ) | ( pg35  &  (~ ng2495)  &  (~ ng2421) ) ;
 assign wire31151 = ( ng26770  &  wire31150 ) | ( ng17424  &  wire31150 ) ;
 assign wire31152 = ( ng2509  &  pg35 ) ;
 assign wire31153 = ( wire5759 ) | ( (~ ng26770)  &  (~ ng17424)  &  wire31152 ) ;
 assign wire31155 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31156 = ( ng3921  &  pg35 ) ;
 assign wire31158 = ( pg35  &  ng11915  &  ng17317 ) | ( pg35  &  ng11915  &  ng26694 ) ;
 assign wire31159 = ( ng1756  &  pg35 ) ;
 assign wire31161 = ( ng872  &  pg35 ) ;
 assign wire31162 = ( ng446  &  pg35 ) ;
 assign wire31165 = ( pg35  &  (~ ng4349)  &  (~ ng12925) ) ;
 assign wire31167 = ( pg35  &  ng4349  &  ng12925 ) ;
 assign wire31170 = ( pg35  &  ng6159  &  (~ ng6154) ) ;
 assign wire31171 = ( ng6154  &  (~ ng6159) ) ;
 assign wire31173 = ( (~ ng23699)  &  wire31171 ) | ( pg35  &  ng6163  &  ng23699 ) ;
 assign wire31174 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31175 = ( ng5248  &  pg35 ) ;
 assign wire31177 = ( (~ ng4392)  &  pg35 ) ;
 assign wire31178 = ( wire5727 ) | ( wire29520  &  wire29521  &  wire31177 ) ;
 assign wire31182 = ( (~ pg11447)  &  (~ pg8789) ) ;
 assign wire31183 = ( pg35  &  (~ pg8783)  &  (~ ng4180) ) ;
 assign wire31184 = ( (~ pg8784)  &  (~ pg8785)  &  (~ pg8787)  &  (~ pg8788) ) ;
 assign wire31189 = ( (~ pg35)  &  ng2946 ) | ( pg35  &  (~ pg8786)  &  ng4180 ) | ( pg35  &  pg8786  &  (~ ng4180) ) ;
 assign wire31190 = ( (~ ng2116)  &  pg35 ) ;
 assign wire31191 = ( ng2116  &  pg35 ) ;
 assign wire31194 = ( pg35  &  (~ ng2485)  &  (~ ng2476) ) | ( pg35  &  (~ ng2485)  &  ng2453 ) ;
 assign wire31195 = ( ng2453  &  pg35 ) ;
 assign wire31196 = ( pg35  &  wire7725 ) | ( pg35  &  ng14367  &  wire28488 ) ;
 assign wire31198 = ( wire5713 ) | ( (~ ng27903)  &  wire31196 ) ;
 assign wire31201 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31202 = ( ng3606  &  pg35 ) ;
 assign wire31204 = ( (~ ng843)  &  ng837 ) ;
 assign wire31205 = ( ng843  &  ng837 ) ;
 assign wire31206 = ( wire5702 ) | ( ng847  &  (~ ng8806)  &  wire31204 ) ;
 assign wire31210 = ( pg35  &  (~ ng1036)  &  (~ ng15737) ) ;
 assign wire31211 = ( ng1036  &  pg35 ) ;
 assign wire31213 = ( ng4104  &  pg35 ) ;
 assign wire31214 = ( (~ ng4104)  &  pg35 ) ;
 assign wire31215 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng4108 ) ;
 assign wire31217 = ( ng1706  &  pg35 ) ;
 assign wire31220 = ( pg35  &  (~ ng5523)  &  ng5511  &  ng5517 ) ;
 assign wire31226 = ( pg35  &  (~ ng1306) ) | ( pg35  &  (~ ng962) ) ;
 assign wire31229 = ( pg35  &  ng17405  &  ng11939 ) | ( pg35  &  ng26737  &  ng11939 ) ;
 assign wire31230 = ( ng2315  &  pg35 ) ;
 assign wire31232 = ( ng2619 ) | ( (~ ng2610) ) ;
 assign wire31233 = ( ng2555  &  pg35 ) ;
 assign wire31237 = ( pg35  &  ng2595  &  ng25498 ) | ( pg35  &  (~ ng2599)  &  (~ ng25498) ) ;
 assign wire31240 = ( (~ ng2652)  &  ng2638 ) | ( ng2610  &  (~ ng2587)  &  ng2638 ) ;
 assign wire31241 = ( ng2652  &  pg35 ) ;
 assign wire31242 = ( (~ pg35)  &  ng2638 ) | ( pg35  &  (~ ng2638)  &  ng22498  &  ng14752 ) ;
 assign wire31244 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31245 = ( ng6235  &  pg35 ) ;
 assign wire31246 = ( wire5661 ) | ( ng10341  &  ng12667  &  wire31244 ) ;
 assign wire31250 = ( ng1840  &  pg35 ) ;
 assign wire31254 = ( pg35  &  ng822  &  ng723  &  (~ ng847) ) ;
 assign wire31255 = ( ng703  &  pg35 ) ;
 assign wire31256 = ( ng703  &  (~ ng837) ) ;
 assign wire31259 = ( wire5649 ) | ( (~ ng14279)  &  wire31255 ) | ( ng14279  &  wire31256 ) ;
 assign wire31268 = ( pg35  &  (~ ng2841)  &  (~ ng4098) ) | ( pg35  &  (~ ng2841)  &  (~ ng4076) ) ;
 assign wire31271 = ( wire5641 ) | ( wire5642 ) | ( wire31268 ) ;
 assign wire31275 = ( ng1862  &  pg35 ) ;
 assign wire31281 = ( ng1945  &  (~ ng1959) ) | ( ng1945  &  ng1917  &  (~ ng1894) ) ;
 assign wire31282 = ( ng1959  &  pg35 ) ;
 assign wire31283 = ( (~ pg35)  &  ng1945 ) | ( pg35  &  (~ ng1945)  &  ng22417  &  ng14678 ) ;
 assign wire31287 = ( pg35  &  ng2375  &  ng2361 ) | ( pg35  &  ng2375  &  ng2287 ) ;
 assign wire31288 = ( ng17405  &  wire31287 ) | ( ng26737  &  wire31287 ) ;
 assign wire31289 = ( pg35  &  (~ ng2375) ) | ( pg35  &  (~ ng2361)  &  (~ ng2287) ) ;
 assign wire31290 = ( ng17405  &  wire31289 ) | ( ng26737  &  wire31289 ) ;
 assign wire31291 = ( ng2375  &  pg35 ) ;
 assign wire31292 = ( wire5623 ) | ( (~ ng17405)  &  (~ ng26737)  &  wire31291 ) ;
 assign wire31295 = ( pg35  &  (~ ng4991)  &  ng4983  &  ng10862 ) ;
 assign wire31297 = ( pg35  &  ng4991  &  (~ ng4983) ) | ( pg35  &  ng4991  &  (~ ng10862) ) ;
 assign wire31298 = ( wire5619 ) | ( ng28349  &  ng13486  &  wire31295 ) ;
 assign wire31301 = ( pg35  &  (~ ng2715)  &  (~ ng2771) ) ;
 assign wire31304 = ( pg35  &  ng2715  &  (~ ng2775) ) ;
 assign wire31308 = ( pg35  &  (~ ng2715)  &  ng1677 ) ;
 assign wire31311 = ( pg35  &  ng2715  &  ng1811 ) ;
 assign wire31313 = ( ng2719  &  pg35 ) ;
 assign wire31316 = ( pg35  &  ng2719  &  (~ ng23618) ) ;
 assign wire31317 = ( ng21277  &  (~ ng23532)  &  wire31301 ) | ( ng21277  &  (~ ng23532)  &  wire31304 ) ;
 assign wire31318 = ( (~ ng21277)  &  (~ ng23618)  &  wire31308 ) | ( (~ ng21277)  &  (~ ng23618)  &  wire31311 ) ;
 assign wire31319 = ( (~ ng21277)  &  wire31316 ) | ( ng21277  &  (~ ng23532)  &  wire31313 ) ;
 assign wire31322 = ( pg35  &  (~ pg11678)  &  (~ ng739) ) | ( pg35  &  (~ ng739)  &  ng736 ) ;
 assign wire31324 = ( pg35  &  (~ pg11678)  &  ng739 ) | ( pg35  &  ng739  &  ng736 ) ;
 assign wire31326 = ( (~ ng5084)  &  pg35 ) ;
 assign wire31327 = ( ng5069  &  (~ ng5080) ) | ( (~ ng5077)  &  (~ ng5080) ) ;
 assign wire31328 = ( (~ pg35)  &  ng5080 ) | ( ng5084  &  ng5080 ) ;
 assign wire31332 = ( ng4785  &  pg35 ) ;
 assign wire31333 = ( wire5595 ) | ( ng28336  &  ng13464  &  wire31332 ) ;
 assign wire31334 = ( (~ ng1902)  &  pg35 ) ;
 assign wire31337 = ( (~ pg35)  &  ng2779 ) | ( pg35  &  ng2791  &  (~ ng12377) ) ;
 assign wire31338 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31339 = ( ng6609  &  pg35 ) ;
 assign wire31342 = ( pg35  &  (~ ng2093)  &  ng2089 ) ;
 assign wire31344 = ( ng2098  &  pg35 ) ;
 assign wire31346 = ( ng25492  &  wire31344 ) | ( ng2093  &  (~ ng2089)  &  (~ ng25492) ) ;
 assign wire31347 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31348 = ( ng3546  &  pg35 ) ;
 assign wire31351 = ( pg35  &  ng2185  &  (~ ng2217) ) | ( pg35  &  (~ ng2217)  &  (~ ng2208) ) ;
 assign wire31353 = ( pg35  &  wire6172 ) | ( pg35  &  ng14367  &  wire30555 ) ;
 assign wire31354 = ( ng2185  &  pg35 ) ;
 assign wire31356 = ( wire5576 ) | ( (~ ng27796)  &  wire31353 ) ;
 assign wire31357 = ( ng29503  &  wire7725 ) | ( ng29503  &  ng14367  &  wire28488 ) ;
 assign wire31359 = ( pg35  &  (~ ng2485)  &  ng110 ) | ( pg35  &  ng110  &  ng2476 ) ;
 assign wire31361 = ( pg35  &  ng2485  &  (~ ng110)  &  (~ ng2476) ) ;
 assign wire31362 = ( ng2491  &  pg35 ) ;
 assign wire31363 = ( wire5573 ) | ( ng26218  &  wire31357  &  wire31359 ) ;
 assign wire31364 = ( (~ ng26218)  &  wire31362 ) | ( (~ wire31357)  &  wire31362 ) | ( ng26218  &  wire31357  &  wire31361 ) ;
 assign wire31366 = ( pg35  &  ng1322  &  (~ ng1351) ) | ( pg35  &  (~ ng1351)  &  ng1333 ) ;
 assign wire31367 = ( ng1345  &  ng1367  &  ng1379  &  wire31366 ) ;
 assign wire31368 = ( (~ ng1389)  &  pg35 ) ;
 assign wire31369 = ( ng1361  &  ng1351  &  ng1373 ) ;
 assign wire31372 = ( pg35  &  ng1322  &  ng1339 ) | ( pg35  &  (~ ng1322)  &  ng1333  &  (~ ng1339) ) ;
 assign wire31373 = ( ng1312  &  pg35 ) ;
 assign wire31374 = ( ng13242  &  wire31373 ) | ( (~ ng13242)  &  wire31368  &  wire31369 ) ;
 assign wire31377 = ( ng1124  &  (~ ng1129) ) ;
 assign wire31378 = ( ng1129  &  pg35 ) ;
 assign wire31379 = ( (~ pg35)  &  ng1124 ) | ( pg35  &  ng1129  &  (~ ng1124) ) ;
 assign wire31380 = ( wire31379 ) | ( (~ ng13307)  &  (~ ng10929)  &  wire31377 ) ;
 assign wire31385 = ( pg35  &  ng1624  &  (~ ng1657) ) | ( pg35  &  (~ ng1657)  &  (~ ng1648) ) ;
 assign wire31387 = ( pg35  &  wire7041 ) | ( pg35  &  ng14367  &  wire29097 ) ;
 assign wire31388 = ( ng1624  &  pg35 ) ;
 assign wire31390 = ( wire5557 ) | ( (~ ng27738)  &  wire31387 ) ;
 assign wire31391 = ( (~ ng1848)  &  pg35 ) ;
 assign wire31392 = ( ng1848  &  pg35 ) ;
 assign wire31395 = ( pg35  &  (~ ng4859)  &  (~ ng13346) ) ;
 assign wire31397 = ( pg35  &  ng4859  &  ng13346 ) ;
 assign wire31398 = ( wire5551 ) | ( ng31009  &  (~ ng10862)  &  wire31395 ) ;
 assign wire31399 = ( ng956  &  pg35 ) ;
 assign wire31400 = ( (~ ng956)  &  ng1141 ) ;
 assign wire31402 = ( (~ pg35)  &  ng1141 ) | ( pg35  &  (~ ng1141)  &  ng956 ) ;
 assign wire31403 = ( wire31402 ) | ( ng10929  &  wire31399 ) | ( ng10909  &  wire31399 ) ;
 assign wire31404 = ( (~ ng2495)  &  pg35 ) ;
 assign wire31406 = ( ng26770  &  (~ ng28846)  &  wire31404 ) | ( ng17424  &  (~ ng28846)  &  wire31404 ) ;
 assign wire31414 = ( pg35  &  ng9694  &  ng26725 ) | ( pg35  &  ng9694  &  ng17401 ) ;
 assign wire31415 = ( ng1874  &  pg35 ) ;
 assign wire31424 = ( ng2351 ) | ( (~ ng2342) ) ;
 assign wire31425 = ( ng2287  &  pg35 ) ;
 assign wire31429 = ( pg35  &  ng2327  &  ng25435 ) | ( pg35  &  (~ ng2331)  &  (~ ng25435) ) ;
 assign wire31431 = ( pg35  &  (~ ng723)  &  (~ ng14279) ) ;
 assign wire31433 = ( pg35  &  ng723  &  (~ ng14279) ) ;
 assign wire31434 = ( (~ pg35)  &  ng827 ) | ( ng827  &  (~ ng20905)  &  wire31431 ) ;
 assign wire31435 = ( (~ ng4349)  &  ng4358  &  (~ ng24380)  &  wire29233 ) ;
 assign wire31437 = ( (~ ng3703)  &  pg35 ) ;
 assign wire31439 = ( ng3703  &  pg35 ) ;
 assign wire31445 = ( (~ pg72)  &  pg35  &  ng4581 ) | ( pg35  &  ng4575  &  ng4581 ) ;
 assign wire31446 = ( (~ pg35)  &  ng4546 ) | ( ng4546  &  (~ ng4581) ) | ( pg73  &  pg35  &  ng4581 ) ;
 assign wire31447 = ( ng1917  &  pg35 ) ;
 assign wire31449 = ( pg35  &  wire6655 ) | ( pg35  &  ng14367  &  wire29571 ) ;
 assign wire31450 = ( ng1926  &  pg35 ) ;
 assign wire31452 = ( wire5505 ) | ( (~ ng27833)  &  wire31449 ) ;
 assign wire31454 = ( pg35  &  (~ ng676)  &  ng20375 ) ;
 assign wire31456 = ( pg35  &  ng676  &  (~ ng20375) ) ;
 assign wire31460 = ( (~ pg35)  &  ng1306 ) | ( pg35  &  (~ pg7946)  &  ng1532 ) ;
 assign wire31462 = ( pg35  &  (~ ng1389)  &  ng1351 ) ;
 assign wire31463 = ( ng1389  &  pg35 ) ;
 assign wire31464 = ( wire5490 ) | ( (~ ng13242)  &  (~ wire5491)  &  wire31462 ) ;
 assign wire31466 = ( pg35  &  (~ ng2250)  &  ng2246 ) ;
 assign wire31468 = ( ng2255  &  pg35 ) ;
 assign wire31470 = ( ng25432  &  wire31468 ) | ( ng2250  &  (~ ng2246)  &  (~ ng25432) ) ;
 assign wire31472 = ( pg35  &  (~ ng5489)  &  (~ ng5495) ) ;
 assign wire31474 = ( pg35  &  ng5489  &  ng5495 ) ;
 assign wire31477 = ( ng10838  &  wire31474 ) | ( pg35  &  ng5499  &  (~ ng10838) ) ;
 assign wire31478 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31479 = ( ng5917  &  pg35 ) ;
 assign wire31484 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31485 = ( ng3917  &  pg35 ) ;
 assign wire31488 = ( pg35  &  (~ ng2527)  &  (~ ng2533) ) ;
 assign wire31490 = ( pg35  &  ng2527  &  ng2533 ) ;
 assign wire31491 = ( ng2537  &  pg35 ) ;
 assign wire31494 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31495 = ( ng5268  &  pg35 ) ;
 assign wire31498 = ( pg35  &  ng3873  &  (~ ng3881)  &  ng3869 ) ;
 assign wire31499 = ( pg35  &  (~ ng3873)  &  ng3881 ) | ( pg35  &  ng3881  &  (~ ng3869) ) ;
 assign wire31501 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31502 = ( ng5256  &  pg35 ) ;
 assign wire31505 = ( ng930  &  (~ ng1193) ) | ( ng930  &  (~ ng969)  &  (~ ng1008) ) ;
 assign wire31508 = ( pg35  &  wire7041 ) | ( pg35  &  ng14367  &  wire29097 ) ;
 assign wire31509 = ( ng1648  &  pg35 ) ;
 assign wire31510 = ( ng1657  &  pg35 ) ;
 assign wire31512 = ( wire5431 ) | ( (~ ng27738)  &  wire31508 ) ;
 assign wire31513 = ( ng4035  &  pg35 ) ;
 assign wire31514 = ( pg35  &  wire7325 ) | ( pg35  &  wire7326 ) | ( pg35  &  wire28766 ) ;
 assign wire31515 = ( wire5428 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire31513 ) ;
 assign wire31521 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31522 = ( ng5603  &  pg35 ) ;
 assign wire31527 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31528 = ( ng3949  &  pg35 ) ;
 assign wire31530 = ( pg35  &  pg8291  &  ng218 ) ;
 assign wire31533 = ( ng4473  &  (~ ng4462) ) | ( ng4473  &  (~ ng4643) ) ;
 assign wire31534 = ( (~ pg35)  &  ng4473 ) | ( pg35  &  ng4473  &  ng4467 ) ;
 assign wire31536 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31537 = ( ng5236  &  pg35 ) ;
 assign wire31540 = ( pg35  &  (~ ng4849)  &  ng4843  &  ng4878 ) ;
 assign wire31542 = ( pg35  &  ng4849  &  (~ ng4843) ) | ( pg35  &  ng4849  &  (~ ng4878) ) ;
 assign wire31543 = ( wire5394 ) | ( ng31009  &  (~ ng10862)  &  wire31540 ) ;
 assign wire31544 = ( ng2227  &  pg35 ) ;
 assign wire31546 = ( wire5391 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire31544 ) ;
 assign wire31550 = ( (~ pg35)  &  ng5109 ) | ( pg35  &  pg9497  &  (~ pg9553)  &  (~ ng5109) ) ;
 assign wire31553 = ( pg35  &  pg12923  &  ng1280 ) ;
 assign wire31555 = ( (~ pg35)  &  ng1266 ) | ( pg35  &  (~ ng1280)  &  (~ ng15695) ) ;
 assign wire31556 = ( ng681  &  pg35 ) ;
 assign wire31557 = ( ng650  &  pg35 ) ;
 assign wire31559 = ( pg35  &  ng26703  &  ng11916 ) | ( pg35  &  ng17321  &  ng11916 ) ;
 assign wire31560 = ( ng2181  &  pg35 ) ;
 assign wire31563 = ( pg35  &  (~ ng1046)  &  ng1008 ) ;
 assign wire31564 = ( ng1046  &  pg35 ) ;
 assign wire31565 = ( wire5370 ) | ( (~ ng13211)  &  (~ wire5848)  &  wire31563 ) ;
 assign wire31570 = ( (~ ng2421) ) | ( (~ ng2495) ) ;
 assign wire31571 = ( pg35  &  ng26770  &  (~ wire31570) ) | ( pg35  &  ng17424  &  (~ wire31570) ) ;
 assign wire31572 = ( ng2441  &  pg35 ) ;
 assign wire31574 = ( ng4821  &  pg35 ) ;
 assign wire31575 = ( pg35  &  wire6832 ) | ( pg35  &  wire6833 ) | ( pg35  &  wire29346 ) ;
 assign wire31578 = ( (~ ng1768)  &  pg35 ) ;
 assign wire31581 = ( (~ pg35)  &  ng2767 ) | ( pg35  &  ng2779  &  (~ ng12377) ) ;
 assign wire31587 = ( (~ pg35)  &  ng936 ) | ( pg35  &  ng936  &  (~ ng907)  &  (~ ng15674) ) ;
 assign wire31589 = ( (~ pg35)  &  ng681 ) | ( pg35  &  ng699  &  ng8806 ) ;
 assign wire31591 = ( pg35  &  (~ ng3119)  &  (~ ng3125) ) ;
 assign wire31593 = ( ng3129  &  pg35 ) ;
 assign wire31595 = ( ng23067  &  wire31593 ) | ( ng3119  &  ng3125  &  (~ ng23067) ) ;
 assign wire31596 = ( ng4698  &  pg35 ) ;
 assign wire31597 = ( wire1421  &  ng4704 ) | ( ng4704  &  ng4818 ) | ( ng4704  &  (~ ng24374) ) ;
 assign wire31600 = ( ng29657  &  wire31597 ) | ( pg35  &  ng29657  &  ng30576 ) ;
 assign wire31604 = ( (~ pg35) ) | ( (~ ng4473)  &  ng4507 ) | ( ng4507  &  ng4459 ) ;
 assign wire31608 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31609 = ( ng5555  &  pg35 ) ;
 assign wire31610 = ( wire5322 ) | ( ng12453  &  ng12558  &  wire31608 ) ;
 assign wire31612 = ( pg35  &  (~ pg9048)  &  ng590 ) | ( pg35  &  ng590  &  ng559 ) ;
 assign wire31613 = ( (~ ng590)  &  pg35 ) ;
 assign wire31615 = ( ng1728 ) | ( (~ ng1772) ) ;
 assign wire31616 = ( pg35  &  ng17317  &  (~ wire31615) ) | ( pg35  &  ng26694  &  (~ wire31615) ) ;
 assign wire31617 = ( ng1752  &  pg35 ) ;
 assign wire31621 = ( pg35  &  (~ ng4375)  &  ng4382 ) ;
 assign wire31622 = ( pg35  &  ng4375  &  (~ ng4382) ) ;
 assign wire31623 = ( wire5310 ) | ( (~ wire29325)  &  wire31621 ) | ( (~ wire29326)  &  wire31621 ) ;
 assign wire31629 = ( (~ ng1802)  &  pg35 ) ;
 assign wire31631 = ( (~ ng28761)  &  ng17317  &  wire31629 ) | ( (~ ng28761)  &  ng26694  &  wire31629 ) ;
 assign wire31634 = ( pg35  &  ng990  &  (~ ng1008) ) | ( pg35  &  ng979  &  (~ ng1008) ) ;
 assign wire31637 = ( ng990  &  ng1008 ) | ( ng979  &  ng1008 ) ;
 assign wire31638 = ( pg35  &  ng1030  &  ng1018  &  (~ ng1046) ) ;
 assign wire31640 = ( pg35  &  ng979  &  ng996 ) | ( pg35  &  ng990  &  (~ ng979)  &  (~ ng996) ) ;
 assign wire31642 = ( wire5302 ) | ( wire31637  &  wire31638 ) ;
 assign wire31645 = ( ng225  &  pg35 ) ;
 assign wire31646 = ( pg14189  &  pg35 ) ;
 assign wire31650 = ( pg35  &  (~ ng5869)  &  ng5857  &  ng5863 ) ;
 assign wire31652 = ( pg35  &  ng153  &  ng23042 ) ;
 assign wire31653 = ( (~ ng153)  &  pg35 ) ;
 assign wire31655 = ( (~ ng2327)  &  pg35 ) ;
 assign wire31658 = ( (~ pg35)  &  ng2799 ) | ( pg35  &  ng2811  &  (~ ng12377) ) ;
 assign wire31659 = ( (~ ng4108)  &  pg35 ) ;
 assign wire31660 = ( ng4108  &  pg35 ) ;
 assign wire31661 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng4098 ) ;
 assign wire31662 = ( wire31661 ) | ( ng4098  &  ng22654  &  wire31659 ) ;
 assign wire31664 = ( pg35  &  ng5869  &  (~ ng5881)  &  ng5873 ) ;
 assign wire31665 = ( pg35  &  (~ ng5869)  &  ng5881 ) | ( pg35  &  ng5881  &  (~ ng5873) ) ;
 assign wire31667 = ( (~ ng1099)  &  pg35 ) ;
 assign wire31668 = ( ng1146  &  pg35 ) ;
 assign wire31671 = ( ng513  &  (~ ng667) ) | ( ng513  &  ng686 ) ;
 assign wire31672 = ( ng518  &  pg35 ) ;
 assign wire31677 = ( pg35  &  (~ ng4332)  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire31678 = ( (~ ng4340)  &  (~ ng4322)  &  (~ ng4311)  &  ng4643 ) ;
 assign wire31679 = ( ng5041  &  pg35 ) ;
 assign wire31681 = ( (~ ng5041)  &  pg35 ) ;
 assign wire31686 = ( (~ pg35)  &  ng1514 ) | ( pg35  &  (~ pg7946)  &  ng1526 ) | ( pg35  &  (~ ng1514)  &  ng1526 ) | ( pg35  &  pg7946  &  ng1514  &  (~ ng1526) ) ;
 assign wire31688 = ( pg35  &  (~ pg9048)  &  ng568 ) | ( pg35  &  ng568  &  ng559 ) ;
 assign wire31689 = ( (~ ng568)  &  pg35 ) ;
 assign wire31690 = ( wire5251 ) | ( (~ ng14708)  &  wire31688 ) | ( wire28793  &  wire31688 ) ;
 assign wire31696 = ( (~ pg72)  &  pg35  &  ng4581 ) | ( pg35  &  ng4578  &  ng4581 ) ;
 assign wire31697 = ( (~ pg35)  &  ng4567 ) | ( (~ ng4581)  &  ng4567 ) | ( pg73  &  pg35  &  ng4581 ) ;
 assign wire31701 = ( (~ pg35)  &  ng6148 ) | ( pg35  &  (~ pg9741)  &  pg9682  &  (~ ng6148) ) ;
 assign wire31702 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31703 = ( ng6283  &  pg35 ) ;
 assign wire31711 = ( (~ ng4322)  &  pg35 ) ;
 assign wire31712 = ( ng4311  &  (~ ng10511)  &  (~ ng8347)  &  wire31711 ) ;
 assign wire31713 = ( ng4322  &  pg35 ) ;
 assign wire31714 = ( (~ ng4311)  &  wire31713 ) | ( ng10511  &  wire31713 ) | ( ng8347  &  wire31713 ) ;
 assign wire31715 = ( wire5217 ) | ( (~ ng30583)  &  ng15591  &  wire31712 ) ;
 assign wire31716 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31717 = ( ng5252  &  pg35 ) ;
 assign wire31719 = ( (~ ng1274)  &  pg35 ) ;
 assign wire31720 = ( pg35  &  pg12923  &  ng1274 ) ;
 assign wire31726 = ( wire5201 ) | ( wire5202 ) | ( wire5203 ) | ( wire5204 ) ;
 assign wire31727 = ( wire5205 ) | ( wire5206 ) | ( wire5207 ) | ( wire5208 ) ;
 assign wire31729 = ( pg35  &  ng5033  &  ng15585 ) ;
 assign wire31731 = ( (~ pg35)  &  ng5029 ) | ( pg35  &  (~ ng5033)  &  (~ ng15585) ) ;
 assign wire31733 = ( pg35  &  ng3352  &  ng3288  &  ng3347 ) ;
 assign wire31734 = ( (~ ng4975)  &  (~ ng4899)  &  ng11283  &  wire31733 ) ;
 assign wire31736 = ( pg35  &  ng3352  &  (~ ng3288)  &  (~ ng3347) ) ;
 assign wire31737 = ( (~ ng4975)  &  (~ ng4899)  &  ng11283  &  wire31736 ) ;
 assign wire31739 = ( pg35  &  ng3343  &  (~ ng3352)  &  ng3288 ) ;
 assign wire31740 = ( (~ ng4975)  &  (~ ng4899)  &  ng11283  &  wire31739 ) ;
 assign wire31742 = ( pg35  &  (~ ng3343)  &  (~ ng3352)  &  (~ ng3288) ) ;
 assign wire31743 = ( (~ ng4975)  &  (~ ng4899)  &  ng11283  &  wire31742 ) ;
 assign wire31744 = ( ng4939  &  pg35 ) ;
 assign wire31746 = ( wire5196 ) | ( ng20887  &  wire31740 ) ;
 assign wire31747 = ( ng20887  &  wire31743 ) | ( pg35  &  ng4939  &  (~ ng20887) ) ;
 assign wire31748 = ( (~ ng23286)  &  wire31734 ) | ( (~ ng23286)  &  wire31737 ) ;
 assign wire31754 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31755 = ( ng5200  &  pg35 ) ;
 assign wire31756 = ( wire5183 ) | ( ng12772  &  ng12492  &  wire31754 ) ;
 assign wire31757 = ( ng4349  &  (~ ng4358)  &  (~ ng24380)  &  wire29233 ) ;
 assign wire31759 = ( (~ ng3352)  &  pg35 ) ;
 assign wire31761 = ( ng3352  &  pg35 ) ;
 assign wire31770 = ( (~ ng1906) ) | ( ng1936 ) ;
 assign wire31771 = ( pg35  &  ng26725  &  (~ wire31770) ) | ( pg35  &  ng17401  &  (~ wire31770) ) ;
 assign wire31772 = ( ng1878  &  pg35 ) ;
 assign wire31779 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31780 = ( ng5567  &  pg35 ) ;
 assign wire31783 = ( (~ pg35)  &  ng1246 ) | ( pg35  &  (~ pg17400)  &  pg10500 ) ;
 assign wire31784 = ( ng753  &  pg35 ) ;
 assign wire31788 = ( pg35  &  ng3171  &  (~ ng3179)  &  ng3167 ) ;
 assign wire31789 = ( pg35  &  (~ ng3171)  &  ng3179 ) | ( pg35  &  ng3179  &  (~ ng3167) ) ;
 assign wire31791 = ( (~ ng2811)  &  pg35 ) ;
 assign wire31792 = ( ng2724  &  (~ ng2729)  &  (~ ng11405)  &  wire31791 ) ;
 assign wire31794 = ( (~ ng111)  &  (~ ng11405)  &  (~ wire29805) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire29805) ) ;
 assign wire31795 = ( ng2807  &  pg35 ) ;
 assign wire31796 = ( wire5142 ) | ( ng11405  &  wire31795 ) | ( wire29805  &  wire31795 ) ;
 assign wire31797 = ( wire31796 ) | ( (~ ng111)  &  wire31792 ) | ( (~ ng29503)  &  wire31792 ) ;
 assign wire31798 = ( pg35  &  ng1668  &  ng1682 ) | ( pg35  &  ng1592  &  ng1682 ) ;
 assign wire31799 = ( ng26673  &  wire31798 ) | ( ng17292  &  wire31798 ) ;
 assign wire31800 = ( pg35  &  (~ ng1682) ) | ( pg35  &  (~ ng1668)  &  (~ ng1592) ) ;
 assign wire31801 = ( ng26673  &  wire31800 ) | ( ng17292  &  wire31800 ) ;
 assign wire31802 = ( ng1682  &  pg35 ) ;
 assign wire31803 = ( wire5136 ) | ( (~ ng26673)  &  (~ ng17292)  &  wire31802 ) ;
 assign wire31806 = ( pg35  &  (~ ng5827)  &  (~ ng5821) ) ;
 assign wire31808 = ( pg35  &  ng5827  &  ng5821 ) ;
 assign wire31811 = ( (~ ng23666)  &  wire31808 ) | ( pg35  &  ng5831  &  ng23666 ) ;
 assign wire31812 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31813 = ( ng3231  &  pg35 ) ;
 assign wire31815 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31816 = ( ng5579  &  pg35 ) ;
 assign wire31818 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31819 = ( ng6625  &  pg35 ) ;
 assign wire31821 = ( ng4392  &  ng4401 ) ;
 assign wire31822 = ( (~ pg35)  &  ng4401 ) | ( pg35  &  ng4411 ) ;
 assign wire31823 = ( ng29503  &  wire5887 ) | ( ng29503  &  ng14367  &  wire31005 ) ;
 assign wire31825 = ( pg35  &  ng110  &  ng2610 ) | ( pg35  &  ng110  &  (~ ng2619) ) ;
 assign wire31827 = ( pg35  &  (~ ng110)  &  (~ ng2610)  &  ng2619 ) ;
 assign wire31828 = ( ng2625  &  pg35 ) ;
 assign wire31829 = ( wire5107 ) | ( ng26236  &  wire31823  &  wire31825 ) ;
 assign wire31830 = ( (~ ng26236)  &  wire31828 ) | ( (~ wire31823)  &  wire31828 ) | ( ng26236  &  wire31823  &  wire31827 ) ;
 assign wire31831 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31832 = ( ng3897  &  pg35 ) ;
 assign wire31834 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31835 = ( ng6641  &  pg35 ) ;
 assign wire31838 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31839 = ( ng3538  &  pg35 ) ;
 assign wire31840 = ( wire5092 ) | ( ng8906  &  ng11571  &  wire31838 ) ;
 assign wire31842 = ( pg35  &  (~ ng6519)  &  (~ ng6513) ) ;
 assign wire31844 = ( pg35  &  ng6519  &  ng6513 ) ;
 assign wire31847 = ( (~ ng23733)  &  wire31844 ) | ( pg35  &  ng6523  &  ng23733 ) ;
 assign wire31848 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31849 = ( ng3263  &  pg35 ) ;
 assign wire31851 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31852 = ( ng3562  &  pg35 ) ;
 assign wire31854 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31855 = ( ng5937  &  pg35 ) ;
 assign wire31858 = ( pg35  &  ng6336  &  ng6395  &  ng6390 ) ;
 assign wire31859 = ( (~ ng4785)  &  ng4709  &  ng11261  &  wire31858 ) ;
 assign wire31861 = ( pg35  &  (~ ng6386)  &  (~ ng6336)  &  (~ ng6395) ) ;
 assign wire31862 = ( (~ ng4785)  &  ng4709  &  ng11261  &  wire31861 ) ;
 assign wire31864 = ( pg35  &  (~ ng6336)  &  ng6395  &  (~ ng6390) ) ;
 assign wire31865 = ( (~ ng4785)  &  ng4709  &  ng11261  &  wire31864 ) ;
 assign wire31867 = ( pg35  &  ng6386  &  ng6336  &  (~ ng6395) ) ;
 assign wire31868 = ( (~ ng4785)  &  ng4709  &  ng11261  &  wire31867 ) ;
 assign wire31870 = ( ng4771  &  pg35 ) ;
 assign wire31871 = ( wire5076 ) | ( ng21012  &  wire31862 ) ;
 assign wire31872 = ( ng21012  &  wire31868 ) | ( pg35  &  ng4771  &  (~ ng21012) ) ;
 assign wire31873 = ( (~ ng23949)  &  wire31859 ) | ( (~ ng23949)  &  wire31865 ) ;
 assign wire31875 = ( (~ ng4966)  &  pg35 ) ;
 assign wire31876 = ( ng4991  &  ng4983  &  ng10862  &  wire31875 ) ;
 assign wire31877 = ( ng4966  &  pg35 ) ;
 assign wire31878 = ( (~ ng4991)  &  wire31877 ) | ( (~ ng4983)  &  wire31877 ) | ( (~ ng10862)  &  wire31877 ) ;
 assign wire31879 = ( wire5070 ) | ( ng28349  &  ng13486  &  wire31876 ) ;
 assign wire31881 = ( pg35  &  (~ ng1199)  &  (~ ng10893)  &  wire29901 ) ;
 assign wire31883 = ( pg35  &  ng1199  &  ng10893 ) | ( pg35  &  ng1199  &  (~ wire29901) ) ;
 assign wire31885 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31886 = ( ng5941  &  pg35 ) ;
 assign wire31890 = ( pg35  &  ng1844 ) | ( pg35  &  ng1710 ) ;
 assign wire31891 = ( pg35  &  ng1858 ) | ( pg35  &  ng1724 ) ;
 assign wire31892 = ( pg35  &  ng2126 ) | ( pg35  &  ng1978 ) ;
 assign wire31893 = ( pg35  &  ng2112 ) | ( pg35  &  ng1992 ) ;
 assign wire31896 = ( pg35  &  ng2403 ) | ( pg35  &  ng2283 ) ;
 assign wire31897 = ( pg35  &  ng2537 ) | ( pg35  &  ng2685 ) ;
 assign wire31898 = ( pg35  &  ng2417 ) | ( pg35  &  ng2551 ) ;
 assign wire31899 = ( pg35  &  ng2269 ) | ( pg35  &  ng2671 ) ;
 assign wire31902 = ( pg35  &  ng2856 ) | ( (~ pg35)  &  ng2848 ) ;
 assign wire31906 = ( pg35  &  (~ ng1959)  &  ng1955 ) ;
 assign wire31908 = ( ng1964  &  pg35 ) ;
 assign wire31910 = ( ng25467  &  wire31908 ) | ( ng1959  &  (~ ng1955)  &  (~ ng25467) ) ;
 assign wire31913 = ( (~ ng1559)  &  pg35 ) ;
 assign wire31915 = ( ng1559  &  pg35 ) ;
 assign wire31917 = ( wire5024 ) | ( (~ ng11171)  &  (~ ng11149)  &  wire31913 ) ;
 assign wire31919 = ( pg35  &  ng4843  &  (~ ng4878) ) ;
 assign wire31920 = ( ng4878  &  (~ ng4843) ) ;
 assign wire31921 = ( wire5021 ) | ( ng31009  &  (~ ng10862)  &  wire31919 ) ;
 assign wire31922 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31923 = ( ng6657  &  pg35 ) ;
 assign wire31926 = ( pg35  &  ng4311  &  ng10511 ) | ( pg35  &  ng4311  &  ng8347 ) ;
 assign wire31928 = ( pg35  &  (~ ng4311)  &  (~ ng10511)  &  (~ ng8347) ) ;
 assign wire31929 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31930 = ( ng3223  &  pg35 ) ;
 assign wire31932 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31933 = ( ng3251  &  pg35 ) ;
 assign wire31935 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31936 = ( ng5619  &  pg35 ) ;
 assign wire31938 = ( (~ pg11678)  &  ng790 ) | ( ng790  &  ng736 ) ;
 assign wire31939 = ( (~ ng794) ) | ( pg11678  &  (~ ng736) ) ;
 assign wire31940 = ( (~ pg11678)  &  ng807 ) | ( ng736  &  ng807 ) ;
 assign wire31942 = ( pg35  &  (~ pg11678)  &  ng554 ) | ( pg35  &  ng554  &  ng736 ) ;
 assign wire31943 = ( (~ ng554)  &  pg35 ) ;
 assign wire31945 = ( ng29503  &  wire7257 ) | ( ng29503  &  ng14367  &  wire28834 ) ;
 assign wire31947 = ( pg35  &  ng110  &  ng1783 ) | ( pg35  &  ng110  &  (~ ng1792) ) ;
 assign wire31949 = ( pg35  &  (~ ng110)  &  (~ ng1783)  &  ng1792 ) ;
 assign wire31950 = ( ng1798  &  pg35 ) ;
 assign wire31951 = ( wire4999 ) | ( ng26166  &  wire31945  &  wire31947 ) ;
 assign wire31952 = ( (~ ng26166)  &  wire31950 ) | ( (~ wire31945)  &  wire31950 ) | ( ng26166  &  wire31945  &  wire31949 ) ;
 assign wire31954 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31955 = ( ng5901  &  pg35 ) ;
 assign wire31956 = ( wire4988 ) | ( ng12609  &  ng12515  &  wire31954 ) ;
 assign wire31958 = ( pg35  &  ng182  &  ng174 ) ;
 assign wire31960 = ( pg35  &  ng168  &  ng174 ) ;
 assign wire31962 = ( pg35  &  ng168  &  ng182 ) ;
 assign wire31965 = ( pg35  &  ng4653  &  (~ ng4688) ) ;
 assign wire31966 = ( ng4688  &  (~ ng4653) ) ;
 assign wire31967 = ( wire4982 ) | ( ng31003  &  (~ ng10831)  &  wire31965 ) ;
 assign wire31968 = ( ng1111  &  (~ ng1105) ) ;
 assign wire31970 = ( ng1105  &  pg35 ) ;
 assign wire31971 = ( (~ pg35)  &  ng1111 ) | ( pg35  &  ng1105  &  (~ ng1111) ) ;
 assign wire31972 = ( wire31971 ) | ( (~ ng10929)  &  (~ ng13260)  &  wire31968 ) ;
 assign wire31973 = ( ng3889  &  pg35 ) ;
 assign wire31974 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31975 = ( wire4972 ) | ( (~ ng11626)  &  wire31973 ) | ( (~ ng8958)  &  wire31973 ) ;
 assign wire31978 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng4093 ) ;
 assign wire31984 = ( (~ pg72)  &  pg35  &  ng4581 ) | ( pg35  &  ng4581  &  ng59 ) ;
 assign wire31985 = ( (~ pg35)  &  ng4501 ) | ( ng4501  &  (~ ng4581) ) | ( pg73  &  pg35  &  ng4581 ) ;
 assign wire31986 = ( ng93  &  (~ ng4349)  &  ng4358  &  ng29503 ) ;
 assign wire31989 = ( pg35  &  (~ ng5990)  &  (~ ng23932) ) ;
 assign wire31991 = ( pg35  &  ng5990  &  ng23932 ) ;
 assign wire31993 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31994 = ( ng6275  &  pg35 ) ;
 assign wire31996 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire31997 = ( ng6239  &  pg35 ) ;
 assign wire31998 = ( wire4952 ) | ( ng10421  &  ng12667  &  wire31996 ) ;
 assign wire32002 = ( (~ pg35)  &  ng5456 ) | ( pg35  &  pg9555  &  (~ pg9615)  &  (~ ng5456) ) ;
 assign wire32003 = ( ng150  &  pg35 ) ;
 assign wire32005 = ( (~ ng150)  &  pg35 ) ;
 assign wire32007 = ( wire1421  &  ng4749 ) | ( ng4818  &  ng4749 ) | ( ng4749  &  (~ ng24374) ) ;
 assign wire32011 = ( pg35  &  ng4743  &  (~ ng29672) ) | ( pg35  &  ng29672  &  ng30576 ) ;
 assign wire32012 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32013 = ( ng5571  &  pg35 ) ;
 assign wire32015 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32016 = ( ng5196  &  pg35 ) ;
 assign wire32017 = ( wire4934 ) | ( ng10266  &  ng12492  &  wire32015 ) ;
 assign wire32018 = ( pg35  &  wire7030 ) | ( pg35  &  ng14367  &  wire29111 ) ;
 assign wire32019 = ( ng2351  &  pg35 ) ;
 assign wire32020 = ( ng2342  &  pg35 ) ;
 assign wire32022 = ( wire4930 ) | ( (~ ng27854)  &  wire32018 ) ;
 assign wire32024 = ( pg35  &  (~ ng4392)  &  ng4430 ) ;
 assign wire32031 = ( (~ ng405)  &  ng437  &  ng392 ) | ( ng405  &  ng437  &  (~ ng392) ) ;
 assign wire32032 = ( ng405  &  ng401  &  ng392 ) | ( (~ ng405)  &  ng424  &  (~ ng392) ) ;
 assign wire32035 = ( ng182  &  (~ ng411)  &  (~ ng392) ) ;
 assign wire32039 = ( (~ ng441)  &  ng182  &  ng392 ) ;
 assign wire32043 = ( (~ ng182)  &  (~ ng411)  &  (~ ng392) ) ;
 assign wire32047 = ( (~ ng441)  &  (~ ng182)  &  ng392 ) ;
 assign wire32051 = ( wire4913 ) | ( wire4914 ) | ( wire4915 ) | ( wire4916 ) ;
 assign wire32052 = ( (~ ng11326)  &  pg35 ) ;
 assign wire32056 = ( (~ ng2518)  &  ng2504 ) | ( ng2476  &  (~ ng2453)  &  ng2504 ) ;
 assign wire32057 = ( ng2518  &  pg35 ) ;
 assign wire32058 = ( (~ pg35)  &  ng2504 ) | ( pg35  &  (~ ng2504)  &  ng22472  &  ng14713 ) ;
 assign wire32061 = ( pg35  &  (~ ng4616)  &  (~ ng30583)  &  (~ wire6408) ) ;
 assign wire32063 = ( pg35  &  ng4616  &  (~ ng30583)  &  (~ wire6408) ) ;
 assign wire32066 = ( pg35  &  (~ ng2518)  &  ng2514 ) ;
 assign wire32068 = ( ng2523  &  pg35 ) ;
 assign wire32070 = ( ng25495  &  wire32068 ) | ( ng2518  &  (~ ng2514)  &  (~ ng25495) ) ;
 assign wire32072 = ( pg35  &  (~ ng2541)  &  (~ ng2547) ) ;
 assign wire32074 = ( pg35  &  ng2541  &  ng2547 ) ;
 assign wire32077 = ( (~ ng25400)  &  wire32074 ) | ( pg35  &  ng2551  &  ng25400 ) ;
 assign wire32078 = ( ng2555 ) | ( (~ ng2599) ) ;
 assign wire32079 = ( ng2579  &  pg35 ) ;
 assign wire32080 = ( pg35  &  ng26793  &  (~ wire32078) ) | ( pg35  &  ng14506  &  (~ wire32078) ) ;
 assign wire32082 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32083 = ( ng3929  &  pg35 ) ;
 assign wire32085 = ( (~ ng2040) ) | ( ng2070 ) ;
 assign wire32086 = ( pg35  &  ng26759  &  (~ wire32085) ) | ( pg35  &  ng14438  &  (~ wire32085) ) ;
 assign wire32087 = ( ng2012  &  pg35 ) ;
 assign wire32091 = ( pg35  &  (~ ng4864)  &  (~ ng4871)  &  (~ ng4836) ) ;
 assign wire32093 = ( ng2108  &  pg35 ) ;
 assign wire32095 = ( ng2629 ) | ( (~ ng2599) ) ;
 assign wire32096 = ( pg35  &  ng26793  &  (~ wire32095) ) | ( pg35  &  ng14506  &  (~ wire32095) ) ;
 assign wire32097 = ( ng2571  &  pg35 ) ;
 assign wire32101 = ( ng2079  &  (~ ng2093) ) | ( ng2079  &  ng2051  &  (~ ng2028) ) ;
 assign wire32102 = ( ng2093  &  pg35 ) ;
 assign wire32103 = ( (~ pg35)  &  ng2079 ) | ( pg35  &  (~ ng2079)  &  ng22457  &  ng14712 ) ;
 assign wire32105 = ( (~ ng1554)  &  pg35 ) ;
 assign wire32107 = ( ng1554  &  pg35 ) ;
 assign wire32109 = ( wire4873 ) | ( (~ ng11171)  &  (~ ng13597)  &  wire32105 ) ;
 assign wire32110 = ( ng3207  &  pg35 ) ;
 assign wire32111 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32112 = ( wire4870 ) | ( (~ ng11473)  &  wire32110 ) | ( (~ ng11514)  &  wire32110 ) ;
 assign wire32117 = ( ng1193  &  pg35 ) ;
 assign wire32118 = ( (~ pg35)  &  ng1189 ) | ( pg35  &  (~ ng1070)  &  ng1193 ) ;
 assign wire32120 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32121 = ( ng3255  &  pg35 ) ;
 assign wire32123 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32124 = ( ng5893  &  pg35 ) ;
 assign wire32125 = ( wire4857 ) | ( ng12609  &  ng12824  &  wire32123 ) ;
 assign wire32126 = ( (~ ng1300)  &  ng1484 ) ;
 assign wire32127 = ( ng1300  &  pg35 ) ;
 assign wire32129 = ( (~ pg35)  &  ng1484 ) | ( pg35  &  (~ ng1484)  &  ng1300 ) ;
 assign wire32130 = ( wire32129 ) | ( (~ ng10939)  &  (~ ng10961)  &  wire32126 ) ;
 assign wire32133 = ( (~ pg35)  &  ng4549 ) | ( ng4549  &  (~ ng4581) ) ;
 assign wire32135 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32136 = ( ng3187  &  pg35 ) ;
 assign wire32137 = ( wire4839 ) | ( ng8864  &  ng11514  &  wire32135 ) ;
 assign wire32138 = ( (~ ng2040) ) | ( ng1996 ) ;
 assign wire32139 = ( (~ ng2070)  &  pg35 ) ;
 assign wire32141 = ( ng26759  &  (~ ng28833)  &  wire32139 ) | ( ng14438  &  (~ ng28833)  &  wire32139 ) ;
 assign wire32145 = ( (~ pg16744)  &  (~ pg16656) ) ;
 assign wire32146 = ( pg35  &  (~ pg13926)  &  (~ pg14451)  &  (~ pg16627) ) ;
 assign wire32151 = ( pg35  &  pg13926  &  (~ pg14451)  &  pg11388 ) ;
 assign wire32154 = ( ng269  &  ng255 ) ;
 assign wire32155 = ( (~ pg73)  &  (~ pg72)  &  pg35 ) ;
 assign wire32158 = ( pg73  &  (~ pg72)  &  pg35 ) ;
 assign wire32166 = ( (~ pg35)  &  ng102 ) | ( wire32154  &  wire32155 ) ;
 assign wire32167 = ( wire4826 ) | ( ng262  &  ng255  &  wire32158 ) ;
 assign wire32170 = ( (~ ng6381)  &  pg17845 ) ;
 assign wire32171 = ( ng6336  &  ng6395  &  ng6271 ) ;
 assign wire32172 = ( ng6381  &  pg17743 ) ;
 assign wire32173 = ( ng6336  &  ng6295  &  ng6395 ) ;
 assign wire32175 = ( pg17760  &  ng6283  &  ng6336  &  ng6395 ) ;
 assign wire32176 = ( ng6381  &  pg17845 ) ;
 assign wire32177 = ( (~ ng6336)  &  ng6395  &  ng6263 ) ;
 assign wire32179 = ( pg17649  &  ng6299  &  (~ ng6336)  &  (~ ng6395) ) ;
 assign wire32180 = ( ng6381  &  pg13085 ) ;
 assign wire32181 = ( ng6235  &  (~ ng6336)  &  (~ ng6395) ) ;
 assign wire32182 = ( ng6243  &  ng6381 ) ;
 assign wire32183 = ( (~ ng6336)  &  (~ ng6395)  &  ng6377 ) ;
 assign wire32185 = ( pg14779  &  ng6267  &  ng6336  &  (~ ng6395) ) ;
 assign wire32186 = ( (~ ng6381)  &  pg13085 ) ;
 assign wire32187 = ( ng6247  &  ng6336  &  (~ ng6395) ) ;
 assign wire32188 = ( ng6381  &  pg14705 ) ;
 assign wire32189 = ( ng6279  &  ng6336  &  (~ ng6395) ) ;
 assign wire32190 = ( ng6381  &  pg12422 ) ;
 assign wire32191 = ( ng6239  &  (~ ng6336)  &  ng6395 ) ;
 assign wire32192 = ( (~ ng6381)  &  pg17685 ) ;
 assign wire32193 = ( ng6251  &  (~ ng6336)  &  ng6395 ) ;
 assign wire32194 = ( wire32170  &  wire32171 ) | ( wire32172  &  wire32173 ) ;
 assign wire32195 = ( (~ ng12423)  &  wire32175 ) | ( wire32176  &  wire32177 ) ;
 assign wire32196 = ( (~ ng12423)  &  wire32179 ) | ( wire32180  &  wire32181 ) ;
 assign wire32197 = ( wire32182  &  wire32183 ) | ( (~ ng12423)  &  wire32185 ) ;
 assign wire32198 = ( wire32186  &  wire32187 ) | ( wire32188  &  wire32189 ) ;
 assign wire32199 = ( wire32190  &  wire32191 ) | ( wire32192  &  wire32193 ) ;
 assign wire32202 = ( wire32199 ) | ( wire32198 ) ;
 assign wire32203 = ( wire32194 ) | ( wire32195 ) | ( wire32196 ) | ( wire32197 ) ;
 assign wire32204 = ( ng6381  &  pg17685 ) ;
 assign wire32205 = ( ng6311  &  ng6336  &  ng6395 ) ;
 assign wire32206 = ( ng6255  &  pg12422 ) ;
 assign wire32207 = ( (~ ng6381)  &  ng6336  &  ng6395 ) ;
 assign wire32208 = ( (~ ng6381)  &  pg14705 ) ;
 assign wire32209 = ( (~ ng6336)  &  (~ ng6395)  &  ng6287 ) ;
 assign wire32211 = ( pg14779  &  ng6275  &  (~ ng6336)  &  (~ ng6395) ) ;
 assign wire32212 = ( ng6377  &  (~ ng6381) ) ;
 assign wire32213 = ( ng6336  &  (~ ng6395)  &  ng6259 ) ;
 assign wire32215 = ( pg17760  &  (~ ng6336)  &  ng6395  &  ng6291 ) ;
 assign wire32217 = ( pg17649  &  ng6307  &  ng6336  &  (~ ng6395) ) ;
 assign wire32218 = ( ng6303  &  pg17743 ) ;
 assign wire32219 = ( (~ ng6381)  &  (~ ng6336)  &  ng6395 ) ;
 assign wire32220 = ( wire32204  &  wire32205 ) | ( wire32206  &  wire32207 ) ;
 assign wire32221 = ( wire32208  &  wire32209 ) | ( ng12423  &  wire32211 ) ;
 assign wire32222 = ( wire32212  &  wire32213 ) | ( ng12423  &  wire32215 ) ;
 assign wire32223 = ( ng12423  &  wire32217 ) | ( wire32218  &  wire32219 ) ;
 assign wire32226 = ( wire32220 ) | ( wire32221 ) | ( wire32222 ) | ( wire32223 ) ;
 assign wire32228 = ( pg35  &  (~ ng6154)  &  ng21012 ) | ( pg35  &  ng11160  &  ng21012 ) ;
 assign wire32230 = ( pg35  &  ng6154  &  (~ ng11160)  &  ng21012 ) ;
 assign wire32231 = ( ng6154  &  pg35 ) ;
 assign wire32234 = ( ng5264  &  pg35 ) ;
 assign wire32235 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32239 = ( ng4349  &  ng4358  &  (~ ng24380)  &  wire29233 ) ;
 assign wire32242 = ( pg35  &  (~ ng4054)  &  wire28765 ) | ( pg35  &  (~ ng4054)  &  wire28766 ) ;
 assign wire32243 = ( ng4054  &  pg35 ) ;
 assign wire32244 = ( wire4783 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire32243 ) ;
 assign wire32251 = ( ng4785  &  (~ ng4776)  &  ng4709 ) ;
 assign wire32252 = ( pg35  &  (~ ng4801)  &  (~ ng4674)  &  (~ ng4681) ) ;
 assign wire32253 = ( (~ ng4646)  &  (~ ng4737)  &  (~ ng4793)  &  (~ ng4688) ) ;
 assign wire32259 = ( pg35  &  (~ ng4801)  &  ng4785  &  (~ ng4709) ) ;
 assign wire32260 = ( (~ ng4674)  &  (~ ng4681)  &  (~ ng4646)  &  (~ ng4793) ) ;
 assign wire32266 = ( pg35  &  (~ ng4801)  &  (~ ng4785)  &  ng4709 ) ;
 assign wire32267 = ( (~ ng4674)  &  (~ ng4681)  &  (~ ng4646)  &  (~ ng4793) ) ;
 assign wire32269 = ( (~ ng4785)  &  ng4698  &  (~ ng4709) ) | ( ng4785  &  ng4743  &  (~ ng4709) ) ;
 assign wire32270 = ( ng4765  &  ng4785  &  ng4709 ) | ( (~ ng4785)  &  ng4754  &  ng4709 ) ;
 assign wire32271 = ( (~ ng4785)  &  ng4722  &  (~ ng4709) ) | ( ng4785  &  ng4717  &  (~ ng4709) ) ;
 assign wire32272 = ( ng4727  &  ng4785  &  ng4709 ) | ( (~ ng4785)  &  ng4732  &  ng4709 ) ;
 assign wire32275 = ( pg35  &  (~ ng4674)  &  (~ ng4688) ) ;
 assign wire32277 = ( (~ ng4681)  &  (~ ng4646)  &  (~ ng11155)  &  wire32275 ) ;
 assign wire32281 = ( pg35  &  (~ ng4674)  &  (~ ng4688) ) ;
 assign wire32283 = ( (~ ng4681)  &  (~ ng4646)  &  (~ ng11155)  &  wire32281 ) ;
 assign wire32288 = ( pg35  &  (~ ng4674)  &  (~ ng4776) ) ;
 assign wire32289 = ( (~ ng4681)  &  (~ ng4646)  &  ng4793  &  (~ ng4688) ) ;
 assign wire32293 = ( pg35  &  (~ ng4674)  &  (~ ng4688) ) ;
 assign wire32301 = ( wire4766 ) | ( wire4767 ) | ( wire4768 ) | ( wire4769 ) ;
 assign wire32304 = ( wire4764 ) | ( wire32301 ) ;
 assign wire32305 = ( wire4759 ) | ( wire4760 ) | ( wire4761 ) | ( wire4765 ) ;
 assign wire32306 = ( ng16663  &  (~ ng16728)  &  wire32277 ) | ( (~ ng16663)  &  ng16728  &  wire32283 ) ;
 assign wire32313 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32314 = ( ng6311  &  pg35 ) ;
 assign wire32316 = ( ng4826  &  pg35 ) ;
 assign wire32317 = ( pg35  &  wire7248 ) | ( pg35  &  wire7249 ) | ( pg35  &  wire28843 ) ;
 assign wire32323 = ( pg35  &  (~ ng1691)  &  ng1687 ) ;
 assign wire32325 = ( ng1696  &  pg35 ) ;
 assign wire32327 = ( ng25382  &  wire32325 ) | ( ng1691  &  (~ ng1687)  &  (~ ng25382) ) ;
 assign wire32328 = ( ng3578  &  pg35 ) ;
 assign wire32329 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32331 = ( ng2380  &  pg35 ) ;
 assign wire32333 = ( ng2648  &  pg35 ) ;
 assign wire32336 = ( pg35  &  (~ ng4601)  &  ng4593  &  ng24411 ) ;
 assign wire32338 = ( pg35  &  ng4601  &  (~ ng4593) ) | ( pg35  &  ng4601  &  (~ ng24411) ) ;
 assign wire32340 = ( pg35  &  ng26793  &  ng9835 ) | ( pg35  &  ng14506  &  ng9835 ) ;
 assign wire32341 = ( ng2567  &  pg35 ) ;
 assign wire32344 = ( pg35  &  ng862  &  (~ ng8721) ) ;
 assign wire32345 = ( ng862  &  pg35 ) ;
 assign wire32348 = ( pg35  &  ng862  &  ng703 ) ;
 assign wire32350 = ( (~ pg35)  &  ng446 ) | ( pg35  &  ng896  &  ng890 ) ;
 assign wire32352 = ( wire32350 ) | ( (~ ng8721)  &  ng11326  &  wire32345 ) ;
 assign wire32353 = ( wire4708 ) | ( wire32352 ) | ( (~ ng8721)  &  wire32348 ) ;
 assign wire32354 = ( pg35  &  ng3817 ) | ( pg35  &  ng3466 ) ;
 assign wire32355 = ( pg35  &  ng4427 ) | ( pg35  &  ng4420 ) | ( pg35  &  ng3115 ) ;
 assign wire32357 = ( pg35  &  ng5124 ) | ( pg35  &  ng5817 ) ;
 assign wire32358 = ( pg35  &  ng6509 ) | ( pg35  &  ng6163 ) | ( pg35  &  ng5471 ) ;
 assign wire32363 = ( (~ ng2273)  &  pg35 ) ;
 assign wire32364 = ( ng2273  &  pg35 ) ;
 assign wire32367 = ( pg35  &  ng6215  &  (~ ng6227)  &  ng6219 ) ;
 assign wire32368 = ( pg35  &  (~ ng6215)  &  ng6227 ) | ( pg35  &  ng6227  &  (~ ng6219) ) ;
 assign wire32377 = ( pg35  &  (~ ng4332)  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire32378 = ( (~ ng4584)  &  ng4340  &  (~ ng4322)  &  (~ ng4311) ) ;
 assign wire32379 = ( (~ ng4616)  &  (~ ng4601)  &  (~ ng4608)  &  (~ ng4593) ) ;
 assign wire32382 = ( pg35  &  ng9649  &  ng26703 ) | ( pg35  &  ng9649  &  ng17321 ) ;
 assign wire32383 = ( ng2165  &  pg35 ) ;
 assign wire32385 = ( ng4141 ) | ( ng4064 ) | ( ng4057 ) | ( ng4082 ) ;
 assign wire32386 = ( ng4112  &  pg35 ) ;
 assign wire32387 = ( wire4681 ) | ( (~ ng13806)  &  wire32386 ) | ( wire32385  &  wire32386 ) ;
 assign wire32388 = ( (~ ng1982)  &  pg35 ) ;
 assign wire32389 = ( ng1982  &  pg35 ) ;
 assign wire32391 = ( ng3215  &  pg35 ) ;
 assign wire32392 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32395 = ( ng1367  &  pg35 ) ;
 assign wire32396 = ( (~ pg35)  &  ng1361 ) | ( pg35  &  (~ ng25917)  &  wire4669 ) ;
 assign wire32398 = ( pg35  &  wire6319 ) | ( pg35  &  ng14367  &  wire30342 ) ;
 assign wire32399 = ( ng2051  &  pg35 ) ;
 assign wire32401 = ( wire4664 ) | ( (~ ng27882)  &  wire32398 ) ;
 assign wire32404 = ( ng1677  &  (~ ng1691) ) | ( ng1677  &  (~ ng1624)  &  ng1648 ) ;
 assign wire32405 = ( ng1691  &  pg35 ) ;
 assign wire32406 = ( (~ pg35)  &  ng1677 ) | ( pg35  &  (~ ng1677)  &  ng22342  &  ng14611 ) ;
 assign wire32408 = ( ng1105  &  pg35 ) ;
 assign wire32409 = ( ng1146  &  ng1111 ) | ( ng1111  &  ng1099 ) ;
 assign wire32412 = ( (~ ng1105)  &  pg35 ) ;
 assign wire32413 = ( ng1146  &  ng1111 ) | ( ng1111  &  ng1099 ) ;
 assign wire32417 = ( pg35  &  (~ ng1146)  &  ng1105  &  (~ ng1099) ) ;
 assign wire32420 = ( pg35  &  (~ ng1146)  &  (~ ng1105)  &  (~ ng1099) ) ;
 assign wire32423 = ( (~ pg35)  &  ng1135 ) | ( pg35  &  ng1111  &  ng13260 ) ;
 assign wire32424 = ( (~ ng13336)  &  (~ ng13260)  &  wire32417 ) | ( ng13336  &  (~ ng13260)  &  wire32420 ) ;
 assign wire32431 = ( pg35  &  (~ ng417)  &  (~ ng8806) ) ;
 assign wire32432 = ( (~ ng8806)  &  ng417 ) ;
 assign wire32434 = ( (~ pg35)  &  ng417 ) | ( pg35  &  ng411  &  ng8806 ) ;
 assign wire32438 = ( (~ ng2587) ) | ( (~ ng2619) ) ;
 assign wire32443 = ( pg35  &  ng4639  &  (~ ng4628)  &  ng4621 ) ;
 assign wire32445 = ( pg35  &  (~ ng4639)  &  ng4628 ) | ( pg35  &  ng4628  &  (~ ng4621) ) ;
 assign wire32447 = ( (~ ng2767)  &  pg35 ) ;
 assign wire32448 = ( (~ ng2724)  &  (~ ng2729)  &  (~ ng11405)  &  wire32447 ) ;
 assign wire32450 = ( (~ ng85)  &  ng12026  &  (~ ng11405) ) | ( (~ ng29503)  &  ng12026  &  (~ ng11405) ) ;
 assign wire32451 = ( ng2771  &  pg35 ) ;
 assign wire32452 = ( wire4630 ) | ( (~ ng12026)  &  wire32451 ) | ( ng11405  &  wire32451 ) ;
 assign wire32453 = ( wire32452 ) | ( (~ ng85)  &  wire32448 ) | ( (~ ng29503)  &  wire32448 ) ;
 assign wire32454 = ( ng3570  &  pg35 ) ;
 assign wire32455 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32458 = ( pg35  &  (~ pg9048)  &  ng622 ) | ( pg35  &  ng559  &  ng622 ) ;
 assign wire32459 = ( (~ ng622)  &  pg35 ) ;
 assign wire32460 = ( wire4623 ) | ( (~ ng33851)  &  wire32458 ) | ( wire30331  &  wire32458 ) ;
 assign wire32462 = ( (~ pg35)  &  ng2927 ) | ( pg35  &  ng4153 ) ;
 assign wire32463 = ( ng4760  &  pg35 ) ;
 assign wire32464 = ( wire1421  &  wire32463 ) | ( ng4818  &  wire32463 ) | ( (~ ng24374)  &  wire32463 ) ;
 assign wire32466 = ( pg35  &  ng101  &  ng24374  &  (~ wire29730) ) ;
 assign wire32468 = ( ng29694  &  wire32466 ) | ( pg35  &  ng4754  &  (~ ng29694) ) ;
 assign wire32470 = ( pg35  &  ng4983  &  (~ ng10862) ) ;
 assign wire32472 = ( pg35  &  (~ ng4983)  &  ng10862 ) ;
 assign wire32473 = ( wire4604 ) | ( ng28349  &  ng13486  &  wire32470 ) ;
 assign wire32475 = ( pg35  &  (~ ng4049)  &  ng4054  &  (~ ng3990) ) ;
 assign wire32476 = ( (~ ng4975)  &  ng4899  &  ng11283  &  wire32475 ) ;
 assign wire32478 = ( pg35  &  (~ ng4045)  &  (~ ng4054)  &  (~ ng3990) ) ;
 assign wire32479 = ( (~ ng4975)  &  ng4899  &  ng11283  &  wire32478 ) ;
 assign wire32481 = ( pg35  &  ng4049  &  ng4054  &  ng3990 ) ;
 assign wire32482 = ( (~ ng4975)  &  ng4899  &  ng11283  &  wire32481 ) ;
 assign wire32484 = ( pg35  &  ng4045  &  (~ ng4054)  &  ng3990 ) ;
 assign wire32485 = ( (~ ng4975)  &  ng4899  &  ng11283  &  wire32484 ) ;
 assign wire32486 = ( ng4961  &  pg35 ) ;
 assign wire32487 = ( ng4961  &  pg35 ) ;
 assign wire32488 = ( wire4600 ) | ( wire28765  &  wire32479 ) | ( wire28766  &  wire32479 ) ;
 assign wire32489 = ( wire28765  &  wire32485 ) | ( wire28766  &  wire32485 ) | ( (~ wire28765)  &  (~ wire28766)  &  wire32487 ) ;
 assign wire32493 = ( pg35  &  (~ ng3484)  &  (~ ng3490) ) ;
 assign wire32495 = ( pg35  &  ng3484  &  ng3490 ) ;
 assign wire32498 = ( ng12692  &  wire32495 ) | ( pg35  &  ng3494  &  (~ ng12692) ) ;
 assign wire32500 = ( pg35  &  ng5703  &  (~ ng5698)  &  (~ ng5644) ) ;
 assign wire32501 = ( (~ ng4785)  &  (~ ng4709)  &  ng11261  &  wire32500 ) ;
 assign wire32503 = ( pg35  &  (~ ng5703)  &  (~ ng5694)  &  (~ ng5644) ) ;
 assign wire32504 = ( (~ ng4785)  &  (~ ng4709)  &  ng11261  &  wire32503 ) ;
 assign wire32506 = ( pg35  &  (~ ng5703)  &  ng5694  &  ng5644 ) ;
 assign wire32507 = ( (~ ng4785)  &  (~ ng4709)  &  ng11261  &  wire32506 ) ;
 assign wire32509 = ( pg35  &  ng5703  &  ng5698  &  ng5644 ) ;
 assign wire32510 = ( (~ ng4785)  &  (~ ng4709)  &  ng11261  &  wire32509 ) ;
 assign wire32511 = ( ng4749  &  pg35 ) ;
 assign wire32513 = ( wire4590 ) | ( ng20739  &  wire32504 ) ;
 assign wire32514 = ( ng20739  &  wire32507 ) | ( pg35  &  ng4749  &  (~ ng20739) ) ;
 assign wire32515 = ( (~ ng23909)  &  wire32501 ) | ( (~ ng23909)  &  wire32510 ) ;
 assign wire32517 = ( ng2421  &  pg35 ) ;
 assign wire32521 = ( (~ ng1802) ) | ( (~ ng1728) ) ;
 assign wire32522 = ( pg35  &  ng17317  &  (~ wire32521) ) | ( pg35  &  ng26694  &  (~ wire32521) ) ;
 assign wire32523 = ( ng1748  &  pg35 ) ;
 assign wire32526 = ( pg35  &  (~ pg11678)  &  ng758 ) | ( pg35  &  ng758  &  ng736 ) ;
 assign wire32527 = ( (~ ng758)  &  pg35 ) ;
 assign wire32529 = ( ng29503  &  wire7041 ) | ( ng29503  &  ng14367  &  wire29097 ) ;
 assign wire32531 = ( pg35  &  ng110  &  (~ ng1657) ) | ( pg35  &  ng110  &  ng1648 ) ;
 assign wire32533 = ( pg35  &  (~ ng110)  &  ng1657  &  (~ ng1648) ) ;
 assign wire32534 = ( ng1664  &  pg35 ) ;
 assign wire32535 = ( wire4574 ) | ( ng26148  &  wire32529  &  wire32531 ) ;
 assign wire32536 = ( (~ ng26148)  &  wire32534 ) | ( (~ wire32529)  &  wire32534 ) | ( ng26148  &  wire32529  &  wire32533 ) ;
 assign wire32538 = ( pg35  &  (~ ng667)  &  ng528 ) | ( pg35  &  ng528  &  ng686 ) ;
 assign wire32539 = ( pg35  &  (~ ng667) ) | ( pg35  &  ng686 ) ;
 assign wire32540 = ( (~ ng513)  &  ng518  &  ng11607  &  wire32539 ) ;
 assign wire32541 = ( wire4570 ) | ( (~ ng11607)  &  wire32538 ) | ( (~ ng12812)  &  wire32538 ) ;
 assign wire32542 = ( pg35  &  ng1964 ) | ( pg35  &  ng1830 ) ;
 assign wire32543 = ( pg35  &  ng2098 ) | ( pg35  &  ng1696 ) ;
 assign wire32544 = ( pg35  &  ng2523 ) | ( pg35  &  ng2657 ) ;
 assign wire32545 = ( pg35  &  ng2255 ) | ( pg35  &  ng2389 ) ;
 assign wire32550 = ( ng962  &  pg35 ) ;
 assign wire32551 = ( ng996  &  pg35 ) ;
 assign wire32554 = ( pg35  &  (~ ng3821)  &  (~ ng3827) ) ;
 assign wire32555 = ( ng3831  &  pg35 ) ;
 assign wire32556 = ( ng3827  &  ng3821 ) ;
 assign wire32560 = ( pg35  &  (~ ng4793)  &  ng10831 ) ;
 assign wire32562 = ( pg35  &  ng4793  &  (~ ng10831) ) ;
 assign wire32563 = ( wire4537 ) | ( ng28336  &  ng13464  &  wire32560 ) ;
 assign wire32565 = ( pg35  &  (~ ng5808)  &  ng20875 ) | ( pg35  &  ng20875  &  ng11139 ) ;
 assign wire32567 = ( pg35  &  ng5808  &  ng20875  &  (~ ng11139) ) ;
 assign wire32568 = ( ng5808  &  pg35 ) ;
 assign wire32571 = ( ng1890  &  pg35 ) ;
 assign wire32572 = ( pg35  &  ng26725  &  ng11937 ) | ( pg35  &  ng17401  &  ng11937 ) ;
 assign wire32574 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32575 = ( ng5897  &  pg35 ) ;
 assign wire32578 = ( pg35  &  ng2841  &  (~ ng4093) ) ;
 assign wire32580 = ( pg35  &  ng2841  &  ng4093 ) ;
 assign wire32582 = ( pg35  &  wire5887 ) | ( pg35  &  ng14367  &  wire31005 ) ;
 assign wire32583 = ( ng2619  &  pg35 ) ;
 assign wire32584 = ( ng2610  &  pg35 ) ;
 assign wire32586 = ( wire4515 ) | ( (~ ng27933)  &  wire32582 ) ;
 assign wire32589 = ( (~ ng1413)  &  pg35 ) ;
 assign wire32590 = ( ng1542  &  (~ ng10918)  &  wire28896  &  wire32589 ) ;
 assign wire32591 = ( ng1413  &  pg35 ) ;
 assign wire32592 = ( (~ ng1542)  &  wire32591 ) | ( ng10918  &  wire32591 ) | ( (~ wire28896)  &  wire32591 ) ;
 assign wire32594 = ( (~ ng2331) ) | ( ng2287 ) ;
 assign wire32595 = ( pg35  &  ng17405  &  (~ wire32594) ) | ( pg35  &  ng26737  &  (~ wire32594) ) ;
 assign wire32596 = ( ng2311  &  pg35 ) ;
 assign wire32599 = ( pg35  &  (~ pg11678)  &  ng794 ) | ( pg35  &  ng794  &  ng736 ) ;
 assign wire32600 = ( (~ ng794)  &  pg35 ) ;
 assign wire32601 = ( wire4499 ) | ( ng34162  &  wire32599 ) | ( (~ wire31938)  &  wire32599 ) ;
 assign wire32602 = ( ng2667  &  pg35 ) ;
 assign wire32604 = ( (~ ng2629)  &  pg35 ) ;
 assign wire32606 = ( (~ ng28880)  &  ng26793  &  wire32604 ) | ( (~ ng28880)  &  ng14506  &  wire32604 ) ;
 assign wire32609 = ( pg35  &  ng26673  &  (~ wire31143) ) | ( pg35  &  ng17292  &  (~ wire31143) ) ;
 assign wire32610 = ( ng1616  &  pg35 ) ;
 assign wire32612 = ( ng255  &  pg35 ) ;
 assign wire32613 = ( pg14201  &  pg35 ) ;
 assign wire32616 = ( pg35  &  (~ pg9048)  &  ng613 ) | ( pg35  &  ng559  &  ng613 ) ;
 assign wire32617 = ( (~ ng613)  &  pg35 ) ;
 assign wire32619 = ( (~ ng817)  &  pg35 ) ;
 assign wire32621 = ( ng817  &  pg35 ) ;
 assign wire32623 = ( wire4470 ) | ( (~ ng8806)  &  (~ ng14279)  &  wire32619 ) ;
 assign wire32624 = ( ng686  &  pg35 ) ;
 assign wire32625 = ( ng691 ) | ( (~ ng703) ) ;
 assign wire32626 = ( pg35  &  ng385  &  ng358  &  (~ ng376) ) ;
 assign wire32628 = ( ng4955  &  pg35 ) ;
 assign wire32629 = ( wire1421  &  ng4961 ) | ( ng4818  &  ng4961 ) | ( ng4961  &  (~ ng24374) ) ;
 assign wire32630 = ( pg35  &  ng71  &  ng24374  &  (~ wire28575) ) ;
 assign wire32632 = ( ng29737  &  wire32629 ) | ( ng29737  &  wire32630 ) ;
 assign wire32633 = ( (~ ng2675)  &  pg35 ) ;
 assign wire32634 = ( ng2675  &  pg35 ) ;
 assign wire32636 = ( ng2533  &  pg35 ) ;
 assign wire32638 = ( ng6299  &  pg35 ) ;
 assign wire32639 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32642 = ( pg35  &  (~ ng1361)  &  ng1351 ) | ( pg35  &  ng1351  &  (~ ng1373) ) ;
 assign wire32644 = ( pg35  &  (~ ng1361)  &  ng1351 ) | ( pg35  &  ng1351  &  (~ ng1373) ) ;
 assign wire32647 = ( wire4429 ) | ( wire4431 ) | ( ng13242  &  wire32644 ) ;
 assign wire32651 = ( pg35  &  ng2070  &  ng2084 ) | ( pg35  &  ng1996  &  ng2084 ) ;
 assign wire32652 = ( ng26759  &  wire32651 ) | ( ng14438  &  wire32651 ) ;
 assign wire32653 = ( pg35  &  (~ ng2084) ) | ( pg35  &  (~ ng2070)  &  (~ ng1996) ) ;
 assign wire32654 = ( ng26759  &  wire32653 ) | ( ng14438  &  wire32653 ) ;
 assign wire32655 = ( ng2084  &  pg35 ) ;
 assign wire32656 = ( wire4421 ) | ( (~ ng26759)  &  (~ ng14438)  &  wire32655 ) ;
 assign wire32661 = ( pg35  &  (~ ng691)  &  ng11607 ) ;
 assign wire32662 = ( ng691  &  pg35 ) ;
 assign wire32664 = ( wire4414 ) | ( wire4417 ) | ( (~ ng11607)  &  wire32662 ) ;
 assign wire32665 = ( (~ ng4521)  &  pg35 ) ;
 assign wire32667 = ( (~ pg35)  &  ng4527 ) | ( pg35  &  ng4515  &  ng4521 ) ;
 assign wire32668 = ( (~ ng1862) ) | ( (~ ng1936) ) ;
 assign wire32669 = ( ng1882  &  pg35 ) ;
 assign wire32670 = ( pg35  &  ng26725  &  (~ wire32668) ) | ( pg35  &  ng17401  &  (~ wire32668) ) ;
 assign wire32672 = ( ng93  &  ng4349  &  ng4358  &  ng29503 ) ;
 assign wire32675 = ( pg35  &  (~ ng6336)  &  (~ ng23949) ) ;
 assign wire32677 = ( pg35  &  ng6336  &  ng23949 ) ;
 assign wire32683 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng4082 ) ;
 assign wire32689 = ( (~ pg35)  &  ng962 ) | ( pg35  &  pg7916  &  ng1178 ) ;
 assign wire32694 = ( ng3965  &  pg35 ) ;
 assign wire32695 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32699 = ( (~ ng914)  &  pg35 ) ;
 assign wire32700 = ( pg35  &  pg12919  &  ng914 ) ;
 assign wire32702 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32703 = ( ng5551  &  pg35 ) ;
 assign wire32706 = ( ng1373  &  pg35 ) ;
 assign wire32707 = ( wire4361 ) | ( ng25917  &  wire32706 ) | ( wire4669  &  wire32706 ) ;
 assign wire32708 = ( (~ ng626) ) | ( pg9048  &  (~ ng559) ) ;
 assign wire32710 = ( pg35  &  (~ pg9048)  &  ng632 ) | ( pg35  &  ng559  &  ng632 ) ;
 assign wire32711 = ( (~ ng632)  &  pg35 ) ;
 assign wire32717 = ( pg72  &  pg35  &  ng4581 ) | ( pg35  &  ng4581  &  ng59 ) ;
 assign wire32718 = ( (~ pg35)  &  ng4495 ) | ( ng4495  &  (~ ng4581) ) | ( (~ pg73)  &  pg35  &  ng4581 ) ;
 assign wire32719 = ( pg35  &  (~ ng2241) ) | ( pg35  &  (~ ng2153)  &  (~ ng2227) ) ;
 assign wire32720 = ( ng26703  &  wire32719 ) | ( ng17321  &  wire32719 ) ;
 assign wire32721 = ( pg35  &  ng2153  &  ng2241 ) | ( pg35  &  ng2227  &  ng2241 ) ;
 assign wire32722 = ( ng26703  &  wire32721 ) | ( ng17321  &  wire32721 ) ;
 assign wire32723 = ( ng2241  &  pg35 ) ;
 assign wire32724 = ( wire4343 ) | ( (~ ng26703)  &  (~ ng17321)  &  wire32723 ) ;
 assign wire32728 = ( pg35  &  ng2307  &  (~ ng2319)  &  (~ ng2351) ) ;
 assign wire32731 = ( pg35  &  (~ ng2342)  &  ng2319  &  ng2311 ) ;
 assign wire32733 = ( pg35  &  ng2342  &  (~ ng2319)  &  ng2295 ) ;
 assign wire32734 = ( (~ ng2342)  &  ng2351  &  ng2303 ) ;
 assign wire32735 = ( ng2370  &  pg35 ) ;
 assign wire32736 = ( ng2315  &  pg35 ) ;
 assign wire32740 = ( ng2299  &  (~ ng25349) ) | ( (~ ng25435)  &  wire32736 ) ;
 assign wire32741 = ( wire4332 ) | ( wire4333 ) | ( wire4334 ) | ( wire4339 ) ;
 assign wire32745 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng2748 ) ;
 assign wire32747 = ( ng2514  &  pg35 ) ;
 assign wire32749 = ( (~ ng2763)  &  pg35 ) ;
 assign wire32750 = ( ng2763  &  pg35 ) ;
 assign wire32751 = ( (~ pg35)  &  ng2759 ) | ( pg35  &  (~ ng2841) ) ;
 assign wire32753 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32754 = ( ng6645  &  pg35 ) ;
 assign wire32757 = ( pg35  &  ng3857  &  ng3863  &  (~ ng3869) ) ;
 assign wire32758 = ( ng2629  &  pg35 ) ;
 assign wire32760 = ( wire4309 ) | ( (~ ng26793)  &  (~ ng14506)  &  wire32758 ) ;
 assign wire32762 = ( pg35  &  (~ ng3639)  &  (~ ng23309) ) ;
 assign wire32764 = ( pg35  &  ng3639  &  ng23309 ) ;
 assign wire32766 = ( ng269  &  pg35 ) ;
 assign wire32767 = ( pg14147  &  pg35 ) ;
 assign wire32769 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32770 = ( ng3957  &  pg35 ) ;
 assign wire32775 = ( (~ pg35)  &  ng1171 ) | ( pg35  &  (~ pg7916)  &  ng1183 ) | ( pg35  &  (~ ng1171)  &  ng1183 ) | ( pg35  &  pg7916  &  ng1171  &  (~ ng1183) ) ;
 assign wire32777 = ( pg35  &  (~ ng4669)  &  (~ ng13330) ) ;
 assign wire32779 = ( pg35  &  ng4669  &  ng13330 ) ;
 assign wire32780 = ( wire4291 ) | ( ng31003  &  (~ ng10831)  &  wire32777 ) ;
 assign wire32781 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32782 = ( ng3602  &  pg35 ) ;
 assign wire32784 = ( ng3227  &  pg35 ) ;
 assign wire32785 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32787 = ( ng1996  &  pg35 ) ;
 assign wire32795 = ( (~ ng2036)  &  pg35 ) ;
 assign wire32798 = ( (~ pg35)  &  ng2791 ) | ( pg35  &  ng2795  &  (~ ng12377) ) ;
 assign wire32802 = ( (~ ng6049)  &  pg35 ) ;
 assign wire32804 = ( ng6049  &  pg35 ) ;
 assign wire32808 = ( (~ pg35)  &  ng4141 ) | ( pg35  &  (~ ng2841) ) ;
 assign wire32810 = ( pg35  &  pg12923  &  ng1252 ) ;
 assign wire32811 = ( (~ ng1252)  &  pg35 ) ;
 assign wire32817 = ( ng5224  &  pg35 ) ;
 assign wire32818 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32823 = ( pg35  &  (~ ng1668)  &  ng112 ) | ( pg35  &  ng1636  &  ng112 ) ;
 assign wire32825 = ( pg35  &  ng1668  &  (~ ng1636)  &  (~ ng112) ) ;
 assign wire32826 = ( ng1644  &  pg35 ) ;
 assign wire32830 = ( pg35  &  ng5170  &  (~ ng5176)  &  ng5164 ) ;
 assign wire32832 = ( ng1536  &  pg35 ) ;
 assign wire32834 = ( (~ pg35)  &  ng1532 ) | ( pg35  &  (~ ng1413)  &  ng1536 ) ;
 assign wire32836 = ( ng5228  &  pg35 ) ;
 assign wire32837 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32841 = ( (~ ng2331) ) | ( ng2361 ) ;
 assign wire32842 = ( pg35  &  ng17405  &  (~ wire32841) ) | ( pg35  &  ng26737  &  (~ wire32841) ) ;
 assign wire32843 = ( ng2303  &  pg35 ) ;
 assign wire32846 = ( (~ pg35)  &  ng336 ) | ( pg35  &  ng305 ) ;
 assign wire32851 = ( pg35  &  (~ ng5644)  &  (~ ng23909) ) ;
 assign wire32853 = ( pg35  &  ng5644  &  ng23909 ) ;
 assign wire32855 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32856 = ( ng3953  &  pg35 ) ;
 assign wire32858 = ( ng164  &  pg35 ) ;
 assign wire32860 = ( (~ ng164)  &  pg35 ) ;
 assign wire32861 = ( wire4204 ) | ( ng23042  &  (~ wire28708)  &  wire32858 ) ;
 assign wire32862 = ( pg35  &  wire7041 ) | ( pg35  &  ng14367  &  wire29097 ) ;
 assign wire32863 = ( ng1648  &  pg35 ) ;
 assign wire32865 = ( wire4200 ) | ( (~ ng27738)  &  wire32862 ) ;
 assign wire32866 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32867 = ( ng6295  &  pg35 ) ;
 assign wire32869 = ( ng1792  &  pg35 ) ;
 assign wire32870 = ( pg35  &  wire7257 ) | ( pg35  &  ng14367  &  wire28834 ) ;
 assign wire32871 = ( ng1783  &  pg35 ) ;
 assign wire32873 = ( wire4193 ) | ( (~ ng27775)  &  wire32870 ) ;
 assign wire32874 = ( pg35  &  ng26793  &  ng11978 ) | ( pg35  &  ng14506  &  ng11978 ) ;
 assign wire32875 = ( ng2583  &  pg35 ) ;
 assign wire32878 = ( pg35  &  wire28555  &  wire28556 ) ;
 assign wire32879 = ( (~ ng6395)  &  pg35 ) ;
 assign wire32881 = ( ng6395  &  pg35 ) ;
 assign wire32884 = ( pg35  &  (~ pg11678)  &  ng763 ) | ( pg35  &  ng763  &  ng736 ) ;
 assign wire32885 = ( (~ ng763)  &  pg35 ) ;
 assign wire32887 = ( ng1592  &  pg35 ) ;
 assign wire32891 = ( pg35  &  ng1632  &  ng25337 ) | ( pg35  &  (~ ng1636)  &  (~ ng25337) ) ;
 assign wire32893 = ( pg35  &  (~ pg11678)  &  ng744 ) | ( pg35  &  ng744  &  ng736 ) ;
 assign wire32894 = ( (~ ng744)  &  pg35 ) ;
 assign wire32898 = ( ng1448  &  pg35 ) ;
 assign wire32899 = ( ng1442  &  ng1454 ) | ( ng1454  &  ng1489 ) ;
 assign wire32902 = ( (~ ng1448)  &  pg35 ) ;
 assign wire32903 = ( ng1442  &  ng1454 ) | ( ng1454  &  ng1489 ) ;
 assign wire32907 = ( pg35  &  ng1448  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire32910 = ( pg35  &  (~ ng1448)  &  (~ ng1442)  &  (~ ng1489) ) ;
 assign wire32913 = ( (~ pg35)  &  ng1478 ) | ( pg35  &  ng1454  &  ng13273 ) ;
 assign wire32914 = ( (~ ng13378)  &  (~ ng13273)  &  wire32907 ) | ( ng13378  &  (~ ng13273)  &  wire32910 ) ;
 assign wire32917 = ( (~ ng2361)  &  pg35 ) ;
 assign wire32919 = ( ng17405  &  (~ ng28799)  &  wire32917 ) | ( ng26737  &  (~ ng28799)  &  wire32917 ) ;
 assign wire32921 = ( ng3566  &  pg35 ) ;
 assign wire32922 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32927 = ( pg35  &  ng3506  &  (~ ng3518)  &  ng3512 ) ;
 assign wire32928 = ( (~ ng3835)  &  pg35 ) ;
 assign wire32929 = ( ng3835  &  pg35 ) ;
 assign wire32933 = ( (~ ng2791)  &  pg35 ) ;
 assign wire32934 = ( (~ ng2724)  &  ng2729  &  (~ ng11405)  &  wire32933 ) ;
 assign wire32936 = ( (~ ng85)  &  (~ ng11405)  &  (~ wire28567) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire28567) ) ;
 assign wire32937 = ( ng2783  &  pg35 ) ;
 assign wire32938 = ( wire4137 ) | ( ng11405  &  wire32937 ) | ( wire28567  &  wire32937 ) ;
 assign wire32939 = ( wire32938 ) | ( (~ ng85)  &  wire32934 ) | ( (~ ng29503)  &  wire32934 ) ;
 assign wire32940 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire32941 = ( ng6243  &  pg35 ) ;
 assign wire32943 = ( ng239  &  pg35 ) ;
 assign wire32944 = ( pg14125  &  pg35 ) ;
 assign wire32948 = ( (~ ng2476) ) | ( ng2485 ) ;
 assign wire32949 = ( (~ ng2465)  &  pg35 ) ;
 assign wire32953 = ( pg35  &  ng2461  &  ng25476 ) | ( pg35  &  ng2421  &  (~ ng25476) ) ;
 assign wire32955 = ( pg35  &  (~ ng3288)  &  (~ ng23286) ) ;
 assign wire32957 = ( pg35  &  ng3288  &  ng23286 ) ;
 assign wire32961 = ( wire4115 ) | ( ng1263  &  ng22862  &  ng25895 ) ;
 assign wire32963 = ( pg35  &  ng4664  &  (~ ng11006) ) ;
 assign wire32965 = ( pg35  &  (~ ng4664)  &  ng11006 ) ;
 assign wire32966 = ( wire4112 ) | ( ng31003  &  (~ ng10831)  &  wire32963 ) ;
 assign wire32969 = ( pg35  &  (~ ng2070)  &  ng112 ) | ( pg35  &  ng112  &  ng2040 ) ;
 assign wire32971 = ( pg35  &  ng2070  &  (~ ng112)  &  (~ ng2040) ) ;
 assign wire32972 = ( ng2047  &  pg35 ) ;
 assign wire32975 = ( ng4434  &  ng4392 ) ;
 assign wire32976 = ( pg35  &  ng4443 ) | ( (~ pg35)  &  ng4434 ) ;
 assign wire32978 = ( pg35  &  (~ pg9048)  &  ng572 ) | ( pg35  &  ng559  &  ng572 ) ;
 assign wire32979 = ( (~ ng572)  &  pg35 ) ;
 assign wire32981 = ( (~ ng3990)  &  pg35 ) ;
 assign wire32983 = ( ng3990  &  pg35 ) ;
 assign wire32985 = ( wire4099 ) | ( (~ ng28484)  &  (~ ng23342)  &  wire32981 ) ;
 assign wire32987 = ( pg35  &  ng837  &  (~ ng812) ) ;
 assign wire32989 = ( pg35  &  ng837  &  ng812 ) ;
 assign wire32991 = ( ng3684  &  pg35 ) ;
 assign wire32992 = ( (~ ng3689)  &  pg16656 ) ;
 assign wire32993 = ( ng3703  &  (~ ng3639)  &  ng3554 ) ;
 assign wire32994 = ( ng3689  &  pg16924 ) ;
 assign wire32995 = ( ng3703  &  (~ ng3639)  &  ng3566 ) ;
 assign wire32997 = ( ng3703  &  (~ ng3639)  &  ng3542 ) ;
 assign wire32999 = ( pg16627  &  (~ ng3703)  &  (~ ng3639)  &  ng3602 ) ;
 assign wire33000 = ( ng3689  &  pg14451 ) ;
 assign wire33001 = ( (~ ng3703)  &  ng3538  &  (~ ng3639) ) ;
 assign wire33002 = ( ng3546  &  ng3689 ) ;
 assign wire33003 = ( (~ ng3703)  &  ng3680  &  (~ ng3639) ) ;
 assign wire33005 = ( pg13926  &  (~ ng3703)  &  ng3570  &  ng3639 ) ;
 assign wire33007 = ( pg16744  &  ng3586  &  ng3703  &  ng3639 ) ;
 assign wire33008 = ( (~ ng3689)  &  pg14451 ) ;
 assign wire33009 = ( (~ ng3703)  &  ng3639  &  ng3550 ) ;
 assign wire33010 = ( ng3689  &  pg16722 ) ;
 assign wire33011 = ( ng3703  &  ng3639  &  ng3598 ) ;
 assign wire33012 = ( ng3689  &  pg13881 ) ;
 assign wire33013 = ( (~ ng3703)  &  ng3639  &  ng3582 ) ;
 assign wire33014 = ( (~ ng3689)  &  pg16924 ) ;
 assign wire33015 = ( ng3574  &  ng3703  &  ng3639 ) ;
 assign wire33016 = ( wire32992  &  wire32993 ) | ( wire32994  &  wire32995 ) ;
 assign wire33017 = ( pg11388  &  ng3689  &  wire32997 ) | ( pg11388  &  ng3689  &  wire32999 ) | ( (~ pg11388)  &  (~ ng3689)  &  wire32999 ) ;
 assign wire33018 = ( wire33000  &  wire33001 ) | ( wire33002  &  wire33003 ) ;
 assign wire33019 = ( pg11388  &  ng3689  &  wire33005 ) | ( (~ pg11388)  &  (~ ng3689)  &  wire33005 ) | ( pg11388  &  ng3689  &  wire33007 ) | ( (~ pg11388)  &  (~ ng3689)  &  wire33007 ) ;
 assign wire33020 = ( wire33008  &  wire33009 ) | ( wire33010  &  wire33011 ) ;
 assign wire33021 = ( wire33012  &  wire33013 ) | ( wire33014  &  wire33015 ) ;
 assign wire33024 = ( wire33021 ) | ( wire33020 ) ;
 assign wire33025 = ( wire33016 ) | ( wire33017 ) | ( wire33018 ) | ( wire33019 ) ;
 assign wire33026 = ( ng3689  &  pg16656 ) ;
 assign wire33027 = ( ng3703  &  ng3639  &  ng3614 ) ;
 assign wire33029 = ( pg16744  &  ng3594  &  ng3703  &  (~ ng3639) ) ;
 assign wire33030 = ( (~ ng3689)  &  pg16722 ) ;
 assign wire33031 = ( ng3606  &  ng3703  &  (~ ng3639) ) ;
 assign wire33033 = ( pg13926  &  (~ ng3703)  &  ng3578  &  (~ ng3639) ) ;
 assign wire33034 = ( (~ ng3689)  &  pg13881 ) ;
 assign wire33035 = ( (~ ng3703)  &  (~ ng3639)  &  ng3590 ) ;
 assign wire33037 = ( pg16627  &  ng3610  &  (~ ng3703)  &  ng3639 ) ;
 assign wire33038 = ( (~ ng3689)  &  pg11388 ) ;
 assign wire33039 = ( ng3703  &  ng3639  &  ng3558 ) ;
 assign wire33040 = ( ng3562  &  (~ ng3689) ) ;
 assign wire33041 = ( (~ ng3703)  &  ng3680  &  ng3639 ) ;
 assign wire33042 = ( wire33026  &  wire33027 ) | ( ng11389  &  wire33029 ) ;
 assign wire33043 = ( wire33030  &  wire33031 ) | ( ng11389  &  wire33033 ) ;
 assign wire33044 = ( wire33034  &  wire33035 ) | ( ng11389  &  wire33037 ) ;
 assign wire33045 = ( wire33038  &  wire33039 ) | ( wire33040  &  wire33041 ) ;
 assign wire33048 = ( wire33042 ) | ( wire33043 ) | ( wire33044 ) | ( wire33045 ) ;
 assign wire33049 = ( pg35  &  wire6966 ) | ( pg35  &  wire6967 ) | ( pg35  &  wire29216 ) ;
 assign wire33054 = ( pg35  &  (~ pg9048)  &  ng586 ) | ( pg35  &  ng559  &  ng586 ) ;
 assign wire33055 = ( (~ ng586)  &  pg35 ) ;
 assign wire33061 = ( pg35  &  (~ ng2610)  &  (~ ng2619) ) | ( pg35  &  (~ ng2619)  &  ng2587 ) ;
 assign wire33062 = ( pg35  &  wire5887 ) | ( pg35  &  ng14367  &  wire31005 ) ;
 assign wire33063 = ( ng2587  &  pg35 ) ;
 assign wire33065 = ( wire4053 ) | ( (~ ng27933)  &  wire33062 ) ;
 assign wire33066 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33067 = ( ng6271  &  pg35 ) ;
 assign wire33069 = ( ng2020  &  pg35 ) ;
 assign wire33070 = ( pg35  &  ng26759  &  (~ wire32138) ) | ( pg35  &  ng14438  &  (~ wire32138) ) ;
 assign wire33072 = ( ng246  &  pg35 ) ;
 assign wire33073 = ( ng460  &  pg35 ) ;
 assign wire33075 = ( ng3247  &  pg35 ) ;
 assign wire33076 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33081 = ( (~ pg35)  &  ng5077 ) | ( pg35  &  (~ ng5073)  &  ng5077  &  (~ ng5084) ) ;
 assign wire33083 = ( (~ pg91)  &  pg35 ) | ( pg35  &  ng2965 ) | ( (~ pg35)  &  ng2955 ) ;
 assign wire33085 = ( pg35  &  (~ ng1322)  &  (~ ng1404) ) ;
 assign wire33087 = ( pg35  &  (~ ng1322)  &  ng1404 ) ;
 assign wire33088 = ( (~ pg35)  &  ng1395 ) | ( ng1395  &  (~ ng13134)  &  wire33085 ) ;
 assign wire33090 = ( pg35  &  (~ pg9048)  &  ng617 ) | ( pg35  &  ng559  &  ng617 ) ;
 assign wire33091 = ( (~ ng617)  &  pg35 ) ;
 assign wire33096 = ( pg35  &  (~ ng1834)  &  (~ ng1840) ) ;
 assign wire33098 = ( pg35  &  ng1834  &  ng1840 ) ;
 assign wire33099 = ( ng1844  &  pg35 ) ;
 assign wire33102 = ( ng1955  &  pg35 ) ;
 assign wire33104 = ( ng671  &  pg35 ) ;
 assign wire33105 = ( ng8806  &  wire33104 ) | ( (~ ng11185)  &  wire33104 ) | ( (~ wire30776)  &  wire33104 ) ;
 assign wire33106 = ( (~ ng671)  &  pg35 ) ;
 assign wire33107 = ( (~ ng8806)  &  ng11185  &  wire30776  &  wire33106 ) ;
 assign wire33109 = ( pg35  &  pg12923  &  ng1270 ) ;
 assign wire33111 = ( (~ pg35)  &  ng1263 ) | ( (~ ng1263)  &  wire33109 ) | ( ng25895  &  wire33109 ) ;
 assign wire33112 = ( ng5925  &  pg35 ) ;
 assign wire33113 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33115 = ( (~ ng2795)  &  pg35 ) ;
 assign wire33116 = ( ng2724  &  ng2729  &  (~ ng11405)  &  wire33115 ) ;
 assign wire33118 = ( (~ ng85)  &  (~ ng11405)  &  (~ wire29883) ) | ( (~ ng29503)  &  (~ ng11405)  &  (~ wire29883) ) ;
 assign wire33119 = ( ng2787  &  pg35 ) ;
 assign wire33120 = ( wire3998 ) | ( ng11405  &  wire33119 ) | ( wire29883  &  wire33119 ) ;
 assign wire33121 = ( wire33120 ) | ( (~ ng85)  &  wire33116 ) | ( (~ ng29503)  &  wire33116 ) ;
 assign wire33122 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33123 = ( ng6601  &  pg35 ) ;
 assign wire33124 = ( wire3994 ) | ( ng12716  &  ng12680  &  wire33122 ) ;
 assign wire33126 = ( ng4141 ) | ( ng4064 ) | ( (~ ng4057) ) | ( ng4082 ) ;
 assign wire33127 = ( ng4145  &  pg35 ) ;
 assign wire33128 = ( ng4119  &  pg35 ) ;
 assign wire33129 = ( wire3991 ) | ( ng13806  &  (~ wire33126)  &  wire33127 ) ;
 assign wire33131 = ( pg35  &  (~ ng5835)  &  (~ ng5841) ) ;
 assign wire33133 = ( pg35  &  ng5835  &  ng5841 ) ;
 assign wire33136 = ( ng10869  &  wire33133 ) | ( pg35  &  ng5845  &  (~ ng10869) ) ;
 assign wire33137 = ( ng3550  &  pg35 ) ;
 assign wire33138 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33139 = ( wire3984 ) | ( (~ ng11483)  &  wire33137 ) | ( (~ ng11571)  &  wire33137 ) ;
 assign wire33140 = ( ng1687  &  pg35 ) ;
 assign wire33143 = ( pg35  &  (~ ng1700)  &  (~ ng1706) ) ;
 assign wire33145 = ( pg35  &  ng1700  &  ng1706 ) ;
 assign wire33146 = ( ng1710  &  pg35 ) ;
 assign wire33150 = ( pg35  &  (~ ng5142)  &  (~ ng5148) ) ;
 assign wire33152 = ( pg35  &  ng5142  &  ng5148 ) ;
 assign wire33155 = ( ng10823  &  wire33152 ) | ( pg35  &  ng5152  &  (~ ng10823) ) ;
 assign wire33156 = ( ng2060  &  pg35 ) ;
 assign wire33157 = ( pg35  &  wire6319 ) | ( pg35  &  ng14367  &  wire30342 ) ;
 assign wire33158 = ( ng2051  &  pg35 ) ;
 assign wire33160 = ( wire3969 ) | ( (~ ng27882)  &  wire33157 ) ;
 assign wire33161 = ( ng5046  &  pg35 ) ;
 assign wire33165 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33166 = ( ng3614  &  pg35 ) ;
 assign wire33168 = ( ng5272  &  pg35 ) ;
 assign wire33169 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33172 = ( pg35  &  ng4349  &  (~ ng4358)  &  (~ ng12925) ) ;
 assign wire33174 = ( pg35  &  (~ ng4349)  &  ng4358 ) | ( pg35  &  ng4358  &  ng12925 ) ;
 assign wire33176 = ( ng5260  &  pg35 ) ;
 assign wire33177 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33180 = ( pg35  &  ng17405  &  ng9700 ) | ( pg35  &  ng26737  &  ng9700 ) ;
 assign wire33181 = ( ng2299  &  pg35 ) ;
 assign wire33183 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33184 = ( ng3905  &  pg35 ) ;
 assign wire33189 = ( pg35  &  (~ pg17577)  &  (~ pg17674)  &  (~ pg14662) ) ;
 assign wire33194 = ( pg35  &  (~ pg17577)  &  pg17674  &  pg14662 ) ;
 assign wire33199 = ( pg35  &  pg17577  &  pg17674  &  pg14662 ) ;
 assign wire33200 = ( (~ pg17674)  &  pg17519  &  pg12238 ) | ( (~ pg14662)  &  pg17519  &  pg12238 ) ;
 assign wire33204 = ( pg35  &  (~ pg17577)  &  pg14662  &  (~ pg17519) ) ;
 assign wire33208 = ( ng1917  &  pg35 ) ;
 assign wire33209 = ( pg35  &  wire6655 ) | ( pg35  &  ng14367  &  wire29571 ) ;
 assign wire33211 = ( wire3924 ) | ( (~ ng27833)  &  wire33209 ) ;
 assign wire33212 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33213 = ( ng5965  &  pg35 ) ;
 assign wire33215 = ( ng5933  &  pg35 ) ;
 assign wire33216 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33218 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33219 = ( ng5611  &  pg35 ) ;
 assign wire33222 = ( ng4555  &  ng4561 ) ;
 assign wire33223 = ( (~ pg73)  &  (~ pg72)  &  ng4558  &  ng4564 ) ;
 assign wire33225 = ( pg73  &  pg35 ) | ( pg72  &  pg35 ) ;
 assign wire33227 = ( wire3910 ) | ( wire3912 ) | ( wire33222  &  wire33223 ) ;
 assign wire33230 = ( pg35  &  ng26673  &  ng9586 ) | ( pg35  &  ng9586  &  ng17292 ) ;
 assign wire33231 = ( ng1604  &  pg35 ) ;
 assign wire33233 = ( pg35  &  ng26759  &  ng9755 ) | ( pg35  &  ng14438  &  ng9755 ) ;
 assign wire33234 = ( ng2008  &  pg35 ) ;
 assign wire33238 = ( ng2433  &  pg35 ) ;
 assign wire33239 = ( pg35  &  ng26770  &  ng9762 ) | ( pg35  &  ng17424  &  ng9762 ) ;
 assign wire33241 = ( ng6637  &  pg35 ) ;
 assign wire33242 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33244 = ( ng3558  &  pg35 ) ;
 assign wire33245 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33246 = ( wire3889 ) | ( (~ ng11527)  &  wire33244 ) | ( (~ ng11571)  &  wire33244 ) ;
 assign wire33248 = ( pg35  &  ng157  &  ng23042 ) ;
 assign wire33249 = ( (~ ng157)  &  pg35 ) ;
 assign wire33250 = ( wire3886 ) | ( (~ ng28353)  &  wire33248 ) | ( wire28711  &  wire33248 ) ;
 assign wire33251 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33252 = ( ng5961  &  pg35 ) ;
 assign wire33254 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33255 = ( ng6629  &  pg35 ) ;
 assign wire33257 = ( (~ ng1216)  &  pg35 ) ;
 assign wire33259 = ( ng1216  &  pg35 ) ;
 assign wire33261 = ( wire3874 ) | ( (~ ng11130)  &  (~ ng11148)  &  wire33257 ) ;
 assign wire33262 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33263 = ( ng5208  &  pg35 ) ;
 assign wire33264 = ( wire3868 ) | ( ng12405  &  ng12492  &  wire33262 ) ;
 assign wire33265 = ( pg35  &  (~ ng1816) ) | ( pg35  &  (~ ng1728)  &  (~ ng1802) ) ;
 assign wire33266 = ( ng17317  &  wire33265 ) | ( ng26694  &  wire33265 ) ;
 assign wire33267 = ( pg35  &  ng1728  &  ng1816 ) | ( pg35  &  ng1816  &  ng1802 ) ;
 assign wire33268 = ( ng17317  &  wire33267 ) | ( ng26694  &  wire33267 ) ;
 assign wire33269 = ( ng1816  &  pg35 ) ;
 assign wire33270 = ( wire3860 ) | ( (~ ng17317)  &  (~ ng26694)  &  wire33269 ) ;
 assign wire33273 = ( pg35  &  (~ ng2399)  &  (~ ng2393) ) ;
 assign wire33275 = ( pg35  &  ng2399  &  ng2393 ) ;
 assign wire33276 = ( ng2403  &  pg35 ) ;
 assign wire33280 = ( ng29503  &  wire6172 ) | ( ng29503  &  ng14367  &  wire30555 ) ;
 assign wire33282 = ( pg35  &  ng110  &  (~ ng2217) ) | ( pg35  &  ng110  &  ng2208 ) ;
 assign wire33284 = ( pg35  &  (~ ng110)  &  ng2217  &  (~ ng2208) ) ;
 assign wire33285 = ( ng2223  &  pg35 ) ;
 assign wire33286 = ( wire3849 ) | ( ng26171  &  wire33280  &  wire33282 ) ;
 assign wire33287 = ( (~ ng26171)  &  wire33285 ) | ( (~ wire33280)  &  wire33285 ) | ( ng26171  &  wire33280  &  wire33284 ) ;
 assign wire33288 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33289 = ( ng5957  &  pg35 ) ;
 assign wire33291 = ( (~ ng832)  &  pg35 ) ;
 assign wire33293 = ( ng832  &  pg35 ) ;
 assign wire33296 = ( (~ ng2461)  &  pg35 ) ;
 assign wire33299 = ( (~ pg35)  &  ng2811 ) | ( pg35  &  ng2823  &  (~ ng12377) ) ;
 assign wire33302 = ( pg35  &  (~ ng1783)  &  (~ ng1792) ) | ( pg35  &  (~ ng1792)  &  ng1760 ) ;
 assign wire33303 = ( ng1760  &  pg35 ) ;
 assign wire33304 = ( pg35  &  wire7257 ) | ( pg35  &  ng14367  &  wire28834 ) ;
 assign wire33306 = ( wire3829 ) | ( (~ ng27775)  &  wire33304 ) ;
 assign wire33307 = ( (~ ng2208) ) | ( ng2217 ) ;
 assign wire33308 = ( ng2193  &  pg35 ) ;
 assign wire33312 = ( pg35  &  (~ ng2197)  &  (~ ng25396) ) | ( pg35  &  ng2153  &  (~ ng25396) ) ;
 assign wire33316 = ( (~ pg35)  &  ng4477 ) | ( pg35  &  ng4581  &  ng59 ) ;
 assign wire33317 = ( (~ pg73)  &  pg35  &  ng4581 ) | ( (~ pg72)  &  pg35  &  ng4581 ) ;
 assign wire33319 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33320 = ( ng3582  &  pg35 ) ;
 assign wire33325 = ( pg35  &  (~ ng4608)  &  (~ ng30583)  &  (~ wire6408) ) ;
 assign wire33327 = ( pg35  &  ng4608  &  (~ ng30583)  &  (~ wire6408) ) ;
 assign wire33330 = ( pg35  &  (~ ng1926)  &  (~ ng1917) ) | ( pg35  &  (~ ng1926)  &  ng1894 ) ;
 assign wire33331 = ( ng1894  &  pg35 ) ;
 assign wire33332 = ( pg35  &  wire6655 ) | ( pg35  &  ng14367  &  wire29571 ) ;
 assign wire33334 = ( wire3805 ) | ( (~ ng27833)  &  wire33332 ) ;
 assign wire33335 = ( ng5011  &  pg35 ) ;
 assign wire33336 = ( pg35  &  wire7046 ) | ( pg35  &  wire7047 ) | ( pg35  &  wire29091 ) ;
 assign wire33343 = ( (~ pg35)  &  ng6494 ) | ( pg35  &  (~ pg9817)  &  pg9743  &  (~ ng6494) ) ;
 assign wire33344 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33345 = ( ng5220  &  pg35 ) ;
 assign wire33349 = ( ng2370  &  (~ ng2384) ) | ( ng2342  &  (~ ng2319)  &  ng2370 ) ;
 assign wire33350 = ( ng2384  &  pg35 ) ;
 assign wire33351 = ( (~ pg35)  &  ng2370 ) | ( pg35  &  (~ ng2370)  &  ng22432  &  ng14679 ) ;
 assign wire33353 = ( (~ ng4521)  &  pg35 ) ;
 assign wire33354 = ( (~ pg35)  &  ng4521 ) | ( (~ ng4527)  &  ng4521  &  ng12228 ) | ( ng4527  &  ng4521  &  (~ ng12228) ) ;
 assign wire33355 = ( ng1489  &  pg35 ) ;
 assign wire33357 = ( (~ ng1442)  &  pg35 ) ;
 assign wire33362 = ( ng2265  &  pg35 ) ;
 assign wire33364 = ( ng1974  &  pg35 ) ;
 assign wire33366 = ( pg35  &  (~ ng1146)  &  (~ ng1099) ) ;
 assign wire33370 = ( (~ pg35)  &  ng1105 ) | ( pg35  &  ng1124  &  ng13307 ) ;
 assign wire33372 = ( ng2465 ) | ( (~ ng2421) ) ;
 assign wire33373 = ( pg35  &  ng26770  &  (~ wire33372) ) | ( pg35  &  ng17424  &  (~ wire33372) ) ;
 assign wire33374 = ( ng2429  &  pg35 ) ;
 assign wire33377 = ( pg35  &  (~ ng1974)  &  (~ ng1968) ) ;
 assign wire33378 = ( ng1968  &  ng1974 ) ;
 assign wire33379 = ( ng1978  &  pg35 ) ;
 assign wire33382 = ( ng3199  &  pg35 ) ;
 assign wire33383 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33384 = ( wire3752 ) | ( (~ ng11514)  &  wire33382 ) | ( (~ ng11435)  &  wire33382 ) ;
 assign wire33385 = ( pg35  &  ng17317  &  ng9640 ) | ( pg35  &  ng26694  &  ng9640 ) ;
 assign wire33386 = ( ng1740  &  pg35 ) ;
 assign wire33392 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33393 = ( ng6617  &  pg35 ) ;
 assign wire33397 = ( (~ ng2250)  &  ng2236 ) | ( (~ ng2185)  &  ng2236  &  ng2208 ) ;
 assign wire33398 = ( ng2250  &  pg35 ) ;
 assign wire33399 = ( (~ pg35)  &  ng2236 ) | ( pg35  &  (~ ng2236)  &  ng22384  &  ng14642 ) ;
 assign wire33401 = ( ng29503  &  wire7030 ) | ( ng29503  &  ng14367  &  wire29111 ) ;
 assign wire33403 = ( pg35  &  ng110  &  ng2342 ) | ( pg35  &  ng110  &  (~ ng2351) ) ;
 assign wire33405 = ( pg35  &  (~ ng110)  &  (~ ng2342)  &  ng2351 ) ;
 assign wire33406 = ( ng2357  &  pg35 ) ;
 assign wire33407 = ( wire3727 ) | ( ng26195  &  wire33401  &  wire33403 ) ;
 assign wire33408 = ( (~ ng26195)  &  wire33406 ) | ( (~ wire33401)  &  wire33406 ) | ( ng26195  &  wire33401  &  wire33405 ) ;
 assign wire33410 = ( pg35  &  (~ ng5115)  &  ng20682 ) | ( pg35  &  ng20682  &  ng11111 ) ;
 assign wire33412 = ( pg35  &  ng5115  &  ng20682  &  (~ ng11111) ) ;
 assign wire33413 = ( ng5115  &  pg35 ) ;
 assign wire33416 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33417 = ( ng5595  &  pg35 ) ;
 assign wire33421 = ( pg35  &  (~ ng2841) ) | ( (~ pg35)  &  ng2729 ) ;
 assign wire33424 = ( pg35  &  ng4653  &  ng4688  &  (~ ng4659) ) ;
 assign wire33426 = ( pg35  &  (~ ng4653)  &  ng4659 ) | ( pg35  &  (~ ng4688)  &  ng4659 ) ;
 assign wire33427 = ( wire3712 ) | ( ng31003  &  (~ ng10831)  &  wire33424 ) ;
 assign wire33428 = ( ng1135  &  pg35 ) ;
 assign wire33429 = ( ng1146  &  ng1094 ) | ( ng1094  &  ng1099 ) ;
 assign wire33432 = ( (~ ng1135)  &  pg35 ) ;
 assign wire33433 = ( ng1146  &  ng1094 ) | ( ng1094  &  ng1099 ) ;
 assign wire33437 = ( pg35  &  ng1135  &  (~ ng1146)  &  (~ ng1099) ) ;
 assign wire33440 = ( pg35  &  (~ ng1135)  &  (~ ng1146)  &  (~ ng1099) ) ;
 assign wire33443 = ( (~ pg35)  &  ng1099 ) | ( pg35  &  ng1094  &  ng13846 ) ;
 assign wire33444 = ( (~ ng13336)  &  (~ ng13846)  &  wire33437 ) | ( ng13336  &  (~ ng13846)  &  wire33440 ) ;
 assign wire33450 = ( (~ pg35)  &  ng1526 ) | ( pg35  &  (~ pg7946)  &  ng1521 ) ;
 assign wire33452 = ( pg35  &  (~ pg11678)  &  ng772 ) | ( pg35  &  ng736  &  ng772 ) ;
 assign wire33453 = ( (~ ng772)  &  pg35 ) ;
 assign wire33455 = ( (~ ng2555) ) | ( ng2599 ) ;
 assign wire33456 = ( pg35  &  ng26793  &  (~ wire33455) ) | ( pg35  &  ng14506  &  (~ wire33455) ) ;
 assign wire33457 = ( ng2563  &  pg35 ) ;
 assign wire33459 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33460 = ( ng3598  &  pg35 ) ;
 assign wire33463 = ( pg35  &  ng294  &  ng23204 ) ;
 assign wire33464 = ( (~ ng294)  &  pg35 ) ;
 assign wire33472 = ( pg35  &  (~ ng1379)  &  (~ ng15748) ) ;
 assign wire33473 = ( ng1379  &  pg35 ) ;
 assign wire33475 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33476 = ( ng5587  &  pg35 ) ;
 assign wire33480 = ( pg13272 ) | ( pg19357 ) | ( ng1333 ) ;
 assign wire33485 = ( ng6291  &  pg35 ) ;
 assign wire33486 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33489 = ( pg35  &  ng2946 ) | ( (~ pg35)  &  ng2941 ) | ( pg35  &  ng2955 ) ;
 assign wire33492 = ( wire33489 ) | ( pg35  &  ng28220 ) | ( pg35  &  ng22585 ) ;
 assign wire33494 = ( pg35  &  (~ ng3106)  &  ng3111 ) ;
 assign wire33495 = ( (~ ng3111)  &  ng3106 ) ;
 assign wire33497 = ( (~ ng23067)  &  wire33495 ) | ( pg35  &  ng3115  &  ng23067 ) ;
 assign wire33499 = ( pg35  &  (~ ng1720)  &  (~ ng1714) ) ;
 assign wire33501 = ( ng1724  &  pg35 ) ;
 assign wire33503 = ( ng25275  &  wire33501 ) | ( ng1720  &  ng1714  &  (~ ng25275) ) ;
 assign wire33505 = ( pg35  &  (~ ng6173)  &  (~ ng6167) ) ;
 assign wire33507 = ( ng6167  &  ng6173 ) ;
 assign wire33509 = ( (~ ng23699)  &  wire33507 ) | ( pg35  &  ng6177  &  ng23699 ) ;
 assign wire33510 = ( (~ ng4593)  &  pg35 ) ;
 assign wire33512 = ( ng4593  &  pg35 ) ;
 assign wire33515 = ( ng1024  &  pg35 ) ;
 assign wire33517 = ( wire3642 ) | ( ng25911  &  wire33515 ) | ( wire7652  &  wire33515 ) ;
 assign wire33519 = ( pg35  &  ng5057  &  (~ wire29550)  &  (~ wire29551) ) ;
 assign wire33520 = ( (~ ng5057)  &  pg35 ) ;
 assign wire33522 = ( (~ ng4776)  &  pg35 ) ;
 assign wire33523 = ( ng4801  &  ng4793  &  ng10831  &  wire33522 ) ;
 assign wire33524 = ( ng4776  &  pg35 ) ;
 assign wire33525 = ( (~ ng4801)  &  wire33524 ) | ( (~ ng4793)  &  wire33524 ) | ( (~ ng10831)  &  wire33524 ) ;
 assign wire33526 = ( wire3632 ) | ( ng28336  &  ng13464  &  wire33523 ) ;
 assign wire33527 = ( ng5591  &  pg35 ) ;
 assign wire33528 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33533 = ( pg35  &  (~ pg11678)  &  ng807 ) | ( pg35  &  ng736  &  ng807 ) ;
 assign wire33534 = ( (~ ng807)  &  pg35 ) ;
 assign wire33536 = ( (~ ng1592) ) | ( ng1636 ) ;
 assign wire33537 = ( pg35  &  ng26673  &  (~ wire33536) ) | ( pg35  &  ng17292  &  (~ wire33536) ) ;
 assign wire33538 = ( ng1600  &  pg35 ) ;
 assign wire33544 = ( pg35  &  ng26759  &  ng11956 ) | ( pg35  &  ng14438  &  ng11956 ) ;
 assign wire33545 = ( ng2024  &  pg35 ) ;
 assign wire33551 = ( (~ pg8919)  &  (~ pg8918)  &  (~ pg11770)  &  (~ pg8920) ) ;
 assign wire33552 = ( (~ pg8915)  &  (~ pg8917)  &  (~ pg8916)  &  (~ ng4235) ) ;
 assign wire33553 = ( (~ pg8870)  &  ng4235 ) | ( pg8870  &  (~ ng4235) ) ;
 assign wire33554 = ( pg35  &  (~ ng4145)  &  (~ ng4253) ) | ( pg35  &  ng4253  &  (~ ng4164) ) ;
 assign wire33555 = ( pg35  &  ng4145  &  (~ ng4253) ) | ( pg35  &  ng4145  &  ng4164 ) | ( pg35  &  ng4253  &  ng4164 ) ;
 assign wire33558 = ( pg35  &  ng2841  &  (~ ng2741) ) ;
 assign wire33560 = ( pg35  &  ng2841  &  ng2741 ) ;
 assign wire33561 = ( (~ pg35)  &  ng2735 ) | ( ng2735  &  (~ ng17297)  &  wire33558 ) ;
 assign wire33562 = ( pg35  &  wire6172 ) | ( pg35  &  ng14367  &  wire30555 ) ;
 assign wire33563 = ( ng2217  &  pg35 ) ;
 assign wire33564 = ( ng2208  &  pg35 ) ;
 assign wire33566 = ( wire3595 ) | ( (~ ng27796)  &  wire33562 ) ;
 assign wire33571 = ( (~ ng1714)  &  pg35 ) ;
 assign wire33572 = ( ng1714  &  pg35 ) ;
 assign wire33579 = ( (~ pg14421)  &  pg11349 ) ;
 assign wire33580 = ( pg35  &  (~ pg16624)  &  (~ pg16603)  &  pg13895 ) ;
 assign wire33585 = ( pg35  &  (~ pg16718)  &  (~ pg16624)  &  (~ pg16603) ) ;
 assign wire33590 = ( pg35  &  (~ pg9048)  &  ng595 ) | ( pg35  &  ng559  &  ng595 ) ;
 assign wire33591 = ( (~ ng595)  &  pg35 ) ;
 assign wire33592 = ( wire3574 ) | ( (~ ng27629)  &  wire33590 ) | ( wire28803  &  wire33590 ) ;
 assign wire33593 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33594 = ( ng3542  &  pg35 ) ;
 assign wire33595 = ( wire3571 ) | ( ng11747  &  ng11571  &  wire33593 ) ;
 assign wire33600 = ( pg12350  &  (~ pg17646) ) ;
 assign wire33601 = ( pg35  &  (~ pg13068)  &  pg14738  &  (~ pg17607) ) ;
 assign wire33606 = ( pg35  &  (~ pg13068)  &  (~ pg14738)  &  (~ pg17607) ) ;
 assign wire33608 = ( (~ ng1728) ) | ( ng1772 ) ;
 assign wire33609 = ( pg35  &  ng17317  &  (~ wire33608) ) | ( pg35  &  ng26694  &  (~ wire33608) ) ;
 assign wire33610 = ( ng1736  &  pg35 ) ;
 assign wire33613 = ( pg35  &  ng2380  &  (~ ng2384) ) ;
 assign wire33615 = ( ng2389  &  pg35 ) ;
 assign wire33617 = ( ng25473  &  wire33615 ) | ( (~ ng2380)  &  ng2384  &  (~ ng25473) ) ;
 assign wire33620 = ( pg35  &  ng2575  &  (~ ng2619)  &  (~ ng2587) ) ;
 assign wire33623 = ( pg35  &  (~ ng2610)  &  ng2579  &  ng2587 ) ;
 assign wire33625 = ( pg35  &  ng2610  &  (~ ng2587)  &  ng2563 ) ;
 assign wire33626 = ( (~ ng2610)  &  ng2571  &  ng2619 ) ;
 assign wire33627 = ( ng2583  &  pg35 ) ;
 assign wire33628 = ( ng2638  &  pg35 ) ;
 assign wire33632 = ( ng2567  &  (~ ng25439) ) | ( (~ ng25498)  &  wire33627 ) ;
 assign wire33633 = ( wire3546 ) | ( wire3547 ) | ( wire3548 ) | ( wire3553 ) ;
 assign wire33635 = ( ng29503  &  wire6319 ) | ( ng29503  &  ng14367  &  wire30342 ) ;
 assign wire33637 = ( pg35  &  ng110  &  ng2051 ) | ( pg35  &  ng110  &  (~ ng2060) ) ;
 assign wire33639 = ( pg35  &  (~ ng110)  &  (~ ng2051)  &  ng2060 ) ;
 assign wire33640 = ( ng2066  &  pg35 ) ;
 assign wire33641 = ( wire3545 ) | ( ng26213  &  wire33635  &  wire33637 ) ;
 assign wire33642 = ( (~ ng26213)  &  wire33640 ) | ( (~ wire33635)  &  wire33640 ) | ( ng26213  &  wire33635  &  wire33639 ) ;
 assign wire33643 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33644 = ( ng5232  &  pg35 ) ;
 assign wire33648 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33649 = ( ng5547  &  pg35 ) ;
 assign wire33650 = ( wire3533 ) | ( ng12798  &  ng12558  &  wire33648 ) ;
 assign wire33651 = ( ng4141 ) | ( (~ ng4064) ) | ( (~ ng4057) ) | ( ng4082 ) ;
 assign wire33652 = ( ng4122  &  pg35 ) ;
 assign wire33653 = ( ng4145  &  pg35 ) ;
 assign wire33654 = ( wire3530 ) | ( (~ ng13806)  &  wire33652 ) | ( wire33651  &  wire33652 ) ;
 assign wire33656 = ( pg35  &  (~ pg19357) ) | ( (~ pg35)  &  ng1404 ) ;
 assign wire33657 = ( pg35  &  pg12923  &  ng1404 ) | ( pg35  &  (~ pg12923)  &  (~ ng1404) ) ;
 assign wire33659 = ( (~ ng1592) ) | ( (~ ng1668) ) ;
 assign wire33660 = ( pg35  &  ng26673  &  (~ wire33659) ) | ( pg35  &  ng17292  &  (~ wire33659) ) ;
 assign wire33661 = ( ng1612  &  pg35 ) ;
 assign wire33665 = ( (~ ng490)  &  pg35 ) ;
 assign wire33666 = ( ng490  &  pg35 ) ;
 assign wire33667 = ( (~ pg35)  &  ng482 ) | ( pg35  &  ng667  &  (~ ng686) ) ;
 assign wire33668 = ( wire33667 ) | ( ng482  &  ng20000  &  wire33665 ) ;
 assign wire33670 = ( pg35  &  (~ ng3457)  &  ng21024 ) | ( pg35  &  ng21024  &  ng10733 ) ;
 assign wire33672 = ( pg35  &  ng3457  &  ng21024  &  (~ ng10733) ) ;
 assign wire33673 = ( ng3457  &  pg35 ) ;
 assign wire33676 = ( (~ ng4709)  &  pg35 ) ;
 assign wire33678 = ( ng4709  &  pg35 ) ;
 assign wire33680 = ( wire3501 ) | ( ng28336  &  (~ ng16173)  &  wire33676 ) ;
 assign wire33681 = ( pg35  &  ng26770  &  ng11960 ) | ( pg35  &  ng17424  &  ng11960 ) ;
 assign wire33682 = ( ng2449  &  pg35 ) ;
 assign wire33684 = ( ng5212  &  pg35 ) ;
 assign wire33685 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33688 = ( pg35  &  ng1821  &  (~ ng1825) ) ;
 assign wire33690 = ( pg35  &  (~ ng1821)  &  ng1825 ) ;
 assign wire33693 = ( (~ ng25426)  &  wire33690 ) | ( pg35  &  ng1830  &  ng25426 ) ;
 assign wire33694 = ( pg35  &  ng4375  &  (~ ng4382) ) ;
 assign wire33695 = ( (~ ng4392)  &  pg35 ) ;
 assign wire33696 = ( wire3485 ) | ( (~ wire29325)  &  wire33694 ) | ( (~ wire29326)  &  wire33694 ) ;
 assign wire33699 = ( pg35  &  (~ pg12919)  &  (~ ng1061) ) | ( pg35  &  pg12919  &  ng1052 ) ;
 assign wire33700 = ( pg35  &  (~ pg19334) ) | ( (~ pg35)  &  ng1061 ) | ( pg35  &  pg12919  &  ng1061 ) ;
 assign wire33703 = ( pg35  &  ng2173  &  (~ ng2185)  &  (~ ng2217) ) ;
 assign wire33706 = ( pg35  &  ng2177  &  ng2185  &  (~ ng2208) ) ;
 assign wire33708 = ( pg35  &  ng2161  &  (~ ng2185)  &  ng2208 ) ;
 assign wire33709 = ( ng2217  &  (~ ng2208)  &  ng2169 ) ;
 assign wire33710 = ( ng2181  &  pg35 ) ;
 assign wire33711 = ( ng2236  &  pg35 ) ;
 assign wire33715 = ( ng2165  &  (~ ng25309) ) | ( (~ ng25396)  &  wire33710 ) ;
 assign wire33716 = ( wire3465 ) | ( wire3466 ) | ( wire3467 ) | ( wire3471 ) ;
 assign wire33720 = ( (~ pg13049)  &  pg12300 ) ;
 assign wire33721 = ( pg35  &  pg14694  &  (~ pg17580)  &  (~ pg17604) ) ;
 assign wire33726 = ( pg35  &  (~ pg14694)  &  (~ pg17580)  &  (~ pg17711) ) ;
 assign wire33728 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33729 = ( ng6287  &  pg35 ) ;
 assign wire33735 = ( (~ ng918)  &  pg35 ) ;
 assign wire33736 = ( pg35  &  pg12919  &  ng918 ) ;
 assign wire33738 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33739 = ( ng5945  &  pg35 ) ;
 assign wire33743 = ( ng2246  &  pg35 ) ;
 assign wire33745 = ( ng29503  &  ng25357  &  wire28614 ) ;
 assign wire33747 = ( pg35  &  ng110  &  (~ ng1926) ) | ( pg35  &  ng110  &  ng1917 ) ;
 assign wire33749 = ( pg35  &  (~ ng110)  &  ng1926  &  (~ ng1917) ) ;
 assign wire33750 = ( ng1932  &  pg35 ) ;
 assign wire33751 = ( wire3442 ) | ( ng22417  &  wire33745  &  wire33747 ) ;
 assign wire33752 = ( (~ ng22417)  &  wire33750 ) | ( (~ wire33745)  &  wire33750 ) | ( ng22417  &  wire33745  &  wire33749 ) ;
 assign wire33754 = ( (~ pg35)  &  ng1589 ) | ( pg35  &  (~ pg17423)  &  pg10527 ) ;
 assign wire33755 = ( ng3941  &  pg35 ) ;
 assign wire33756 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33758 = ( ng1802 ) | ( (~ ng1772) ) ;
 assign wire33759 = ( pg35  &  ng17317  &  (~ wire33758) ) | ( pg35  &  ng26694  &  (~ wire33758) ) ;
 assign wire33760 = ( ng1744  &  pg35 ) ;
 assign wire33765 = ( pg35  &  ng2652  &  (~ ng2648) ) ;
 assign wire33767 = ( pg35  &  (~ ng2652)  &  ng2648 ) ;
 assign wire33770 = ( (~ ng25514)  &  wire33767 ) | ( pg35  &  ng2657  &  ng25514 ) ;
 assign wire33771 = ( wire1421  &  ng4939 ) | ( ng4939  &  ng4818 ) | ( ng4939  &  (~ ng24374) ) ;
 assign wire33773 = ( pg35  &  ng71  &  ng24374  &  (~ wire28575) ) ;
 assign wire33775 = ( ng29702  &  wire33773 ) | ( pg35  &  ng4933  &  (~ ng29702) ) ;
 assign wire33777 = ( pg35  &  (~ pg9048)  &  ng608 ) | ( pg35  &  ng559  &  ng608 ) ;
 assign wire33778 = ( (~ ng608)  &  pg35 ) ;
 assign wire33779 = ( wire3418 ) | ( ng31509  &  wire33777 ) | ( (~ wire30328)  &  wire33777 ) ;
 assign wire33780 = ( pg35  &  ng26725  &  (~ wire30477) ) | ( pg35  &  ng17401  &  (~ wire30477) ) ;
 assign wire33781 = ( ng1886  &  pg35 ) ;
 assign wire33784 = ( pg35  &  (~ ng1030)  &  ng1008 ) | ( pg35  &  (~ ng1018)  &  ng1008 ) ;
 assign wire33786 = ( pg35  &  (~ ng1030)  &  ng1008 ) | ( pg35  &  (~ ng1018)  &  ng1008 ) ;
 assign wire33789 = ( wire3407 ) | ( wire3409 ) | ( (~ ng7598)  &  wire33784 ) ;
 assign wire33794 = ( pg35  &  (~ ng703)  &  ng854 ) ;
 assign wire33795 = ( ng392  &  pg35 ) ;
 assign wire33798 = ( pg35  &  (~ ng146)  &  (~ ng13756) ) ;
 assign wire33800 = ( pg35  &  ng146  &  ng13756 ) ;
 assign wire33803 = ( pg35  &  (~ ng2661)  &  (~ ng2667) ) ;
 assign wire33804 = ( ng2667  &  ng2661 ) ;
 assign wire33805 = ( ng2671  &  pg35 ) ;
 assign wire33812 = ( ng5909  &  pg35 ) ;
 assign wire33813 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33814 = ( wire3389 ) | ( (~ ng12609)  &  wire33812 ) | ( (~ ng12571)  &  wire33812 ) ;
 assign wire33817 = ( (~ ng4349)  &  (~ ng4322)  &  (~ ng4358) ) ;
 assign wire33818 = ( pg90  &  pg35  &  (~ ng4332)  &  (~ ng2994) ) ;
 assign wire33820 = ( pg73  &  (~ ng4322) ) | ( pg72  &  (~ ng4322) ) ;
 assign wire33821 = ( pg35  &  (~ ng4332)  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire33823 = ( pg73  &  ng4322 ) | ( pg72  &  ng4322 ) ;
 assign wire33824 = ( pg35  &  (~ ng4332)  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire33826 = ( ng4311  &  (~ ng4322) ) ;
 assign wire33827 = ( pg35  &  ng4332  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire33830 = ( pg35  &  (~ ng4332)  &  (~ ng4349)  &  (~ ng4358) ) ;
 assign wire33832 = ( pg35  &  (~ ng4340)  &  ng4358 ) ;
 assign wire33834 = ( pg35  &  (~ ng4340)  &  ng4349  &  (~ ng4358) ) ;
 assign wire33836 = ( wire3384 ) | ( (~ pg35)  &  ng4366 ) ;
 assign wire33837 = ( wire33817  &  wire33818 ) | ( wire33820  &  wire33821 ) ;
 assign wire33838 = ( wire33823  &  wire33824 ) | ( wire33826  &  wire33827 ) ;
 assign wire33839 = ( wire3385 ) | ( ng4322  &  (~ ng4515)  &  wire33830 ) ;
 assign wire33842 = ( wire33836 ) | ( wire33837 ) | ( wire33838 ) | ( wire33839 ) ;
 assign wire33846 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33847 = ( ng5607  &  pg35 ) ;
 assign wire33850 = ( (~ ng632)  &  pg35 ) ;
 assign wire33851 = ( (~ pg9048)  &  (~ ng562) ) | ( ng559  &  (~ ng562) ) ;
 assign wire33854 = ( (~ pg9048)  &  (~ ng562) ) | ( ng559  &  (~ ng562) ) ;
 assign wire33857 = ( (~ pg9048)  &  ng562 ) | ( ng559  &  ng562 ) ;
 assign wire33860 = ( (~ pg9048)  &  ng562 ) | ( ng559  &  ng562 ) ;
 assign wire33862 = ( wire3370 ) | ( ng14708  &  wire33850  &  wire33851 ) ;
 assign wire33865 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33866 = ( ng3590  &  pg35 ) ;
 assign wire33869 = ( pg35  &  (~ ng2051)  &  (~ ng2060) ) | ( pg35  &  (~ ng2060)  &  ng2028 ) ;
 assign wire33870 = ( ng2028  &  pg35 ) ;
 assign wire33871 = ( pg35  &  wire6319 ) | ( pg35  &  ng14367  &  wire30342 ) ;
 assign wire33873 = ( wire3351 ) | ( (~ ng27882)  &  wire33871 ) ;
 assign wire33875 = ( pg35  &  (~ ng2675)  &  (~ ng2681) ) ;
 assign wire33877 = ( ng2685  &  pg35 ) ;
 assign wire33879 = ( ng25439  &  wire33877 ) | ( ng2675  &  ng2681  &  (~ ng25439) ) ;
 assign wire33886 = ( pg35  &  ng3161  &  ng3155  &  (~ ng3167) ) ;
 assign wire33887 = ( ng2331 ) | ( (~ ng2287) ) ;
 assign wire33888 = ( pg35  &  ng17405  &  (~ wire33887) ) | ( pg35  &  ng26737  &  (~ wire33887) ) ;
 assign wire33889 = ( ng2295  &  pg35 ) ;
 assign wire33895 = ( pg35  &  wire6172 ) | ( pg35  &  ng14367  &  wire30555 ) ;
 assign wire33896 = ( ng2208  &  pg35 ) ;
 assign wire33898 = ( wire3327 ) | ( (~ ng27796)  &  wire33895 ) ;
 assign wire33902 = ( ng6263  &  pg35 ) ;
 assign wire33903 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33908 = ( (~ pg35)  &  ng4423 ) | ( pg35  &  ng4575  &  ng4581 ) ;
 assign wire33909 = ( (~ pg73)  &  pg35  &  ng4581 ) | ( (~ pg72)  &  pg35  &  ng4581 ) ;
 assign wire33912 = ( ng3554  &  pg35 ) ;
 assign wire33913 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33916 = ( pg35  &  (~ pg11678)  &  ng749 ) | ( pg35  &  ng736  &  ng749 ) ;
 assign wire33917 = ( (~ ng749)  &  pg35 ) ;
 assign wire33918 = ( wire3292 ) | ( (~ ng24875)  &  wire33916 ) | ( wire28810  &  wire33916 ) ;
 assign wire33919 = ( ng5615  &  pg35 ) ;
 assign wire33920 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33922 = ( ng2089  &  pg35 ) ;
 assign wire33924 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33925 = ( ng3909  &  pg35 ) ;
 assign wire33926 = ( wire3281 ) | ( ng11626  &  ng11584  &  wire33924 ) ;
 assign wire33927 = ( (~ pg35)  &  ng2902 ) | ( pg35  &  ng2917 ) ;
 assign wire33931 = ( pg35  &  (~ ng2485)  &  (~ ng2453)  &  ng2441 ) ;
 assign wire33934 = ( pg35  &  ng2445  &  (~ ng2476)  &  ng2453 ) ;
 assign wire33936 = ( pg35  &  ng2476  &  (~ ng2453)  &  ng2429 ) ;
 assign wire33937 = ( ng2449  &  pg35 ) ;
 assign wire33938 = ( ng2504  &  pg35 ) ;
 assign wire33939 = ( ng2485  &  ng2437  &  (~ ng2476) ) ;
 assign wire33943 = ( ng2433  &  (~ ng25400) ) | ( (~ ng25476)  &  wire33937 ) ;
 assign wire33944 = ( wire3267 ) | ( wire3268 ) | ( wire3269 ) | ( wire3274 ) ;
 assign wire33949 = ( pg35  &  (~ pg16693)  &  (~ pg14518)  &  (~ pg16659) ) ;
 assign wire33950 = ( (~ pg16775)  &  (~ pg13966) ) ;
 assign wire33954 = ( pg35  &  (~ pg16693)  &  (~ pg14518)  &  pg11418 ) ;
 assign wire33955 = ( (~ pg16659)  &  pg13966 ) ;
 assign wire33956 = ( ng2287  &  pg35 ) ;
 assign wire33960 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33961 = ( ng6585  &  pg35 ) ;
 assign wire33962 = ( wire3256 ) | ( ng10491  &  ng12716  &  wire33960 ) ;
 assign wire33963 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33964 = ( ng6633  &  pg35 ) ;
 assign wire33970 = ( pg72  &  pg35  &  ng4581 ) | ( pg35  &  ng4575  &  ng4581 ) ;
 assign wire33971 = ( (~ pg35)  &  ng4543 ) | ( ng4543  &  (~ ng4581) ) | ( (~ pg73)  &  pg35  &  ng4581 ) ;
 assign wire33973 = ( pg35  &  (~ pg11678)  &  ng767 ) | ( pg35  &  ng736  &  ng767 ) ;
 assign wire33974 = ( (~ ng767)  &  pg35 ) ;
 assign wire33975 = ( wire3240 ) | ( ng28504  &  wire33973 ) | ( (~ wire28813)  &  wire33973 ) ;
 assign wire33976 = ( ng6259  &  pg35 ) ;
 assign wire33977 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33979 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33980 = ( ng3945  &  pg35 ) ;
 assign wire33983 = ( pg35  &  ng2841  &  (~ ng2748) ) ;
 assign wire33985 = ( pg35  &  ng2841  &  ng2748 ) ;
 assign wire33988 = ( pg35  &  (~ ng2279)  &  (~ ng2273) ) ;
 assign wire33990 = ( pg35  &  ng2279  &  ng2273 ) ;
 assign wire33993 = ( (~ ng25309)  &  wire33990 ) | ( pg35  &  ng2283  &  ng25309 ) ;
 assign wire33996 = ( (~ pg35)  &  ng1379 ) | ( pg35  &  ng1384  &  ng13242 ) ;
 assign wire33997 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire33998 = ( ng5559  &  pg35 ) ;
 assign wire34000 = ( pg35  &  ng4284 ) | ( pg35  &  (~ ng4180) ) ;
 assign wire34001 = ( ng5905  &  pg35 ) ;
 assign wire34004 = ( pg35  &  (~ ng5462)  &  ng5467 ) ;
 assign wire34005 = ( (~ ng5467)  &  ng5462 ) ;
 assign wire34007 = ( (~ ng23630)  &  wire34005 ) | ( pg35  &  ng5471  &  ng23630 ) ;
 assign wire34008 = ( ng2227 ) | ( (~ ng2197) ) ;
 assign wire34009 = ( ng2169  &  pg35 ) ;
 assign wire34010 = ( pg35  &  ng26703  &  (~ wire34008) ) | ( pg35  &  ng17321  &  (~ wire34008) ) ;
 assign wire34016 = ( (~ ng20841)  &  ng21193  &  (~ ng20982)  &  (~ ng19968) ) ;
 assign wire34017 = ( (~ ng20014)  &  (~ ng19919)  &  (~ ng21127)  &  (~ ng21256) ) ;
 assign wire34022 = ( (~ ng20841)  &  (~ ng21193)  &  ng20982  &  (~ ng19968) ) ;
 assign wire34023 = ( (~ ng20014)  &  (~ ng19919)  &  (~ ng21127)  &  (~ ng21256) ) ;
 assign wire34028 = ( (~ ng20841)  &  (~ ng21193)  &  (~ ng20982)  &  (~ ng19968) ) ;
 assign wire34029 = ( (~ ng20014)  &  (~ ng19919)  &  ng21127  &  (~ ng21256) ) ;
 assign wire34034 = ( (~ ng20841)  &  (~ ng21193)  &  (~ ng20982)  &  (~ ng19968) ) ;
 assign wire34035 = ( (~ ng20014)  &  (~ ng19919)  &  (~ ng21127)  &  ng21256 ) ;
 assign wire34038 = ( (~ ng20841)  &  (~ ng19968)  &  (~ ng20014)  &  (~ ng19919) ) ;
 assign wire34041 = ( ng20841  &  (~ ng19968)  &  (~ ng20014)  &  (~ ng19919) ) ;
 assign wire34044 = ( (~ ng20841)  &  ng19968  &  (~ ng20014)  &  (~ ng19919) ) ;
 assign wire34047 = ( (~ ng20841)  &  (~ ng19968)  &  ng20014  &  (~ ng19919) ) ;
 assign wire34050 = ( (~ ng20841)  &  (~ ng19968)  &  (~ ng20014)  &  ng19919 ) ;
 assign wire34051 = ( wire34016  &  wire34017 ) | ( wire34022  &  wire34023 ) ;
 assign wire34052 = ( wire34028  &  wire34029 ) | ( wire34034  &  wire34035 ) ;
 assign wire34053 = ( ni24685  &  wire34038 ) | ( ni24685  &  wire34041 ) ;
 assign wire34054 = ( ni24685  &  wire34044 ) | ( ni24685  &  wire34047 ) ;
 assign wire34057 = ( wire34051 ) | ( wire34054 ) | ( ni24685  &  wire34050 ) ;
 assign wire34059 = ( (~ ng4064)  &  (~ ng4057)  &  ng4076 ) ;
 assign wire34061 = ( ng4141  &  (~ ng4125) ) | ( (~ ng4125)  &  ng4082 ) ;
 assign wire34062 = ( pg134  &  pg113 ) | ( pg99  &  pg113  &  ng37 ) ;
 assign wire34063 = ( pg134  &  pg113 ) | ( pg99  &  pg113  &  ng37 ) ;
 assign wire34064 = ( (~ pg35) ) | ( (~ ng3817)  &  (~ ng5471) ) ;
 assign wire34065 = ( (~ pg35) ) | ( (~ ng3466)  &  (~ ng6163) ) ;
 assign wire34066 = ( (~ pg35) ) | ( (~ ng5124)  &  (~ ng5817) ) ;
 assign wire34067 = ( (~ pg35) ) | ( (~ ng6509)  &  (~ ng3115) ) ;
 assign wire34070 = ( ng26365  &  wire34064  &  wire34067 ) ;
 assign wire34071 = ( (~ pg35) ) | ( (~ ng5124)  &  (~ ng5471) ) ;
 assign wire34072 = ( (~ pg35) ) | ( (~ ng4427)  &  (~ ng5817)  &  (~ ng4420) ) ;
 assign wire34073 = ( (~ pg35) ) | ( (~ ng3466)  &  (~ ng6163) ) ;
 assign wire34074 = ( (~ pg35) ) | ( (~ ng6509)  &  (~ ng3115) ) ;
 assign wire34076 = ( wire34071  &  wire34072  &  wire34073  &  wire34074 ) ;
 assign wire34078 = ( pg35  &  ng3466  &  (~ ng6509) ) ;
 assign wire34079 = ( (~ pg35) ) | ( (~ ng3817)  &  (~ ng6163)  &  (~ ng3115) ) ;
 assign wire34082 = ( (~ pg35) ) | ( (~ ng3466)  &  (~ ng6509) ) ;
 assign wire34083 = ( pg35  &  (~ ng3817)  &  (~ ng6163)  &  ng3115 ) ;
 assign wire34085 = ( (~ pg35) ) | ( (~ ng5124)  &  (~ ng6163) ) ;
 assign wire34086 = ( (~ pg35) ) | ( (~ ng6509)  &  (~ ng5817) ) ;
 assign wire34088 = ( (~ pg35) ) | ( (~ ng6163)  &  (~ ng5471) ) ;
 assign wire34089 = ( (~ pg35) ) | ( (~ ng6509)  &  (~ ng5817) ) ;
 assign wire34091 = ( (~ pg35) ) | ( (~ ng6163)  &  (~ ng5471) ) ;
 assign wire34092 = ( (~ pg35) ) | ( (~ ng5124)  &  (~ ng6509) ) ;
 assign wire34094 = ( (~ pg35)  &  wire34071  &  wire34072 ) | ( (~ ng6509)  &  wire34071  &  wire34072 ) ;
 assign wire34095 = ( (~ pg35)  &  wire34071  &  wire34072 ) | ( (~ ng6163)  &  wire34071  &  wire34072 ) ;
 assign wire34096 = ( wire3183 ) | ( wire34065  &  wire34066  &  wire34070 ) ;
 assign wire34099 = ( wire32354  &  wire34076 ) | ( wire32355  &  wire34076 ) | ( (~ wire32354)  &  (~ wire32355)  &  wire34094 ) ;
 assign wire34101 = ( wire3184 ) | ( wire3185 ) | ( wire3186 ) | ( wire3187 ) ;
 assign wire34104 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29957) ) | ( ng28180  &  (~ wire30003) ) ;
 assign wire34105 = ( ng27511  &  ng17653  &  (~ ni17529) ) | ( ng27511  &  ng17653  &  (~ wire30041) ) ;
 assign wire34106 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30000) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30000)  &  (~ wire30045) ) ;
 assign wire34109 = ( (~ ng31327)  &  wire34104  &  wire34105  &  wire34106 ) ;
 assign wire34111 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29957) ) | ( ng28180  &  (~ wire30003) ) ;
 assign wire34112 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34113 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30000) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30000)  &  (~ wire30045) ) ;
 assign wire34116 = ( (~ ng31327)  &  wire34111  &  wire34112  &  wire34113 ) ;
 assign wire34118 = ( (~ ng28180) ) | ( ng13156  &  wire29957  &  wire30003 ) ;
 assign wire34120 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34121 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire29997)  &  (~ wire30045) ) ;
 assign wire34124 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29957) ) | ( ng28180  &  (~ wire30003) ) ;
 assign wire34126 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34127 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire29997)  &  (~ wire30045) ) ;
 assign wire34130 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29957) ) | ( ng28180  &  (~ wire30003) ) ;
 assign wire34132 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34133 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire29997)  &  (~ wire30045) ) ;
 assign wire34136 = ( (~ ng28180)  &  (~ ng13156) ) | ( (~ ng28180)  &  (~ wire29957) ) | ( (~ ng28180)  &  (~ wire30003) ) ;
 assign wire34138 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34139 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire29997)  &  (~ wire30045) ) ;
 assign wire34142 = ( ng28180  &  ng13156  &  wire29957  &  wire30003 ) ;
 assign wire34144 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire30041) ) ;
 assign wire34145 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire29997)  &  (~ wire30045) ) ;
 assign wire34149 = ( ng28180  &  ni17529  &  wire29997  &  (~ wire30000) ) ;
 assign wire34150 = ( (~ ng27511) ) | ( (~ ni18740) ) | ( (~ wire29959)  &  (~ wire30002) ) ;
 assign wire34151 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34154 = ( ng28180  &  ng13156  &  wire29957  &  wire30045 ) ;
 assign wire34156 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire29997) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ wire29997)  &  (~ wire30003) ) ;
 assign wire34159 = ( ng28180  &  ni17529  &  (~ wire30000)  &  wire30042 ) ;
 assign wire34160 = ( (~ ng30614)  &  (~ wire29984)  &  (~ wire29985)  &  wire34159 ) ;
 assign wire34161 = ( (~ ng31021)  &  (~ ng31376)  &  wire34109 ) | ( ng31021  &  (~ ng31376)  &  wire34116 ) ;
 assign wire34166 = ( wire3170 ) | ( wire3171 ) | ( wire34161 ) ;
 assign wire34167 = ( wire3172 ) | ( wire3173 ) | ( wire3174 ) | ( wire3175 ) ;
 assign wire34169 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire29996) ) ;
 assign wire34170 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34173 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire29996) ) ;
 assign wire34174 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34177 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire29996) ) ;
 assign wire34178 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34181 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire29996) ) ;
 assign wire34182 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34185 = ( (~ ng27511) ) | ( (~ ng17653)  &  (~ ni17529) ) | ( (~ ng17653)  &  (~ wire29996) ) ;
 assign wire34186 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34188 = ( (~ ng13156) ) | ( (~ wire29957) ) | ( (~ wire29962)  &  (~ wire30003) ) ;
 assign wire34189 = ( (~ ng13156)  &  wire34188 ) | ( (~ wire29963)  &  wire34188 ) | ( (~ wire29966)  &  wire34188 ) ;
 assign wire34193 = ( (~ ng30937)  &  (~ wire29984)  &  (~ wire29985)  &  wire34149 ) ;
 assign wire34198 = ( wire3159 ) | ( wire3160 ) | ( wire3167 ) ;
 assign wire34199 = ( wire3161 ) | ( wire3162 ) | ( wire3163 ) | ( wire3164 ) ;
 assign wire34201 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ wire30003)  &  (~ wire30042) ) ;
 assign wire34202 = ( (~ ng13156)  &  wire34201 ) | ( (~ wire29957)  &  wire34201 ) | ( (~ wire30045)  &  wire34201 ) ;
 assign wire34203 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29937) ) | ( ng28180  &  (~ wire30000) ) ;
 assign wire34204 = ( (~ ni18740)  &  ni18785  &  wire29966 ) | ( ni18785  &  (~ wire29962)  &  wire29966 ) ;
 assign wire34206 = ( (~ wire29984)  &  (~ wire29985)  &  wire34203  &  wire34204 ) ;
 assign wire34207 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34208 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34211 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34212 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34215 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34216 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34219 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34220 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34225 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34226 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34229 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29937) ) | ( ng28180  &  (~ wire30000) ) ;
 assign wire34230 = ( (~ wire29984)  &  (~ wire29985)  &  wire34229 ) ;
 assign wire34231 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ wire30003)  &  (~ wire30042) ) ;
 assign wire34232 = ( (~ ng13156) ) | ( (~ wire29957) ) | ( (~ wire29962)  &  (~ wire30045) ) ;
 assign wire34234 = ( (~ ni18785)  &  wire34231  &  wire34232 ) | ( (~ wire29966)  &  wire34231  &  wire34232 ) ;
 assign wire34235 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ wire30003)  &  (~ wire30042) ) ;
 assign wire34236 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34239 = ( ng28180  &  (~ ng13156) ) | ( ng28180  &  (~ wire29937) ) | ( ng28180  &  (~ wire30000) ) ;
 assign wire34241 = ( (~ ng13156) ) | ( (~ wire29957) ) | ( (~ wire30003)  &  (~ wire30045) ) ;
 assign wire34242 = ( (~ ng13156)  &  wire34241 ) | ( (~ wire29963)  &  wire34241 ) | ( (~ wire29966)  &  wire34241 ) ;
 assign wire34244 = ( (~ ng31566)  &  (~ wire29984)  &  (~ wire29985)  &  wire34159 ) ;
 assign wire34248 = ( ng33496 ) | ( wire3148 ) | ( wire3149 ) | ( wire3150 ) ;
 assign wire34256 = ( (~ pg113) ) | ( (~ pg99)  &  (~ pg134) ) | ( (~ pg134)  &  (~ ng37) ) ;
 assign wire34258 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ ni17529)  &  (~ wire30045) ) | ( (~ wire30042)  &  (~ wire30045) ) ;
 assign wire34259 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34262 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ wire30003)  &  (~ wire30042) ) ;
 assign wire34263 = ( (~ ng13156) ) | ( (~ wire29957) ) | ( (~ wire29962)  &  (~ wire30045) ) ;
 assign wire34265 = ( (~ ni18785)  &  wire34262  &  wire34263 ) | ( (~ wire29966)  &  wire34262  &  wire34263 ) ;
 assign wire34266 = ( (~ ni18740)  &  (~ ni17529) ) | ( (~ ni17529)  &  (~ wire30003) ) | ( (~ ni18740)  &  (~ wire30042) ) | ( (~ wire30003)  &  (~ wire30042) ) ;
 assign wire34267 = ( (~ ni18740)  &  (~ ni18785) ) | ( (~ ni18785)  &  (~ wire29962) ) | ( (~ ni18740)  &  (~ wire29966) ) | ( (~ wire29962)  &  (~ wire29966) ) ;
 assign wire34271 = ( (~ ng31566)  &  (~ wire29984)  &  (~ wire29985)  &  wire34159 ) ;
 assign wire34275 = ( ng33496 ) | ( wire3137 ) | ( wire3138 ) | ( wire3139 ) ;
 assign wire34278 = ( pg73  &  ng4332  &  (~ ng4366)  &  (~ ng4311) ) | ( (~ pg73)  &  (~ ng4332)  &  (~ ng4366)  &  (~ ng4311) ) ;
 assign wire34279 = ( ng2941  &  ng2936 ) | ( ng2912  &  ng2917 ) ;
 assign wire34280 = ( ng2960  &  ng2965 ) | ( ng2902  &  ng2907 ) ;
 assign wire34281 = ( ng2975  &  ng2970 ) | ( ng2950  &  ng2955 ) ;
 assign wire34290 = ( (~ pg113) ) | ( (~ pg99)  &  (~ pg134) ) | ( (~ pg134)  &  (~ ng37) ) ;
 assign wire34292 = ( (~ wire1457) ) | ( (~ wire1411) ) ;
 assign wire34294 = ( (~ pg113) ) | ( (~ pg99)  &  (~ pg134) ) | ( (~ pg134)  &  (~ ng37) ) ;
 assign wire34296 = ( (~ wire1457) ) | ( (~ wire1411) ) ;


endmodule

