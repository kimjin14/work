module apex2 (
	i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, 
	i_27_, i_14_, i_3_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, 
	i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, 
	i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, 
	i_37_, o_1_, o_2_, o_0_);

input i_30_;
input i_20_;
input i_9_;
input i_10_;
input i_7_;
input i_8_;
input i_5_;
input i_6_;
input i_27_;
input i_14_;
input i_3_;
input i_28_;
input i_13_;
input i_4_;
input i_25_;
input i_12_;
input i_1_;
input i_26_;
input i_11_;
input i_2_;
input i_23_;
input i_18_;
input i_24_;
input i_17_;
input i_0_;
input i_21_;
input i_16_;
input i_22_;
input i_15_;
input i_32_;
input i_31_;
input i_34_;
input i_33_;
input i_19_;
input i_36_;
input i_35_;
input i_38_;
input i_29_;
input i_37_;
output o_1_;
output o_2_;
output o_0_;
wire wire59;
wire n_n1827;
wire n_n1829;
wire n_n1812;
wire n_n1866;
wire n_n1865;
wire n_n1558;
wire n_n1559;
wire n_n1542;
wire wire204;
wire wire232;
wire wire296;
wire wire462;
wire wire493;
wire wire58;
wire n_n1441;
wire wire43;
wire n_n1443;
wire wire302;
wire n_n1433;
wire n_n1425;
wire wire54;
wire n_n1396;
wire wire10;
wire n_n1404;
wire n_n1390;
wire wire415;
wire n_n1372;
wire n_n1369;
wire n_n1429;
wire n_n1454;
wire wire42;
wire n_n1489;
wire n_n1353;
wire n_n1361;
wire wire428;
wire n_n1423;
wire n_n1295;
wire n_n1439;
wire wire3;
wire n_n1438;
wire n_n1397;
wire n_n1274;
wire n_n1334;
wire n_n1368;
wire n_n1216;
wire wire290;
wire n_n1391;
wire n_n1478;
wire n_n1307;
wire n_n1374;
wire n_n805;
wire n_n1504;
wire n_n841;
wire n_n853;
wire n_n793;
wire n_n1315;
wire n_n1092;
wire n_n1406;
wire n_n1466;
wire wire224;
wire n_n1278;
wire n_n787;
wire n_n1197;
wire n_n762;
wire n_n1038;
wire n_n1314;
wire n_n1375;
wire wire13;
wire n_n1141;
wire n_n544;
wire n_n1486;
wire n_n1408;
wire n_n1318;
wire n_n504;
wire wire297;
wire n_n416;
wire wire243;
wire n_n1305;
wire n_n1118;
wire n_n358;
wire n_n1048;
wire wire76;
wire n_n307;
wire n_n1263;
wire n_n620;
wire n_n1288;
wire n_n1018;
wire n_n1400;
wire n_n819;
wire n_n394;
wire n_n458;
wire n_n391;
wire n_n1055;
wire n_n372;
wire n_n1179;
wire wire257;
wire n_n300;
wire n_n1225;
wire n_n461;
wire n_n294;
wire n_n301;
wire n_n880;
wire n_n1100;
wire wire51;
wire wire260;
wire n_n437;
wire n_n571;
wire n_n1258;
wire wire263;
wire n_n825;
wire n_n1437;
wire n_n1340;
wire n_n180;
wire n_n132;
wire n_n152;
wire n_n1300;
wire n_n1472;
wire wire50;
wire wire52;
wire wire85;
wire wire223;
wire wire264;
wire wire266;
wire wire388;
wire wire446;
wire wire529;
wire n_n1871;
wire n_n1147;
wire n_n1089;
wire wire79;
wire wire298;
wire wire410;
wire wire516;
wire wire530;
wire n_n1580;
wire n_n1326;
wire wire245;
wire wire277;
wire wire340;
wire wire432;
wire wire533;
wire wire532;
wire n_n1579;
wire wire80;
wire wire536;
wire wire535;
wire n_n1581;
wire n_n1519;
wire n_n1419;
wire n_n1302;
wire n_n1401;
wire wire283;
wire n_n1192;
wire n_n1257;
wire n_n1323;
wire n_n1279;
wire n_n1133;
wire n_n1128;
wire n_n1303;
wire n_n1285;
wire n_n586;
wire n_n1523;
wire n_n1322;
wire n_n269;
wire wire259;
wire n_n242;
wire n_n1202;
wire wire258;
wire n_n355;
wire n_n1345;
wire n_n371;
wire wire53;
wire n_n316;
wire n_n735;
wire n_n315;
wire n_n984;
wire n_n1458;
wire n_n1213;
wire n_n177;
wire n_n1241;
wire n_n179;
wire n_n245;
wire n_n1431;
wire wire62;
wire wire70;
wire wire72;
wire wire212;
wire wire239;
wire wire250;
wire wire288;
wire wire539;
wire wire537;
wire n_n1881;
wire n_n576;
wire n_n1499;
wire wire47;
wire wire307;
wire wire541;
wire wire540;
wire n_n195;
wire n_n1563;
wire wire86;
wire wire244;
wire wire275;
wire wire483;
wire wire500;
wire wire543;
wire n_n1548;
wire n_n1568;
wire n_n1497;
wire n_n1384;
wire n_n1393;
wire n_n1282;
wire n_n839;
wire n_n1311;
wire n_n263;
wire n_n363;
wire n_n584;
wire n_n1033;
wire n_n309;
wire n_n317;
wire n_n712;
wire n_n284;
wire n_n1028;
wire n_n178;
wire n_n460;
wire wire9;
wire wire57;
wire wire77;
wire wire83;
wire wire372;
wire wire380;
wire wire395;
wire wire503;
wire n_n1387;
wire n_n1306;
wire n_n1359;
wire n_n1080;
wire n_n1254;
wire wire411;
wire n_n1144;
wire n_n1585;
wire n_n1422;
wire wire8;
wire wire38;
wire wire90;
wire wire112;
wire wire127;
wire wire546;
wire n_n1556;
wire n_n1459;
wire n_n1377;
wire n_n1312;
wire n_n820;
wire n_n706;
wire wire205;
wire n_n1191;
wire n_n608;
wire n_n1058;
wire n_n916;
wire n_n629;
wire n_n338;
wire wire261;
wire n_n129;
wire n_n26;
wire wire463;
wire wire548;
wire wire547;
wire n_n1574;
wire n_n1575;
wire n_n1578;
wire n_n1576;
wire n_n1577;
wire n_n1571;
wire n_n1573;
wire n_n1572;
wire n_n1545;
wire n_n1251;
wire n_n998;
wire wire124;
wire wire132;
wire wire236;
wire wire355;
wire wire550;
wire n_n1583;
wire n_n1582;
wire wire252;
wire wire555;
wire n_n1584;
wire wire214;
wire wire227;
wire wire265;
wire wire267;
wire wire559;
wire n_n329;
wire wire312;
wire wire468;
wire wire126;
wire wire128;
wire wire196;
wire wire452;
wire wire363;
wire wire420;
wire wire455;
wire wire566;
wire wire568;
wire n_n1511;
wire n_n130;
wire wire475;
wire n_n849;
wire n_n1059;
wire wire222;
wire n_n18;
wire n_n21;
wire wire299;
wire wire342;
wire wire478;
wire wire572;
wire wire48;
wire wire385;
wire wire67;
wire wire418;
wire wire578;
wire wire576;
wire wire253;
wire wire330;
wire wire405;
wire wire583;
wire n_n1847;
wire wire585;
wire n_n1889;
wire wire4;
wire wire56;
wire wire226;
wire wire282;
wire n_n1856;
wire wire81;
wire wire377;
wire n_n1825;
wire n_n1854;
wire wire71;
wire n_n1861;
wire wire319;
wire wire599;
wire wire598;
wire wire597;
wire n_n1718;
wire wire317;
wire wire365;
wire wire601;
wire wire600;
wire wire233;
wire wire246;
wire wire492;
wire wire63;
wire wire268;
wire wire361;
wire wire431;
wire wire508;
wire wire301;
wire wire441;
wire wire608;
wire wire360;
wire wire610;
wire n_n1149;
wire wire447;
wire wire21;
wire wire235;
wire n_n1846;
wire wire61;
wire wire616;
wire wire615;
wire wire614;
wire n_n1892;
wire wire35;
wire n_n1837;
wire wire249;
wire wire311;
wire wire329;
wire wire344;
wire n_n1862;
wire wire218;
wire wire310;
wire wire315;
wire wire387;
wire wire408;
wire n_n1870;
wire wire78;
wire wire271;
wire wire278;
wire wire346;
wire wire627;
wire wire320;
wire wire416;
wire wire630;
wire wire629;
wire n_n1719;
wire wire248;
wire wire634;
wire wire632;
wire wire88;
wire n_n1697;
wire n_n1720;
wire n_n1716;
wire n_n1715;
wire n_n1723;
wire wire55;
wire n_n1684;
wire wire440;
wire wire644;
wire wire643;
wire n_n1896;
wire wire12;
wire wire254;
wire wire381;
wire wire430;
wire wire429;
wire n_n1852;
wire n_n1843;
wire wire75;
wire wire654;
wire wire276;
wire wire423;
wire wire656;
wire wire664;
wire wire663;
wire wire29;
wire wire273;
wire wire491;
wire n_n1690;
wire wire668;
wire wire383;
wire wire669;
wire wire390;
wire wire671;
wire wire675;
wire wire674;
wire wire676;
wire n_n1844;
wire wire270;
wire wire677;
wire n_n1821;
wire wire272;
wire wire379;
wire wire482;
wire wire74;
wire wire688;
wire wire687;
wire wire68;
wire wire206;
wire wire519;
wire wire692;
wire wire691;
wire n_n1882;
wire wire524;
wire wire694;
wire wire693;
wire n_n1714;
wire wire470;
wire wire697;
wire n_n1703;
wire wire295;
wire wire286;
wire wire700;
wire wire306;
wire wire398;
wire wire464;
wire wire705;
wire wire704;
wire n_n1704;
wire wire708;
wire n_n1705;
wire wire712;
wire wire289;
wire wire327;
wire wire335;
wire wire456;
wire wire41;
wire wire305;
wire wire717;
wire wire716;
wire wire256;
wire n_n1701;
wire n_n1702;
wire wire274;
wire wire351;
wire wire724;
wire wire723;
wire wire394;
wire wire322;
wire wire727;
wire n_n1713;
wire wire731;
wire wire730;
wire wire284;
wire wire734;
wire wire66;
wire wire502;
wire n_n1875;
wire n_n1873;
wire n_n1831;
wire n_n1816;
wire wire739;
wire n_n1818;
wire n_n1834;
wire n_n1835;
wire wire744;
wire wire745;
wire n_n1884;
wire wire457;
wire wire262;
wire wire465;
wire wire510;
wire wire755;
wire wire82;
wire n_n1712;
wire wire760;
wire wire515;
wire wire768;
wire wire771;
wire n_n1877;
wire wire784;
wire wire788;
wire wire792;
wire n_n1887;
wire wire353;
wire wire484;
wire wire489;
wire wire437;
wire wire18;
wire wire435;
wire wire422;
wire wire434;
wire wire349;
wire wire404;
wire wire413;
wire wire37;
wire wire44;
wire wire211;
wire wire65;
wire wire436;
wire wire803;
wire wire802;
wire wire95;
wire wire96;
wire wire143;
wire wire147;
wire wire202;
wire wire458;
wire wire221;
wire wire231;
wire wire251;
wire wire314;
wire wire334;
wire wire338;
wire wire343;
wire wire345;
wire wire356;
wire wire367;
wire wire373;
wire wire384;
wire wire402;
wire wire406;
wire wire425;
wire wire438;
wire wire454;
wire wire495;
wire wire498;
wire wire517;
wire wire521;
wire wire522;
wire wire526;
wire wire544;
wire wire557;
wire wire582;
wire wire590;
wire wire593;
wire wire604;
wire wire603;
wire wire606;
wire wire624;
wire wire635;
wire wire638;
wire wire657;
wire wire661;
wire wire666;
wire wire679;
wire wire683;
wire wire698;
wire wire710;
wire wire713;
wire wire721;
wire wire735;
wire wire741;
wire wire740;
wire wire759;
wire wire758;
wire wire767;
wire wire22;
wire wire34;
wire wire101;
wire wire102;
wire wire105;
wire wire107;
wire wire110;
wire wire111;
wire wire117;
wire wire118;
wire wire119;
wire wire120;
wire wire121;
wire wire123;
wire wire125;
wire wire129;
wire wire130;
wire wire133;
wire wire134;
wire wire142;
wire wire150;
wire wire151;
wire wire153;
wire wire154;
wire wire158;
wire wire160;
wire wire161;
wire wire163;
wire wire164;
wire wire166;
wire wire167;
wire wire169;
wire wire172;
wire wire174;
wire wire176;
wire wire177;
wire wire178;
wire wire183;
wire wire184;
wire wire185;
wire wire187;
wire wire189;
wire wire190;
wire wire191;
wire wire192;
wire wire194;
wire wire195;
wire wire197;
wire wire198;
wire wire200;
wire wire201;
wire wire234;
wire wire304;
wire wire336;
wire wire339;
wire wire350;
wire wire412;
wire wire417;
wire wire424;
wire wire427;
wire wire439;
wire wire451;
wire wire469;
wire wire471;
wire wire494;
wire wire497;
wire wire507;
wire wire512;
wire wire812;
wire wire813;
wire wire818;
wire wire825;
wire wire829;
wire wire833;
wire wire834;
wire wire841;
wire wire843;
wire wire849;
wire wire850;
wire wire857;
wire wire863;
wire wire864;
wire wire868;
wire wire875;
wire wire877;
wire wire878;
wire wire881;
wire wire884;
wire wire891;
wire wire903;
wire wire904;
wire wire906;
wire wire910;
wire wire911;
wire wire916;
wire wire918;
wire wire919;
wire wire920;
wire wire924;
wire wire925;
wire wire926;
wire wire928;
wire wire933;
wire wire935;
wire wire937;
wire wire939;
wire wire940;
wire wire941;
wire wire942;
wire wire943;
wire wire945;
wire wire948;
wire wire950;
wire wire953;
wire wire955;
wire wire956;
wire wire957;
wire wire958;
wire wire959;
wire wire960;
wire wire961;
wire wire965;
wire wire966;
wire wire967;
wire wire968;
wire wire969;
wire wire977;
wire wire978;
wire wire981;
wire wire983;
wire wire987;
wire wire988;
wire wire990;
wire wire991;
wire wire992;
wire wire993;
wire wire994;
wire wire996;
wire wire999;
wire wire1000;
wire wire1002;
wire wire1007;
wire wire1008;
wire wire1009;
wire wire1010;
wire wire1011;
wire wire1012;
wire wire1014;
wire wire1015;
wire wire1017;
wire wire1019;
wire wire1020;
wire wire1021;
wire wire1022;
wire wire1023;
wire wire1024;
wire wire1029;
wire wire1030;
wire wire1032;
wire wire1033;
wire wire1040;
wire wire1041;
wire wire1043;
wire wire1044;
wire wire1045;
wire wire1048;
wire wire1050;
wire wire1051;
wire wire1052;
wire wire1053;
wire wire1054;
wire wire1055;
wire wire1056;
wire wire1057;
wire wire1058;
wire wire1059;
wire wire1060;
wire wire1061;
wire wire1062;
wire wire1064;
wire wire1066;
wire wire1069;
wire wire1070;
wire wire1077;
wire wire1080;
wire wire1081;
wire wire1082;
wire wire1086;
wire wire1087;
wire wire1089;
wire wire1091;
wire wire1095;
wire wire1097;
wire wire1100;
wire wire1101;
wire wire1105;
wire wire1106;
wire wire1108;
wire wire1111;
wire wire1112;
wire wire1113;
wire wire1114;
wire wire1121;
wire wire1123;
wire wire1125;
wire wire1126;
wire wire1127;
wire wire1128;
wire wire1129;
wire wire1130;
wire wire1131;
wire wire1132;
wire wire1133;
wire wire1134;
wire wire1135;
wire wire1136;
wire wire1137;
wire wire1139;
wire wire1140;
wire wire1141;
wire wire1142;
wire wire1143;
wire wire1146;
wire wire1147;
wire wire1148;
wire wire1150;
wire wire1152;
wire wire1156;
wire wire1157;
wire wire1159;
wire wire1161;
wire wire1162;
wire wire1163;
wire wire1164;
wire wire1167;
wire wire1168;
wire wire1169;
wire wire1170;
wire wire1172;
wire wire1173;
wire wire1176;
wire wire1180;
wire wire1181;
wire wire1184;
wire wire1186;
wire wire1187;
wire wire1189;
wire wire1190;
wire wire1191;
wire wire1197;
wire wire1198;
wire wire1201;
wire wire1202;
wire wire1203;
wire wire1208;
wire wire1211;
wire wire1212;
wire wire1214;
wire wire1215;
wire wire1218;
wire wire1227;
wire wire1230;
wire wire1234;
wire wire1235;
wire wire1236;
wire wire1238;
wire wire1239;
wire wire1240;
wire wire1241;
wire wire1242;
wire wire1247;
wire wire1249;
wire wire1253;
wire wire1256;
wire wire1257;
wire wire1258;
wire wire1259;
wire wire1260;
wire wire1263;
wire wire1264;
wire wire1265;
wire wire1266;
wire wire1267;
wire wire1268;
wire wire1271;
wire wire1274;
wire wire1277;
wire wire1279;
wire wire1280;
wire wire1281;
wire wire1283;
wire wire1284;
wire wire1286;
wire wire1288;
wire wire1289;
wire wire1290;
wire wire1291;
wire wire1293;
wire wire1296;
wire wire1303;
wire wire1305;
wire wire1308;
wire wire1309;
wire wire1314;
wire wire1316;
wire wire1317;
wire wire1318;
wire wire1319;
wire wire1320;
wire wire1323;
wire wire1324;
wire wire1325;
wire wire1330;
wire wire1337;
wire wire1338;
wire wire1340;
wire wire1341;
wire wire1342;
wire wire1343;
wire wire1347;
wire wire1349;
wire wire1350;
wire wire1351;
wire wire1356;
wire wire1357;
wire wire1367;
wire wire1372;
wire wire1377;
wire wire1379;
wire wire1382;
wire wire1383;
wire wire1384;
wire wire1392;
wire wire1397;
wire wire1399;
wire wire1403;
wire wire1404;
wire wire1405;
wire wire1406;
wire wire1408;
wire wire1409;
wire wire1412;
wire wire1413;
wire wire1414;
wire wire1416;
wire wire1417;
wire wire1419;
wire wire1421;
wire wire1423;
wire wire1426;
wire wire1428;
wire wire1429;
wire wire1430;
wire wire1431;
wire wire1432;
wire wire1433;
wire wire1434;
wire wire1435;
wire wire1436;
wire wire1437;
wire wire1439;
wire wire1443;
wire wire1449;
wire wire1450;
wire wire1456;
wire wire1457;
wire wire1460;
wire wire1461;
wire wire1463;
wire wire1464;
wire wire1465;
wire wire1470;
wire wire1473;
wire wire1474;
wire wire1476;
wire wire1477;
wire wire1480;
wire wire1481;
wire wire1482;
wire wire1483;
wire wire1484;
wire wire1485;
wire wire1486;
wire wire1490;
wire wire1491;
wire wire1492;
wire wire1493;
wire wire1495;
wire wire1498;
wire wire1499;
wire wire1500;
wire wire1501;
wire wire1502;
wire wire1503;
wire wire1506;
wire wire1507;
wire wire1508;
wire wire1509;
wire wire1511;
wire wire1514;
wire wire1523;
wire wire1525;
wire wire1531;
wire wire1532;
wire wire1534;
wire wire1535;
wire wire1539;
wire wire1542;
wire wire1546;
wire wire1548;
wire wire1549;
wire wire1550;
wire wire1551;
wire wire1552;
wire wire1553;
wire wire1554;
wire wire1559;
wire wire1561;
wire wire1564;
wire wire1565;
wire wire1566;
wire wire1567;
wire wire1568;
wire wire1570;
wire wire1572;
wire wire1573;
wire wire1574;
wire wire1576;
wire wire1577;
wire wire1580;
wire wire1581;
wire wire1582;
wire wire1583;
wire wire1585;
wire wire1586;
wire wire1587;
wire wire1589;
wire wire1591;
wire wire1592;
wire wire1593;
wire wire1597;
wire wire1600;
wire wire1603;
wire wire1604;
wire wire1607;
wire wire1608;
wire wire1611;
wire wire1615;
wire wire1618;
wire wire1619;
wire wire1622;
wire wire1623;
wire wire1624;
wire wire1625;
wire wire1628;
wire wire1632;
wire wire1634;
wire wire1635;
wire wire1636;
wire wire1637;
wire wire1638;
wire wire1640;
wire wire1649;
wire wire1650;
wire wire1651;
wire wire1652;
wire wire1653;
wire wire1654;
wire wire1656;
wire wire1657;
wire wire1659;
wire wire1661;
wire wire1663;
wire wire1665;
wire wire1668;
wire wire1669;
wire wire1670;
wire wire1672;
wire wire1675;
wire wire1676;
wire wire1677;
wire wire1678;
wire wire1682;
wire wire1683;
wire wire1684;
wire wire1685;
wire wire1686;
wire wire1688;
wire wire1689;
wire wire1690;
wire wire1691;
wire wire1692;
wire wire1693;
wire wire1694;
wire wire1695;
wire wire1696;
wire wire1697;
wire wire1698;
wire wire1699;
wire wire1700;
wire wire1701;
wire wire1702;
wire wire1703;
wire wire1704;
wire wire1706;
wire wire1709;
wire wire1710;
wire wire1715;
wire wire1716;
wire wire1717;
wire wire1718;
wire wire1719;
wire wire1721;
wire wire1722;
wire wire1726;
wire wire1730;
wire wire1731;
wire wire1738;
wire wire1746;
wire wire1747;
wire wire1748;
wire wire1749;
wire wire1750;
wire wire1753;
wire wire1756;
wire wire1757;
wire wire1758;
wire wire1759;
wire wire1766;
wire wire1767;
wire wire1768;
wire wire6876;
wire wire6879;
wire wire6880;
wire wire6881;
wire wire6882;
wire wire6884;
wire wire6885;
wire wire6889;
wire wire6890;
wire wire6891;
wire wire6892;
wire wire6893;
wire wire6894;
wire wire6898;
wire wire6899;
wire wire6901;
wire wire6903;
wire wire6905;
wire wire6906;
wire wire6908;
wire wire6910;
wire wire6912;
wire wire6913;
wire wire6915;
wire wire6917;
wire wire6919;
wire wire6920;
wire wire6922;
wire wire6923;
wire wire6924;
wire wire6926;
wire wire6927;
wire wire6928;
wire wire6930;
wire wire6931;
wire wire6933;
wire wire6934;
wire wire6935;
wire wire6936;
wire wire6937;
wire wire6938;
wire wire6939;
wire wire6941;
wire wire6942;
wire wire6943;
wire wire6947;
wire wire6948;
wire wire6949;
wire wire6951;
wire wire6952;
wire wire6953;
wire wire6955;
wire wire6957;
wire wire6958;
wire wire6959;
wire wire6960;
wire wire6961;
wire wire6962;
wire wire6963;
wire wire6967;
wire wire6971;
wire wire6973;
wire wire6977;
wire wire6979;
wire wire6982;
wire wire6984;
wire wire6989;
wire wire6990;
wire wire6993;
wire wire6994;
wire wire6996;
wire wire6997;
wire wire6998;
wire wire7000;
wire wire7001;
wire wire7004;
wire wire7005;
wire wire7006;
wire wire7007;
wire wire7009;
wire wire7010;
wire wire7011;
wire wire7014;
wire wire7017;
wire wire7018;
wire wire7019;
wire wire7022;
wire wire7025;
wire wire7026;
wire wire7027;
wire wire7028;
wire wire7029;
wire wire7031;
wire wire7033;
wire wire7036;
wire wire7037;
wire wire7040;
wire wire7041;
wire wire7043;
wire wire7044;
wire wire7045;
wire wire7046;
wire wire7050;
wire wire7051;
wire wire7052;
wire wire7053;
wire wire7054;
wire wire7055;
wire wire7057;
wire wire7058;
wire wire7059;
wire wire7060;
wire wire7062;
wire wire7063;
wire wire7064;
wire wire7068;
wire wire7069;
wire wire7070;
wire wire7072;
wire wire7073;
wire wire7074;
wire wire7075;
wire wire7076;
wire wire7079;
wire wire7080;
wire wire7082;
wire wire7083;
wire wire7084;
wire wire7085;
wire wire7086;
wire wire7087;
wire wire7089;
wire wire7090;
wire wire7093;
wire wire7094;
wire wire7095;
wire wire7096;
wire wire7097;
wire wire7098;
wire wire7099;
wire wire7102;
wire wire7103;
wire wire7104;
wire wire7105;
wire wire7108;
wire wire7110;
wire wire7111;
wire wire7114;
wire wire7115;
wire wire7116;
wire wire7117;
wire wire7119;
wire wire7120;
wire wire7121;
wire wire7123;
wire wire7126;
wire wire7130;
wire wire7134;
wire wire7135;
wire wire7136;
wire wire7137;
wire wire7139;
wire wire7140;
wire wire7141;
wire wire7142;
wire wire7143;
wire wire7145;
wire wire7148;
wire wire7151;
wire wire7152;
wire wire7153;
wire wire7157;
wire wire7158;
wire wire7159;
wire wire7160;
wire wire7161;
wire wire7162;
wire wire7163;
wire wire7165;
wire wire7166;
wire wire7167;
wire wire7169;
wire wire7172;
wire wire7173;
wire wire7174;
wire wire7175;
wire wire7176;
wire wire7177;
wire wire7178;
wire wire7179;
wire wire7181;
wire wire7183;
wire wire7185;
wire wire7186;
wire wire7187;
wire wire7188;
wire wire7189;
wire wire7190;
wire wire7191;
wire wire7192;
wire wire7195;
wire wire7197;
wire wire7199;
wire wire7203;
wire wire7204;
wire wire7205;
wire wire7208;
wire wire7210;
wire wire7211;
wire wire7212;
wire wire7214;
wire wire7215;
wire wire7216;
wire wire7217;
wire wire7218;
wire wire7219;
wire wire7221;
wire wire7224;
wire wire7226;
wire wire7228;
wire wire7229;
wire wire7230;
wire wire7234;
wire wire7235;
wire wire7238;
wire wire7239;
wire wire7240;
wire wire7242;
wire wire7243;
wire wire7244;
wire wire7247;
wire wire7248;
wire wire7250;
wire wire7252;
wire wire7254;
wire wire7255;
wire wire7256;
wire wire7257;
wire wire7258;
wire wire7259;
wire wire7261;
wire wire7264;
wire wire7265;
wire wire7266;
wire wire7267;
wire wire7268;
wire wire7269;
wire wire7271;
wire wire7272;
wire wire7273;
wire wire7274;
wire wire7275;
wire wire7276;
wire wire7277;
wire wire7281;
wire wire7282;
wire wire7284;
wire wire7285;
wire wire7286;
wire wire7288;
wire wire7290;
wire wire7295;
wire wire7296;
wire wire7297;
wire wire7298;
wire wire7299;
wire wire7301;
wire wire7306;
wire wire7308;
wire wire7309;
wire wire7310;
wire wire7311;
wire wire7312;
wire wire7316;
wire wire7317;
wire wire7319;
wire wire7320;
wire wire7321;
wire wire7322;
wire wire7323;
wire wire7324;
wire wire7325;
wire wire7327;
wire wire7328;
wire wire7329;
wire wire7330;
wire wire7331;
wire wire7332;
wire wire7333;
wire wire7334;
wire wire7335;
wire wire7336;
wire wire7337;
wire wire7339;
wire wire7340;
wire wire7341;
wire wire7342;
wire wire7343;
wire wire7344;
wire wire7345;
wire wire7348;
wire wire7349;
wire wire7350;
wire wire7351;
wire wire7352;
wire wire7353;
wire wire7354;
wire wire7355;
wire wire7356;
wire wire7357;
wire wire7358;
wire wire7361;
wire wire7362;
wire wire7363;
wire wire7364;
wire wire7365;
wire wire7366;
wire wire7367;
wire wire7368;
wire wire7370;
wire wire7371;
wire wire7372;
wire wire7373;
wire wire7374;
wire wire7375;
wire wire7377;
wire wire7379;
wire wire7380;
wire wire7383;
wire wire7385;
wire wire7386;
wire wire7387;
wire wire7388;
wire wire7390;
wire wire7393;
wire wire7394;
wire wire7395;
wire wire7397;
wire wire7399;
wire wire7400;
wire wire7402;
wire wire7406;
wire wire7407;
wire wire7409;
wire wire7411;
wire wire7412;
wire wire7413;
wire wire7415;
wire wire7417;
wire wire7419;
wire wire7420;
wire wire7423;
wire wire7424;
wire wire7425;
wire wire7426;
wire wire7427;
wire wire7428;
wire wire7430;
wire wire7431;
wire wire7432;
wire wire7433;
wire wire7435;
wire wire7437;
wire wire7439;
wire wire7441;
wire wire7443;
wire wire7445;
wire wire7446;
wire wire7447;
wire wire7448;
wire wire7452;
wire wire7454;
wire wire7456;
wire wire7457;
wire wire7458;
wire wire7459;
wire wire7461;
wire wire7462;
wire wire7464;
wire wire7465;
wire wire7466;
wire wire7469;
wire wire7470;
wire wire7473;
wire wire7474;
wire wire7477;
wire wire7479;
wire wire7483;
wire wire7485;
wire wire7487;
wire wire7488;
wire wire7491;
wire wire7492;
wire wire7493;
wire wire7494;
wire wire7495;
wire wire7500;
wire wire7502;
wire wire7503;
wire wire7504;
wire wire7507;
wire wire7508;
wire wire7510;
wire wire7511;
wire wire7512;
wire wire7516;
wire wire7519;
wire wire7521;
wire wire7522;
wire wire7523;
wire wire7525;
wire wire7526;
wire wire7529;
wire wire7531;
wire wire7532;
wire wire7534;
wire wire7536;
wire wire7537;
wire wire7538;
wire wire7541;
wire wire7543;
wire wire7545;
wire wire7547;
wire wire7548;
wire wire7549;
wire wire7552;
wire wire7553;
wire wire7554;
wire wire7555;
wire wire7559;
wire wire7561;
wire wire7562;
wire wire7565;
wire wire7566;
wire wire7567;
wire wire7570;
wire wire7572;
wire wire7574;
wire wire7576;
wire wire7577;
wire wire7578;
wire wire7580;
wire wire7582;
wire wire7585;
wire wire7586;
wire wire7587;
wire wire7588;
wire wire7591;
wire wire7592;
wire wire7595;
wire wire7596;
wire wire7598;
wire wire7600;
wire wire7602;
wire wire7603;
wire wire7609;
wire wire7612;
wire wire7615;
wire wire7616;
wire wire7618;
wire wire7619;
wire wire7621;
wire wire7622;
wire wire7626;
wire wire7627;
wire wire7629;
wire wire7631;
wire wire7632;
wire wire7636;
wire wire7638;
wire wire7639;
wire wire7640;
wire wire7642;
wire wire7644;
wire wire7646;
wire wire7647;
wire wire7648;
wire wire7651;
wire wire7652;
wire wire7653;
wire wire7655;
wire wire7657;
wire wire7661;
wire wire7666;
wire wire7669;
wire wire7670;
wire wire7673;
wire wire7676;
wire wire7677;
wire wire7678;
wire wire7680;
wire wire7682;
wire wire7686;
wire wire7689;
wire wire7690;
wire wire7691;
wire wire7696;
wire wire7699;
wire wire7701;
wire wire7702;
wire wire7703;
wire wire7704;
wire wire7705;
wire wire7706;
wire wire7708;
wire wire7711;
wire wire7714;
wire wire7716;
wire wire7717;
wire wire7718;
wire wire7721;
wire wire7722;
wire wire7723;
wire wire7724;
wire wire7725;
wire wire7726;
wire wire7727;
wire wire7728;
wire wire7731;
wire wire7732;
wire wire7733;
wire wire7734;
wire wire7735;
wire wire7736;
wire wire7737;
wire wire7738;
wire wire7740;
wire wire7741;
wire wire7743;
wire wire7744;
wire wire7746;
wire wire7747;
wire wire7749;
wire wire7750;
wire wire7751;
wire wire7753;
wire wire7757;
wire wire7761;
wire wire7763;
wire wire7765;
wire wire7766;
wire wire7769;
wire wire7771;
wire wire7772;
wire wire7773;
wire wire7774;
wire wire7776;
wire wire7777;
wire wire7778;
wire wire7781;
wire wire7782;
wire wire7784;
wire wire7785;
wire wire7787;
wire wire7789;
wire wire7791;
wire wire7793;
wire wire7794;
wire wire7795;
wire wire7798;
wire wire7802;
wire wire7803;
wire wire7806;
wire wire7807;
wire wire7808;
wire wire7810;
wire wire7811;
wire wire7812;
wire wire7813;
wire wire7817;
wire wire7819;
wire wire7820;
wire wire7821;
wire wire7822;
wire wire7823;
wire wire7825;
wire wire7826;
wire wire7827;
wire wire7828;
wire wire7829;
wire wire7830;
wire wire7831;
wire wire7832;
wire wire7834;
wire wire7835;
wire wire7836;
wire wire7837;
wire wire7838;
wire wire7839;
wire wire7840;
wire wire7842;
wire wire7843;
wire wire7844;
wire wire7845;
wire wire7846;
wire wire7847;
wire wire7849;
wire wire7851;
wire wire7852;
wire wire7853;
wire wire7854;
wire wire7855;
wire wire7856;
wire wire7857;
wire wire7858;
wire wire7859;
wire wire7860;
wire wire7862;
wire wire7863;
wire wire7864;
wire wire7866;
wire wire7867;
wire wire7868;
wire wire7869;
wire wire7870;
wire wire7871;
wire wire7874;
wire wire7875;
wire wire7878;
wire wire7879;
wire wire7881;
wire wire7882;
wire wire7885;
wire wire7886;
wire wire7887;
wire wire7888;
wire wire7889;
wire wire7890;
wire wire7892;
wire wire7893;
wire wire7895;
wire wire7896;
wire wire7897;
wire wire7898;
wire wire7899;
wire wire7900;
wire wire7901;
wire wire7902;
wire wire7903;
wire wire7906;
wire wire7907;
wire wire7909;
wire wire7910;
wire wire7911;
wire wire7912;
wire wire7913;
wire wire7914;
wire wire7915;
wire wire7916;
wire wire7917;
wire wire7918;
wire wire7920;
wire wire7921;
wire wire7923;
wire wire7926;
wire wire7927;
wire wire7930;
wire wire7931;
wire wire7932;
wire wire7935;
wire wire7936;
wire wire7938;
wire wire7940;
wire wire7941;
wire wire7942;
wire wire7945;
wire wire7946;
wire wire7947;
wire wire7949;
wire wire7952;
wire wire7953;
wire wire7954;
wire wire7957;
wire wire7958;
wire wire7959;
wire wire7960;
wire wire7961;
wire wire7963;
wire wire7964;
wire wire7965;
wire wire7968;
wire wire7969;
wire wire7971;
wire wire7976;
wire wire7978;
wire wire7979;
wire wire7980;
wire wire7981;
wire wire7984;
wire wire7986;
wire wire7989;
wire wire7990;
wire wire7991;
wire wire7994;
wire wire7997;
wire wire7999;
wire wire8002;
wire wire8003;
wire wire8006;
wire wire8007;
wire wire8008;
wire wire8010;
wire wire8014;
wire wire8016;
wire wire8019;
wire wire8021;
wire wire8022;
wire wire8023;
wire wire8026;
wire wire8027;
wire wire8028;
wire wire8029;
wire wire8030;
wire wire8031;
wire wire8035;
wire wire8036;
wire wire8037;
wire wire8039;
wire wire8041;
wire wire8042;
wire wire8043;
wire wire8046;
wire wire8047;
wire wire8049;
wire wire8052;
wire wire8054;
wire wire8056;
wire wire8057;
wire wire8061;
wire wire8062;
wire wire8065;
wire wire8067;
wire wire8071;
wire wire8072;
wire wire8077;
wire wire8079;
wire wire8082;
wire wire8084;
wire wire8085;
wire wire8086;
wire wire8090;
wire wire8091;
wire wire8093;
wire wire8094;
wire wire8096;
assign o_1_ = ( n_n1684 ) | ( wire7250 ) | ( wire7252 ) | ( wire7257 ) ;
 assign o_2_ = ( n_n1816 ) | ( wire7714 ) | ( wire7746 ) | ( wire7747 ) ;
 assign o_0_ = ( n_n1558 ) | ( n_n1559 ) | ( n_n1542 ) | ( wire8096 ) ;
 assign wire59 = ( (~ i_33_)  &  i_37_ ) ;
 assign n_n1827 = ( n_n1862 ) | ( wire7370 ) | ( wire7371 ) | ( wire7383 ) ;
 assign n_n1829 = ( n_n1870 ) | ( wire7407 ) | ( i_38_  &  wire627 ) ;
 assign n_n1812 = ( wire7432 ) | ( wire7433 ) | ( wire7435 ) | ( wire7441 ) ;
 assign n_n1866 = ( wire990 ) | ( wire991 ) | ( wire992 ) | ( wire993 ) ;
 assign n_n1865 = ( wire983 ) | ( wire987 ) | ( wire7727 ) | ( wire7728 ) ;
 assign n_n1558 = ( wire960 ) | ( wire961 ) | ( i_36_  &  wire548 ) ;
 assign n_n1559 = ( wire7771 ) | ( i_36_  &  wire566 ) ;
 assign n_n1542 = ( n_n1548 ) | ( n_n1545 ) | ( wire7923 ) | ( wire8079 ) ;
 assign wire204 = ( (~ i_11_)  &  (~ i_19_) ) ;
 assign wire232 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign wire296 = ( (~ i_23_)  &  (~ i_21_) ) ;
 assign wire462 = ( n_n1443  &  wire79  &  n_n460 ) ;
 assign wire493 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  wire227 ) ;
 assign wire58 = ( (~ i_28_)  &  (~ i_26_) ) ;
 assign n_n1441 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_) ) ;
 assign wire43 = ( (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n1443 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire302 = ( (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1433 = ( (~ i_32_)  &  (~ i_31_)  &  i_34_ ) ;
 assign n_n1425 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_26_) ) ;
 assign wire54 = ( (~ i_23_)  &  (~ i_24_) ) ;
 assign n_n1396 = ( i_25_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire10 = ( (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n1404 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign n_n1390 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign wire415 = ( (~ i_14_)  &  (~ i_12_) ) ;
 assign n_n1372 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign n_n1369 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign n_n1429 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign n_n1454 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire42 = ( (~ i_28_)  &  (~ i_29_) ) ;
 assign n_n1489 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign n_n1353 = ( i_9_  &  (~ i_10_)  &  (~ i_8_) ) ;
 assign n_n1361 = ( (~ i_35_)  &  i_38_ ) ;
 assign wire428 = ( (~ i_25_)  &  (~ i_24_) ) ;
 assign n_n1423 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_24_) ) ;
 assign n_n1295 = ( i_34_  &  i_37_ ) ;
 assign n_n1439 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire3 = ( i_30_ ) | ( i_32_ ) ;
 assign n_n1438 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign n_n1397 = ( (~ i_34_)  &  i_35_ ) ;
 assign n_n1274 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_17_) ) ;
 assign n_n1334 = ( i_31_  &  i_34_ ) ;
 assign n_n1368 = ( (~ i_28_)  &  i_29_ ) ;
 assign n_n1216 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_) ) ;
 assign wire290 = ( (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1391 = ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1478 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_) ) ;
 assign n_n1307 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign n_n1374 = ( i_34_  &  i_33_ ) ;
 assign n_n805 = ( i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n1504 = ( i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign n_n841 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n853 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_) ) ;
 assign n_n793 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_) ) ;
 assign n_n1315 = ( (~ i_9_)  &  i_7_  &  (~ i_12_) ) ;
 assign n_n1092 = ( i_20_  &  (~ i_23_)  &  (~ i_21_) ) ;
 assign n_n1406 = ( (~ i_27_)  &  (~ i_28_)  &  i_29_ ) ;
 assign n_n1466 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_) ) ;
 assign wire224 = ( (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n1278 = ( (~ i_7_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n787 = ( i_3_  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign n_n1197 = ( (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign n_n762 = ( (~ i_30_)  &  (~ i_32_)  &  n_n1197 ) ;
 assign n_n1038 = ( i_9_  &  (~ i_8_)  &  (~ i_3_) ) ;
 assign n_n1314 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n1375 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire13 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n_n1141 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_12_) ) ;
 assign n_n544 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7086 ) ;
 assign n_n1486 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign n_n1408 = ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1318 = ( (~ i_35_)  &  i_37_ ) ;
 assign n_n504 = ( (~ i_33_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire297 = ( (~ i_18_)  &  n_n1278  &  wire404 ) ;
 assign n_n416 = ( (~ i_8_)  &  (~ i_18_)  &  n_n1278  &  wire404 ) ;
 assign wire243 = ( (~ i_32_)  &  (~ i_29_) ) ;
 assign n_n1305 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n1118 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n358 = ( n_n1278  &  n_n1408  &  n_n1279 ) ;
 assign n_n1048 = ( i_9_  &  (~ i_13_)  &  i_18_ ) ;
 assign wire76 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  n_n1144 ) ;
 assign n_n307 = ( n_n1307  &  n_n1048  &  n_n1144 ) ;
 assign n_n1263 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n620 = ( n_n1307  &  n_n1263  &  n_n1306 ) ;
 assign n_n1288 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign n_n1018 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign n_n1400 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_17_) ) ;
 assign n_n819 = ( i_9_  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign n_n394 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7425 ) ;
 assign n_n458 = ( n_n1443  &  n_n1278  &  n_n1279 ) ;
 assign n_n391 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7426 ) ;
 assign n_n1055 = ( i_9_  &  (~ i_13_)  &  i_11_ ) ;
 assign n_n372 = ( n_n1055  &  n_n461  &  wire7411 ) ;
 assign n_n1179 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire257 = ( (~ i_24_)  &  (~ i_22_)  &  wire7265 ) ;
 assign n_n300 = ( (~ i_24_)  &  (~ i_22_)  &  n_n1179  &  wire7265 ) ;
 assign n_n1225 = ( (~ i_28_)  &  i_34_  &  (~ i_29_) ) ;
 assign n_n461 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_) ) ;
 assign n_n294 = ( n_n461  &  wire7411  &  wire7412 ) ;
 assign n_n301 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n880 = ( i_36_  &  (~ i_35_) ) ;
 assign n_n1100 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_) ) ;
 assign wire51 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279 ) ;
 assign wire260 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n437 = ( (~ i_5_)  &  (~ i_6_)  &  wire260  &  n_n1279 ) ;
 assign n_n571 = ( i_35_  &  i_37_ ) ;
 assign n_n1258 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_) ) ;
 assign wire263 = ( (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n825 = ( (~ i_17_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign n_n1437 = ( i_34_  &  (~ i_33_)  &  (~ i_35_) ) ;
 assign n_n1340 = ( (~ i_32_)  &  i_34_  &  (~ i_33_) ) ;
 assign n_n180 = ( (~ i_9_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n132 = ( (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n152 = ( (~ i_4_)  &  (~ i_1_)  &  (~ i_0_) ) ;
 assign n_n1300 = ( (~ i_33_)  &  i_38_ ) ;
 assign n_n1472 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire50 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  n_n1279 ) ;
 assign wire52 = ( (~ i_28_)  &  (~ i_22_)  &  n_n1454 ) ;
 assign wire85 = ( (~ i_32_)  &  n_n1307  &  n_n1100 ) ;
 assign wire223 = ( (~ i_9_)  &  (~ i_10_)  &  n_n1307  &  n_n1303 ) ;
 assign wire264 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire266 = ( i_34_  &  i_38_ ) ;
 assign wire388 = ( (~ i_33_)  &  i_38_  &  wire61 ) ;
 assign wire446 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire529 = ( wire262 ) | ( wire436 ) | ( i_19_  &  wire18 ) ;
 assign n_n1871 = ( wire1215 ) | ( wire1218 ) | ( wire7511 ) | ( wire7512 ) ;
 assign n_n1147 = ( (~ i_7_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1089 = ( (~ i_7_)  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign wire79 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_)  &  i_36_ ) ;
 assign wire298 = ( (~ i_24_)  &  i_34_ ) ;
 assign wire410 = ( n_n1375  &  n_n1400  &  wire244  &  wire7789 ) ;
 assign wire516 = ( n_n1441  &  n_n1400  &  n_n1472  &  wire7785 ) ;
 assign wire530 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign n_n1580 = ( wire935 ) | ( wire7793 ) | ( wire7794 ) | ( wire7795 ) ;
 assign n_n1326 = ( (~ i_28_)  &  (~ i_34_)  &  i_29_ ) ;
 assign wire245 = ( (~ i_23_)  &  (~ i_24_)  &  i_21_  &  i_34_ ) ;
 assign wire277 = ( (~ i_30_)  &  (~ i_28_) ) ;
 assign wire340 = ( i_14_  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire432 = ( (~ i_20_)  &  n_n1406  &  n_n1213  &  wire7000 ) ;
 assign wire533 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire532 = ( wire43  &  n_n1315 ) | ( wire263  &  n_n1323 ) ;
 assign n_n1579 = ( wire7806 ) | ( wire7807 ) | ( wire7808 ) ;
 assign wire80 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire536 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign wire535 = ( n_n1315  &  n_n1263 ) | ( n_n1285  &  n_n1322 ) ;
 assign n_n1581 = ( wire916 ) | ( wire918 ) | ( wire7812 ) | ( wire7813 ) ;
 assign n_n1519 = ( i_12_  &  (~ i_24_)  &  i_17_ ) ;
 assign n_n1419 = ( (~ i_34_)  &  i_35_  &  i_38_ ) ;
 assign n_n1302 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n1401 = ( i_7_  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign wire283 = ( (~ i_8_)  &  (~ i_2_) ) ;
 assign n_n1192 = ( i_9_  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign n_n1257 = ( (~ i_28_)  &  i_33_  &  (~ i_29_) ) ;
 assign n_n1323 = ( (~ i_9_)  &  i_7_  &  (~ i_13_) ) ;
 assign n_n1279 = ( (~ i_4_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n_n1133 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n1128 = ( (~ i_28_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n1303 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign n_n1285 = ( (~ i_9_)  &  i_7_  &  (~ i_14_) ) ;
 assign n_n586 = ( (~ i_13_)  &  i_12_  &  i_11_ ) ;
 assign n_n1523 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign n_n1322 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n269 = ( n_n1307  &  n_n1314  &  n_n1306 ) ;
 assign wire259 = ( (~ i_8_)  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n242 = ( n_n1278  &  n_n1279  &  wire259 ) ;
 assign n_n1202 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_ ) ;
 assign wire258 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n355 = ( n_n1278  &  n_n1279  &  wire258 ) ;
 assign n_n1345 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign n_n371 = ( n_n819  &  n_n1279  &  wire7413 ) ;
 assign wire53 = ( (~ i_28_)  &  n_n1197  &  n_n1523 ) ;
 assign n_n316 = ( (~ i_28_)  &  (~ i_32_)  &  n_n1197  &  n_n1523 ) ;
 assign n_n735 = ( (~ i_13_)  &  i_18_  &  i_19_ ) ;
 assign n_n315 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7423 ) ;
 assign n_n984 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_ ) ;
 assign n_n1458 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_) ) ;
 assign n_n1213 = ( (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign n_n177 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign n_n1241 = ( i_34_  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n179 = ( (~ i_23_)  &  (~ i_18_)  &  (~ i_17_) ) ;
 assign n_n245 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign n_n1431 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_) ) ;
 assign wire62 = ( n_n1406  &  n_n1213  &  wire7491 ) ;
 assign wire70 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_22_)  &  wire7266 ) ;
 assign wire72 = ( (~ i_12_)  &  n_n1307  &  n_n1303 ) ;
 assign wire212 = ( n_n1278  &  n_n1279  &  wire7492 ) ;
 assign wire239 = ( (~ i_25_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire250 = ( i_38_  &  n_n1278  &  n_n1279 ) ;
 assign wire288 = ( (~ i_28_)  &  i_34_  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire539 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire537 = ( n_n1439  &  n_n1340 ) | ( n_n1423  &  wire7409 ) ;
 assign n_n1881 = ( wire7493 ) | ( wire7494 ) | ( wire7495 ) ;
 assign n_n576 = ( (~ i_32_)  &  i_36_  &  (~ i_35_) ) ;
 assign n_n1499 = ( (~ i_28_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire47 = ( (~ i_23_)  &  (~ i_34_)  &  i_35_ ) ;
 assign wire307 = ( n_n576  &  wire44  &  wire7749  &  wire7847 ) ;
 assign wire541 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire540 = ( n_n329  &  wire468 ) | ( wire67  &  wire367 ) ;
 assign n_n195 = ( n_n1408  &  n_n1118  &  n_n1279 ) ;
 assign n_n1563 = ( wire863 ) | ( wire864 ) | ( wire7874 ) | ( wire7875 ) ;
 assign wire86 = ( i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign wire244 = ( i_34_  &  i_36_ ) ;
 assign wire275 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_  &  wire47 ) ;
 assign wire483 = ( n_n1216  &  n_n1133  &  wire86 ) ;
 assign wire500 = ( n_n1018  &  n_n1128  &  wire86 ) ;
 assign wire543 = ( wire221  &  wire495 ) | ( wire41  &  wire7189 ) ;
 assign n_n1548 = ( n_n1563 ) | ( wire877 ) | ( wire7866 ) | ( wire7882 ) ;
 assign n_n1568 = ( wire7916 ) | ( wire7917 ) | ( wire7920 ) ;
 assign n_n1497 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign n_n1384 = ( i_14_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign n_n1393 = ( (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign n_n1282 = ( (~ i_23_)  &  (~ i_17_)  &  (~ i_21_) ) ;
 assign n_n839 = ( (~ i_9_)  &  (~ i_6_)  &  i_13_ ) ;
 assign n_n1311 = ( (~ i_32_)  &  (~ i_34_)  &  (~ i_33_) ) ;
 assign n_n263 = ( n_n1429  &  n_n1307  &  n_n1303 ) ;
 assign n_n363 = ( n_n1404  &  n_n1307  &  n_n1303 ) ;
 assign n_n584 = ( (~ i_13_)  &  i_12_  &  i_18_ ) ;
 assign n_n1033 = ( i_9_  &  (~ i_8_)  &  i_11_ ) ;
 assign n_n309 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7420 ) ;
 assign n_n317 = ( (~ i_4_)  &  (~ i_2_)  &  wire7419  &  wire7424 ) ;
 assign n_n712 = ( i_10_  &  i_7_  &  (~ i_11_) ) ;
 assign n_n284 = ( n_n819  &  n_n1279  &  n_n735 ) ;
 assign n_n1028 = ( i_9_  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign n_n178 = ( (~ i_13_)  &  (~ i_11_)  &  (~ i_16_) ) ;
 assign n_n460 = ( (~ i_28_)  &  (~ i_32_)  &  i_29_ ) ;
 assign wire9 = ( (~ i_24_)  &  i_38_ ) ;
 assign wire57 = ( (~ i_30_)  &  (~ i_29_) ) ;
 assign wire77 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire83 = ( (~ i_28_)  &  i_22_ ) ;
 assign wire372 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  i_29_ ) ;
 assign wire380 = ( (~ i_33_)  &  i_38_  &  n_n1486 ) ;
 assign wire395 = ( (~ i_24_)  &  i_38_  &  wire71 ) ;
 assign wire503 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_33_)  &  i_38_ ) ;
 assign n_n1387 = ( i_14_  &  (~ i_13_)  &  (~ i_16_) ) ;
 assign n_n1306 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign n_n1359 = ( i_9_  &  (~ i_10_)  &  (~ i_24_) ) ;
 assign n_n1080 = ( (~ i_27_)  &  (~ i_23_)  &  i_21_ ) ;
 assign n_n1254 = ( (~ i_23_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign wire411 = ( (~ i_8_)  &  (~ i_12_) ) ;
 assign n_n1144 = ( (~ i_8_)  &  (~ i_6_)  &  (~ i_12_) ) ;
 assign n_n1585 = ( wire196 ) | ( wire812 ) | ( wire7926 ) | ( wire7927 ) ;
 assign n_n1422 = ( (~ i_32_)  &  i_34_  &  (~ i_35_) ) ;
 assign wire8 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire38 = ( n_n1390  &  n_n1384 ) | ( n_n1400  &  n_n1387 ) ;
 assign wire90 = ( wire1661 ) | ( i_22_  &  wire803 ) ;
 assign wire112 = ( n_n1489  &  wire340  &  wire7682 ) ;
 assign wire127 = ( wire372  &  wire7029 ) ;
 assign wire546 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1556 = ( n_n1585 ) | ( wire90 ) | ( wire7938 ) ;
 assign n_n1459 = ( (~ i_30_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign n_n1377 = ( i_7_  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign n_n1312 = ( (~ i_23_)  &  (~ i_24_)  &  i_21_ ) ;
 assign n_n820 = ( (~ i_30_)  &  (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign n_n706 = ( (~ i_9_)  &  wire204  &  n_n1307  &  n_n1303 ) ;
 assign wire205 = ( (~ i_24_)  &  (~ i_22_) ) ;
 assign n_n1191 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign n_n608 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire7051 ) ;
 assign n_n1058 = ( i_9_  &  (~ i_3_)  &  i_11_ ) ;
 assign n_n916 = ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign n_n629 = ( (~ i_20_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n338 = ( i_19_  &  wire288  &  wire12 ) ;
 assign wire261 = ( (~ i_9_)  &  i_13_  &  n_n1307  &  n_n1303 ) ;
 assign n_n129 = ( (~ i_9_)  &  n_n1307  &  n_n1303  &  wire6881 ) ;
 assign n_n26 = ( i_3_  &  (~ i_4_)  &  (~ i_0_) ) ;
 assign wire463 = ( wire296  &  n_n1443  &  n_n1369  &  n_n1368 ) ;
 assign wire548 = ( wire965 ) | ( wire966 ) | ( wire967 ) | ( wire968 ) ;
 assign wire547 = ( n_n841  &  wire338 ) | ( wire232  &  wire7753 ) ;
 assign n_n1574 = ( wire451 ) | ( wire7952 ) | ( wire7953 ) | ( wire7954 ) ;
 assign n_n1575 = ( wire412 ) | ( wire7963 ) | ( wire7964 ) | ( wire7965 ) ;
 assign n_n1578 = ( wire7978 ) | ( wire7979 ) | ( wire7980 ) | ( wire7981 ) ;
 assign n_n1576 = ( wire195 ) | ( wire7989 ) | ( wire7990 ) | ( wire7991 ) ;
 assign n_n1577 = ( wire8002 ) | ( wire8003 ) | ( i_21_  &  wire688 ) ;
 assign n_n1571 = ( wire174 ) | ( wire176 ) | ( wire177 ) | ( wire8016 ) ;
 assign n_n1573 = ( wire8035 ) | ( wire8036 ) | ( wire8037 ) ;
 assign n_n1572 = ( wire8046 ) | ( wire8047 ) | ( i_21_  &  wire730 ) ;
 assign n_n1545 = ( n_n1571 ) | ( wire8049 ) | ( wire8052 ) | ( wire8054 ) ;
 assign n_n1251 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_16_) ) ;
 assign n_n998 = ( (~ i_25_)  &  (~ i_24_)  &  i_19_ ) ;
 assign wire124 = ( n_n1397  &  n_n1258  &  n_n1257  &  n_n1387 ) ;
 assign wire132 = ( n_n1397  &  n_n1257  &  n_n1384  &  n_n1251 ) ;
 assign wire236 = ( (~ i_28_)  &  i_31_  &  n_n1369 ) ;
 assign wire355 = ( (~ i_28_)  &  i_0_  &  i_29_  &  n_n1369 ) ;
 assign wire550 = ( wire10  &  n_n1282 ) | ( wire290  &  n_n1254 ) ;
 assign n_n1583 = ( wire129 ) | ( wire8061 ) | ( wire8062 ) ;
 assign n_n1582 = ( wire118 ) | ( wire119 ) | ( wire120 ) | ( wire8067 ) ;
 assign wire252 = ( i_34_  &  i_33_  &  n_n1396  &  n_n1375 ) ;
 assign wire555 = ( n_n1315  &  n_n1314 ) | ( n_n1322  &  wire557 ) ;
 assign n_n1584 = ( wire8071 ) | ( wire8072 ) | ( wire236  &  wire555 ) ;
 assign wire214 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  (~ i_29_) ) ;
 assign wire227 = ( (~ i_32_)  &  (~ i_34_)  &  i_36_  &  i_35_ ) ;
 assign wire265 = ( (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire267 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  (~ i_29_) ) ;
 assign wire559 = ( n_n1443  &  n_n1118  &  n_n1279 ) | ( n_n1408  &  n_n1118  &  n_n1279 ) ;
 assign n_n329 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire6920 ) ;
 assign wire312 = ( n_n1443  &  n_n1118  &  n_n1279 ) ;
 assign wire468 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_24_)  &  n_n1128 ) ;
 assign wire126 = ( n_n1438  &  wire6948  &  wire6949 ) ;
 assign wire128 = ( n_n1438  &  wire6948  &  wire7653 ) ;
 assign wire196 = ( n_n1489  &  n_n1393  &  wire1649 ) | ( n_n1489  &  n_n1393  &  wire1650 ) ;
 assign wire452 = ( (~ i_26_)  &  (~ i_24_)  &  (~ i_34_) ) ;
 assign wire363 = ( n_n1369  &  n_n1368  &  n_n1282  &  wire7761 ) ;
 assign wire420 = ( (~ i_14_)  &  i_13_  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire455 = ( wire232  &  wire44  &  wire7749  &  wire7769 ) ;
 assign wire566 = ( wire956 ) | ( wire957 ) | ( wire958 ) | ( wire959 ) ;
 assign wire568 = ( n_n301  &  wire363 ) | ( wire7776  &  wire7777 ) ;
 assign n_n1511 = ( (~ i_28_)  &  i_31_  &  i_34_ ) ;
 assign n_n130 = ( (~ i_17_)  &  (~ i_16_)  &  (~ i_19_) ) ;
 assign wire475 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1353  &  n_n1307 ) ;
 assign n_n849 = ( (~ i_24_)  &  n_n1353  &  n_n1307  &  wire7050 ) ;
 assign n_n1059 = ( (~ i_34_)  &  (~ i_33_)  &  i_35_  &  i_38_ ) ;
 assign wire222 = ( (~ i_20_)  &  n_n1406  &  n_n1213 ) ;
 assign n_n18 = ( (~ i_20_)  &  n_n1406  &  n_n1213  &  wire6893 ) ;
 assign n_n21 = ( (~ i_20_)  &  n_n1406  &  n_n1213  &  wire6890 ) ;
 assign wire299 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_23_)  &  wire7942 ) ;
 assign wire342 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_16_)  &  wire6993 ) ;
 assign wire478 = ( n_n1441  &  n_n1438  &  n_n880  &  wire7831 ) ;
 assign wire572 = ( wire43  &  n_n1315 ) | ( wire263  &  n_n1323 ) ;
 assign wire48 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  n_n1400 ) ;
 assign wire385 = ( i_36_  &  (~ i_35_)  &  n_n1459 ) ;
 assign wire67 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  n_n1213 ) ;
 assign wire418 = ( wire79  &  wire7822 ) ;
 assign wire578 = ( i_3_  &  (~ i_18_) ) | ( (~ i_11_)  &  (~ i_19_) ) ;
 assign wire576 = ( wire221  &  wire367 ) | ( wire41  &  wire384 ) ;
 assign wire253 = ( (~ i_35_)  &  i_38_  &  n_n1439  &  n_n1340 ) ;
 assign wire330 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire71 ) ;
 assign wire405 = ( i_10_  &  i_12_ ) ;
 assign wire583 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign n_n1847 = ( wire1281 ) | ( wire1283 ) | ( wire253  &  wire583 ) ;
 assign wire585 = ( i_14_  &  i_13_ ) | ( i_12_  &  i_17_ ) ;
 assign n_n1889 = ( wire1125 ) | ( wire7615 ) ;
 assign wire4 = ( n_n1307  &  wire361 ) | ( n_n787  &  wire353 ) ;
 assign wire56 = ( (~ i_35_)  &  i_38_  &  n_n1425  &  wire7276 ) ;
 assign wire226 = ( (~ i_31_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire282 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_)  &  wire7272 ) ;
 assign n_n1856 = ( wire1449 ) | ( wire1450 ) | ( wire7282 ) ;
 assign wire81 = ( (~ i_35_)  &  i_38_  &  n_n1454 ) ;
 assign wire377 = ( (~ i_30_)  &  (~ i_28_)  &  n_n1197  &  n_n1523 ) ;
 assign n_n1825 = ( n_n1856 ) | ( wire1457 ) | ( wire7267 ) | ( wire7290 ) ;
 assign n_n1854 = ( wire1428 ) | ( wire1429 ) | ( wire1430 ) | ( wire1431 ) ;
 assign wire71 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign n_n1861 = ( wire1382 ) | ( wire1383 ) | ( wire1384 ) | ( wire7345 ) ;
 assign wire319 = ( (~ i_28_)  &  i_29_  &  n_n1369  &  n_n1274 ) ;
 assign wire599 = ( n_n1425  &  wire6951 ) | ( wire277  &  wire6952 ) ;
 assign wire598 = ( n_n1406  &  wire245 ) | ( n_n1396  &  wire6958 ) ;
 assign wire597 = ( i_21_  &  wire372 ) | ( n_n1302  &  wire6957 ) ;
 assign n_n1718 = ( wire6961 ) | ( wire6962 ) | ( wire6963 ) ;
 assign wire317 = ( i_34_  &  i_37_  &  n_n1018  &  n_n1302 ) ;
 assign wire365 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  i_37_ ) ;
 assign wire601 = ( n_n355  &  wire48 ) | ( n_n358  &  wire221 ) ;
 assign wire600 = ( n_n195  &  wire273 ) | ( n_n437  &  wire256 ) ;
 assign wire233 = ( n_n1406  &  n_n1213  &  n_n629  &  wire6876 ) ;
 assign wire246 = ( (~ i_34_)  &  (~ i_33_)  &  i_35_  &  i_37_ ) ;
 assign wire492 = ( i_35_  &  i_37_  &  n_n1375  &  n_n1311 ) ;
 assign wire63 = ( (~ i_20_)  &  (~ i_23_)  &  n_n1369  &  n_n460 ) ;
 assign wire268 = ( (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire361 = ( (~ i_9_)  &  (~ i_6_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire431 = ( (~ i_11_)  &  (~ i_17_)  &  (~ i_16_)  &  (~ i_19_) ) ;
 assign wire508 = ( n_n1303  &  n_n245  &  wire44  &  wire6899 ) ;
 assign wire301 = ( n_n1141  &  n_n1213  &  wire7053  &  wire7976 ) ;
 assign wire441 = ( (~ i_24_)  &  i_21_  &  (~ i_34_)  &  n_n1425 ) ;
 assign wire608 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire360 = ( (~ i_31_)  &  n_n1307  &  n_n1144 ) ;
 assign wire610 = ( n_n1443  &  wire437 ) | ( n_n1429  &  wire437 ) | ( n_n1443  &  wire891 ) ;
 assign n_n1149 = ( (~ i_32_)  &  wire226 ) ;
 assign wire447 = ( (~ i_28_)  &  (~ i_24_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire21 = ( wire434 ) | ( n_n1118  &  n_n1058  &  wire7415 ) ;
 assign wire235 = ( n_n1197  &  n_n1523  &  wire7466 ) ;
 assign n_n1846 = ( wire1264 ) | ( wire1265 ) | ( wire1266 ) | ( wire1267 ) ;
 assign wire61 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire616 = ( wire1111 ) | ( i_30_  &  n_n1225 ) | ( i_32_  &  n_n1225 ) ;
 assign wire615 = ( i_14_  &  i_13_ ) | ( i_12_  &  i_17_ ) ;
 assign wire614 = ( wire1108 ) | ( i_12_  &  (~ i_24_)  &  i_17_ ) ;
 assign n_n1892 = ( wire1105 ) | ( wire1106 ) | ( wire616  &  wire614 ) ;
 assign wire35 = ( i_30_  &  i_27_ ) | ( i_27_  &  i_32_ ) | ( i_16_  &  i_32_ ) ;
 assign n_n1837 = ( n_n1892 ) | ( wire1097 ) | ( wire7631 ) | ( wire7632 ) ;
 assign wire249 = ( n_n1425  &  wire7276  &  wire7301 ) ;
 assign wire311 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  i_38_ ) ;
 assign wire329 = ( (~ i_24_)  &  i_38_  &  wire77  &  wire78 ) ;
 assign wire344 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign n_n1862 = ( wire1372 ) | ( wire1377 ) | ( wire7357 ) | ( wire7358 ) ;
 assign wire218 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  n_n839 ) ;
 assign wire310 = ( n_n1307  &  n_n1100  &  n_n1311  &  wire7377 ) ;
 assign wire315 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_24_)  &  n_n805 ) ;
 assign wire387 = ( (~ i_34_)  &  i_35_  &  i_38_  &  n_n1302 ) ;
 assign wire408 = ( (~ i_10_)  &  n_n1307  &  n_n841 ) ;
 assign n_n1870 = ( wire1337 ) | ( wire7400 ) | ( n_n1489  &  wire784 ) ;
 assign wire78 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_22_) ) ;
 assign wire271 = ( i_34_  &  (~ i_35_)  &  i_38_  &  n_n1466 ) ;
 assign wire278 = ( (~ i_30_)  &  (~ i_24_) ) ;
 assign wire346 = ( i_13_  &  (~ i_32_)  &  n_n1307  &  n_n1100 ) ;
 assign wire627 = ( wire1330 ) | ( wire52  &  wire223 ) | ( wire52  &  wire261 ) ;
 assign wire320 = ( i_31_  &  i_34_  &  n_n1375 ) ;
 assign wire416 = ( (~ i_14_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire630 = ( n_n1406  &  wire245 ) | ( n_n1396  &  wire6958 ) ;
 assign wire629 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1719 = ( wire1715 ) | ( wire1716 ) | ( wire1717 ) | ( wire6977 ) ;
 assign wire248 = ( i_34_  &  (~ i_35_)  &  i_37_ ) ;
 assign wire634 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) | ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign wire632 = ( wire312  &  wire6937 ) | ( n_n329  &  wire6938 ) ;
 assign wire88 = ( n_n245  &  wire44  &  wire6899 ) ;
 assign n_n1697 = ( wire1564 ) | ( wire1565 ) | ( wire1566 ) | ( wire1567 ) ;
 assign n_n1720 = ( wire1697 ) | ( wire1701 ) | ( wire6989 ) | ( wire6990 ) ;
 assign n_n1716 = ( wire1688 ) | ( wire1689 ) | ( wire1690 ) | ( wire7001 ) ;
 assign n_n1715 = ( wire1682 ) | ( wire1683 ) | ( wire7010 ) | ( wire7011 ) ;
 assign n_n1723 = ( wire1659 ) | ( wire1661 ) | ( i_22_  &  wire803 ) ;
 assign wire55 = ( (~ i_28_)  &  i_29_  &  n_n1369  &  wire7033 ) ;
 assign n_n1684 = ( wire7044 ) | ( wire7045 ) ;
 assign wire440 = ( i_21_  &  (~ i_19_)  &  n_n712 ) ;
 assign wire644 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire643 = ( n_n355  &  wire48 ) | ( n_n358  &  wire221 ) ;
 assign n_n1896 = ( wire1086 ) | ( wire1087 ) | ( wire447  &  wire35 ) ;
 assign wire12 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire254 = ( (~ i_35_)  &  i_38_  &  n_n1305  &  n_n1497 ) ;
 assign wire381 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1288 ) ;
 assign wire430 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire429 = ( (~ i_25_)  &  (~ i_34_)  &  i_35_  &  i_38_ ) ;
 assign n_n1852 = ( wire7452 ) | ( (~ i_31_)  &  wire1288 ) | ( (~ i_31_)  &  wire1289 ) ;
 assign n_n1843 = ( wire1314 ) | ( wire1316 ) | ( n_n316  &  wire755 ) ;
 assign wire75 = ( (~ i_35_)  &  i_38_  &  n_n1423  &  wire7409 ) ;
 assign wire654 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire276 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire78 ) ;
 assign wire423 = ( n_n461  &  wire7411  &  wire7427 ) ;
 assign wire656 = ( n_n372 ) | ( n_n294 ) | ( n_n371 ) | ( n_n284 ) ;
 assign wire664 = ( (~ i_14_)  &  wire233 ) | ( wire314  &  wire7136 ) ;
 assign wire663 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) | ( (~ i_14_)  &  i_13_  &  (~ i_16_) ) ;
 assign wire29 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire273 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  n_n1225 ) ;
 assign wire491 = ( n_n1307  &  n_n1314  &  n_n1144 ) ;
 assign n_n1690 = ( wire7062 ) | ( wire7094 ) | ( i_37_  &  wire768 ) ;
 assign wire668 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire383 = ( n_n461  &  wire79  &  n_n460  &  n_n1254 ) ;
 assign wire669 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire390 = ( (~ i_33_)  &  (~ i_35_)  &  i_38_  &  wire61 ) ;
 assign wire671 = ( n_n372 ) | ( n_n294 ) | ( n_n371 ) | ( n_n284 ) ;
 assign wire675 = ( n_n372 ) | ( n_n294 ) | ( n_n371 ) | ( n_n284 ) ;
 assign wire674 = ( wire435 ) | ( i_19_  &  wire1323 ) | ( i_19_  &  wire1324 ) ;
 assign wire676 = ( n_n372 ) | ( n_n294 ) | ( n_n371 ) | ( n_n284 ) ;
 assign n_n1844 = ( wire1256 ) | ( wire1257 ) | ( wire1258 ) | ( wire1259 ) ;
 assign wire270 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_)  &  n_n1179 ) ;
 assign wire677 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign n_n1821 = ( n_n1846 ) | ( n_n1844 ) | ( wire7477 ) ;
 assign wire272 = ( n_n1307  &  n_n1288  &  n_n1100 ) ;
 assign wire379 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_)  &  n_n1419 ) ;
 assign wire482 = ( (~ i_35_)  &  i_37_  &  n_n1216  &  n_n1241 ) ;
 assign wire74 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  n_n1400 ) ;
 assign wire688 = ( wire189 ) | ( (~ i_16_)  &  wire190 ) | ( (~ i_16_)  &  wire191 ) ;
 assign wire687 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire68 = ( i_9_  &  i_12_ ) ;
 assign wire206 = ( i_38_  &  n_n1307  &  n_n1306 ) ;
 assign wire519 = ( (~ i_12_)  &  n_n1307  &  n_n1303  &  wire9 ) ;
 assign wire692 = ( n_n1439  &  n_n1340 ) | ( n_n1423  &  wire7409 ) ;
 assign wire691 = ( wire71 ) | ( wire430 ) ;
 assign n_n1882 = ( wire7502 ) | ( wire7503 ) | ( wire7504 ) ;
 assign wire524 = ( i_34_  &  i_37_  &  n_n1216  &  wire57 ) ;
 assign wire694 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire693 = ( n_n1401  &  wire6960 ) | ( n_n1391  &  wire7017 ) ;
 assign n_n1714 = ( wire1587 ) | ( wire7110 ) | ( wire7111 ) ;
 assign wire470 = ( (~ i_33_)  &  i_37_  &  n_n1429 ) ;
 assign wire697 = ( wire1542 ) | ( wire7169 ) | ( n_n1437  &  wire698 ) ;
 assign n_n1703 = ( wire7172 ) | ( i_37_  &  wire697 ) ;
 assign wire295 = ( n_n1345  &  n_n576  &  n_n1282  &  wire8010 ) ;
 assign wire286 = ( n_n1307  &  n_n1100  &  wire344  &  wire7523 ) ;
 assign wire700 = ( wire1214 ) | ( (~ i_24_)  &  wire223  &  wire266 ) ;
 assign wire306 = ( n_n1375  &  n_n1213  &  wire7006 ) ;
 assign wire398 = ( (~ i_32_)  &  (~ i_31_)  &  i_34_  &  wire6984 ) ;
 assign wire464 = ( (~ i_23_)  &  (~ i_24_)  &  n_n1433  &  n_n1489 ) ;
 assign wire705 = ( n_n358  &  wire7173 ) | ( n_n355  &  wire7174 ) ;
 assign wire704 = ( n_n1404  &  wire508 ) | ( wire367  &  wire7177 ) ;
 assign n_n1704 = ( wire1525 ) | ( wire7183 ) | ( i_37_  &  wire704 ) ;
 assign wire708 = ( n_n242  &  wire48 ) | ( n_n458  &  wire221 ) ;
 assign n_n1705 = ( wire1511 ) | ( wire7192 ) | ( wire708  &  wire7188 ) ;
 assign wire712 = ( n_n363  &  wire273 ) | ( n_n620  &  wire256 ) ;
 assign wire289 = ( i_13_  &  (~ i_31_)  &  n_n1307  &  n_n841 ) ;
 assign wire327 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  n_n1359 ) ;
 assign wire335 = ( (~ i_10_)  &  n_n819  &  n_n1279 ) ;
 assign wire456 = ( (~ i_25_)  &  (~ i_26_)  &  (~ i_24_)  &  wire7356 ) ;
 assign wire41 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_2_)  &  n_n841 ) ;
 assign wire305 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_31_ ) ;
 assign wire717 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) | ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire716 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire256 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  wire6928 ) ;
 assign n_n1701 = ( wire1498 ) | ( wire1499 ) | ( wire1500 ) | ( wire1501 ) ;
 assign n_n1702 = ( wire1490 ) | ( wire1491 ) | ( wire1493 ) | ( wire7221 ) ;
 assign wire274 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_)  &  wire44 ) ;
 assign wire351 = ( n_n1307  &  n_n1100  &  wire268  &  wire7121 ) ;
 assign wire724 = ( n_n1408  &  wire7827 ) | ( n_n916  &  wire7828 ) ;
 assign wire723 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire394 = ( n_n1118  &  n_n1279  &  n_n1359 ) ;
 assign wire322 = ( i_34_  &  i_33_  &  wire6996  &  wire6997 ) ;
 assign wire727 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1713 = ( wire1581 ) | ( wire7116 ) | ( wire7117 ) ;
 assign wire731 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire730 = ( wire151 ) | ( (~ i_17_)  &  wire153 ) | ( (~ i_17_)  &  wire154 ) ;
 assign wire284 = ( (~ i_8_)  &  (~ i_31_) ) ;
 assign wire734 = ( wire345  &  wire735 ) | ( wire83  &  wire7686 ) ;
 assign wire66 = ( (~ i_31_)  &  n_n805  &  wire7547 ) ;
 assign wire502 = ( n_n1340  &  n_n1128  &  wire12 ) ;
 assign n_n1875 = ( wire1190 ) | ( wire1191 ) | ( wire7548 ) | ( wire7549 ) ;
 assign n_n1873 = ( wire1202 ) | ( wire1203 ) | ( wire7537 ) | ( wire7538 ) ;
 assign n_n1831 = ( n_n1875 ) | ( wire1184 ) | ( wire7554 ) | ( wire7570 ) ;
 assign n_n1816 = ( n_n1831 ) | ( n_n1877 ) | ( wire7596 ) | ( wire7598 ) ;
 assign wire739 = ( n_n1523  &  (~ n_n1251) ) | ( wire740  &  wire7639 ) ;
 assign n_n1818 = ( n_n1889 ) | ( n_n1837 ) | ( wire7622 ) | ( wire7642 ) ;
 assign n_n1834 = ( n_n1884 ) | ( wire1043 ) | ( wire7669 ) | ( wire7680 ) ;
 assign n_n1835 = ( n_n1887 ) | ( wire1002 ) | ( wire7705 ) | ( wire7708 ) ;
 assign wire744 = ( wire262 ) | ( wire436 ) | ( i_19_  &  wire18 ) ;
 assign wire745 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1884 = ( wire1053 ) | ( wire1054 ) | ( wire7661 ) ;
 assign wire457 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire262 = ( i_9_  &  (~ i_3_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire465 = ( n_n1433  &  n_n1466  &  wire12 ) ;
 assign wire510 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  wire71 ) ;
 assign wire755 = ( n_n394 ) | ( n_n391 ) | ( n_n315 ) | ( n_n317 ) ;
 assign wire82 = ( (~ i_27_)  &  i_25_  &  n_n1257  &  wire47 ) ;
 assign n_n1712 = ( wire1473 ) | ( wire1474 ) | ( wire7244 ) ;
 assign wire760 = ( wire249 ) | ( n_n1300  &  wire282 ) | ( n_n1300  &  wire1048 ) ;
 assign wire515 = ( n_n1307  &  n_n1263  &  n_n1144 ) ;
 assign wire768 = ( wire1634 ) | ( (~ i_0_)  &  wire1636 ) | ( (~ i_0_)  &  wire7057 ) ;
 assign wire771 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1877 = ( wire7587 ) | ( wire7588 ) | ( wire7591 ) ;
 assign wire784 = ( wire1338 ) | ( wire425  &  wire7399 ) | ( wire454  &  wire7399 ) ;
 assign wire788 = ( wire1069 ) | ( wire257  &  wire250 ) | ( wire257  &  wire206 ) ;
 assign wire792 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign n_n1887 = ( wire7699 ) | ( i_38_  &  wire1019 ) | ( i_38_  &  wire7696 ) ;
 assign wire353 = ( (~ i_9_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_18_) ) ;
 assign wire484 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  wire7145 ) ;
 assign wire489 = ( (~ i_9_)  &  (~ i_18_)  &  n_n787  &  wire7148 ) ;
 assign wire437 = ( i_10_  &  i_7_  &  i_3_  &  (~ i_18_) ) ;
 assign wire18 = ( i_9_  &  (~ i_3_)  &  (~ i_13_) ) | ( i_9_  &  (~ i_13_)  &  i_18_ ) ;
 assign wire435 = ( n_n1118  &  n_n1279  &  wire7428 ) ;
 assign wire422 = ( n_n1118  &  n_n1058  &  wire7415 ) ;
 assign wire434 = ( n_n1307  &  n_n1033  &  wire7050  &  wire7417 ) ;
 assign wire349 = ( (~ i_13_)  &  i_11_  &  i_18_  &  (~ i_22_) ) ;
 assign wire404 = ( (~ i_9_)  &  i_3_  &  (~ i_4_)  &  (~ i_2_) ) ;
 assign wire413 = ( (~ i_8_)  &  (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire37 = ( n_n1192  &  wire7342 ) | ( n_n1038  &  wire7343 ) ;
 assign wire44 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_29_ ) ;
 assign wire211 = ( (~ i_7_)  &  (~ i_32_) ) ;
 assign wire65 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1213  &  wire7053 ) ;
 assign wire436 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire803 = ( wire1663 ) | ( wire54  &  wire398 ) | ( wire54  &  wire1665 ) ;
 assign wire802 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire95 = ( i_30_  &  i_23_ ) | ( i_27_  &  i_32_ ) | ( i_23_  &  i_32_ ) ;
 assign wire96 = ( i_30_  &  i_27_ ) | ( i_30_  &  i_16_ ) | ( i_16_  &  i_32_ ) ;
 assign wire143 = ( i_30_  &  i_16_  &  i_34_ ) ;
 assign wire147 = ( (~ i_32_)  &  n_n1307  &  n_n1100  &  wire7178 ) ;
 assign wire202 = ( (~ i_8_)  &  n_n1213  &  wire7053 ) ;
 assign wire458 = ( (~ i_29_)  &  n_n1441  &  n_n1400 ) ;
 assign wire221 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_)  &  n_n1018 ) ;
 assign wire231 = ( wire404  &  wire7274 ) ;
 assign wire251 = ( n_n1441  &  wire77  &  wire7055 ) ;
 assign wire314 = ( n_n1369  &  n_n1100  &  n_n460 ) ;
 assign wire334 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_) ) ;
 assign wire338 = ( (~ i_5_)  &  i_3_  &  (~ i_4_)  &  (~ i_18_) ) ;
 assign wire343 = ( i_9_  &  (~ i_3_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire345 = ( i_14_  &  (~ i_28_)  &  i_13_  &  i_22_ ) ;
 assign wire356 = ( n_n1406  &  n_n461  &  n_n1213  &  wire7890 ) ;
 assign wire367 = ( n_n1443  &  n_n1307  &  n_n853 ) ;
 assign wire373 = ( (~ i_34_)  &  i_35_  &  n_n1375  &  n_n1322 ) ;
 assign wire384 = ( n_n1375  &  n_n1400  &  n_n301 ) ;
 assign wire402 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire406 = ( i_10_  &  wire1432 ) | ( i_10_  &  wire1433 ) | ( i_10_  &  wire1434 ) ;
 assign wire425 = ( (~ i_13_)  &  wire1342 ) | ( (~ i_13_)  &  wire1343 ) ;
 assign wire438 = ( (~ i_32_)  &  wire226  &  wire7576 ) ;
 assign wire454 = ( i_19_  &  wire1340 ) | ( i_19_  &  wire1341 ) ;
 assign wire495 = ( n_n1307  &  n_n1408  &  n_n839 ) ;
 assign wire498 = ( n_n787  &  n_n1118  &  n_n180  &  n_n179 ) ;
 assign wire517 = ( n_n1375  &  wire13  &  n_n1322  &  n_n820 ) ;
 assign wire521 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n841 ) ;
 assign wire522 = ( n_n1307  &  n_n841  &  n_n177  &  n_n178 ) ;
 assign wire526 = ( wire431  &  wire508 ) | ( wire274  &  wire7254 ) ;
 assign wire544 = ( n_n1443  &  wire437 ) | ( n_n1429  &  wire437 ) | ( n_n1429  &  wire891 ) ;
 assign wire557 = ( (~ i_9_)  &  i_7_  &  (~ i_14_) ) | ( (~ i_9_)  &  i_7_  &  (~ i_13_) ) ;
 assign wire582 = ( wire349 ) | ( (~ i_13_)  &  (~ i_22_)  &  wire7259 ) ;
 assign wire590 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire593 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire604 = ( n_n245  &  wire361 ) | ( n_n26  &  wire353 ) ;
 assign wire603 = ( n_n21  &  wire6892 ) | ( n_n18  &  wire6894 ) ;
 assign wire606 = ( n_n504  &  n_n1118 ) | ( n_n1278  &  wire6913 ) ;
 assign wire624 = ( n_n1307  &  wire361 ) | ( n_n787  &  wire353 ) ;
 assign wire635 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_) ) | ( (~ i_9_)  &  (~ i_6_)  &  i_13_ ) ;
 assign wire638 = ( wire1570 ) | ( n_n301  &  wire1572 ) | ( n_n301  &  wire1573 ) ;
 assign wire657 = ( n_n307 ) | ( n_n309 ) | ( wire1323 ) | ( wire1324 ) ;
 assign wire661 = ( i_7_  &  (~ i_14_)  &  (~ i_12_) ) | ( i_7_  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire666 = ( wire43  &  n_n1274 ) | ( (~ i_23_)  &  wire402 ) ;
 assign wire679 = ( i_12_  &  wire349 ) | ( n_n586  &  wire7473 ) ;
 assign wire683 = ( wire402 ) | ( wire1604 ) ;
 assign wire698 = ( wire221  &  wire367 ) | ( wire41  &  wire384 ) ;
 assign wire710 = ( n_n1307  &  n_n853  &  n_n1408 ) | ( n_n1307  &  n_n1408  &  n_n839 ) ;
 assign wire713 = ( n_n712  &  wire7898 ) | ( wire8021  &  wire8022 ) ;
 assign wire721 = ( n_n1318  &  n_n1118 ) | ( n_n1278  &  wire7217 ) ;
 assign wire735 = ( i_30_ ) | ( i_32_ ) ;
 assign wire741 = ( i_30_ ) | ( i_32_ ) | ( i_31_ ) ;
 assign wire740 = ( i_20_ ) | ( i_21_ ) ;
 assign wire759 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire758 = ( n_n1314  &  n_n1141 ) | ( n_n1322  &  wire7243 ) ;
 assign wire767 = ( (~ i_13_)  &  i_12_  &  i_11_ ) | ( (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire22 = ( wire1766  &  wire8085 ) | ( n_n129  &  n_n130  &  wire8085 ) ;
 assign wire34 = ( n_n1375  &  wire227  &  wire1767 ) | ( n_n1375  &  wire227  &  wire1768 ) ;
 assign wire101 = ( wire105  &  wire8090 ) | ( wire107  &  wire8090 ) ;
 assign wire102 = ( wire462  &  wire338  &  wire8091 ) ;
 assign wire105 = ( wire232  &  n_n178  &  wire8086 ) ;
 assign wire107 = ( n_n180  &  n_n1303  &  wire338 ) ;
 assign wire110 = ( n_n1429  &  n_n1326  &  wire6947 ) | ( n_n1408  &  n_n1326  &  wire6947 ) ;
 assign wire111 = ( n_n1396  &  n_n1404  &  n_n1374  &  n_n1375 ) ;
 assign wire117 = ( (~ i_28_)  &  n_n1438  &  wire6948  &  wire8065 ) ;
 assign wire118 = ( n_n1429  &  wire62 ) | ( wire62  &  wire8 ) ;
 assign wire119 = ( n_n1408  &  wire82 ) | ( n_n1408  &  wire121 ) ;
 assign wire120 = ( i_31_  &  i_34_  &  wire123 ) | ( i_31_  &  i_34_  &  wire125 ) ;
 assign wire121 = ( i_34_  &  i_33_  &  n_n1312  &  wire6996 ) ;
 assign wire123 = ( n_n1315  &  n_n1314  &  wire80 ) ;
 assign wire125 = ( wire80  &  n_n1323  &  n_n1322 ) ;
 assign wire129 = ( wire441  &  wire8056 ) | ( wire245  &  wire277  &  wire8056 ) ;
 assign wire130 = ( n_n1369  &  n_n1315  &  n_n1263  &  wire8057 ) ;
 assign wire133 = ( n_n1443  &  n_n1406  &  n_n1213  &  wire7491 ) ;
 assign wire134 = ( n_n1404  &  n_n1326  &  wire6947 ) ;
 assign wire142 = ( wire10  &  n_n793  &  n_n1315  &  wire7942 ) ;
 assign wire150 = ( n_n1397  &  n_n1092  &  n_n1406  &  n_n1408 ) ;
 assign wire151 = ( wire47  &  wire7058  &  wire8042 ) ;
 assign wire153 = ( n_n793  &  n_n1285  &  wire8043 ) ;
 assign wire154 = ( wire47  &  n_n1387  &  wire7058 ) ;
 assign wire158 = ( n_n1375  &  n_n1141  &  n_n1263  &  n_n820 ) ;
 assign wire160 = ( n_n1489  &  n_n1089  &  n_n1251  &  wire227 ) ;
 assign wire161 = ( n_n1429  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire163 = ( wire245  &  n_n984  &  n_n916  &  wire7828 ) ;
 assign wire164 = ( wire320  &  wire169 ) | ( n_n1443  &  wire320  &  wire713 ) ;
 assign wire166 = ( (~ i_14_)  &  wire265  &  wire202  &  wire8008 ) ;
 assign wire167 = ( (~ i_14_)  &  (~ i_16_)  &  wire295 ) ;
 assign wire169 = ( i_3_  &  (~ i_18_)  &  n_n1429  &  wire8022 ) ;
 assign wire172 = ( n_n1408  &  wire245  &  n_n984  &  wire7827 ) ;
 assign wire174 = ( i_36_  &  wire8007 ) | ( i_36_  &  n_n363  &  wire67 ) ;
 assign wire176 = ( (~ i_13_)  &  wire265  &  wire202  &  wire8008 ) ;
 assign wire177 = ( (~ i_13_)  &  (~ i_16_)  &  wire295 ) ;
 assign wire178 = ( n_n1404  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire183 = ( wire10  &  n_n1315  &  n_n1511  &  wire7802 ) ;
 assign wire184 = ( n_n1504  &  n_n1375  &  n_n1323  &  n_n1322 ) ;
 assign wire185 = ( n_n1216  &  n_n1092  &  wire687  &  wire7803 ) ;
 assign wire187 = ( n_n1504  &  n_n1315  &  n_n1314  &  n_n1375 ) ;
 assign wire189 = ( i_14_  &  (~ i_28_)  &  n_n1438  &  wire6948 ) ;
 assign wire190 = ( n_n1285  &  n_n1511  &  wire7997 ) ;
 assign wire191 = ( n_n1216  &  n_n1384  &  wire7999 ) ;
 assign wire192 = ( wire47  &  wire668  &  wire7058  &  wire7984 ) ;
 assign wire194 = ( n_n1504  &  n_n1375  &  n_n1285  &  n_n1322 ) ;
 assign wire195 = ( n_n880  &  n_n1459  &  wire200 ) | ( n_n880  &  n_n1459  &  wire201 ) ;
 assign wire197 = ( n_n1089  &  wire79  &  n_n1431  &  n_n1254 ) ;
 assign wire198 = ( n_n1504  &  n_n1315  &  n_n1375  &  n_n1263 ) ;
 assign wire200 = ( n_n1441  &  n_n1390  &  wire7105 ) ;
 assign wire201 = ( n_n1441  &  n_n1400  &  wire258 ) ;
 assign wire234 = ( n_n1216  &  n_n1374  &  n_n1387  &  wire7971 ) ;
 assign wire304 = ( n_n1147  &  wire79  &  n_n1431  &  n_n1254 ) ;
 assign wire336 = ( n_n1390  &  n_n1375  &  n_n1089  &  wire7787 ) ;
 assign wire339 = ( i_21_  &  n_n1425  &  wire340  &  wire6951 ) ;
 assign wire350 = ( n_n1216  &  n_n1141  &  n_n1263  &  wire7784 ) ;
 assign wire412 = ( (~ i_13_)  &  wire517 ) | ( (~ i_13_)  &  wire65  &  wire7961 ) ;
 assign wire417 = ( n_n1489  &  n_n1147  &  n_n1251  &  wire227 ) ;
 assign wire424 = ( wire43  &  n_n1258  &  wire227  &  wire7949 ) ;
 assign wire427 = ( n_n1390  &  wire86  &  wire7105  &  wire7940 ) ;
 assign wire439 = ( n_n1314  &  n_n1141  &  n_n820 ) ;
 assign wire451 = ( (~ i_14_)  &  wire517 ) | ( (~ i_14_)  &  wire65  &  wire7945 ) ;
 assign wire469 = ( wire10  &  n_n1258  &  wire227  &  wire7949 ) ;
 assign wire471 = ( n_n1443  &  n_n1397  &  n_n1092  &  n_n1406 ) ;
 assign wire494 = ( n_n1497  &  n_n1459  &  wire7930 ) ;
 assign wire497 = ( n_n1459  &  wire6982  &  wire7931 ) ;
 assign wire507 = ( n_n1396  &  wire546  &  wire6958 ) ;
 assign wire512 = ( n_n1406  &  wire8  &  wire7025 ) ;
 assign wire812 = ( (~ i_7_)  &  i_36_  &  wire464 ) | ( (~ i_7_)  &  i_36_  &  wire818 ) ;
 assign wire813 = ( n_n1489  &  wire340  &  wire452 ) ;
 assign wire818 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_31_)  &  wire214 ) ;
 assign wire825 = ( wire420  &  wire44  &  wire7749  &  wire7900 ) ;
 assign wire829 = ( n_n1369  &  n_n1128  &  wire515 ) ;
 assign wire833 = ( wire44  &  wire7749  &  wire7900  &  wire7901 ) ;
 assign wire834 = ( i_36_  &  wire7903 ) | ( i_36_  &  wire43  &  wire356 ) ;
 assign wire841 = ( (~ i_31_)  &  n_n1307  &  n_n1144  &  wire7887 ) ;
 assign wire843 = ( i_36_  &  wire7892 ) | ( i_36_  &  wire10  &  wire356 ) ;
 assign wire849 = ( (~ i_13_)  &  wire223  &  wire7878 ) ;
 assign wire850 = ( wire275  &  wire857 ) | ( i_21_  &  wire275  &  wire544 ) ;
 assign wire857 = ( i_21_  &  (~ i_19_)  &  n_n1443  &  n_n712 ) ;
 assign wire863 = ( wire265  &  wire868 ) | ( n_n195  &  wire265  &  wire67 ) ;
 assign wire864 = ( i_36_  &  wire7871 ) | ( i_36_  &  wire384  &  wire7868 ) ;
 assign wire868 = ( (~ i_14_)  &  n_n461  &  wire411  &  wire7819 ) ;
 assign wire875 = ( wire881  &  wire7862 ) | ( wire7858  &  wire7859  &  wire7862 ) ;
 assign wire877 = ( i_34_  &  i_36_  &  wire147 ) | ( i_34_  &  i_36_  &  wire878 ) ;
 assign wire878 = ( (~ i_14_)  &  wire80  &  n_n1322  &  wire261 ) ;
 assign wire881 = ( wire232  &  n_n1406  &  n_n1213  &  wire7860 ) ;
 assign wire884 = ( n_n1307  &  n_n841  &  wire458  &  wire7846 ) ;
 assign wire891 = ( i_10_  &  i_7_  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire903 = ( n_n461  &  wire411  &  wire7819  &  wire7820 ) ;
 assign wire904 = ( n_n1307  &  n_n841  &  wire458  &  wire7821 ) ;
 assign wire906 = ( n_n1375  &  n_n1213  &  wire910 ) | ( n_n1375  &  n_n1213  &  wire911 ) ;
 assign wire910 = ( n_n1307  &  n_n1408  &  n_n576  &  n_n839 ) ;
 assign wire911 = ( n_n1443  &  n_n1118  &  n_n1279  &  wire265 ) ;
 assign wire916 = ( n_n1404  &  wire82 ) | ( n_n1404  &  wire920 ) ;
 assign wire918 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_)  &  wire432 ) ;
 assign wire919 = ( n_n1390  &  n_n1472  &  n_n1147  &  wire7791 ) ;
 assign wire920 = ( i_34_  &  i_33_  &  n_n1312  &  wire6996 ) ;
 assign wire924 = ( n_n1438  &  n_n1326  &  wire7798 ) ;
 assign wire925 = ( n_n1216  &  wire13  &  wire260  &  wire7784 ) ;
 assign wire926 = ( (~ i_30_)  &  (~ i_28_)  &  wire245  &  wire340 ) ;
 assign wire928 = ( n_n1216  &  n_n1092  &  wire533  &  wire7803 ) ;
 assign wire933 = ( n_n1438  &  n_n1092  &  wire7782 ) ;
 assign wire935 = ( wire79  &  wire940 ) | ( wire79  &  wire941 ) ;
 assign wire937 = ( n_n1390  &  n_n1375  &  n_n1147  &  wire7787 ) ;
 assign wire939 = ( n_n1390  &  n_n1472  &  n_n1089  &  wire7791 ) ;
 assign wire940 = ( (~ i_7_)  &  (~ i_8_)  &  n_n1489  &  wire260 ) ;
 assign wire941 = ( n_n1489  &  n_n1141  &  n_n1263 ) ;
 assign wire942 = ( wire232  &  wire44  &  wire7749  &  wire7773 ) ;
 assign wire943 = ( wire498  &  wire7774 ) | ( wire522  &  wire7774 ) ;
 assign wire945 = ( n_n1443  &  wire948 ) | ( (~ i_10_)  &  n_n1443  &  wire455 ) ;
 assign wire948 = ( n_n576  &  wire484  &  wire7778 ) | ( n_n576  &  wire489  &  wire7778 ) ;
 assign wire950 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire953 = ( wire80  &  wire86  &  wire498 ) | ( wire80  &  wire86  &  wire522 ) ;
 assign wire955 = ( wire420  &  wire455 ) ;
 assign wire956 = ( wire484  &  wire7765 ) | ( wire489  &  wire7765 ) ;
 assign wire957 = ( n_n787  &  n_n180  &  n_n179  &  wire7766 ) ;
 assign wire958 = ( (~ i_13_)  &  wire223  &  wire373 ) ;
 assign wire959 = ( n_n1397  &  n_n301  &  n_n1258  &  wire272 ) ;
 assign wire960 = ( wire232  &  wire44  &  wire7749  &  wire7751 ) ;
 assign wire961 = ( i_36_  &  (~ i_35_)  &  wire463  &  wire547 ) ;
 assign wire965 = ( n_n177  &  n_n178  &  wire7757 ) ;
 assign wire966 = ( (~ i_14_)  &  wire261  &  wire373 ) ;
 assign wire967 = ( wire273  &  wire1766 ) | ( n_n129  &  n_n130  &  wire273 ) ;
 assign wire968 = ( n_n1397  &  n_n1258  &  n_n916  &  wire272 ) ;
 assign wire969 = ( i_3_  &  (~ i_18_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire977 = ( n_n1197  &  wire981 ) | ( n_n1197  &  wire335  &  wire7736 ) ;
 assign wire978 = ( (~ i_10_)  &  (~ i_31_)  &  n_n1307  &  n_n841 ) ;
 assign wire981 = ( n_n1486  &  n_n1118  &  n_n1279  &  n_n1359 ) ;
 assign wire983 = ( wire988  &  wire7724 ) | ( wire61  &  wire343  &  wire7724 ) ;
 assign wire987 = ( n_n805  &  n_n1466  &  n_n849 ) ;
 assign wire988 = ( wire349  &  wire7723 ) | ( wire7258  &  wire7259  &  wire7723 ) ;
 assign wire990 = ( n_n416  &  n_n1300  &  wire457 ) | ( n_n1300  &  n_n706  &  wire457 ) ;
 assign wire991 = ( (~ i_24_)  &  wire297  &  wire7716 ) | ( (~ i_24_)  &  wire1406  &  wire7716 ) ;
 assign wire992 = ( n_n805  &  wire994 ) | ( n_n805  &  n_n1302  &  n_n849 ) ;
 assign wire993 = ( wire66  &  wire996 ) | ( wire66  &  wire7718 ) ;
 assign wire994 = ( n_n1307  &  n_n1359  &  wire7050  &  wire7717 ) ;
 assign wire996 = ( (~ i_32_)  &  n_n1307  &  n_n839 ) ;
 assign wire999 = ( (~ i_33_)  &  i_38_  &  wire61  &  wire7701 ) ;
 assign wire1000 = ( n_n1497  &  n_n1459  &  wire7702 ) ;
 assign wire1002 = ( n_n1489  &  wire1007 ) | ( n_n1489  &  wire226  &  wire7704 ) ;
 assign wire1007 = ( (~ i_31_)  &  n_n1454  &  n_n1179 ) ;
 assign wire1008 = ( i_30_  &  i_12_  &  i_17_ ) | ( i_12_  &  i_17_  &  i_32_ ) ;
 assign wire1009 = ( i_30_  &  i_14_  &  i_13_ ) | ( i_14_  &  i_13_  &  i_32_ ) ;
 assign wire1010 = ( n_n1437  &  wire7308  &  wire7690 ) ;
 assign wire1011 = ( n_n1523  &  wire7266  &  wire7691 ) ;
 assign wire1012 = ( n_n1504  &  wire345 ) | ( n_n1504  &  wire1015 ) ;
 assign wire1014 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1489  &  n_n1059 ) ;
 assign wire1015 = ( (~ i_28_)  &  i_12_  &  i_17_  &  i_22_ ) ;
 assign wire1017 = ( n_n1423  &  n_n1422  &  n_n1459 ) ;
 assign wire1019 = ( (~ i_2_)  &  wire1020 ) | ( (~ i_2_)  &  wire1021 ) ;
 assign wire1020 = ( (~ i_7_)  &  (~ i_22_)  &  n_n1454  &  n_n1431 ) ;
 assign wire1021 = ( (~ i_7_)  &  (~ i_8_)  &  n_n1425  &  wire7276 ) ;
 assign wire1022 = ( (~ i_7_)  &  (~ i_28_)  &  n_n1472  &  wire429 ) ;
 assign wire1023 = ( n_n1489  &  wire428  &  n_n805  &  wire284 ) ;
 assign wire1024 = ( n_n1489  &  wire13  &  n_n1059 ) | ( n_n1489  &  wire13  &  wire429 ) ;
 assign wire1029 = ( wire226  &  wire61  &  wire7670 ) ;
 assign wire1030 = ( n_n1353  &  n_n1197  &  n_n1497  &  wire57 ) ;
 assign wire1032 = ( (~ wire3)  &  n_n1197  &  n_n1486  &  n_n1359 ) ;
 assign wire1033 = ( n_n1369  &  n_n1368  &  wire792  &  wire7033 ) ;
 assign wire1040 = ( n_n1305  &  wire250  &  n_n1497 ) | ( n_n1305  &  n_n1497  &  wire206 ) ;
 assign wire1041 = ( n_n1353  &  n_n1423  &  n_n805  &  wire57 ) ;
 assign wire1043 = ( i_9_  &  i_12_  &  wire760 ) ;
 assign wire1044 = ( wire430  &  wire519 ) ;
 assign wire1045 = ( (~ i_24_)  &  i_38_  &  wire72  &  wire71 ) ;
 assign wire1048 = ( (~ i_7_)  &  (~ i_8_)  &  n_n1425  &  wire205 ) ;
 assign wire1050 = ( n_n1454  &  n_n1361  &  n_n1345  &  wire7655 ) ;
 assign wire1051 = ( wire78  &  wire12  &  wire7657 ) ;
 assign wire1052 = ( n_n1369  &  n_n1368  &  wire745  &  wire7033 ) ;
 assign wire1053 = ( n_n1353  &  wire1055 ) | ( n_n1353  &  wire1056 ) ;
 assign wire1054 = ( n_n1359  &  wire1057 ) | ( n_n1359  &  wire1058 ) | ( n_n1359  &  wire1059 ) ;
 assign wire1055 = ( (~ i_30_)  &  n_n805  &  wire7547 ) ;
 assign wire1056 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1489 ) ;
 assign wire1057 = ( (~ i_35_)  &  i_38_  &  n_n1489  &  n_n1340 ) ;
 assign wire1058 = ( (~ i_35_)  &  i_38_  &  n_n1478  &  n_n1472 ) ;
 assign wire1059 = ( (~ i_30_)  &  (~ i_32_)  &  n_n805  &  n_n1466 ) ;
 assign wire1060 = ( n_n1425  &  n_n1179  &  wire7276  &  wire7644 ) ;
 assign wire1061 = ( wire1066  &  wire7646 ) | ( n_n1425  &  n_n1197  &  wire7646 ) ;
 assign wire1062 = ( n_n1278  &  n_n1279  &  wire7492  &  wire7647 ) ;
 assign wire1064 = ( (~ i_32_)  &  wire788 ) ;
 assign wire1066 = ( (~ i_30_)  &  (~ i_35_)  &  i_38_  &  n_n1478 ) ;
 assign wire1069 = ( n_n1278  &  n_n1279  &  n_n1523  &  wire7266 ) ;
 assign wire1070 = ( wire58  &  wire1077 ) | ( wire58  &  wire741  &  wire7638 ) ;
 assign wire1077 = ( i_12_  &  (~ i_24_)  &  i_17_  &  i_31_ ) ;
 assign wire1080 = ( n_n1497  &  wire35 ) | ( n_n1497  &  wire1082 ) | ( n_n1497  &  wire7636 ) ;
 assign wire1081 = ( i_23_  &  wire447 ) ;
 assign wire1082 = ( i_27_  &  i_31_ ) | ( i_23_  &  i_31_ ) | ( i_16_  &  i_31_ ) ;
 assign wire1086 = ( n_n1439  &  wire143 ) | ( n_n1439  &  wire1089 ) ;
 assign wire1087 = ( i_23_  &  wire1091 ) | ( i_23_  &  wire3  &  n_n1497 ) ;
 assign wire1089 = ( i_27_  &  i_31_  &  i_34_ ) | ( i_16_  &  i_31_  &  i_34_ ) ;
 assign wire1091 = ( (~ i_28_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire1095 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1504  &  (~ n_n1251) ) ;
 assign wire1097 = ( (~ i_24_)  &  wire1100 ) | ( (~ i_24_)  &  n_n1511  &  wire7629 ) ;
 assign wire1100 = ( (~ i_28_)  &  i_22_  &  wire143 ) | ( (~ i_28_)  &  i_22_  &  wire1101 ) ;
 assign wire1101 = ( i_14_  &  i_34_  &  i_33_ ) ;
 assign wire1105 = ( i_29_  &  wire61  &  wire615 ) ;
 assign wire1106 = ( i_21_  &  (~ i_22_)  &  wire372 ) ;
 assign wire1108 = ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire1111 = ( (~ i_28_)  &  i_31_  &  i_34_  &  (~ i_29_) ) ;
 assign wire1112 = ( (~ i_7_)  &  (~ i_28_)  &  n_n1472  &  wire7616 ) ;
 assign wire1113 = ( wire95  &  wire7618 ) | ( wire96  &  wire7618 ) ;
 assign wire1114 = ( n_n1519  &  wire7619 ) | ( wire1121  &  wire7619 ) ;
 assign wire1121 = ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire1123 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1504  &  wire585 ) ;
 assign wire1125 = ( i_34_  &  wire1128 ) | ( i_34_  &  wire1129 ) | ( i_34_  &  wire1130 ) ;
 assign wire1126 = ( (~ i_7_)  &  (~ i_8_)  &  n_n1489  &  n_n1300 ) ;
 assign wire1127 = ( i_30_  &  wire345 ) | ( i_32_  &  wire345 ) ;
 assign wire1128 = ( i_12_  &  (~ i_24_)  &  i_17_  &  wire7612 ) ;
 assign wire1129 = ( (~ i_24_)  &  i_38_  &  n_n1466  &  wire77 ) ;
 assign wire1130 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1489  &  wire239 ) ;
 assign wire1131 = ( (~ i_30_)  &  (~ i_29_)  &  n_n1478  &  wire7600 ) ;
 assign wire1132 = ( (~ i_24_)  &  i_38_  &  wire71  &  wire7602 ) ;
 assign wire1133 = ( (~ i_33_)  &  i_38_  &  n_n1486  &  wire7603 ) ;
 assign wire1134 = ( i_20_  &  (~ i_22_)  &  wire372 ) ;
 assign wire1135 = ( wire83  &  wire1137 ) | ( n_n1504  &  wire83  &  (~ n_n1251) ) ;
 assign wire1136 = ( (~ i_7_)  &  (~ i_32_)  &  n_n1489  &  wire503 ) ;
 assign wire1137 = ( i_14_  &  (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire1139 = ( n_n1307  &  n_n1144  &  wire1146 ) | ( n_n1307  &  n_n1144  &  wire1147 ) ;
 assign wire1140 = ( i_9_  &  i_12_  &  wire235 ) | ( i_9_  &  i_12_  &  wire1148 ) ;
 assign wire1141 = ( n_n1307  &  wire438  &  wire7050 ) | ( n_n1307  &  wire1150  &  wire7050 ) ;
 assign wire1142 = ( n_n1278  &  n_n1279  &  wire78  &  wire7492 ) ;
 assign wire1143 = ( n_n1406  &  n_n1213  &  wire8  &  wire7491 ) ;
 assign wire1146 = ( wire226  &  wire457 ) ;
 assign wire1147 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1128 ) ;
 assign wire1148 = ( n_n1438  &  n_n1197  &  wire61 ) ;
 assign wire1150 = ( n_n1478  &  n_n1133  &  wire12 ) ;
 assign wire1152 = ( n_n1353  &  wire78  &  wire12  &  wire7582 ) ;
 assign wire1156 = ( (~ i_24_)  &  wire223  &  wire380 ) | ( (~ i_24_)  &  wire380  &  wire261 ) ;
 assign wire1157 = ( n_n1307  &  wire502  &  wire7050 ) | ( n_n1307  &  wire465  &  wire7050 ) ;
 assign wire1159 = ( n_n1425  &  n_n1197  &  wire205  &  wire7572 ) ;
 assign wire1161 = ( n_n1118  &  n_n1279  &  wire226  &  wire457 ) ;
 assign wire1162 = ( wire224  &  n_n1279  &  wire438 ) | ( wire224  &  n_n1279  &  wire1164 ) ;
 assign wire1163 = ( i_9_  &  i_12_  &  wire1167 ) | ( i_9_  &  i_12_  &  wire7578 ) ;
 assign wire1164 = ( n_n1478  &  n_n1133  &  wire12 ) ;
 assign wire1167 = ( (~ i_10_)  &  wire1169 ) | ( (~ i_10_)  &  wire1170 ) ;
 assign wire1168 = ( n_n1425  &  n_n1361  &  wire284  &  wire7276 ) ;
 assign wire1169 = ( n_n1197  &  n_n1523  &  n_n1431 ) ;
 assign wire1170 = ( n_n1425  &  n_n1179  &  wire7276 ) ;
 assign wire1172 = ( wire1180  &  wire7559 ) | ( wire1181  &  wire7559 ) ;
 assign wire1173 = ( n_n1179  &  wire71  &  wire278  &  wire262 ) ;
 assign wire1176 = ( n_n1278  &  n_n1288  &  n_n1279  &  n_n1059 ) ;
 assign wire1180 = ( (~ i_24_)  &  wire71  &  wire436 ) ;
 assign wire1181 = ( n_n1486  &  n_n998  &  wire18 ) ;
 assign wire1184 = ( (~ i_29_)  &  wire1189 ) | ( (~ i_29_)  &  wire360  &  wire315 ) ;
 assign wire1186 = ( n_n1307  &  n_n1288  &  n_n1306 ) ;
 assign wire1187 = ( (~ i_12_)  &  wire42  &  n_n1307  &  n_n1303 ) ;
 assign wire1189 = ( (~ i_24_)  &  wire223  &  wire311 ) ;
 assign wire1190 = ( wire1197  &  wire7543 ) | ( n_n1028  &  wire7541  &  wire7543 ) ;
 assign wire1191 = ( (~ i_24_)  &  (~ i_29_)  &  wire261  &  wire311 ) ;
 assign wire1197 = ( (~ i_13_)  &  wire1198 ) | ( (~ i_13_)  &  wire1342 ) | ( (~ i_13_)  &  wire1343 ) ;
 assign wire1198 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  i_19_ ) ;
 assign wire1201 = ( n_n1278  &  n_n1279  &  n_n1059  &  wire7532 ) ;
 assign wire1202 = ( wire425  &  wire7534 ) | ( wire454  &  wire7534 ) ;
 assign wire1203 = ( (~ i_24_)  &  wire223  &  wire266  &  n_n1302 ) ;
 assign wire1208 = ( (~ i_24_)  &  wire266  &  n_n1302  &  wire261 ) ;
 assign wire1211 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_29_)  &  wire700 ) ;
 assign wire1212 = ( i_13_  &  wire286 ) ;
 assign wire1214 = ( i_38_  &  n_n1278  &  n_n1279  &  n_n1202 ) ;
 assign wire1215 = ( n_n1437  &  n_n1472  &  wire529  &  wire7308 ) ;
 assign wire1218 = ( (~ i_24_)  &  n_n1466  &  wire266  &  wire261 ) ;
 assign wire1227 = ( wire9  &  wire77  &  wire78  &  wire68 ) ;
 assign wire1230 = ( n_n1197  &  n_n1523  &  n_n1431  &  wire7488 ) ;
 assign wire1234 = ( n_n1406  &  n_n1213  &  wire539  &  wire7491 ) ;
 assign wire1235 = ( n_n1278  &  n_n1279  &  wire288  &  wire7492 ) ;
 assign wire1236 = ( (~ i_32_)  &  n_n1307  &  n_n1306 ) ;
 assign wire1238 = ( wire521  &  wire7479 ) | ( wire404  &  wire7274  &  wire7479 ) ;
 assign wire1239 = ( (~ i_11_)  &  (~ i_19_)  &  wire429  &  wire272 ) ;
 assign wire1240 = ( n_n1466  &  n_n416  &  n_n1419 ) | ( n_n1466  &  n_n1419  &  n_n706 ) ;
 assign wire1241 = ( (~ i_24_)  &  wire446  &  wire4  &  wire78 ) ;
 assign wire1242 = ( n_n394  &  wire254 ) | ( n_n391  &  wire254 ) ;
 assign wire1247 = ( wire1253  &  wire7474 ) | ( i_10_  &  wire679  &  wire7474 ) ;
 assign wire1249 = ( i_19_  &  n_n307  &  wire288  &  wire12 ) ;
 assign wire1253 = ( i_10_  &  i_12_  &  wire7258  &  wire7259 ) ;
 assign wire1256 = ( wire1260  &  wire7469 ) | ( n_n735  &  wire405  &  wire7469 ) ;
 assign wire1257 = ( n_n307  &  wire7470 ) | ( n_n309  &  wire7470 ) ;
 assign wire1258 = ( wire12  &  wire422  &  wire7431 ) | ( wire12  &  wire434  &  wire7431 ) ;
 assign wire1259 = ( n_n1055  &  n_n461  &  wire253  &  wire7411 ) ;
 assign wire1260 = ( i_10_  &  wire1263 ) | ( i_10_  &  (~ i_3_)  &  wire767 ) ;
 assign wire1263 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire1264 = ( wire1323  &  wire7465 ) | ( wire1324  &  wire7465 ) ;
 assign wire1265 = ( wire235  &  wire406 ) | ( n_n586  &  wire235  &  wire7271 ) ;
 assign wire1266 = ( wire288  &  wire12  &  wire422 ) | ( wire288  &  wire12  &  wire434 ) ;
 assign wire1267 = ( i_19_  &  wire288  &  n_n309  &  wire12 ) ;
 assign wire1268 = ( n_n307  &  wire7459 ) | ( n_n309  &  wire7459 ) ;
 assign wire1271 = ( wire71  &  wire12  &  wire422 ) | ( wire71  &  wire12  &  wire434 ) ;
 assign wire1274 = ( wire423  &  wire7456 ) | ( wire435  &  wire7456 ) | ( wire1277  &  wire7456 ) ;
 assign wire1277 = ( i_19_  &  wire1279 ) | ( i_19_  &  wire1280 ) ;
 assign wire1279 = ( n_n461  &  n_n1028  &  wire7411 ) ;
 assign wire1280 = ( n_n1118  &  n_n1048  &  n_n1279 ) ;
 assign wire1281 = ( wire349  &  wire7454 ) | ( wire7258  &  wire7259  &  wire7454 ) ;
 assign wire1283 = ( wire71  &  wire12  &  wire423 ) | ( wire71  &  wire12  &  wire435 ) ;
 assign wire1284 = ( wire521  &  wire7446 ) | ( wire404  &  wire7274  &  wire7446 ) ;
 assign wire1286 = ( n_n416  &  n_n1419  &  n_n1302 ) | ( n_n1419  &  n_n1302  &  n_n706 ) ;
 assign wire1288 = ( n_n1523  &  n_n1458  &  wire4  &  wire7448 ) ;
 assign wire1289 = ( (~ i_24_)  &  wire271  &  wire231 ) | ( (~ i_24_)  &  wire271  &  wire521 ) ;
 assign wire1290 = ( wire422  &  wire7443 ) | ( wire434  &  wire7443 ) | ( wire1293  &  wire7443 ) ;
 assign wire1291 = ( n_n394  &  wire381 ) | ( n_n391  &  wire381 ) | ( n_n317  &  wire381 ) ;
 assign wire1293 = ( i_19_  &  n_n307 ) | ( i_19_  &  n_n309 ) ;
 assign wire1296 = ( wire21  &  wire276 ) | ( i_19_  &  wire276  &  wire657 ) ;
 assign wire1303 = ( (~ i_28_)  &  n_n1197  &  n_n1523  &  wire674 ) ;
 assign wire1305 = ( wire78  &  wire12  &  wire423 ) | ( wire78  &  wire12  &  wire435 ) ;
 assign wire1308 = ( wire1323  &  wire7430 ) | ( wire1324  &  wire7430 ) ;
 assign wire1309 = ( wire12  &  wire423  &  wire7431 ) | ( wire12  &  wire435  &  wire7431 ) ;
 assign wire1314 = ( n_n294  &  wire253 ) | ( n_n371  &  wire253 ) | ( n_n284  &  wire253 ) ;
 assign wire1316 = ( wire288  &  wire12  &  wire423 ) | ( wire288  &  wire12  &  wire435 ) ;
 assign wire1317 = ( n_n372  &  wire75 ) | ( n_n294  &  wire75 ) | ( n_n371  &  wire75 ) ;
 assign wire1318 = ( wire53  &  wire422 ) | ( wire53  &  wire434 ) | ( wire53  &  wire1320 ) ;
 assign wire1319 = ( n_n338  &  wire1323 ) | ( n_n338  &  wire1324 ) ;
 assign wire1320 = ( i_19_  &  n_n307 ) | ( i_19_  &  n_n309 ) ;
 assign wire1323 = ( n_n461  &  n_n1028  &  wire7411 ) ;
 assign wire1324 = ( n_n1118  &  n_n1048  &  n_n1279 ) ;
 assign wire1325 = ( wire425  &  wire7402 ) | ( wire454  &  wire7402 ) ;
 assign wire1330 = ( n_n1489  &  n_n1422  &  n_n998  &  wire18 ) ;
 assign wire1337 = ( n_n1523  &  wire346  &  wire7266 ) ;
 assign wire1338 = ( wire239  &  n_n1422  &  wire262 ) | ( wire239  &  n_n1422  &  wire436 ) ;
 assign wire1340 = ( i_9_  &  (~ i_8_)  &  (~ i_13_)  &  i_18_ ) ;
 assign wire1341 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  (~ i_13_) ) ;
 assign wire1342 = ( i_9_  &  (~ i_8_)  &  i_11_  &  i_18_ ) ;
 assign wire1343 = ( i_9_  &  (~ i_8_)  &  (~ i_3_)  &  i_11_ ) ;
 assign wire1347 = ( n_n1197  &  wire7393 ) | ( n_n1197  &  n_n1486  &  n_n849 ) ;
 assign wire1349 = ( n_n1307  &  n_n841  &  n_n1128  &  wire7388 ) ;
 assign wire1350 = ( n_n1307  &  n_n1359  &  wire7050  &  wire7390 ) ;
 assign wire1351 = ( n_n1307  &  n_n853  &  n_n1133  &  n_n1497 ) ;
 assign wire1356 = ( wire377  &  wire7375 ) | ( (~ i_13_)  &  wire377  &  wire37 ) ;
 assign wire1357 = ( wire223  &  n_n1419  &  n_n1302 ) ;
 assign wire1367 = ( (~ i_24_)  &  wire297  &  wire7364 ) | ( (~ i_24_)  &  wire1406  &  wire7364 ) ;
 assign wire1372 = ( wire1379  &  wire7352 ) | ( (~ i_22_)  &  wire343  &  wire7352 ) ;
 assign wire1377 = ( (~ i_28_)  &  n_n1197  &  n_n1523  &  wire289 ) ;
 assign wire1379 = ( i_9_  &  wire349 ) | ( i_9_  &  wire7258  &  wire7259 ) ;
 assign wire1382 = ( n_n1466  &  wire223  &  n_n1419 ) | ( n_n1466  &  n_n1419  &  wire346 ) ;
 assign wire1383 = ( wire56  &  wire7344 ) | ( (~ i_13_)  &  wire56  &  wire37 ) ;
 assign wire1384 = ( n_n805  &  n_n1466  &  wire394 ) ;
 assign wire1392 = ( wire1397  &  wire7332 ) | ( n_n1439  &  n_n416  &  wire7332 ) ;
 assign wire1397 = ( (~ i_24_)  &  wire297  &  n_n1288 ) | ( (~ i_24_)  &  n_n1288  &  wire1406 ) ;
 assign wire1399 = ( n_n1423  &  n_n416  &  wire7317 ) | ( n_n1423  &  n_n706  &  wire7317 ) ;
 assign wire1403 = ( (~ i_32_)  &  wire1404 ) | ( (~ i_32_)  &  wire1405 ) ;
 assign wire1404 = ( (~ i_24_)  &  wire297  &  wire7324 ) | ( (~ i_24_)  &  wire1406  &  wire7324 ) ;
 assign wire1405 = ( wire297  &  n_n1300  &  wire61 ) | ( n_n1300  &  wire61  &  wire1426 ) ;
 assign wire1406 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n1100 ) ;
 assign wire1408 = ( (~ i_33_)  &  i_38_  &  wire1412 ) | ( (~ i_33_)  &  i_38_  &  wire1413 ) ;
 assign wire1409 = ( (~ i_24_)  &  wire446  &  wire4  &  wire71 ) ;
 assign wire1412 = ( n_n1425  &  wire1414 ) | ( n_n1425  &  wire1435 ) | ( n_n1425  &  wire1436 ) ;
 assign wire1413 = ( n_n1431  &  wire406  &  wire7272 ) ;
 assign wire1414 = ( wire205  &  wire1416  &  wire7297 ) | ( wire205  &  wire1417  &  wire7297 ) ;
 assign wire1416 = ( (~ i_13_)  &  i_12_  &  i_18_  &  i_19_ ) ;
 assign wire1417 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire1419 = ( wire297  &  n_n1419  &  wire344 ) | ( n_n1419  &  wire344  &  wire1426 ) ;
 assign wire1421 = ( n_n1128  &  wire1423 ) | ( n_n1128  &  wire624  &  wire7310 ) ;
 assign wire1423 = ( (~ i_24_)  &  wire231  &  wire7311 ) | ( (~ i_24_)  &  wire521  &  wire7311 ) ;
 assign wire1426 = ( (~ i_11_)  &  (~ i_19_)  &  n_n1307  &  n_n1100 ) ;
 assign wire1428 = ( i_10_  &  i_18_  &  n_n586  &  wire329 ) ;
 assign wire1429 = ( (~ i_24_)  &  wire231  &  wire7296 ) | ( (~ i_24_)  &  wire521  &  wire7296 ) ;
 assign wire1430 = ( (~ i_30_)  &  wire311  &  wire1435 ) | ( (~ i_30_)  &  wire311  &  wire1436 ) ;
 assign wire1431 = ( wire249  &  wire406 ) | ( n_n586  &  wire249  &  wire7271 ) ;
 assign wire1432 = ( (~ i_13_)  &  i_12_  &  i_18_  &  i_19_ ) ;
 assign wire1433 = ( (~ i_13_)  &  i_12_  &  i_11_  &  i_18_ ) ;
 assign wire1434 = ( (~ i_3_)  &  (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire1435 = ( (~ i_24_)  &  (~ i_22_)  &  wire7297  &  wire7298 ) ;
 assign wire1436 = ( i_10_  &  (~ i_3_)  &  n_n586  &  wire7299 ) ;
 assign wire1437 = ( wire1443  &  wire7285 ) | ( wire262  &  wire7284  &  wire7285 ) ;
 assign wire1439 = ( wire377  &  wire7288 ) | ( n_n1038  &  wire377  &  wire593 ) ;
 assign wire1443 = ( wire68  &  wire349 ) | ( wire68  &  wire7258  &  wire7259 ) ;
 assign wire1449 = ( (~ i_24_)  &  wire231  &  wire7275 ) | ( (~ i_24_)  &  wire521  &  wire7275 ) ;
 assign wire1450 = ( wire56  &  wire7281 ) | ( n_n1038  &  wire56  &  wire590 ) ;
 assign wire1456 = ( n_n762  &  wire1460 ) | ( n_n762  &  wire582  &  wire7261 ) ;
 assign wire1457 = ( i_38_  &  wire1461 ) | ( i_38_  &  n_n416  &  wire257 ) ;
 assign wire1460 = ( i_12_  &  wire61  &  wire262 ) ;
 assign wire1461 = ( n_n1454  &  wire1463  &  wire7264 ) | ( n_n1454  &  wire1464  &  wire7264 ) ;
 assign wire1463 = ( (~ i_18_)  &  (~ i_32_)  &  n_n1278  &  wire404 ) ;
 assign wire1464 = ( (~ i_32_)  &  wire204  &  n_n1307  &  n_n1100 ) ;
 assign wire1465 = ( wire59  &  wire1470 ) | ( wire59  &  wire526  &  wire7255 ) ;
 assign wire1470 = ( n_n245  &  n_n178  &  n_n18  &  wire6906 ) ;
 assign wire1473 = ( wire1477  &  wire7242 ) | ( wire260  &  wire77  &  wire7242 ) ;
 assign wire1474 = ( (~ i_33_)  &  wire1480 ) | ( (~ i_33_)  &  wire524  &  wire758 ) ;
 assign wire1476 = ( n_n1257  &  wire47  &  wire29  &  wire6998 ) ;
 assign wire1477 = ( (~ i_30_)  &  n_n1141  &  n_n1263 ) ;
 assign wire1480 = ( n_n1489  &  n_n1018  &  wire759  &  wire7108 ) ;
 assign wire1481 = ( wire44  &  wire6899  &  wire7224 ) ;
 assign wire1482 = ( wire224  &  n_n152  &  wire7214  &  wire7226 ) ;
 assign wire1483 = ( wire484  &  wire7228 ) | ( wire489  &  wire7228 ) ;
 assign wire1484 = ( wire498  &  wire7229 ) | ( wire522  &  wire7229 ) ;
 assign wire1485 = ( wire1576  &  wire7230 ) | ( wire1577  &  wire7230 ) ;
 assign wire1486 = ( n_n1216  &  wire351  &  wire6928 ) ;
 assign wire1490 = ( wire1507  &  wire7212 ) | ( wire1508  &  wire7212 ) ;
 assign wire1491 = ( wire224  &  n_n152  &  wire7214  &  wire7215 ) ;
 assign wire1492 = ( n_n1397  &  n_n1258  &  wire272  &  wire7216 ) ;
 assign wire1493 = ( n_n1408  &  wire1495 ) | ( n_n1408  &  wire721  &  wire7218 ) ;
 assign wire1495 = ( wire484  &  wire7219 ) | ( wire489  &  wire7219 ) ;
 assign wire1498 = ( n_n1278  &  wire404  &  wire7195 ) ;
 assign wire1499 = ( wire1507  &  wire7199 ) | ( wire1508  &  wire7199 ) ;
 assign wire1500 = ( wire365  &  wire1502 ) | ( wire365  &  wire1503 ) ;
 assign wire1501 = ( i_37_  &  wire1506 ) | ( i_37_  &  wire7205 ) ;
 assign wire1502 = ( n_n1408  &  n_n1422  &  wire484 ) | ( n_n1408  &  n_n1422  &  wire489 ) ;
 assign wire1503 = ( (~ i_14_)  &  n_n1397  &  n_n1322  &  wire261 ) ;
 assign wire1506 = ( n_n1397  &  n_n1258  &  n_n916  &  wire272 ) ;
 assign wire1507 = ( n_n1118  &  n_n179  &  wire404 ) ;
 assign wire1508 = ( n_n1307  &  n_n841  &  wire7197 ) ;
 assign wire1509 = ( wire1514  &  wire7187 ) | ( wire222  &  wire7185  &  wire7187 ) ;
 assign wire1511 = ( wire248  &  wire7191 ) | ( wire248  &  wire221  &  wire710 ) ;
 assign wire1514 = ( n_n1369  &  n_n460  &  wire6885  &  wire7186 ) ;
 assign wire1523 = ( n_n1307  &  n_n841  &  wire458  &  wire7176 ) ;
 assign wire1525 = ( n_n1295  &  wire1531 ) | ( n_n1295  &  wire1532 ) | ( n_n1295  &  wire7181 ) ;
 assign wire1531 = ( wire260  &  wire223  &  wire80 ) ;
 assign wire1532 = ( (~ i_14_)  &  wire80  &  n_n1322  &  wire261 ) ;
 assign wire1534 = ( wire1539  &  wire7160 ) | ( wire222  &  wire7158  &  wire7160 ) ;
 assign wire1535 = ( n_n1306  &  wire222  &  wire7161  &  wire7163 ) ;
 assign wire1539 = ( n_n1369  &  n_n460  &  wire6885  &  wire7159 ) ;
 assign wire1542 = ( n_n1278  &  n_n1279  &  wire259  &  wire7167 ) ;
 assign wire1546 = ( wire484  &  wire7151 ) | ( wire489  &  wire7151 ) ;
 assign wire1548 = ( wire482  &  wire498 ) | ( wire482  &  wire522 ) ;
 assign wire1549 = ( wire59  &  wire1550 ) | ( wire59  &  wire1551 ) | ( wire59  &  wire1552 ) ;
 assign wire1550 = ( n_n1278  &  n_n152  &  wire1553 ) | ( n_n1278  &  n_n152  &  wire1554 ) ;
 assign wire1551 = ( (~ i_13_)  &  wire223  &  wire373 ) ;
 assign wire1552 = ( n_n1397  &  n_n301  &  n_n1258  &  wire272 ) ;
 assign wire1553 = ( wire44  &  wire6899  &  wire7153 ) ;
 assign wire1554 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire259 ) ;
 assign wire1559 = ( wire317  &  wire1561 ) | ( n_n129  &  n_n130  &  wire317 ) ;
 assign wire1561 = ( n_n1278  &  n_n132  &  wire404  &  wire6882 ) ;
 assign wire1564 = ( n_n245  &  wire44  &  wire6899  &  wire7120 ) ;
 assign wire1565 = ( n_n1375  &  n_n1202  &  wire351 ) | ( n_n1375  &  n_n1202  &  wire1574 ) ;
 assign wire1566 = ( wire1576  &  wire7126 ) | ( wire1577  &  wire7126 ) ;
 assign wire1567 = ( n_n245  &  wire1568 ) | ( n_n1274  &  n_n245  &  wire638 ) ;
 assign wire1568 = ( (~ i_14_)  &  i_13_  &  i_37_  &  wire233 ) ;
 assign wire1570 = ( n_n1369  &  n_n1100  &  n_n460  &  wire7130 ) ;
 assign wire1572 = ( n_n1369  &  n_n1368  &  n_n841  &  n_n504 ) ;
 assign wire1573 = ( wire59  &  n_n1369  &  n_n1100  &  n_n460 ) ;
 assign wire1574 = ( n_n1278  &  n_n179  &  wire404  &  wire7123 ) ;
 assign wire1576 = ( (~ i_9_)  &  n_n1307  &  n_n1303  &  wire431 ) ;
 assign wire1577 = ( n_n1278  &  wire404  &  wire413 ) ;
 assign wire1580 = ( wire47  &  wire727  &  wire7058  &  wire7059 ) ;
 assign wire1581 = ( n_n1443  &  wire322 ) | ( n_n1443  &  wire1583 ) ;
 assign wire1582 = ( n_n1429  &  n_n1374  &  wire6996  &  wire6997 ) ;
 assign wire1583 = ( wire59  &  n_n1375  &  n_n1213  &  wire7006 ) ;
 assign wire1585 = ( n_n1390  &  n_n1375  &  wire7105 ) ;
 assign wire1586 = ( n_n1375  &  n_n1400  &  wire259 ) ;
 assign wire1587 = ( n_n504  &  wire57  &  wire1592 ) | ( n_n504  &  wire57  &  wire1593 ) ;
 assign wire1589 = ( n_n1080  &  wire694  &  wire7009 ) ;
 assign wire1591 = ( n_n1489  &  n_n1018  &  wire8  &  wire7108 ) ;
 assign wire1592 = ( n_n1441  &  n_n1390  &  wire7105 ) ;
 assign wire1593 = ( n_n1441  &  n_n1400  &  wire259 ) ;
 assign wire1597 = ( (~ i_0_)  &  wire1600 ) | ( (~ i_0_)  &  wire7099 ) ;
 assign wire1600 = ( wire59  &  wire1603 ) | ( wire59  &  wire65  &  wire683 ) ;
 assign wire1603 = ( n_n1441  &  n_n1443  &  wire77  &  wire7055 ) ;
 assign wire1604 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1607 = ( n_n1314  &  n_n1141  &  wire246  &  wire7080 ) ;
 assign wire1608 = ( wire1615  &  wire7084 ) | ( wire666  &  wire7082  &  wire7084 ) ;
 assign wire1611 = ( i_37_  &  n_n1018  &  n_n1225  &  n_n363 ) ;
 assign wire1615 = ( (~ i_8_)  &  n_n1213  &  wire7053  &  wire7083 ) ;
 assign wire1618 = ( n_n793  &  wire771  &  wire7063  &  wire7064 ) ;
 assign wire1619 = ( wire1623  &  wire7072 ) | ( wire1624  &  wire7072 ) | ( wire1625  &  wire7072 ) ;
 assign wire1622 = ( n_n1443  &  wire47  &  wire7058  &  wire7059 ) ;
 assign wire1623 = ( wire10  &  n_n1369  &  n_n1274  &  n_n1431 ) ;
 assign wire1624 = ( wire202  &  wire7069 ) | ( n_n1431  &  wire7068  &  wire7069 ) ;
 assign wire1625 = ( (~ i_8_)  &  n_n1213  &  wire7053  &  wire7070 ) ;
 assign wire1628 = ( n_n1375  &  n_n1322  &  wire246  &  wire7046 ) ;
 assign wire1632 = ( n_n1429  &  wire47  &  wire7058  &  wire7059 ) ;
 assign wire1634 = ( n_n1216  &  n_n620  &  wire6928 ) ;
 assign wire1635 = ( n_n1213  &  wire211  &  wire7053  &  wire7054 ) ;
 assign wire1636 = ( n_n1404  &  wire251 ) | ( n_n1404  &  wire1638 ) ;
 assign wire1637 = ( n_n1441  &  n_n1408  &  wire77  &  wire7055 ) ;
 assign wire1638 = ( (~ i_20_)  &  n_n1213  &  wire211  &  wire7053 ) ;
 assign wire1640 = ( n_n1334  &  n_n1375  &  n_n1400  &  n_n1401 ) ;
 assign wire1649 = ( i_25_  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_34_) ) ;
 assign wire1650 = ( i_25_  &  (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire1651 = ( n_n1396  &  n_n1374  &  n_n1375  &  n_n1408 ) ;
 assign wire1652 = ( n_n1443  &  n_n1326  &  wire6947 ) ;
 assign wire1653 = ( n_n1390  &  wire305  &  wire717 ) ;
 assign wire1654 = ( n_n1441  &  n_n1400  &  wire7031 ) ;
 assign wire1656 = ( n_n1406  &  wire8  &  wire7025 ) ;
 assign wire1657 = ( n_n1443  &  n_n1369  &  n_n1368  &  wire7033 ) ;
 assign wire1659 = ( n_n1441  &  n_n1400  &  wire7028 ) ;
 assign wire1661 = ( n_n1406  &  wire802  &  wire7025 ) ;
 assign wire1663 = ( (~ i_24_)  &  (~ i_34_)  &  n_n1425  &  wire7026 ) ;
 assign wire1665 = ( wire29  &  wire44 ) | ( wire44  &  wire7027 ) ;
 assign wire1668 = ( n_n1397  &  n_n1258  &  n_n1401  &  n_n1499 ) ;
 assign wire1669 = ( n_n1408  &  wire322 ) | ( n_n1408  &  wire82 ) ;
 assign wire1670 = ( i_20_  &  wire1675 ) | ( i_20_  &  wire1676 ) ;
 assign wire1672 = ( n_n1216  &  n_n1391  &  wire6959  &  wire7017 ) ;
 assign wire1675 = ( (~ i_28_)  &  i_25_  &  n_n1438  &  wire6948 ) ;
 assign wire1676 = ( n_n1216  &  wire1677  &  wire6959 ) | ( n_n1216  &  wire1678  &  wire6959 ) ;
 assign wire1677 = ( i_7_  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire1678 = ( i_7_  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire1682 = ( n_n1429  &  wire252 ) | ( n_n1429  &  n_n1080  &  wire7009 ) ;
 assign wire1683 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_)  &  wire432 ) ;
 assign wire1684 = ( n_n1443  &  n_n1080  &  wire7009 ) ;
 assign wire1685 = ( n_n1390  &  n_n1375  &  wire6993 ) ;
 assign wire1686 = ( n_n1375  &  n_n1400  &  wire258 ) ;
 assign wire1688 = ( n_n1499  &  wire1692 ) | ( n_n1499  &  wire1693 ) ;
 assign wire1689 = ( n_n1404  &  wire322 ) | ( n_n1404  &  wire82 ) ;
 assign wire1690 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_)  &  wire432 ) ;
 assign wire1691 = ( n_n1443  &  n_n1396  &  n_n1374  &  n_n1375 ) ;
 assign wire1692 = ( (~ i_34_)  &  i_35_  &  n_n1251  &  wire661 ) ;
 assign wire1693 = ( (~ i_34_)  &  i_35_  &  n_n1258  &  n_n1377 ) ;
 assign wire1694 = ( n_n1441  &  n_n1390  &  wire6993 ) ;
 assign wire1695 = ( n_n1441  &  n_n1400  &  wire258 ) ;
 assign wire1696 = ( n_n1318  &  n_n1497  &  n_n1311  &  n_n1459 ) ;
 assign wire1697 = ( i_21_  &  n_n1425  &  wire6951  &  wire6979 ) ;
 assign wire1698 = ( n_n1390  &  n_n1334  &  n_n1391  &  n_n1375 ) ;
 assign wire1699 = ( n_n1334  &  n_n1375  &  n_n1400  &  n_n1377 ) ;
 assign wire1700 = ( n_n1318  &  n_n1340  &  n_n1459  &  wire6982 ) ;
 assign wire1701 = ( n_n1433  &  wire54  &  n_n1489  &  wire416 ) ;
 assign wire1702 = ( n_n1433  &  n_n1312  &  wire6984 ) ;
 assign wire1703 = ( n_n1396  &  n_n1404  &  n_n1374  &  n_n1375 ) ;
 assign wire1704 = ( n_n1429  &  n_n1326  &  wire6947 ) ;
 assign wire1706 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire6955 ) ;
 assign wire1709 = ( n_n1406  &  n_n1408  &  wire245 ) ;
 assign wire1710 = ( n_n1216  &  n_n1401  &  wire6959  &  wire6960 ) ;
 assign wire1715 = ( wire302  &  n_n1489  &  wire452  &  wire416 ) ;
 assign wire1716 = ( wire1721  &  wire6971 ) | ( wire1722  &  wire6971 ) ;
 assign wire1717 = ( n_n1390  &  n_n1372  &  n_n1334  &  n_n1375 ) ;
 assign wire1718 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire6973 ) ;
 assign wire1719 = ( n_n1326  &  wire629  &  wire6947 ) ;
 assign wire1721 = ( (~ i_23_)  &  (~ i_24_)  &  n_n1489  &  wire6967 ) ;
 assign wire1722 = ( (~ i_14_)  &  (~ i_23_)  &  n_n1439  &  n_n1438 ) ;
 assign wire1726 = ( n_n1375  &  n_n1213  &  wire1730 ) | ( n_n1375  &  n_n1213  &  wire1731 ) ;
 assign wire1730 = ( n_n1307  &  n_n1408  &  wire635  &  wire6939 ) ;
 assign wire1731 = ( n_n1443  &  n_n504  &  n_n1118  &  n_n1279 ) ;
 assign wire1738 = ( n_n1429  &  n_n1307  &  n_n1303  &  wire317 ) ;
 assign wire1746 = ( n_n245  &  n_n18  &  wire6906  &  wire6908 ) ;
 assign wire1747 = ( n_n26  &  wire1748 ) | ( n_n26  &  wire1749 ) | ( n_n26  &  wire1750 ) ;
 assign wire1748 = ( wire1753  &  wire6912 ) | ( n_n21  &  wire6910  &  wire6912 ) ;
 assign wire1749 = ( n_n180  &  n_n21  &  wire606 ) ;
 assign wire1750 = ( n_n1369  &  n_n460  &  wire6885  &  wire6915 ) ;
 assign wire1753 = ( (~ i_14_)  &  wire413  &  wire44  &  wire6899 ) ;
 assign wire1756 = ( wire1766  &  wire6884 ) | ( n_n129  &  n_n130  &  wire6884 ) ;
 assign wire1757 = ( n_n1318  &  wire1759 ) | ( wire10  &  n_n1318  &  wire603 ) ;
 assign wire1758 = ( wire492  &  wire1767 ) | ( wire492  &  wire1768 ) ;
 assign wire1759 = ( wire604  &  wire6889 ) ;
 assign wire1766 = ( n_n1278  &  n_n132  &  wire404  &  wire6882 ) ;
 assign wire1767 = ( n_n1307  &  n_n1100  &  n_n177  &  n_n178 ) ;
 assign wire1768 = ( n_n1278  &  n_n787  &  n_n180  &  n_n179 ) ;
 assign wire6876 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_6_) ) ;
 assign wire6879 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire6880 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  wire6879 ) ;
 assign wire6881 = ( (~ i_11_)  &  (~ i_13_) ) ;
 assign wire6882 = ( (~ i_13_)  &  (~ i_8_) ) ;
 assign wire6884 = ( wire267  &  wire246 ) ;
 assign wire6885 = ( (~ i_23_)  &  (~ i_20_) ) ;
 assign wire6889 = ( n_n1369  &  n_n1408  &  n_n460  &  wire6885 ) ;
 assign wire6890 = ( (~ i_17_)  &  (~ i_18_) ) ;
 assign wire6891 = ( (~ i_9_)  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire6892 = ( i_3_  &  (~ i_4_)  &  (~ i_0_)  &  wire6891 ) ;
 assign wire6893 = ( (~ i_19_)  &  (~ i_17_) ) ;
 assign wire6894 = ( (~ i_11_)  &  n_n841  &  n_n245 ) ;
 assign wire6898 = ( wire1756 ) | ( wire1758 ) | ( wire233  &  wire6880 ) ;
 assign wire6899 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire6901 = ( (~ i_9_)  &  (~ i_14_)  &  i_37_  &  wire431 ) ;
 assign wire6903 = ( n_n841  &  n_n504  &  n_n245  &  n_n178 ) ;
 assign wire6905 = ( n_n1443  &  n_n504  &  n_n245  &  wire361 ) ;
 assign wire6906 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_32_) ) ;
 assign wire6908 = ( (~ i_14_)  &  (~ i_11_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire6910 = ( (~ i_14_)  &  (~ i_16_)  &  (~ i_32_) ) ;
 assign wire6912 = ( (~ i_9_)  &  i_37_  &  n_n1278 ) ;
 assign wire6913 = ( (~ i_32_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire6915 = ( n_n1443  &  n_n504  &  wire353 ) ;
 assign wire6917 = ( n_n18  &  wire6903 ) | ( wire63  &  wire6905 ) ;
 assign wire6919 = ( wire1746 ) | ( wire6917 ) | ( wire508  &  wire6901 ) ;
 assign wire6920 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire6922 = ( n_n1369  &  n_n504  &  n_n1288 ) ;
 assign wire6923 = ( (~ i_34_)  &  i_35_  &  (~ i_29_) ) ;
 assign wire6924 = ( i_37_  &  n_n793  &  wire6923 ) ;
 assign wire6926 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  wire365 ) ;
 assign wire6927 = ( i_34_  &  i_37_  &  n_n1216  &  n_n1305 ) ;
 assign wire6928 = ( (~ i_32_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire6930 = ( n_n329  &  wire6922 ) | ( n_n363  &  wire6924 ) ;
 assign wire6931 = ( n_n620  &  wire6926 ) | ( n_n269  &  wire6927 ) ;
 assign wire6933 = ( wire6931 ) | ( (~ i_35_)  &  i_37_  &  wire600 ) ;
 assign wire6934 = ( wire1738 ) | ( wire6930 ) | ( n_n1295  &  wire601 ) ;
 assign wire6935 = ( (~ i_35_)  &  i_37_  &  wire634 ) ;
 assign wire6936 = ( wire267  &  wire246 ) ;
 assign wire6937 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_)  &  n_n1018 ) ;
 assign wire6938 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_29_)  &  n_n1216 ) ;
 assign wire6939 = ( (~ i_32_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire6941 = ( n_n269  &  wire492 ) | ( n_n263  &  wire6936 ) ;
 assign wire6942 = ( wire6941 ) | ( wire41  &  wire458  &  wire6935 ) ;
 assign wire6943 = ( wire1726 ) | ( wire248  &  wire632 ) ;
 assign wire6947 = ( (~ i_27_)  &  (~ i_23_)  &  i_22_  &  i_35_ ) ;
 assign wire6948 = ( (~ i_34_)  &  i_33_  &  i_35_ ) ;
 assign wire6949 = ( (~ i_28_)  &  i_25_  &  (~ i_29_) ) ;
 assign wire6951 = ( (~ i_34_)  &  (~ i_24_) ) ;
 assign wire6952 = ( (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire6953 = ( i_25_  &  i_20_ ) ;
 assign wire6955 = ( (~ i_14_)  &  i_2_  &  (~ i_16_) ) ;
 assign wire6957 = ( (~ i_7_)  &  (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire6958 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_33_ ) ;
 assign wire6959 = ( (~ i_23_)  &  i_31_  &  i_34_ ) ;
 assign wire6960 = ( (~ i_17_)  &  i_20_ ) ;
 assign wire6961 = ( wire1710 ) | ( n_n1393  &  wire599  &  wire6953 ) ;
 assign wire6962 = ( wire1706 ) | ( n_n1438  &  wire597 ) ;
 assign wire6963 = ( wire1709 ) | ( n_n1429  &  wire598 ) ;
 assign wire6967 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_33_) ) ;
 assign wire6971 = ( (~ i_7_)  &  i_34_  &  i_37_ ) ;
 assign wire6973 = ( (~ i_13_)  &  i_2_  &  (~ i_16_) ) ;
 assign wire6977 = ( wire1718 ) | ( wire1719 ) | ( n_n1443  &  wire630 ) ;
 assign wire6979 = ( (~ i_32_)  &  (~ i_31_)  &  i_29_ ) ;
 assign wire6982 = ( (~ i_28_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire6984 = ( (~ i_30_)  &  (~ i_28_)  &  i_29_ ) ;
 assign wire6989 = ( wire1696 ) | ( wire1698 ) | ( wire1703 ) ;
 assign wire6990 = ( wire1699 ) | ( wire1700 ) | ( wire1702 ) | ( wire1704 ) ;
 assign wire6993 = ( (~ i_8_)  &  (~ i_14_)  &  (~ i_12_) ) ;
 assign wire6994 = ( (~ i_30_)  &  (~ i_35_)  &  (~ i_29_)  &  i_37_ ) ;
 assign wire6996 = ( (~ i_27_)  &  (~ i_28_)  &  i_25_ ) ;
 assign wire6997 = ( i_20_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire6998 = ( i_25_  &  (~ i_27_) ) ;
 assign wire7000 = ( (~ i_21_)  &  i_2_ ) ;
 assign wire7001 = ( wire1691 ) | ( wire1694  &  wire6994 ) | ( wire1695  &  wire6994 ) ;
 assign wire7004 = ( (~ i_30_)  &  i_34_  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7005 = ( (~ i_7_)  &  (~ i_8_)  &  wire260 ) ;
 assign wire7006 = ( (~ i_30_)  &  (~ i_32_)  &  i_31_ ) ;
 assign wire7007 = ( wire8  &  i_37_ ) ;
 assign wire7009 = ( (~ i_28_)  &  (~ i_34_)  &  i_35_  &  i_29_ ) ;
 assign wire7010 = ( wire524  &  wire7005 ) | ( wire306  &  wire7007 ) ;
 assign wire7011 = ( wire1684 ) | ( wire1685  &  wire7004 ) | ( wire1686  &  wire7004 ) ;
 assign wire7014 = ( (~ i_7_)  &  (~ i_14_)  &  (~ i_28_)  &  i_37_ ) ;
 assign wire7017 = ( (~ i_16_)  &  i_20_ ) ;
 assign wire7018 = ( wire1668 ) | ( n_n1202  &  n_n1459  &  wire7014 ) ;
 assign wire7019 = ( wire1672 ) | ( n_n1404  &  n_n1406  &  wire245 ) ;
 assign wire7022 = ( wire1669 ) | ( wire1670 ) | ( wire7018 ) | ( wire7019 ) ;
 assign wire7025 = ( (~ i_23_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire7026 = ( (~ i_32_)  &  (~ i_31_)  &  i_29_ ) ;
 assign wire7027 = ( (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) | ( (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7028 = ( i_7_  &  (~ i_13_)  &  (~ i_16_)  &  i_31_ ) ;
 assign wire7029 = ( (~ i_30_)  &  i_22_  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire7031 = ( i_7_  &  (~ i_14_)  &  (~ i_16_)  &  i_31_ ) ;
 assign wire7033 = ( (~ i_23_)  &  i_21_  &  (~ i_22_) ) ;
 assign wire7036 = ( wire1657 ) | ( n_n1396  &  wire716  &  wire6958 ) ;
 assign wire7037 = ( wire127 ) | ( wire1653 ) | ( wire1654 ) | ( wire1656 ) ;
 assign wire7040 = ( wire196 ) | ( n_n1429  &  wire55 ) | ( wire8  &  wire55 ) ;
 assign wire7041 = ( wire126 ) | ( wire1640 ) | ( wire1651 ) | ( wire1652 ) ;
 assign wire7043 = ( wire7036 ) | ( wire7037 ) | ( wire7040 ) | ( wire7041 ) ;
 assign wire7044 = ( n_n1718 ) | ( n_n1719 ) | ( n_n1720 ) | ( wire7043 ) ;
 assign wire7045 = ( n_n1716 ) | ( n_n1715 ) | ( n_n1723 ) | ( wire7022 ) ;
 assign wire7046 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire7050 = ( (~ i_12_)  &  (~ i_6_) ) ;
 assign wire7051 = ( (~ i_14_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign wire7052 = ( (~ i_32_)  &  i_34_  &  (~ i_35_)  &  wire365 ) ;
 assign wire7053 = ( (~ i_30_)  &  (~ i_27_)  &  (~ i_28_) ) ;
 assign wire7054 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7055 = ( (~ i_20_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7057 = ( wire1637 ) | ( wire1635 ) ;
 assign wire7058 = ( (~ i_27_)  &  (~ i_28_)  &  i_33_ ) ;
 assign wire7059 = ( i_25_  &  i_20_ ) ;
 assign wire7060 = ( wire1628 ) | ( wire80  &  wire248  &  wire515 ) ;
 assign wire7062 = ( wire1632 ) | ( wire7060 ) | ( n_n608  &  wire7052 ) ;
 assign wire7063 = ( (~ i_30_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire7064 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire7068 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7069 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire7070 = ( (~ i_20_)  &  (~ i_14_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7072 = ( (~ i_0_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7073 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1369  &  n_n1318 ) ;
 assign wire7074 = ( (~ i_35_)  &  i_37_  &  n_n1441  &  wire243 ) ;
 assign wire7075 = ( wire1618 ) | ( wire515  &  wire7073 ) ;
 assign wire7076 = ( wire1622 ) | ( n_n608  &  wire7074 ) ;
 assign wire7079 = ( n_n793  &  wire29  &  wire7063 ) ;
 assign wire7080 = ( (~ i_30_)  &  (~ i_27_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire7082 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_32_)  &  n_n1369 ) ;
 assign wire7083 = ( (~ i_20_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7084 = ( (~ i_0_)  &  (~ i_33_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7085 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1302 ) ;
 assign wire7086 = ( (~ i_13_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_16_) ) ;
 assign wire7087 = ( (~ i_35_)  &  i_37_  &  n_n1441  &  n_n1305 ) ;
 assign wire7089 = ( wire1607 ) | ( n_n571  &  n_n1311  &  wire7079 ) ;
 assign wire7090 = ( wire491  &  wire7085 ) | ( n_n544  &  wire7087 ) ;
 assign wire7093 = ( wire1608 ) | ( wire1611 ) | ( wire7089 ) | ( wire7090 ) ;
 assign wire7094 = ( wire1619 ) | ( wire7075 ) | ( wire7076 ) | ( wire7093 ) ;
 assign wire7095 = ( (~ i_35_)  &  i_37_  &  n_n1375  &  n_n1340 ) ;
 assign wire7096 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1288 ) ;
 assign wire7097 = ( (~ i_35_)  &  i_37_  &  n_n1375  &  n_n1213 ) ;
 assign wire7098 = ( (~ i_33_)  &  (~ i_35_)  &  i_37_  &  wire402 ) ;
 assign wire7099 = ( wire470  &  wire251 ) | ( wire202  &  wire7098 ) ;
 assign wire7102 = ( n_n544  &  wire7095 ) | ( n_n437  &  wire7096 ) ;
 assign wire7103 = ( wire491  &  wire482 ) | ( n_n195  &  wire7097 ) ;
 assign wire7104 = ( wire7103 ) | ( wire7102 ) ;
 assign wire7105 = ( (~ i_8_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire7108 = ( (~ i_32_)  &  i_31_  &  i_34_  &  i_37_ ) ;
 assign wire7110 = ( wire1589 ) | ( n_n984  &  wire47  &  wire693 ) ;
 assign wire7111 = ( wire1591 ) | ( n_n1141  &  n_n1263  &  wire524 ) ;
 assign wire7114 = ( (~ i_30_)  &  i_34_  &  n_n504 ) ;
 assign wire7115 = ( i_20_  &  n_n984  &  wire47 ) ;
 assign wire7116 = ( wire1580 ) | ( wire1677  &  wire7115 ) | ( wire1678  &  wire7115 ) ;
 assign wire7117 = ( wire1582 ) | ( wire1585  &  wire7114 ) | ( wire1586  &  wire7114 ) ;
 assign wire7119 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_6_)  &  (~ i_32_) ) ;
 assign wire7120 = ( n_n1443  &  n_n504  &  wire7119 ) ;
 assign wire7121 = ( (~ i_11_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign wire7123 = ( (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7126 = ( (~ i_14_)  &  i_37_  &  n_n793  &  wire6923 ) ;
 assign wire7130 = ( (~ i_14_)  &  i_13_  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7134 = ( (~ i_35_)  &  i_37_  &  n_n841  &  n_n245 ) ;
 assign wire7135 = ( n_n1369  &  n_n1274  &  n_n1368  &  wire663 ) ;
 assign wire7136 = ( (~ i_14_)  &  (~ i_16_)  &  n_n1274 ) ;
 assign wire7137 = ( i_37_  &  (~ i_10_) ) ;
 assign wire7139 = ( i_34_  &  i_37_  &  n_n1216  &  n_n1305 ) ;
 assign wire7140 = ( n_n1408  &  n_n839  &  wire6939 ) ;
 assign wire7141 = ( wire7134  &  wire7135 ) | ( wire88  &  wire7140 ) ;
 assign wire7142 = ( wire7141 ) | ( wire1767  &  wire7139 ) | ( wire1768  &  wire7139 ) ;
 assign wire7143 = ( wire1559 ) | ( n_n245  &  wire664  &  wire7137 ) ;
 assign wire7145 = ( (~ i_9_)  &  (~ i_6_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7148 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire7151 = ( n_n1443  &  n_n1375  &  n_n1318  &  n_n1340 ) ;
 assign wire7152 = ( n_n853  &  n_n1408  &  wire6939 ) ;
 assign wire7153 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_)  &  (~ i_32_) ) ;
 assign wire7157 = ( wire1546 ) | ( wire1548 ) | ( wire88  &  wire7152 ) ;
 assign wire7158 = ( (~ i_13_)  &  (~ i_16_)  &  n_n1144 ) ;
 assign wire7159 = ( (~ i_6_)  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire7160 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  n_n504 ) ;
 assign wire7161 = ( (~ i_5_)  &  (~ i_4_)  &  (~ i_0_)  &  (~ i_32_) ) ;
 assign wire7162 = ( (~ i_7_)  &  (~ i_6_)  &  (~ i_12_)  &  wire7161 ) ;
 assign wire7163 = ( (~ i_13_)  &  (~ i_16_)  &  (~ i_33_)  &  i_37_ ) ;
 assign wire7165 = ( (~ i_34_)  &  i_35_  &  n_n793  &  n_n1305 ) ;
 assign wire7166 = ( n_n1307  &  n_n1100  &  n_n1340 ) ;
 assign wire7167 = ( (~ i_34_)  &  i_35_  &  n_n1258  &  n_n1302 ) ;
 assign wire7169 = ( n_n458  &  wire7165 ) | ( wire384  &  wire7166 ) ;
 assign wire7172 = ( wire1534 ) | ( wire1535 ) | ( wire508  &  wire470 ) ;
 assign wire7173 = ( (~ i_32_)  &  (~ i_29_)  &  n_n793 ) ;
 assign wire7174 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1258 ) ;
 assign wire7175 = ( (~ i_34_)  &  i_35_  &  i_37_ ) ;
 assign wire7176 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_16_)  &  n_n504 ) ;
 assign wire7177 = ( n_n1375  &  n_n1458  &  n_n1213 ) ;
 assign wire7178 = ( n_n1375  &  n_n1400  &  n_n916 ) ;
 assign wire7179 = ( n_n1375  &  n_n1400  &  wire334 ) ;
 assign wire7181 = ( wire85  &  wire7178 ) | ( wire85  &  wire7179 ) ;
 assign wire7183 = ( wire1523 ) | ( wire705  &  wire7175 ) ;
 assign wire7185 = ( (~ i_14_)  &  (~ i_16_)  &  n_n1144 ) ;
 assign wire7186 = ( (~ i_6_)  &  (~ i_14_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire7187 = ( (~ i_35_)  &  i_37_  &  n_n245 ) ;
 assign wire7188 = ( i_34_  &  (~ i_33_)  &  i_37_ ) ;
 assign wire7189 = ( n_n1375  &  n_n1400  &  n_n916 ) ;
 assign wire7190 = ( n_n1375  &  n_n1400  &  wire334 ) ;
 assign wire7191 = ( n_n1307  &  n_n841  &  wire7189 ) | ( n_n1307  &  n_n841  &  wire7190 ) ;
 assign wire7192 = ( wire1509 ) | ( wire222  &  wire268  &  wire7162 ) ;
 assign wire7195 = ( n_n1216  &  n_n179  &  wire268  &  wire6928 ) ;
 assign wire7197 = ( (~ i_11_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_19_) ) ;
 assign wire7199 = ( (~ i_14_)  &  (~ i_16_)  &  wire80  &  wire248 ) ;
 assign wire7203 = ( n_n1278  &  n_n152  &  wire258 ) ;
 assign wire7204 = ( (~ i_14_)  &  n_n1397  &  n_n1375  &  n_n1322 ) ;
 assign wire7205 = ( wire319  &  wire7203 ) | ( wire223  &  wire7204 ) ;
 assign wire7208 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_24_)  &  i_37_ ) ;
 assign wire7210 = ( n_n1322  &  n_n1241  &  wire7208 ) ;
 assign wire7211 = ( (~ i_14_)  &  (~ i_28_)  &  (~ i_16_)  &  (~ i_29_) ) ;
 assign wire7212 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  wire7211 ) ;
 assign wire7214 = ( n_n1406  &  n_n1213  &  n_n629 ) ;
 assign wire7215 = ( (~ i_14_)  &  (~ i_32_)  &  (~ i_35_)  &  i_37_ ) ;
 assign wire7216 = ( (~ i_10_)  &  (~ i_14_)  &  (~ i_16_)  &  i_37_ ) ;
 assign wire7217 = ( i_37_  &  (~ i_32_) ) ;
 assign wire7218 = ( n_n152  &  wire44  &  wire6899 ) ;
 assign wire7219 = ( (~ i_35_)  &  i_37_  &  n_n1441  &  wire243 ) ;
 assign wire7221 = ( wire1492 ) | ( (~ i_13_)  &  wire223  &  wire7210 ) ;
 assign wire7224 = ( n_n1443  &  n_n504  &  n_n1118  &  n_n152 ) ;
 assign wire7226 = ( (~ i_13_)  &  i_37_  &  n_n1458 ) ;
 assign wire7228 = ( n_n1441  &  n_n1443  &  n_n1318  &  n_n1305 ) ;
 assign wire7229 = ( (~ i_35_)  &  i_37_  &  n_n1369  &  n_n1302 ) ;
 assign wire7230 = ( (~ i_14_)  &  i_37_  &  n_n1018  &  n_n1225 ) ;
 assign wire7234 = ( wire1481 ) | ( wire1482 ) | ( wire1483 ) | ( wire1486 ) ;
 assign wire7235 = ( wire1484 ) | ( wire1485 ) | ( wire7234 ) ;
 assign wire7238 = ( n_n1705 ) | ( wire1549 ) | ( wire7157 ) ;
 assign wire7239 = ( n_n1703 ) | ( n_n1704 ) | ( wire7142 ) | ( wire7143 ) ;
 assign wire7240 = ( n_n1697 ) | ( n_n1701 ) | ( n_n1702 ) | ( wire7235 ) ;
 assign wire7242 = ( (~ i_34_)  &  i_35_  &  wire365 ) ;
 assign wire7243 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_13_) ) ;
 assign wire7244 = ( wire1476 ) | ( wire59  &  n_n1429  &  wire306 ) ;
 assign wire7247 = ( wire6933 ) | ( wire6934 ) | ( wire6942 ) | ( wire6943 ) ;
 assign wire7248 = ( n_n1714 ) | ( n_n1713 ) | ( n_n1712 ) ;
 assign wire7250 = ( wire1597 ) | ( wire7104 ) | ( wire7247 ) | ( wire7248 ) ;
 assign wire7252 = ( n_n1690 ) | ( wire7238 ) | ( wire7239 ) | ( wire7240 ) ;
 assign wire7254 = ( n_n1278  &  n_n26  &  wire413 ) ;
 assign wire7255 = ( (~ i_13_)  &  (~ i_9_) ) ;
 assign wire7256 = ( wire1747 ) | ( wire1757 ) | ( wire6898 ) | ( wire6919 ) ;
 assign wire7257 = ( wire7256 ) | ( wire1465 ) ;
 assign wire7258 = ( (~ i_22_)  &  (~ i_13_) ) ;
 assign wire7259 = ( (~ i_3_)  &  i_19_ ) | ( i_18_  &  i_19_ ) ;
 assign wire7261 = ( i_9_  &  i_12_  &  n_n1497 ) ;
 assign wire7264 = ( (~ i_22_)  &  (~ i_28_) ) ;
 assign wire7265 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_) ) ;
 assign wire7266 = ( (~ i_28_)  &  (~ i_33_)  &  i_38_ ) ;
 assign wire7267 = ( wire1456 ) | ( n_n416  &  wire70 ) | ( wire70  &  n_n706 ) ;
 assign wire7268 = ( (~ i_26_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7269 = ( n_n1128  &  n_n1458  &  wire7268 ) ;
 assign wire7271 = ( (~ i_3_)  &  i_10_ ) ;
 assign wire7272 = ( (~ i_7_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire7273 = ( (~ i_33_)  &  i_38_  &  n_n586  &  wire7271 ) ;
 assign wire7274 = ( (~ i_8_)  &  (~ i_5_)  &  (~ i_6_)  &  (~ i_18_) ) ;
 assign wire7275 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_29_)  &  wire226 ) ;
 assign wire7276 = ( (~ i_25_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire7277 = ( i_9_  &  (~ i_8_)  &  i_12_ ) ;
 assign wire7281 = ( n_n584  &  n_n1033 ) | ( n_n735  &  wire7277 ) ;
 assign wire7282 = ( wire4  &  wire7269 ) | ( wire282  &  wire7273 ) ;
 assign wire7284 = ( (~ i_22_)  &  i_12_ ) ;
 assign wire7285 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  n_n1431 ) ;
 assign wire7286 = ( (~ i_24_)  &  (~ i_22_)  &  i_38_  &  wire7265 ) ;
 assign wire7288 = ( n_n584  &  n_n1033 ) | ( n_n735  &  wire7277 ) ;
 assign wire7290 = ( wire1437 ) | ( wire1439 ) | ( n_n706  &  wire7286 ) ;
 assign wire7295 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign wire7296 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_  &  wire7295 ) ;
 assign wire7297 = ( i_10_  &  (~ i_7_)  &  (~ i_8_) ) ;
 assign wire7298 = ( (~ i_3_)  &  (~ i_13_)  &  i_12_  &  i_19_ ) ;
 assign wire7299 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_24_)  &  (~ i_22_) ) ;
 assign wire7301 = ( (~ i_7_)  &  (~ i_32_)  &  i_38_ ) ;
 assign wire7306 = ( i_10_  &  i_19_  &  n_n584 ) ;
 assign wire7308 = ( (~ i_28_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7309 = ( n_n1437  &  n_n1133  &  wire7308 ) ;
 assign wire7310 = ( (~ i_32_)  &  i_34_  &  (~ i_35_)  &  wire239 ) ;
 assign wire7311 = ( i_34_  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7312 = ( wire329  &  wire7306 ) | ( wire4  &  wire7309 ) ;
 assign wire7316 = ( wire1408 ) | ( wire1419 ) | ( wire1421 ) | ( wire7312 ) ;
 assign wire7317 = ( i_34_  &  i_38_  &  (~ i_29_) ) ;
 assign wire7319 = ( i_9_  &  (~ i_10_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7320 = ( n_n1118  &  n_n1279  &  wire7319 ) ;
 assign wire7321 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  n_n1478 ) ;
 assign wire7322 = ( n_n819  &  n_n1279  &  n_n1191 ) ;
 assign wire7323 = ( (~ i_33_)  &  i_38_  &  wire447 ) ;
 assign wire7324 = ( i_34_  &  i_38_  &  n_n1466 ) ;
 assign wire7325 = ( wire52  &  wire7320 ) | ( wire7321  &  wire7322 ) ;
 assign wire7327 = ( wire1399 ) | ( wire7325 ) | ( n_n706  &  wire7323 ) ;
 assign wire7328 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7329 = ( wire58  &  n_n819  &  n_n1279  &  n_n1191 ) ;
 assign wire7330 = ( (~ i_31_)  &  (~ i_35_)  &  i_38_  &  n_n1478 ) ;
 assign wire7331 = ( n_n1307  &  n_n841  &  n_n1191 ) ;
 assign wire7332 = ( i_34_  &  (~ i_33_)  &  i_38_ ) ;
 assign wire7333 = ( i_9_  &  (~ i_10_)  &  n_n1118  &  n_n1279 ) ;
 assign wire7334 = ( (~ i_31_)  &  n_n1307  &  n_n839 ) ;
 assign wire7335 = ( wire7328  &  wire7329 ) | ( wire7330  &  wire7331 ) ;
 assign wire7336 = ( wire390  &  wire7333 ) | ( n_n300  &  wire7334 ) ;
 assign wire7337 = ( wire261  &  wire379 ) | ( wire276  &  wire289 ) ;
 assign wire7339 = ( wire7335 ) | ( wire7336 ) | ( wire7337 ) ;
 assign wire7340 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  wire7264 ) ;
 assign wire7341 = ( (~ i_31_)  &  n_n1307  &  n_n853 ) ;
 assign wire7342 = ( i_18_  &  i_11_ ) ;
 assign wire7343 = ( i_19_  &  (~ i_2_) ) ;
 assign wire7344 = ( wire283  &  wire343 ) | ( i_9_  &  wire283  &  n_n735 ) ;
 assign wire7345 = ( wire475  &  wire7340 ) | ( n_n300  &  wire7341 ) ;
 assign wire7348 = ( n_n1861 ) | ( wire1403 ) | ( wire7327 ) ;
 assign wire7349 = ( n_n1825 ) | ( wire1392 ) | ( wire7339 ) ;
 assign wire7350 = ( n_n1854 ) | ( wire1409 ) | ( wire7316 ) | ( wire7348 ) ;
 assign wire7351 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign wire7352 = ( (~ i_35_)  &  i_38_  &  n_n1454  &  wire7351 ) ;
 assign wire7353 = ( (~ i_10_)  &  n_n1466  &  n_n1419 ) ;
 assign wire7354 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1288 ) ;
 assign wire7355 = ( (~ i_32_)  &  (~ i_35_)  &  i_38_  &  wire78 ) ;
 assign wire7356 = ( (~ i_28_)  &  i_38_  &  (~ i_29_) ) ;
 assign wire7357 = ( wire85  &  wire7353 ) | ( wire335  &  wire7354 ) ;
 assign wire7358 = ( n_n706  &  wire456 ) | ( wire327  &  wire7355 ) ;
 assign wire7361 = ( (~ i_28_)  &  (~ i_26_)  &  n_n1191  &  wire226 ) ;
 assign wire7362 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1128 ) ;
 assign wire7363 = ( (~ i_28_)  &  (~ i_33_)  &  (~ i_29_)  &  n_n805 ) ;
 assign wire7364 = ( (~ i_32_)  &  (~ i_29_)  &  wire311 ) ;
 assign wire7365 = ( (~ i_31_)  &  n_n1307  &  n_n839 ) ;
 assign wire7366 = ( wire41  &  wire7361 ) | ( i_13_  &  wire41  &  wire7362 ) ;
 assign wire7367 = ( wire475  &  wire390 ) | ( wire394  &  wire7363 ) ;
 assign wire7368 = ( wire261  &  wire387 ) | ( n_n316  &  wire7365 ) ;
 assign wire7370 = ( wire7368 ) | ( n_n1454  &  n_n416  &  wire7356 ) ;
 assign wire7371 = ( wire1367 ) | ( wire7366 ) | ( wire7367 ) ;
 assign wire7372 = ( (~ i_25_)  &  (~ i_24_)  &  n_n805  &  n_n1128 ) ;
 assign wire7373 = ( n_n1307  &  n_n1133  &  n_n839 ) ;
 assign wire7374 = ( (~ i_31_)  &  n_n1307  &  n_n853 ) ;
 assign wire7375 = ( wire283  &  wire343 ) | ( i_9_  &  wire283  &  n_n735 ) ;
 assign wire7377 = ( (~ i_28_)  &  i_35_  &  i_38_  &  (~ i_29_) ) ;
 assign wire7379 = ( wire408  &  wire7372 ) | ( wire315  &  wire7373 ) ;
 assign wire7380 = ( i_13_  &  wire310 ) | ( n_n316  &  wire7374 ) ;
 assign wire7383 = ( wire1356 ) | ( wire1357 ) | ( wire7379 ) | ( wire7380 ) ;
 assign wire7385 = ( n_n1197  &  n_n1133  &  n_n1497 ) ;
 assign wire7386 = ( (~ i_35_)  &  i_38_  &  (~ i_29_)  &  n_n1478 ) ;
 assign wire7387 = ( n_n1307  &  n_n853  &  n_n1128 ) ;
 assign wire7388 = ( (~ i_10_)  &  (~ i_26_)  &  (~ i_24_) ) | ( i_13_  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire7390 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire7393 = ( wire1349 ) | ( wire1350 ) | ( wire1351 ) ;
 assign wire7394 = ( wire218  &  wire7385 ) | ( wire270  &  wire7387 ) ;
 assign wire7395 = ( wire327  &  wire510 ) | ( n_n849  &  wire7386 ) ;
 assign wire7397 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_)  &  wire311 ) ;
 assign wire7399 = ( (~ i_24_)  &  i_38_  &  n_n1437 ) ;
 assign wire7400 = ( wire388  &  wire261 ) | ( wire85  &  wire7397 ) ;
 assign wire7402 = ( (~ i_30_)  &  (~ i_24_)  &  n_n805  &  n_n1466 ) ;
 assign wire7406 = ( wire1325 ) | ( wire9  &  wire78  &  wire346 ) ;
 assign wire7407 = ( wire1347 ) | ( wire7394 ) | ( wire7395 ) | ( wire7406 ) ;
 assign wire7409 = ( (~ i_32_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire7411 = ( (~ i_3_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign wire7412 = ( i_9_  &  (~ i_13_)  &  i_19_ ) ;
 assign wire7413 = ( (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire7415 = ( (~ i_13_)  &  (~ i_4_)  &  (~ i_12_)  &  (~ i_2_) ) ;
 assign wire7417 = ( i_18_  &  (~ i_13_) ) ;
 assign wire7419 = ( (~ i_3_)  &  (~ i_13_)  &  (~ i_12_) ) ;
 assign wire7420 = ( i_9_  &  (~ i_8_)  &  (~ i_5_)  &  (~ i_6_) ) ;
 assign wire7423 = ( i_9_  &  (~ i_13_)  &  i_18_  &  i_19_ ) ;
 assign wire7424 = ( i_9_  &  (~ i_5_)  &  (~ i_6_)  &  i_19_ ) ;
 assign wire7425 = ( i_9_  &  (~ i_5_)  &  (~ i_6_)  &  i_11_ ) ;
 assign wire7426 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire7427 = ( i_9_  &  (~ i_8_)  &  (~ i_13_)  &  i_11_ ) ;
 assign wire7428 = ( i_9_  &  (~ i_13_)  &  i_11_  &  i_18_ ) ;
 assign wire7430 = ( (~ i_35_)  &  i_38_  &  n_n1225  &  n_n998 ) ;
 assign wire7431 = ( (~ i_28_)  &  (~ i_25_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire7432 = ( wire1308 ) | ( n_n284  &  wire75 ) ;
 assign wire7433 = ( wire1309 ) | ( n_n300  &  wire654 ) ;
 assign wire7435 = ( n_n1843 ) | ( wire1317 ) | ( wire1318 ) | ( wire1319 ) ;
 assign wire7437 = ( wire1305 ) | ( n_n300  &  wire675 ) ;
 assign wire7439 = ( wire53  &  wire423 ) | ( n_n316  &  wire656 ) ;
 assign wire7441 = ( wire1296 ) | ( wire1303 ) | ( wire7437 ) | ( wire7439 ) ;
 assign wire7443 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire430 ) ;
 assign wire7445 = ( wire1291 ) | ( n_n315  &  wire254 ) | ( n_n317  &  wire254 ) ;
 assign wire7446 = ( wire61  &  wire226 ) ;
 assign wire7447 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_)  &  wire429 ) ;
 assign wire7448 = ( i_38_  &  (~ i_28_) ) ;
 assign wire7452 = ( wire1284 ) | ( wire1286 ) | ( wire297  &  wire7447 ) ;
 assign wire7454 = ( n_n1438  &  n_n1197  &  n_n1497  &  wire405 ) ;
 assign wire7456 = ( (~ i_24_)  &  (~ i_35_)  &  i_38_  &  wire430 ) ;
 assign wire7457 = ( i_10_  &  (~ i_3_)  &  n_n1438  &  n_n586 ) ;
 assign wire7458 = ( wire381  &  wire671 ) | ( wire390  &  wire7457 ) ;
 assign wire7459 = ( (~ i_35_)  &  i_38_  &  n_n1486  &  n_n998 ) ;
 assign wire7461 = ( wire1268 ) | ( n_n315  &  wire381 ) ;
 assign wire7462 = ( wire1271 ) | ( wire254  &  wire676 ) ;
 assign wire7464 = ( n_n1847 ) | ( wire1274 ) | ( wire7458 ) ;
 assign wire7465 = ( (~ i_35_)  &  i_38_  &  n_n1486  &  n_n998 ) ;
 assign wire7466 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign wire7469 = ( n_n1425  &  n_n1361  &  wire284  &  wire7276 ) ;
 assign wire7470 = ( (~ i_35_)  &  i_38_  &  n_n1225  &  n_n998 ) ;
 assign wire7473 = ( (~ i_22_)  &  (~ i_3_) ) ;
 assign wire7474 = ( n_n1454  &  n_n1179  &  n_n1345 ) ;
 assign wire7477 = ( wire1247 ) | ( wire1249 ) | ( wire75  &  wire677 ) ;
 assign wire7479 = ( (~ i_28_)  &  (~ i_22_)  &  n_n1454  &  wire264 ) ;
 assign wire7483 = ( wire1238 ) | ( wire1239 ) | ( wire1241 ) | ( wire1242 ) ;
 assign wire7485 = ( wire1240 ) | ( wire1290 ) | ( wire7445 ) | ( wire7483 ) ;
 assign wire7487 = ( n_n1821 ) | ( wire7461 ) | ( wire7462 ) | ( wire7464 ) ;
 assign wire7488 = ( i_9_  &  (~ i_10_)  &  (~ i_2_) ) ;
 assign wire7491 = ( i_20_  &  (~ i_21_)  &  (~ i_22_) ) ;
 assign wire7492 = ( (~ i_8_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7493 = ( wire1230 ) | ( n_n1225  &  wire72  &  wire239 ) ;
 assign wire7494 = ( wire1234 ) | ( wire250  &  wire537 ) ;
 assign wire7495 = ( wire1235 ) | ( wire70  &  wire72 ) | ( wire70  &  wire1236 ) ;
 assign wire7500 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_)  &  n_n1454 ) ;
 assign wire7502 = ( wire212  &  wire691 ) | ( wire250  &  wire7500 ) ;
 assign wire7503 = ( wire1227 ) | ( wire206  &  wire692 ) ;
 assign wire7504 = ( wire124 ) | ( wire132 ) | ( wire288  &  wire519 ) ;
 assign wire7507 = ( (~ i_28_)  &  (~ i_26_)  &  n_n1300  &  n_n1191 ) ;
 assign wire7508 = ( n_n1454  &  wire224  &  n_n1279  &  wire7264 ) ;
 assign wire7510 = ( (~ i_24_)  &  (~ i_22_)  &  wire264  &  wire7265 ) ;
 assign wire7511 = ( wire85  &  wire7507 ) | ( wire446  &  wire7508 ) ;
 assign wire7512 = ( wire223  &  wire388 ) | ( wire50  &  wire7510 ) ;
 assign wire7516 = ( (~ i_10_)  &  i_34_  &  wire239 ) | ( i_13_  &  i_34_  &  wire239 ) ;
 assign wire7519 = ( (~ i_8_)  &  (~ i_25_)  &  wire214 ) ;
 assign wire7521 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire61 ) ;
 assign wire7522 = ( (~ i_31_)  &  n_n1118  &  n_n1279 ) ;
 assign wire7523 = ( (~ i_24_)  &  i_34_  &  i_38_ ) ;
 assign wire7525 = ( wire272  &  wire7516 ) | ( wire250  &  wire7519 ) ;
 assign wire7526 = ( n_n1149  &  wire7521 ) | ( wire53  &  wire7522 ) ;
 assign wire7529 = ( wire1208 ) | ( wire1212 ) | ( wire7525 ) | ( wire7526 ) ;
 assign wire7531 = ( (~ i_31_)  &  (~ i_29_)  &  n_n1118  &  n_n1279 ) ;
 assign wire7532 = ( (~ i_8_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire7534 = ( (~ i_30_)  &  (~ i_29_)  &  n_n1478  &  wire12 ) ;
 assign wire7536 = ( n_n1307  &  wire264  &  n_n1144 ) ;
 assign wire7537 = ( wire1201 ) | ( n_n1423  &  n_n805  &  wire7531 ) ;
 assign wire7538 = ( (~ i_10_)  &  wire286 ) | ( wire257  &  wire7536 ) ;
 assign wire7541 = ( i_19_  &  i_18_ ) ;
 assign wire7543 = ( (~ i_30_)  &  (~ i_24_)  &  n_n1197  &  n_n1486 ) ;
 assign wire7545 = ( (~ i_6_)  &  (~ i_12_)  &  n_n1307  &  wire61 ) ;
 assign wire7547 = ( (~ i_28_)  &  (~ i_24_)  &  (~ i_33_)  &  (~ i_29_) ) ;
 assign wire7548 = ( wire51  &  wire502 ) | ( n_n1149  &  wire7545 ) ;
 assign wire7549 = ( wire53  &  wire360 ) | ( wire50  &  wire66 ) ;
 assign wire7552 = ( n_n1489  &  n_n1458  &  wire7268 ) ;
 assign wire7553 = ( wire395  &  wire346 ) | ( wire744  &  wire7552 ) ;
 assign wire7554 = ( wire7553 ) | ( n_n1059  &  wire1186 ) | ( n_n1059  &  wire1187 ) ;
 assign wire7555 = ( i_38_  &  (~ i_25_) ) ;
 assign wire7559 = ( (~ i_30_)  &  (~ i_32_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7561 = ( n_n1454  &  n_n1307  &  wire7050  &  wire7264 ) ;
 assign wire7562 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  n_n1466 ) ;
 assign wire7565 = ( wire1173 ) | ( wire72  &  wire214  &  wire7555 ) ;
 assign wire7566 = ( wire446  &  wire7561 ) | ( wire206  &  wire7562 ) ;
 assign wire7567 = ( wire1176 ) | ( wire224  &  n_n1279  &  wire465 ) ;
 assign wire7570 = ( wire1172 ) | ( wire7565 ) | ( wire7566 ) | ( wire7567 ) ;
 assign wire7572 = ( i_9_  &  (~ i_10_)  &  (~ i_8_)  &  i_12_ ) ;
 assign wire7574 = ( wire503  &  (~ i_10_) ) ;
 assign wire7576 = ( (~ i_28_)  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_29_) ) ;
 assign wire7577 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_22_)  &  (~ i_31_) ) ;
 assign wire7578 = ( wire1168 ) | ( n_n1454  &  n_n1179  &  wire7577 ) ;
 assign wire7580 = ( wire1159 ) | ( wire1161 ) | ( wire272  &  wire7574 ) ;
 assign wire7582 = ( i_12_  &  (~ i_30_) ) ;
 assign wire7585 = ( (~ i_10_)  &  (~ i_32_)  &  n_n1307  &  n_n1100 ) ;
 assign wire7586 = ( n_n1118  &  n_n1279  &  n_n1128 ) ;
 assign wire7587 = ( wire1152 ) | ( i_13_  &  wire503  &  wire272 ) ;
 assign wire7588 = ( wire395  &  wire7585 ) | ( wire81  &  wire7586 ) ;
 assign wire7591 = ( wire1156 ) | ( wire1157 ) | ( wire76  &  wire66 ) ;
 assign wire7592 = ( wire1143 ) | ( wire1142 ) ;
 assign wire7595 = ( wire1139 ) | ( wire1140 ) | ( wire1141 ) | ( wire7592 ) ;
 assign wire7596 = ( wire1162 ) | ( wire1163 ) | ( wire7580 ) | ( wire7595 ) ;
 assign wire7598 = ( n_n1871 ) | ( n_n1873 ) | ( wire1211 ) | ( wire7529 ) ;
 assign wire7600 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_24_)  &  i_38_ ) ;
 assign wire7602 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign wire7603 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_24_) ) ;
 assign wire7609 = ( wire1131 ) | ( wire1133 ) | ( wire1134 ) | ( wire1136 ) ;
 assign wire7612 = ( i_30_  &  (~ i_28_)  &  i_22_ ) | ( (~ i_28_)  &  i_22_  &  i_32_ ) ;
 assign wire7615 = ( wire1123 ) | ( wire298  &  wire1126 ) | ( wire298  &  wire1127 ) ;
 assign wire7616 = ( (~ i_24_)  &  i_34_  &  (~ i_33_)  &  i_38_ ) ;
 assign wire7618 = ( (~ i_28_)  &  i_22_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire7619 = ( (~ i_28_)  &  i_22_  &  i_31_  &  i_34_ ) ;
 assign wire7621 = ( wire1112 ) | ( wire1113 ) | ( wire1114 ) ;
 assign wire7622 = ( wire1132 ) | ( wire1135 ) | ( wire7609 ) | ( wire7621 ) ;
 assign wire7626 = ( (~ i_28_)  &  (~ i_24_)  &  i_22_  &  i_34_ ) ;
 assign wire7627 = ( i_30_  &  (~ i_28_)  &  (~ i_26_) ) | ( (~ i_28_)  &  (~ i_26_)  &  i_32_ ) ;
 assign wire7629 = ( i_27_  &  i_22_ ) | ( i_16_  &  i_22_ ) ;
 assign wire7631 = ( wire35  &  wire7626 ) | ( n_n1519  &  wire7627 ) ;
 assign wire7632 = ( wire1095 ) | ( wire214  &  wire95 ) | ( wire214  &  wire96 ) ;
 assign wire7636 = ( i_30_  &  i_16_ ) | ( i_14_  &  i_33_ ) ;
 assign wire7638 = ( i_14_  &  i_13_  &  (~ i_24_) ) ;
 assign wire7639 = ( (~ i_24_)  &  (~ i_22_)  &  i_34_ ) ;
 assign wire7640 = ( wire1070 ) | ( (~ i_28_)  &  i_29_  &  wire739 ) ;
 assign wire7642 = ( n_n1896 ) | ( wire1080 ) | ( wire1081 ) | ( wire7640 ) ;
 assign wire7644 = ( i_9_  &  (~ i_10_)  &  (~ i_2_) ) ;
 assign wire7646 = ( (~ i_10_)  &  (~ i_24_)  &  (~ i_22_)  &  n_n1192 ) ;
 assign wire7647 = ( (~ i_28_)  &  (~ i_25_)  &  i_34_  &  (~ i_29_) ) ;
 assign wire7648 = ( (~ i_8_)  &  n_n1278  &  n_n1279 ) ;
 assign wire7651 = ( wire1060 ) | ( wire1062 ) | ( wire78  &  wire519 ) ;
 assign wire7652 = ( wire1061 ) | ( wire7651 ) | ( wire70  &  wire7648 ) ;
 assign wire7653 = ( i_14_  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire7655 = ( (~ i_8_)  &  (~ i_2_)  &  (~ i_22_) ) ;
 assign wire7657 = ( (~ i_30_)  &  (~ i_2_)  &  (~ i_32_)  &  (~ i_31_) ) ;
 assign wire7661 = ( wire1050 ) | ( wire1051 ) | ( wire1052 ) ;
 assign wire7666 = ( wire1041 ) | ( n_n1454  &  n_n1288  &  wire206 ) ;
 assign wire7669 = ( wire1040 ) | ( wire1044 ) | ( wire1045 ) | ( wire7666 ) ;
 assign wire7670 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign wire7673 = ( (~ i_2_)  &  (~ i_24_)  &  (~ i_22_)  &  n_n1425 ) ;
 assign wire7676 = ( wire1032 ) | ( n_n1374  &  n_n1375  &  wire38 ) ;
 assign wire7677 = ( wire1029 ) | ( (~ i_32_)  &  wire226  &  wire7673 ) ;
 assign wire7678 = ( wire128 ) | ( wire1030 ) | ( wire1033 ) ;
 assign wire7680 = ( wire7676 ) | ( wire7677 ) | ( wire7678 ) ;
 assign wire7682 = ( (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire7686 = ( i_30_  &  i_12_  &  i_17_ ) | ( i_12_  &  i_17_  &  i_32_ ) ;
 assign wire7689 = ( wire112 ) | ( wire1022 ) | ( n_n1397  &  wire734 ) ;
 assign wire7690 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_31_)  &  (~ i_29_) ) ;
 assign wire7691 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_8_)  &  (~ i_2_) ) ;
 assign wire7696 = ( wire1017 ) | ( n_n1439  &  n_n1438  &  n_n1437 ) ;
 assign wire7699 = ( wire1010 ) | ( wire1011 ) | ( wire1012 ) | ( wire1014 ) ;
 assign wire7701 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_2_)  &  (~ i_32_) ) ;
 assign wire7702 = ( (~ i_32_)  &  (~ i_33_)  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7703 = ( (~ i_30_)  &  (~ i_8_)  &  (~ i_31_) ) ;
 assign wire7704 = ( (~ i_8_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire7705 = ( wire1000 ) | ( wire214  &  wire1008 ) | ( wire214  &  wire1009 ) ;
 assign wire7706 = ( wire999 ) | ( wire71  &  wire12  &  wire7703 ) ;
 assign wire7708 = ( wire1023 ) | ( wire1024 ) | ( wire7689 ) | ( wire7706 ) ;
 assign wire7711 = ( n_n1881 ) | ( n_n1882 ) | ( wire1064 ) | ( wire7652 ) ;
 assign wire7714 = ( n_n1818 ) | ( n_n1834 ) | ( n_n1835 ) | ( wire7711 ) ;
 assign wire7716 = ( (~ i_32_)  &  (~ i_33_)  &  i_38_  &  n_n1486 ) ;
 assign wire7717 = ( (~ i_28_)  &  (~ i_25_)  &  (~ i_32_)  &  (~ i_29_) ) ;
 assign wire7718 = ( (~ i_10_)  &  n_n1307  &  n_n841 ) | ( i_13_  &  n_n1307  &  n_n841 ) ;
 assign wire7721 = ( (~ i_24_)  &  i_34_  &  (~ i_35_)  &  i_38_ ) ;
 assign wire7722 = ( wire7721  &  wire344 ) ;
 assign wire7723 = ( i_9_  &  (~ i_28_)  &  (~ i_26_)  &  (~ i_24_) ) ;
 assign wire7724 = ( (~ i_30_)  &  (~ i_2_)  &  (~ i_32_)  &  n_n1197 ) ;
 assign wire7725 = ( n_n1307  &  n_n853  &  n_n1133 ) ;
 assign wire7726 = ( i_9_  &  (~ i_10_)  &  n_n1307  &  wire7050 ) ;
 assign wire7727 = ( wire335  &  wire7722 ) | ( wire315  &  wire7725 ) ;
 assign wire7728 = ( (~ i_10_)  &  wire310 ) | ( n_n316  &  wire7726 ) ;
 assign wire7731 = ( (~ i_10_)  &  (~ i_24_)  &  n_n819  &  n_n1279 ) ;
 assign wire7732 = ( (~ i_35_)  &  i_38_  &  (~ i_29_)  &  n_n1478 ) ;
 assign wire7733 = ( i_34_  &  (~ i_35_)  &  i_38_  &  wire344 ) ;
 assign wire7734 = ( n_n1307  &  n_n1128  &  n_n839 ) ;
 assign wire7735 = ( (~ i_32_)  &  n_n1307  &  n_n853 ) ;
 assign wire7736 = ( (~ i_26_)  &  (~ i_24_)  &  n_n1288 ) ;
 assign wire7737 = ( wire394  &  wire7732 ) | ( wire327  &  wire7733 ) ;
 assign wire7738 = ( wire510  &  wire7731 ) | ( wire270  &  wire7734 ) ;
 assign wire7740 = ( wire977 ) | ( wire330  &  wire289 ) | ( wire330  &  wire978 ) ;
 assign wire7741 = ( wire7737 ) | ( wire7738 ) | ( wire66  &  wire7735 ) ;
 assign wire7743 = ( n_n1866 ) | ( n_n1865 ) | ( wire7740 ) | ( wire7741 ) ;
 assign wire7744 = ( wire7743 ) | ( n_n1827 ) ;
 assign wire7746 = ( n_n1852 ) | ( wire7485 ) | ( wire7487 ) | ( wire7744 ) ;
 assign wire7747 = ( n_n1829 ) | ( n_n1812 ) | ( wire7349 ) | ( wire7350 ) ;
 assign wire7749 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire7750 = ( (~ i_13_)  &  (~ i_32_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7751 = ( wire431  &  wire7750 ) | ( wire969  &  wire7750 ) ;
 assign wire7753 = ( (~ i_8_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire7757 = ( n_n1216  &  n_n1307  &  n_n1100  &  wire6928 ) ;
 assign wire7761 = ( (~ i_7_)  &  (~ i_8_)  &  i_36_ ) ;
 assign wire7763 = ( (~ i_14_)  &  i_13_  &  (~ i_16_)  &  wire232 ) ;
 assign wire7765 = ( n_n1443  &  n_n1375  &  n_n1422 ) ;
 assign wire7766 = ( n_n1216  &  n_n1278  &  wire6928 ) ;
 assign wire7769 = ( (~ i_7_)  &  (~ i_32_)  &  i_36_ ) ;
 assign wire7771 = ( wire953 ) | ( wire955 ) | ( wire363  &  wire7763 ) ;
 assign wire7772 = ( (~ i_8_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7773 = ( wire420  &  wire7772 ) | ( wire950  &  wire7772 ) ;
 assign wire7774 = ( (~ i_28_)  &  (~ i_29_)  &  n_n1369  &  n_n880 ) ;
 assign wire7776 = ( (~ i_14_)  &  i_13_  &  n_n825 ) ;
 assign wire7777 = ( n_n1406  &  n_n1213  &  n_n576 ) ;
 assign wire7778 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  (~ i_29_) ) ;
 assign wire7781 = ( wire942 ) | ( wire943 ) | ( wire232  &  wire568 ) ;
 assign wire7782 = ( (~ i_28_)  &  (~ i_24_)  &  i_34_  &  i_29_ ) ;
 assign wire7784 = ( (~ i_30_)  &  i_34_  &  i_36_  &  (~ i_29_) ) ;
 assign wire7785 = ( i_36_  &  (~ i_7_) ) ;
 assign wire7787 = ( (~ i_30_)  &  (~ i_32_)  &  i_34_  &  i_36_ ) ;
 assign wire7789 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_32_) ) ;
 assign wire7791 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_36_ ) ;
 assign wire7793 = ( wire933 ) | ( n_n1216  &  wire530  &  wire7784 ) ;
 assign wire7794 = ( wire937 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire516 ) ;
 assign wire7795 = ( wire939 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire410 ) ;
 assign wire7798 = ( i_20_  &  (~ i_26_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire7802 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  i_21_ ) ;
 assign wire7803 = ( i_29_  &  i_34_ ) ;
 assign wire7806 = ( wire926 ) | ( wire532  &  n_n1511  &  wire7802 ) ;
 assign wire7807 = ( wire928 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire410 ) ;
 assign wire7808 = ( wire924 ) | ( wire925 ) | ( n_n1404  &  wire432 ) ;
 assign wire7810 = ( i_31_  &  i_34_  &  wire80 ) ;
 assign wire7811 = ( (~ i_30_)  &  (~ i_28_)  &  (~ i_29_)  &  wire79 ) ;
 assign wire7812 = ( wire535  &  wire7810 ) | ( wire536  &  wire7811 ) ;
 assign wire7813 = ( wire919 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire516 ) ;
 assign wire7817 = ( (~ i_9_)  &  i_2_  &  wire578 ) ;
 assign wire7819 = ( (~ i_28_)  &  i_29_  &  n_n1369  &  n_n1254 ) ;
 assign wire7820 = ( (~ i_13_)  &  (~ i_31_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7821 = ( i_36_  &  (~ i_35_)  &  n_n916 ) ;
 assign wire7822 = ( (~ i_28_)  &  (~ i_23_)  &  (~ i_17_)  &  (~ i_21_) ) ;
 assign wire7823 = ( n_n355  &  wire418 ) | ( wire463  &  wire7817 ) ;
 assign wire7825 = ( wire7823 ) | ( wire86  &  wire576 ) ;
 assign wire7826 = ( wire903 ) | ( wire904 ) | ( wire906 ) ;
 assign wire7827 = ( i_10_  &  i_7_  &  i_13_ ) ;
 assign wire7828 = ( i_10_  &  i_7_  &  (~ i_12_) ) ;
 assign wire7829 = ( (~ i_28_)  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire7830 = ( (~ i_27_)  &  (~ i_23_)  &  i_21_  &  wire7829 ) ;
 assign wire7831 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_21_) ) ;
 assign wire7832 = ( (~ i_32_)  &  i_36_  &  n_n1441  &  wire7831 ) ;
 assign wire7834 = ( n_n1429  &  n_n1216  &  wire6959 ) ;
 assign wire7835 = ( i_36_  &  n_n793  &  wire6923 ) ;
 assign wire7836 = ( wire644  &  wire7830 ) | ( n_n458  &  wire7832 ) ;
 assign wire7837 = ( wire440  &  wire7834 ) | ( n_n363  &  wire7835 ) ;
 assign wire7838 = ( wire493  &  n_n620 ) | ( n_n242  &  wire418 ) ;
 assign wire7839 = ( wire7837 ) | ( wire7836 ) ;
 assign wire7840 = ( wire7838 ) | ( i_34_  &  i_36_  &  wire643 ) ;
 assign wire7842 = ( (~ i_27_)  &  (~ i_28_)  &  i_31_  &  (~ i_29_) ) ;
 assign wire7843 = ( (~ i_23_)  &  (~ i_34_)  &  i_35_  &  wire541 ) ;
 assign wire7844 = ( wire437  &  wire7842 ) | ( wire891  &  wire7842 ) ;
 assign wire7845 = ( (~ i_32_)  &  i_36_  &  n_n1441  &  wire7831 ) ;
 assign wire7846 = ( i_36_  &  (~ i_35_)  &  n_n301 ) ;
 assign wire7847 = ( (~ i_5_)  &  (~ i_6_)  &  (~ i_4_)  &  (~ i_31_) ) ;
 assign wire7849 = ( wire7843  &  wire7844 ) | ( n_n358  &  wire7845 ) ;
 assign wire7851 = ( wire7849 ) | ( n_n576  &  wire540 ) ;
 assign wire7852 = ( wire884 ) | ( wire7851 ) | ( n_n1429  &  wire307 ) ;
 assign wire7853 = ( wire7825 ) | ( wire7826 ) | ( wire7839 ) | ( wire7840 ) ;
 assign wire7854 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_)  &  i_36_ ) ;
 assign wire7855 = ( wire7854  &  wire214 ) ;
 assign wire7856 = ( n_n1441  &  wire265  &  wire7831 ) ;
 assign wire7857 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_31_) ) ;
 assign wire7858 = ( (~ i_14_)  &  n_n1213 ) | ( (~ i_13_)  &  n_n1213 ) ;
 assign wire7859 = ( (~ i_5_)  &  (~ i_6_)  &  n_n1279  &  wire7857 ) ;
 assign wire7860 = ( (~ i_13_)  &  (~ i_10_) ) ;
 assign wire7862 = ( (~ i_32_)  &  i_36_  &  (~ i_35_)  &  n_n825 ) ;
 assign wire7863 = ( wire267  &  wire227 ) ;
 assign wire7864 = ( n_n355  &  wire7855 ) | ( n_n358  &  wire7863 ) ;
 assign wire7866 = ( wire875 ) | ( wire7864 ) | ( wire559  &  wire7856 ) ;
 assign wire7867 = ( n_n1369  &  n_n1128  &  n_n576 ) ;
 assign wire7868 = ( (~ i_32_)  &  i_34_  &  n_n1307  &  n_n1100 ) ;
 assign wire7869 = ( (~ i_32_)  &  (~ i_34_)  &  i_35_  &  wire267 ) ;
 assign wire7870 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_17_)  &  wire214 ) ;
 assign wire7871 = ( n_n458  &  wire7869 ) | ( n_n242  &  wire7870 ) ;
 assign wire7874 = ( wire500  &  wire312 ) | ( n_n437  &  wire7867 ) ;
 assign wire7875 = ( n_n1404  &  wire307 ) | ( wire483  &  n_n329 ) ;
 assign wire7878 = ( i_34_  &  i_36_  &  wire80  &  n_n1322 ) ;
 assign wire7879 = ( n_n437  &  wire483 ) | ( n_n195  &  wire500 ) ;
 assign wire7881 = ( wire849 ) | ( wire7879 ) | ( wire86  &  wire543 ) ;
 assign wire7882 = ( wire7881 ) | ( wire850 ) ;
 assign wire7885 = ( i_36_  &  (~ i_35_)  &  n_n1433  &  n_n1375 ) ;
 assign wire7886 = ( i_21_  &  n_n1216  &  wire6959 ) ;
 assign wire7887 = ( n_n1263  &  wire80  &  wire86 ) ;
 assign wire7888 = ( i_34_  &  i_36_  &  n_n1375  &  n_n1400 ) ;
 assign wire7889 = ( i_34_  &  n_n1288  &  n_n1018 ) ;
 assign wire7890 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_12_)  &  (~ i_21_) ) ;
 assign wire7892 = ( n_n355  &  wire458 ) | ( n_n458  &  wire7889 ) ;
 assign wire7893 = ( n_n608  &  wire7885 ) | ( n_n242  &  wire7888 ) ;
 assign wire7895 = ( wire841 ) | ( wire7893 ) | ( wire610  &  wire7886 ) ;
 assign wire7896 = ( i_31_  &  (~ i_34_)  &  i_35_  &  wire267 ) ;
 assign wire7897 = ( i_36_  &  (~ i_35_)  &  n_n1369  &  n_n1128 ) ;
 assign wire7898 = ( (~ i_23_)  &  (~ i_24_)  &  (~ i_19_) ) ;
 assign wire7899 = ( i_31_  &  i_34_  &  n_n1429  &  n_n1375 ) ;
 assign wire7900 = ( i_2_  &  (~ i_9_) ) ;
 assign wire7901 = ( (~ i_10_)  &  (~ i_13_)  &  (~ i_17_)  &  (~ i_16_) ) ;
 assign wire7902 = ( (~ i_32_)  &  n_n1375  &  n_n1213 ) ;
 assign wire7903 = ( n_n242  &  wire458 ) | ( n_n458  &  wire7902 ) ;
 assign wire7906 = ( wire669  &  wire7896 ) | ( wire491  &  wire7897 ) ;
 assign wire7907 = ( wire833 ) | ( n_n712  &  wire7898  &  wire7899 ) ;
 assign wire7909 = ( wire7906 ) | ( wire7907 ) | ( n_n1147  &  wire383 ) ;
 assign wire7910 = ( (~ i_32_)  &  i_36_  &  n_n1375  &  n_n1213 ) ;
 assign wire7911 = ( n_n1314  &  wire80  &  wire86 ) ;
 assign wire7912 = ( i_36_  &  n_n793  &  wire6923 ) ;
 assign wire7913 = ( (~ i_32_)  &  (~ i_31_)  &  (~ i_29_)  &  n_n1441 ) ;
 assign wire7914 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_29_)  &  n_n1433 ) ;
 assign wire7915 = ( n_n608  &  wire7913 ) | ( n_n544  &  wire7914 ) ;
 assign wire7916 = ( n_n358  &  wire7910 ) | ( n_n263  &  wire7912 ) ;
 assign wire7917 = ( wire493  &  n_n269 ) | ( wire360  &  wire7911 ) ;
 assign wire7918 = ( wire825 ) | ( n_n1089  &  wire383 ) ;
 assign wire7920 = ( wire7918 ) | ( n_n880  &  wire829 ) | ( n_n880  &  wire7915 ) ;
 assign wire7921 = ( wire834 ) | ( wire843 ) | ( wire7895 ) | ( wire7909 ) ;
 assign wire7923 = ( n_n1568 ) | ( wire7852 ) | ( wire7853 ) | ( wire7921 ) ;
 assign wire7926 = ( n_n1438  &  wire6948  &  wire6949 ) | ( n_n1438  &  wire6948  &  wire7653 ) ;
 assign wire7927 = ( wire813 ) | ( n_n1374  &  n_n1375  &  wire38 ) ;
 assign wire7930 = ( (~ i_32_)  &  (~ i_34_)  &  i_36_  &  (~ i_35_) ) ;
 assign wire7931 = ( (~ i_32_)  &  i_34_  &  i_36_  &  (~ i_35_) ) ;
 assign wire7932 = ( (~ i_27_)  &  (~ i_28_)  &  (~ i_26_)  &  i_33_ ) ;
 assign wire7935 = ( wire512 ) | ( wire38  &  wire7932 ) ;
 assign wire7936 = ( wire112 ) | ( wire507 ) | ( wire372  &  wire7029 ) ;
 assign wire7938 = ( wire494 ) | ( wire497 ) | ( wire7935 ) | ( wire7936 ) ;
 assign wire7940 = ( (~ i_31_)  &  (~ i_30_) ) ;
 assign wire7941 = ( (~ i_30_)  &  (~ i_31_)  &  n_n1375  &  wire86 ) ;
 assign wire7942 = ( i_21_  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire7945 = ( (~ i_2_)  &  i_36_  &  n_n825 ) ;
 assign wire7946 = ( (~ i_8_)  &  (~ i_12_)  &  n_n1345 ) ;
 assign wire7947 = ( i_36_  &  (~ i_35_)  &  n_n1369  &  n_n1254 ) ;
 assign wire7949 = ( (~ i_30_)  &  (~ i_7_)  &  (~ i_28_)  &  (~ i_29_) ) ;
 assign wire7952 = ( wire299  &  wire572 ) | ( wire342  &  wire7941 ) ;
 assign wire7953 = ( wire471 ) | ( n_n1429  &  wire478 ) ;
 assign wire7954 = ( wire469 ) | ( (~ i_13_)  &  wire7946  &  wire7947 ) ;
 assign wire7957 = ( (~ i_2_)  &  i_36_  &  n_n1443 ) ;
 assign wire7958 = ( n_n1441  &  wire77  &  wire7831 ) ;
 assign wire7959 = ( n_n1441  &  n_n1390  &  wire6993 ) ;
 assign wire7960 = ( (~ i_30_)  &  (~ i_31_)  &  wire258  &  wire86 ) ;
 assign wire7961 = ( (~ i_2_)  &  i_36_  &  n_n825 ) ;
 assign wire7963 = ( wire7957  &  wire7958 ) | ( wire385  &  wire7959 ) ;
 assign wire7964 = ( wire417 ) | ( n_n1375  &  n_n1400  &  wire7960 ) ;
 assign wire7965 = ( wire424 ) | ( n_n1375  &  wire427 ) | ( n_n1375  &  wire439 ) ;
 assign wire7968 = ( (~ i_31_)  &  (~ i_30_) ) ;
 assign wire7969 = ( i_20_  &  (~ i_28_)  &  (~ i_21_)  &  i_29_ ) ;
 assign wire7971 = ( (~ i_23_)  &  (~ i_17_)  &  i_21_ ) ;
 assign wire7976 = ( i_36_  &  (~ i_21_) ) ;
 assign wire7978 = ( wire234 ) | ( n_n1202  &  wire7968  &  wire7969 ) ;
 assign wire7979 = ( wire350 ) | ( n_n984  &  n_n1213  &  wire608 ) ;
 assign wire7980 = ( wire336 ) | ( wire304 ) ;
 assign wire7981 = ( wire339 ) | ( (~ i_13_)  &  (~ i_16_)  &  wire301 ) ;
 assign wire7984 = ( i_21_  &  i_25_ ) ;
 assign wire7986 = ( (~ i_30_)  &  (~ i_31_)  &  wire259  &  wire86 ) ;
 assign wire7989 = ( wire192 ) | ( wire194 ) ;
 assign wire7990 = ( wire197 ) | ( n_n1375  &  n_n1400  &  wire7986 ) ;
 assign wire7991 = ( wire198 ) | ( (~ i_14_)  &  (~ i_16_)  &  wire301 ) ;
 assign wire7994 = ( i_36_  &  (~ i_35_)  &  wire259  &  n_n1459 ) ;
 assign wire7997 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  (~ i_17_) ) ;
 assign wire7999 = ( (~ i_23_)  &  i_34_  &  i_33_ ) ;
 assign wire8002 = ( wire185 ) | ( wire183 ) ;
 assign wire8003 = ( wire184 ) | ( wire187 ) | ( wire74  &  wire7994 ) ;
 assign wire8006 = ( (~ i_28_)  &  (~ i_32_)  &  (~ i_29_)  &  wire79 ) ;
 assign wire8007 = ( n_n263  &  wire273 ) | ( n_n269  &  wire256 ) ;
 assign wire8008 = ( (~ i_2_)  &  (~ i_17_)  &  (~ i_21_)  &  (~ i_16_) ) ;
 assign wire8010 = ( (~ i_27_)  &  (~ i_26_)  &  (~ i_2_)  &  (~ i_24_) ) ;
 assign wire8014 = ( wire178 ) | ( (~ i_14_)  &  wire7946  &  wire7947 ) ;
 assign wire8016 = ( wire172 ) | ( wire8014 ) | ( n_n620  &  wire8006 ) ;
 assign wire8019 = ( i_36_  &  (~ i_35_)  &  n_n1441  &  n_n1133 ) ;
 assign wire8021 = ( (~ i_18_)  &  i_3_ ) ;
 assign wire8022 = ( i_10_  &  i_7_  &  (~ i_23_)  &  (~ i_24_) ) ;
 assign wire8023 = ( wire163 ) | ( n_n544  &  wire8019 ) ;
 assign wire8026 = ( wire166 ) | ( wire167 ) | ( i_36_  &  wire712 ) ;
 assign wire8027 = ( (~ i_27_)  &  (~ i_23_)  &  (~ i_24_)  &  i_34_ ) ;
 assign wire8028 = ( (~ i_28_)  &  i_31_  &  (~ i_29_)  &  wire8027 ) ;
 assign wire8029 = ( (~ i_2_)  &  i_36_  &  n_n1408 ) ;
 assign wire8030 = ( n_n1441  &  wire77  &  wire7831 ) ;
 assign wire8031 = ( (~ i_13_)  &  (~ i_17_)  &  (~ i_16_)  &  wire305 ) ;
 assign wire8035 = ( wire8029  &  wire8030 ) | ( wire723  &  wire8031 ) ;
 assign wire8036 = ( wire160 ) | ( n_n1288  &  wire79  &  n_n269 ) ;
 assign wire8037 = ( wire158 ) | ( wire161 ) | ( wire724  &  wire8028 ) ;
 assign wire8039 = ( (~ i_13_)  &  (~ i_12_)  &  (~ i_16_)  &  wire305 ) ;
 assign wire8041 = ( i_36_  &  n_n1375  &  n_n1213 ) ;
 assign wire8042 = ( i_14_  &  (~ i_13_)  &  (~ i_12_)  &  (~ i_16_) ) ;
 assign wire8043 = ( (~ i_16_)  &  i_31_  &  (~ i_34_)  &  i_35_ ) ;
 assign wire8046 = ( n_n1404  &  wire478 ) | ( n_n263  &  wire8041 ) ;
 assign wire8047 = ( wire142 ) | ( wire150 ) | ( wire731  &  wire8039 ) ;
 assign wire8049 = ( n_n1576 ) | ( n_n1578 ) ;
 assign wire8052 = ( n_n1572 ) | ( wire164 ) | ( wire8023 ) | ( wire8026 ) ;
 assign wire8054 = ( n_n1574 ) | ( n_n1575 ) | ( n_n1577 ) | ( n_n1573 ) ;
 assign wire8056 = ( i_25_  &  (~ i_32_)  &  (~ i_31_)  &  i_33_ ) ;
 assign wire8057 = ( i_31_  &  (~ i_28_) ) ;
 assign wire8061 = ( wire133 ) | ( wire355  &  wire550 ) ;
 assign wire8062 = ( wire124 ) | ( wire132 ) | ( wire130 ) | ( wire134 ) ;
 assign wire8065 = ( i_21_  &  i_25_ ) ;
 assign wire8067 = ( wire117 ) | ( wire415  &  n_n1254  &  wire355 ) ;
 assign wire8071 = ( wire110 ) | ( wire43  &  n_n1282  &  wire355 ) ;
 assign wire8072 = ( wire111 ) | ( wire1651 ) | ( wire1652 ) ;
 assign wire8077 = ( n_n1580 ) | ( n_n1579 ) | ( n_n1581 ) | ( n_n1583 ) ;
 assign wire8079 = ( n_n1556 ) | ( n_n1582 ) | ( n_n1584 ) | ( wire8077 ) ;
 assign wire8082 = ( (~ i_7_)  &  (~ i_11_)  &  (~ i_19_) ) ;
 assign wire8084 = ( (~ i_23_)  &  (~ i_21_)  &  wire232  &  wire8082 ) ;
 assign wire8085 = ( i_36_  &  n_n793  &  wire6923 ) ;
 assign wire8086 = ( (~ i_7_)  &  (~ i_8_)  &  (~ i_19_) ) ;
 assign wire8090 = ( (~ i_17_)  &  i_36_  &  n_n1406  &  n_n1213 ) ;
 assign wire8091 = ( (~ i_9_)  &  (~ i_7_)  &  (~ i_6_)  &  (~ i_23_) ) ;
 assign wire8093 = ( wire34 ) | ( wire462  &  wire8084 ) ;
 assign wire8094 = ( wire22 ) | ( (~ i_21_)  &  wire101 ) | ( (~ i_21_)  &  wire102 ) ;
 assign wire8096 = ( wire945 ) | ( wire7781 ) | ( wire8093 ) | ( wire8094 ) ;


endmodule

