module ex5p (
	i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, 
	o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_, 
	o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, 
	o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, 
	o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_, 
	o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_, 
	o_53_, o_46_, o_61_, o_9_, o_62_, o_49_, o_7_, o_8_, o_5_, o_59_, 
	o_6_, o_3_, o_4_);

input i_7_;
input i_5_;
input i_6_;
input i_3_;
input i_4_;
input i_1_;
input i_2_;
input i_0_;
output o_1_;
output o_19_;
output o_2_;
output o_0_;
output o_29_;
output o_60_;
output o_39_;
output o_38_;
output o_25_;
output o_12_;
output o_37_;
output o_26_;
output o_11_;
output o_50_;
output o_36_;
output o_27_;
output o_14_;
output o_35_;
output o_28_;
output o_13_;
output o_34_;
output o_21_;
output o_16_;
output o_40_;
output o_33_;
output o_22_;
output o_15_;
output o_32_;
output o_23_;
output o_18_;
output o_31_;
output o_24_;
output o_17_;
output o_56_;
output o_43_;
output o_30_;
output o_55_;
output o_44_;
output o_58_;
output o_41_;
output o_57_;
output o_42_;
output o_20_;
output o_52_;
output o_47_;
output o_51_;
output o_48_;
output o_54_;
output o_45_;
output o_10_;
output o_53_;
output o_46_;
output o_61_;
output o_9_;
output o_62_;
output o_49_;
output o_7_;
output o_8_;
output o_5_;
output o_59_;
output o_6_;
output o_3_;
output o_4_;
wire n_n1154;
wire n_n1245;
wire n_n1215;
wire n_n1274;
wire n_n1305;
wire n_n744;
wire wire248;
wire n_n1121;
wire n_n1180;
wire n_n1211;
wire n_n1271;
wire n_n1302;
wire wire246;
wire wire354;
wire n_n1168;
wire n_n1321;
wire n_n1169;
wire wire73;
wire wire92;
wire wire93;
wire wire94;
wire wire146;
wire wire147;
wire wire186;
wire wire208;
wire wire249;
wire n_n0;
wire n_n1120;
wire n_n1008;
wire n_n1009;
wire n_n872;
wire n_n958;
wire n_n949;
wire wire108;
wire wire115;
wire wire152;
wire wire187;
wire wire192;
wire wire222;
wire wire226;
wire wire228;
wire wire240;
wire wire252;
wire wire280;
wire wire301;
wire wire324;
wire wire327;
wire wire330;
wire wire331;
wire wire346;
wire n_n1193;
wire n_n1225;
wire n_n1197;
wire n_n936;
wire n_n1194;
wire n_n136;
wire n_n1028;
wire n_n137;
wire n_n1029;
wire n_n935;
wire wire184;
wire wire218;
wire wire326;
wire wire348;
wire n_n1261;
wire n_n573;
wire n_n616;
wire n_n617;
wire n_n602;
wire wire88;
wire wire114;
wire wire196;
wire wire298;
wire wire318;
wire wire319;
wire n_n7;
wire n_n5;
wire wire82;
wire n_n1196;
wire n_n1287;
wire n_n1163;
wire n_n1049;
wire n_n864;
wire n_n1318;
wire n_n1189;
wire n_n1061;
wire n_n756;
wire n_n1083;
wire n_n215;
wire n_n1135;
wire wire250;
wire wire285;
wire wire297;
wire wire309;
wire wire333;
wire wire337;
wire wire341;
wire wire343;
wire n_n1181;
wire n_n6;
wire n_n427;
wire n_n459;
wire n_n973;
wire n_n1134;
wire n_n904;
wire n_n996;
wire wire87;
wire wire200;
wire wire261;
wire n_n1255;
wire n_n1256;
wire n_n1229;
wire n_n953;
wire n_n1203;
wire n_n845;
wire wire110;
wire wire177;
wire wire182;
wire wire189;
wire wire310;
wire wire339;
wire n_n4;
wire wire102;
wire n_n13;
wire n_n1056;
wire wire84;
wire wire129;
wire wire153;
wire wire155;
wire wire201;
wire wire221;
wire n_n2;
wire n_n950;
wire n_n805;
wire n_n804;
wire n_n803;
wire n_n1208;
wire wire104;
wire wire116;
wire wire159;
wire wire162;
wire wire164;
wire wire178;
wire wire288;
wire wire293;
wire n_n11;
wire wire66;
wire n_n923;
wire n_n814;
wire n_n822;
wire n_n1122;
wire n_n1288;
wire n_n963;
wire n_n1006;
wire n_n1204;
wire wire76;
wire wire86;
wire wire111;
wire wire130;
wire wire136;
wire wire154;
wire wire253;
wire wire274;
wire wire276;
wire wire291;
wire wire305;
wire wire345;
wire n_n17;
wire n_n128;
wire n_n1002;
wire wire156;
wire wire193;
wire wire255;
wire wire284;
wire wire313;
wire wire332;
wire n_n3;
wire n_n1010;
wire n_n1283;
wire n_n95;
wire n_n1334;
wire n_n580;
wire n_n1017;
wire n_n1314;
wire n_n1282;
wire n_n925;
wire n_n990;
wire wire179;
wire wire230;
wire wire237;
wire wire238;
wire wire279;
wire wire180;
wire n_n1300;
wire n_n490;
wire n_n387;
wire n_n1258;
wire n_n534;
wire n_n926;
wire n_n1018;
wire n_n1022;
wire wire83;
wire wire183;
wire wire229;
wire wire247;
wire wire257;
wire wire300;
wire n_n1254;
wire n_n813;
wire n_n961;
wire n_n1330;
wire n_n642;
wire n_n1316;
wire n_n574;
wire n_n921;
wire n_n371;
wire wire109;
wire wire112;
wire wire254;
wire wire259;
wire wire314;
wire n_n19;
wire n_n660;
wire n_n673;
wire n_n563;
wire wire99;
wire wire127;
wire wire137;
wire wire197;
wire wire235;
wire wire315;
wire wire325;
wire n_n906;
wire wire141;
wire wire165;
wire wire223;
wire wire267;
wire n_n895;
wire n_n745;
wire wire85;
wire wire181;
wire wire209;
wire wire283;
wire wire292;
wire n_n1216;
wire n_n1244;
wire n_n554;
wire n_n810;
wire n_n809;
wire n_n1269;
wire n_n800;
wire wire150;
wire wire195;
wire wire287;
wire wire308;
wire wire321;
wire wire322;
wire wire340;
wire wire342;
wire n_n1224;
wire n_n711;
wire n_n1284;
wire n_n1076;
wire wire95;
wire wire107;
wire wire217;
wire wire231;
wire wire260;
wire wire295;
wire wire347;
wire n_n581;
wire n_n742;
wire n_n1243;
wire n_n1034;
wire n_n824;
wire wire97;
wire wire101;
wire wire271;
wire wire320;
wire n_n817;
wire n_n960;
wire n_n1165;
wire n_n989;
wire n_n821;
wire n_n1322;
wire wire139;
wire wire207;
wire wire277;
wire n_n1139;
wire n_n553;
wire n_n1138;
wire n_n930;
wire n_n1021;
wire wire113;
wire wire148;
wire wire158;
wire wire161;
wire wire194;
wire wire198;
wire n_n476;
wire wire263;
wire wire264;
wire wire265;
wire n_n1147;
wire n_n1238;
wire n_n1155;
wire n_n1253;
wire n_n1231;
wire n_n738;
wire n_n468;
wire n_n716;
wire wire266;
wire wire278;
wire wire290;
wire wire323;
wire wire268;
wire n_n1239;
wire n_n1268;
wire n_n948;
wire wire135;
wire wire173;
wire n_n1015;
wire wire233;
wire wire281;
wire n_n1167;
wire n_n10;
wire n_n955;
wire n_n883;
wire n_n901;
wire wire269;
wire wire306;
wire n_n1;
wire n_n582;
wire n_n1148;
wire n_n1104;
wire n_n8;
wire n_n1119;
wire n_n1133;
wire n_n1303;
wire n_n1170;
wire n_n826;
wire n_n1023;
wire n_n1024;
wire n_n786;
wire n_n1025;
wire n_n1273;
wire n_n1301;
wire n_n1077;
wire n_n1228;
wire n_n1137;
wire n_n1319;
wire n_n1074;
wire n_n14;
wire wire270;
wire n_n15;
wire n_n859;
wire n_n12;
wire n_n1192;
wire n_n934;
wire n_n1285;
wire wire243;
wire wire273;
wire n_n1153;
wire n_n1230;
wire wire71;
wire n_n1257;
wire n_n1040;
wire n_n937;
wire wire69;
wire n_n802;
wire n_n1226;
wire n_n1298;
wire wire77;
wire n_n823;
wire n_n9;
wire wire67;
wire n_n962;
wire n_n1329;
wire wire128;
wire n_n609;
wire wire286;
wire n_n1272;
wire wire160;
wire n_n1320;
wire n_n858;
wire wire64;
wire n_n1020;
wire n_n1315;
wire n_n16;
wire wire72;
wire wire236;
wire wire163;
wire wire242;
wire n_n1223;
wire n_n931;
wire wire353;
wire n_n1227;
wire n_n1275;
wire wire132;
wire wire98;
wire n_n18;
wire n_n910;
wire n_n909;
wire n_n911;
wire n_n792;
wire n_n1013;
wire wire225;
wire n_n1136;
wire n_n825;
wire wire70;
wire n_n799;
wire wire134;
wire wire78;
wire wire302;
wire wire211;
wire n_n1213;
wire n_n1166;
wire n_n1037;
wire n_n1014;
wire wire219;
wire wire215;
wire n_n1032;
wire wire303;
wire n_n797;
wire wire316;
wire n_n1033;
wire wire191;
wire wire106;
wire wire133;
wire wire138;
wire wire140;
wire wire216;
wire wire174;
wire wire412;
wire wire413;
wire wire414;
wire wire421;
wire wire426;
wire wire434;
wire wire450;
wire wire456;
wire wire461;
wire wire462;
wire wire466;
wire wire468;
wire wire471;
wire wire473;
wire wire476;
wire wire483;
wire wire487;
wire wire488;
wire wire493;
wire wire500;
wire wire504;
wire wire505;
wire wire507;
wire wire512;
wire wire515;
wire wire532;
wire wire534;
wire wire545;
wire wire546;
wire wire549;
wire wire551;
wire wire561;
wire wire564;
wire wire568;
wire wire588;
wire wire592;
wire wire3176;
wire wire3177;
wire wire3178;
wire wire3179;
wire wire3180;
wire wire3184;
wire wire3188;
wire wire3189;
wire wire3190;
wire wire3191;
wire wire3195;
wire wire3196;
wire wire3203;
wire wire3204;
wire wire3205;
wire wire3206;
wire wire3209;
wire wire3210;
wire wire3213;
wire wire3216;
wire wire3217;
wire wire3218;
wire wire3221;
wire wire3222;
wire wire3225;
wire wire3236;
wire wire3237;
wire wire3238;
wire wire3239;
wire wire3243;
wire wire3244;
wire wire3245;
wire wire3248;
wire wire3250;
wire wire3251;
wire wire3255;
wire wire3256;
wire wire3257;
wire wire3261;
wire wire3262;
wire wire3264;
wire wire3266;
wire wire3267;
wire wire3268;
wire wire3269;
wire wire3273;
wire wire3274;
wire wire3277;
wire wire3278;
wire wire3279;
wire wire3282;
wire wire3283;
wire wire3285;
wire wire3286;
wire wire3287;
wire wire3288;
wire wire3290;
wire wire3292;
wire wire3294;
wire wire3296;
wire wire3299;
wire wire3304;
wire wire3305;
wire wire3309;
wire wire3311;
wire wire3312;
wire wire3313;
wire wire3316;
wire wire3317;
wire wire3318;
wire wire3319;
wire wire3320;
wire wire3321;
wire wire3322;
wire wire3327;
wire wire3328;
wire wire3329;
wire wire3332;
wire wire3333;
wire wire3334;
wire wire3340;
wire wire3341;
wire wire3342;
wire wire3344;
wire wire3345;
wire wire3348;
wire wire3349;
wire wire3350;
wire wire3351;
wire wire3353;
wire wire3355;
wire wire3358;
wire wire3359;
wire wire3360;
wire wire3361;
wire wire3363;
wire wire3366;
wire wire3367;
wire wire3368;
wire wire3369;
wire wire3370;
wire wire3373;
wire wire3375;
wire wire3377;
wire wire3378;
wire wire3379;
wire wire3381;
wire wire3383;
wire wire3384;
wire wire3387;
wire wire3388;
wire wire3390;
wire wire3393;
wire wire3395;
wire wire3400;
wire wire3404;
wire wire3405;
wire wire3406;
wire wire3407;
wire wire3408;
wire wire3410;
wire wire3411;
wire wire3413;
wire wire3414;
wire wire3417;
wire wire3418;
wire wire3420;
wire wire3422;
wire wire3424;
wire wire3425;
wire wire3428;
wire wire3430;
wire wire3432;
wire wire3433;
wire wire3434;
wire wire3435;
wire wire3436;
wire wire3437;
wire wire3439;
wire wire3440;
wire wire3441;
wire wire3442;
wire wire3443;
wire wire3446;
wire wire3447;
wire wire3448;
wire wire3452;
wire wire3453;
wire wire3454;
wire wire3455;
wire wire3458;
wire wire3460;
wire wire3462;
wire wire3464;
wire wire3465;
wire wire3467;
wire wire3470;
wire wire3471;
wire wire3472;
wire wire3474;
wire wire3475;
wire wire3477;
wire wire3480;
wire wire3481;
wire wire3482;
wire wire3485;
wire wire3486;
wire wire3487;
wire wire3488;
wire wire3491;
wire wire3492;
wire wire3493;
wire wire3494;
wire wire3495;
wire wire3496;
wire wire3497;
wire wire3498;
wire wire3502;
wire wire3503;
wire wire3505;
wire wire3506;
wire wire3507;
wire wire3510;
wire wire3511;
wire wire3515;
wire wire3516;
wire wire3517;
wire wire3518;
wire wire3519;
wire wire3520;
wire wire3521;
wire wire3526;
wire wire3527;
wire wire3528;
wire wire3533;
wire wire3535;
wire wire3541;
wire wire3542;
wire wire3545;
wire wire3546;
wire wire3548;
wire wire3552;
wire wire3554;
wire wire3556;
wire wire3557;
wire wire3558;
wire wire3560;
wire wire3561;
wire wire3566;
wire wire3567;
wire wire3568;
wire wire3569;
wire wire3573;
wire wire3577;
wire wire3579;
wire wire3581;
wire wire3582;
wire wire3585;
wire wire3586;
wire wire3587;
wire wire3588;
wire wire3589;
wire wire3590;
wire wire3592;
wire wire3598;
wire wire3599;
wire wire3600;
wire wire3601;
wire wire3604;
wire wire3605;
wire wire3607;
wire wire3609;
wire wire3610;
wire wire3612;
wire wire3613;
wire wire3614;
wire wire3615;
wire wire3616;
wire wire3618;
wire wire3619;
wire wire3621;
wire wire3623;
wire wire3624;
wire wire3628;
wire wire3630;
wire wire3631;
wire wire3632;
wire wire3635;
wire wire3636;
wire wire3638;
wire wire3639;
wire wire3641;
wire wire3643;
wire wire3644;
wire wire3645;
wire wire3652;
wire wire3653;
wire wire3654;
wire wire3655;
wire wire3658;
wire wire3659;
wire wire3660;
wire wire3663;
wire wire3667;
wire wire3668;
wire wire3669;
wire wire3671;
wire wire3672;
wire wire3674;
wire wire3676;
wire wire3679;
wire wire3682;
wire wire3686;
wire wire3687;
wire wire3688;
wire wire3689;
wire wire3690;
wire wire3691;
wire wire3692;
wire wire3693;
wire wire3695;
wire wire3702;
wire wire3703;
wire wire3704;
wire wire3705;
wire wire3706;
wire wire3710;
wire wire3712;
wire wire3713;
wire wire3714;
wire wire3715;
wire wire3716;
wire wire3717;
wire wire3719;
wire wire3722;
wire wire3723;
wire wire3724;
wire wire3725;
wire wire3730;
wire wire3731;
wire wire3732;
wire wire3733;
wire wire3736;
wire wire3739;
wire wire3743;
wire wire3744;
wire wire3745;
wire wire3749;
wire wire3750;
wire wire3751;
wire wire3754;
wire wire3756;
wire wire3758;
wire wire3759;
wire wire3760;
wire wire3763;
wire wire3764;
wire wire3765;
wire wire3767;
wire wire3770;
wire wire3772;
wire wire3774;
wire wire3775;
wire wire3777;
wire wire3781;
wire wire3782;
wire wire3784;
wire wire3786;
wire wire3789;
wire wire3790;
wire wire3792;
wire wire3795;
wire wire3796;
wire wire3797;
wire wire3798;
wire wire3800;
wire wire3801;
wire wire3802;
wire wire3804;
wire wire3806;
wire wire3807;
wire wire3808;
wire wire3809;
wire wire3810;
wire wire3813;
wire wire3816;
wire wire3818;
wire wire3820;
wire wire3821;
wire wire3822;
wire wire3823;
wire wire3827;
wire wire3829;
wire wire3830;
wire wire3831;
wire wire3832;
wire wire3841;
wire wire3842;
wire wire3843;
wire wire3844;
wire wire3847;
wire wire3850;
wire wire3853;
wire wire3854;
wire wire3855;
wire wire3856;
wire wire3857;
wire wire3860;
wire wire3864;
wire wire3868;
wire wire3870;
wire wire3871;
wire wire3872;
wire wire3873;
wire wire3874;
wire wire3875;
wire wire3876;
wire wire3877;
wire wire3882;
wire wire3883;
wire wire3885;
wire wire3886;
wire wire3890;
wire wire3892;
wire wire3897;
wire wire3899;
wire wire3900;
wire wire3903;
wire wire3905;
wire wire3908;
wire wire3909;
wire wire3910;
wire wire3911;
wire wire3915;
wire wire3916;
wire wire3920;
wire wire3921;
wire wire3922;
wire wire3925;
wire wire3926;
wire wire3928;
wire wire3929;
wire wire3935;
wire wire3936;
wire wire3937;
wire wire3938;
wire wire3939;
wire wire3940;
wire wire3941;
wire wire3942;
wire wire3944;
wire wire3945;
wire wire3950;
wire wire3951;
wire wire3952;
wire wire3955;
wire wire3957;
wire wire3958;
wire wire3962;
wire wire3965;
wire wire3966;
wire wire3967;
wire wire3968;
wire wire3969;
wire wire3973;
wire wire3975;
wire wire3976;
wire wire3978;
wire wire3982;
wire wire3983;
wire wire3985;
wire wire3986;
wire wire3993;
wire wire3994;
wire wire3995;
wire wire3997;
wire wire3998;
wire wire4001;
wire wire4003;
wire wire4004;
wire wire4005;
wire wire4006;
wire wire4007;
wire wire4008;
wire wire4009;
wire wire4013;
wire wire4014;
wire wire4015;
wire wire4016;
wire wire4019;
wire wire4020;
wire wire4023;
wire wire4024;
wire wire4025;
wire wire4027;
wire wire4029;
wire wire4031;
wire wire4037;
wire wire4038;
wire wire4039;
wire wire4042;
wire wire4044;
wire wire4046;
wire wire4047;
wire wire4050;
wire wire4051;
wire wire4053;
wire wire4055;
wire wire4056;
wire wire4057;
wire wire4058;
wire wire4063;
wire wire4065;
wire wire4066;
wire wire4068;
wire wire4069;
wire wire4071;
wire wire4074;
wire wire4076;
wire wire4079;
wire wire4081;
wire wire4082;
wire wire4083;
wire wire4084;
wire wire4086;
wire wire4090;
wire wire4091;
wire wire4092;
wire wire4093;
wire wire4094;
wire wire4097;
wire wire4098;
wire wire4099;
wire wire4100;
wire wire4101;
wire wire4105;
wire wire4106;
wire wire4108;
wire wire4109;
wire wire4112;
wire wire4113;
wire wire4115;
wire wire4117;
wire wire4119;
wire wire4122;
wire wire4123;
wire wire4125;
wire wire4126;
wire wire4127;
wire wire4128;
wire wire4129;
wire wire4138;
wire wire4139;
wire wire4140;
wire wire4141;
wire wire4142;
wire wire4144;
wire wire4145;
wire wire4149;
wire wire4150;
wire wire4151;
wire wire4152;
wire wire4153;
wire wire4154;
wire wire4160;
wire wire4161;
wire wire4162;
wire wire4163;
wire wire4166;
wire wire4167;
wire wire4168;
wire wire4169;
assign o_1_ = ( wire3179 ) | ( wire3180 ) | ( wire3184 ) ;
 assign o_19_ = ( n_n744 ) | ( wire248 ) | ( n_n0  &  wire71 ) ;
 assign o_2_ = ( wire3188 ) | ( wire3189 ) | ( wire3190 ) | ( wire3191 ) ;
 assign o_0_ = ( wire3204 ) | ( wire3205 ) | ( wire3209 ) ;
 assign o_29_ = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign o_60_ = ( wire3266 ) | ( wire3267 ) | ( wire3268 ) | ( wire3269 ) ;
 assign o_39_ = ( n_n136 ) | ( wire3332 ) | ( wire3333 ) | ( wire3334 ) ;
 assign o_38_ = ( wire3377 ) | ( wire3378 ) | ( wire3381 ) ;
 assign o_25_ = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign o_12_ = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) ;
 assign o_37_ = ( wire3417 ) | ( wire3418 ) | ( wire3424 ) | ( wire3428 ) ;
 assign o_26_ = ( n_n7  &  n_n5  &  n_n17 ) | ( n_n7  &  n_n17  &  n_n19 ) ;
 assign o_11_ = ( i_7_  &  i_6_  &  n_n6  &  n_n8 ) ;
 assign o_50_ = ( wire3452 ) | ( wire3453 ) | ( wire3454 ) | ( wire3455 ) ;
 assign o_36_ = ( wire339 ) | ( wire3480 ) | ( wire3481 ) | ( wire3482 ) ;
 assign o_27_ = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign o_14_ = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign o_35_ = ( wire339 ) | ( wire3502 ) | ( wire3503 ) ;
 assign o_28_ = ( i_7_  &  i_6_  &  n_n5  &  n_n11 ) ;
 assign o_13_ = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) ;
 assign o_34_ = ( n_n136 ) | ( wire3526 ) | ( wire3527 ) | ( wire3528 ) ;
 assign o_21_ = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign o_16_ = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign o_40_ = ( wire3566 ) | ( wire3567 ) | ( wire3568 ) | ( wire3569 ) ;
 assign o_33_ = ( wire3598 ) | ( wire3599 ) | ( wire3600 ) | ( wire3601 ) ;
 assign o_22_ = ( n_n7  &  n_n4  &  n_n17 ) | ( n_n4  &  n_n11  &  n_n17 ) ;
 assign o_15_ = ( i_7_  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign o_32_ = ( wire3614 ) | ( wire3615 ) | ( wire3618 ) ;
 assign o_23_ = ( n_n1017 ) | ( wire3619 ) ;
 assign o_18_ = ( i_7_  &  i_6_  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign o_31_ = ( wire318 ) | ( wire3605 ) | ( wire3632 ) | ( wire3635 ) ;
 assign o_24_ = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign o_17_ = ( wire180 ) | ( wire3636 ) ;
 assign o_56_ = ( wire322 ) | ( wire3639 ) | ( wire3660 ) | ( wire3663 ) ;
 assign o_43_ = ( n_n371 ) | ( wire3705 ) | ( wire3706 ) | ( wire3710 ) ;
 assign o_30_ = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign o_55_ = ( wire3730 ) | ( wire3731 ) | ( wire3732 ) | ( wire3733 ) ;
 assign o_44_ = ( wire339 ) | ( wire3743 ) | ( wire3744 ) | ( wire3745 ) ;
 assign o_58_ = ( wire3763 ) | ( wire3764 ) | ( wire3767 ) ;
 assign o_41_ = ( wire321 ) | ( wire322 ) | ( wire3790 ) | ( wire3795 ) ;
 assign o_57_ = ( wire3829 ) | ( wire3830 ) | ( wire3831 ) | ( wire3832 ) ;
 assign o_42_ = ( wire314 ) | ( wire3876 ) | ( wire3882 ) | ( wire3885 ) ;
 assign o_20_ = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign o_52_ = ( wire3908 ) | ( wire3909 ) | ( wire3910 ) | ( wire3911 ) ;
 assign o_47_ = ( wire3921 ) | ( wire3922 ) | ( wire3925 ) | ( wire3928 ) ;
 assign o_51_ = ( wire3966 ) | ( wire3967 ) | ( wire3968 ) | ( wire3969 ) ;
 assign o_48_ = ( n_n476 ) | ( wire263 ) | ( wire264 ) | ( wire3986 ) ;
 assign o_54_ = ( wire4013 ) | ( wire4014 ) | ( wire4015 ) | ( wire4016 ) ;
 assign o_45_ = ( wire137 ) | ( n_n883 ) | ( wire3355 ) | ( wire4031 ) ;
 assign o_10_ = ( n_n17  &  n_n3  &  n_n8 ) | ( n_n17  &  n_n3  &  n_n12 ) ;
 assign o_53_ = ( wire4055 ) | ( wire4056 ) | ( wire4057 ) | ( wire4058 ) ;
 assign o_46_ = ( wire263 ) | ( wire4068 ) | ( wire4069 ) ;
 assign o_61_ = ( wire3344 ) | ( wire3345 ) | ( wire4093 ) | ( wire4097 ) ;
 assign o_9_ = ( i_7_  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign o_62_ = ( wire267 ) | ( wire347 ) | ( wire4108 ) | ( wire4112 ) ;
 assign o_49_ = ( n_n476 ) | ( wire263 ) | ( wire4117 ) ;
 assign o_7_ = ( i_7_  &  i_6_  &  n_n2  &  n_n8 ) ;
 assign o_8_ = ( i_7_  &  i_6_  &  n_n19  &  n_n8 ) ;
 assign o_5_ = ( wire4126 ) | ( wire4127 ) | ( wire4128 ) | ( wire4129 ) ;
 assign o_59_ = ( wire4160 ) | ( wire4161 ) | ( wire4162 ) | ( wire4163 ) ;
 assign o_6_ = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign o_4_ = ( wire4166 ) | ( wire4167 ) | ( wire4168 ) | ( wire4169 ) ;
 assign n_n1154 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign n_n1245 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign n_n1215 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign n_n1274 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1305 = ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign n_n744 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n10 ) ;
 assign wire248 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign n_n1121 = ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n8 ) ;
 assign n_n1180 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign n_n1211 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n8 ) ;
 assign n_n1271 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign n_n1302 = ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n8 ) ;
 assign wire246 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n8 ) ;
 assign wire354 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n8 ) ;
 assign n_n1168 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign n_n1321 = ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign n_n1169 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign wire73 = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n19 ) ;
 assign wire92 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign wire93 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire94 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire146 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign wire147 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire186 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n5 ) ;
 assign wire208 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire249 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign n_n0 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n1120 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n8 ) ;
 assign n_n1008 = ( n_n1083 ) | ( wire236 ) | ( wire3213 ) ;
 assign n_n1009 = ( n_n19  &  wire163 ) | ( n_n17  &  n_n19  &  n_n12 ) ;
 assign n_n872 = ( i_7_  &  i_6_  &  n_n6  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n18 ) ;
 assign n_n958 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign n_n949 = ( i_7_  &  i_6_  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n4 ) ;
 assign wire108 = ( n_n1137 ) | ( n_n6  &  n_n14  &  n_n12 ) ;
 assign wire115 = ( wire85 ) | ( n_n1021 ) | ( n_n1020 ) ;
 assign wire152 = ( n_n1136 ) | ( n_n6  &  n_n15  &  n_n12 ) ;
 assign wire187 = ( n_n864 ) | ( n_n5  &  wire69 ) ;
 assign wire192 = ( n_n602 ) | ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) ;
 assign wire222 = ( i_7_  &  i_6_  &  n_n6  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n8 ) ;
 assign wire226 = ( n_n930 ) | ( n_n2  &  wire72 ) ;
 assign wire228 = ( wire104 ) | ( n_n1226 ) | ( wire77 ) ;
 assign wire240 = ( wire3221 ) | ( wire3222 ) | ( n_n3  &  wire70 ) ;
 assign wire252 = ( n_n1197 ) | ( wire88 ) | ( n_n955 ) | ( wire3225 ) ;
 assign wire280 = ( n_n950 ) | ( n_n1208 ) | ( wire551 ) ;
 assign wire301 = ( o_18_ ) | ( n_n1271 ) | ( wire254 ) | ( wire269 ) ;
 assign wire324 = ( wire194 ) | ( n_n859 ) | ( n_n5  &  wire72 ) ;
 assign wire327 = ( n_n1121 ) | ( wire94 ) | ( wire134 ) ;
 assign wire330 = ( n_n387 ) | ( wire3237 ) | ( wire3238 ) ;
 assign wire331 = ( wire147 ) | ( wire300 ) | ( wire127 ) ;
 assign wire346 = ( n_n1133 ) | ( wire3239 ) | ( n_n6  &  wire69 ) ;
 assign n_n1193 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign n_n1225 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n1197 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign n_n936 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire69 ) ;
 assign n_n1194 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign n_n136 = ( wire285 ) | ( wire3288 ) | ( wire3290 ) | ( wire3292 ) ;
 assign n_n1028 = ( i_7_  &  i_6_  &  n_n1  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n12 ) ;
 assign n_n137 = ( wire196 ) | ( n_n1316 ) | ( wire306 ) | ( wire3296 ) ;
 assign n_n1029 = ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n935 = ( o_13_ ) | ( n_n1253 ) | ( wire588 ) ;
 assign wire184 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire218 = ( wire209 ) | ( n_n809 ) | ( n_n1223 ) | ( wire3299 ) ;
 assign wire326 = ( wire197 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire348 = ( n_n1203 ) | ( n_n1056 ) | ( wire476 ) ;
 assign n_n1261 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) ;
 assign n_n573 = ( wire287 ) | ( n_n1268 ) | ( wire132 ) ;
 assign n_n616 = ( i_7_  &  i_6_  &  n_n2  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign n_n617 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n10 ) ;
 assign n_n602 = ( o_6_ ) | ( n_n1024 ) | ( n_n1025 ) | ( wire568 ) ;
 assign wire88 = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) ;
 assign wire114 = ( wire76 ) | ( n_n1017 ) ;
 assign wire196 = ( wire128 ) | ( n_n0  &  n_n7  &  n_n17 ) ;
 assign wire298 = ( n_n1028 ) | ( wire162 ) | ( wire243 ) ;
 assign wire318 = ( n_n822 ) | ( n_n826 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire319 = ( n_n800 ) | ( wire195 ) | ( wire138 ) | ( wire3361 ) ;
 assign n_n7 = ( (~ i_5_)  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n5 = ( (~ i_1_)  &  i_2_  &  i_0_ ) ;
 assign wire82 = ( i_7_  &  i_6_  &  n_n8 ) ;
 assign n_n1196 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign n_n1287 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign n_n1163 = ( i_7_  &  i_6_  &  n_n5  &  n_n12 ) ;
 assign n_n1049 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n864 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n18 ) ;
 assign n_n1318 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign n_n1189 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) ;
 assign n_n1061 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign n_n756 = ( i_7_  &  i_6_  &  n_n19  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n10 ) ;
 assign n_n1083 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n12 ) ;
 assign n_n215 = ( n_n845 ) | ( wire128 ) ;
 assign n_n1135 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign wire250 = ( n_n921 ) | ( n_n11  &  wire66  &  n_n1 ) ;
 assign wire285 = ( n_n1121 ) | ( n_n468 ) | ( wire140 ) | ( wire3274 ) ;
 assign wire297 = ( n_n5  &  n_n13 ) | ( n_n5  &  wire70 ) ;
 assign wire309 = ( o_28_ ) | ( wire98 ) | ( n_n1166 ) ;
 assign wire333 = ( wire229 ) | ( wire215 ) | ( wire3387 ) | ( wire3388 ) ;
 assign wire337 = ( n_n1076 ) | ( n_n1077 ) | ( n_n1136 ) ;
 assign wire341 = ( wire237 ) | ( wire139 ) | ( wire3393 ) ;
 assign wire343 = ( n_n895 ) | ( wire173 ) | ( wire3222 ) ;
 assign n_n1181 = ( i_7_  &  i_6_  &  n_n7  &  n_n5 ) ;
 assign n_n6 = ( i_1_  &  (~ i_2_)  &  i_0_ ) ;
 assign n_n427 = ( n_n716 ) | ( wire278 ) | ( wire140 ) | ( wire3274 ) ;
 assign n_n459 = ( n_n906 ) | ( n_n1329 ) | ( wire128 ) ;
 assign n_n973 = ( i_7_  &  i_6_  &  n_n6  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign n_n1134 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign n_n904 = ( n_n1121 ) | ( wire94 ) | ( wire353 ) | ( wire134 ) ;
 assign n_n996 = ( n_n1037 ) | ( wire3312 ) | ( n_n2  &  wire71 ) ;
 assign wire87 = ( o_7_ ) | ( n_n1268 ) | ( n_n1033 ) | ( wire483 ) ;
 assign wire200 = ( wire216 ) | ( wire3304 ) | ( wire3305 ) | ( wire3309 ) ;
 assign wire261 = ( n_n909 ) | ( n_n0  &  n_n10  &  wire67 ) ;
 assign n_n1255 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n1256 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n1229 = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n3 ) ;
 assign n_n953 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign n_n1203 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign n_n845 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign wire110 = ( n_n1029 ) | ( n_n1  &  wire70 ) ;
 assign wire177 = ( n_n826 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire182 = ( n_n858 ) | ( wire3462 ) | ( wire3464 ) ;
 assign wire189 = ( o_20_ ) | ( n_n1211 ) | ( wire279 ) | ( n_n813 ) ;
 assign wire310 = ( n_n822 ) | ( n_n821 ) | ( wire421 ) ;
 assign wire339 = ( wire116 ) | ( wire137 ) | ( n_n883 ) | ( wire3355 ) ;
 assign n_n4 = ( (~ i_1_)  &  (~ i_2_)  &  i_0_ ) ;
 assign wire102 = ( i_7_  &  i_6_  &  n_n12 ) ;
 assign n_n13 = ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign n_n1056 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire84 = ( wire3304 ) | ( wire3305 ) ;
 assign wire129 = ( n_n1283 ) | ( n_n580 ) | ( wire260 ) ;
 assign wire153 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign wire155 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire201 = ( wire148 ) | ( wire487 ) | ( wire488 ) | ( wire3311 ) ;
 assign wire221 = ( n_n996 ) | ( n_n2  &  n_n11  &  n_n17 ) ;
 assign n_n2 = ( i_1_  &  (~ i_2_)  &  (~ i_0_) ) ;
 assign n_n950 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n8 ) ;
 assign n_n805 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n10 ) ;
 assign n_n804 = ( i_1_  &  i_2_  &  (~ i_0_)  &  wire71 ) ;
 assign n_n803 = ( n_n1238 ) | ( n_n1239 ) | ( wire450 ) ;
 assign n_n1208 = ( i_7_  &  i_6_  &  n_n4  &  n_n8 ) ;
 assign wire104 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign wire116 = ( wire3465 ) | ( wire3467 ) | ( n_n3  &  wire69 ) ;
 assign wire159 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire162 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign wire164 = ( wire88 ) | ( n_n4  &  n_n11  &  n_n16 ) ;
 assign wire178 = ( n_n1245 ) | ( wire195 ) | ( wire277 ) | ( wire3361 ) ;
 assign wire288 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire293 = ( n_n4  &  n_n11  &  n_n15 ) | ( n_n4  &  n_n15  &  n_n12 ) ;
 assign n_n11 = ( (~ i_5_)  &  i_3_  &  (~ i_4_) ) ;
 assign wire66 = ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n923 = ( n_n1287 ) | ( n_n1285 ) | ( wire243 ) ;
 assign n_n814 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign n_n822 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n5 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n5 ) ;
 assign n_n1122 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign n_n1288 = ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) ;
 assign n_n963 = ( (~ i_1_)  &  i_2_  &  i_0_  &  wire72 ) ;
 assign n_n1006 = ( n_n1135 ) | ( wire337 ) | ( n_n1137 ) ;
 assign n_n1204 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) ;
 assign wire76 = ( i_7_  &  i_6_  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign wire86 = ( n_n1211 ) | ( wire279 ) | ( n_n813 ) ;
 assign wire111 = ( n_n961 ) | ( n_n5  &  n_n9  &  wire67 ) ;
 assign wire130 = ( i_7_  &  i_6_  &  n_n1  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n12 ) ;
 assign wire136 = ( n_n6  &  n_n18 ) | ( n_n6  &  wire70 ) ;
 assign wire154 = ( o_14_ ) | ( n_n1192 ) | ( wire534 ) | ( wire3535 ) ;
 assign wire253 = ( wire3312 ) | ( n_n2  &  wire71 ) ;
 assign wire274 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) ;
 assign wire276 = ( n_n1238 ) | ( n_n1239 ) | ( wire434 ) ;
 assign wire291 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) ;
 assign wire305 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire345 = ( n_n1253 ) | ( n_n934 ) | ( n_n797 ) ;
 assign n_n17 = ( i_7_  &  i_6_ ) ;
 assign n_n128 = ( wire94 ) | ( n_n973 ) | ( n_n6  &  n_n18 ) ;
 assign n_n1002 = ( n_n1061 ) | ( wire274 ) | ( wire242 ) | ( wire3573 ) ;
 assign wire156 = ( wire186 ) | ( n_n958 ) | ( wire592 ) ;
 assign wire193 = ( o_6_ ) | ( wire298 ) | ( wire110 ) | ( wire568 ) ;
 assign wire255 = ( n_n1074 ) | ( n_n609 ) | ( wire286 ) | ( wire316 ) ;
 assign wire284 = ( n_n1083 ) | ( wire236 ) | ( wire3577 ) ;
 assign wire313 = ( n_n1134 ) | ( n_n673 ) | ( n_n1136 ) ;
 assign wire332 = ( wire114 ) | ( n_n1015 ) | ( n_n1320 ) | ( wire3216 ) ;
 assign n_n3 = ( i_1_  &  i_2_  &  (~ i_0_) ) ;
 assign n_n1010 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign n_n1283 = ( i_7_  &  i_6_  &  n_n1  &  n_n12 ) ;
 assign n_n95 = ( o_25_ ) | ( n_n930 ) | ( n_n1272 ) | ( wire132 ) ;
 assign n_n1334 = ( i_7_  &  i_6_  &  n_n0  &  n_n7 ) ;
 assign n_n580 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n12 ) ;
 assign n_n1017 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign n_n1314 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign n_n1282 = ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n925 = ( i_7_  &  i_6_  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign n_n990 = ( o_24_ ) | ( n_n1334 ) | ( wire128 ) | ( n_n1013 ) ;
 assign wire179 = ( o_6_ ) | ( n_n923 ) | ( n_n921 ) | ( wire3621 ) ;
 assign wire230 = ( o_18_ ) | ( wire130 ) ;
 assign wire237 = ( wire174 ) | ( wire3395 ) | ( n_n0  &  wire70 ) ;
 assign wire238 = ( n_n804 ) | ( n_n803 ) | ( wire283 ) | ( wire3359 ) ;
 assign wire279 = ( i_7_  &  i_6_  &  n_n7  &  n_n4 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) ;
 assign wire180 = ( i_7_  &  i_6_  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign n_n1300 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n8 ) ;
 assign n_n490 = ( n_n809 ) | ( wire322 ) | ( wire3638 ) ;
 assign n_n387 = ( n_n1231 ) | ( wire135 ) | ( wire545 ) | ( wire546 ) ;
 assign n_n1258 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign n_n534 = ( wire254 ) | ( n_n1275 ) | ( wire132 ) ;
 assign n_n926 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign n_n1018 = ( wire266 ) | ( n_n0  &  n_n17  &  n_n12 ) ;
 assign n_n1022 = ( o_9_ ) | ( n_n1302 ) | ( n_n1301 ) ;
 assign wire83 = ( n_n1021 ) | ( n_n0  &  wire64  &  n_n18 ) ;
 assign wire183 = ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign wire229 = ( wire246 ) | ( wire109 ) | ( wire112 ) ;
 assign wire247 = ( n_n13  &  n_n3  &  n_n14 ) | ( n_n3  &  n_n14  &  n_n9 ) ;
 assign wire257 = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire300 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) ;
 assign n_n1254 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) ;
 assign n_n813 = ( i_7_  &  i_6_  &  n_n4  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n8 ) ;
 assign n_n961 = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign n_n1330 = ( i_7_  &  i_6_  &  n_n0  &  n_n8 ) ;
 assign n_n642 = ( wire146 ) | ( wire268 ) | ( n_n1040 ) ;
 assign n_n1316 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign n_n574 = ( wire147 ) | ( n_n1261 ) | ( n_n616 ) | ( n_n617 ) ;
 assign n_n921 = ( i_7_  &  i_6_  &  n_n10  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n10  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n10  &  n_n1 ) ;
 assign n_n371 = ( wire3671 ) | ( wire3672 ) | ( wire3674 ) | ( wire3676 ) ;
 assign wire109 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n8 ) ;
 assign wire112 = ( i_7_  &  i_6_  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign wire254 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire259 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign wire314 = ( wire153 ) | ( wire85 ) | ( n_n1021 ) | ( n_n1020 ) ;
 assign n_n19 = ( i_1_  &  i_2_  &  i_0_ ) ;
 assign n_n660 = ( wire237 ) | ( wire139 ) | ( wire306 ) | ( wire3393 ) ;
 assign n_n673 = ( o_11_ ) | ( n_n1147 ) | ( wire532 ) ;
 assign n_n563 = ( n_n1334 ) | ( wire128 ) | ( wire3296 ) ;
 assign wire99 = ( o_28_ ) | ( wire78 ) | ( n_n1166 ) ;
 assign wire127 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign wire137 = ( n_n1049 ) | ( wire77 ) ;
 assign wire197 = ( n_n822 ) | ( wire291 ) | ( n_n821 ) | ( wire500 ) ;
 assign wire235 = ( n_n1169 ) | ( n_n1170 ) | ( n_n826 ) ;
 assign wire315 = ( n_n814 ) | ( wire154 ) | ( wire97 ) | ( n_n817 ) ;
 assign wire325 = ( o_10_ ) | ( wire112 ) | ( n_n802 ) ;
 assign n_n906 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n7 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n7 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n7 ) ;
 assign wire141 = ( n_n814 ) | ( wire97 ) | ( n_n817 ) ;
 assign wire165 = ( n_n1274 ) | ( wire87 ) | ( wire281 ) | ( n_n1032 ) ;
 assign wire223 = ( n_n1025 ) | ( n_n1  &  n_n9  &  wire64 ) ;
 assign wire267 = ( n_n996 ) | ( wire345 ) | ( n_n1257 ) | ( n_n1040 ) ;
 assign n_n895 = ( n_n949 ) | ( n_n950 ) | ( n_n1208 ) | ( wire551 ) ;
 assign n_n745 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign wire85 = ( wire266 ) | ( n_n0  &  wire102 ) | ( n_n0  &  wire69 ) ;
 assign wire181 = ( wire229 ) | ( wire3387 ) | ( wire3388 ) ;
 assign wire209 = ( i_7_  &  i_6_  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign wire283 = ( n_n1228 ) | ( n_n1227 ) | ( wire3358 ) ;
 assign wire292 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) ;
 assign n_n1216 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) ;
 assign n_n1244 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign n_n554 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign n_n810 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign n_n809 = ( i_7_  &  i_6_  &  n_n13  &  n_n3 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n3 ) ;
 assign n_n1269 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) ;
 assign n_n800 = ( wire277 ) | ( n_n7  &  n_n3  &  n_n14 ) ;
 assign wire150 = ( wire487 ) | ( wire488 ) | ( wire3311 ) ;
 assign wire195 = ( wire112 ) | ( n_n802 ) ;
 assign wire287 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire308 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire321 = ( n_n845 ) | ( n_n858 ) | ( wire3462 ) | ( wire3464 ) ;
 assign wire322 = ( wire189 ) | ( n_n814 ) | ( wire97 ) | ( n_n817 ) ;
 assign wire340 = ( n_n574 ) | ( wire138 ) | ( n_n2  &  wire70 ) ;
 assign wire342 = ( wire187 ) | ( wire99 ) | ( wire191 ) ;
 assign n_n1224 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n12 ) ;
 assign n_n711 = ( n_n937 ) | ( wire3802 ) | ( n_n2  &  wire69 ) ;
 assign n_n1284 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n12 ) ;
 assign n_n1076 = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n12 ) ;
 assign wire95 = ( wire3465 ) | ( n_n3  &  wire69 ) ;
 assign wire107 = ( wire3384 ) | ( n_n1  &  wire69 ) ;
 assign wire217 = ( wire246 ) | ( wire109 ) | ( n_n1243 ) ;
 assign wire231 = ( wire132 ) | ( n_n7  &  n_n2  &  n_n16 ) ;
 assign wire260 = ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n1 ) ;
 assign wire295 = ( o_13_ ) | ( n_n1253 ) | ( n_n934 ) | ( wire588 ) ;
 assign wire347 = ( n_n1002 ) | ( wire3485 ) | ( wire3486 ) | ( wire3804 ) ;
 assign n_n581 = ( wire260 ) | ( n_n17  &  n_n1  &  n_n12 ) ;
 assign n_n742 = ( wire248 ) | ( n_n0  &  n_n17  &  n_n8 ) ;
 assign n_n1243 = ( i_7_  &  i_6_  &  n_n7  &  n_n3 ) ;
 assign n_n1034 = ( o_7_ ) | ( n_n1268 ) | ( wire483 ) ;
 assign n_n824 = ( o_12_ ) | ( wire504 ) | ( wire505 ) ;
 assign wire97 = ( wire288 ) | ( n_n1204 ) | ( wire412 ) | ( wire413 ) ;
 assign wire101 = ( i_7_  &  (~ i_6_)  &  n_n8 ) ;
 assign wire271 = ( i_7_  &  i_6_  &  n_n7  &  n_n5 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n5 ) ;
 assign wire320 = ( wire186 ) | ( n_n958 ) | ( wire180 ) | ( wire592 ) ;
 assign n_n817 = ( i_7_  &  i_6_  &  n_n4  &  n_n11 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign n_n960 = ( wire271 ) | ( n_n5  &  n_n8  &  n_n14 ) ;
 assign n_n1165 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n989 = ( n_n1008 ) | ( wire136 ) | ( wire198 ) | ( wire3886 ) ;
 assign n_n821 = ( i_7_  &  i_6_  &  n_n4  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign n_n1322 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) ;
 assign wire139 = ( n_n1301 ) | ( wire106 ) | ( wire3390 ) ;
 assign wire207 = ( i_7_  &  i_6_  &  n_n1  &  n_n8 ) ;
 assign wire277 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) ;
 assign n_n1139 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign n_n553 = ( i_7_  &  i_6_  &  n_n1  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n8 ) ;
 assign n_n1138 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign n_n930 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign n_n1021 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n1 ) ;
 assign wire113 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n8 ) ;
 assign wire148 = ( n_n554 ) | ( n_n1  &  wire72 ) ;
 assign wire158 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n8 ) ;
 assign wire161 = ( i_7_  &  i_6_  &  n_n11  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n19 ) ;
 assign wire194 = ( n_n1180 ) | ( n_n961 ) | ( wire271 ) | ( n_n962 ) ;
 assign wire198 = ( wire134 ) | ( n_n19  &  n_n8  &  n_n14 ) ;
 assign n_n476 = ( n_n574 ) | ( n_n799 ) | ( wire138 ) | ( wire3973 ) ;
 assign wire263 = ( n_n490 ) | ( n_n883 ) | ( wire3355 ) | ( wire3978 ) ;
 assign wire264 = ( n_n990 ) | ( n_n0  &  wire72 ) ;
 assign wire265 = ( i_7_  &  i_6_  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) ;
 assign n_n1147 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n9 ) ;
 assign n_n1238 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign n_n1155 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) ;
 assign n_n1253 = ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n2 ) ;
 assign n_n1231 = ( i_7_  &  i_6_  &  n_n3  &  n_n10 ) ;
 assign n_n738 = ( wire93 ) | ( wire466 ) ;
 assign n_n468 = ( wire3273 ) | ( n_n6  &  n_n18 ) | ( n_n6  &  wire70 ) ;
 assign n_n716 = ( n_n1083 ) | ( wire236 ) | ( wire473 ) ;
 assign wire266 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign wire278 = ( n_n1009 ) | ( wire471 ) ;
 assign wire290 = ( wire546 ) | ( n_n3  &  n_n10  &  wire67 ) ;
 assign wire323 = ( wire354 ) | ( wire92 ) | ( wire158 ) | ( wire160 ) ;
 assign wire268 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n18 ) ;
 assign n_n1239 = ( i_7_  &  i_6_  &  n_n3  &  n_n8 ) ;
 assign n_n1268 = ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign n_n948 = ( n_n1215 ) | ( n_n1216 ) | ( wire561 ) ;
 assign wire135 = ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n3 ) ;
 assign wire173 = ( wire3221 ) | ( n_n3  &  wire70 ) ;
 assign n_n1015 = ( wire265 ) | ( n_n0  &  n_n11  &  n_n14 ) ;
 assign wire233 = ( wire138 ) | ( n_n2  &  wire70 ) ;
 assign wire281 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) ;
 assign n_n1167 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n11 ) ;
 assign n_n10 = ( i_5_  &  (~ i_3_)  &  i_4_ ) ;
 assign n_n955 = ( n_n1194 ) | ( n_n1196 ) | ( wire242 ) ;
 assign n_n883 = ( wire461 ) | ( wire3341 ) | ( wire3342 ) | ( wire3345 ) ;
 assign n_n901 = ( wire222 ) | ( wire3348 ) ;
 assign wire269 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign wire306 = ( n_n1321 ) | ( wire76 ) | ( n_n1322 ) | ( n_n1320 ) ;
 assign n_n1 = ( (~ i_1_)  &  i_2_  &  (~ i_0_) ) ;
 assign n_n582 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1148 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n8 ) ;
 assign n_n1104 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n12 ) ;
 assign n_n8 = ( i_5_  &  (~ i_3_)  &  (~ i_4_) ) ;
 assign n_n1119 = ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n8 ) ;
 assign n_n1133 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign n_n1303 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign n_n1170 = ( i_7_  &  i_6_  &  n_n5  &  n_n10 ) ;
 assign n_n826 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n10 ) ;
 assign n_n1023 = ( wire3218 ) | ( n_n1  &  n_n14  &  n_n9 ) ;
 assign n_n1024 = ( i_7_  &  i_6_  &  n_n1  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign n_n786 = ( n_n1139 ) | ( n_n1147 ) | ( wire532 ) ;
 assign n_n1025 = ( (~ i_7_)  &  i_6_  &  n_n10  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n10  &  n_n1 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n10  &  n_n1 ) ;
 assign n_n1273 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign n_n1301 = ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n8 ) ;
 assign n_n1077 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign o_3_ = ( (~ i_7_)  &  (~ i_6_)  &  n_n12 ) ;
 assign n_n1228 = ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n3 ) ;
 assign n_n1137 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign n_n1319 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n11 ) ;
 assign n_n1074 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n8 ) ;
 assign n_n14 = ( (~ i_7_)  &  (~ i_6_) ) ;
 assign wire270 = ( o_12_ ) | ( n_n825 ) | ( wire504 ) | ( wire505 ) ;
 assign n_n15 = ( i_7_  &  (~ i_6_) ) ;
 assign n_n859 = ( n_n1169 ) | ( n_n1170 ) | ( wire549 ) ;
 assign n_n12 = ( i_5_  &  i_3_  &  (~ i_4_) ) ;
 assign n_n1192 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign n_n934 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign n_n1285 = ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n12 ) ;
 assign wire243 = ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n12 ) ;
 assign wire273 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) ;
 assign n_n1153 = ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign n_n1230 = ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n3 ) ;
 assign wire71 = ( (~ i_7_)  &  (~ i_6_)  &  n_n10 ) | ( i_7_  &  i_6_  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n9 ) ;
 assign n_n1257 = ( i_7_  &  i_6_  &  n_n2  &  n_n11 ) ;
 assign n_n1040 = ( i_7_  &  i_6_  &  n_n13  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n2 ) ;
 assign n_n937 = ( i_7_  &  i_6_  &  n_n2  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n18 ) ;
 assign wire69 = ( i_7_  &  i_6_  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n18 ) ;
 assign n_n802 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n8 ) ;
 assign n_n1226 = ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign n_n1298 = ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n9 ) ;
 assign wire77 = ( i_7_  &  i_6_  &  n_n11  &  n_n3 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n3 ) ;
 assign n_n823 = ( n_n1180 ) | ( n_n1181 ) | ( wire507 ) ;
 assign n_n9 = ( (~ i_5_)  &  (~ i_3_)  &  i_4_ ) ;
 assign wire67 = ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) | ( (~ i_7_)  &  (~ i_6_) ) ;
 assign n_n962 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign n_n1329 = ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign wire128 = ( i_7_  &  i_6_  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign n_n609 = ( wire3349 ) | ( n_n5  &  n_n13 ) | ( n_n5  &  wire70 ) ;
 assign wire286 = ( i_7_  &  i_6_  &  n_n5  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n18 ) ;
 assign n_n1272 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign wire160 = ( i_7_  &  i_6_  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n6 ) ;
 assign n_n1320 = ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n11 ) ;
 assign n_n858 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n8 ) ;
 assign wire64 = ( i_7_  &  i_6_ ) | ( (~ i_7_)  &  i_6_ ) | ( i_7_  &  (~ i_6_) ) ;
 assign n_n1020 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n18 ) ;
 assign n_n1315 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign n_n16 = ( (~ i_7_)  &  i_6_ ) ;
 assign wire72 = ( i_7_  &  (~ i_6_)  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n10 ) | ( i_7_  &  i_6_  &  n_n9 ) ;
 assign wire236 = ( i_7_  &  i_6_  &  n_n11  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n19 ) ;
 assign wire163 = ( i_5_  &  i_3_  &  i_4_ ) | ( (~ i_5_)  &  i_3_  &  i_4_ ) ;
 assign wire242 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign n_n1223 = ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n3 ) ;
 assign n_n931 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire72 ) ;
 assign wire353 = ( i_1_  &  (~ i_2_)  &  i_0_  &  n_n18 ) ;
 assign n_n1227 = ( i_7_  &  i_6_  &  n_n11  &  n_n3 ) ;
 assign n_n1275 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) ;
 assign wire132 = ( i_7_  &  i_6_  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire98 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n18 = ( i_5_  &  i_3_  &  i_4_ ) ;
 assign n_n910 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n10 ) ;
 assign n_n909 = ( i_7_  &  i_6_  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign n_n911 = ( n_n1321 ) | ( n_n1322 ) | ( n_n1320 ) ;
 assign n_n792 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n18 ) ;
 assign n_n1013 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n9 ) ;
 assign wire225 = ( n_n1076 ) | ( n_n6  &  n_n11  &  n_n17 ) ;
 assign n_n1136 = ( i_7_  &  i_6_  &  n_n6  &  n_n11 ) ;
 assign n_n825 = ( i_7_  &  i_6_  &  n_n5  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign wire70 = ( i_7_  &  i_6_  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n18 ) ;
 assign n_n799 = ( i_1_  &  (~ i_2_)  &  (~ i_0_)  &  wire70 ) ;
 assign wire134 = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) ;
 assign wire78 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n11 ) ;
 assign wire302 = ( n_n1009 ) | ( wire515 ) | ( wire3283 ) ;
 assign wire211 = ( n_n1238 ) | ( n_n1239 ) | ( n_n937 ) | ( wire3238 ) ;
 assign n_n1213 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n4 ) ;
 assign n_n1166 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign n_n1037 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign n_n1014 = ( (~ i_1_)  &  (~ i_2_)  &  (~ i_0_)  &  wire72 ) ;
 assign wire219 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n12 ) ;
 assign wire215 = ( n_n1229 ) | ( wire292 ) | ( n_n1230 ) ;
 assign n_n1032 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n2 ) ;
 assign wire303 = ( wire568 ) | ( n_n11  &  wire66  &  n_n1 ) ;
 assign n_n797 = ( i_7_  &  i_6_  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire316 = ( i_7_  &  i_6_  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n6 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n6 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n6 ) ;
 assign n_n1033 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire191 = ( n_n1163 ) | ( wire98 ) | ( wire564 ) ;
 assign wire106 = ( i_7_  &  i_6_  &  n_n7  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n1 ) ;
 assign wire133 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n19  &  n_n9 ) ;
 assign wire138 = ( n_n1256 ) | ( wire127 ) | ( n_n797 ) | ( wire3363 ) ;
 assign wire140 = ( wire113 ) | ( n_n19  &  wire71 ) ;
 assign wire216 = ( wire249 ) | ( n_n792 ) | ( wire493 ) ;
 assign wire174 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n12 ) ;
 assign wire412 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) ;
 assign wire413 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n11 ) ;
 assign wire414 = ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n3 ) ;
 assign wire421 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign wire426 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n18 ) ;
 assign wire434 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign wire450 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign wire456 = ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n9 ) ;
 assign wire461 = ( i_7_  &  i_6_  &  wire93 ) | ( (~ i_7_)  &  i_6_  &  wire93 ) | ( i_7_  &  i_6_  &  wire466 ) | ( (~ i_7_)  &  i_6_  &  wire466 ) ;
 assign wire462 = ( wire93  &  n_n10 ) | ( n_n10  &  wire466 ) ;
 assign wire466 = ( n_n6  &  n_n10 ) | ( n_n6  &  n_n9  &  wire64 ) ;
 assign wire468 = ( (~ i_7_)  &  (~ i_6_)  &  n_n6  &  n_n13 ) ;
 assign wire471 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n10 ) ;
 assign wire473 = ( i_7_  &  i_6_  &  n_n19  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n10 ) ;
 assign wire476 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire483 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n9 ) ;
 assign wire487 = ( i_7_  &  i_6_  &  n_n10  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n10  &  n_n1 ) ;
 assign wire488 = ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign wire493 = ( i_7_  &  i_6_  &  n_n0  &  n_n18 ) ;
 assign wire500 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n18 ) ;
 assign wire504 = ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n9 ) ;
 assign wire505 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) ;
 assign wire507 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign wire512 = ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire515 = ( i_7_  &  (~ i_6_)  &  n_n19  &  n_n12 ) ;
 assign wire532 = ( n_n6  &  n_n10 ) | ( n_n6  &  n_n9  &  wire64 ) ;
 assign wire534 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n13 ) ;
 assign wire545 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n10 ) ;
 assign wire546 = ( i_7_  &  i_6_  &  n_n3  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n9 ) ;
 assign wire549 = ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n10 ) ;
 assign wire551 = ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire561 = ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) ;
 assign wire564 = ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n13 ) ;
 assign wire568 = ( i_7_  &  i_6_  &  n_n10  &  n_n1 ) ;
 assign wire588 = ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n2 ) ;
 assign wire592 = ( i_7_  &  i_6_  &  n_n4  &  n_n18 ) ;
 assign wire3176 = ( (~ i_5_)  &  i_3_  &  i_4_  &  n_n14 ) | ( (~ i_5_)  &  (~ i_3_)  &  i_4_  &  n_n14 ) ;
 assign wire3177 = ( n_n11  &  n_n14 ) | ( n_n7  &  n_n5  &  n_n14 ) ;
 assign wire3178 = ( n_n7  &  n_n6  &  n_n14 ) | ( n_n7  &  n_n3  &  n_n14 ) ;
 assign wire3179 = ( n_n0  &  n_n7  &  n_n14 ) | ( n_n7  &  n_n4  &  n_n14 ) ;
 assign wire3180 = ( n_n7  &  n_n2  &  n_n14 ) | ( n_n7  &  n_n19  &  n_n14 ) ;
 assign wire3184 = ( n_n1305 ) | ( wire3176 ) | ( wire3177 ) | ( wire3178 ) ;
 assign wire3188 = ( n_n5  &  n_n8  &  n_n14 ) | ( n_n19  &  n_n8  &  n_n14 ) ;
 assign wire3189 = ( n_n4  &  n_n8  &  n_n14 ) | ( n_n2  &  n_n8  &  n_n14 ) ;
 assign wire3190 = ( n_n0  &  n_n8  &  n_n14 ) | ( n_n1  &  n_n8  &  n_n14 ) ;
 assign wire3191 = ( n_n6  &  n_n8  &  n_n14 ) | ( n_n3  &  n_n8  &  n_n14 ) ;
 assign wire3195 = ( i_7_  &  (~ i_6_)  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11 ) ;
 assign wire3196 = ( n_n4  &  n_n11  &  wire66 ) | ( n_n11  &  wire66  &  n_n1 ) ;
 assign wire3203 = ( n_n1168 ) | ( n_n1321 ) | ( wire3196 ) ;
 assign wire3204 = ( o_20_ ) | ( n_n1010 ) | ( wire135 ) | ( n_n1320 ) ;
 assign wire3205 = ( n_n1169 ) | ( wire73 ) | ( wire92 ) | ( wire93 ) ;
 assign wire3206 = ( wire94 ) | ( wire146 ) | ( wire147 ) | ( wire186 ) ;
 assign wire3209 = ( wire208 ) | ( wire249 ) | ( wire3203 ) | ( wire3206 ) ;
 assign wire3210 = ( o_21_ ) | ( n_n1197 ) | ( n_n953 ) ;
 assign wire3213 = ( i_7_  &  i_6_  &  n_n19  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n19  &  n_n8 ) ;
 assign wire3216 = ( n_n1013 ) | ( n_n0  &  wire72 ) ;
 assign wire3217 = ( n_n845 ) | ( n_n858 ) ;
 assign wire3218 = ( i_7_  &  i_6_  &  n_n1  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n8 ) ;
 assign wire3221 = ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n3 ) ;
 assign wire3222 = ( o_15_ ) | ( n_n1215 ) | ( n_n1216 ) | ( wire561 ) ;
 assign wire3225 = ( wire180 ) | ( n_n4  &  n_n11  &  wire66 ) ;
 assign wire3236 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign wire3237 = ( n_n1238 ) | ( n_n1239 ) | ( n_n937 ) ;
 assign wire3238 = ( wire246 ) | ( wire109 ) | ( n_n1243 ) | ( wire3236 ) ;
 assign wire3239 = ( n_n6  &  n_n13 ) | ( n_n6  &  n_n17  &  n_n12 ) ;
 assign wire3243 = ( n_n1009 ) | ( n_n4  &  wire67  &  n_n18 ) ;
 assign wire3244 = ( n_n1135 ) | ( n_n1134 ) | ( n_n1137 ) | ( n_n1136 ) ;
 assign wire3245 = ( o_7_ ) | ( wire186 ) | ( n_n1120 ) | ( wire592 ) ;
 assign wire3248 = ( wire93 ) | ( n_n872 ) | ( wire159 ) | ( wire219 ) ;
 assign wire3250 = ( n_n1008 ) | ( n_n1203 ) | ( wire273 ) | ( wire3210 ) ;
 assign wire3251 = ( wire354 ) | ( wire92 ) | ( wire222 ) | ( wire160 ) ;
 assign wire3255 = ( n_n949 ) | ( wire162 ) | ( wire243 ) | ( wire3245 ) ;
 assign wire3256 = ( wire187 ) | ( wire226 ) | ( wire3248 ) ;
 assign wire3257 = ( n_n936 ) | ( wire295 ) | ( wire3243 ) | ( wire3244 ) ;
 assign wire3261 = ( wire228 ) | ( wire99 ) | ( wire191 ) | ( wire3251 ) ;
 assign wire3262 = ( wire280 ) | ( wire327 ) | ( wire331 ) | ( wire346 ) ;
 assign wire3264 = ( wire301 ) | ( n_n387 ) | ( wire3237 ) | ( wire3238 ) ;
 assign wire3266 = ( wire240 ) | ( wire252 ) | ( wire324 ) | ( wire3250 ) ;
 assign wire3267 = ( wire3262 ) | ( wire3261 ) ;
 assign wire3268 = ( wire332 ) | ( wire3217 ) | ( wire3255 ) | ( wire3256 ) ;
 assign wire3269 = ( wire115 ) | ( wire192 ) | ( wire3257 ) | ( wire3264 ) ;
 assign wire3273 = ( i_7_  &  i_6_  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire3274 = ( wire133 ) | ( n_n17  &  n_n19  &  n_n8 ) ;
 assign wire3277 = ( o_11_ ) | ( n_n5  &  n_n17  &  n_n18 ) ;
 assign wire3278 = ( n_n5  &  n_n12  &  n_n16 ) | ( n_n5  &  n_n16  &  n_n18 ) ;
 assign wire3279 = ( n_n1163 ) | ( wire564 ) | ( wire3278 ) ;
 assign wire3282 = ( n_n1009 ) | ( n_n19  &  n_n15  &  n_n12 ) ;
 assign wire3283 = ( n_n756 ) | ( n_n1104 ) | ( wire236 ) ;
 assign wire3285 = ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n11 ) | ( i_7_  &  (~ i_6_)  &  n_n6  &  n_n11 ) ;
 assign wire3286 = ( o_28_ ) | ( n_n1165 ) | ( wire78 ) ;
 assign wire3287 = ( n_n1169 ) | ( n_n1170 ) | ( n_n826 ) | ( wire3285 ) ;
 assign wire3288 = ( wire297 ) | ( wire3279 ) | ( wire3286 ) ;
 assign wire3290 = ( n_n1009 ) | ( n_n786 ) | ( wire515 ) | ( wire3283 ) ;
 assign wire3292 = ( wire337 ) | ( wire323 ) | ( wire3277 ) | ( wire3287 ) ;
 assign wire3294 = ( i_7_  &  i_6_  &  n_n4  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n8 ) ;
 assign wire3296 = ( n_n906 ) | ( n_n1329 ) | ( n_n910 ) | ( n_n909 ) ;
 assign wire3299 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign wire3304 = ( i_7_  &  i_6_  &  n_n0  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n12 ) ;
 assign wire3305 = ( i_7_  &  i_6_  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign wire3309 = ( n_n1302 ) | ( n_n553 ) | ( wire106 ) ;
 assign wire3311 = ( i_7_  &  i_6_  &  n_n11  &  n_n1 ) | ( (~ i_7_)  &  i_6_  &  n_n11  &  n_n1 ) | ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n1 ) ;
 assign wire3312 = ( i_7_  &  i_6_  &  n_n2  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n10 ) ;
 assign wire3313 = ( n_n4  &  n_n10 ) | ( n_n4  &  n_n11  &  wire66 ) ;
 assign wire3316 = ( n_n4  &  n_n8  &  n_n15 ) | ( n_n4  &  n_n15  &  n_n12 ) ;
 assign wire3317 = ( o_20_ ) | ( n_n2  &  wire69 ) ;
 assign wire3318 = ( n_n1029 ) | ( n_n1  &  wire70 ) ;
 assign wire3319 = ( wire3313 ) | ( wire184 ) ;
 assign wire3320 = ( n_n1211 ) | ( n_n1193 ) | ( n_n1225 ) | ( n_n1197 ) ;
 assign wire3321 = ( o_14_ ) | ( n_n1192 ) | ( wire534 ) | ( wire3316 ) ;
 assign wire3322 = ( n_n1028 ) | ( wire512 ) | ( wire3294 ) ;
 assign wire3327 = ( n_n935 ) | ( wire77 ) | ( n_n1213 ) | ( wire3322 ) ;
 assign wire3328 = ( wire3317 ) | ( wire3318 ) | ( wire3319 ) | ( wire3320 ) ;
 assign wire3329 = ( wire218 ) | ( wire348 ) | ( wire3321 ) ;
 assign wire3332 = ( wire3327 ) | ( wire3328 ) | ( wire3329 ) ;
 assign wire3333 = ( n_n137 ) | ( wire200 ) | ( wire150 ) | ( wire148 ) ;
 assign wire3334 = ( wire330 ) | ( wire326 ) | ( wire221 ) | ( wire165 ) ;
 assign wire3340 = ( i_7_  &  i_6_  &  n_n6  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n6  &  n_n12 ) ;
 assign wire3341 = ( n_n1135 ) | ( n_n1134 ) | ( n_n1136 ) ;
 assign wire3342 = ( n_n973 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3344 = ( wire461 ) | ( wire3341 ) | ( wire3342 ) ;
 assign wire3345 = ( n_n904 ) | ( wire308 ) | ( wire462 ) ;
 assign wire3348 = ( n_n1147 ) | ( n_n1153 ) | ( wire160 ) | ( wire456 ) ;
 assign wire3349 = ( i_7_  &  i_6_  &  n_n5  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n12 ) ;
 assign wire3350 = ( n_n1154 ) | ( n_n1169 ) | ( n_n1170 ) ;
 assign wire3351 = ( o_28_ ) | ( wire286 ) | ( wire78 ) | ( n_n1166 ) ;
 assign wire3353 = ( wire222 ) | ( wire3348 ) | ( wire3351 ) ;
 assign wire3355 = ( n_n427 ) | ( n_n609 ) | ( wire3350 ) | ( wire3353 ) ;
 assign wire3358 = ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n12 ) ;
 assign wire3359 = ( wire135 ) | ( n_n805 ) ;
 assign wire3360 = ( wire189 ) | ( wire218 ) ;
 assign wire3361 = ( n_n1244 ) | ( n_n2  &  wire70 ) ;
 assign wire3363 = ( (~ i_7_)  &  i_6_  &  n_n13  &  n_n2 ) | ( i_7_  &  (~ i_6_)  &  n_n13  &  n_n2 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n13  &  n_n2 ) ;
 assign wire3366 = ( wire88 ) | ( n_n2  &  n_n10  &  wire67 ) ;
 assign wire3367 = ( n_n1194 ) | ( n_n1261 ) | ( n_n1010 ) | ( n_n1320 ) ;
 assign wire3368 = ( wire147 ) | ( n_n616 ) | ( wire274 ) | ( wire242 ) ;
 assign wire3369 = ( n_n1321 ) | ( wire265 ) | ( wire3216 ) | ( wire3366 ) ;
 assign wire3370 = ( n_n602 ) | ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) ;
 assign wire3373 = ( n_n1334 ) | ( wire83 ) | ( wire85 ) | ( wire128 ) ;
 assign wire3375 = ( wire114 ) | ( wire298 ) | ( wire3367 ) | ( wire3368 ) ;
 assign wire3377 = ( wire3369 ) | ( wire3370 ) | ( wire3373 ) ;
 assign wire3378 = ( wire218 ) | ( wire189 ) | ( wire238 ) | ( wire3375 ) ;
 assign wire3379 = ( n_n573 ) | ( wire318 ) | ( wire319 ) ;
 assign wire3381 = ( wire3344 ) | ( wire3345 ) | ( wire3355 ) | ( wire3379 ) ;
 assign wire3383 = ( n_n1257 ) | ( n_n13  &  n_n2  &  wire64 ) ;
 assign wire3384 = ( i_7_  &  i_6_  &  n_n1  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n1  &  n_n18 ) ;
 assign wire3387 = ( wire146 ) | ( n_n3  &  wire72 ) ;
 assign wire3388 = ( n_n1238 ) | ( wire268 ) | ( n_n1239 ) | ( wire434 ) ;
 assign wire3390 = ( (~ i_7_)  &  i_6_  &  n_n1  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n1  &  n_n8 ) ;
 assign wire3393 = ( wire249 ) | ( wire183 ) | ( wire207 ) | ( wire426 ) ;
 assign wire3395 = ( (~ i_7_)  &  i_6_  &  n_n0  &  n_n13 ) | ( i_7_  &  (~ i_6_)  &  n_n0  &  n_n13 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n0  &  n_n13 ) ;
 assign wire3400 = ( i_7_  &  i_6_  &  n_n11  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n11  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n11  &  n_n19 ) ;
 assign wire3404 = ( n_n921 ) | ( n_n1  &  wire71 ) | ( n_n1  &  wire3195 ) ;
 assign wire3405 = ( o_21_ ) | ( n_n1168 ) | ( n_n1196 ) | ( n_n953 ) ;
 assign wire3406 = ( n_n1287 ) | ( n_n1163 ) | ( n_n1318 ) | ( n_n1189 ) ;
 assign wire3407 = ( n_n756 ) | ( n_n1135 ) | ( n_n1203 ) | ( wire273 ) ;
 assign wire3408 = ( n_n1049 ) | ( n_n1227 ) | ( wire3358 ) ;
 assign wire3410 = ( wire93 ) | ( wire186 ) | ( wire3400 ) ;
 assign wire3411 = ( n_n1009 ) | ( n_n864 ) | ( n_n1061 ) | ( n_n1083 ) ;
 assign wire3413 = ( wire3407 ) | ( wire3406 ) ;
 assign wire3414 = ( wire297 ) | ( wire309 ) | ( wire3408 ) ;
 assign wire3417 = ( n_n845 ) | ( wire129 ) | ( wire107 ) | ( wire128 ) ;
 assign wire3418 = ( wire337 ) | ( n_n1015 ) | ( n_n1320 ) | ( wire3216 ) ;
 assign wire3420 = ( wire345 ) | ( wire3383 ) | ( wire3410 ) | ( wire3411 ) ;
 assign wire3422 = ( wire324 ) | ( wire343 ) | ( wire3404 ) | ( wire3405 ) ;
 assign wire3424 = ( n_n573 ) | ( n_n574 ) | ( wire3413 ) | ( wire3414 ) ;
 assign wire3425 = ( wire3420 ) | ( wire333 ) ;
 assign wire3428 = ( wire285 ) | ( wire341 ) | ( wire3422 ) | ( wire3425 ) ;
 assign wire3430 = ( wire129 ) | ( wire107 ) | ( n_n582 ) ;
 assign wire3432 = ( wire228 ) | ( n_n1231 ) | ( wire135 ) ;
 assign wire3433 = ( n_n1169 ) | ( n_n1147 ) | ( n_n1170 ) | ( wire549 ) ;
 assign wire3434 = ( wire354 ) | ( wire92 ) | ( wire222 ) | ( wire160 ) ;
 assign wire3435 = ( wire93 ) | ( wire466 ) | ( wire3433 ) ;
 assign wire3436 = ( wire187 ) | ( wire99 ) | ( wire191 ) | ( wire3434 ) ;
 assign wire3437 = ( wire88 ) | ( n_n5  &  wire72 ) ;
 assign wire3439 = ( n_n1203 ) | ( wire194 ) | ( wire273 ) | ( wire3210 ) ;
 assign wire3440 = ( wire320 ) | ( n_n955 ) | ( wire3437 ) ;
 assign wire3441 = ( wire155 ) | ( n_n0  &  n_n11  &  n_n16 ) ;
 assign wire3442 = ( n_n1135 ) | ( n_n1134 ) | ( n_n1137 ) ;
 assign wire3443 = ( n_n973 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3446 = ( wire155 ) | ( n_n1319 ) | ( n_n911 ) | ( wire3443 ) ;
 assign wire3447 = ( n_n936 ) | ( wire261 ) | ( wire295 ) | ( wire3442 ) ;
 assign wire3448 = ( n_n904 ) | ( n_n906 ) | ( n_n1329 ) | ( wire128 ) ;
 assign wire3452 = ( n_n996 ) | ( wire87 ) | ( wire3446 ) | ( wire3448 ) ;
 assign wire3453 = ( wire343 ) | ( wire201 ) | ( wire3430 ) | ( wire3432 ) ;
 assign wire3454 = ( wire3435 ) | ( wire3436 ) | ( wire3439 ) | ( wire3440 ) ;
 assign wire3455 = ( wire330 ) | ( n_n427 ) | ( wire200 ) | ( wire3447 ) ;
 assign wire3458 = ( o_13_ ) | ( n_n1254 ) | ( n_n1253 ) ;
 assign wire3460 = ( wire292 ) | ( n_n1230 ) | ( n_n1040 ) | ( wire3458 ) ;
 assign wire3462 = ( wire248 ) | ( n_n0  &  wire82 ) | ( n_n0  &  wire71 ) ;
 assign wire3464 = ( n_n744 ) | ( wire153 ) | ( wire155 ) ;
 assign wire3465 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign wire3467 = ( o_15_ ) | ( n_n1223 ) | ( wire414 ) ;
 assign wire3470 = ( i_7_  &  i_6_  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n10 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n10 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n10 ) ;
 assign wire3471 = ( o_21_ ) | ( n_n1255 ) | ( n_n1256 ) | ( n_n1229 ) ;
 assign wire3472 = ( n_n1029 ) | ( wire3470 ) | ( n_n1  &  wire70 ) ;
 assign wire3474 = ( n_n1197 ) | ( wire88 ) | ( n_n845 ) | ( n_n955 ) ;
 assign wire3475 = ( n_n602 ) | ( n_n1022 ) | ( n_n1023 ) | ( wire3472 ) ;
 assign wire3477 = ( wire298 ) | ( wire84 ) | ( wire216 ) | ( wire3471 ) ;
 assign wire3480 = ( wire189 ) | ( wire310 ) | ( wire3477 ) ;
 assign wire3481 = ( wire221 ) | ( wire165 ) | ( wire181 ) | ( wire3460 ) ;
 assign wire3482 = ( wire177 ) | ( wire182 ) | ( wire3474 ) | ( wire3475 ) ;
 assign wire3485 = ( o_20_ ) | ( n_n4  &  n_n8  &  n_n15 ) ;
 assign wire3486 = ( n_n1211 ) | ( wire279 ) | ( wire512 ) | ( wire3294 ) ;
 assign wire3487 = ( n_n13 ) | ( n_n7  &  n_n2  &  n_n14 ) ;
 assign wire3488 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n12 ) ;
 assign wire3491 = ( n_n1229 ) | ( n_n1056 ) | ( wire3488 ) ;
 assign wire3492 = ( wire155 ) | ( wire3304 ) | ( wire3305 ) | ( wire3487 ) ;
 assign wire3493 = ( wire153 ) | ( n_n1283 ) | ( n_n580 ) | ( wire260 ) ;
 assign wire3494 = ( wire164 ) | ( n_n955 ) | ( wire3225 ) | ( wire3491 ) ;
 assign wire3495 = ( n_n845 ) | ( wire128 ) | ( wire3485 ) | ( wire3486 ) ;
 assign wire3496 = ( wire87 ) | ( n_n1032 ) | ( wire216 ) | ( wire3309 ) ;
 assign wire3497 = ( n_n996 ) | ( wire150 ) | ( wire148 ) | ( n_n1257 ) ;
 assign wire3498 = ( wire3493 ) | ( wire3492 ) ;
 assign wire3502 = ( wire181 ) | ( wire3460 ) | ( wire3494 ) | ( wire3495 ) ;
 assign wire3503 = ( wire318 ) | ( wire3496 ) | ( wire3497 ) | ( wire3498 ) ;
 assign wire3505 = ( n_n4  &  n_n17  &  n_n8 ) | ( n_n2  &  n_n17  &  n_n8 ) ;
 assign wire3506 = ( n_n805 ) | ( n_n3  &  wire71 ) ;
 assign wire3507 = ( wire104 ) | ( wire412 ) | ( wire413 ) ;
 assign wire3510 = ( o_20_ ) | ( wire135 ) | ( wire3505 ) ;
 assign wire3511 = ( n_n1028 ) | ( n_n930 ) | ( n_n2  &  wire72 ) ;
 assign wire3515 = ( wire159 ) | ( wire162 ) | ( wire288 ) | ( wire293 ) ;
 assign wire3516 = ( wire331 ) | ( n_n797 ) | ( wire3363 ) ;
 assign wire3517 = ( wire95 ) | ( wire3467 ) | ( wire3510 ) ;
 assign wire3518 = ( n_n950 ) | ( wire77 ) | ( n_n1213 ) | ( wire3511 ) ;
 assign wire3519 = ( n_n803 ) | ( wire164 ) | ( wire3506 ) | ( wire3507 ) ;
 assign wire3520 = ( n_n602 ) | ( n_n1022 ) | ( n_n1023 ) | ( wire3515 ) ;
 assign wire3521 = ( wire310 ) | ( wire216 ) | ( wire3304 ) | ( wire3305 ) ;
 assign wire3526 = ( wire178 ) | ( wire270 ) | ( n_n823 ) | ( wire3521 ) ;
 assign wire3527 = ( wire3516 ) | ( wire3517 ) | ( wire3518 ) | ( wire3519 ) ;
 assign wire3528 = ( wire301 ) | ( n_n137 ) | ( wire3520 ) ;
 assign wire3533 = ( wire77 ) | ( n_n3  &  wire72 ) ;
 assign wire3535 = ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign wire3541 = ( wire94 ) | ( n_n1  &  wire71 ) ;
 assign wire3542 = ( o_6_ ) | ( n_n921 ) | ( n_n5  &  wire72 ) ;
 assign wire3545 = ( n_n1274 ) | ( n_n1121 ) | ( n_n1180 ) | ( n_n1321 ) ;
 assign wire3546 = ( n_n814 ) | ( n_n1122 ) | ( n_n1288 ) | ( n_n1204 ) ;
 assign wire3548 = ( n_n1287 ) | ( n_n822 ) | ( n_n1285 ) | ( wire243 ) ;
 assign wire3552 = ( wire76 ) | ( wire130 ) | ( wire274 ) | ( wire291 ) ;
 assign wire3554 = ( wire86 ) | ( wire95 ) | ( wire3467 ) ;
 assign wire3556 = ( n_n1049 ) | ( n_n1010 ) | ( n_n1320 ) | ( wire3548 ) ;
 assign wire3557 = ( wire111 ) | ( wire136 ) | ( wire253 ) | ( wire276 ) ;
 assign wire3558 = ( wire3541 ) | ( wire3542 ) | ( wire3552 ) ;
 assign wire3560 = ( wire87 ) | ( wire215 ) | ( n_n1032 ) | ( wire3533 ) ;
 assign wire3561 = ( wire345 ) | ( wire229 ) | ( n_n642 ) ;
 assign wire3566 = ( wire196 ) | ( wire3545 ) | ( wire3546 ) | ( wire3560 ) ;
 assign wire3567 = ( wire154 ) | ( wire305 ) | ( wire3554 ) | ( wire3561 ) ;
 assign wire3568 = ( wire3435 ) | ( wire3436 ) | ( wire3556 ) | ( wire3557 ) ;
 assign wire3569 = ( wire341 ) | ( n_n427 ) | ( n_n1006 ) | ( wire3558 ) ;
 assign wire3573 = ( i_7_  &  i_6_  &  n_n4  &  n_n12 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n12 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n12 ) ;
 assign wire3577 = ( n_n19  &  wire163 ) | ( n_n19  &  n_n10  &  wire64 ) ;
 assign wire3579 = ( wire133 ) | ( n_n19  &  n_n8  &  n_n14 ) ;
 assign wire3581 = ( n_n953 ) | ( (~ n_n17) ) | ( n_n4  &  n_n13  &  n_n17 ) ;
 assign wire3582 = ( n_n961 ) | ( n_n962 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3585 = ( n_n128 ) | ( n_n859 ) | ( n_n5  &  wire72 ) ;
 assign wire3586 = ( n_n1083 ) | ( wire156 ) | ( wire236 ) | ( wire3577 ) ;
 assign wire3587 = ( n_n1121 ) | ( wire133 ) | ( wire140 ) | ( wire3582 ) ;
 assign wire3588 = ( wire276 ) | ( wire83 ) | ( wire85 ) | ( wire3581 ) ;
 assign wire3589 = ( n_n602 ) | ( n_n215 ) | ( n_n1022 ) | ( n_n1023 ) ;
 assign wire3590 = ( wire215 ) | ( wire3485 ) | ( wire3486 ) | ( wire3533 ) ;
 assign wire3592 = ( wire348 ) | ( n_n1002 ) | ( wire95 ) | ( wire3467 ) ;
 assign wire3598 = ( wire345 ) | ( wire229 ) | ( n_n642 ) | ( wire3592 ) ;
 assign wire3599 = ( wire221 ) | ( wire165 ) | ( wire3585 ) | ( wire3586 ) ;
 assign wire3600 = ( wire193 ) | ( wire255 ) | ( wire313 ) | ( wire3587 ) ;
 assign wire3601 = ( wire332 ) | ( wire3588 ) | ( wire3589 ) | ( wire3590 ) ;
 assign wire3604 = ( wire180 ) | ( wire273 ) ;
 assign wire3605 = ( n_n1197 ) | ( wire88 ) | ( n_n955 ) | ( wire3604 ) ;
 assign wire3607 = ( wire295 ) | ( wire290 ) | ( n_n2  &  wire69 ) ;
 assign wire3609 = ( n_n1010 ) | ( wire208 ) ;
 assign wire3610 = ( n_n1283 ) | ( n_n1334 ) | ( n_n580 ) ;
 assign wire3612 = ( wire331 ) | ( n_n931 ) | ( wire3609 ) | ( wire3610 ) ;
 assign wire3613 = ( n_n95 ) | ( n_n858 ) | ( wire3462 ) | ( wire3464 ) ;
 assign wire3614 = ( wire200 ) | ( wire150 ) | ( wire148 ) | ( wire3612 ) ;
 assign wire3615 = ( wire343 ) | ( wire211 ) | ( wire3432 ) | ( wire3607 ) ;
 assign wire3616 = ( wire318 ) | ( wire3605 ) | ( wire3613 ) ;
 assign wire3618 = ( wire3344 ) | ( wire3345 ) | ( wire3355 ) | ( wire3616 ) ;
 assign wire3619 = ( n_n0  &  n_n18 ) | ( n_n0  &  n_n17  &  n_n12 ) ;
 assign wire3621 = ( n_n1  &  wire71 ) | ( n_n11  &  n_n1  &  n_n16 ) ;
 assign wire3623 = ( n_n1010 ) | ( wire279 ) | ( n_n17  &  n_n9 ) ;
 assign wire3624 = ( wire153 ) | ( n_n950 ) | ( n_n1208 ) | ( wire551 ) ;
 assign wire3628 = ( o_18_ ) | ( wire130 ) | ( wire237 ) | ( wire3624 ) ;
 assign wire3630 = ( wire218 ) | ( wire238 ) | ( wire3623 ) ;
 assign wire3631 = ( wire179 ) | ( wire139 ) | ( wire3393 ) | ( wire3628 ) ;
 assign wire3632 = ( n_n573 ) | ( wire319 ) | ( n_n990 ) | ( n_n574 ) ;
 assign wire3635 = ( n_n883 ) | ( wire3355 ) | ( wire3630 ) | ( wire3631 ) ;
 assign wire3636 = ( i_7_  &  i_6_  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  i_6_  &  n_n4  &  n_n9 ) | ( i_7_  &  (~ i_6_)  &  n_n4  &  n_n9 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n4  &  n_n9 ) ;
 assign wire3638 = ( i_7_  &  i_6_  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  i_6_  &  n_n3  &  n_n18 ) | ( i_7_  &  (~ i_6_)  &  n_n3  &  n_n18 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n3  &  n_n18 ) ;
 assign wire3639 = ( wire3638 ) | ( n_n13  &  n_n3  &  wire64 ) ;
 assign wire3641 = ( wire197 ) | ( wire154 ) ;
 assign wire3643 = ( wire146 ) | ( n_n1  &  wire67  &  n_n18 ) ;
 assign wire3644 = ( wire183 ) | ( n_n0  &  wire69 ) ;
 assign wire3645 = ( wire300 ) | ( wire247 ) ;
 assign wire3652 = ( wire226 ) | ( n_n1300 ) | ( n_n1258 ) | ( wire257 ) ;
 assign wire3653 = ( n_n1018 ) | ( n_n1022 ) | ( wire3643 ) | ( wire3644 ) ;
 assign wire3654 = ( n_n215 ) | ( wire250 ) | ( n_n923 ) | ( wire3621 ) ;
 assign wire3655 = ( wire228 ) | ( wire230 ) | ( n_n387 ) | ( wire3645 ) ;
 assign wire3658 = ( wire254 ) | ( n_n1275 ) | ( wire132 ) | ( wire3654 ) ;
 assign wire3659 = ( wire83 ) | ( wire229 ) | ( wire3652 ) | ( wire3655 ) ;
 assign wire3660 = ( wire177 ) | ( wire332 ) | ( wire3641 ) | ( wire3653 ) ;
 assign wire3663 = ( n_n883 ) | ( wire3355 ) | ( wire3658 ) | ( wire3659 ) ;
 assign wire3667 = ( n_n1122 ) | ( n_n1165 ) | ( wire78 ) ;
 assign wire3668 = ( n_n1137 ) | ( n_n962 ) | ( wire468 ) | ( wire3340 ) ;
 assign wire3669 = ( n_n864 ) | ( wire158 ) | ( wire316 ) ;
 assign wire3671 = ( wire297 ) | ( n_n963 ) | ( n_n859 ) | ( wire3279 ) ;
 assign wire3672 = ( wire93 ) | ( wire140 ) | ( wire466 ) | ( wire3274 ) ;
 assign wire3674 = ( n_n128 ) | ( wire3282 ) | ( wire3283 ) | ( wire3667 ) ;
 assign wire3676 = ( wire152 ) | ( n_n673 ) | ( wire3668 ) | ( wire3669 ) ;
 assign wire3679 = ( n_n4  &  n_n15  &  n_n12 ) | ( n_n2  &  n_n15  &  n_n12 ) ;
 assign wire3682 = ( n_n1  &  wire71 ) | ( n_n10  &  n_n1  &  wire64 ) ;
 assign wire3686 = ( n_n1300 ) | ( n_n1238 ) | ( n_n1239 ) | ( n_n1315 ) ;
 assign wire3687 = ( o_9_ ) | ( wire259 ) | ( n_n1301 ) ;
 assign wire3688 = ( o_13_ ) | ( o_7_ ) | ( n_n1253 ) | ( n_n1268 ) ;
 assign wire3689 = ( o_6_ ) | ( n_n1225 ) | ( wire3679 ) ;
 assign wire3690 = ( n_n1334 ) | ( n_n1254 ) | ( n_n1330 ) | ( n_n1316 ) ;
 assign wire3691 = ( n_n1028 ) | ( wire77 ) | ( n_n1213 ) ;
 assign wire3692 = ( n_n1197 ) | ( wire88 ) | ( n_n822 ) ;
 assign wire3693 = ( wire183 ) | ( n_n813 ) | ( wire207 ) ;
 assign wire3695 = ( n_n1010 ) | ( n_n961 ) | ( wire109 ) | ( wire112 ) ;
 assign wire3702 = ( wire159 ) | ( wire162 ) | ( wire3682 ) | ( wire3693 ) ;
 assign wire3703 = ( wire3686 ) | ( wire3687 ) | ( wire3695 ) ;
 assign wire3704 = ( wire218 ) | ( wire3688 ) | ( wire3689 ) ;
 assign wire3705 = ( wire305 ) | ( n_n387 ) | ( n_n642 ) | ( wire3690 ) ;
 assign wire3706 = ( n_n574 ) | ( wire254 ) | ( wire3691 ) | ( wire3692 ) ;
 assign wire3710 = ( wire314 ) | ( wire3702 ) | ( wire3703 ) | ( wire3704 ) ;
 assign wire3712 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n19 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n19 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n19 ) ;
 assign wire3713 = ( n_n1135 ) | ( n_n1137 ) | ( wire3712 ) ;
 assign wire3714 = ( i_7_  &  i_6_  &  n_n7  &  n_n2 ) | ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n2 ) ;
 assign wire3715 = ( wire269 ) | ( wire3714 ) ;
 assign wire3716 = ( o_18_ ) | ( wire130 ) | ( n_n1033 ) ;
 assign wire3717 = ( wire250 ) | ( n_n923 ) | ( wire3621 ) | ( wire3715 ) ;
 assign wire3719 = ( o_30_ ) | ( o_7_ ) | ( wire127 ) ;
 assign wire3722 = ( n_n1121 ) | ( wire257 ) | ( wire133 ) | ( wire140 ) ;
 assign wire3723 = ( n_n1049 ) | ( wire99 ) | ( wire235 ) | ( wire77 ) ;
 assign wire3724 = ( wire189 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire3725 = ( n_n673 ) | ( n_n1076 ) | ( n_n1136 ) | ( wire3713 ) ;
 assign wire3730 = ( wire197 ) | ( wire325 ) | ( wire3725 ) ;
 assign wire3731 = ( wire284 ) | ( n_n660 ) | ( wire3719 ) | ( wire3722 ) ;
 assign wire3732 = ( wire315 ) | ( wire3716 ) | ( wire3717 ) ;
 assign wire3733 = ( wire255 ) | ( n_n563 ) | ( wire3723 ) | ( wire3724 ) ;
 assign wire3736 = ( n_n906 ) | ( n_n1017 ) ;
 assign wire3739 = ( wire196 ) | ( n_n1022 ) | ( wire223 ) | ( n_n1023 ) ;
 assign wire3743 = ( wire333 ) | ( wire177 ) | ( wire154 ) | ( wire197 ) ;
 assign wire3744 = ( wire86 ) | ( wire193 ) | ( wire267 ) | ( wire3736 ) ;
 assign wire3745 = ( wire314 ) | ( wire141 ) | ( wire165 ) | ( wire3739 ) ;
 assign wire3749 = ( wire108 ) | ( wire337 ) | ( wire3435 ) | ( wire3436 ) ;
 assign wire3750 = ( n_n1022 ) | ( n_n1023 ) | ( n_n1024 ) | ( n_n1025 ) ;
 assign wire3751 = ( wire298 ) | ( n_n1021 ) | ( n_n1020 ) | ( wire303 ) ;
 assign wire3754 = ( n_n1029 ) | ( n_n1017 ) | ( n_n1  &  wire70 ) ;
 assign wire3756 = ( n_n845 ) | ( wire209 ) | ( wire292 ) ;
 assign wire3758 = ( n_n1215 ) | ( n_n744 ) | ( n_n745 ) | ( wire3754 ) ;
 assign wire3759 = ( n_n895 ) | ( n_n858 ) | ( wire3462 ) ;
 assign wire3760 = ( wire85 ) | ( wire283 ) | ( wire3756 ) ;
 assign wire3763 = ( wire3439 ) | ( wire3440 ) | ( wire3760 ) ;
 assign wire3764 = ( wire267 ) | ( wire3750 ) | ( wire3751 ) ;
 assign wire3765 = ( wire165 ) | ( wire181 ) | ( wire3758 ) | ( wire3759 ) ;
 assign wire3767 = ( wire285 ) | ( wire284 ) | ( wire3749 ) | ( wire3765 ) ;
 assign wire3770 = ( (~ i_7_)  &  i_6_  &  n_n2  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n8 ) ;
 assign wire3772 = ( o_7_ ) | ( n_n554 ) | ( n_n1268 ) ;
 assign wire3774 = ( n_n1271 ) | ( n_n1189 ) | ( n_n1  &  wire72 ) ;
 assign wire3775 = ( n_n1216 ) | ( n_n1244 ) | ( wire3770 ) ;
 assign wire3777 = ( wire186 ) | ( n_n1061 ) | ( wire209 ) | ( n_n1223 ) ;
 assign wire3781 = ( n_n1245 ) | ( wire287 ) | ( wire308 ) | ( wire277 ) ;
 assign wire3782 = ( n_n810 ) | ( n_n809 ) | ( wire3772 ) | ( wire3777 ) ;
 assign wire3784 = ( n_n904 ) | ( wire129 ) | ( wire107 ) ;
 assign wire3786 = ( wire112 ) | ( wire150 ) | ( n_n802 ) | ( wire3781 ) ;
 assign wire3789 = ( wire324 ) | ( wire3774 ) | ( wire3775 ) | ( wire3784 ) ;
 assign wire3790 = ( wire342 ) | ( wire3341 ) | ( wire3342 ) | ( wire3786 ) ;
 assign wire3792 = ( n_n427 ) | ( wire340 ) | ( wire3782 ) ;
 assign wire3795 = ( wire200 ) | ( wire238 ) | ( wire3789 ) | ( wire3792 ) ;
 assign wire3796 = ( i_7_  &  i_6_  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  i_6_  &  n_n5  &  n_n8 ) | ( i_7_  &  (~ i_6_)  &  n_n5  &  n_n8 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n5  &  n_n8 ) ;
 assign wire3797 = ( wire3796 ) | ( n_n5  &  n_n14  &  wire72 ) ;
 assign wire3798 = ( wire271 ) | ( n_n4  &  n_n13  &  n_n17 ) ;
 assign wire3800 = ( n_n5  &  n_n10  &  n_n15 ) | ( n_n5  &  n_n15  &  n_n12 ) ;
 assign wire3801 = ( o_28_ ) | ( wire78 ) | ( n_n1166 ) | ( wire3800 ) ;
 assign wire3802 = ( (~ i_7_)  &  i_6_  &  n_n7  &  n_n3 ) | ( i_7_  &  (~ i_6_)  &  n_n7  &  n_n3 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n7  &  n_n3 ) ;
 assign wire3804 = ( o_21_ ) | ( n_n953 ) | ( n_n1203 ) | ( n_n1056 ) ;
 assign wire3806 = ( n_n3  &  n_n12  &  n_n16 ) | ( n_n1  &  n_n12  &  n_n16 ) ;
 assign wire3807 = ( i_7_  &  (~ i_6_)  &  n_n2  &  n_n11 ) | ( (~ i_7_)  &  (~ i_6_)  &  n_n2  &  n_n11 ) ;
 assign wire3808 = ( n_n13  &  n_n3  &  n_n15 ) | ( n_n3  &  n_n15  &  n_n9 ) ;
 assign wire3809 = ( n_n1135 ) | ( n_n1137 ) | ( n_n3  &  wire71 ) ;
 assign wire3810 = ( wire127 ) | ( wire247 ) ;
 assign wire3813 = ( n_n1076 ) | ( wire3465 ) | ( n_n3  &  wire69 ) ;
 assign wire3816 = ( wire260 ) | ( wire3806 ) | ( wire3807 ) | ( wire3808 ) ;
 assign wire3818 = ( wire297 ) | ( n_n1147 ) | ( wire532 ) | ( wire3279 ) ;
 assign wire3820 = ( wire107 ) | ( wire217 ) | ( wire3809 ) | ( wire3810 ) ;
 assign wire3821 = ( wire250 ) | ( n_n923 ) | ( wire3621 ) | ( wire3816 ) ;
 assign wire3822 = ( wire156 ) | ( wire270 ) | ( wire3797 ) | ( wire3798 ) ;
 assign wire3823 = ( wire283 ) | ( n_n859 ) | ( wire3359 ) | ( wire3801 ) ;
 assign wire3827 = ( wire196 ) | ( wire323 ) | ( wire3277 ) | ( wire3296 ) ;
 assign wire3829 = ( wire327 ) | ( n_n711 ) | ( wire231 ) | ( wire3823 ) ;
 assign wire3830 = ( n_n660 ) | ( wire295 ) | ( wire3813 ) | ( wire3818 ) ;
 assign wire3831 = ( n_n427 ) | ( wire347 ) | ( wire3820 ) ;
 assign wire3832 = ( wire3821 ) | ( wire3822 ) | ( wire3827 ) ;
 assign wire3841 = ( wire158 ) | ( n_n825 ) | ( wire134 ) | ( wire78 ) ;
 assign wire3842 = ( o_8_ ) | ( wire346 ) | ( wire133 ) | ( wire140 ) ;
 assign wire3843 = ( wire187 ) | ( wire235 ) | ( wire308 ) | ( wire316 ) ;
 assign wire3844 = ( wire94 ) | ( n_n872 ) | ( wire191 ) | ( wire3841 ) ;
 assign wire3847 = ( wire152 ) | ( n_n673 ) | ( wire302 ) | ( wire3842 ) ;
 assign wire3850 = ( n_n1243 ) | ( n_n0  &  wire71 ) ;
 assign wire3853 = ( wire109 ) | ( wire293 ) ;
 assign wire3854 = ( o_9_ ) | ( n_n1300 ) | ( n_n1301 ) | ( n_n1315 ) ;
 assign wire3855 = ( wire271 ) | ( wire259 ) ;
 assign wire3856 = ( n_n1287 ) | ( n_n814 ) | ( n_n1316 ) | ( wire101 ) ;
 assign wire3857 = ( o_20_ ) | ( wire159 ) | ( wire135 ) | ( wire219 ) ;
 assign wire3860 = ( wire183 ) | ( n_n813 ) | ( wire207 ) ;
 assign wire3864 = ( n_n744 ) | ( wire184 ) | ( n_n805 ) | ( wire104 ) ;
 assign wire3868 = ( wire287 ) | ( wire305 ) ;
 assign wire3870 = ( n_n803 ) | ( wire97 ) | ( n_n3  &  wire71 ) ;
 assign wire3871 = ( n_n935 ) | ( wire77 ) | ( n_n1213 ) | ( wire3857 ) ;
 assign wire3872 = ( n_n1197 ) | ( wire88 ) | ( wire253 ) | ( wire3860 ) ;
 assign wire3873 = ( wire107 ) | ( n_n581 ) | ( n_n742 ) | ( n_n1034 ) ;
 assign wire3874 = ( n_n824 ) | ( wire3850 ) | ( wire3864 ) ;
 assign wire3875 = ( wire3853 ) | ( wire3854 ) | ( wire3855 ) | ( wire3856 ) ;
 assign wire3876 = ( n_n845 ) | ( wire95 ) | ( wire320 ) | ( wire3467 ) ;
 assign wire3877 = ( wire250 ) | ( n_n711 ) | ( wire3621 ) | ( wire3868 ) ;
 assign wire3882 = ( wire3870 ) | ( wire3871 ) | ( wire3877 ) ;
 assign wire3883 = ( wire3872 ) | ( wire3873 ) | ( wire3874 ) | ( wire3875 ) ;
 assign wire3885 = ( wire3843 ) | ( wire3844 ) | ( wire3847 ) | ( wire3883 ) ;
 assign wire3886 = ( n_n1009 ) | ( n_n19  &  n_n8  &  n_n15 ) ;
 assign wire3890 = ( wire93 ) | ( n_n1155 ) | ( wire160 ) ;
 assign wire3892 = ( wire222 ) | ( wire297 ) | ( wire3279 ) | ( wire3890 ) ;
 assign wire3897 = ( n_n1169 ) | ( n_n1314 ) | ( n_n1165 ) | ( n_n821 ) ;
 assign wire3899 = ( n_n1180 ) | ( wire271 ) | ( n_n817 ) ;
 assign wire3900 = ( wire162 ) | ( wire291 ) | ( n_n961 ) | ( wire500 ) ;
 assign wire3903 = ( wire99 ) | ( n_n1322 ) | ( wire207 ) | ( wire3899 ) ;
 assign wire3905 = ( wire114 ) | ( n_n814 ) | ( wire97 ) | ( wire3897 ) ;
 assign wire3908 = ( wire129 ) | ( wire107 ) | ( n_n989 ) | ( wire3900 ) ;
 assign wire3909 = ( wire154 ) | ( wire139 ) | ( wire3903 ) | ( wire3905 ) ;
 assign wire3910 = ( n_n573 ) | ( wire238 ) | ( n_n574 ) | ( wire3360 ) ;
 assign wire3911 = ( wire319 ) | ( n_n1006 ) | ( n_n563 ) | ( wire3892 ) ;
 assign wire3915 = ( o_10_ ) | ( n_n3  &  n_n12  &  n_n16 ) ;
 assign wire3916 = ( o_27_ ) | ( n_n1215 ) | ( wire277 ) ;
 assign wire3920 = ( wire261 ) | ( wire217 ) | ( wire3915 ) | ( wire3916 ) ;
 assign wire3921 = ( n_n459 ) | ( wire129 ) | ( wire107 ) ;
 assign wire3922 = ( n_n895 ) | ( wire283 ) | ( n_n911 ) | ( wire3441 ) ;
 assign wire3925 = ( wire200 ) | ( wire201 ) | ( wire3439 ) | ( wire3440 ) ;
 assign wire3926 = ( n_n573 ) | ( wire340 ) | ( wire3920 ) ;
 assign wire3928 = ( wire285 ) | ( wire284 ) | ( wire3749 ) | ( wire3926 ) ;
 assign wire3929 = ( n_n10  &  n_n1 ) | ( n_n17  &  n_n12 ) ;
 assign wire3935 = ( n_n1135 ) | ( n_n1134 ) | ( n_n1137 ) | ( n_n1136 ) ;
 assign wire3936 = ( wire104 ) | ( n_n1083 ) ;
 assign wire3937 = ( n_n926 ) | ( n_n1238 ) | ( n_n1239 ) ;
 assign wire3938 = ( wire113 ) | ( n_n930 ) ;
 assign wire3939 = ( wire161 ) | ( wire158 ) ;
 assign wire3940 = ( o_9_ ) | ( o_8_ ) | ( n_n1302 ) | ( n_n872 ) ;
 assign wire3941 = ( n_n953 ) | ( n_n1288 ) | ( n_n1322 ) | ( n_n1139 ) ;
 assign wire3942 = ( n_n1203 ) | ( n_n1138 ) | ( wire273 ) | ( wire3929 ) ;
 assign wire3944 = ( wire354 ) | ( n_n1226 ) | ( wire77 ) | ( wire160 ) ;
 assign wire3945 = ( n_n1021 ) | ( n_n553 ) ;
 assign wire3950 = ( wire346 ) | ( wire3941 ) ;
 assign wire3951 = ( n_n963 ) | ( wire76 ) | ( n_n1017 ) | ( n_n859 ) ;
 assign wire3952 = ( o_18_ ) | ( wire130 ) | ( wire156 ) ;
 assign wire3955 = ( n_n923 ) | ( wire217 ) | ( wire3942 ) ;
 assign wire3957 = ( wire148 ) | ( wire198 ) | ( wire3935 ) | ( wire3936 ) ;
 assign wire3958 = ( wire3937 ) | ( wire3938 ) | ( wire3939 ) | ( wire3940 ) ;
 assign wire3962 = ( n_n387 ) | ( n_n711 ) | ( wire295 ) | ( wire194 ) ;
 assign wire3965 = ( n_n534 ) | ( n_n895 ) | ( wire173 ) | ( wire3222 ) ;
 assign wire3966 = ( wire252 ) | ( wire331 ) | ( n_n563 ) | ( n_n931 ) ;
 assign wire3967 = ( wire342 ) | ( wire3950 ) | ( wire3951 ) | ( wire3952 ) ;
 assign wire3968 = ( wire3944 ) | ( wire3945 ) | ( wire3955 ) | ( wire3962 ) ;
 assign wire3969 = ( wire3957 ) | ( wire3958 ) | ( wire3965 ) ;
 assign wire3973 = ( n_n1268 ) | ( n_n1272 ) | ( wire132 ) ;
 assign wire3975 = ( wire112 ) | ( wire209 ) | ( n_n802 ) | ( n_n1223 ) ;
 assign wire3976 = ( n_n1245 ) | ( n_n1244 ) | ( wire277 ) | ( wire3975 ) ;
 assign wire3978 = ( wire177 ) | ( wire238 ) | ( wire3641 ) | ( wire3976 ) ;
 assign wire3982 = ( o_9_ ) | ( n_n1302 ) | ( n_n553 ) ;
 assign wire3983 = ( n_n1010 ) | ( n_n1021 ) | ( wire265 ) ;
 assign wire3985 = ( wire76 ) | ( n_n1017 ) | ( wire3982 ) | ( wire3983 ) ;
 assign wire3986 = ( wire150 ) | ( wire148 ) | ( wire3430 ) | ( wire3985 ) ;
 assign wire3993 = ( wire183 ) | ( n_n0  &  wire69 ) ;
 assign wire3994 = ( n_n1300 ) | ( wire266 ) | ( n_n1315 ) ;
 assign wire3995 = ( o_7_ ) | ( n_n1147 ) | ( n_n1238 ) | ( n_n1155 ) ;
 assign wire3997 = ( n_n1009 ) | ( n_n1256 ) | ( wire127 ) | ( wire471 ) ;
 assign wire3998 = ( wire147 ) | ( wire184 ) | ( wire545 ) | ( wire546 ) ;
 assign wire4001 = ( n_n1049 ) | ( n_n1021 ) | ( wire77 ) | ( n_n1020 ) ;
 assign wire4003 = ( n_n1083 ) | ( n_n468 ) | ( wire236 ) | ( wire473 ) ;
 assign wire4004 = ( n_n1022 ) | ( n_n1253 ) | ( n_n1231 ) | ( wire3997 ) ;
 assign wire4005 = ( wire3993 ) | ( wire3994 ) | ( wire3998 ) ;
 assign wire4006 = ( wire229 ) | ( n_n642 ) | ( wire270 ) | ( wire3797 ) ;
 assign wire4007 = ( wire156 ) | ( n_n859 ) | ( wire3798 ) | ( wire3801 ) ;
 assign wire4008 = ( wire323 ) | ( wire140 ) | ( wire3579 ) | ( wire3995 ) ;
 assign wire4009 = ( wire297 ) | ( n_n738 ) | ( wire3279 ) | ( wire4001 ) ;
 assign wire4013 = ( wire4009 ) | ( wire4008 ) ;
 assign wire4014 = ( wire3716 ) | ( wire3717 ) | ( wire4003 ) | ( wire4004 ) ;
 assign wire4015 = ( wire347 ) | ( wire321 ) ;
 assign wire4016 = ( n_n1006 ) | ( wire4005 ) | ( wire4006 ) | ( wire4007 ) ;
 assign wire4019 = ( n_n1017 ) | ( n_n1024 ) | ( n_n1025 ) ;
 assign wire4020 = ( n_n1022 ) | ( n_n1298 ) | ( wire3218 ) | ( wire4019 ) ;
 assign wire4023 = ( n_n744 ) | ( n_n906 ) | ( n_n745 ) | ( wire268 ) ;
 assign wire4024 = ( wire325 ) | ( n_n858 ) | ( wire3462 ) ;
 assign wire4025 = ( wire298 ) | ( wire110 ) | ( wire303 ) | ( wire4023 ) ;
 assign wire4027 = ( wire177 ) | ( wire154 ) | ( wire197 ) | ( wire4024 ) ;
 assign wire4029 = ( wire115 ) | ( wire165 ) | ( wire4020 ) | ( wire4025 ) ;
 assign wire4031 = ( wire267 ) | ( wire322 ) | ( wire4027 ) | ( wire4029 ) ;
 assign wire4037 = ( o_30_ ) | ( n_n1261 ) | ( n_n756 ) | ( n_n1268 ) ;
 assign wire4038 = ( n_n949 ) | ( wire162 ) | ( wire243 ) ;
 assign wire4039 = ( n_n950 ) | ( wire159 ) | ( wire219 ) ;
 assign wire4042 = ( n_n616 ) | ( n_n617 ) | ( n_n1083 ) | ( wire127 ) ;
 assign wire4044 = ( wire104 ) | ( wire257 ) | ( n_n1226 ) | ( wire77 ) ;
 assign wire4046 = ( wire99 ) | ( wire235 ) | ( n_n948 ) | ( wire173 ) ;
 assign wire4047 = ( wire161 ) | ( wire135 ) | ( wire4037 ) | ( wire4042 ) ;
 assign wire4050 = ( n_n1121 ) | ( wire325 ) | ( wire140 ) | ( wire3274 ) ;
 assign wire4051 = ( wire4038 ) | ( wire4039 ) | ( wire4044 ) ;
 assign wire4053 = ( wire301 ) | ( wire197 ) | ( wire270 ) | ( n_n823 ) ;
 assign wire4055 = ( n_n673 ) | ( wire225 ) | ( wire3713 ) | ( wire4050 ) ;
 assign wire4056 = ( wire4046 ) | ( wire4047 ) | ( wire4051 ) ;
 assign wire4057 = ( n_n845 ) | ( wire332 ) | ( wire315 ) | ( n_n858 ) ;
 assign wire4058 = ( wire115 ) | ( wire192 ) | ( wire255 ) | ( wire4053 ) ;
 assign wire4063 = ( n_n1321 ) | ( wire147 ) | ( wire265 ) | ( wire281 ) ;
 assign wire4065 = ( wire110 ) | ( n_n1010 ) | ( n_n1320 ) | ( wire4063 ) ;
 assign wire4066 = ( wire76 ) | ( n_n1017 ) | ( wire85 ) | ( wire231 ) ;
 assign wire4068 = ( wire3750 ) | ( wire3751 ) | ( wire4066 ) ;
 assign wire4069 = ( n_n990 ) | ( wire233 ) | ( n_n1014 ) | ( wire4065 ) ;
 assign wire4071 = ( n_n10 ) | ( n_n7  &  n_n6  &  n_n14 ) ;
 assign wire4074 = ( wire88 ) | ( n_n5  &  wire72 ) ;
 assign wire4076 = ( n_n1163 ) | ( n_n1282 ) | ( wire4071 ) ;
 assign wire4079 = ( wire208 ) | ( n_n1167 ) | ( wire269 ) ;
 assign wire4081 = ( n_n1203 ) | ( wire273 ) | ( wire3210 ) | ( wire4076 ) ;
 assign wire4082 = ( wire306 ) | ( wire237 ) ;
 assign wire4083 = ( wire309 ) | ( wire111 ) | ( n_n960 ) | ( n_n955 ) ;
 assign wire4084 = ( wire130 ) | ( n_n925 ) | ( wire4074 ) | ( wire4079 ) ;
 assign wire4086 = ( wire320 ) | ( wire139 ) | ( wire3393 ) ;
 assign wire4090 = ( n_n95 ) | ( n_n1334 ) | ( wire128 ) | ( wire3296 ) ;
 assign wire4091 = ( wire331 ) | ( wire179 ) | ( n_n931 ) | ( wire4086 ) ;
 assign wire4092 = ( n_n901 ) | ( wire4081 ) | ( wire4082 ) | ( wire4083 ) ;
 assign wire4093 = ( wire343 ) | ( wire211 ) | ( wire3432 ) | ( wire3607 ) ;
 assign wire4094 = ( n_n427 ) | ( wire4084 ) | ( wire4090 ) ;
 assign wire4097 = ( wire4091 ) | ( wire4092 ) | ( wire4094 ) ;
 assign wire4098 = ( wire76 ) | ( n_n1010 ) | ( n_n1320 ) ;
 assign wire4099 = ( n_n1321 ) | ( wire95 ) | ( wire265 ) | ( wire3467 ) ;
 assign wire4100 = ( n_n1049 ) | ( wire77 ) | ( wire4098 ) ;
 assign wire4101 = ( wire156 ) | ( wire270 ) | ( wire3797 ) | ( wire3798 ) ;
 assign wire4105 = ( wire83 ) | ( wire85 ) | ( wire4020 ) | ( wire4101 ) ;
 assign wire4106 = ( wire333 ) | ( n_n859 ) | ( wire3801 ) | ( wire4099 ) ;
 assign wire4108 = ( wire108 ) | ( wire337 ) | ( wire264 ) | ( wire3892 ) ;
 assign wire4109 = ( wire193 ) | ( wire165 ) | ( n_n989 ) | ( wire4100 ) ;
 assign wire4112 = ( wire4105 ) | ( wire4106 ) | ( wire4109 ) ;
 assign wire4113 = ( n_n0 ) | ( n_n17  &  n_n1  &  n_n8 ) ;
 assign wire4115 = ( wire162 ) | ( n_n582 ) | ( wire4113 ) ;
 assign wire4117 = ( wire129 ) | ( wire107 ) | ( wire139 ) | ( wire4115 ) ;
 assign wire4119 = ( n_n4  &  n_n12  &  n_n16 ) | ( n_n2  &  n_n12  &  n_n16 ) ;
 assign wire4122 = ( n_n0  &  n_n8  &  n_n16 ) | ( n_n3  &  n_n8  &  n_n16 ) ;
 assign wire4123 = ( n_n5  &  n_n12  &  n_n16 ) | ( n_n19  &  n_n12  &  n_n16 ) ;
 assign wire4125 = ( n_n5  &  n_n8  &  n_n16 ) | ( n_n4  &  n_n8  &  n_n16 ) ;
 assign wire4126 = ( n_n1300 ) | ( n_n1315 ) | ( wire4119 ) ;
 assign wire4127 = ( n_n1269 ) | ( n_n1224 ) | ( n_n1284 ) | ( n_n1148 ) ;
 assign wire4128 = ( wire4123 ) | ( wire4122 ) ;
 assign wire4129 = ( n_n1119 ) | ( n_n1133 ) | ( wire4125 ) ;
 assign wire4138 = ( n_n1135 ) | ( n_n826 ) | ( n_n1137 ) ;
 assign wire4139 = ( n_n1024 ) | ( n_n10  &  n_n1  &  wire67 ) ;
 assign wire4140 = ( o_11_ ) | ( n_n1302 ) | ( n_n1163 ) | ( n_n1256 ) ;
 assign wire4141 = ( n_n1258 ) | ( n_n1138 ) | ( n_n1167 ) | ( n_n1303 ) ;
 assign wire4142 = ( n_n1170 ) | ( n_n1273 ) | ( n_n1301 ) | ( n_n1077 ) ;
 assign wire4144 = ( n_n1076 ) | ( n_n910 ) | ( n_n909 ) ;
 assign wire4145 = ( n_n1274 ) | ( wire281 ) | ( n_n1298 ) | ( wire3218 ) ;
 assign wire4149 = ( n_n911 ) | ( n_n797 ) | ( wire3363 ) | ( wire3441 ) ;
 assign wire4150 = ( wire226 ) | ( wire309 ) | ( wire4144 ) ;
 assign wire4151 = ( wire147 ) | ( wire300 ) | ( wire4138 ) | ( wire4145 ) ;
 assign wire4152 = ( wire4139 ) | ( wire4140 ) | ( wire4141 ) | ( wire4142 ) ;
 assign wire4153 = ( n_n459 ) | ( wire216 ) | ( wire3304 ) | ( wire3305 ) ;
 assign wire4154 = ( n_n800 ) | ( wire195 ) | ( wire231 ) | ( wire3361 ) ;
 assign wire4160 = ( wire323 ) | ( n_n786 ) | ( wire4154 ) ;
 assign wire4161 = ( wire4149 ) | ( wire4150 ) | ( wire4151 ) | ( wire4152 ) ;
 assign wire4162 = ( wire218 ) | ( wire189 ) | ( wire238 ) | ( wire315 ) ;
 assign wire4163 = ( wire326 ) | ( wire193 ) | ( n_n989 ) | ( wire4153 ) ;
 assign wire4166 = ( n_n4  &  n_n11  &  n_n16 ) | ( n_n11  &  n_n1  &  n_n16 ) ;
 assign wire4167 = ( n_n5  &  n_n11  &  n_n16 ) | ( n_n2  &  n_n11  &  n_n16 ) ;
 assign wire4168 = ( n_n6  &  n_n11  &  n_n16 ) | ( n_n11  &  n_n3  &  n_n16 ) ;
 assign wire4169 = ( n_n0  &  n_n11  &  n_n16 ) | ( n_n11  &  n_n19  &  n_n16 ) ;


endmodule

